magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -66 377 2370 897
<< pwell >>
rect 1865 217 2298 283
rect 8 43 2298 217
rect -26 -43 2330 43
<< mvnmos >>
rect 91 107 191 191
rect 247 107 347 191
rect 389 107 489 191
rect 545 107 645 191
rect 687 107 787 191
rect 844 107 944 191
rect 1114 107 1214 191
rect 1380 107 1480 191
rect 1536 107 1636 191
rect 1678 107 1778 191
rect 1944 173 2044 257
rect 2119 107 2219 257
<< mvpmos >>
rect 87 587 187 671
rect 262 587 362 737
rect 404 587 504 737
rect 560 587 660 737
rect 702 587 802 737
rect 858 587 958 737
rect 1154 525 1254 675
rect 1445 593 1545 743
rect 1624 593 1724 677
rect 1766 593 1866 677
rect 1938 443 2038 527
rect 2117 443 2217 743
<< mvndiff >>
rect 1891 232 1944 257
rect 1891 198 1899 232
rect 1933 198 1944 232
rect 34 166 91 191
rect 34 132 46 166
rect 80 132 91 166
rect 34 107 91 132
rect 191 166 247 191
rect 191 132 202 166
rect 236 132 247 166
rect 191 107 247 132
rect 347 107 389 191
rect 489 166 545 191
rect 489 132 500 166
rect 534 132 545 166
rect 489 107 545 132
rect 645 107 687 191
rect 787 166 844 191
rect 787 132 798 166
rect 832 132 844 166
rect 787 107 844 132
rect 944 166 997 191
rect 944 132 955 166
rect 989 132 997 166
rect 944 107 997 132
rect 1057 166 1114 191
rect 1057 132 1069 166
rect 1103 132 1114 166
rect 1057 107 1114 132
rect 1214 166 1267 191
rect 1214 132 1225 166
rect 1259 132 1267 166
rect 1214 107 1267 132
rect 1327 168 1380 191
rect 1327 134 1335 168
rect 1369 134 1380 168
rect 1327 107 1380 134
rect 1480 166 1536 191
rect 1480 132 1491 166
rect 1525 132 1536 166
rect 1480 107 1536 132
rect 1636 107 1678 191
rect 1778 166 1831 191
rect 1891 173 1944 198
rect 2044 245 2119 257
rect 2044 211 2074 245
rect 2108 211 2119 245
rect 2044 173 2119 211
rect 1778 132 1789 166
rect 1823 132 1831 166
rect 2066 153 2119 173
rect 1778 107 1831 132
rect 2066 119 2074 153
rect 2108 119 2119 153
rect 2066 107 2119 119
rect 2219 245 2272 257
rect 2219 211 2230 245
rect 2264 211 2272 245
rect 2219 153 2272 211
rect 2219 119 2230 153
rect 2264 119 2272 153
rect 2219 107 2272 119
<< mvpdiff >>
rect 209 725 262 737
rect 209 691 217 725
rect 251 691 262 725
rect 209 671 262 691
rect 30 646 87 671
rect 30 612 42 646
rect 76 612 87 646
rect 30 587 87 612
rect 187 633 262 671
rect 187 599 217 633
rect 251 599 262 633
rect 187 587 262 599
rect 362 587 404 737
rect 504 729 560 737
rect 504 695 515 729
rect 549 695 560 729
rect 504 629 560 695
rect 504 595 515 629
rect 549 595 560 629
rect 504 587 560 595
rect 660 587 702 737
rect 802 729 858 737
rect 802 695 813 729
rect 847 695 858 729
rect 802 639 858 695
rect 802 605 813 639
rect 847 605 858 639
rect 802 587 858 605
rect 958 652 1015 737
rect 1388 735 1445 743
rect 1388 701 1400 735
rect 1434 701 1445 735
rect 958 618 969 652
rect 1003 618 1015 652
rect 958 587 1015 618
rect 1097 667 1154 675
rect 1097 633 1109 667
rect 1143 633 1154 667
rect 1097 567 1154 633
rect 1097 533 1109 567
rect 1143 533 1154 567
rect 1097 525 1154 533
rect 1254 667 1311 675
rect 1254 633 1265 667
rect 1299 633 1311 667
rect 1254 567 1311 633
rect 1388 635 1445 701
rect 1388 601 1400 635
rect 1434 601 1445 635
rect 1388 593 1445 601
rect 1545 735 1602 743
rect 1545 701 1556 735
rect 1590 701 1602 735
rect 2060 735 2117 743
rect 1545 677 1602 701
rect 2060 701 2072 735
rect 2106 701 2117 735
rect 1545 635 1624 677
rect 1545 601 1556 635
rect 1590 601 1624 635
rect 1545 593 1624 601
rect 1724 593 1766 677
rect 1866 652 1923 677
rect 1866 618 1877 652
rect 1911 618 1923 652
rect 1866 593 1923 618
rect 2060 638 2117 701
rect 2060 604 2072 638
rect 2106 604 2117 638
rect 1254 533 1265 567
rect 1299 533 1311 567
rect 1254 525 1311 533
rect 2060 541 2117 604
rect 2060 527 2072 541
rect 1881 502 1938 527
rect 1881 468 1893 502
rect 1927 468 1938 502
rect 1881 443 1938 468
rect 2038 507 2072 527
rect 2106 507 2117 541
rect 2038 443 2117 507
rect 2217 735 2274 743
rect 2217 701 2228 735
rect 2262 701 2274 735
rect 2217 652 2274 701
rect 2217 618 2228 652
rect 2262 618 2274 652
rect 2217 568 2274 618
rect 2217 534 2228 568
rect 2262 534 2274 568
rect 2217 485 2274 534
rect 2217 451 2228 485
rect 2262 451 2274 485
rect 2217 443 2274 451
<< mvndiffc >>
rect 1899 198 1933 232
rect 46 132 80 166
rect 202 132 236 166
rect 500 132 534 166
rect 798 132 832 166
rect 955 132 989 166
rect 1069 132 1103 166
rect 1225 132 1259 166
rect 1335 134 1369 168
rect 1491 132 1525 166
rect 2074 211 2108 245
rect 1789 132 1823 166
rect 2074 119 2108 153
rect 2230 211 2264 245
rect 2230 119 2264 153
<< mvpdiffc >>
rect 217 691 251 725
rect 42 612 76 646
rect 217 599 251 633
rect 515 695 549 729
rect 515 595 549 629
rect 813 695 847 729
rect 813 605 847 639
rect 1400 701 1434 735
rect 969 618 1003 652
rect 1109 633 1143 667
rect 1109 533 1143 567
rect 1265 633 1299 667
rect 1400 601 1434 635
rect 1556 701 1590 735
rect 2072 701 2106 735
rect 1556 601 1590 635
rect 1877 618 1911 652
rect 2072 604 2106 638
rect 1265 533 1299 567
rect 1893 468 1927 502
rect 2072 507 2106 541
rect 2228 701 2262 735
rect 2228 618 2262 652
rect 2228 534 2262 568
rect 2228 451 2262 485
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2304 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2304 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
<< poly >>
rect 262 737 362 763
rect 404 737 504 763
rect 560 737 660 763
rect 702 737 802 763
rect 858 737 958 763
rect 1445 743 1545 769
rect 2117 743 2217 769
rect 87 671 187 697
rect 1154 675 1254 701
rect 87 565 187 587
rect 262 565 362 587
rect 87 539 362 565
rect 87 505 133 539
rect 167 505 251 539
rect 285 505 362 539
rect 87 499 362 505
rect 404 539 504 587
rect 404 505 424 539
rect 458 505 504 539
rect 87 485 305 499
rect 87 471 187 485
rect 87 437 133 471
rect 167 437 187 471
rect 404 471 504 505
rect 404 457 424 471
rect 347 443 424 457
rect 87 317 187 437
rect 247 437 424 443
rect 458 437 504 471
rect 247 391 504 437
rect 560 499 660 587
rect 560 465 606 499
rect 640 465 660 499
rect 560 431 660 465
rect 560 397 606 431
rect 640 397 660 431
rect 87 217 191 317
rect 91 191 191 217
rect 247 191 347 391
rect 560 381 660 397
rect 702 491 802 587
rect 858 565 958 587
rect 702 457 722 491
rect 756 457 802 491
rect 702 423 802 457
rect 702 389 722 423
rect 756 389 802 423
rect 702 355 802 389
rect 389 331 489 349
rect 389 297 409 331
rect 443 297 489 331
rect 389 263 489 297
rect 389 229 409 263
rect 443 229 489 263
rect 389 191 489 229
rect 531 323 645 339
rect 531 289 547 323
rect 581 289 645 323
rect 702 321 722 355
rect 756 321 802 355
rect 702 317 802 321
rect 531 217 645 289
rect 545 191 645 217
rect 687 217 802 317
rect 844 483 958 565
rect 1624 677 1724 703
rect 1766 677 1866 703
rect 1154 503 1254 525
rect 1445 503 1545 593
rect 1624 505 1724 593
rect 844 449 887 483
rect 921 449 958 483
rect 844 415 958 449
rect 844 381 887 415
rect 921 381 958 415
rect 844 347 958 381
rect 844 313 887 347
rect 921 313 958 347
rect 844 279 958 313
rect 844 245 887 279
rect 921 245 958 279
rect 844 217 958 245
rect 1114 463 1545 503
rect 1644 493 1724 505
rect 1114 403 1602 463
rect 1644 459 1664 493
rect 1698 459 1724 493
rect 1644 439 1724 459
rect 1114 353 1214 403
rect 1445 397 1602 403
rect 1522 391 1622 397
rect 1114 319 1134 353
rect 1168 319 1214 353
rect 1114 285 1214 319
rect 1114 251 1134 285
rect 1168 251 1214 285
rect 687 191 787 217
rect 844 191 944 217
rect 1114 191 1214 251
rect 1380 335 1480 355
rect 1380 301 1421 335
rect 1455 301 1480 335
rect 1380 267 1480 301
rect 1522 291 1636 391
rect 1766 351 1866 593
rect 1938 527 2038 553
rect 1380 233 1421 267
rect 1455 233 1480 267
rect 1380 191 1480 233
rect 1536 191 1636 291
rect 1678 331 1866 351
rect 1678 297 1724 331
rect 1758 297 1866 331
rect 1678 263 1866 297
rect 1938 417 2038 443
rect 2117 417 2217 443
rect 1938 393 2219 417
rect 1938 359 1990 393
rect 2024 359 2219 393
rect 1938 283 2219 359
rect 1678 229 1724 263
rect 1758 229 1866 263
rect 1944 257 2044 283
rect 2119 257 2219 283
rect 1678 213 1866 229
rect 1678 191 1778 213
rect 1944 147 2044 173
rect 91 81 191 107
rect 247 81 347 107
rect 389 81 489 107
rect 545 81 645 107
rect 687 81 787 107
rect 844 81 944 107
rect 1114 81 1214 107
rect 1380 81 1480 107
rect 1536 81 1636 107
rect 1678 81 1778 107
rect 2119 81 2219 107
<< polycont >>
rect 133 505 167 539
rect 251 505 285 539
rect 424 505 458 539
rect 133 437 167 471
rect 424 437 458 471
rect 606 465 640 499
rect 606 397 640 431
rect 722 457 756 491
rect 722 389 756 423
rect 409 297 443 331
rect 409 229 443 263
rect 547 289 581 323
rect 722 321 756 355
rect 887 449 921 483
rect 887 381 921 415
rect 887 313 921 347
rect 887 245 921 279
rect 1664 459 1698 493
rect 1134 319 1168 353
rect 1134 251 1168 285
rect 1421 301 1455 335
rect 1421 233 1455 267
rect 1724 297 1758 331
rect 1990 359 2024 393
rect 1724 229 1758 263
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2304 831
rect 112 735 302 741
rect 112 701 118 735
rect 152 701 190 735
rect 224 725 262 735
rect 251 701 262 725
rect 296 701 302 735
rect 112 691 217 701
rect 251 691 302 701
rect 26 646 76 679
rect 26 612 42 646
rect 26 269 76 612
rect 112 633 302 691
rect 515 729 565 745
rect 549 695 565 729
rect 112 599 217 633
rect 251 599 302 633
rect 117 539 359 555
rect 117 505 133 539
rect 167 505 251 539
rect 285 505 359 539
rect 117 471 359 505
rect 117 437 133 471
rect 167 437 359 471
rect 408 539 474 652
rect 408 505 424 539
rect 458 505 474 539
rect 515 629 565 695
rect 549 595 565 629
rect 673 735 863 745
rect 673 701 679 735
rect 713 701 751 735
rect 785 729 823 735
rect 785 701 813 729
rect 857 701 863 735
rect 673 695 813 701
rect 847 695 863 701
rect 673 639 863 695
rect 673 605 813 639
rect 847 605 863 639
rect 899 727 1073 761
rect 515 569 565 595
rect 899 569 933 727
rect 515 535 933 569
rect 969 652 1003 691
rect 408 471 474 505
rect 408 437 424 471
rect 458 437 474 471
rect 590 465 606 499
rect 640 465 667 499
rect 117 401 359 437
rect 590 431 667 465
rect 117 367 554 401
rect 590 397 606 431
rect 640 397 667 431
rect 590 381 667 397
rect 520 339 554 367
rect 393 297 409 331
rect 443 297 459 331
rect 393 269 459 297
rect 520 323 597 339
rect 520 289 547 323
rect 581 289 597 323
rect 26 263 459 269
rect 26 235 409 263
rect 26 166 96 235
rect 393 229 409 235
rect 443 253 459 263
rect 633 253 667 381
rect 703 491 772 499
rect 703 457 722 491
rect 756 457 772 491
rect 703 423 772 457
rect 703 389 722 423
rect 756 389 772 423
rect 703 355 772 389
rect 703 321 722 355
rect 756 321 772 355
rect 703 305 772 321
rect 806 269 840 535
rect 443 229 667 253
rect 393 219 667 229
rect 703 235 840 269
rect 874 483 933 499
rect 874 449 887 483
rect 921 449 933 483
rect 874 415 933 449
rect 874 381 887 415
rect 921 381 933 415
rect 874 347 933 381
rect 874 313 887 347
rect 921 313 933 347
rect 874 279 933 313
rect 874 245 887 279
rect 921 245 933 279
rect 26 132 46 166
rect 80 132 96 166
rect 26 99 96 132
rect 132 166 322 199
rect 703 183 737 235
rect 874 229 933 245
rect 969 269 1003 618
rect 1039 481 1073 727
rect 1109 735 1143 741
rect 1109 667 1143 701
rect 1109 567 1143 633
rect 1109 517 1143 533
rect 1179 735 1450 753
rect 1179 719 1400 735
rect 1179 481 1213 719
rect 1351 701 1400 719
rect 1434 701 1450 735
rect 1039 447 1213 481
rect 1249 667 1315 683
rect 1249 633 1265 667
rect 1299 633 1315 667
rect 1249 567 1315 633
rect 1249 533 1265 567
rect 1299 533 1315 567
rect 1249 517 1315 533
rect 1351 635 1450 701
rect 1351 601 1400 635
rect 1434 601 1450 635
rect 1351 585 1450 601
rect 1540 735 1606 751
rect 1540 701 1556 735
rect 1590 701 1606 735
rect 1540 635 1606 701
rect 1540 601 1556 635
rect 1590 601 1606 635
rect 1737 735 1927 741
rect 1737 701 1743 735
rect 1777 701 1815 735
rect 1849 701 1887 735
rect 1921 701 1927 735
rect 1737 652 1927 701
rect 1737 618 1877 652
rect 1911 618 1927 652
rect 1737 601 1927 618
rect 1979 735 2169 751
rect 1979 701 1985 735
rect 2019 701 2057 735
rect 2106 701 2129 735
rect 2163 701 2169 735
rect 1979 638 2169 701
rect 1979 604 2072 638
rect 2106 604 2169 638
rect 1540 585 1606 601
rect 1118 353 1184 369
rect 1118 319 1134 353
rect 1168 319 1184 353
rect 1118 285 1184 319
rect 1118 269 1134 285
rect 969 251 1134 269
rect 1168 251 1184 285
rect 969 235 1184 251
rect 969 195 1003 235
rect 132 132 202 166
rect 236 132 322 166
rect 132 113 322 132
rect 132 79 138 113
rect 172 79 210 113
rect 244 79 282 113
rect 316 79 322 113
rect 484 166 737 183
rect 484 132 500 166
rect 534 149 737 166
rect 773 166 891 195
rect 534 132 550 149
rect 484 99 550 132
rect 773 132 798 166
rect 832 132 891 166
rect 773 113 891 132
rect 132 73 322 79
rect 773 79 779 113
rect 813 79 851 113
rect 885 79 891 113
rect 939 166 1005 195
rect 939 132 955 166
rect 989 132 1005 166
rect 939 103 1005 132
rect 1041 166 1159 199
rect 1249 195 1283 517
rect 1351 195 1385 585
rect 1572 565 1606 585
rect 1572 531 1784 565
rect 1979 541 2169 604
rect 1568 493 1714 495
rect 1568 459 1664 493
rect 1698 459 1714 493
rect 1568 443 1714 459
rect 1568 351 1602 443
rect 1750 401 1784 531
rect 1877 502 1943 535
rect 1979 507 2072 541
rect 2106 507 2169 541
rect 2212 735 2280 751
rect 2212 701 2228 735
rect 2262 701 2280 735
rect 2212 652 2280 701
rect 2212 618 2228 652
rect 2262 618 2280 652
rect 2212 568 2280 618
rect 2212 534 2228 568
rect 2262 534 2280 568
rect 1877 468 1893 502
rect 1927 471 1943 502
rect 2212 485 2280 534
rect 1927 468 2110 471
rect 1877 437 2110 468
rect 1041 132 1069 166
rect 1103 132 1159 166
rect 1041 113 1159 132
rect 773 73 891 79
rect 1041 79 1047 113
rect 1081 79 1119 113
rect 1153 79 1159 113
rect 1041 73 1159 79
rect 1209 166 1283 195
rect 1209 132 1225 166
rect 1259 132 1283 166
rect 1209 87 1283 132
rect 1319 168 1385 195
rect 1319 134 1335 168
rect 1369 134 1385 168
rect 1319 123 1385 134
rect 1421 335 1602 351
rect 1455 317 1602 335
rect 1638 393 2040 401
rect 1638 367 1990 393
rect 1421 267 1455 301
rect 1638 249 1672 367
rect 1974 359 1990 367
rect 2024 359 2040 393
rect 1974 351 2040 359
rect 1421 87 1455 233
rect 1491 215 1672 249
rect 1708 297 1724 331
rect 1758 315 1774 331
rect 2076 315 2110 437
rect 1758 297 2110 315
rect 1708 281 2110 297
rect 2212 451 2228 485
rect 2262 451 2280 485
rect 1708 263 1774 281
rect 1708 229 1724 263
rect 1758 229 1774 263
rect 1708 215 1774 229
rect 1883 232 1949 281
rect 2212 245 2280 451
rect 1491 166 1541 215
rect 1883 198 1899 232
rect 1933 198 1949 232
rect 1525 132 1541 166
rect 1491 99 1541 132
rect 1649 166 1839 179
rect 1883 169 1949 198
rect 1985 211 2074 245
rect 2108 211 2175 245
rect 1649 132 1789 166
rect 1823 132 1839 166
rect 1649 113 1839 132
rect 1209 53 1455 87
rect 1649 79 1655 113
rect 1689 79 1727 113
rect 1761 79 1799 113
rect 1833 79 1839 113
rect 1649 73 1839 79
rect 1985 153 2175 211
rect 1985 119 2074 153
rect 2108 119 2175 153
rect 1985 113 2175 119
rect 1985 79 1991 113
rect 2025 79 2063 113
rect 2097 79 2135 113
rect 2169 79 2175 113
rect 2212 211 2230 245
rect 2264 211 2280 245
rect 2212 153 2280 211
rect 2212 119 2230 153
rect 2264 119 2280 153
rect 2212 103 2280 119
rect 1985 73 2175 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2304 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 118 701 152 735
rect 190 725 224 735
rect 190 701 217 725
rect 217 701 224 725
rect 262 701 296 735
rect 679 701 713 735
rect 751 701 785 735
rect 823 729 857 735
rect 823 701 847 729
rect 847 701 857 729
rect 1109 701 1143 735
rect 1743 701 1777 735
rect 1815 701 1849 735
rect 1887 701 1921 735
rect 1985 701 2019 735
rect 2057 701 2072 735
rect 2072 701 2091 735
rect 2129 701 2163 735
rect 138 79 172 113
rect 210 79 244 113
rect 282 79 316 113
rect 779 79 813 113
rect 851 79 885 113
rect 1047 79 1081 113
rect 1119 79 1153 113
rect 1655 79 1689 113
rect 1727 79 1761 113
rect 1799 79 1833 113
rect 1991 79 2025 113
rect 2063 79 2097 113
rect 2135 79 2169 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
<< metal1 >>
rect 0 831 2304 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2304 831
rect 0 791 2304 797
rect 0 735 2304 763
rect 0 701 118 735
rect 152 701 190 735
rect 224 701 262 735
rect 296 701 679 735
rect 713 701 751 735
rect 785 701 823 735
rect 857 701 1109 735
rect 1143 701 1743 735
rect 1777 701 1815 735
rect 1849 701 1887 735
rect 1921 701 1985 735
rect 2019 701 2057 735
rect 2091 701 2129 735
rect 2163 701 2304 735
rect 0 689 2304 701
rect 0 113 2304 125
rect 0 79 138 113
rect 172 79 210 113
rect 244 79 282 113
rect 316 79 779 113
rect 813 79 851 113
rect 885 79 1047 113
rect 1081 79 1119 113
rect 1153 79 1655 113
rect 1689 79 1727 113
rect 1761 79 1799 113
rect 1833 79 1991 113
rect 2025 79 2063 113
rect 2097 79 2135 113
rect 2169 79 2304 113
rect 0 51 2304 79
rect 0 17 2304 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2304 17
rect 0 -23 2304 -17
<< labels >>
rlabel comment s 0 0 0 0 4 sdlxtp_1
flabel metal1 s 0 51 2304 125 0 FreeSans 340 0 0 0 VGND
port 5 nsew ground bidirectional
flabel metal1 s 0 0 2304 23 0 FreeSans 340 0 0 0 VNB
port 6 nsew ground bidirectional
flabel metal1 s 0 689 2304 763 0 FreeSans 340 0 0 0 VPWR
port 8 nsew power bidirectional
flabel metal1 s 0 791 2304 814 0 FreeSans 340 0 0 0 VPB
port 7 nsew power bidirectional
flabel locali s 415 464 449 498 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 415 538 449 572 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 415 612 449 646 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 127 464 161 498 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 223 464 257 498 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 319 464 353 498 0 FreeSans 340 0 0 0 SCE
port 4 nsew signal input
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 703 390 737 424 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 703 464 737 498 0 FreeSans 340 0 0 0 SCD
port 3 nsew signal input
flabel locali s 895 242 929 276 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 895 390 929 424 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 895 464 929 498 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 2239 168 2273 202 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 2239 242 2273 276 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 2239 316 2273 350 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 2239 390 2273 424 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 2239 464 2273 498 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 2239 538 2273 572 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
flabel locali s 2239 612 2273 646 0 FreeSans 340 0 0 0 Q
port 9 nsew signal output
rlabel locali s 773 73 891 195 1 VGND
port 5 nsew ground bidirectional
rlabel locali s 1041 73 1159 199 1 VGND
port 5 nsew ground bidirectional
rlabel locali s 1649 73 1839 179 1 VGND
port 5 nsew ground bidirectional
rlabel locali s 1985 73 2175 245 1 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 51 2304 125 1 VGND
port 5 nsew ground bidirectional
rlabel metal1 s 0 -23 2304 23 1 VNB
port 6 nsew ground bidirectional
rlabel metal1 s 0 791 2304 837 1 VPB
port 7 nsew power bidirectional
rlabel locali s 673 605 863 745 1 VPWR
port 8 nsew power bidirectional
rlabel locali s 1109 517 1143 741 1 VPWR
port 8 nsew power bidirectional
rlabel locali s 1737 601 1927 741 1 VPWR
port 8 nsew power bidirectional
rlabel locali s 1979 507 2169 751 1 VPWR
port 8 nsew power bidirectional
rlabel metal1 s 0 689 2304 763 1 VPWR
port 8 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 2304 814
string GDS_END 719052
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 695106
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
