magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect 24304 8658 24606 9485
rect 23686 5549 24606 8658
rect 211 50 515 4583
rect 1440 4640 10026 4641
rect 1020 4512 10026 4640
rect 1020 1443 13547 4512
rect 1020 1353 10090 1443
rect 23882 2258 24606 5549
rect 23882 1042 24186 2258
rect 14745 976 24186 1042
rect 14745 740 24185 976
<< pwell >>
rect 22740 9368 23626 9398
rect 22740 8719 24185 9368
rect 22740 5489 23626 8719
rect 670 1293 892 4797
rect 22740 4745 23822 5489
rect 23542 2102 23822 4745
rect 13702 1293 23822 2102
rect 670 1102 23822 1293
rect 670 841 14651 1102
<< mvpsubdiff >>
rect 22766 9342 23600 9372
rect 22766 9318 24159 9342
rect 22766 9295 23638 9318
rect 22766 9261 22818 9295
rect 22852 9261 22886 9295
rect 22920 9261 22954 9295
rect 22988 9261 23022 9295
rect 23056 9261 23090 9295
rect 23124 9261 23158 9295
rect 23192 9261 23226 9295
rect 23260 9261 23294 9295
rect 23328 9261 23362 9295
rect 23396 9261 23430 9295
rect 23464 9261 23498 9295
rect 23532 9261 23566 9295
rect 23600 9284 23638 9295
rect 23672 9284 23706 9318
rect 23740 9284 23774 9318
rect 23808 9284 23842 9318
rect 23876 9284 23910 9318
rect 23944 9284 23978 9318
rect 24012 9284 24046 9318
rect 24080 9284 24114 9318
rect 24148 9284 24159 9318
rect 23600 9261 24159 9284
rect 22766 9245 24159 9261
rect 22766 9226 23638 9245
rect 22766 9192 22818 9226
rect 22852 9192 22886 9226
rect 22920 9192 22954 9226
rect 22988 9192 23022 9226
rect 23056 9192 23090 9226
rect 23124 9192 23158 9226
rect 23192 9192 23226 9226
rect 23260 9192 23294 9226
rect 23328 9192 23362 9226
rect 23396 9192 23430 9226
rect 23464 9192 23498 9226
rect 23532 9192 23566 9226
rect 23600 9211 23638 9226
rect 23672 9211 23706 9245
rect 23740 9211 23774 9245
rect 23808 9211 23842 9245
rect 23876 9211 23910 9245
rect 23944 9211 23978 9245
rect 24012 9211 24046 9245
rect 24080 9211 24114 9245
rect 24148 9211 24159 9245
rect 23600 9192 24159 9211
rect 22766 9172 24159 9192
rect 22766 9157 23638 9172
rect 22766 9123 22818 9157
rect 22852 9123 22886 9157
rect 22920 9123 22954 9157
rect 22988 9123 23022 9157
rect 23056 9123 23090 9157
rect 23124 9123 23158 9157
rect 23192 9123 23226 9157
rect 23260 9123 23294 9157
rect 23328 9123 23362 9157
rect 23396 9123 23430 9157
rect 23464 9123 23498 9157
rect 23532 9123 23566 9157
rect 23600 9138 23638 9157
rect 23672 9138 23706 9172
rect 23740 9138 23774 9172
rect 23808 9138 23842 9172
rect 23876 9138 23910 9172
rect 23944 9138 23978 9172
rect 24012 9138 24046 9172
rect 24080 9138 24114 9172
rect 24148 9138 24159 9172
rect 23600 9123 24159 9138
rect 22766 9099 24159 9123
rect 22766 9088 23638 9099
rect 22766 9054 22818 9088
rect 22852 9054 22886 9088
rect 22920 9054 22954 9088
rect 22988 9054 23022 9088
rect 23056 9054 23090 9088
rect 23124 9054 23158 9088
rect 23192 9054 23226 9088
rect 23260 9054 23294 9088
rect 23328 9054 23362 9088
rect 23396 9054 23430 9088
rect 23464 9054 23498 9088
rect 23532 9054 23566 9088
rect 23600 9065 23638 9088
rect 23672 9065 23706 9099
rect 23740 9065 23774 9099
rect 23808 9065 23842 9099
rect 23876 9065 23910 9099
rect 23944 9065 23978 9099
rect 24012 9065 24046 9099
rect 24080 9065 24114 9099
rect 24148 9065 24159 9099
rect 23600 9054 24159 9065
rect 22766 9025 24159 9054
rect 22766 9019 23638 9025
rect 22766 8985 22818 9019
rect 22852 8985 22886 9019
rect 22920 8985 22954 9019
rect 22988 8985 23022 9019
rect 23056 8985 23090 9019
rect 23124 8985 23158 9019
rect 23192 8985 23226 9019
rect 23260 8985 23294 9019
rect 23328 8985 23362 9019
rect 23396 8985 23430 9019
rect 23464 8985 23498 9019
rect 23532 8985 23566 9019
rect 23600 8991 23638 9019
rect 23672 8991 23706 9025
rect 23740 8991 23774 9025
rect 23808 8991 23842 9025
rect 23876 8991 23910 9025
rect 23944 8991 23978 9025
rect 24012 8991 24046 9025
rect 24080 8991 24114 9025
rect 24148 8991 24159 9025
rect 23600 8985 24159 8991
rect 22766 8951 24159 8985
rect 22766 8950 23638 8951
rect 22766 8916 22818 8950
rect 22852 8916 22886 8950
rect 22920 8916 22954 8950
rect 22988 8916 23022 8950
rect 23056 8916 23090 8950
rect 23124 8916 23158 8950
rect 23192 8916 23226 8950
rect 23260 8916 23294 8950
rect 23328 8916 23362 8950
rect 23396 8916 23430 8950
rect 23464 8916 23498 8950
rect 23532 8916 23566 8950
rect 23600 8917 23638 8950
rect 23672 8917 23706 8951
rect 23740 8917 23774 8951
rect 23808 8917 23842 8951
rect 23876 8917 23910 8951
rect 23944 8917 23978 8951
rect 24012 8917 24046 8951
rect 24080 8917 24114 8951
rect 24148 8917 24159 8951
rect 23600 8916 24159 8917
rect 22766 8881 24159 8916
rect 22766 8847 22818 8881
rect 22852 8847 22886 8881
rect 22920 8847 22954 8881
rect 22988 8847 23022 8881
rect 23056 8847 23090 8881
rect 23124 8847 23158 8881
rect 23192 8847 23226 8881
rect 23260 8847 23294 8881
rect 23328 8847 23362 8881
rect 23396 8847 23430 8881
rect 23464 8847 23498 8881
rect 23532 8847 23566 8881
rect 23600 8877 24159 8881
rect 23600 8847 23638 8877
rect 22766 8843 23638 8847
rect 23672 8843 23706 8877
rect 23740 8843 23774 8877
rect 23808 8843 23842 8877
rect 23876 8843 23910 8877
rect 23944 8843 23978 8877
rect 24012 8843 24046 8877
rect 24080 8843 24114 8877
rect 24148 8843 24159 8877
rect 22766 8812 24159 8843
rect 22766 8778 22818 8812
rect 22852 8778 22886 8812
rect 22920 8778 22954 8812
rect 22988 8778 23022 8812
rect 23056 8778 23090 8812
rect 23124 8778 23158 8812
rect 23192 8778 23226 8812
rect 23260 8778 23294 8812
rect 23328 8778 23362 8812
rect 23396 8778 23430 8812
rect 23464 8778 23498 8812
rect 23532 8778 23566 8812
rect 23600 8803 24159 8812
rect 23600 8778 23638 8803
rect 22766 8769 23638 8778
rect 23672 8769 23706 8803
rect 23740 8769 23774 8803
rect 23808 8769 23842 8803
rect 23876 8769 23910 8803
rect 23944 8769 23978 8803
rect 24012 8769 24046 8803
rect 24080 8769 24114 8803
rect 24148 8769 24159 8803
rect 22766 8745 24159 8769
rect 22766 8743 23600 8745
rect 22766 8709 22818 8743
rect 22852 8709 22886 8743
rect 22920 8709 22954 8743
rect 22988 8709 23022 8743
rect 23056 8709 23090 8743
rect 23124 8709 23158 8743
rect 23192 8709 23226 8743
rect 23260 8709 23294 8743
rect 23328 8709 23362 8743
rect 23396 8709 23430 8743
rect 23464 8709 23498 8743
rect 23532 8709 23566 8743
rect 22766 8674 23600 8709
rect 22766 8640 22818 8674
rect 22852 8640 22886 8674
rect 22920 8640 22954 8674
rect 22988 8640 23022 8674
rect 23056 8640 23090 8674
rect 23124 8640 23158 8674
rect 23192 8640 23226 8674
rect 23260 8640 23294 8674
rect 23328 8640 23362 8674
rect 23396 8640 23430 8674
rect 23464 8640 23498 8674
rect 23532 8640 23566 8674
rect 22766 8605 23600 8640
rect 22766 8571 22818 8605
rect 22852 8571 22886 8605
rect 22920 8571 22954 8605
rect 22988 8571 23022 8605
rect 23056 8571 23090 8605
rect 23124 8571 23158 8605
rect 23192 8571 23226 8605
rect 23260 8571 23294 8605
rect 23328 8571 23362 8605
rect 23396 8571 23430 8605
rect 23464 8571 23498 8605
rect 23532 8571 23566 8605
rect 22766 8536 23600 8571
rect 22766 8502 22818 8536
rect 22852 8502 22886 8536
rect 22920 8502 22954 8536
rect 22988 8502 23022 8536
rect 23056 8502 23090 8536
rect 23124 8502 23158 8536
rect 23192 8502 23226 8536
rect 23260 8502 23294 8536
rect 23328 8502 23362 8536
rect 23396 8502 23430 8536
rect 23464 8502 23498 8536
rect 23532 8502 23566 8536
rect 22766 8467 23600 8502
rect 22766 8433 22818 8467
rect 22852 8433 22886 8467
rect 22920 8433 22954 8467
rect 22988 8433 23022 8467
rect 23056 8433 23090 8467
rect 23124 8433 23158 8467
rect 23192 8433 23226 8467
rect 23260 8433 23294 8467
rect 23328 8433 23362 8467
rect 23396 8433 23430 8467
rect 23464 8433 23498 8467
rect 23532 8433 23566 8467
rect 22766 8398 23600 8433
rect 22766 8364 22818 8398
rect 22852 8364 22886 8398
rect 22920 8364 22954 8398
rect 22988 8364 23022 8398
rect 23056 8364 23090 8398
rect 23124 8364 23158 8398
rect 23192 8364 23226 8398
rect 23260 8364 23294 8398
rect 23328 8364 23362 8398
rect 23396 8364 23430 8398
rect 23464 8364 23498 8398
rect 23532 8364 23566 8398
rect 22766 8329 23600 8364
rect 22766 8295 22818 8329
rect 22852 8295 22886 8329
rect 22920 8295 22954 8329
rect 22988 8295 23022 8329
rect 23056 8295 23090 8329
rect 23124 8295 23158 8329
rect 23192 8295 23226 8329
rect 23260 8295 23294 8329
rect 23328 8295 23362 8329
rect 23396 8295 23430 8329
rect 23464 8295 23498 8329
rect 23532 8295 23566 8329
rect 22766 8260 23600 8295
rect 22766 8226 22818 8260
rect 22852 8226 22886 8260
rect 22920 8226 22954 8260
rect 22988 8226 23022 8260
rect 23056 8226 23090 8260
rect 23124 8226 23158 8260
rect 23192 8226 23226 8260
rect 23260 8226 23294 8260
rect 23328 8226 23362 8260
rect 23396 8226 23430 8260
rect 23464 8226 23498 8260
rect 23532 8226 23566 8260
rect 22766 8191 23600 8226
rect 22766 8157 22818 8191
rect 22852 8157 22886 8191
rect 22920 8157 22954 8191
rect 22988 8157 23022 8191
rect 23056 8157 23090 8191
rect 23124 8157 23158 8191
rect 23192 8157 23226 8191
rect 23260 8157 23294 8191
rect 23328 8157 23362 8191
rect 23396 8157 23430 8191
rect 23464 8157 23498 8191
rect 23532 8157 23566 8191
rect 22766 8122 23600 8157
rect 22766 8088 22818 8122
rect 22852 8088 22886 8122
rect 22920 8088 22954 8122
rect 22988 8088 23022 8122
rect 23056 8088 23090 8122
rect 23124 8088 23158 8122
rect 23192 8088 23226 8122
rect 23260 8088 23294 8122
rect 23328 8088 23362 8122
rect 23396 8088 23430 8122
rect 23464 8088 23498 8122
rect 23532 8088 23566 8122
rect 22766 8053 23600 8088
rect 22766 8019 22818 8053
rect 22852 8019 22886 8053
rect 22920 8019 22954 8053
rect 22988 8019 23022 8053
rect 23056 8019 23090 8053
rect 23124 8019 23158 8053
rect 23192 8019 23226 8053
rect 23260 8019 23294 8053
rect 23328 8019 23362 8053
rect 23396 8019 23430 8053
rect 23464 8019 23498 8053
rect 23532 8019 23566 8053
rect 22766 7984 23600 8019
rect 22766 7950 22818 7984
rect 22852 7950 22886 7984
rect 22920 7950 22954 7984
rect 22988 7950 23022 7984
rect 23056 7950 23090 7984
rect 23124 7950 23158 7984
rect 23192 7950 23226 7984
rect 23260 7950 23294 7984
rect 23328 7950 23362 7984
rect 23396 7950 23430 7984
rect 23464 7950 23498 7984
rect 23532 7950 23566 7984
rect 22766 7915 23600 7950
rect 22766 7881 22818 7915
rect 22852 7881 22886 7915
rect 22920 7881 22954 7915
rect 22988 7881 23022 7915
rect 23056 7881 23090 7915
rect 23124 7881 23158 7915
rect 23192 7881 23226 7915
rect 23260 7881 23294 7915
rect 23328 7881 23362 7915
rect 23396 7881 23430 7915
rect 23464 7881 23498 7915
rect 23532 7881 23566 7915
rect 22766 7846 23600 7881
rect 22766 7812 22818 7846
rect 22852 7812 22886 7846
rect 22920 7812 22954 7846
rect 22988 7812 23022 7846
rect 23056 7812 23090 7846
rect 23124 7812 23158 7846
rect 23192 7812 23226 7846
rect 23260 7812 23294 7846
rect 23328 7812 23362 7846
rect 23396 7812 23430 7846
rect 23464 7812 23498 7846
rect 23532 7812 23566 7846
rect 22766 7777 23600 7812
rect 22766 7743 22818 7777
rect 22852 7743 22886 7777
rect 22920 7743 22954 7777
rect 22988 7743 23022 7777
rect 23056 7743 23090 7777
rect 23124 7743 23158 7777
rect 23192 7743 23226 7777
rect 23260 7743 23294 7777
rect 23328 7743 23362 7777
rect 23396 7743 23430 7777
rect 23464 7743 23498 7777
rect 23532 7743 23566 7777
rect 22766 7708 23600 7743
rect 22766 7674 22818 7708
rect 22852 7674 22886 7708
rect 22920 7674 22954 7708
rect 22988 7674 23022 7708
rect 23056 7674 23090 7708
rect 23124 7674 23158 7708
rect 23192 7674 23226 7708
rect 23260 7674 23294 7708
rect 23328 7674 23362 7708
rect 23396 7674 23430 7708
rect 23464 7674 23498 7708
rect 23532 7674 23566 7708
rect 22766 7639 23600 7674
rect 22766 7605 22818 7639
rect 22852 7605 22886 7639
rect 22920 7605 22954 7639
rect 22988 7605 23022 7639
rect 23056 7605 23090 7639
rect 23124 7605 23158 7639
rect 23192 7605 23226 7639
rect 23260 7605 23294 7639
rect 23328 7605 23362 7639
rect 23396 7605 23430 7639
rect 23464 7605 23498 7639
rect 23532 7605 23566 7639
rect 22766 7570 23600 7605
rect 22766 7536 22818 7570
rect 22852 7536 22886 7570
rect 22920 7536 22954 7570
rect 22988 7536 23022 7570
rect 23056 7536 23090 7570
rect 23124 7536 23158 7570
rect 23192 7536 23226 7570
rect 23260 7536 23294 7570
rect 23328 7536 23362 7570
rect 23396 7536 23430 7570
rect 23464 7536 23498 7570
rect 23532 7536 23566 7570
rect 22766 7501 23600 7536
rect 22766 7467 22818 7501
rect 22852 7467 22886 7501
rect 22920 7467 22954 7501
rect 22988 7467 23022 7501
rect 23056 7467 23090 7501
rect 23124 7467 23158 7501
rect 23192 7467 23226 7501
rect 23260 7467 23294 7501
rect 23328 7467 23362 7501
rect 23396 7467 23430 7501
rect 23464 7467 23498 7501
rect 23532 7467 23566 7501
rect 22766 7432 23600 7467
rect 22766 7398 22818 7432
rect 22852 7398 22886 7432
rect 22920 7398 22954 7432
rect 22988 7398 23022 7432
rect 23056 7398 23090 7432
rect 23124 7398 23158 7432
rect 23192 7398 23226 7432
rect 23260 7398 23294 7432
rect 23328 7398 23362 7432
rect 23396 7398 23430 7432
rect 23464 7398 23498 7432
rect 23532 7398 23566 7432
rect 22766 7363 23600 7398
rect 22766 7329 22818 7363
rect 22852 7329 22886 7363
rect 22920 7329 22954 7363
rect 22988 7329 23022 7363
rect 23056 7329 23090 7363
rect 23124 7329 23158 7363
rect 23192 7329 23226 7363
rect 23260 7329 23294 7363
rect 23328 7329 23362 7363
rect 23396 7329 23430 7363
rect 23464 7329 23498 7363
rect 23532 7329 23566 7363
rect 22766 7294 23600 7329
rect 22766 7260 22818 7294
rect 22852 7260 22886 7294
rect 22920 7260 22954 7294
rect 22988 7260 23022 7294
rect 23056 7260 23090 7294
rect 23124 7260 23158 7294
rect 23192 7260 23226 7294
rect 23260 7260 23294 7294
rect 23328 7260 23362 7294
rect 23396 7260 23430 7294
rect 23464 7260 23498 7294
rect 23532 7260 23566 7294
rect 22766 7225 23600 7260
rect 22766 7191 22818 7225
rect 22852 7191 22886 7225
rect 22920 7191 22954 7225
rect 22988 7191 23022 7225
rect 23056 7191 23090 7225
rect 23124 7191 23158 7225
rect 23192 7191 23226 7225
rect 23260 7191 23294 7225
rect 23328 7191 23362 7225
rect 23396 7191 23430 7225
rect 23464 7191 23498 7225
rect 23532 7191 23566 7225
rect 22766 7156 23600 7191
rect 22766 7122 22818 7156
rect 22852 7122 22886 7156
rect 22920 7122 22954 7156
rect 22988 7122 23022 7156
rect 23056 7122 23090 7156
rect 23124 7122 23158 7156
rect 23192 7122 23226 7156
rect 23260 7122 23294 7156
rect 23328 7122 23362 7156
rect 23396 7122 23430 7156
rect 23464 7122 23498 7156
rect 23532 7122 23566 7156
rect 22766 7087 23600 7122
rect 22766 7053 22818 7087
rect 22852 7053 22886 7087
rect 22920 7053 22954 7087
rect 22988 7053 23022 7087
rect 23056 7053 23090 7087
rect 23124 7053 23158 7087
rect 23192 7053 23226 7087
rect 23260 7053 23294 7087
rect 23328 7053 23362 7087
rect 23396 7053 23430 7087
rect 23464 7053 23498 7087
rect 23532 7053 23566 7087
rect 22766 7018 23600 7053
rect 22766 6984 22818 7018
rect 22852 6984 22886 7018
rect 22920 6984 22954 7018
rect 22988 6984 23022 7018
rect 23056 6984 23090 7018
rect 23124 6984 23158 7018
rect 23192 6984 23226 7018
rect 23260 6984 23294 7018
rect 23328 6984 23362 7018
rect 23396 6984 23430 7018
rect 23464 6984 23498 7018
rect 23532 6984 23566 7018
rect 22766 6949 23600 6984
rect 22766 6915 22818 6949
rect 22852 6915 22886 6949
rect 22920 6915 22954 6949
rect 22988 6915 23022 6949
rect 23056 6915 23090 6949
rect 23124 6915 23158 6949
rect 23192 6915 23226 6949
rect 23260 6915 23294 6949
rect 23328 6915 23362 6949
rect 23396 6915 23430 6949
rect 23464 6915 23498 6949
rect 23532 6915 23566 6949
rect 22766 6880 23600 6915
rect 22766 6846 22818 6880
rect 22852 6846 22886 6880
rect 22920 6846 22954 6880
rect 22988 6846 23022 6880
rect 23056 6846 23090 6880
rect 23124 6846 23158 6880
rect 23192 6846 23226 6880
rect 23260 6846 23294 6880
rect 23328 6846 23362 6880
rect 23396 6846 23430 6880
rect 23464 6846 23498 6880
rect 23532 6846 23566 6880
rect 22766 6811 23600 6846
rect 22766 5485 22818 6811
rect 22766 5463 23600 5485
rect 22766 5440 23796 5463
rect 22766 4794 22842 5440
rect 22944 5406 22979 5440
rect 23013 5406 23048 5440
rect 23082 5406 23117 5440
rect 23151 5406 23186 5440
rect 23220 5406 23255 5440
rect 23289 5406 23324 5440
rect 23358 5406 23393 5440
rect 23427 5406 23462 5440
rect 23496 5406 23531 5440
rect 23565 5406 23600 5440
rect 23634 5406 23669 5440
rect 23703 5406 23738 5440
rect 23772 5406 23796 5440
rect 22944 5372 23796 5406
rect 22944 5338 22979 5372
rect 23013 5338 23048 5372
rect 23082 5338 23117 5372
rect 23151 5338 23186 5372
rect 23220 5338 23255 5372
rect 23289 5338 23324 5372
rect 23358 5338 23393 5372
rect 23427 5338 23462 5372
rect 23496 5338 23531 5372
rect 23565 5338 23600 5372
rect 23634 5338 23669 5372
rect 23703 5338 23738 5372
rect 23772 5338 23796 5372
rect 22944 5304 23796 5338
rect 22944 5270 22979 5304
rect 23013 5270 23048 5304
rect 23082 5270 23117 5304
rect 23151 5270 23186 5304
rect 23220 5270 23255 5304
rect 23289 5270 23324 5304
rect 23358 5270 23393 5304
rect 23427 5270 23462 5304
rect 23496 5270 23531 5304
rect 23565 5270 23600 5304
rect 23634 5270 23669 5304
rect 23703 5270 23738 5304
rect 23772 5270 23796 5304
rect 22944 5236 23796 5270
rect 22944 5202 22979 5236
rect 23013 5202 23048 5236
rect 23082 5202 23117 5236
rect 23151 5202 23186 5236
rect 23220 5202 23255 5236
rect 23289 5202 23324 5236
rect 23358 5202 23393 5236
rect 23427 5202 23462 5236
rect 23496 5202 23531 5236
rect 23565 5202 23600 5236
rect 23634 5202 23669 5236
rect 23703 5202 23738 5236
rect 23772 5202 23796 5236
rect 22944 5168 23796 5202
rect 22944 5134 22979 5168
rect 23013 5134 23048 5168
rect 23082 5134 23117 5168
rect 23151 5134 23186 5168
rect 23220 5134 23255 5168
rect 23289 5134 23324 5168
rect 23358 5134 23393 5168
rect 23427 5134 23462 5168
rect 23496 5134 23531 5168
rect 23565 5134 23600 5168
rect 23634 5134 23669 5168
rect 23703 5134 23738 5168
rect 23772 5134 23796 5168
rect 22944 5100 23796 5134
rect 22944 5066 22979 5100
rect 23013 5066 23048 5100
rect 23082 5066 23117 5100
rect 23151 5066 23186 5100
rect 23220 5066 23255 5100
rect 23289 5066 23324 5100
rect 23358 5066 23393 5100
rect 23427 5066 23462 5100
rect 23496 5066 23531 5100
rect 23565 5066 23600 5100
rect 23634 5066 23669 5100
rect 23703 5066 23738 5100
rect 23772 5066 23796 5100
rect 22944 5032 23796 5066
rect 22944 4998 22979 5032
rect 23013 4998 23048 5032
rect 23082 4998 23117 5032
rect 23151 4998 23186 5032
rect 23220 4998 23255 5032
rect 23289 4998 23324 5032
rect 23358 4998 23393 5032
rect 23427 4998 23462 5032
rect 23496 4998 23531 5032
rect 23565 4998 23600 5032
rect 23634 4998 23669 5032
rect 23703 4998 23738 5032
rect 23772 4998 23796 5032
rect 22944 4964 23796 4998
rect 22944 4930 22979 4964
rect 23013 4930 23048 4964
rect 23082 4930 23117 4964
rect 23151 4930 23186 4964
rect 23220 4930 23255 4964
rect 23289 4930 23324 4964
rect 23358 4930 23393 4964
rect 23427 4930 23462 4964
rect 23496 4930 23531 4964
rect 23565 4930 23600 4964
rect 23634 4930 23669 4964
rect 23703 4930 23738 4964
rect 23772 4930 23796 4964
rect 22944 4896 23796 4930
rect 22944 4862 22979 4896
rect 23013 4862 23048 4896
rect 23082 4862 23117 4896
rect 23151 4862 23186 4896
rect 23220 4862 23255 4896
rect 23289 4862 23324 4896
rect 23358 4862 23393 4896
rect 23427 4862 23462 4896
rect 23496 4862 23531 4896
rect 23565 4862 23600 4896
rect 23634 4862 23669 4896
rect 23703 4862 23738 4896
rect 23772 4862 23796 4896
rect 22944 4828 23796 4862
rect 22944 4794 22979 4828
rect 23013 4794 23048 4828
rect 23082 4794 23117 4828
rect 23151 4794 23186 4828
rect 23220 4794 23255 4828
rect 23289 4794 23324 4828
rect 23358 4794 23393 4828
rect 23427 4794 23462 4828
rect 23496 4794 23531 4828
rect 23565 4794 23600 4828
rect 23634 4794 23669 4828
rect 23703 4794 23738 4828
rect 23772 4794 23796 4828
rect 22766 4771 23796 4794
rect 696 4737 866 4771
rect 730 4703 764 4737
rect 798 4703 832 4737
rect 696 4665 866 4703
rect 730 4631 764 4665
rect 798 4631 832 4665
rect 696 4593 866 4631
rect 730 4559 764 4593
rect 798 4559 832 4593
rect 23568 4737 23796 4771
rect 23568 4703 23597 4737
rect 23631 4703 23665 4737
rect 23699 4703 23733 4737
rect 23767 4703 23796 4737
rect 23568 4668 23796 4703
rect 23568 4634 23597 4668
rect 23631 4634 23665 4668
rect 23699 4634 23733 4668
rect 23767 4634 23796 4668
rect 23568 4599 23796 4634
rect 696 4521 866 4559
rect 730 4487 764 4521
rect 798 4487 832 4521
rect 696 4449 866 4487
rect 730 4415 764 4449
rect 798 4415 832 4449
rect 696 4377 866 4415
rect 730 4343 764 4377
rect 798 4343 832 4377
rect 696 4305 866 4343
rect 730 4271 764 4305
rect 798 4271 832 4305
rect 696 4233 866 4271
rect 730 4199 764 4233
rect 798 4199 832 4233
rect 696 4161 866 4199
rect 730 4127 764 4161
rect 798 4127 832 4161
rect 696 4089 866 4127
rect 730 4055 764 4089
rect 798 4055 832 4089
rect 696 4017 866 4055
rect 730 3983 764 4017
rect 798 3983 832 4017
rect 696 3946 866 3983
rect 730 3912 764 3946
rect 798 3912 832 3946
rect 696 3875 866 3912
rect 730 3841 764 3875
rect 798 3841 832 3875
rect 696 3804 866 3841
rect 730 3770 764 3804
rect 798 3770 832 3804
rect 696 3733 866 3770
rect 730 3699 764 3733
rect 798 3699 832 3733
rect 696 3662 866 3699
rect 730 3628 764 3662
rect 798 3628 832 3662
rect 696 3591 866 3628
rect 730 3557 764 3591
rect 798 3557 832 3591
rect 696 3520 866 3557
rect 730 3486 764 3520
rect 798 3486 832 3520
rect 696 3449 866 3486
rect 730 3415 764 3449
rect 798 3415 832 3449
rect 696 3378 866 3415
rect 730 3344 764 3378
rect 798 3344 832 3378
rect 696 3286 866 3344
rect 730 3252 764 3286
rect 798 3252 832 3286
rect 696 3217 866 3252
rect 696 3216 764 3217
rect 730 3183 764 3216
rect 798 3183 832 3217
rect 730 3182 866 3183
rect 696 3148 866 3182
rect 696 3146 764 3148
rect 730 3114 764 3146
rect 798 3114 832 3148
rect 730 3112 866 3114
rect 696 3079 866 3112
rect 696 3076 764 3079
rect 730 3045 764 3076
rect 798 3045 832 3079
rect 730 3042 866 3045
rect 696 3010 866 3042
rect 696 3006 764 3010
rect 730 2976 764 3006
rect 798 2976 832 3010
rect 730 2972 866 2976
rect 696 2941 866 2972
rect 696 2937 764 2941
rect 730 2903 764 2937
rect 696 2868 764 2903
rect 730 2834 764 2868
rect 696 2799 764 2834
rect 730 2765 764 2799
rect 696 2730 764 2765
rect 730 2696 764 2730
rect 696 2661 764 2696
rect 730 2627 764 2661
rect 696 2592 764 2627
rect 730 2558 764 2592
rect 696 2523 764 2558
rect 730 2489 764 2523
rect 696 2454 764 2489
rect 730 2420 764 2454
rect 696 2385 764 2420
rect 730 2351 764 2385
rect 696 2316 764 2351
rect 730 2282 764 2316
rect 696 2247 764 2282
rect 730 2213 764 2247
rect 696 2178 764 2213
rect 730 2144 764 2178
rect 696 2109 764 2144
rect 730 2075 764 2109
rect 696 2040 764 2075
rect 730 2006 764 2040
rect 696 1971 764 2006
rect 730 1937 764 1971
rect 696 1902 764 1937
rect 730 1868 764 1902
rect 696 1833 764 1868
rect 730 1799 764 1833
rect 696 1764 764 1799
rect 730 1730 764 1764
rect 696 1695 764 1730
rect 730 1661 764 1695
rect 696 1626 764 1661
rect 730 1592 764 1626
rect 696 1557 764 1592
rect 730 1523 764 1557
rect 696 1488 764 1523
rect 730 1454 764 1488
rect 696 1419 764 1454
rect 730 1385 764 1419
rect 696 1350 764 1385
rect 730 1316 764 1350
rect 696 1281 764 1316
rect 730 1247 764 1281
rect 23568 4565 23597 4599
rect 23631 4565 23665 4599
rect 23699 4565 23733 4599
rect 23767 4565 23796 4599
rect 23568 4530 23796 4565
rect 23568 4496 23597 4530
rect 23631 4496 23665 4530
rect 23699 4496 23733 4530
rect 23767 4496 23796 4530
rect 23568 4461 23796 4496
rect 23568 4427 23597 4461
rect 23631 4427 23665 4461
rect 23699 4427 23733 4461
rect 23767 4427 23796 4461
rect 23568 4392 23796 4427
rect 23568 4358 23597 4392
rect 23631 4358 23665 4392
rect 23699 4358 23733 4392
rect 23767 4358 23796 4392
rect 23568 4323 23796 4358
rect 23568 4289 23597 4323
rect 23631 4289 23665 4323
rect 23699 4289 23733 4323
rect 23767 4289 23796 4323
rect 23568 4254 23796 4289
rect 23568 4220 23597 4254
rect 23631 4220 23665 4254
rect 23699 4220 23733 4254
rect 23767 4220 23796 4254
rect 23568 4185 23796 4220
rect 23568 4151 23597 4185
rect 23631 4151 23665 4185
rect 23699 4151 23733 4185
rect 23767 4151 23796 4185
rect 23568 4116 23796 4151
rect 23568 2110 23597 4116
rect 23767 2110 23796 4116
rect 23568 2076 23796 2110
rect 13728 2052 14489 2076
rect 13728 2018 13751 2052
rect 13785 2018 13819 2052
rect 13853 2018 13887 2052
rect 13921 2018 13955 2052
rect 13989 2018 14023 2052
rect 14057 2018 14091 2052
rect 14125 2018 14159 2052
rect 14193 2018 14227 2052
rect 14261 2018 14295 2052
rect 14329 2018 14363 2052
rect 14397 2042 14489 2052
rect 14523 2042 14567 2076
rect 14601 2061 23796 2076
rect 14601 2042 14701 2061
rect 14397 2018 14701 2042
rect 13728 2008 14701 2018
rect 13728 1980 14545 2008
rect 13728 1946 13751 1980
rect 13785 1946 13819 1980
rect 13853 1946 13887 1980
rect 13921 1946 13955 1980
rect 13989 1946 14023 1980
rect 14057 1946 14091 1980
rect 14125 1946 14159 1980
rect 14193 1946 14227 1980
rect 14261 1946 14295 1980
rect 14329 1946 14363 1980
rect 14397 1974 14545 1980
rect 14579 1974 14701 2008
rect 14397 1968 14701 1974
rect 14397 1946 14455 1968
rect 13728 1934 14455 1946
rect 14489 1939 14701 1968
rect 14489 1934 14523 1939
rect 13728 1908 14523 1934
rect 13728 1874 13751 1908
rect 13785 1874 13819 1908
rect 13853 1874 13887 1908
rect 13921 1874 13955 1908
rect 13989 1874 14023 1908
rect 14057 1874 14091 1908
rect 14125 1874 14159 1908
rect 14193 1874 14227 1908
rect 14261 1874 14295 1908
rect 14329 1874 14363 1908
rect 14397 1905 14523 1908
rect 14557 1916 14701 1939
rect 14557 1905 14591 1916
rect 14397 1897 14591 1905
rect 14397 1874 14455 1897
rect 13728 1863 14455 1874
rect 14489 1882 14591 1897
rect 14625 1882 14701 1916
rect 14489 1870 14701 1882
rect 14489 1863 14523 1870
rect 13728 1836 14523 1863
rect 14557 1846 14701 1870
rect 14557 1836 14591 1846
rect 13728 1802 13751 1836
rect 13785 1802 13819 1836
rect 13853 1802 13887 1836
rect 13921 1802 13955 1836
rect 13989 1802 14023 1836
rect 14057 1802 14091 1836
rect 14125 1802 14159 1836
rect 14193 1802 14227 1836
rect 14261 1802 14295 1836
rect 14329 1802 14363 1836
rect 14397 1826 14591 1836
rect 14397 1802 14455 1826
rect 13728 1792 14455 1802
rect 14489 1812 14591 1826
rect 14625 1812 14701 1846
rect 14489 1801 14701 1812
rect 14489 1792 14523 1801
rect 13728 1767 14523 1792
rect 14557 1776 14701 1801
rect 14557 1767 14591 1776
rect 13728 1764 14591 1767
rect 13728 1730 13751 1764
rect 13785 1730 13819 1764
rect 13853 1730 13887 1764
rect 13921 1730 13955 1764
rect 13989 1730 14023 1764
rect 14057 1730 14091 1764
rect 14125 1730 14159 1764
rect 14193 1730 14227 1764
rect 14261 1730 14295 1764
rect 14329 1730 14363 1764
rect 14397 1755 14591 1764
rect 14397 1730 14455 1755
rect 13728 1721 14455 1730
rect 14489 1742 14591 1755
rect 14625 1742 14701 1776
rect 14489 1732 14701 1742
rect 14489 1721 14523 1732
rect 13728 1698 14523 1721
rect 14557 1706 14701 1732
rect 14557 1698 14591 1706
rect 13728 1692 14591 1698
rect 13728 1658 13751 1692
rect 13785 1658 13819 1692
rect 13853 1658 13887 1692
rect 13921 1658 13955 1692
rect 13989 1658 14023 1692
rect 14057 1658 14091 1692
rect 14125 1658 14159 1692
rect 14193 1658 14227 1692
rect 14261 1658 14295 1692
rect 14329 1658 14363 1692
rect 14397 1684 14591 1692
rect 14397 1658 14455 1684
rect 13728 1650 14455 1658
rect 14489 1672 14591 1684
rect 14625 1672 14701 1706
rect 14489 1663 14701 1672
rect 14489 1650 14523 1663
rect 13728 1629 14523 1650
rect 14557 1636 14701 1663
rect 14557 1629 14591 1636
rect 13728 1620 14591 1629
rect 13728 1586 13751 1620
rect 13785 1586 13819 1620
rect 13853 1586 13887 1620
rect 13921 1586 13955 1620
rect 13989 1586 14023 1620
rect 14057 1586 14091 1620
rect 14125 1586 14159 1620
rect 14193 1586 14227 1620
rect 14261 1586 14295 1620
rect 14329 1586 14363 1620
rect 14397 1613 14591 1620
rect 14397 1586 14455 1613
rect 13728 1579 14455 1586
rect 14489 1602 14591 1613
rect 14625 1602 14701 1636
rect 14489 1594 14701 1602
rect 14489 1579 14523 1594
rect 13728 1560 14523 1579
rect 14557 1566 14701 1594
rect 14557 1560 14591 1566
rect 13728 1548 14591 1560
rect 13728 1514 13751 1548
rect 13785 1514 13819 1548
rect 13853 1514 13887 1548
rect 13921 1514 13955 1548
rect 13989 1514 14023 1548
rect 14057 1514 14091 1548
rect 14125 1514 14159 1548
rect 14193 1514 14227 1548
rect 14261 1514 14295 1548
rect 14329 1514 14363 1548
rect 14397 1541 14591 1548
rect 14397 1514 14455 1541
rect 13728 1507 14455 1514
rect 14489 1532 14591 1541
rect 14625 1532 14701 1566
rect 14489 1525 14701 1532
rect 14489 1507 14523 1525
rect 13728 1491 14523 1507
rect 14557 1496 14701 1525
rect 14557 1491 14591 1496
rect 13728 1475 14591 1491
rect 13728 1441 13751 1475
rect 13785 1441 13819 1475
rect 13853 1441 13887 1475
rect 13921 1441 13955 1475
rect 13989 1441 14023 1475
rect 14057 1441 14091 1475
rect 14125 1441 14159 1475
rect 14193 1441 14227 1475
rect 14261 1441 14295 1475
rect 14329 1441 14363 1475
rect 14397 1469 14591 1475
rect 14397 1441 14455 1469
rect 13728 1435 14455 1441
rect 14489 1462 14591 1469
rect 14625 1462 14701 1496
rect 14489 1456 14701 1462
rect 14489 1435 14523 1456
rect 13728 1422 14523 1435
rect 14557 1426 14701 1456
rect 14557 1422 14591 1426
rect 13728 1402 14591 1422
rect 13728 1368 13751 1402
rect 13785 1368 13819 1402
rect 13853 1368 13887 1402
rect 13921 1368 13955 1402
rect 13989 1368 14023 1402
rect 14057 1368 14091 1402
rect 14125 1368 14159 1402
rect 14193 1368 14227 1402
rect 14261 1368 14295 1402
rect 14329 1368 14363 1402
rect 14397 1397 14591 1402
rect 14397 1368 14455 1397
rect 13728 1363 14455 1368
rect 14489 1392 14591 1397
rect 14625 1392 14701 1426
rect 14489 1387 14701 1392
rect 14489 1363 14523 1387
rect 13728 1353 14523 1363
rect 14557 1356 14701 1387
rect 14557 1353 14591 1356
rect 13728 1329 14591 1353
rect 13728 1267 13751 1329
rect 866 1261 13751 1267
rect 14397 1325 14591 1329
rect 14397 1291 14455 1325
rect 14489 1322 14591 1325
rect 14625 1322 14701 1356
rect 14489 1318 14701 1322
rect 14489 1291 14523 1318
rect 14397 1284 14523 1291
rect 14557 1286 14701 1318
rect 14557 1284 14591 1286
rect 696 1212 764 1247
rect 730 1178 764 1212
rect 696 1143 764 1178
rect 730 1109 764 1143
rect 696 1074 764 1109
rect 934 1227 969 1261
rect 1003 1227 1038 1261
rect 1072 1227 1107 1261
rect 1141 1227 1176 1261
rect 1210 1227 1245 1261
rect 1279 1227 1314 1261
rect 1348 1227 1383 1261
rect 1417 1227 1452 1261
rect 1486 1227 1521 1261
rect 1555 1227 1590 1261
rect 1624 1227 1659 1261
rect 1693 1227 1728 1261
rect 1762 1227 1797 1261
rect 1831 1227 1866 1261
rect 1900 1227 1935 1261
rect 1969 1227 2004 1261
rect 2038 1227 2073 1261
rect 2107 1227 2142 1261
rect 2176 1227 2211 1261
rect 2245 1227 2280 1261
rect 2314 1227 2349 1261
rect 2383 1227 2418 1261
rect 2452 1227 2487 1261
rect 2521 1227 2556 1261
rect 2590 1227 2625 1261
rect 2659 1227 2694 1261
rect 2728 1227 2763 1261
rect 2797 1227 2832 1261
rect 2866 1227 2901 1261
rect 2935 1227 2970 1261
rect 3004 1227 3039 1261
rect 3073 1227 3108 1261
rect 3142 1227 3177 1261
rect 3211 1227 3246 1261
rect 3280 1227 3315 1261
rect 3349 1227 3384 1261
rect 3418 1227 3453 1261
rect 3487 1227 3522 1261
rect 3556 1227 3591 1261
rect 3625 1227 3660 1261
rect 3694 1227 3729 1261
rect 3763 1227 3798 1261
rect 3832 1227 3867 1261
rect 3901 1227 3936 1261
rect 3970 1227 4005 1261
rect 4039 1227 4074 1261
rect 4108 1227 4143 1261
rect 4177 1227 4212 1261
rect 4246 1227 4281 1261
rect 4315 1227 4350 1261
rect 4384 1227 4419 1261
rect 4453 1227 4488 1261
rect 4522 1227 4557 1261
rect 4591 1227 4626 1261
rect 4660 1227 4695 1261
rect 4729 1227 4764 1261
rect 4798 1227 4833 1261
rect 4867 1227 4902 1261
rect 4936 1227 4971 1261
rect 5005 1227 5040 1261
rect 5074 1227 5109 1261
rect 5143 1227 5178 1261
rect 5212 1227 5247 1261
rect 5281 1227 5316 1261
rect 5350 1227 5385 1261
rect 5419 1227 5454 1261
rect 5488 1227 5523 1261
rect 934 1193 5523 1227
rect 934 1159 969 1193
rect 1003 1159 1038 1193
rect 1072 1159 1107 1193
rect 1141 1159 1176 1193
rect 1210 1159 1245 1193
rect 1279 1159 1314 1193
rect 1348 1159 1383 1193
rect 1417 1159 1452 1193
rect 1486 1159 1521 1193
rect 1555 1159 1590 1193
rect 1624 1159 1659 1193
rect 1693 1159 1728 1193
rect 1762 1159 1797 1193
rect 1831 1159 1866 1193
rect 1900 1159 1935 1193
rect 1969 1159 2004 1193
rect 2038 1159 2073 1193
rect 2107 1159 2142 1193
rect 2176 1159 2211 1193
rect 2245 1159 2280 1193
rect 2314 1159 2349 1193
rect 2383 1159 2418 1193
rect 2452 1159 2487 1193
rect 2521 1159 2556 1193
rect 2590 1159 2625 1193
rect 2659 1159 2694 1193
rect 2728 1159 2763 1193
rect 2797 1159 2832 1193
rect 2866 1159 2901 1193
rect 2935 1159 2970 1193
rect 3004 1159 3039 1193
rect 3073 1159 3108 1193
rect 3142 1159 3177 1193
rect 3211 1159 3246 1193
rect 3280 1159 3315 1193
rect 3349 1159 3384 1193
rect 3418 1159 3453 1193
rect 3487 1159 3522 1193
rect 3556 1159 3591 1193
rect 3625 1159 3660 1193
rect 3694 1159 3729 1193
rect 3763 1159 3798 1193
rect 3832 1159 3867 1193
rect 3901 1159 3936 1193
rect 3970 1159 4005 1193
rect 4039 1159 4074 1193
rect 4108 1159 4143 1193
rect 4177 1159 4212 1193
rect 4246 1159 4281 1193
rect 4315 1159 4350 1193
rect 4384 1159 4419 1193
rect 4453 1159 4488 1193
rect 4522 1159 4557 1193
rect 4591 1159 4626 1193
rect 4660 1159 4695 1193
rect 4729 1159 4764 1193
rect 4798 1159 4833 1193
rect 4867 1159 4902 1193
rect 4936 1159 4971 1193
rect 5005 1159 5040 1193
rect 5074 1159 5109 1193
rect 5143 1159 5178 1193
rect 5212 1159 5247 1193
rect 5281 1159 5316 1193
rect 5350 1159 5385 1193
rect 5419 1159 5454 1193
rect 5488 1159 5523 1193
rect 934 1125 5523 1159
rect 934 1091 969 1125
rect 1003 1091 1038 1125
rect 1072 1091 1107 1125
rect 1141 1091 1176 1125
rect 1210 1091 1245 1125
rect 1279 1091 1314 1125
rect 1348 1091 1383 1125
rect 1417 1091 1452 1125
rect 1486 1091 1521 1125
rect 1555 1091 1590 1125
rect 1624 1091 1659 1125
rect 1693 1091 1728 1125
rect 1762 1091 1797 1125
rect 1831 1091 1866 1125
rect 1900 1091 1935 1125
rect 1969 1091 2004 1125
rect 2038 1091 2073 1125
rect 2107 1091 2142 1125
rect 2176 1091 2211 1125
rect 2245 1091 2280 1125
rect 2314 1091 2349 1125
rect 2383 1091 2418 1125
rect 2452 1091 2487 1125
rect 2521 1091 2556 1125
rect 2590 1091 2625 1125
rect 2659 1091 2694 1125
rect 2728 1091 2763 1125
rect 2797 1091 2832 1125
rect 2866 1091 2901 1125
rect 2935 1091 2970 1125
rect 3004 1091 3039 1125
rect 3073 1091 3108 1125
rect 3142 1091 3177 1125
rect 3211 1091 3246 1125
rect 3280 1091 3315 1125
rect 3349 1091 3384 1125
rect 3418 1091 3453 1125
rect 3487 1091 3522 1125
rect 3556 1091 3591 1125
rect 3625 1091 3660 1125
rect 3694 1091 3729 1125
rect 3763 1091 3798 1125
rect 3832 1091 3867 1125
rect 3901 1091 3936 1125
rect 3970 1091 4005 1125
rect 4039 1091 4074 1125
rect 4108 1091 4143 1125
rect 4177 1091 4212 1125
rect 4246 1091 4281 1125
rect 4315 1091 4350 1125
rect 4384 1091 4419 1125
rect 4453 1091 4488 1125
rect 4522 1091 4557 1125
rect 4591 1091 4626 1125
rect 4660 1091 4695 1125
rect 4729 1091 4764 1125
rect 4798 1091 4833 1125
rect 4867 1091 4902 1125
rect 4936 1091 4971 1125
rect 5005 1091 5040 1125
rect 5074 1091 5109 1125
rect 5143 1091 5178 1125
rect 5212 1091 5247 1125
rect 5281 1091 5316 1125
rect 5350 1091 5385 1125
rect 5419 1091 5454 1125
rect 5488 1091 5523 1125
rect 14397 1253 14591 1284
rect 14397 1219 14455 1253
rect 14489 1252 14591 1253
rect 14625 1252 14701 1286
rect 14489 1249 14701 1252
rect 14489 1219 14523 1249
rect 14397 1215 14523 1219
rect 14557 1216 14701 1249
rect 14557 1215 14591 1216
rect 14397 1182 14591 1215
rect 14625 1182 14701 1216
rect 14397 1181 14701 1182
rect 14397 1147 14455 1181
rect 14489 1179 14701 1181
rect 14489 1147 14523 1179
rect 14397 1145 14523 1147
rect 14557 1146 14701 1179
rect 14557 1145 14591 1146
rect 14397 1112 14591 1145
rect 14625 1143 14701 1146
rect 19563 2027 19598 2061
rect 19632 2027 19667 2061
rect 19701 2027 19736 2061
rect 19770 2027 19805 2061
rect 19839 2027 19874 2061
rect 19908 2027 19943 2061
rect 19977 2027 20012 2061
rect 20046 2027 20081 2061
rect 20115 2027 20150 2061
rect 20184 2027 20219 2061
rect 20253 2027 20288 2061
rect 20322 2027 20357 2061
rect 20391 2027 20426 2061
rect 20460 2027 20495 2061
rect 20529 2027 20564 2061
rect 20598 2027 20633 2061
rect 20667 2027 20702 2061
rect 20736 2027 20771 2061
rect 20805 2027 20840 2061
rect 20874 2027 20909 2061
rect 20943 2027 20978 2061
rect 21012 2027 21047 2061
rect 21081 2027 21116 2061
rect 21150 2027 21185 2061
rect 21219 2027 21254 2061
rect 21288 2027 21323 2061
rect 21357 2027 21392 2061
rect 21426 2027 21461 2061
rect 21495 2027 21530 2061
rect 21564 2027 21599 2061
rect 21633 2027 21668 2061
rect 21702 2027 21737 2061
rect 21771 2027 21806 2061
rect 21840 2027 21875 2061
rect 21909 2027 21944 2061
rect 21978 2027 22013 2061
rect 22047 2027 22082 2061
rect 22116 2027 22151 2061
rect 22185 2027 22220 2061
rect 22254 2027 22289 2061
rect 22323 2027 22358 2061
rect 22392 2027 22427 2061
rect 22461 2027 22496 2061
rect 22530 2027 22565 2061
rect 22599 2027 22634 2061
rect 22668 2027 22703 2061
rect 22737 2027 22772 2061
rect 22806 2027 22841 2061
rect 22875 2027 22910 2061
rect 22944 2027 22979 2061
rect 23013 2027 23048 2061
rect 23082 2027 23117 2061
rect 23151 2027 23186 2061
rect 23220 2027 23255 2061
rect 23289 2027 23324 2061
rect 23358 2027 23393 2061
rect 23427 2027 23462 2061
rect 23496 2027 23531 2061
rect 23565 2027 23600 2061
rect 23634 2027 23669 2061
rect 23703 2027 23738 2061
rect 23772 2027 23796 2061
rect 19563 1993 23796 2027
rect 19563 1959 19598 1993
rect 19632 1959 19667 1993
rect 19701 1959 19736 1993
rect 19770 1959 19805 1993
rect 19839 1959 19874 1993
rect 19908 1959 19943 1993
rect 19977 1959 20012 1993
rect 20046 1959 20081 1993
rect 20115 1959 20150 1993
rect 20184 1959 20219 1993
rect 20253 1959 20288 1993
rect 20322 1959 20357 1993
rect 20391 1959 20426 1993
rect 20460 1959 20495 1993
rect 20529 1959 20564 1993
rect 20598 1959 20633 1993
rect 20667 1959 20702 1993
rect 20736 1959 20771 1993
rect 20805 1959 20840 1993
rect 20874 1959 20909 1993
rect 20943 1959 20978 1993
rect 21012 1959 21047 1993
rect 21081 1959 21116 1993
rect 21150 1959 21185 1993
rect 21219 1959 21254 1993
rect 21288 1959 21323 1993
rect 21357 1959 21392 1993
rect 21426 1959 21461 1993
rect 21495 1959 21530 1993
rect 21564 1959 21599 1993
rect 21633 1959 21668 1993
rect 21702 1959 21737 1993
rect 21771 1959 21806 1993
rect 21840 1959 21875 1993
rect 21909 1959 21944 1993
rect 21978 1959 22013 1993
rect 22047 1959 22082 1993
rect 22116 1959 22151 1993
rect 22185 1959 22220 1993
rect 22254 1959 22289 1993
rect 22323 1959 22358 1993
rect 22392 1959 22427 1993
rect 22461 1959 22496 1993
rect 22530 1959 22565 1993
rect 22599 1959 22634 1993
rect 22668 1959 22703 1993
rect 22737 1959 22772 1993
rect 22806 1959 22841 1993
rect 22875 1959 22910 1993
rect 22944 1959 22979 1993
rect 23013 1959 23048 1993
rect 23082 1959 23117 1993
rect 23151 1959 23186 1993
rect 23220 1959 23255 1993
rect 23289 1959 23324 1993
rect 23358 1959 23393 1993
rect 23427 1959 23462 1993
rect 23496 1959 23531 1993
rect 23565 1959 23600 1993
rect 23634 1959 23669 1993
rect 23703 1959 23738 1993
rect 23772 1959 23796 1993
rect 19563 1925 23796 1959
rect 19563 1891 19598 1925
rect 19632 1891 19667 1925
rect 19701 1891 19736 1925
rect 19770 1891 19805 1925
rect 19839 1891 19874 1925
rect 19908 1891 19943 1925
rect 19977 1891 20012 1925
rect 20046 1891 20081 1925
rect 20115 1891 20150 1925
rect 20184 1891 20219 1925
rect 20253 1891 20288 1925
rect 20322 1891 20357 1925
rect 20391 1891 20426 1925
rect 20460 1891 20495 1925
rect 20529 1891 20564 1925
rect 20598 1891 20633 1925
rect 20667 1891 20702 1925
rect 20736 1891 20771 1925
rect 20805 1891 20840 1925
rect 20874 1891 20909 1925
rect 20943 1891 20978 1925
rect 21012 1891 21047 1925
rect 21081 1891 21116 1925
rect 21150 1891 21185 1925
rect 21219 1891 21254 1925
rect 21288 1891 21323 1925
rect 21357 1891 21392 1925
rect 21426 1891 21461 1925
rect 21495 1891 21530 1925
rect 21564 1891 21599 1925
rect 21633 1891 21668 1925
rect 21702 1891 21737 1925
rect 21771 1891 21806 1925
rect 21840 1891 21875 1925
rect 21909 1891 21944 1925
rect 21978 1891 22013 1925
rect 22047 1891 22082 1925
rect 22116 1891 22151 1925
rect 22185 1891 22220 1925
rect 22254 1891 22289 1925
rect 22323 1891 22358 1925
rect 22392 1891 22427 1925
rect 22461 1891 22496 1925
rect 22530 1891 22565 1925
rect 22599 1891 22634 1925
rect 22668 1891 22703 1925
rect 22737 1891 22772 1925
rect 22806 1891 22841 1925
rect 22875 1891 22910 1925
rect 22944 1891 22979 1925
rect 23013 1891 23048 1925
rect 23082 1891 23117 1925
rect 23151 1891 23186 1925
rect 23220 1891 23255 1925
rect 23289 1891 23324 1925
rect 23358 1891 23393 1925
rect 23427 1891 23462 1925
rect 23496 1891 23531 1925
rect 23565 1891 23600 1925
rect 23634 1891 23669 1925
rect 23703 1891 23738 1925
rect 23772 1891 23796 1925
rect 19563 1857 23796 1891
rect 19563 1823 19598 1857
rect 19632 1823 19667 1857
rect 19701 1823 19736 1857
rect 19770 1823 19805 1857
rect 19839 1823 19874 1857
rect 19908 1823 19943 1857
rect 19977 1823 20012 1857
rect 20046 1823 20081 1857
rect 20115 1823 20150 1857
rect 20184 1823 20219 1857
rect 20253 1823 20288 1857
rect 20322 1823 20357 1857
rect 20391 1823 20426 1857
rect 20460 1823 20495 1857
rect 20529 1823 20564 1857
rect 20598 1823 20633 1857
rect 20667 1823 20702 1857
rect 20736 1823 20771 1857
rect 20805 1823 20840 1857
rect 20874 1823 20909 1857
rect 20943 1823 20978 1857
rect 21012 1823 21047 1857
rect 21081 1823 21116 1857
rect 21150 1823 21185 1857
rect 21219 1823 21254 1857
rect 21288 1823 21323 1857
rect 21357 1823 21392 1857
rect 21426 1823 21461 1857
rect 21495 1823 21530 1857
rect 21564 1823 21599 1857
rect 21633 1823 21668 1857
rect 21702 1823 21737 1857
rect 21771 1823 21806 1857
rect 21840 1823 21875 1857
rect 21909 1823 21944 1857
rect 21978 1823 22013 1857
rect 22047 1823 22082 1857
rect 22116 1823 22151 1857
rect 22185 1823 22220 1857
rect 22254 1823 22289 1857
rect 22323 1823 22358 1857
rect 22392 1823 22427 1857
rect 22461 1823 22496 1857
rect 22530 1823 22565 1857
rect 22599 1823 22634 1857
rect 22668 1823 22703 1857
rect 22737 1823 22772 1857
rect 22806 1823 22841 1857
rect 22875 1823 22910 1857
rect 22944 1823 22979 1857
rect 23013 1823 23048 1857
rect 23082 1823 23117 1857
rect 23151 1823 23186 1857
rect 23220 1823 23255 1857
rect 23289 1823 23324 1857
rect 23358 1823 23393 1857
rect 23427 1823 23462 1857
rect 23496 1823 23531 1857
rect 23565 1823 23600 1857
rect 23634 1823 23669 1857
rect 23703 1823 23738 1857
rect 23772 1823 23796 1857
rect 19563 1789 23796 1823
rect 19563 1755 19598 1789
rect 19632 1755 19667 1789
rect 19701 1755 19736 1789
rect 19770 1755 19805 1789
rect 19839 1755 19874 1789
rect 19908 1755 19943 1789
rect 19977 1755 20012 1789
rect 20046 1755 20081 1789
rect 20115 1755 20150 1789
rect 20184 1755 20219 1789
rect 20253 1755 20288 1789
rect 20322 1755 20357 1789
rect 20391 1755 20426 1789
rect 20460 1755 20495 1789
rect 20529 1755 20564 1789
rect 20598 1755 20633 1789
rect 20667 1755 20702 1789
rect 20736 1755 20771 1789
rect 20805 1755 20840 1789
rect 20874 1755 20909 1789
rect 20943 1755 20978 1789
rect 21012 1755 21047 1789
rect 21081 1755 21116 1789
rect 21150 1755 21185 1789
rect 21219 1755 21254 1789
rect 21288 1755 21323 1789
rect 21357 1755 21392 1789
rect 21426 1755 21461 1789
rect 21495 1755 21530 1789
rect 21564 1755 21599 1789
rect 21633 1755 21668 1789
rect 21702 1755 21737 1789
rect 21771 1755 21806 1789
rect 21840 1755 21875 1789
rect 21909 1755 21944 1789
rect 21978 1755 22013 1789
rect 22047 1755 22082 1789
rect 22116 1755 22151 1789
rect 22185 1755 22220 1789
rect 22254 1755 22289 1789
rect 22323 1755 22358 1789
rect 22392 1755 22427 1789
rect 22461 1755 22496 1789
rect 22530 1755 22565 1789
rect 22599 1755 22634 1789
rect 22668 1755 22703 1789
rect 22737 1755 22772 1789
rect 22806 1755 22841 1789
rect 22875 1755 22910 1789
rect 22944 1755 22979 1789
rect 23013 1755 23048 1789
rect 23082 1755 23117 1789
rect 23151 1755 23186 1789
rect 23220 1755 23255 1789
rect 23289 1755 23324 1789
rect 23358 1755 23393 1789
rect 23427 1755 23462 1789
rect 23496 1755 23531 1789
rect 23565 1755 23600 1789
rect 23634 1755 23669 1789
rect 23703 1755 23738 1789
rect 23772 1755 23796 1789
rect 19563 1721 23796 1755
rect 19563 1687 19598 1721
rect 19632 1687 19667 1721
rect 19701 1687 19736 1721
rect 19770 1687 19805 1721
rect 19839 1687 19874 1721
rect 19908 1687 19943 1721
rect 19977 1687 20012 1721
rect 20046 1687 20081 1721
rect 20115 1687 20150 1721
rect 20184 1687 20219 1721
rect 20253 1687 20288 1721
rect 20322 1687 20357 1721
rect 20391 1687 20426 1721
rect 20460 1687 20495 1721
rect 20529 1687 20564 1721
rect 20598 1687 20633 1721
rect 20667 1687 20702 1721
rect 20736 1687 20771 1721
rect 20805 1687 20840 1721
rect 20874 1687 20909 1721
rect 20943 1687 20978 1721
rect 21012 1687 21047 1721
rect 21081 1687 21116 1721
rect 21150 1687 21185 1721
rect 21219 1687 21254 1721
rect 21288 1687 21323 1721
rect 21357 1687 21392 1721
rect 21426 1687 21461 1721
rect 21495 1687 21530 1721
rect 21564 1687 21599 1721
rect 21633 1687 21668 1721
rect 21702 1687 21737 1721
rect 21771 1687 21806 1721
rect 21840 1687 21875 1721
rect 21909 1687 21944 1721
rect 21978 1687 22013 1721
rect 22047 1687 22082 1721
rect 22116 1687 22151 1721
rect 22185 1687 22220 1721
rect 22254 1687 22289 1721
rect 22323 1687 22358 1721
rect 22392 1687 22427 1721
rect 22461 1687 22496 1721
rect 22530 1687 22565 1721
rect 22599 1687 22634 1721
rect 22668 1687 22703 1721
rect 22737 1687 22772 1721
rect 22806 1687 22841 1721
rect 22875 1687 22910 1721
rect 22944 1687 22979 1721
rect 23013 1687 23048 1721
rect 23082 1687 23117 1721
rect 23151 1687 23186 1721
rect 23220 1687 23255 1721
rect 23289 1687 23324 1721
rect 23358 1687 23393 1721
rect 23427 1687 23462 1721
rect 23496 1687 23531 1721
rect 23565 1687 23600 1721
rect 23634 1687 23669 1721
rect 23703 1687 23738 1721
rect 23772 1687 23796 1721
rect 19563 1653 23796 1687
rect 19563 1619 19598 1653
rect 19632 1619 19667 1653
rect 19701 1619 19736 1653
rect 19770 1619 19805 1653
rect 19839 1619 19874 1653
rect 19908 1619 19943 1653
rect 19977 1619 20012 1653
rect 20046 1619 20081 1653
rect 20115 1619 20150 1653
rect 20184 1619 20219 1653
rect 20253 1619 20288 1653
rect 20322 1619 20357 1653
rect 20391 1619 20426 1653
rect 20460 1619 20495 1653
rect 20529 1619 20564 1653
rect 20598 1619 20633 1653
rect 20667 1619 20702 1653
rect 20736 1619 20771 1653
rect 20805 1619 20840 1653
rect 20874 1619 20909 1653
rect 20943 1619 20978 1653
rect 21012 1619 21047 1653
rect 21081 1619 21116 1653
rect 21150 1619 21185 1653
rect 21219 1619 21254 1653
rect 21288 1619 21323 1653
rect 21357 1619 21392 1653
rect 21426 1619 21461 1653
rect 21495 1619 21530 1653
rect 21564 1619 21599 1653
rect 21633 1619 21668 1653
rect 21702 1619 21737 1653
rect 21771 1619 21806 1653
rect 21840 1619 21875 1653
rect 21909 1619 21944 1653
rect 21978 1619 22013 1653
rect 22047 1619 22082 1653
rect 22116 1619 22151 1653
rect 22185 1619 22220 1653
rect 22254 1619 22289 1653
rect 22323 1619 22358 1653
rect 22392 1619 22427 1653
rect 22461 1619 22496 1653
rect 22530 1619 22565 1653
rect 22599 1619 22634 1653
rect 22668 1619 22703 1653
rect 22737 1619 22772 1653
rect 22806 1619 22841 1653
rect 22875 1619 22910 1653
rect 22944 1619 22979 1653
rect 23013 1619 23048 1653
rect 23082 1619 23117 1653
rect 23151 1619 23186 1653
rect 23220 1619 23255 1653
rect 23289 1619 23324 1653
rect 23358 1619 23393 1653
rect 23427 1619 23462 1653
rect 23496 1619 23531 1653
rect 23565 1619 23600 1653
rect 23634 1619 23669 1653
rect 23703 1619 23738 1653
rect 23772 1619 23796 1653
rect 19563 1585 23796 1619
rect 19563 1551 19598 1585
rect 19632 1551 19667 1585
rect 19701 1551 19736 1585
rect 19770 1551 19805 1585
rect 19839 1551 19874 1585
rect 19908 1551 19943 1585
rect 19977 1551 20012 1585
rect 20046 1551 20081 1585
rect 20115 1551 20150 1585
rect 20184 1551 20219 1585
rect 20253 1551 20288 1585
rect 20322 1551 20357 1585
rect 20391 1551 20426 1585
rect 20460 1551 20495 1585
rect 20529 1551 20564 1585
rect 20598 1551 20633 1585
rect 20667 1551 20702 1585
rect 20736 1551 20771 1585
rect 20805 1551 20840 1585
rect 20874 1551 20909 1585
rect 20943 1551 20978 1585
rect 21012 1551 21047 1585
rect 21081 1551 21116 1585
rect 21150 1551 21185 1585
rect 21219 1551 21254 1585
rect 21288 1551 21323 1585
rect 21357 1551 21392 1585
rect 21426 1551 21461 1585
rect 21495 1551 21530 1585
rect 21564 1551 21599 1585
rect 21633 1551 21668 1585
rect 21702 1551 21737 1585
rect 21771 1551 21806 1585
rect 21840 1551 21875 1585
rect 21909 1551 21944 1585
rect 21978 1551 22013 1585
rect 22047 1551 22082 1585
rect 22116 1551 22151 1585
rect 22185 1551 22220 1585
rect 22254 1551 22289 1585
rect 22323 1551 22358 1585
rect 22392 1551 22427 1585
rect 22461 1551 22496 1585
rect 22530 1551 22565 1585
rect 22599 1551 22634 1585
rect 22668 1551 22703 1585
rect 22737 1551 22772 1585
rect 22806 1551 22841 1585
rect 22875 1551 22910 1585
rect 22944 1551 22979 1585
rect 23013 1551 23048 1585
rect 23082 1551 23117 1585
rect 23151 1551 23186 1585
rect 23220 1551 23255 1585
rect 23289 1551 23324 1585
rect 23358 1551 23393 1585
rect 23427 1551 23462 1585
rect 23496 1551 23531 1585
rect 23565 1551 23600 1585
rect 23634 1551 23669 1585
rect 23703 1551 23738 1585
rect 23772 1551 23796 1585
rect 19563 1517 23796 1551
rect 19563 1483 19598 1517
rect 19632 1483 19667 1517
rect 19701 1483 19736 1517
rect 19770 1483 19805 1517
rect 19839 1483 19874 1517
rect 19908 1483 19943 1517
rect 19977 1483 20012 1517
rect 20046 1483 20081 1517
rect 20115 1483 20150 1517
rect 20184 1483 20219 1517
rect 20253 1483 20288 1517
rect 20322 1483 20357 1517
rect 20391 1483 20426 1517
rect 20460 1483 20495 1517
rect 20529 1483 20564 1517
rect 20598 1483 20633 1517
rect 20667 1483 20702 1517
rect 20736 1483 20771 1517
rect 20805 1483 20840 1517
rect 20874 1483 20909 1517
rect 20943 1483 20978 1517
rect 21012 1483 21047 1517
rect 21081 1483 21116 1517
rect 21150 1483 21185 1517
rect 21219 1483 21254 1517
rect 21288 1483 21323 1517
rect 21357 1483 21392 1517
rect 21426 1483 21461 1517
rect 21495 1483 21530 1517
rect 21564 1483 21599 1517
rect 21633 1483 21668 1517
rect 21702 1483 21737 1517
rect 21771 1483 21806 1517
rect 21840 1483 21875 1517
rect 21909 1483 21944 1517
rect 21978 1483 22013 1517
rect 22047 1483 22082 1517
rect 22116 1483 22151 1517
rect 22185 1483 22220 1517
rect 22254 1483 22289 1517
rect 22323 1483 22358 1517
rect 22392 1483 22427 1517
rect 22461 1483 22496 1517
rect 22530 1483 22565 1517
rect 22599 1483 22634 1517
rect 22668 1483 22703 1517
rect 22737 1483 22772 1517
rect 22806 1483 22841 1517
rect 22875 1483 22910 1517
rect 22944 1483 22979 1517
rect 23013 1483 23048 1517
rect 23082 1483 23117 1517
rect 23151 1483 23186 1517
rect 23220 1483 23255 1517
rect 23289 1483 23324 1517
rect 23358 1483 23393 1517
rect 23427 1483 23462 1517
rect 23496 1483 23531 1517
rect 23565 1483 23600 1517
rect 23634 1483 23669 1517
rect 23703 1483 23738 1517
rect 23772 1483 23796 1517
rect 19563 1449 23796 1483
rect 19563 1415 19598 1449
rect 19632 1415 19667 1449
rect 19701 1415 19736 1449
rect 19770 1415 19805 1449
rect 19839 1415 19874 1449
rect 19908 1415 19943 1449
rect 19977 1415 20012 1449
rect 20046 1415 20081 1449
rect 20115 1415 20150 1449
rect 20184 1415 20219 1449
rect 20253 1415 20288 1449
rect 20322 1415 20357 1449
rect 20391 1415 20426 1449
rect 20460 1415 20495 1449
rect 20529 1415 20564 1449
rect 20598 1415 20633 1449
rect 20667 1415 20702 1449
rect 20736 1415 20771 1449
rect 20805 1415 20840 1449
rect 20874 1415 20909 1449
rect 20943 1415 20978 1449
rect 21012 1415 21047 1449
rect 21081 1415 21116 1449
rect 21150 1415 21185 1449
rect 21219 1415 21254 1449
rect 21288 1415 21323 1449
rect 21357 1415 21392 1449
rect 21426 1415 21461 1449
rect 21495 1415 21530 1449
rect 21564 1415 21599 1449
rect 21633 1415 21668 1449
rect 21702 1415 21737 1449
rect 21771 1415 21806 1449
rect 21840 1415 21875 1449
rect 21909 1415 21944 1449
rect 21978 1415 22013 1449
rect 22047 1415 22082 1449
rect 22116 1415 22151 1449
rect 22185 1415 22220 1449
rect 22254 1415 22289 1449
rect 22323 1415 22358 1449
rect 22392 1415 22427 1449
rect 22461 1415 22496 1449
rect 22530 1415 22565 1449
rect 22599 1415 22634 1449
rect 22668 1415 22703 1449
rect 22737 1415 22772 1449
rect 22806 1415 22841 1449
rect 22875 1415 22910 1449
rect 22944 1415 22979 1449
rect 23013 1415 23048 1449
rect 23082 1415 23117 1449
rect 23151 1415 23186 1449
rect 23220 1415 23255 1449
rect 23289 1415 23324 1449
rect 23358 1415 23393 1449
rect 23427 1415 23462 1449
rect 23496 1415 23531 1449
rect 23565 1415 23600 1449
rect 23634 1415 23669 1449
rect 23703 1415 23738 1449
rect 23772 1415 23796 1449
rect 19563 1381 23796 1415
rect 19563 1347 19598 1381
rect 19632 1347 19667 1381
rect 19701 1347 19736 1381
rect 19770 1347 19805 1381
rect 19839 1347 19874 1381
rect 19908 1347 19943 1381
rect 19977 1347 20012 1381
rect 20046 1347 20081 1381
rect 20115 1347 20150 1381
rect 20184 1347 20219 1381
rect 20253 1347 20288 1381
rect 20322 1347 20357 1381
rect 20391 1347 20426 1381
rect 20460 1347 20495 1381
rect 20529 1347 20564 1381
rect 20598 1347 20633 1381
rect 20667 1347 20702 1381
rect 20736 1347 20771 1381
rect 20805 1347 20840 1381
rect 20874 1347 20909 1381
rect 20943 1347 20978 1381
rect 21012 1347 21047 1381
rect 21081 1347 21116 1381
rect 21150 1347 21185 1381
rect 21219 1347 21254 1381
rect 21288 1347 21323 1381
rect 21357 1347 21392 1381
rect 21426 1347 21461 1381
rect 21495 1347 21530 1381
rect 21564 1347 21599 1381
rect 21633 1347 21668 1381
rect 21702 1347 21737 1381
rect 21771 1347 21806 1381
rect 21840 1347 21875 1381
rect 21909 1347 21944 1381
rect 21978 1347 22013 1381
rect 22047 1347 22082 1381
rect 22116 1347 22151 1381
rect 22185 1347 22220 1381
rect 22254 1347 22289 1381
rect 22323 1347 22358 1381
rect 22392 1347 22427 1381
rect 22461 1347 22496 1381
rect 22530 1347 22565 1381
rect 22599 1347 22634 1381
rect 22668 1347 22703 1381
rect 22737 1347 22772 1381
rect 22806 1347 22841 1381
rect 22875 1347 22910 1381
rect 22944 1347 22979 1381
rect 23013 1347 23048 1381
rect 23082 1347 23117 1381
rect 23151 1347 23186 1381
rect 23220 1347 23255 1381
rect 23289 1347 23324 1381
rect 23358 1347 23393 1381
rect 23427 1347 23462 1381
rect 23496 1347 23531 1381
rect 23565 1347 23600 1381
rect 23634 1347 23669 1381
rect 23703 1347 23738 1381
rect 23772 1347 23796 1381
rect 19563 1313 23796 1347
rect 19563 1279 19598 1313
rect 19632 1279 19667 1313
rect 19701 1279 19736 1313
rect 19770 1279 19805 1313
rect 19839 1279 19874 1313
rect 19908 1279 19943 1313
rect 19977 1279 20012 1313
rect 20046 1279 20081 1313
rect 20115 1279 20150 1313
rect 20184 1279 20219 1313
rect 20253 1279 20288 1313
rect 20322 1279 20357 1313
rect 20391 1279 20426 1313
rect 20460 1279 20495 1313
rect 20529 1279 20564 1313
rect 20598 1279 20633 1313
rect 20667 1279 20702 1313
rect 20736 1279 20771 1313
rect 20805 1279 20840 1313
rect 20874 1279 20909 1313
rect 20943 1279 20978 1313
rect 21012 1279 21047 1313
rect 21081 1279 21116 1313
rect 21150 1279 21185 1313
rect 21219 1279 21254 1313
rect 21288 1279 21323 1313
rect 21357 1279 21392 1313
rect 21426 1279 21461 1313
rect 21495 1279 21530 1313
rect 21564 1279 21599 1313
rect 21633 1279 21668 1313
rect 21702 1279 21737 1313
rect 21771 1279 21806 1313
rect 21840 1279 21875 1313
rect 21909 1279 21944 1313
rect 21978 1279 22013 1313
rect 22047 1279 22082 1313
rect 22116 1279 22151 1313
rect 22185 1279 22220 1313
rect 22254 1279 22289 1313
rect 22323 1279 22358 1313
rect 22392 1279 22427 1313
rect 22461 1279 22496 1313
rect 22530 1279 22565 1313
rect 22599 1279 22634 1313
rect 22668 1279 22703 1313
rect 22737 1279 22772 1313
rect 22806 1279 22841 1313
rect 22875 1279 22910 1313
rect 22944 1279 22979 1313
rect 23013 1279 23048 1313
rect 23082 1279 23117 1313
rect 23151 1279 23186 1313
rect 23220 1279 23255 1313
rect 23289 1279 23324 1313
rect 23358 1279 23393 1313
rect 23427 1279 23462 1313
rect 23496 1279 23531 1313
rect 23565 1279 23600 1313
rect 23634 1279 23669 1313
rect 23703 1279 23738 1313
rect 23772 1279 23796 1313
rect 19563 1245 23796 1279
rect 19563 1211 19598 1245
rect 19632 1211 19667 1245
rect 19701 1211 19736 1245
rect 19770 1211 19805 1245
rect 19839 1211 19874 1245
rect 19908 1211 19943 1245
rect 19977 1211 20012 1245
rect 20046 1211 20081 1245
rect 20115 1211 20150 1245
rect 20184 1211 20219 1245
rect 20253 1211 20288 1245
rect 20322 1211 20357 1245
rect 20391 1211 20426 1245
rect 20460 1211 20495 1245
rect 20529 1211 20564 1245
rect 20598 1211 20633 1245
rect 20667 1211 20702 1245
rect 20736 1211 20771 1245
rect 20805 1211 20840 1245
rect 20874 1211 20909 1245
rect 20943 1211 20978 1245
rect 21012 1211 21047 1245
rect 21081 1211 21116 1245
rect 21150 1211 21185 1245
rect 21219 1211 21254 1245
rect 21288 1211 21323 1245
rect 21357 1211 21392 1245
rect 21426 1211 21461 1245
rect 21495 1211 21530 1245
rect 21564 1211 21599 1245
rect 21633 1211 21668 1245
rect 21702 1211 21737 1245
rect 21771 1211 21806 1245
rect 21840 1211 21875 1245
rect 21909 1211 21944 1245
rect 21978 1211 22013 1245
rect 22047 1211 22082 1245
rect 22116 1211 22151 1245
rect 22185 1211 22220 1245
rect 22254 1211 22289 1245
rect 22323 1211 22358 1245
rect 22392 1211 22427 1245
rect 22461 1211 22496 1245
rect 22530 1211 22565 1245
rect 22599 1211 22634 1245
rect 22668 1211 22703 1245
rect 22737 1211 22772 1245
rect 22806 1211 22841 1245
rect 22875 1211 22910 1245
rect 22944 1211 22979 1245
rect 23013 1211 23048 1245
rect 23082 1211 23117 1245
rect 23151 1211 23186 1245
rect 23220 1211 23255 1245
rect 23289 1211 23324 1245
rect 23358 1211 23393 1245
rect 23427 1211 23462 1245
rect 23496 1211 23531 1245
rect 23565 1211 23600 1245
rect 23634 1211 23669 1245
rect 23703 1211 23738 1245
rect 23772 1211 23796 1245
rect 19563 1177 23796 1211
rect 19563 1143 19598 1177
rect 19632 1143 19667 1177
rect 19701 1143 19736 1177
rect 19770 1143 19805 1177
rect 19839 1143 19874 1177
rect 19908 1143 19943 1177
rect 19977 1143 20012 1177
rect 20046 1143 20081 1177
rect 20115 1143 20150 1177
rect 20184 1143 20219 1177
rect 20253 1143 20288 1177
rect 20322 1143 20357 1177
rect 20391 1143 20426 1177
rect 20460 1143 20495 1177
rect 20529 1143 20564 1177
rect 20598 1143 20633 1177
rect 20667 1143 20702 1177
rect 20736 1143 20771 1177
rect 20805 1143 20840 1177
rect 20874 1143 20909 1177
rect 20943 1143 20978 1177
rect 21012 1143 21047 1177
rect 21081 1143 21116 1177
rect 21150 1143 21185 1177
rect 21219 1143 21254 1177
rect 21288 1143 21323 1177
rect 21357 1143 21392 1177
rect 21426 1143 21461 1177
rect 21495 1143 21530 1177
rect 21564 1143 21599 1177
rect 21633 1143 21668 1177
rect 21702 1143 21737 1177
rect 21771 1143 21806 1177
rect 21840 1143 21875 1177
rect 21909 1143 21944 1177
rect 21978 1143 22013 1177
rect 22047 1143 22082 1177
rect 22116 1143 22151 1177
rect 22185 1143 22220 1177
rect 22254 1143 22289 1177
rect 22323 1143 22358 1177
rect 22392 1143 22427 1177
rect 22461 1143 22496 1177
rect 22530 1143 22565 1177
rect 22599 1143 22634 1177
rect 22668 1143 22703 1177
rect 22737 1143 22772 1177
rect 22806 1143 22841 1177
rect 22875 1143 22910 1177
rect 22944 1143 22979 1177
rect 23013 1143 23048 1177
rect 23082 1143 23117 1177
rect 23151 1143 23186 1177
rect 23220 1143 23255 1177
rect 23289 1143 23324 1177
rect 23358 1143 23393 1177
rect 23427 1143 23462 1177
rect 23496 1143 23531 1177
rect 23565 1143 23600 1177
rect 23634 1143 23669 1177
rect 23703 1143 23738 1177
rect 23772 1143 23796 1177
rect 14625 1128 23796 1143
rect 14397 1109 14625 1112
rect 14397 1091 14455 1109
rect 730 1040 764 1074
rect 696 1005 764 1040
rect 730 1003 764 1005
rect 866 1075 14455 1091
rect 14489 1075 14523 1109
rect 14557 1076 14625 1109
rect 14557 1075 14591 1076
rect 866 1042 14591 1075
rect 866 1039 14625 1042
rect 866 1037 14523 1039
rect 866 1003 901 1037
rect 935 1003 970 1037
rect 1004 1003 1039 1037
rect 1073 1003 1108 1037
rect 1142 1003 1177 1037
rect 1211 1003 1246 1037
rect 1280 1003 1315 1037
rect 1349 1003 1384 1037
rect 1418 1003 1453 1037
rect 1487 1003 1522 1037
rect 1556 1003 1591 1037
rect 1625 1003 1660 1037
rect 1694 1003 1729 1037
rect 1763 1003 1798 1037
rect 1832 1003 1867 1037
rect 1901 1003 1936 1037
rect 1970 1003 2005 1037
rect 2039 1003 2074 1037
rect 2108 1003 2143 1037
rect 2177 1003 2212 1037
rect 2246 1003 2281 1037
rect 2315 1003 2350 1037
rect 2384 1003 2419 1037
rect 730 971 2419 1003
rect 696 969 2419 971
rect 14489 1005 14523 1037
rect 14557 1006 14625 1039
rect 14557 1005 14591 1006
rect 14489 972 14591 1005
rect 14489 969 14625 972
rect 696 935 764 969
rect 798 935 833 969
rect 867 935 902 969
rect 936 935 971 969
rect 1005 935 1040 969
rect 1074 935 1109 969
rect 1143 935 1178 969
rect 1212 935 1247 969
rect 1281 935 1316 969
rect 1350 935 1385 969
rect 1419 935 1454 969
rect 1488 935 1523 969
rect 1557 935 1592 969
rect 1626 935 1661 969
rect 1695 935 1730 969
rect 1764 935 1799 969
rect 1833 935 1868 969
rect 1902 935 1937 969
rect 1971 935 2006 969
rect 2040 935 2075 969
rect 2109 935 2144 969
rect 2178 935 2213 969
rect 2247 935 2282 969
rect 2316 935 2351 969
rect 14557 935 14625 969
rect 696 901 2351 935
rect 14523 901 14591 935
rect 696 867 730 901
rect 764 867 799 901
rect 833 867 868 901
rect 902 867 937 901
rect 971 867 1006 901
rect 1040 867 1075 901
rect 1109 867 1144 901
rect 1178 867 1213 901
rect 1247 867 1282 901
rect 1316 867 1351 901
rect 1385 867 1420 901
rect 1454 867 1489 901
rect 1523 867 1558 901
rect 1592 867 1627 901
rect 1661 867 1696 901
rect 1730 867 1765 901
rect 1799 867 1834 901
rect 1868 867 1903 901
rect 1937 867 1972 901
rect 2006 867 2041 901
rect 2075 867 2110 901
rect 2144 867 2179 901
rect 2213 867 2248 901
rect 2282 867 2317 901
rect 14523 867 14625 901
<< mvnsubdiff >>
rect 24370 9395 24540 9419
rect 24370 9121 24540 9157
rect 24404 9087 24438 9121
rect 24472 9087 24506 9121
rect 24370 9051 24540 9087
rect 24404 9017 24438 9051
rect 24472 9017 24506 9051
rect 24370 8981 24540 9017
rect 24404 8947 24438 8981
rect 24472 8947 24506 8981
rect 24370 8912 24540 8947
rect 24404 8878 24438 8912
rect 24472 8878 24506 8912
rect 24370 8843 24540 8878
rect 24404 8809 24438 8843
rect 24472 8809 24506 8843
rect 24370 8774 24540 8809
rect 24404 8740 24438 8774
rect 24472 8740 24506 8774
rect 24370 8705 24540 8740
rect 24404 8671 24438 8705
rect 24472 8671 24506 8705
rect 24370 8636 24540 8671
rect 23752 8568 24370 8592
rect 23752 8534 23755 8568
rect 23789 8534 23823 8568
rect 23857 8534 23891 8568
rect 23925 8534 23959 8568
rect 23993 8534 24027 8568
rect 24061 8534 24095 8568
rect 24129 8534 24163 8568
rect 24197 8534 24231 8568
rect 24265 8534 24299 8568
rect 24333 8534 24367 8568
rect 24537 8534 24540 8602
rect 23752 8499 24540 8534
rect 23752 8465 23755 8499
rect 23789 8465 23823 8499
rect 23857 8465 23891 8499
rect 23925 8465 23959 8499
rect 23993 8465 24027 8499
rect 24061 8465 24095 8499
rect 24129 8465 24163 8499
rect 24197 8465 24231 8499
rect 24265 8465 24299 8499
rect 24333 8465 24367 8499
rect 24401 8465 24435 8499
rect 24469 8465 24503 8499
rect 24537 8465 24540 8499
rect 23752 8430 24540 8465
rect 23752 8396 23755 8430
rect 23789 8396 23823 8430
rect 23857 8396 23891 8430
rect 23925 8396 23959 8430
rect 23993 8396 24027 8430
rect 24061 8396 24095 8430
rect 24129 8396 24163 8430
rect 24197 8396 24231 8430
rect 24265 8396 24299 8430
rect 24333 8396 24367 8430
rect 24401 8396 24435 8430
rect 24469 8396 24503 8430
rect 24537 8396 24540 8430
rect 23752 8361 24540 8396
rect 23752 8327 23755 8361
rect 23789 8327 23823 8361
rect 23857 8327 23891 8361
rect 23925 8327 23959 8361
rect 23993 8327 24027 8361
rect 24061 8327 24095 8361
rect 24129 8327 24163 8361
rect 24197 8327 24231 8361
rect 24265 8327 24299 8361
rect 24333 8327 24367 8361
rect 24401 8327 24435 8361
rect 24469 8327 24503 8361
rect 24537 8327 24540 8361
rect 23752 8292 24540 8327
rect 23752 8258 23755 8292
rect 23789 8258 23823 8292
rect 23857 8258 23891 8292
rect 23925 8258 23959 8292
rect 23993 8258 24027 8292
rect 24061 8258 24095 8292
rect 24129 8258 24163 8292
rect 24197 8258 24231 8292
rect 24265 8258 24299 8292
rect 24333 8258 24367 8292
rect 24401 8258 24435 8292
rect 24469 8258 24503 8292
rect 24537 8258 24540 8292
rect 23752 8223 24540 8258
rect 23752 8189 23755 8223
rect 23789 8189 23823 8223
rect 23857 8189 23891 8223
rect 23925 8189 23959 8223
rect 23993 8189 24027 8223
rect 24061 8189 24095 8223
rect 24129 8189 24163 8223
rect 24197 8189 24231 8223
rect 24265 8189 24299 8223
rect 24333 8189 24367 8223
rect 24401 8189 24435 8223
rect 24469 8189 24503 8223
rect 24537 8189 24540 8223
rect 23752 8154 24540 8189
rect 23752 8120 23755 8154
rect 23789 8120 23823 8154
rect 23857 8120 23891 8154
rect 23925 8120 23959 8154
rect 23993 8120 24027 8154
rect 24061 8120 24095 8154
rect 24129 8120 24163 8154
rect 24197 8120 24231 8154
rect 24265 8120 24299 8154
rect 24333 8120 24367 8154
rect 24401 8120 24435 8154
rect 24469 8120 24503 8154
rect 24537 8120 24540 8154
rect 23752 8085 24540 8120
rect 23752 8051 23755 8085
rect 23789 8051 23823 8085
rect 23857 8051 23891 8085
rect 23925 8051 23959 8085
rect 23993 8051 24027 8085
rect 24061 8051 24095 8085
rect 24129 8051 24163 8085
rect 24197 8051 24231 8085
rect 24265 8051 24299 8085
rect 24333 8051 24367 8085
rect 24401 8051 24435 8085
rect 24469 8051 24503 8085
rect 24537 8051 24540 8085
rect 23752 8016 24540 8051
rect 23752 7982 23755 8016
rect 23789 7982 23823 8016
rect 23857 7982 23891 8016
rect 23925 7982 23959 8016
rect 23993 7982 24027 8016
rect 24061 7982 24095 8016
rect 24129 7982 24163 8016
rect 24197 7982 24231 8016
rect 24265 7982 24299 8016
rect 24333 7982 24367 8016
rect 24401 7982 24435 8016
rect 24469 7982 24503 8016
rect 24537 7982 24540 8016
rect 23752 7947 24540 7982
rect 23752 7913 23755 7947
rect 23789 7913 23823 7947
rect 23857 7913 23891 7947
rect 23925 7913 23959 7947
rect 23993 7913 24027 7947
rect 24061 7913 24095 7947
rect 24129 7913 24163 7947
rect 24197 7913 24231 7947
rect 24265 7913 24299 7947
rect 24333 7913 24367 7947
rect 24401 7913 24435 7947
rect 24469 7913 24503 7947
rect 24537 7913 24540 7947
rect 23752 7878 24540 7913
rect 23752 7844 23755 7878
rect 23789 7844 23823 7878
rect 23857 7844 23891 7878
rect 23925 7844 23959 7878
rect 23993 7844 24027 7878
rect 24061 7844 24095 7878
rect 24129 7844 24163 7878
rect 24197 7844 24231 7878
rect 24265 7844 24299 7878
rect 24333 7844 24367 7878
rect 24401 7844 24435 7878
rect 24469 7844 24503 7878
rect 24537 7844 24540 7878
rect 23752 7809 24540 7844
rect 23752 7775 23755 7809
rect 23789 7775 23823 7809
rect 23857 7775 23891 7809
rect 23925 7775 23959 7809
rect 23993 7775 24027 7809
rect 24061 7775 24095 7809
rect 24129 7775 24163 7809
rect 24197 7775 24231 7809
rect 24265 7775 24299 7809
rect 24333 7775 24367 7809
rect 24401 7775 24435 7809
rect 24469 7775 24503 7809
rect 24537 7775 24540 7809
rect 23752 7740 24540 7775
rect 23752 7706 23755 7740
rect 23789 7706 23823 7740
rect 23857 7706 23891 7740
rect 23925 7706 23959 7740
rect 23993 7706 24027 7740
rect 24061 7706 24095 7740
rect 24129 7706 24163 7740
rect 24197 7706 24231 7740
rect 24265 7706 24299 7740
rect 24333 7706 24367 7740
rect 24401 7706 24435 7740
rect 24469 7706 24503 7740
rect 24537 7706 24540 7740
rect 23752 7671 24540 7706
rect 23752 7637 23755 7671
rect 23789 7637 23823 7671
rect 23857 7637 23891 7671
rect 23925 7637 23959 7671
rect 23993 7637 24027 7671
rect 24061 7637 24095 7671
rect 24129 7637 24163 7671
rect 24197 7637 24231 7671
rect 24265 7637 24299 7671
rect 24333 7637 24367 7671
rect 24401 7637 24435 7671
rect 24469 7637 24503 7671
rect 24537 7637 24540 7671
rect 23752 7602 24540 7637
rect 23752 7568 23755 7602
rect 23789 7568 23823 7602
rect 23857 7568 23891 7602
rect 23925 7568 23959 7602
rect 23993 7568 24027 7602
rect 24061 7568 24095 7602
rect 24129 7568 24163 7602
rect 24197 7568 24231 7602
rect 24265 7568 24299 7602
rect 24333 7568 24367 7602
rect 24401 7568 24435 7602
rect 24469 7568 24503 7602
rect 24537 7568 24540 7602
rect 23752 7533 24540 7568
rect 23752 7499 23755 7533
rect 23789 7499 23823 7533
rect 23857 7499 23891 7533
rect 23925 7499 23959 7533
rect 23993 7499 24027 7533
rect 24061 7499 24095 7533
rect 24129 7499 24163 7533
rect 24197 7499 24231 7533
rect 24265 7499 24299 7533
rect 24333 7499 24367 7533
rect 24401 7499 24435 7533
rect 24469 7499 24503 7533
rect 24537 7499 24540 7533
rect 23752 7464 24540 7499
rect 23752 7430 23755 7464
rect 23789 7430 23823 7464
rect 23857 7430 23891 7464
rect 23925 7430 23959 7464
rect 23993 7430 24027 7464
rect 24061 7430 24095 7464
rect 24129 7430 24163 7464
rect 24197 7430 24231 7464
rect 24265 7430 24299 7464
rect 24333 7430 24367 7464
rect 24401 7430 24435 7464
rect 24469 7430 24503 7464
rect 24537 7430 24540 7464
rect 23752 7395 24540 7430
rect 23752 7361 23755 7395
rect 23789 7361 23823 7395
rect 23857 7361 23891 7395
rect 23925 7361 23959 7395
rect 23993 7361 24027 7395
rect 24061 7361 24095 7395
rect 24129 7361 24163 7395
rect 24197 7361 24231 7395
rect 24265 7361 24299 7395
rect 24333 7361 24367 7395
rect 24401 7361 24435 7395
rect 24469 7361 24503 7395
rect 24537 7361 24540 7395
rect 23752 7326 24540 7361
rect 23752 7292 23755 7326
rect 23789 7292 23823 7326
rect 23857 7292 23891 7326
rect 23925 7292 23959 7326
rect 23993 7292 24027 7326
rect 24061 7292 24095 7326
rect 24129 7292 24163 7326
rect 24197 7292 24231 7326
rect 24265 7292 24299 7326
rect 24333 7292 24367 7326
rect 24401 7292 24435 7326
rect 24469 7292 24503 7326
rect 24537 7292 24540 7326
rect 23752 7257 24540 7292
rect 23752 7223 23755 7257
rect 23789 7223 23823 7257
rect 23857 7223 23891 7257
rect 23925 7223 23959 7257
rect 23993 7223 24027 7257
rect 24061 7223 24095 7257
rect 24129 7223 24163 7257
rect 24197 7223 24231 7257
rect 24265 7223 24299 7257
rect 24333 7223 24367 7257
rect 24401 7223 24435 7257
rect 24469 7223 24503 7257
rect 24537 7223 24540 7257
rect 23752 7188 24540 7223
rect 23752 7154 23755 7188
rect 23789 7154 23823 7188
rect 23857 7154 23891 7188
rect 23925 7154 23959 7188
rect 23993 7154 24027 7188
rect 24061 7154 24095 7188
rect 24129 7154 24163 7188
rect 24197 7154 24231 7188
rect 24265 7154 24299 7188
rect 24333 7154 24367 7188
rect 24401 7154 24435 7188
rect 24469 7154 24503 7188
rect 24537 7154 24540 7188
rect 23752 7119 24540 7154
rect 23752 7085 23755 7119
rect 23789 7085 23823 7119
rect 23857 7085 23891 7119
rect 23925 7085 23959 7119
rect 23993 7085 24027 7119
rect 24061 7085 24095 7119
rect 24129 7085 24163 7119
rect 24197 7085 24231 7119
rect 24265 7085 24299 7119
rect 24333 7085 24367 7119
rect 24401 7085 24435 7119
rect 24469 7085 24503 7119
rect 24537 7085 24540 7119
rect 23752 7050 24540 7085
rect 23752 7016 23755 7050
rect 23789 7016 23823 7050
rect 23857 7016 23891 7050
rect 23925 7016 23959 7050
rect 23993 7016 24027 7050
rect 24061 7016 24095 7050
rect 24129 7016 24163 7050
rect 24197 7016 24231 7050
rect 24265 7016 24299 7050
rect 24333 7016 24367 7050
rect 24401 7016 24435 7050
rect 24469 7016 24503 7050
rect 24537 7016 24540 7050
rect 23752 6981 24540 7016
rect 23752 6947 23755 6981
rect 23789 6947 23823 6981
rect 23857 6947 23891 6981
rect 23925 6947 23959 6981
rect 23993 6947 24027 6981
rect 24061 6947 24095 6981
rect 24129 6947 24163 6981
rect 24197 6947 24231 6981
rect 24265 6947 24299 6981
rect 24333 6947 24367 6981
rect 24401 6947 24435 6981
rect 24469 6947 24503 6981
rect 24537 6947 24540 6981
rect 23752 6912 24540 6947
rect 23752 6878 23755 6912
rect 23789 6878 23823 6912
rect 23857 6878 23891 6912
rect 23925 6878 23959 6912
rect 23993 6878 24027 6912
rect 24061 6878 24095 6912
rect 24129 6878 24163 6912
rect 24197 6878 24231 6912
rect 24265 6878 24299 6912
rect 24333 6878 24367 6912
rect 24401 6878 24435 6912
rect 24469 6878 24503 6912
rect 24537 6878 24540 6912
rect 23752 6843 24540 6878
rect 23752 6809 23755 6843
rect 23789 6809 23823 6843
rect 23857 6809 23891 6843
rect 23925 6809 23959 6843
rect 23993 6809 24027 6843
rect 24061 6809 24095 6843
rect 24129 6809 24163 6843
rect 24197 6809 24231 6843
rect 24265 6809 24299 6843
rect 24333 6809 24367 6843
rect 24401 6809 24435 6843
rect 24469 6809 24503 6843
rect 24537 6809 24540 6843
rect 23752 6774 24540 6809
rect 23752 6740 23755 6774
rect 23789 6740 23823 6774
rect 23857 6740 23891 6774
rect 23925 6740 23959 6774
rect 23993 6740 24027 6774
rect 24061 6740 24095 6774
rect 24129 6740 24163 6774
rect 24197 6740 24231 6774
rect 24265 6740 24299 6774
rect 24333 6740 24367 6774
rect 24401 6740 24435 6774
rect 24469 6740 24503 6774
rect 24537 6740 24540 6774
rect 23752 6705 24540 6740
rect 23752 6671 23755 6705
rect 23789 6671 23823 6705
rect 23857 6671 23891 6705
rect 23925 6671 23959 6705
rect 23993 6671 24027 6705
rect 24061 6671 24095 6705
rect 24129 6671 24163 6705
rect 24197 6671 24231 6705
rect 24265 6671 24299 6705
rect 24333 6671 24367 6705
rect 24401 6671 24435 6705
rect 24469 6671 24503 6705
rect 24537 6671 24540 6705
rect 23752 6636 24540 6671
rect 23752 6602 23755 6636
rect 23789 6602 23823 6636
rect 23857 6602 23891 6636
rect 23925 6602 23959 6636
rect 23993 6602 24027 6636
rect 24061 6602 24095 6636
rect 24129 6602 24163 6636
rect 24197 6602 24231 6636
rect 24265 6602 24299 6636
rect 24333 6602 24367 6636
rect 24401 6602 24435 6636
rect 24469 6602 24503 6636
rect 24537 6602 24540 6636
rect 23752 6567 24540 6602
rect 23752 6533 23755 6567
rect 23789 6533 23823 6567
rect 23857 6533 23891 6567
rect 23925 6533 23959 6567
rect 23993 6533 24027 6567
rect 24061 6533 24095 6567
rect 24129 6533 24163 6567
rect 24197 6533 24231 6567
rect 24265 6533 24299 6567
rect 24333 6533 24367 6567
rect 24401 6533 24435 6567
rect 24469 6533 24503 6567
rect 24537 6533 24540 6567
rect 23752 6498 24540 6533
rect 23752 6464 23755 6498
rect 23789 6464 23823 6498
rect 23857 6464 23891 6498
rect 23925 6464 23959 6498
rect 23993 6464 24027 6498
rect 24061 6464 24095 6498
rect 24129 6464 24163 6498
rect 24197 6464 24231 6498
rect 24265 6464 24299 6498
rect 24333 6464 24367 6498
rect 24401 6464 24435 6498
rect 24469 6464 24503 6498
rect 24537 6464 24540 6498
rect 23752 6429 24540 6464
rect 23752 6395 23755 6429
rect 23789 6395 23823 6429
rect 23857 6395 23891 6429
rect 23925 6395 23959 6429
rect 23993 6395 24027 6429
rect 24061 6395 24095 6429
rect 24129 6395 24163 6429
rect 24197 6395 24231 6429
rect 24265 6395 24299 6429
rect 24333 6395 24367 6429
rect 24401 6395 24435 6429
rect 24469 6395 24503 6429
rect 24537 6395 24540 6429
rect 23752 6360 24540 6395
rect 23752 6326 23755 6360
rect 23789 6326 23823 6360
rect 23857 6326 23891 6360
rect 23925 6326 23959 6360
rect 23993 6326 24027 6360
rect 24061 6326 24095 6360
rect 24129 6326 24163 6360
rect 24197 6326 24231 6360
rect 24265 6326 24299 6360
rect 24333 6326 24367 6360
rect 24401 6326 24435 6360
rect 24469 6326 24503 6360
rect 24537 6326 24540 6360
rect 23752 6291 24540 6326
rect 23752 6257 23755 6291
rect 23789 6257 23823 6291
rect 23857 6257 23891 6291
rect 23925 6257 23959 6291
rect 23993 6257 24027 6291
rect 24061 6257 24095 6291
rect 24129 6257 24163 6291
rect 24197 6257 24231 6291
rect 24265 6257 24299 6291
rect 24333 6257 24367 6291
rect 24401 6257 24435 6291
rect 24469 6257 24503 6291
rect 24537 6257 24540 6291
rect 23752 6222 24540 6257
rect 23752 6188 23755 6222
rect 23789 6188 23823 6222
rect 23857 6188 23891 6222
rect 23925 6188 23959 6222
rect 23993 6188 24027 6222
rect 24061 6188 24095 6222
rect 24129 6188 24163 6222
rect 24197 6188 24231 6222
rect 24265 6188 24299 6222
rect 24333 6188 24367 6222
rect 24401 6188 24435 6222
rect 24469 6188 24503 6222
rect 24537 6188 24540 6222
rect 23752 6153 24540 6188
rect 23752 6119 23755 6153
rect 23789 6119 23823 6153
rect 23857 6119 23891 6153
rect 23925 6119 23959 6153
rect 23993 6119 24027 6153
rect 24061 6119 24095 6153
rect 24129 6119 24163 6153
rect 24197 6119 24231 6153
rect 24265 6119 24299 6153
rect 24333 6119 24367 6153
rect 24401 6119 24435 6153
rect 24469 6119 24503 6153
rect 24537 6119 24540 6153
rect 23752 6084 24540 6119
rect 23752 6050 23755 6084
rect 23789 6050 23823 6084
rect 23857 6050 23891 6084
rect 23925 6050 23959 6084
rect 23993 6050 24027 6084
rect 24061 6050 24095 6084
rect 24129 6050 24163 6084
rect 24197 6050 24231 6084
rect 24265 6050 24299 6084
rect 24333 6050 24367 6084
rect 24401 6050 24435 6084
rect 24469 6050 24503 6084
rect 24537 6050 24540 6084
rect 23752 6015 24540 6050
rect 23752 5981 23755 6015
rect 23789 5981 23823 6015
rect 23857 5981 23891 6015
rect 23925 5981 23959 6015
rect 23993 5981 24027 6015
rect 24061 5981 24095 6015
rect 24129 5981 24163 6015
rect 24197 5981 24231 6015
rect 24265 5981 24299 6015
rect 24333 5981 24367 6015
rect 24401 5981 24435 6015
rect 24469 5981 24503 6015
rect 24537 5981 24540 6015
rect 23752 5946 24540 5981
rect 23752 5912 23755 5946
rect 23789 5912 23823 5946
rect 23857 5912 23891 5946
rect 23925 5912 23959 5946
rect 23993 5912 24027 5946
rect 24061 5912 24095 5946
rect 24129 5912 24163 5946
rect 24197 5912 24231 5946
rect 24265 5912 24299 5946
rect 24333 5912 24367 5946
rect 24401 5912 24435 5946
rect 24469 5912 24503 5946
rect 24537 5912 24540 5946
rect 23752 5877 24540 5912
rect 23752 5639 23755 5877
rect 24537 5639 24540 5877
rect 23752 5615 24540 5639
rect 23949 5591 24540 5615
rect 23949 5557 24153 5591
rect 24187 5557 24221 5591
rect 24255 5557 24289 5591
rect 24323 5557 24357 5591
rect 24391 5557 24425 5591
rect 24459 5557 24493 5591
rect 24527 5557 24540 5591
rect 23949 5532 24540 5557
rect 278 4483 448 4517
rect 312 4449 346 4483
rect 380 4449 414 4483
rect 278 4413 448 4449
rect 312 4379 346 4413
rect 380 4379 414 4413
rect 278 4343 448 4379
rect 312 4309 346 4343
rect 380 4309 414 4343
rect 278 4273 448 4309
rect 312 4239 346 4273
rect 380 4239 414 4273
rect 278 4203 448 4239
rect 312 4169 346 4203
rect 380 4169 414 4203
rect 278 4134 448 4169
rect 312 4100 346 4134
rect 380 4100 414 4134
rect 278 4065 448 4100
rect 312 4031 346 4065
rect 380 4031 414 4065
rect 278 3996 448 4031
rect 312 3962 346 3996
rect 380 3962 414 3996
rect 278 3927 448 3962
rect 312 3893 346 3927
rect 380 3893 414 3927
rect 278 3858 448 3893
rect 312 3824 346 3858
rect 380 3824 414 3858
rect 278 3789 448 3824
rect 312 3755 346 3789
rect 380 3755 414 3789
rect 278 3720 448 3755
rect 312 3686 346 3720
rect 380 3686 414 3720
rect 278 3651 448 3686
rect 312 3617 346 3651
rect 380 3617 414 3651
rect 278 3582 448 3617
rect 312 3548 346 3582
rect 380 3548 414 3582
rect 278 3513 448 3548
rect 312 3479 346 3513
rect 380 3479 414 3513
rect 278 3444 448 3479
rect 312 3410 346 3444
rect 380 3410 414 3444
rect 278 3375 448 3410
rect 312 3341 346 3375
rect 380 3341 414 3375
rect 278 3306 448 3341
rect 312 3272 346 3306
rect 380 3272 414 3306
rect 278 3237 448 3272
rect 312 3203 346 3237
rect 380 3203 414 3237
rect 278 3168 448 3203
rect 312 3134 346 3168
rect 380 3134 414 3168
rect 278 3099 448 3134
rect 312 3065 346 3099
rect 380 3065 414 3099
rect 278 3030 448 3065
rect 312 2996 346 3030
rect 380 2996 414 3030
rect 278 2961 448 2996
rect 312 2927 346 2961
rect 380 2927 414 2961
rect 278 2892 448 2927
rect 312 2858 346 2892
rect 380 2858 414 2892
rect 278 2823 448 2858
rect 312 2789 346 2823
rect 380 2789 414 2823
rect 278 2754 448 2789
rect 312 2720 346 2754
rect 380 2720 414 2754
rect 278 2685 448 2720
rect 312 2651 346 2685
rect 380 2651 414 2685
rect 278 2616 448 2651
rect 312 2582 346 2616
rect 380 2582 414 2616
rect 278 2547 448 2582
rect 312 2513 346 2547
rect 380 2513 414 2547
rect 278 2478 448 2513
rect 312 2444 346 2478
rect 380 2444 414 2478
rect 278 2409 448 2444
rect 312 2375 346 2409
rect 380 2375 414 2409
rect 278 2340 448 2375
rect 312 2306 346 2340
rect 380 2306 414 2340
rect 278 2271 448 2306
rect 312 2237 346 2271
rect 380 2237 414 2271
rect 278 2202 448 2237
rect 312 2168 346 2202
rect 380 2168 414 2202
rect 278 2133 448 2168
rect 312 2099 346 2133
rect 380 2099 414 2133
rect 278 2064 448 2099
rect 312 2030 346 2064
rect 380 2030 414 2064
rect 278 1995 448 2030
rect 312 1961 346 1995
rect 380 1961 414 1995
rect 278 1926 448 1961
rect 312 1892 346 1926
rect 380 1892 414 1926
rect 278 1857 448 1892
rect 312 1823 346 1857
rect 380 1823 414 1857
rect 278 1788 448 1823
rect 312 1754 346 1788
rect 380 1754 414 1788
rect 278 1719 448 1754
rect 312 1685 346 1719
rect 380 1685 414 1719
rect 278 1650 448 1685
rect 312 1616 346 1650
rect 380 1616 414 1650
rect 278 1581 448 1616
rect 312 1547 346 1581
rect 380 1547 414 1581
rect 278 1512 448 1547
rect 312 1478 346 1512
rect 380 1478 414 1512
rect 278 1443 448 1478
rect 312 1409 346 1443
rect 380 1409 414 1443
rect 278 1374 448 1409
rect 312 1340 346 1374
rect 380 1340 414 1374
rect 278 1305 448 1340
rect 312 1271 346 1305
rect 380 1271 414 1305
rect 278 1236 448 1271
rect 312 1202 346 1236
rect 380 1202 414 1236
rect 278 1167 448 1202
rect 312 1133 346 1167
rect 380 1133 414 1167
rect 278 1098 448 1133
rect 312 1064 346 1098
rect 380 1064 414 1098
rect 278 1029 448 1064
rect 312 995 346 1029
rect 380 995 414 1029
rect 278 960 448 995
rect 312 926 346 960
rect 380 926 414 960
rect 278 891 448 926
rect 312 857 346 891
rect 380 857 414 891
rect 1086 4550 1609 4574
rect 1120 4516 1154 4550
rect 1188 4516 1222 4550
rect 1256 4516 1290 4550
rect 1324 4516 1358 4550
rect 1392 4516 1426 4550
rect 1460 4540 1609 4550
rect 1460 4516 1507 4540
rect 1086 4506 1507 4516
rect 1541 4506 1609 4540
rect 6335 4540 6370 4574
rect 6404 4540 6439 4574
rect 6473 4540 6508 4574
rect 6542 4540 6577 4574
rect 6611 4540 6646 4574
rect 6680 4540 6715 4574
rect 6749 4540 6784 4574
rect 6818 4540 6853 4574
rect 6887 4540 6922 4574
rect 6956 4540 6991 4574
rect 7025 4540 7060 4574
rect 7094 4540 7129 4574
rect 7163 4540 7198 4574
rect 7232 4540 7267 4574
rect 7301 4540 7336 4574
rect 7370 4540 7405 4574
rect 7439 4540 7474 4574
rect 7508 4540 7543 4574
rect 7577 4540 7612 4574
rect 7646 4540 7681 4574
rect 7715 4540 7750 4574
rect 7784 4540 7819 4574
rect 7853 4540 7888 4574
rect 7922 4540 7957 4574
rect 7991 4540 8026 4574
rect 8060 4540 8095 4574
rect 8129 4540 8164 4574
rect 8198 4540 8233 4574
rect 8267 4540 8302 4574
rect 8336 4540 8371 4574
rect 8405 4540 8440 4574
rect 8474 4540 8509 4574
rect 8543 4540 8578 4574
rect 8612 4540 8647 4574
rect 8681 4540 8716 4574
rect 8750 4540 8785 4574
rect 8819 4540 8854 4574
rect 8888 4540 8923 4574
rect 8957 4540 8992 4574
rect 9026 4540 9061 4574
rect 9095 4540 9130 4574
rect 9164 4540 9199 4574
rect 9233 4540 9268 4574
rect 9302 4540 9337 4574
rect 9371 4540 9406 4574
rect 9440 4540 9475 4574
rect 9509 4540 9544 4574
rect 9578 4540 9613 4574
rect 9647 4540 9682 4574
rect 9716 4540 9751 4574
rect 9785 4540 9820 4574
rect 9854 4540 9889 4574
rect 9923 4540 9958 4574
rect 9992 4540 10026 4574
rect 6335 4506 10026 4540
rect 1086 4481 1575 4506
rect 1120 4447 1154 4481
rect 1188 4447 1222 4481
rect 1256 4447 1290 4481
rect 1324 4447 1358 4481
rect 1392 4447 1426 4481
rect 1460 4472 1575 4481
rect 8681 4472 8716 4506
rect 8750 4472 8785 4506
rect 8819 4472 8854 4506
rect 8888 4472 8923 4506
rect 8957 4472 8992 4506
rect 9026 4472 9061 4506
rect 9095 4472 9130 4506
rect 9164 4472 9199 4506
rect 9233 4472 9268 4506
rect 9302 4472 9337 4506
rect 9371 4472 9406 4506
rect 9440 4472 9475 4506
rect 9509 4472 9544 4506
rect 9578 4472 9613 4506
rect 9647 4472 9682 4506
rect 9716 4472 9751 4506
rect 9785 4472 9820 4506
rect 9854 4472 9889 4506
rect 9923 4472 9958 4506
rect 9992 4472 10026 4506
rect 1460 4471 1643 4472
rect 1460 4447 1507 4471
rect 1086 4437 1507 4447
rect 1541 4437 1643 4471
rect 1086 4436 1643 4437
rect 1086 4412 1575 4436
rect 1120 4378 1154 4412
rect 1188 4378 1222 4412
rect 1256 4378 1290 4412
rect 1324 4378 1358 4412
rect 1392 4378 1426 4412
rect 1460 4402 1575 4412
rect 1609 4404 1643 4436
rect 8681 4438 10026 4472
rect 8681 4404 8716 4438
rect 8750 4404 8785 4438
rect 8819 4404 8854 4438
rect 8888 4404 8923 4438
rect 8957 4404 8992 4438
rect 9026 4404 9061 4438
rect 9095 4404 9130 4438
rect 9164 4404 9199 4438
rect 9233 4404 9268 4438
rect 9302 4404 9337 4438
rect 9371 4404 9406 4438
rect 9440 4404 9475 4438
rect 9509 4404 9544 4438
rect 9578 4404 9613 4438
rect 9647 4404 9682 4438
rect 9716 4404 9751 4438
rect 9785 4404 9820 4438
rect 9854 4404 9889 4438
rect 9923 4404 9958 4438
rect 9992 4405 10026 4438
rect 9992 4404 11589 4405
rect 1609 4402 8643 4404
rect 1460 4378 1507 4402
rect 1086 4368 1507 4378
rect 1541 4368 8643 4402
rect 1086 4366 1643 4368
rect 1086 4343 1575 4366
rect 1120 4309 1154 4343
rect 1188 4309 1222 4343
rect 1256 4309 1290 4343
rect 1324 4309 1358 4343
rect 1392 4309 1426 4343
rect 1460 4333 1575 4343
rect 1460 4309 1507 4333
rect 1086 4299 1507 4309
rect 1541 4332 1575 4333
rect 1609 4334 1643 4366
rect 1677 4359 8643 4368
rect 1677 4334 1711 4359
rect 1609 4332 1711 4334
rect 1541 4325 1711 4332
rect 1745 4325 1780 4359
rect 1814 4325 1849 4359
rect 1883 4325 1918 4359
rect 1952 4325 1987 4359
rect 2021 4325 2056 4359
rect 2090 4325 2125 4359
rect 2159 4325 2194 4359
rect 2228 4325 2263 4359
rect 2297 4325 2332 4359
rect 2366 4325 2401 4359
rect 1541 4299 2401 4325
rect 1086 4298 2401 4299
rect 1086 4296 1643 4298
rect 1086 4274 1575 4296
rect 1120 4240 1154 4274
rect 1188 4240 1222 4274
rect 1256 4240 1290 4274
rect 1324 4240 1358 4274
rect 1392 4240 1426 4274
rect 1460 4264 1575 4274
rect 1460 4240 1507 4264
rect 1086 4230 1507 4240
rect 1541 4262 1575 4264
rect 1609 4264 1643 4296
rect 1677 4291 2401 4298
rect 1677 4264 1711 4291
rect 1609 4262 1711 4264
rect 1541 4257 1711 4262
rect 1745 4257 1780 4291
rect 1814 4257 1849 4291
rect 1883 4257 1918 4291
rect 1952 4257 1987 4291
rect 2021 4257 2056 4291
rect 2090 4257 2125 4291
rect 2159 4257 2194 4291
rect 2228 4257 2263 4291
rect 2297 4257 2332 4291
rect 2366 4257 2401 4291
rect 1541 4230 2401 4257
rect 1086 4228 2401 4230
rect 1086 4226 1643 4228
rect 1086 4205 1575 4226
rect 1120 4171 1154 4205
rect 1188 4171 1222 4205
rect 1256 4171 1290 4205
rect 1324 4171 1358 4205
rect 1392 4171 1426 4205
rect 1460 4195 1575 4205
rect 1460 4171 1507 4195
rect 1086 4161 1507 4171
rect 1541 4192 1575 4195
rect 1609 4194 1643 4226
rect 1677 4223 2401 4228
rect 1677 4194 1711 4223
rect 1609 4192 1711 4194
rect 1541 4189 1711 4192
rect 1745 4189 1780 4223
rect 1814 4189 1849 4223
rect 1883 4189 1918 4223
rect 1952 4189 1987 4223
rect 2021 4189 2056 4223
rect 2090 4189 2125 4223
rect 2159 4189 2194 4223
rect 2228 4189 2263 4223
rect 2297 4189 2332 4223
rect 2366 4189 2401 4223
rect 4135 4336 8643 4359
rect 8681 4371 11589 4404
rect 8681 4370 10312 4371
rect 8681 4336 8711 4370
rect 8745 4336 8779 4370
rect 8813 4336 8847 4370
rect 8881 4336 8915 4370
rect 8949 4336 8983 4370
rect 9017 4336 9051 4370
rect 9085 4336 9119 4370
rect 9153 4336 9187 4370
rect 9221 4336 9255 4370
rect 9289 4336 9323 4370
rect 9357 4336 9391 4370
rect 9425 4336 9459 4370
rect 9493 4336 9527 4370
rect 9561 4336 9595 4370
rect 9629 4336 9663 4370
rect 9697 4336 9731 4370
rect 9765 4336 9799 4370
rect 9833 4336 9867 4370
rect 9901 4336 9935 4370
rect 9969 4336 10003 4370
rect 10037 4336 10071 4370
rect 10105 4336 10139 4370
rect 10173 4336 10207 4370
rect 10241 4337 10312 4370
rect 10346 4337 10380 4371
rect 10414 4337 10448 4371
rect 10482 4337 10516 4371
rect 10550 4337 10584 4371
rect 10618 4337 10652 4371
rect 10686 4337 10720 4371
rect 10754 4337 10788 4371
rect 10822 4337 10856 4371
rect 10890 4337 10924 4371
rect 10958 4337 10992 4371
rect 11026 4337 11060 4371
rect 11094 4337 11128 4371
rect 11162 4337 11196 4371
rect 11230 4337 11264 4371
rect 11298 4337 11332 4371
rect 11366 4337 11400 4371
rect 11434 4337 11468 4371
rect 11502 4337 11536 4371
rect 11570 4337 11589 4371
rect 10241 4336 11589 4337
rect 4135 4334 11589 4336
rect 4135 4300 4179 4334
rect 4213 4300 4248 4334
rect 4282 4300 4317 4334
rect 4351 4300 4386 4334
rect 4420 4300 4455 4334
rect 4489 4300 4524 4334
rect 4558 4300 4593 4334
rect 4627 4300 4662 4334
rect 4696 4300 4731 4334
rect 4765 4300 4800 4334
rect 4834 4300 4869 4334
rect 4903 4300 4938 4334
rect 4972 4300 5007 4334
rect 5041 4300 5076 4334
rect 5110 4300 5145 4334
rect 5179 4300 5214 4334
rect 5248 4300 5283 4334
rect 5317 4300 5352 4334
rect 5386 4300 5421 4334
rect 5455 4300 5490 4334
rect 4135 4266 5490 4300
rect 4135 4232 4179 4266
rect 4213 4232 4248 4266
rect 4282 4232 4317 4266
rect 4351 4232 4386 4266
rect 4420 4232 4455 4266
rect 4489 4232 4524 4266
rect 4558 4232 4593 4266
rect 4627 4232 4662 4266
rect 4696 4232 4731 4266
rect 4765 4232 4800 4266
rect 4834 4232 4869 4266
rect 4903 4232 4938 4266
rect 4972 4232 5007 4266
rect 5041 4232 5076 4266
rect 5110 4232 5145 4266
rect 5179 4232 5214 4266
rect 5248 4232 5283 4266
rect 5317 4232 5352 4266
rect 5386 4232 5421 4266
rect 5455 4232 5490 4266
rect 4135 4198 5490 4232
rect 4135 4189 4179 4198
rect 1541 4161 1677 4189
rect 1086 4158 1677 4161
rect 1086 4156 1643 4158
rect 1086 4136 1575 4156
rect 1120 4102 1154 4136
rect 1188 4102 1222 4136
rect 1256 4102 1290 4136
rect 1324 4102 1358 4136
rect 1392 4102 1426 4136
rect 1460 4126 1575 4136
rect 1460 4102 1507 4126
rect 1086 4092 1507 4102
rect 1541 4122 1575 4126
rect 1609 4124 1643 4156
rect 1609 4122 1677 4124
rect 1541 4092 1677 4122
rect 4155 4164 4179 4189
rect 4213 4164 4248 4198
rect 4282 4164 4317 4198
rect 4351 4164 4386 4198
rect 4420 4164 4455 4198
rect 4489 4164 4524 4198
rect 4558 4164 4593 4198
rect 4627 4164 4662 4198
rect 4696 4164 4731 4198
rect 4765 4164 4800 4198
rect 4834 4164 4869 4198
rect 4903 4164 4938 4198
rect 4972 4164 5007 4198
rect 5041 4164 5076 4198
rect 5110 4164 5145 4198
rect 5179 4164 5214 4198
rect 5248 4164 5283 4198
rect 5317 4164 5352 4198
rect 5386 4164 5421 4198
rect 5455 4164 5490 4198
rect 4155 4130 5490 4164
rect 4155 4096 4179 4130
rect 4213 4096 4248 4130
rect 4282 4096 4317 4130
rect 4351 4096 4386 4130
rect 4420 4096 4455 4130
rect 4489 4096 4524 4130
rect 4558 4096 4593 4130
rect 4627 4096 4662 4130
rect 4696 4096 4731 4130
rect 4765 4096 4800 4130
rect 4834 4096 4869 4130
rect 4903 4096 4938 4130
rect 4972 4096 5007 4130
rect 5041 4096 5076 4130
rect 5110 4096 5145 4130
rect 5179 4096 5214 4130
rect 5248 4096 5283 4130
rect 5317 4096 5352 4130
rect 5386 4096 5421 4130
rect 5455 4096 5490 4130
rect 1086 4088 1677 4092
rect 1086 4086 1643 4088
rect 1086 4067 1575 4086
rect 1120 4033 1154 4067
rect 1188 4033 1222 4067
rect 1256 4033 1290 4067
rect 1324 4033 1358 4067
rect 1392 4033 1426 4067
rect 1460 4057 1575 4067
rect 1460 4033 1507 4057
rect 1086 4023 1507 4033
rect 1541 4052 1575 4057
rect 1609 4054 1643 4086
rect 1609 4052 1677 4054
rect 1541 4023 1677 4052
rect 1086 4018 1677 4023
rect 1086 4016 1643 4018
rect 1086 3998 1575 4016
rect 1120 3964 1154 3998
rect 1188 3964 1222 3998
rect 1256 3964 1290 3998
rect 1324 3964 1358 3998
rect 1392 3964 1426 3998
rect 1460 3988 1575 3998
rect 1460 3964 1507 3988
rect 1086 3954 1507 3964
rect 1541 3982 1575 3988
rect 1609 3984 1643 4016
rect 4155 4062 5490 4096
rect 4155 4028 4179 4062
rect 4213 4028 4248 4062
rect 4282 4028 4317 4062
rect 4351 4028 4386 4062
rect 4420 4028 4455 4062
rect 4489 4028 4524 4062
rect 4558 4028 4593 4062
rect 4627 4028 4662 4062
rect 4696 4028 4731 4062
rect 4765 4028 4800 4062
rect 4834 4028 4869 4062
rect 4903 4028 4938 4062
rect 4972 4028 5007 4062
rect 5041 4028 5076 4062
rect 5110 4028 5145 4062
rect 5179 4028 5214 4062
rect 5248 4028 5283 4062
rect 5317 4028 5352 4062
rect 5386 4028 5421 4062
rect 5455 4028 5490 4062
rect 4155 3994 5490 4028
rect 1609 3982 1677 3984
rect 1541 3954 1677 3982
rect 1086 3948 1677 3954
rect 1086 3946 1643 3948
rect 1086 3929 1575 3946
rect 1120 3895 1154 3929
rect 1188 3895 1222 3929
rect 1256 3895 1290 3929
rect 1324 3895 1358 3929
rect 1392 3895 1426 3929
rect 1460 3919 1575 3929
rect 1460 3895 1507 3919
rect 1086 3885 1507 3895
rect 1541 3912 1575 3919
rect 1609 3914 1643 3946
rect 1609 3912 1677 3914
rect 1541 3885 1677 3912
rect 1086 3878 1677 3885
rect 1086 3876 1643 3878
rect 1086 3860 1575 3876
rect 1120 3826 1154 3860
rect 1188 3826 1222 3860
rect 1256 3826 1290 3860
rect 1324 3826 1358 3860
rect 1392 3826 1426 3860
rect 1460 3850 1575 3860
rect 1460 3826 1507 3850
rect 1086 3816 1507 3826
rect 1541 3842 1575 3850
rect 1609 3844 1643 3876
rect 4155 3960 4179 3994
rect 4213 3960 4248 3994
rect 4282 3960 4317 3994
rect 4351 3960 4386 3994
rect 4420 3960 4455 3994
rect 4489 3960 4524 3994
rect 4558 3960 4593 3994
rect 4627 3960 4662 3994
rect 4696 3960 4731 3994
rect 4765 3960 4800 3994
rect 4834 3960 4869 3994
rect 4903 3960 4938 3994
rect 4972 3960 5007 3994
rect 5041 3960 5076 3994
rect 5110 3960 5145 3994
rect 5179 3960 5214 3994
rect 5248 3960 5283 3994
rect 5317 3960 5352 3994
rect 5386 3960 5421 3994
rect 5455 3960 5490 3994
rect 4155 3926 5490 3960
rect 4155 3892 4179 3926
rect 4213 3892 4248 3926
rect 4282 3892 4317 3926
rect 4351 3892 4386 3926
rect 4420 3892 4455 3926
rect 4489 3892 4524 3926
rect 4558 3892 4593 3926
rect 4627 3892 4662 3926
rect 4696 3892 4731 3926
rect 4765 3892 4800 3926
rect 4834 3892 4869 3926
rect 4903 3892 4938 3926
rect 4972 3892 5007 3926
rect 5041 3892 5076 3926
rect 5110 3892 5145 3926
rect 5179 3892 5214 3926
rect 5248 3892 5283 3926
rect 5317 3892 5352 3926
rect 5386 3892 5421 3926
rect 5455 3892 5490 3926
rect 8584 4301 11589 4334
rect 8584 4300 10312 4301
rect 8584 4266 8643 4300
rect 8677 4266 8711 4300
rect 8745 4266 8779 4300
rect 8813 4266 8847 4300
rect 8881 4266 8915 4300
rect 8949 4266 8983 4300
rect 9017 4266 9051 4300
rect 9085 4266 9119 4300
rect 9153 4266 9187 4300
rect 9221 4266 9255 4300
rect 9289 4266 9323 4300
rect 9357 4266 9391 4300
rect 9425 4266 9459 4300
rect 9493 4266 9527 4300
rect 9561 4266 9595 4300
rect 9629 4266 9663 4300
rect 9697 4266 9731 4300
rect 9765 4266 9799 4300
rect 9833 4266 9867 4300
rect 9901 4266 9935 4300
rect 9969 4266 10003 4300
rect 10037 4266 10071 4300
rect 10105 4266 10139 4300
rect 10173 4266 10207 4300
rect 10241 4267 10312 4300
rect 10346 4267 10380 4301
rect 10414 4267 10448 4301
rect 10482 4267 10516 4301
rect 10550 4267 10584 4301
rect 10618 4267 10652 4301
rect 10686 4267 10720 4301
rect 10754 4267 10788 4301
rect 10822 4267 10856 4301
rect 10890 4267 10924 4301
rect 10958 4267 10992 4301
rect 11026 4267 11060 4301
rect 11094 4267 11128 4301
rect 11162 4267 11196 4301
rect 11230 4267 11264 4301
rect 11298 4267 11332 4301
rect 11366 4267 11400 4301
rect 11434 4267 11468 4301
rect 11502 4267 11536 4301
rect 11570 4267 11589 4301
rect 10241 4266 11589 4267
rect 8584 4231 11589 4266
rect 8584 4230 10312 4231
rect 8584 4196 8643 4230
rect 8677 4196 8711 4230
rect 8745 4196 8779 4230
rect 8813 4196 8847 4230
rect 8881 4196 8915 4230
rect 8949 4196 8983 4230
rect 9017 4196 9051 4230
rect 9085 4196 9119 4230
rect 9153 4196 9187 4230
rect 9221 4196 9255 4230
rect 9289 4196 9323 4230
rect 9357 4196 9391 4230
rect 9425 4196 9459 4230
rect 9493 4196 9527 4230
rect 9561 4196 9595 4230
rect 9629 4196 9663 4230
rect 9697 4196 9731 4230
rect 9765 4196 9799 4230
rect 9833 4196 9867 4230
rect 9901 4196 9935 4230
rect 9969 4196 10003 4230
rect 10037 4196 10071 4230
rect 10105 4196 10139 4230
rect 10173 4196 10207 4230
rect 10241 4197 10312 4230
rect 10346 4197 10380 4231
rect 10414 4197 10448 4231
rect 10482 4197 10516 4231
rect 10550 4197 10584 4231
rect 10618 4197 10652 4231
rect 10686 4197 10720 4231
rect 10754 4197 10788 4231
rect 10822 4197 10856 4231
rect 10890 4197 10924 4231
rect 10958 4197 10992 4231
rect 11026 4197 11060 4231
rect 11094 4197 11128 4231
rect 11162 4197 11196 4231
rect 11230 4197 11264 4231
rect 11298 4197 11332 4231
rect 11366 4197 11400 4231
rect 11434 4197 11468 4231
rect 11502 4197 11536 4231
rect 11570 4197 11589 4231
rect 10241 4196 11589 4197
rect 8584 4161 11589 4196
rect 8584 4160 10312 4161
rect 8584 4126 8643 4160
rect 8677 4126 8711 4160
rect 8745 4126 8779 4160
rect 8813 4126 8847 4160
rect 8881 4126 8915 4160
rect 8949 4126 8983 4160
rect 9017 4126 9051 4160
rect 9085 4126 9119 4160
rect 9153 4126 9187 4160
rect 9221 4126 9255 4160
rect 9289 4126 9323 4160
rect 9357 4126 9391 4160
rect 9425 4126 9459 4160
rect 9493 4126 9527 4160
rect 9561 4126 9595 4160
rect 9629 4126 9663 4160
rect 9697 4126 9731 4160
rect 9765 4126 9799 4160
rect 9833 4126 9867 4160
rect 9901 4126 9935 4160
rect 9969 4126 10003 4160
rect 10037 4126 10071 4160
rect 10105 4126 10139 4160
rect 10173 4126 10207 4160
rect 10241 4127 10312 4160
rect 10346 4127 10380 4161
rect 10414 4127 10448 4161
rect 10482 4127 10516 4161
rect 10550 4127 10584 4161
rect 10618 4127 10652 4161
rect 10686 4127 10720 4161
rect 10754 4127 10788 4161
rect 10822 4127 10856 4161
rect 10890 4127 10924 4161
rect 10958 4127 10992 4161
rect 11026 4127 11060 4161
rect 11094 4127 11128 4161
rect 11162 4127 11196 4161
rect 11230 4127 11264 4161
rect 11298 4127 11332 4161
rect 11366 4127 11400 4161
rect 11434 4127 11468 4161
rect 11502 4127 11536 4161
rect 11570 4127 11589 4161
rect 10241 4126 11589 4127
rect 8584 4091 11589 4126
rect 8584 4090 10312 4091
rect 8584 4056 8643 4090
rect 8677 4056 8711 4090
rect 8745 4056 8779 4090
rect 8813 4056 8847 4090
rect 8881 4056 8915 4090
rect 8949 4056 8983 4090
rect 9017 4056 9051 4090
rect 9085 4056 9119 4090
rect 9153 4056 9187 4090
rect 9221 4056 9255 4090
rect 9289 4056 9323 4090
rect 9357 4056 9391 4090
rect 9425 4056 9459 4090
rect 9493 4056 9527 4090
rect 9561 4056 9595 4090
rect 9629 4056 9663 4090
rect 9697 4056 9731 4090
rect 9765 4056 9799 4090
rect 9833 4056 9867 4090
rect 9901 4056 9935 4090
rect 9969 4056 10003 4090
rect 10037 4056 10071 4090
rect 10105 4056 10139 4090
rect 10173 4056 10207 4090
rect 10241 4057 10312 4090
rect 10346 4057 10380 4091
rect 10414 4057 10448 4091
rect 10482 4057 10516 4091
rect 10550 4057 10584 4091
rect 10618 4057 10652 4091
rect 10686 4057 10720 4091
rect 10754 4057 10788 4091
rect 10822 4057 10856 4091
rect 10890 4057 10924 4091
rect 10958 4057 10992 4091
rect 11026 4057 11060 4091
rect 11094 4057 11128 4091
rect 11162 4057 11196 4091
rect 11230 4057 11264 4091
rect 11298 4057 11332 4091
rect 11366 4057 11400 4091
rect 11434 4057 11468 4091
rect 11502 4057 11536 4091
rect 11570 4057 11589 4091
rect 10241 4056 11589 4057
rect 8584 4021 11589 4056
rect 8584 4020 10312 4021
rect 8584 3986 8643 4020
rect 8677 3986 8711 4020
rect 8745 3986 8779 4020
rect 8813 3986 8847 4020
rect 8881 3986 8915 4020
rect 8949 3986 8983 4020
rect 9017 3986 9051 4020
rect 9085 3986 9119 4020
rect 9153 3986 9187 4020
rect 9221 3986 9255 4020
rect 9289 3986 9323 4020
rect 9357 3986 9391 4020
rect 9425 3986 9459 4020
rect 9493 3986 9527 4020
rect 9561 3986 9595 4020
rect 9629 3986 9663 4020
rect 9697 3986 9731 4020
rect 9765 3986 9799 4020
rect 9833 3986 9867 4020
rect 9901 3986 9935 4020
rect 9969 3986 10003 4020
rect 10037 3986 10071 4020
rect 10105 3986 10139 4020
rect 10173 3986 10207 4020
rect 10241 3987 10312 4020
rect 10346 3987 10380 4021
rect 10414 3987 10448 4021
rect 10482 3987 10516 4021
rect 10550 3987 10584 4021
rect 10618 3987 10652 4021
rect 10686 3987 10720 4021
rect 10754 3987 10788 4021
rect 10822 3987 10856 4021
rect 10890 3987 10924 4021
rect 10958 3987 10992 4021
rect 11026 3987 11060 4021
rect 11094 3987 11128 4021
rect 11162 3987 11196 4021
rect 11230 3987 11264 4021
rect 11298 3987 11332 4021
rect 11366 3987 11400 4021
rect 11434 3987 11468 4021
rect 11502 3987 11536 4021
rect 11570 3987 11589 4021
rect 10241 3986 11589 3987
rect 8584 3951 11589 3986
rect 8584 3950 10312 3951
rect 8584 3916 8643 3950
rect 8677 3916 8711 3950
rect 8745 3916 8779 3950
rect 8813 3916 8847 3950
rect 8881 3916 8915 3950
rect 8949 3916 8983 3950
rect 9017 3916 9051 3950
rect 9085 3916 9119 3950
rect 9153 3916 9187 3950
rect 9221 3916 9255 3950
rect 9289 3916 9323 3950
rect 9357 3916 9391 3950
rect 9425 3916 9459 3950
rect 9493 3916 9527 3950
rect 9561 3916 9595 3950
rect 9629 3916 9663 3950
rect 9697 3916 9731 3950
rect 9765 3916 9799 3950
rect 9833 3916 9867 3950
rect 9901 3916 9935 3950
rect 9969 3916 10003 3950
rect 10037 3916 10071 3950
rect 10105 3916 10139 3950
rect 10173 3916 10207 3950
rect 10241 3917 10312 3950
rect 10346 3917 10380 3951
rect 10414 3917 10448 3951
rect 10482 3917 10516 3951
rect 10550 3917 10584 3951
rect 10618 3917 10652 3951
rect 10686 3917 10720 3951
rect 10754 3917 10788 3951
rect 10822 3917 10856 3951
rect 10890 3917 10924 3951
rect 10958 3917 10992 3951
rect 11026 3917 11060 3951
rect 11094 3917 11128 3951
rect 11162 3917 11196 3951
rect 11230 3917 11264 3951
rect 11298 3917 11332 3951
rect 11366 3917 11400 3951
rect 11434 3917 11468 3951
rect 11502 3917 11536 3951
rect 11570 3917 11589 3951
rect 10241 3916 11589 3917
rect 8584 3892 11589 3916
rect 4155 3881 11589 3892
rect 4155 3880 10312 3881
rect 4155 3867 8643 3880
rect 1609 3842 1677 3844
rect 1541 3816 1677 3842
rect 1086 3808 1677 3816
rect 1086 3806 1643 3808
rect 1086 3791 1575 3806
rect 1120 3757 1154 3791
rect 1188 3757 1222 3791
rect 1256 3757 1290 3791
rect 1324 3757 1358 3791
rect 1392 3757 1426 3791
rect 1460 3781 1575 3791
rect 1460 3757 1507 3781
rect 1086 3747 1507 3757
rect 1541 3772 1575 3781
rect 1609 3774 1643 3806
rect 1609 3772 1677 3774
rect 1541 3747 1677 3772
rect 1086 3738 1677 3747
rect 1086 3736 1643 3738
rect 1086 3722 1575 3736
rect 1120 3688 1154 3722
rect 1188 3688 1222 3722
rect 1256 3688 1290 3722
rect 1324 3688 1358 3722
rect 1392 3688 1426 3722
rect 1460 3712 1575 3722
rect 1460 3688 1507 3712
rect 1086 3678 1507 3688
rect 1541 3702 1575 3712
rect 1609 3704 1643 3736
rect 1609 3702 1677 3704
rect 1541 3678 1677 3702
rect 1086 3668 1677 3678
rect 1086 3666 1643 3668
rect 1086 3653 1575 3666
rect 1460 3643 1575 3653
rect 1460 3609 1507 3643
rect 1541 3632 1575 3643
rect 1609 3634 1643 3666
rect 1609 3632 1677 3634
rect 1541 3609 1677 3632
rect 1460 3598 1677 3609
rect 1460 3596 1643 3598
rect 1460 3574 1575 3596
rect 1460 3540 1507 3574
rect 1541 3562 1575 3574
rect 1609 3564 1643 3596
rect 1609 3562 1677 3564
rect 1541 3540 1677 3562
rect 1460 3528 1677 3540
rect 1460 3526 1643 3528
rect 1460 3505 1575 3526
rect 1460 3471 1507 3505
rect 1541 3492 1575 3505
rect 1609 3494 1643 3526
rect 1609 3492 1677 3494
rect 1541 3471 1677 3492
rect 1460 3458 1677 3471
rect 1460 3456 1643 3458
rect 1460 3436 1575 3456
rect 1460 3402 1507 3436
rect 1541 3422 1575 3436
rect 1609 3424 1643 3456
rect 1609 3422 1677 3424
rect 1541 3402 1677 3422
rect 1460 3388 1677 3402
rect 1460 3386 1643 3388
rect 1460 3367 1575 3386
rect 1460 3333 1507 3367
rect 1541 3352 1575 3367
rect 1609 3354 1643 3386
rect 1609 3352 1677 3354
rect 1541 3333 1677 3352
rect 1460 3318 1677 3333
rect 1460 3316 1643 3318
rect 1460 3298 1575 3316
rect 1460 3264 1507 3298
rect 1541 3282 1575 3298
rect 1609 3284 1643 3316
rect 1609 3282 1677 3284
rect 1541 3264 1677 3282
rect 1460 3258 1677 3264
rect 8677 3846 8711 3880
rect 8745 3846 8779 3880
rect 8813 3846 8847 3880
rect 8881 3846 8915 3880
rect 8949 3846 8983 3880
rect 9017 3846 9051 3880
rect 9085 3846 9119 3880
rect 9153 3846 9187 3880
rect 9221 3846 9255 3880
rect 9289 3846 9323 3880
rect 9357 3846 9391 3880
rect 9425 3846 9459 3880
rect 9493 3846 9527 3880
rect 9561 3846 9595 3880
rect 9629 3846 9663 3880
rect 9697 3846 9731 3880
rect 9765 3846 9799 3880
rect 9833 3846 9867 3880
rect 9901 3846 9935 3880
rect 9969 3846 10003 3880
rect 10037 3846 10071 3880
rect 10105 3846 10139 3880
rect 10173 3846 10207 3880
rect 10241 3847 10312 3880
rect 10346 3847 10380 3881
rect 10414 3847 10448 3881
rect 10482 3847 10516 3881
rect 10550 3847 10584 3881
rect 10618 3847 10652 3881
rect 10686 3847 10720 3881
rect 10754 3847 10788 3881
rect 10822 3847 10856 3881
rect 10890 3847 10924 3881
rect 10958 3847 10992 3881
rect 11026 3847 11060 3881
rect 11094 3847 11128 3881
rect 11162 3847 11196 3881
rect 11230 3847 11264 3881
rect 11298 3847 11332 3881
rect 11366 3847 11400 3881
rect 11434 3847 11468 3881
rect 11502 3847 11536 3881
rect 11570 3847 11589 3881
rect 10241 3846 11589 3847
rect 8643 3811 11589 3846
rect 8643 3810 10312 3811
rect 8677 3776 8711 3810
rect 8745 3776 8779 3810
rect 8813 3776 8847 3810
rect 8881 3776 8915 3810
rect 8949 3776 8983 3810
rect 9017 3776 9051 3810
rect 9085 3776 9119 3810
rect 9153 3776 9187 3810
rect 9221 3776 9255 3810
rect 9289 3776 9323 3810
rect 9357 3776 9391 3810
rect 9425 3776 9459 3810
rect 9493 3776 9527 3810
rect 9561 3776 9595 3810
rect 9629 3776 9663 3810
rect 9697 3776 9731 3810
rect 9765 3776 9799 3810
rect 9833 3776 9867 3810
rect 9901 3776 9935 3810
rect 9969 3776 10003 3810
rect 10037 3776 10071 3810
rect 10105 3776 10139 3810
rect 10173 3776 10207 3810
rect 10241 3777 10312 3810
rect 10346 3777 10380 3811
rect 10414 3777 10448 3811
rect 10482 3777 10516 3811
rect 10550 3777 10584 3811
rect 10618 3777 10652 3811
rect 10686 3777 10720 3811
rect 10754 3777 10788 3811
rect 10822 3777 10856 3811
rect 10890 3777 10924 3811
rect 10958 3777 10992 3811
rect 11026 3777 11060 3811
rect 11094 3777 11128 3811
rect 11162 3777 11196 3811
rect 11230 3777 11264 3811
rect 11298 3777 11332 3811
rect 11366 3777 11400 3811
rect 11434 3777 11468 3811
rect 11502 3777 11536 3811
rect 11570 3777 11589 3811
rect 10241 3776 11589 3777
rect 8643 3741 11589 3776
rect 8643 3740 10312 3741
rect 8677 3706 8711 3740
rect 8745 3706 8779 3740
rect 8813 3706 8847 3740
rect 8881 3706 8915 3740
rect 8949 3706 8983 3740
rect 9017 3706 9051 3740
rect 9085 3706 9119 3740
rect 9153 3706 9187 3740
rect 9221 3706 9255 3740
rect 9289 3706 9323 3740
rect 9357 3706 9391 3740
rect 9425 3706 9459 3740
rect 9493 3706 9527 3740
rect 9561 3706 9595 3740
rect 9629 3706 9663 3740
rect 9697 3706 9731 3740
rect 9765 3706 9799 3740
rect 9833 3706 9867 3740
rect 9901 3706 9935 3740
rect 9969 3706 10003 3740
rect 10037 3706 10071 3740
rect 10105 3706 10139 3740
rect 10173 3706 10207 3740
rect 10241 3707 10312 3740
rect 10346 3707 10380 3741
rect 10414 3707 10448 3741
rect 10482 3707 10516 3741
rect 10550 3707 10584 3741
rect 10618 3707 10652 3741
rect 10686 3707 10720 3741
rect 10754 3707 10788 3741
rect 10822 3707 10856 3741
rect 10890 3707 10924 3741
rect 10958 3707 10992 3741
rect 11026 3707 11060 3741
rect 11094 3707 11128 3741
rect 11162 3707 11196 3741
rect 11230 3707 11264 3741
rect 11298 3707 11332 3741
rect 11366 3707 11400 3741
rect 11434 3707 11468 3741
rect 11502 3707 11536 3741
rect 11570 3707 11589 3741
rect 10241 3706 11589 3707
rect 8643 3671 11589 3706
rect 8643 3670 10312 3671
rect 8677 3636 8711 3670
rect 8745 3636 8779 3670
rect 8813 3636 8847 3670
rect 8881 3636 8915 3670
rect 8949 3636 8983 3670
rect 9017 3636 9051 3670
rect 9085 3636 9119 3670
rect 9153 3636 9187 3670
rect 9221 3636 9255 3670
rect 9289 3636 9323 3670
rect 9357 3636 9391 3670
rect 9425 3636 9459 3670
rect 9493 3636 9527 3670
rect 9561 3636 9595 3670
rect 9629 3636 9663 3670
rect 9697 3636 9731 3670
rect 9765 3636 9799 3670
rect 9833 3636 9867 3670
rect 9901 3636 9935 3670
rect 9969 3636 10003 3670
rect 10037 3636 10071 3670
rect 10105 3636 10139 3670
rect 10173 3636 10207 3670
rect 10241 3637 10312 3670
rect 10346 3637 10380 3671
rect 10414 3637 10448 3671
rect 10482 3637 10516 3671
rect 10550 3637 10584 3671
rect 10618 3637 10652 3671
rect 10686 3637 10720 3671
rect 10754 3637 10788 3671
rect 10822 3637 10856 3671
rect 10890 3637 10924 3671
rect 10958 3637 10992 3671
rect 11026 3637 11060 3671
rect 11094 3637 11128 3671
rect 11162 3637 11196 3671
rect 11230 3637 11264 3671
rect 11298 3637 11332 3671
rect 11366 3637 11400 3671
rect 11434 3637 11468 3671
rect 11502 3637 11536 3671
rect 11570 3637 11589 3671
rect 10241 3636 11589 3637
rect 8643 3601 11589 3636
rect 8643 3600 10312 3601
rect 8677 3566 8711 3600
rect 8745 3566 8779 3600
rect 8813 3566 8847 3600
rect 8881 3566 8915 3600
rect 8949 3566 8983 3600
rect 9017 3566 9051 3600
rect 9085 3566 9119 3600
rect 9153 3566 9187 3600
rect 9221 3566 9255 3600
rect 9289 3566 9323 3600
rect 9357 3566 9391 3600
rect 9425 3566 9459 3600
rect 9493 3566 9527 3600
rect 9561 3566 9595 3600
rect 9629 3566 9663 3600
rect 9697 3566 9731 3600
rect 9765 3566 9799 3600
rect 9833 3566 9867 3600
rect 9901 3566 9935 3600
rect 9969 3566 10003 3600
rect 10037 3566 10071 3600
rect 10105 3566 10139 3600
rect 10173 3566 10207 3600
rect 10241 3567 10312 3600
rect 10346 3567 10380 3601
rect 10414 3567 10448 3601
rect 10482 3567 10516 3601
rect 10550 3567 10584 3601
rect 10618 3567 10652 3601
rect 10686 3567 10720 3601
rect 10754 3567 10788 3601
rect 10822 3567 10856 3601
rect 10890 3567 10924 3601
rect 10958 3567 10992 3601
rect 11026 3567 11060 3601
rect 11094 3567 11128 3601
rect 11162 3567 11196 3601
rect 11230 3567 11264 3601
rect 11298 3567 11332 3601
rect 11366 3567 11400 3601
rect 11434 3567 11468 3601
rect 11502 3567 11536 3601
rect 11570 3567 11589 3601
rect 10241 3566 11589 3567
rect 8643 3531 11589 3566
rect 8643 3530 10312 3531
rect 8677 3496 8711 3530
rect 8745 3496 8779 3530
rect 8813 3496 8847 3530
rect 8881 3496 8915 3530
rect 8949 3496 8983 3530
rect 9017 3496 9051 3530
rect 9085 3496 9119 3530
rect 9153 3496 9187 3530
rect 9221 3496 9255 3530
rect 9289 3496 9323 3530
rect 9357 3496 9391 3530
rect 9425 3496 9459 3530
rect 9493 3496 9527 3530
rect 9561 3496 9595 3530
rect 9629 3496 9663 3530
rect 9697 3496 9731 3530
rect 9765 3496 9799 3530
rect 9833 3496 9867 3530
rect 9901 3496 9935 3530
rect 9969 3496 10003 3530
rect 10037 3496 10071 3530
rect 10105 3496 10139 3530
rect 10173 3496 10207 3530
rect 10241 3497 10312 3530
rect 10346 3497 10380 3531
rect 10414 3497 10448 3531
rect 10482 3497 10516 3531
rect 10550 3497 10584 3531
rect 10618 3497 10652 3531
rect 10686 3497 10720 3531
rect 10754 3497 10788 3531
rect 10822 3497 10856 3531
rect 10890 3497 10924 3531
rect 10958 3497 10992 3531
rect 11026 3497 11060 3531
rect 11094 3497 11128 3531
rect 11162 3497 11196 3531
rect 11230 3497 11264 3531
rect 11298 3497 11332 3531
rect 11366 3497 11400 3531
rect 11434 3497 11468 3531
rect 11502 3497 11536 3531
rect 11570 3497 11589 3531
rect 10241 3496 11589 3497
rect 8643 3461 11589 3496
rect 8643 3460 10312 3461
rect 8677 3426 8711 3460
rect 8745 3426 8779 3460
rect 8813 3426 8847 3460
rect 8881 3426 8915 3460
rect 8949 3426 8983 3460
rect 9017 3426 9051 3460
rect 9085 3426 9119 3460
rect 9153 3426 9187 3460
rect 9221 3426 9255 3460
rect 9289 3426 9323 3460
rect 9357 3426 9391 3460
rect 9425 3426 9459 3460
rect 9493 3426 9527 3460
rect 9561 3426 9595 3460
rect 9629 3426 9663 3460
rect 9697 3426 9731 3460
rect 9765 3426 9799 3460
rect 9833 3426 9867 3460
rect 9901 3426 9935 3460
rect 9969 3426 10003 3460
rect 10037 3426 10071 3460
rect 10105 3426 10139 3460
rect 10173 3426 10207 3460
rect 10241 3427 10312 3460
rect 10346 3427 10380 3461
rect 10414 3427 10448 3461
rect 10482 3427 10516 3461
rect 10550 3427 10584 3461
rect 10618 3427 10652 3461
rect 10686 3427 10720 3461
rect 10754 3427 10788 3461
rect 10822 3427 10856 3461
rect 10890 3427 10924 3461
rect 10958 3427 10992 3461
rect 11026 3427 11060 3461
rect 11094 3427 11128 3461
rect 11162 3427 11196 3461
rect 11230 3427 11264 3461
rect 11298 3427 11332 3461
rect 11366 3427 11400 3461
rect 11434 3427 11468 3461
rect 11502 3427 11536 3461
rect 11570 3427 11589 3461
rect 10241 3426 11589 3427
rect 8643 3391 11589 3426
rect 8643 3390 10312 3391
rect 8677 3356 8711 3390
rect 8745 3356 8779 3390
rect 8813 3356 8847 3390
rect 8881 3356 8915 3390
rect 8949 3356 8983 3390
rect 9017 3356 9051 3390
rect 9085 3356 9119 3390
rect 9153 3356 9187 3390
rect 9221 3356 9255 3390
rect 9289 3356 9323 3390
rect 9357 3356 9391 3390
rect 9425 3356 9459 3390
rect 9493 3356 9527 3390
rect 9561 3356 9595 3390
rect 9629 3356 9663 3390
rect 9697 3356 9731 3390
rect 9765 3356 9799 3390
rect 9833 3356 9867 3390
rect 9901 3356 9935 3390
rect 9969 3356 10003 3390
rect 10037 3356 10071 3390
rect 10105 3356 10139 3390
rect 10173 3356 10207 3390
rect 10241 3357 10312 3390
rect 10346 3357 10380 3391
rect 10414 3357 10448 3391
rect 10482 3357 10516 3391
rect 10550 3357 10584 3391
rect 10618 3357 10652 3391
rect 10686 3357 10720 3391
rect 10754 3357 10788 3391
rect 10822 3357 10856 3391
rect 10890 3357 10924 3391
rect 10958 3357 10992 3391
rect 11026 3357 11060 3391
rect 11094 3357 11128 3391
rect 11162 3357 11196 3391
rect 11230 3357 11264 3391
rect 11298 3357 11332 3391
rect 11366 3357 11400 3391
rect 11434 3357 11468 3391
rect 11502 3357 11536 3391
rect 11570 3357 11589 3391
rect 10241 3356 11589 3357
rect 8643 3321 11589 3356
rect 8643 3320 10312 3321
rect 8677 3286 8711 3320
rect 8745 3286 8779 3320
rect 8813 3286 8847 3320
rect 8881 3286 8915 3320
rect 8949 3286 8983 3320
rect 9017 3286 9051 3320
rect 9085 3286 9119 3320
rect 9153 3286 9187 3320
rect 9221 3286 9255 3320
rect 9289 3286 9323 3320
rect 9357 3286 9391 3320
rect 9425 3286 9459 3320
rect 9493 3286 9527 3320
rect 9561 3286 9595 3320
rect 9629 3286 9663 3320
rect 9697 3286 9731 3320
rect 9765 3286 9799 3320
rect 9833 3286 9867 3320
rect 9901 3286 9935 3320
rect 9969 3286 10003 3320
rect 10037 3286 10071 3320
rect 10105 3286 10139 3320
rect 10173 3286 10207 3320
rect 10241 3287 10312 3320
rect 10346 3287 10380 3321
rect 10414 3287 10448 3321
rect 10482 3287 10516 3321
rect 10550 3287 10584 3321
rect 10618 3287 10652 3321
rect 10686 3287 10720 3321
rect 10754 3287 10788 3321
rect 10822 3287 10856 3321
rect 10890 3287 10924 3321
rect 10958 3287 10992 3321
rect 11026 3287 11060 3321
rect 11094 3287 11128 3321
rect 11162 3287 11196 3321
rect 11230 3287 11264 3321
rect 11298 3287 11332 3321
rect 11366 3287 11400 3321
rect 11434 3287 11468 3321
rect 11502 3287 11536 3321
rect 11570 3287 11589 3321
rect 10241 3286 11589 3287
rect 1460 3248 1740 3258
rect 1460 3246 1643 3248
rect 1460 3229 1575 3246
rect 1460 3195 1507 3229
rect 1541 3212 1575 3229
rect 1609 3214 1643 3246
rect 1677 3224 1740 3248
rect 1774 3224 1809 3258
rect 1843 3224 1878 3258
rect 1912 3224 1947 3258
rect 1981 3224 2016 3258
rect 2050 3224 2085 3258
rect 2119 3224 2154 3258
rect 2188 3224 2223 3258
rect 2257 3224 2292 3258
rect 2326 3224 2361 3258
rect 2395 3224 2430 3258
rect 2464 3224 2499 3258
rect 2533 3224 2568 3258
rect 2602 3224 2637 3258
rect 2671 3224 2706 3258
rect 2740 3224 2775 3258
rect 2809 3224 2844 3258
rect 1677 3214 2844 3224
rect 1609 3212 2844 3214
rect 1541 3195 2844 3212
rect 1460 3190 2844 3195
rect 1460 3178 1740 3190
rect 1460 3176 1643 3178
rect 1460 3160 1575 3176
rect 1460 3126 1507 3160
rect 1541 3142 1575 3160
rect 1609 3144 1643 3176
rect 1677 3156 1740 3178
rect 1774 3156 1809 3190
rect 1843 3156 1878 3190
rect 1912 3156 1947 3190
rect 1981 3156 2016 3190
rect 2050 3156 2085 3190
rect 2119 3156 2154 3190
rect 2188 3156 2223 3190
rect 2257 3156 2292 3190
rect 2326 3156 2361 3190
rect 2395 3156 2430 3190
rect 2464 3156 2499 3190
rect 2533 3156 2568 3190
rect 2602 3156 2637 3190
rect 2671 3156 2706 3190
rect 2740 3156 2775 3190
rect 2809 3156 2844 3190
rect 1677 3144 2844 3156
rect 1609 3142 2844 3144
rect 1541 3126 2844 3142
rect 1460 3122 2844 3126
rect 1460 3108 1740 3122
rect 1460 3107 1643 3108
rect 1460 3091 1575 3107
rect 1460 3057 1507 3091
rect 1541 3073 1575 3091
rect 1609 3074 1643 3107
rect 1677 3088 1740 3108
rect 1774 3088 1809 3122
rect 1843 3088 1878 3122
rect 1912 3088 1947 3122
rect 1981 3088 2016 3122
rect 2050 3088 2085 3122
rect 2119 3088 2154 3122
rect 2188 3088 2223 3122
rect 2257 3088 2292 3122
rect 2326 3088 2361 3122
rect 2395 3088 2430 3122
rect 2464 3088 2499 3122
rect 2533 3088 2568 3122
rect 2602 3088 2637 3122
rect 2671 3088 2706 3122
rect 2740 3088 2775 3122
rect 2809 3088 2844 3122
rect 4782 3088 4806 3258
rect 8643 3251 11589 3286
rect 8643 3250 10312 3251
rect 8677 3216 8711 3250
rect 8745 3216 8779 3250
rect 8813 3216 8847 3250
rect 8881 3216 8915 3250
rect 8949 3216 8983 3250
rect 9017 3216 9051 3250
rect 9085 3216 9119 3250
rect 9153 3216 9187 3250
rect 9221 3216 9255 3250
rect 9289 3216 9323 3250
rect 9357 3216 9391 3250
rect 9425 3216 9459 3250
rect 9493 3216 9527 3250
rect 9561 3216 9595 3250
rect 9629 3216 9663 3250
rect 9697 3216 9731 3250
rect 9765 3216 9799 3250
rect 9833 3216 9867 3250
rect 9901 3216 9935 3250
rect 9969 3216 10003 3250
rect 10037 3216 10071 3250
rect 10105 3216 10139 3250
rect 10173 3216 10207 3250
rect 10241 3217 10312 3250
rect 10346 3217 10380 3251
rect 10414 3217 10448 3251
rect 10482 3217 10516 3251
rect 10550 3217 10584 3251
rect 10618 3217 10652 3251
rect 10686 3217 10720 3251
rect 10754 3217 10788 3251
rect 10822 3217 10856 3251
rect 10890 3217 10924 3251
rect 10958 3217 10992 3251
rect 11026 3217 11060 3251
rect 11094 3217 11128 3251
rect 11162 3217 11196 3251
rect 11230 3217 11264 3251
rect 11298 3217 11332 3251
rect 11366 3217 11400 3251
rect 11434 3217 11468 3251
rect 11502 3217 11536 3251
rect 11570 3217 11589 3251
rect 10241 3216 11589 3217
rect 8643 3181 11589 3216
rect 8643 3180 10312 3181
rect 8677 3146 8711 3180
rect 8745 3146 8779 3180
rect 8813 3146 8847 3180
rect 8881 3146 8915 3180
rect 8949 3146 8983 3180
rect 9017 3146 9051 3180
rect 9085 3146 9119 3180
rect 9153 3146 9187 3180
rect 9221 3146 9255 3180
rect 9289 3146 9323 3180
rect 9357 3146 9391 3180
rect 9425 3146 9459 3180
rect 9493 3146 9527 3180
rect 9561 3146 9595 3180
rect 9629 3146 9663 3180
rect 9697 3146 9731 3180
rect 9765 3146 9799 3180
rect 9833 3146 9867 3180
rect 9901 3146 9935 3180
rect 9969 3146 10003 3180
rect 10037 3146 10071 3180
rect 10105 3146 10139 3180
rect 10173 3146 10207 3180
rect 10241 3147 10312 3180
rect 10346 3147 10380 3181
rect 10414 3147 10448 3181
rect 10482 3147 10516 3181
rect 10550 3147 10584 3181
rect 10618 3147 10652 3181
rect 10686 3147 10720 3181
rect 10754 3147 10788 3181
rect 10822 3147 10856 3181
rect 10890 3147 10924 3181
rect 10958 3147 10992 3181
rect 11026 3147 11060 3181
rect 11094 3147 11128 3181
rect 11162 3147 11196 3181
rect 11230 3147 11264 3181
rect 11298 3147 11332 3181
rect 11366 3147 11400 3181
rect 11434 3147 11468 3181
rect 11502 3147 11536 3181
rect 11570 3147 11589 3181
rect 10241 3146 11589 3147
rect 8643 3111 11589 3146
rect 8643 3110 10312 3111
rect 1609 3073 1677 3074
rect 1541 3057 1677 3073
rect 1460 3038 1677 3057
rect 1460 3022 1575 3038
rect 1460 2988 1507 3022
rect 1541 3004 1575 3022
rect 1609 3004 1643 3038
rect 1541 2988 1677 3004
rect 1460 2969 1677 2988
rect 1460 2953 1575 2969
rect 1460 2919 1507 2953
rect 1541 2935 1575 2953
rect 1609 2935 1643 2969
rect 1541 2919 1677 2935
rect 1460 2900 1677 2919
rect 1460 2884 1575 2900
rect 1460 2850 1507 2884
rect 1541 2866 1575 2884
rect 1609 2866 1643 2900
rect 1541 2850 1677 2866
rect 1460 2831 1677 2850
rect 1460 2815 1575 2831
rect 1460 2781 1507 2815
rect 1541 2797 1575 2815
rect 1609 2797 1643 2831
rect 1541 2781 1677 2797
rect 1460 2762 1677 2781
rect 1460 2746 1575 2762
rect 1460 2712 1507 2746
rect 1541 2728 1575 2746
rect 1609 2728 1643 2762
rect 1541 2712 1677 2728
rect 1460 2693 1677 2712
rect 1460 2677 1575 2693
rect 1460 2643 1507 2677
rect 1541 2659 1575 2677
rect 1609 2659 1643 2693
rect 1541 2643 1677 2659
rect 1460 2624 1677 2643
rect 1460 2609 1575 2624
rect 1460 2575 1507 2609
rect 1541 2590 1575 2609
rect 1609 2590 1643 2624
rect 1541 2575 1677 2590
rect 1460 2555 1677 2575
rect 1460 2541 1575 2555
rect 1460 2507 1507 2541
rect 1541 2521 1575 2541
rect 1609 2521 1643 2555
rect 1541 2507 1677 2521
rect 1460 2486 1677 2507
rect 1460 2473 1575 2486
rect 1460 2439 1507 2473
rect 1541 2452 1575 2473
rect 1609 2452 1643 2486
rect 1541 2439 1677 2452
rect 1460 2417 1677 2439
rect 1460 2405 1575 2417
rect 1460 2371 1507 2405
rect 1541 2383 1575 2405
rect 1609 2383 1643 2417
rect 1541 2371 1677 2383
rect 1460 2361 1677 2371
rect 8677 3076 8711 3110
rect 8745 3076 8779 3110
rect 8813 3076 8847 3110
rect 8881 3076 8915 3110
rect 8949 3076 8983 3110
rect 9017 3076 9051 3110
rect 9085 3076 9119 3110
rect 9153 3076 9187 3110
rect 9221 3076 9255 3110
rect 9289 3076 9323 3110
rect 9357 3076 9391 3110
rect 9425 3076 9459 3110
rect 9493 3076 9527 3110
rect 9561 3076 9595 3110
rect 9629 3076 9663 3110
rect 9697 3076 9731 3110
rect 9765 3076 9799 3110
rect 9833 3076 9867 3110
rect 9901 3076 9935 3110
rect 9969 3076 10003 3110
rect 10037 3076 10071 3110
rect 10105 3076 10139 3110
rect 10173 3076 10207 3110
rect 10241 3077 10312 3110
rect 10346 3077 10380 3111
rect 10414 3077 10448 3111
rect 10482 3077 10516 3111
rect 10550 3077 10584 3111
rect 10618 3077 10652 3111
rect 10686 3077 10720 3111
rect 10754 3077 10788 3111
rect 10822 3077 10856 3111
rect 10890 3077 10924 3111
rect 10958 3077 10992 3111
rect 11026 3077 11060 3111
rect 11094 3077 11128 3111
rect 11162 3077 11196 3111
rect 11230 3077 11264 3111
rect 11298 3077 11332 3111
rect 11366 3077 11400 3111
rect 11434 3077 11468 3111
rect 11502 3077 11536 3111
rect 11570 3077 11589 3111
rect 10241 3076 11589 3077
rect 8643 3041 11589 3076
rect 8643 3040 10312 3041
rect 8677 3006 8711 3040
rect 8745 3006 8779 3040
rect 8813 3006 8847 3040
rect 8881 3006 8915 3040
rect 8949 3006 8983 3040
rect 9017 3006 9051 3040
rect 9085 3006 9119 3040
rect 9153 3006 9187 3040
rect 9221 3006 9255 3040
rect 9289 3006 9323 3040
rect 9357 3006 9391 3040
rect 9425 3006 9459 3040
rect 9493 3006 9527 3040
rect 9561 3006 9595 3040
rect 9629 3006 9663 3040
rect 9697 3006 9731 3040
rect 9765 3006 9799 3040
rect 9833 3006 9867 3040
rect 9901 3006 9935 3040
rect 9969 3006 10003 3040
rect 10037 3006 10071 3040
rect 10105 3006 10139 3040
rect 10173 3006 10207 3040
rect 10241 3007 10312 3040
rect 10346 3007 10380 3041
rect 10414 3007 10448 3041
rect 10482 3007 10516 3041
rect 10550 3007 10584 3041
rect 10618 3007 10652 3041
rect 10686 3007 10720 3041
rect 10754 3007 10788 3041
rect 10822 3007 10856 3041
rect 10890 3007 10924 3041
rect 10958 3007 10992 3041
rect 11026 3007 11060 3041
rect 11094 3007 11128 3041
rect 11162 3007 11196 3041
rect 11230 3007 11264 3041
rect 11298 3007 11332 3041
rect 11366 3007 11400 3041
rect 11434 3007 11468 3041
rect 11502 3007 11536 3041
rect 11570 3007 11589 3041
rect 10241 3006 11589 3007
rect 8643 2971 11589 3006
rect 8643 2970 10312 2971
rect 8677 2936 8711 2970
rect 8745 2936 8779 2970
rect 8813 2936 8847 2970
rect 8881 2936 8915 2970
rect 8949 2936 8983 2970
rect 9017 2936 9051 2970
rect 9085 2936 9119 2970
rect 9153 2936 9187 2970
rect 9221 2936 9255 2970
rect 9289 2936 9323 2970
rect 9357 2936 9391 2970
rect 9425 2936 9459 2970
rect 9493 2936 9527 2970
rect 9561 2936 9595 2970
rect 9629 2936 9663 2970
rect 9697 2936 9731 2970
rect 9765 2936 9799 2970
rect 9833 2936 9867 2970
rect 9901 2936 9935 2970
rect 9969 2936 10003 2970
rect 10037 2936 10071 2970
rect 10105 2936 10139 2970
rect 10173 2936 10207 2970
rect 10241 2937 10312 2970
rect 10346 2937 10380 2971
rect 10414 2937 10448 2971
rect 10482 2937 10516 2971
rect 10550 2937 10584 2971
rect 10618 2937 10652 2971
rect 10686 2937 10720 2971
rect 10754 2937 10788 2971
rect 10822 2937 10856 2971
rect 10890 2937 10924 2971
rect 10958 2937 10992 2971
rect 11026 2937 11060 2971
rect 11094 2937 11128 2971
rect 11162 2937 11196 2971
rect 11230 2937 11264 2971
rect 11298 2937 11332 2971
rect 11366 2937 11400 2971
rect 11434 2937 11468 2971
rect 11502 2937 11536 2971
rect 11570 2937 11589 2971
rect 10241 2936 11589 2937
rect 8643 2901 11589 2936
rect 8643 2900 10312 2901
rect 8677 2866 8711 2900
rect 8745 2866 8779 2900
rect 8813 2866 8847 2900
rect 8881 2866 8915 2900
rect 8949 2866 8983 2900
rect 9017 2866 9051 2900
rect 9085 2866 9119 2900
rect 9153 2866 9187 2900
rect 9221 2866 9255 2900
rect 9289 2866 9323 2900
rect 9357 2866 9391 2900
rect 9425 2866 9459 2900
rect 9493 2866 9527 2900
rect 9561 2866 9595 2900
rect 9629 2866 9663 2900
rect 9697 2866 9731 2900
rect 9765 2866 9799 2900
rect 9833 2866 9867 2900
rect 9901 2866 9935 2900
rect 9969 2866 10003 2900
rect 10037 2866 10071 2900
rect 10105 2866 10139 2900
rect 10173 2866 10207 2900
rect 10241 2867 10312 2900
rect 10346 2867 10380 2901
rect 10414 2867 10448 2901
rect 10482 2867 10516 2901
rect 10550 2867 10584 2901
rect 10618 2867 10652 2901
rect 10686 2867 10720 2901
rect 10754 2867 10788 2901
rect 10822 2867 10856 2901
rect 10890 2867 10924 2901
rect 10958 2867 10992 2901
rect 11026 2867 11060 2901
rect 11094 2867 11128 2901
rect 11162 2867 11196 2901
rect 11230 2867 11264 2901
rect 11298 2867 11332 2901
rect 11366 2867 11400 2901
rect 11434 2867 11468 2901
rect 11502 2867 11536 2901
rect 11570 2867 11589 2901
rect 10241 2866 11589 2867
rect 8643 2831 11589 2866
rect 8643 2830 10312 2831
rect 8677 2796 8711 2830
rect 8745 2796 8779 2830
rect 8813 2796 8847 2830
rect 8881 2796 8915 2830
rect 8949 2796 8983 2830
rect 9017 2796 9051 2830
rect 9085 2796 9119 2830
rect 9153 2796 9187 2830
rect 9221 2796 9255 2830
rect 9289 2796 9323 2830
rect 9357 2796 9391 2830
rect 9425 2796 9459 2830
rect 9493 2796 9527 2830
rect 9561 2796 9595 2830
rect 9629 2796 9663 2830
rect 9697 2796 9731 2830
rect 9765 2796 9799 2830
rect 9833 2796 9867 2830
rect 9901 2796 9935 2830
rect 9969 2796 10003 2830
rect 10037 2796 10071 2830
rect 10105 2796 10139 2830
rect 10173 2796 10207 2830
rect 10241 2797 10312 2830
rect 10346 2797 10380 2831
rect 10414 2797 10448 2831
rect 10482 2797 10516 2831
rect 10550 2797 10584 2831
rect 10618 2797 10652 2831
rect 10686 2797 10720 2831
rect 10754 2797 10788 2831
rect 10822 2797 10856 2831
rect 10890 2797 10924 2831
rect 10958 2797 10992 2831
rect 11026 2797 11060 2831
rect 11094 2797 11128 2831
rect 11162 2797 11196 2831
rect 11230 2797 11264 2831
rect 11298 2797 11332 2831
rect 11366 2797 11400 2831
rect 11434 2797 11468 2831
rect 11502 2797 11536 2831
rect 11570 2797 11589 2831
rect 10241 2796 11589 2797
rect 8643 2761 11589 2796
rect 8677 2727 8711 2761
rect 8745 2727 8779 2761
rect 8813 2727 8847 2761
rect 8881 2727 8915 2761
rect 8949 2727 8983 2761
rect 9017 2727 9051 2761
rect 9085 2727 9119 2761
rect 9153 2727 9187 2761
rect 9221 2727 9255 2761
rect 9289 2727 9323 2761
rect 9357 2727 9391 2761
rect 9425 2727 9459 2761
rect 9493 2727 9527 2761
rect 9561 2727 9595 2761
rect 9629 2727 9663 2761
rect 9697 2727 9731 2761
rect 9765 2727 9799 2761
rect 9833 2727 9867 2761
rect 9901 2727 9935 2761
rect 9969 2727 10003 2761
rect 10037 2727 10071 2761
rect 10105 2727 10139 2761
rect 10173 2727 10207 2761
rect 10241 2727 10312 2761
rect 10346 2727 10380 2761
rect 10414 2727 10448 2761
rect 10482 2727 10516 2761
rect 10550 2727 10584 2761
rect 10618 2727 10652 2761
rect 10686 2727 10720 2761
rect 10754 2727 10788 2761
rect 10822 2727 10856 2761
rect 10890 2727 10924 2761
rect 10958 2727 10992 2761
rect 11026 2727 11060 2761
rect 11094 2727 11128 2761
rect 11162 2727 11196 2761
rect 11230 2727 11264 2761
rect 11298 2727 11332 2761
rect 11366 2727 11400 2761
rect 11434 2727 11468 2761
rect 11502 2727 11536 2761
rect 11570 2730 11589 2761
rect 12582 4363 13390 4387
rect 12582 4329 12595 4363
rect 12629 4329 12663 4363
rect 12697 4329 12731 4363
rect 12765 4329 12799 4363
rect 12833 4329 12867 4363
rect 12901 4329 12935 4363
rect 12969 4329 13003 4363
rect 13037 4329 13071 4363
rect 13105 4329 13139 4363
rect 13173 4329 13207 4363
rect 13241 4329 13275 4363
rect 13309 4329 13343 4363
rect 13377 4329 13390 4363
rect 12582 4293 13390 4329
rect 12582 4259 12595 4293
rect 12629 4259 12663 4293
rect 12697 4259 12731 4293
rect 12765 4259 12799 4293
rect 12833 4259 12867 4293
rect 12901 4259 12935 4293
rect 12969 4259 13003 4293
rect 13037 4259 13071 4293
rect 13105 4259 13139 4293
rect 13173 4259 13207 4293
rect 13241 4259 13275 4293
rect 13309 4259 13343 4293
rect 13377 4259 13390 4293
rect 12582 4223 13390 4259
rect 12582 4189 12595 4223
rect 12629 4189 12663 4223
rect 12697 4189 12731 4223
rect 12765 4189 12799 4223
rect 12833 4189 12867 4223
rect 12901 4189 12935 4223
rect 12969 4189 13003 4223
rect 13037 4189 13071 4223
rect 13105 4189 13139 4223
rect 13173 4189 13207 4223
rect 13241 4189 13275 4223
rect 13309 4189 13343 4223
rect 13377 4189 13390 4223
rect 12582 4153 13390 4189
rect 12582 4119 12595 4153
rect 12629 4119 12663 4153
rect 12697 4119 12731 4153
rect 12765 4119 12799 4153
rect 12833 4119 12867 4153
rect 12901 4119 12935 4153
rect 12969 4119 13003 4153
rect 13037 4119 13071 4153
rect 13105 4119 13139 4153
rect 13173 4119 13207 4153
rect 13241 4119 13275 4153
rect 13309 4119 13343 4153
rect 13377 4119 13390 4153
rect 12582 4083 13390 4119
rect 12582 4049 12595 4083
rect 12629 4049 12663 4083
rect 12697 4049 12731 4083
rect 12765 4049 12799 4083
rect 12833 4049 12867 4083
rect 12901 4049 12935 4083
rect 12969 4049 13003 4083
rect 13037 4049 13071 4083
rect 13105 4049 13139 4083
rect 13173 4049 13207 4083
rect 13241 4049 13275 4083
rect 13309 4049 13343 4083
rect 13377 4049 13390 4083
rect 12582 4013 13390 4049
rect 12582 3979 12595 4013
rect 12629 3979 12663 4013
rect 12697 3979 12731 4013
rect 12765 3979 12799 4013
rect 12833 3979 12867 4013
rect 12901 3979 12935 4013
rect 12969 3979 13003 4013
rect 13037 3979 13071 4013
rect 13105 3979 13139 4013
rect 13173 3979 13207 4013
rect 13241 3979 13275 4013
rect 13309 3979 13343 4013
rect 13377 3979 13390 4013
rect 12582 3943 13390 3979
rect 12582 3909 12595 3943
rect 12629 3909 12663 3943
rect 12697 3909 12731 3943
rect 12765 3909 12799 3943
rect 12833 3909 12867 3943
rect 12901 3909 12935 3943
rect 12969 3909 13003 3943
rect 13037 3909 13071 3943
rect 13105 3909 13139 3943
rect 13173 3909 13207 3943
rect 13241 3909 13275 3943
rect 13309 3909 13343 3943
rect 13377 3909 13390 3943
rect 12582 3873 13390 3909
rect 12582 3839 12595 3873
rect 12629 3839 12663 3873
rect 12697 3839 12731 3873
rect 12765 3839 12799 3873
rect 12833 3839 12867 3873
rect 12901 3839 12935 3873
rect 12969 3839 13003 3873
rect 13037 3839 13071 3873
rect 13105 3839 13139 3873
rect 13173 3839 13207 3873
rect 13241 3839 13275 3873
rect 13309 3839 13343 3873
rect 13377 3839 13390 3873
rect 12582 3803 13390 3839
rect 12582 3769 12595 3803
rect 12629 3769 12663 3803
rect 12697 3769 12731 3803
rect 12765 3769 12799 3803
rect 12833 3769 12867 3803
rect 12901 3769 12935 3803
rect 12969 3769 13003 3803
rect 13037 3769 13071 3803
rect 13105 3769 13139 3803
rect 13173 3769 13207 3803
rect 13241 3769 13275 3803
rect 13309 3769 13343 3803
rect 13377 3769 13390 3803
rect 12582 3733 13390 3769
rect 12582 3699 12595 3733
rect 12629 3699 12663 3733
rect 12697 3699 12731 3733
rect 12765 3699 12799 3733
rect 12833 3699 12867 3733
rect 12901 3699 12935 3733
rect 12969 3699 13003 3733
rect 13037 3699 13071 3733
rect 13105 3699 13139 3733
rect 13173 3699 13207 3733
rect 13241 3699 13275 3733
rect 13309 3699 13343 3733
rect 13377 3699 13390 3733
rect 12582 3663 13390 3699
rect 12582 3629 12595 3663
rect 12629 3629 12663 3663
rect 12697 3629 12731 3663
rect 12765 3629 12799 3663
rect 12833 3629 12867 3663
rect 12901 3629 12935 3663
rect 12969 3629 13003 3663
rect 13037 3629 13071 3663
rect 13105 3629 13139 3663
rect 13173 3629 13207 3663
rect 13241 3629 13275 3663
rect 13309 3629 13343 3663
rect 13377 3629 13390 3663
rect 12582 3593 13390 3629
rect 12582 3559 12595 3593
rect 12629 3559 12663 3593
rect 12697 3559 12731 3593
rect 12765 3559 12799 3593
rect 12833 3559 12867 3593
rect 12901 3559 12935 3593
rect 12969 3559 13003 3593
rect 13037 3559 13071 3593
rect 13105 3559 13139 3593
rect 13173 3559 13207 3593
rect 13241 3559 13275 3593
rect 13309 3559 13343 3593
rect 13377 3559 13390 3593
rect 12582 3523 13390 3559
rect 12582 3489 12595 3523
rect 12629 3489 12663 3523
rect 12697 3489 12731 3523
rect 12765 3489 12799 3523
rect 12833 3489 12867 3523
rect 12901 3489 12935 3523
rect 12969 3489 13003 3523
rect 13037 3489 13071 3523
rect 13105 3489 13139 3523
rect 13173 3489 13207 3523
rect 13241 3489 13275 3523
rect 13309 3489 13343 3523
rect 13377 3489 13390 3523
rect 12582 3453 13390 3489
rect 12582 3419 12595 3453
rect 12629 3419 12663 3453
rect 12697 3419 12731 3453
rect 12765 3419 12799 3453
rect 12833 3419 12867 3453
rect 12901 3419 12935 3453
rect 12969 3419 13003 3453
rect 13037 3419 13071 3453
rect 13105 3419 13139 3453
rect 13173 3419 13207 3453
rect 13241 3419 13275 3453
rect 13309 3419 13343 3453
rect 13377 3419 13390 3453
rect 12582 3383 13390 3419
rect 12582 3349 12595 3383
rect 12629 3349 12663 3383
rect 12697 3349 12731 3383
rect 12765 3349 12799 3383
rect 12833 3349 12867 3383
rect 12901 3349 12935 3383
rect 12969 3349 13003 3383
rect 13037 3349 13071 3383
rect 13105 3349 13139 3383
rect 13173 3349 13207 3383
rect 13241 3349 13275 3383
rect 13309 3349 13343 3383
rect 13377 3349 13390 3383
rect 12582 3313 13390 3349
rect 12582 3279 12595 3313
rect 12629 3279 12663 3313
rect 12697 3279 12731 3313
rect 12765 3279 12799 3313
rect 12833 3279 12867 3313
rect 12901 3279 12935 3313
rect 12969 3279 13003 3313
rect 13037 3279 13071 3313
rect 13105 3279 13139 3313
rect 13173 3279 13207 3313
rect 13241 3279 13275 3313
rect 13309 3279 13343 3313
rect 13377 3279 13390 3313
rect 12582 3243 13390 3279
rect 12582 3209 12595 3243
rect 12629 3209 12663 3243
rect 12697 3209 12731 3243
rect 12765 3209 12799 3243
rect 12833 3209 12867 3243
rect 12901 3209 12935 3243
rect 12969 3209 13003 3243
rect 13037 3209 13071 3243
rect 13105 3209 13139 3243
rect 13173 3209 13207 3243
rect 13241 3209 13275 3243
rect 13309 3209 13343 3243
rect 13377 3209 13390 3243
rect 12582 3173 13390 3209
rect 12582 3139 12595 3173
rect 12629 3139 12663 3173
rect 12697 3139 12731 3173
rect 12765 3139 12799 3173
rect 12833 3139 12867 3173
rect 12901 3139 12935 3173
rect 12969 3139 13003 3173
rect 13037 3139 13071 3173
rect 13105 3139 13139 3173
rect 13173 3139 13207 3173
rect 13241 3139 13275 3173
rect 13309 3139 13343 3173
rect 13377 3139 13390 3173
rect 12582 3103 13390 3139
rect 12582 3069 12595 3103
rect 12629 3069 12663 3103
rect 12697 3069 12731 3103
rect 12765 3069 12799 3103
rect 12833 3069 12867 3103
rect 12901 3069 12935 3103
rect 12969 3069 13003 3103
rect 13037 3069 13071 3103
rect 13105 3069 13139 3103
rect 13173 3069 13207 3103
rect 13241 3069 13275 3103
rect 13309 3069 13343 3103
rect 13377 3069 13390 3103
rect 12582 3033 13390 3069
rect 12582 2999 12595 3033
rect 12629 2999 12663 3033
rect 12697 2999 12731 3033
rect 12765 2999 12799 3033
rect 12833 2999 12867 3033
rect 12901 2999 12935 3033
rect 12969 2999 13003 3033
rect 13037 2999 13071 3033
rect 13105 2999 13139 3033
rect 13173 2999 13207 3033
rect 13241 2999 13275 3033
rect 13309 2999 13343 3033
rect 13377 2999 13390 3033
rect 12582 2964 13390 2999
rect 12582 2930 12595 2964
rect 12629 2930 12663 2964
rect 12697 2930 12731 2964
rect 12765 2930 12799 2964
rect 12833 2930 12867 2964
rect 12901 2930 12935 2964
rect 12969 2930 13003 2964
rect 13037 2930 13071 2964
rect 13105 2930 13139 2964
rect 13173 2930 13207 2964
rect 13241 2930 13275 2964
rect 13309 2930 13343 2964
rect 13377 2930 13390 2964
rect 12582 2895 13390 2930
rect 12582 2861 12595 2895
rect 12629 2861 12663 2895
rect 12697 2861 12731 2895
rect 12765 2861 12799 2895
rect 12833 2861 12867 2895
rect 12901 2861 12935 2895
rect 12969 2861 13003 2895
rect 13037 2861 13071 2895
rect 13105 2861 13139 2895
rect 13173 2861 13207 2895
rect 13241 2861 13275 2895
rect 13309 2861 13343 2895
rect 13377 2861 13390 2895
rect 12582 2826 13390 2861
rect 12582 2792 12595 2826
rect 12629 2792 12663 2826
rect 12697 2792 12731 2826
rect 12765 2792 12799 2826
rect 12833 2792 12867 2826
rect 12901 2792 12935 2826
rect 12969 2792 13003 2826
rect 13037 2792 13071 2826
rect 13105 2792 13139 2826
rect 13173 2792 13207 2826
rect 13241 2792 13275 2826
rect 13309 2792 13343 2826
rect 13377 2792 13390 2826
rect 12582 2757 13390 2792
rect 12582 2730 12595 2757
rect 11570 2727 12595 2730
rect 8643 2699 12595 2727
rect 13377 2730 13390 2757
rect 13377 2723 13458 2730
rect 8643 2692 11652 2699
rect 8677 2658 8711 2692
rect 8745 2658 8779 2692
rect 8813 2658 8847 2692
rect 8881 2658 8915 2692
rect 8949 2658 8983 2692
rect 9017 2658 9051 2692
rect 9085 2658 9119 2692
rect 9153 2658 9187 2692
rect 9221 2658 9255 2692
rect 9289 2658 9323 2692
rect 9357 2658 9391 2692
rect 9425 2658 9459 2692
rect 9493 2658 9527 2692
rect 9561 2658 9595 2692
rect 9629 2658 9663 2692
rect 9697 2658 9731 2692
rect 9765 2658 9799 2692
rect 9833 2658 9867 2692
rect 9901 2658 9935 2692
rect 9969 2658 10003 2692
rect 10037 2658 10071 2692
rect 10105 2658 10139 2692
rect 10173 2658 10207 2692
rect 10241 2658 10312 2692
rect 10346 2658 10380 2692
rect 10414 2658 10448 2692
rect 10482 2658 10516 2692
rect 10550 2658 10584 2692
rect 10618 2658 10652 2692
rect 10686 2658 10720 2692
rect 10754 2658 10788 2692
rect 10822 2658 10856 2692
rect 10890 2658 10924 2692
rect 10958 2658 10992 2692
rect 11026 2658 11060 2692
rect 11094 2658 11128 2692
rect 11162 2658 11196 2692
rect 11230 2658 11264 2692
rect 11298 2658 11332 2692
rect 11366 2658 11400 2692
rect 11434 2658 11468 2692
rect 11502 2658 11536 2692
rect 11570 2665 11652 2692
rect 11686 2665 11720 2699
rect 11754 2665 11788 2699
rect 11822 2665 11856 2699
rect 11890 2665 11924 2699
rect 11958 2665 11992 2699
rect 12026 2665 12060 2699
rect 12094 2665 12128 2699
rect 12162 2665 12196 2699
rect 12230 2665 12264 2699
rect 12298 2665 12332 2699
rect 12366 2665 12400 2699
rect 12434 2665 12468 2699
rect 12502 2689 12595 2699
rect 12502 2665 12573 2689
rect 11570 2658 12573 2665
rect 8643 2655 12573 2658
rect 13355 2655 13458 2723
rect 8643 2629 13458 2655
rect 8643 2623 11652 2629
rect 8677 2589 8711 2623
rect 8745 2589 8779 2623
rect 8813 2589 8847 2623
rect 8881 2589 8915 2623
rect 8949 2589 8983 2623
rect 9017 2589 9051 2623
rect 9085 2589 9119 2623
rect 9153 2589 9187 2623
rect 9221 2589 9255 2623
rect 9289 2589 9323 2623
rect 9357 2589 9391 2623
rect 9425 2589 9459 2623
rect 9493 2589 9527 2623
rect 9561 2589 9595 2623
rect 9629 2589 9663 2623
rect 9697 2589 9731 2623
rect 9765 2589 9799 2623
rect 9833 2589 9867 2623
rect 9901 2589 9935 2623
rect 9969 2589 10003 2623
rect 10037 2589 10071 2623
rect 10105 2589 10139 2623
rect 10173 2589 10207 2623
rect 10241 2589 10312 2623
rect 10346 2589 10380 2623
rect 10414 2589 10448 2623
rect 10482 2589 10516 2623
rect 10550 2589 10584 2623
rect 10618 2589 10652 2623
rect 10686 2589 10720 2623
rect 10754 2589 10788 2623
rect 10822 2589 10856 2623
rect 10890 2589 10924 2623
rect 10958 2589 10992 2623
rect 11026 2589 11060 2623
rect 11094 2589 11128 2623
rect 11162 2589 11196 2623
rect 11230 2589 11264 2623
rect 11298 2589 11332 2623
rect 11366 2589 11400 2623
rect 11434 2589 11468 2623
rect 11502 2589 11536 2623
rect 11570 2595 11652 2623
rect 11686 2595 11720 2629
rect 11754 2595 11788 2629
rect 11822 2595 11856 2629
rect 11890 2595 11924 2629
rect 11958 2595 11992 2629
rect 12026 2595 12060 2629
rect 12094 2595 12128 2629
rect 12162 2595 12196 2629
rect 12230 2595 12264 2629
rect 12298 2595 12332 2629
rect 12366 2595 12400 2629
rect 12434 2595 12468 2629
rect 12502 2620 13458 2629
rect 12502 2595 12573 2620
rect 11570 2589 12573 2595
rect 8643 2586 12573 2589
rect 12607 2586 12641 2620
rect 12675 2586 12709 2620
rect 12743 2586 12777 2620
rect 12811 2586 12845 2620
rect 12879 2586 12913 2620
rect 12947 2586 12981 2620
rect 13015 2586 13049 2620
rect 13083 2586 13117 2620
rect 13151 2586 13185 2620
rect 13219 2586 13253 2620
rect 13287 2586 13321 2620
rect 13355 2586 13458 2620
rect 8643 2559 13458 2586
rect 8643 2554 11652 2559
rect 8677 2520 8711 2554
rect 8745 2520 8779 2554
rect 8813 2520 8847 2554
rect 8881 2520 8915 2554
rect 8949 2520 8983 2554
rect 9017 2520 9051 2554
rect 9085 2520 9119 2554
rect 9153 2520 9187 2554
rect 9221 2520 9255 2554
rect 9289 2520 9323 2554
rect 9357 2520 9391 2554
rect 9425 2520 9459 2554
rect 9493 2520 9527 2554
rect 9561 2520 9595 2554
rect 9629 2520 9663 2554
rect 9697 2520 9731 2554
rect 9765 2520 9799 2554
rect 9833 2520 9867 2554
rect 9901 2520 9935 2554
rect 9969 2520 10003 2554
rect 10037 2520 10071 2554
rect 10105 2520 10139 2554
rect 10173 2520 10207 2554
rect 10241 2520 10312 2554
rect 10346 2520 10380 2554
rect 10414 2520 10448 2554
rect 10482 2520 10516 2554
rect 10550 2520 10584 2554
rect 10618 2520 10652 2554
rect 10686 2520 10720 2554
rect 10754 2520 10788 2554
rect 10822 2520 10856 2554
rect 10890 2520 10924 2554
rect 10958 2520 10992 2554
rect 11026 2520 11060 2554
rect 11094 2520 11128 2554
rect 11162 2520 11196 2554
rect 11230 2520 11264 2554
rect 11298 2520 11332 2554
rect 11366 2520 11400 2554
rect 11434 2520 11468 2554
rect 11502 2520 11536 2554
rect 11570 2525 11652 2554
rect 11686 2525 11720 2559
rect 11754 2525 11788 2559
rect 11822 2525 11856 2559
rect 11890 2525 11924 2559
rect 11958 2525 11992 2559
rect 12026 2525 12060 2559
rect 12094 2525 12128 2559
rect 12162 2525 12196 2559
rect 12230 2525 12264 2559
rect 12298 2525 12332 2559
rect 12366 2525 12400 2559
rect 12434 2525 12468 2559
rect 12502 2551 13458 2559
rect 12502 2525 12573 2551
rect 11570 2520 12573 2525
rect 8643 2517 12573 2520
rect 12607 2517 12641 2551
rect 12675 2517 12709 2551
rect 12743 2517 12777 2551
rect 12811 2517 12845 2551
rect 12879 2517 12913 2551
rect 12947 2517 12981 2551
rect 13015 2517 13049 2551
rect 13083 2517 13117 2551
rect 13151 2517 13185 2551
rect 13219 2517 13253 2551
rect 13287 2517 13321 2551
rect 13355 2517 13458 2551
rect 8643 2489 13458 2517
rect 8643 2485 11652 2489
rect 8677 2451 8711 2485
rect 8745 2451 8779 2485
rect 8813 2451 8847 2485
rect 8881 2451 8915 2485
rect 8949 2451 8983 2485
rect 9017 2451 9051 2485
rect 9085 2451 9119 2485
rect 9153 2451 9187 2485
rect 9221 2451 9255 2485
rect 9289 2451 9323 2485
rect 9357 2451 9391 2485
rect 9425 2451 9459 2485
rect 9493 2451 9527 2485
rect 9561 2451 9595 2485
rect 9629 2451 9663 2485
rect 9697 2451 9731 2485
rect 9765 2451 9799 2485
rect 9833 2451 9867 2485
rect 9901 2451 9935 2485
rect 9969 2451 10003 2485
rect 10037 2451 10071 2485
rect 10105 2451 10139 2485
rect 10173 2451 10207 2485
rect 10241 2451 10312 2485
rect 10346 2451 10380 2485
rect 10414 2451 10448 2485
rect 10482 2451 10516 2485
rect 10550 2451 10584 2485
rect 10618 2451 10652 2485
rect 10686 2451 10720 2485
rect 10754 2451 10788 2485
rect 10822 2451 10856 2485
rect 10890 2451 10924 2485
rect 10958 2451 10992 2485
rect 11026 2451 11060 2485
rect 11094 2451 11128 2485
rect 11162 2451 11196 2485
rect 11230 2451 11264 2485
rect 11298 2451 11332 2485
rect 11366 2451 11400 2485
rect 11434 2451 11468 2485
rect 11502 2451 11536 2485
rect 11570 2455 11652 2485
rect 11686 2455 11720 2489
rect 11754 2455 11788 2489
rect 11822 2455 11856 2489
rect 11890 2455 11924 2489
rect 11958 2455 11992 2489
rect 12026 2455 12060 2489
rect 12094 2455 12128 2489
rect 12162 2455 12196 2489
rect 12230 2455 12264 2489
rect 12298 2455 12332 2489
rect 12366 2455 12400 2489
rect 12434 2455 12468 2489
rect 12502 2482 13458 2489
rect 12502 2455 12573 2482
rect 11570 2451 12573 2455
rect 8643 2448 12573 2451
rect 12607 2448 12641 2482
rect 12675 2448 12709 2482
rect 12743 2448 12777 2482
rect 12811 2448 12845 2482
rect 12879 2448 12913 2482
rect 12947 2448 12981 2482
rect 13015 2448 13049 2482
rect 13083 2448 13117 2482
rect 13151 2448 13185 2482
rect 13219 2448 13253 2482
rect 13287 2448 13321 2482
rect 13355 2448 13458 2482
rect 8643 2419 13458 2448
rect 8643 2416 11652 2419
rect 8677 2382 8711 2416
rect 8745 2382 8779 2416
rect 8813 2382 8847 2416
rect 8881 2382 8915 2416
rect 8949 2382 8983 2416
rect 9017 2382 9051 2416
rect 9085 2382 9119 2416
rect 9153 2382 9187 2416
rect 9221 2382 9255 2416
rect 9289 2382 9323 2416
rect 9357 2382 9391 2416
rect 9425 2382 9459 2416
rect 9493 2382 9527 2416
rect 9561 2382 9595 2416
rect 9629 2382 9663 2416
rect 9697 2382 9731 2416
rect 9765 2382 9799 2416
rect 9833 2382 9867 2416
rect 9901 2382 9935 2416
rect 9969 2382 10003 2416
rect 10037 2382 10071 2416
rect 10105 2382 10139 2416
rect 10173 2382 10207 2416
rect 10241 2382 10312 2416
rect 10346 2382 10380 2416
rect 10414 2382 10448 2416
rect 10482 2382 10516 2416
rect 10550 2382 10584 2416
rect 10618 2382 10652 2416
rect 10686 2382 10720 2416
rect 10754 2382 10788 2416
rect 10822 2382 10856 2416
rect 10890 2382 10924 2416
rect 10958 2382 10992 2416
rect 11026 2382 11060 2416
rect 11094 2382 11128 2416
rect 11162 2382 11196 2416
rect 11230 2382 11264 2416
rect 11298 2382 11332 2416
rect 11366 2382 11400 2416
rect 11434 2382 11468 2416
rect 11502 2382 11536 2416
rect 11570 2385 11652 2416
rect 11686 2385 11720 2419
rect 11754 2385 11788 2419
rect 11822 2385 11856 2419
rect 11890 2385 11924 2419
rect 11958 2385 11992 2419
rect 12026 2385 12060 2419
rect 12094 2385 12128 2419
rect 12162 2385 12196 2419
rect 12230 2385 12264 2419
rect 12298 2385 12332 2419
rect 12366 2385 12400 2419
rect 12434 2385 12468 2419
rect 12502 2413 13458 2419
rect 12502 2385 12573 2413
rect 11570 2382 12573 2385
rect 8643 2379 12573 2382
rect 12607 2379 12641 2413
rect 12675 2379 12709 2413
rect 12743 2379 12777 2413
rect 12811 2379 12845 2413
rect 12879 2379 12913 2413
rect 12947 2379 12981 2413
rect 13015 2379 13049 2413
rect 13083 2379 13117 2413
rect 13151 2379 13185 2413
rect 13219 2379 13253 2413
rect 13287 2379 13321 2413
rect 13355 2379 13458 2413
rect 1460 2348 1740 2361
rect 1460 2337 1575 2348
rect 1460 2303 1507 2337
rect 1541 2314 1575 2337
rect 1609 2314 1643 2348
rect 1677 2327 1740 2348
rect 1774 2327 1809 2361
rect 1843 2327 1878 2361
rect 1912 2327 1947 2361
rect 1981 2327 2016 2361
rect 2050 2327 2085 2361
rect 2119 2327 2154 2361
rect 2188 2327 2223 2361
rect 2257 2327 2292 2361
rect 2326 2327 2361 2361
rect 2395 2327 2430 2361
rect 2464 2327 2499 2361
rect 2533 2327 2568 2361
rect 2602 2327 2637 2361
rect 2671 2327 2706 2361
rect 2740 2327 2775 2361
rect 2809 2327 2844 2361
rect 1677 2314 2844 2327
rect 1541 2303 2844 2314
rect 1460 2293 2844 2303
rect 1460 2279 1740 2293
rect 1460 2269 1575 2279
rect 1460 2235 1507 2269
rect 1541 2245 1575 2269
rect 1609 2245 1643 2279
rect 1677 2259 1740 2279
rect 1774 2259 1809 2293
rect 1843 2259 1878 2293
rect 1912 2259 1947 2293
rect 1981 2259 2016 2293
rect 2050 2259 2085 2293
rect 2119 2259 2154 2293
rect 2188 2259 2223 2293
rect 2257 2259 2292 2293
rect 2326 2259 2361 2293
rect 2395 2259 2430 2293
rect 2464 2259 2499 2293
rect 2533 2259 2568 2293
rect 2602 2259 2637 2293
rect 2671 2259 2706 2293
rect 2740 2259 2775 2293
rect 2809 2259 2844 2293
rect 1677 2245 2844 2259
rect 1541 2235 2844 2245
rect 1460 2225 2844 2235
rect 1460 2210 1740 2225
rect 1460 2201 1575 2210
rect 1460 2167 1507 2201
rect 1541 2176 1575 2201
rect 1609 2176 1643 2210
rect 1677 2191 1740 2210
rect 1774 2191 1809 2225
rect 1843 2191 1878 2225
rect 1912 2191 1947 2225
rect 1981 2191 2016 2225
rect 2050 2191 2085 2225
rect 2119 2191 2154 2225
rect 2188 2191 2223 2225
rect 2257 2191 2292 2225
rect 2326 2191 2361 2225
rect 2395 2191 2430 2225
rect 2464 2191 2499 2225
rect 2533 2191 2568 2225
rect 2602 2191 2637 2225
rect 2671 2191 2706 2225
rect 2740 2191 2775 2225
rect 2809 2191 2844 2225
rect 4782 2191 4806 2361
rect 8643 2349 13458 2379
rect 8643 2347 11652 2349
rect 8677 2313 8711 2347
rect 8745 2313 8779 2347
rect 8813 2313 8847 2347
rect 8881 2313 8915 2347
rect 8949 2313 8983 2347
rect 9017 2313 9051 2347
rect 9085 2313 9119 2347
rect 9153 2313 9187 2347
rect 9221 2313 9255 2347
rect 9289 2313 9323 2347
rect 9357 2313 9391 2347
rect 9425 2313 9459 2347
rect 9493 2313 9527 2347
rect 9561 2313 9595 2347
rect 9629 2313 9663 2347
rect 9697 2313 9731 2347
rect 9765 2313 9799 2347
rect 9833 2313 9867 2347
rect 9901 2313 9935 2347
rect 9969 2313 10003 2347
rect 10037 2313 10071 2347
rect 10105 2313 10139 2347
rect 10173 2313 10207 2347
rect 10241 2313 10312 2347
rect 10346 2313 10380 2347
rect 10414 2313 10448 2347
rect 10482 2313 10516 2347
rect 10550 2313 10584 2347
rect 10618 2313 10652 2347
rect 10686 2313 10720 2347
rect 10754 2313 10788 2347
rect 10822 2313 10856 2347
rect 10890 2313 10924 2347
rect 10958 2313 10992 2347
rect 11026 2313 11060 2347
rect 11094 2313 11128 2347
rect 11162 2313 11196 2347
rect 11230 2313 11264 2347
rect 11298 2313 11332 2347
rect 11366 2313 11400 2347
rect 11434 2313 11468 2347
rect 11502 2313 11536 2347
rect 11570 2315 11652 2347
rect 11686 2315 11720 2349
rect 11754 2315 11788 2349
rect 11822 2315 11856 2349
rect 11890 2315 11924 2349
rect 11958 2315 11992 2349
rect 12026 2315 12060 2349
rect 12094 2315 12128 2349
rect 12162 2315 12196 2349
rect 12230 2315 12264 2349
rect 12298 2315 12332 2349
rect 12366 2315 12400 2349
rect 12434 2315 12468 2349
rect 12502 2344 13458 2349
rect 12502 2315 12573 2344
rect 11570 2313 12573 2315
rect 8643 2310 12573 2313
rect 12607 2310 12641 2344
rect 12675 2310 12709 2344
rect 12743 2310 12777 2344
rect 12811 2310 12845 2344
rect 12879 2310 12913 2344
rect 12947 2310 12981 2344
rect 13015 2310 13049 2344
rect 13083 2310 13117 2344
rect 13151 2310 13185 2344
rect 13219 2310 13253 2344
rect 13287 2310 13321 2344
rect 13355 2310 13458 2344
rect 8643 2279 13458 2310
rect 8643 2278 11652 2279
rect 8677 2244 8711 2278
rect 8745 2244 8779 2278
rect 8813 2244 8847 2278
rect 8881 2244 8915 2278
rect 8949 2244 8983 2278
rect 9017 2244 9051 2278
rect 9085 2244 9119 2278
rect 9153 2244 9187 2278
rect 9221 2244 9255 2278
rect 9289 2244 9323 2278
rect 9357 2244 9391 2278
rect 9425 2244 9459 2278
rect 9493 2244 9527 2278
rect 9561 2244 9595 2278
rect 9629 2244 9663 2278
rect 9697 2244 9731 2278
rect 9765 2244 9799 2278
rect 9833 2244 9867 2278
rect 9901 2244 9935 2278
rect 9969 2244 10003 2278
rect 10037 2244 10071 2278
rect 10105 2244 10139 2278
rect 10173 2244 10207 2278
rect 10241 2244 10312 2278
rect 10346 2244 10380 2278
rect 10414 2244 10448 2278
rect 10482 2244 10516 2278
rect 10550 2244 10584 2278
rect 10618 2244 10652 2278
rect 10686 2244 10720 2278
rect 10754 2244 10788 2278
rect 10822 2244 10856 2278
rect 10890 2244 10924 2278
rect 10958 2244 10992 2278
rect 11026 2244 11060 2278
rect 11094 2244 11128 2278
rect 11162 2244 11196 2278
rect 11230 2244 11264 2278
rect 11298 2244 11332 2278
rect 11366 2244 11400 2278
rect 11434 2244 11468 2278
rect 11502 2244 11536 2278
rect 11570 2245 11652 2278
rect 11686 2245 11720 2279
rect 11754 2245 11788 2279
rect 11822 2245 11856 2279
rect 11890 2245 11924 2279
rect 11958 2245 11992 2279
rect 12026 2245 12060 2279
rect 12094 2245 12128 2279
rect 12162 2245 12196 2279
rect 12230 2245 12264 2279
rect 12298 2245 12332 2279
rect 12366 2245 12400 2279
rect 12434 2245 12468 2279
rect 12502 2275 13458 2279
rect 12502 2245 12573 2275
rect 11570 2244 12573 2245
rect 8643 2241 12573 2244
rect 12607 2241 12641 2275
rect 12675 2241 12709 2275
rect 12743 2241 12777 2275
rect 12811 2241 12845 2275
rect 12879 2241 12913 2275
rect 12947 2241 12981 2275
rect 13015 2241 13049 2275
rect 13083 2241 13117 2275
rect 13151 2241 13185 2275
rect 13219 2241 13253 2275
rect 13287 2241 13321 2275
rect 13355 2241 13458 2275
rect 8643 2209 13458 2241
rect 1541 2167 1677 2176
rect 1460 2141 1677 2167
rect 1460 2133 1575 2141
rect 1460 2099 1507 2133
rect 1541 2107 1575 2133
rect 1609 2107 1643 2141
rect 1541 2099 1677 2107
rect 1460 2072 1677 2099
rect 1460 2065 1575 2072
rect 1460 2031 1507 2065
rect 1541 2038 1575 2065
rect 1609 2038 1643 2072
rect 1541 2031 1677 2038
rect 1460 2003 1677 2031
rect 1460 1997 1575 2003
rect 1460 1963 1507 1997
rect 1541 1969 1575 1997
rect 1609 1969 1643 2003
rect 1541 1963 1677 1969
rect 1460 1934 1677 1963
rect 1460 1929 1575 1934
rect 1460 1895 1507 1929
rect 1541 1900 1575 1929
rect 1609 1900 1643 1934
rect 1541 1895 1677 1900
rect 1460 1865 1677 1895
rect 1460 1861 1575 1865
rect 1460 1827 1507 1861
rect 1541 1831 1575 1861
rect 1609 1831 1643 1865
rect 1541 1827 1677 1831
rect 1460 1796 1677 1827
rect 1460 1793 1575 1796
rect 1460 1759 1507 1793
rect 1541 1762 1575 1793
rect 1609 1762 1643 1796
rect 1541 1759 1677 1762
rect 1460 1727 1677 1759
rect 1460 1725 1575 1727
rect 1460 1691 1507 1725
rect 1541 1693 1575 1725
rect 1609 1693 1643 1727
rect 1541 1691 1677 1693
rect 1460 1658 1677 1691
rect 1460 1657 1575 1658
rect 1460 1623 1507 1657
rect 1541 1624 1575 1657
rect 1609 1624 1643 1658
rect 1541 1623 1677 1624
rect 1460 1589 1677 1623
rect 8677 2175 8711 2209
rect 8745 2175 8779 2209
rect 8813 2175 8847 2209
rect 8881 2175 8915 2209
rect 8949 2175 8983 2209
rect 9017 2175 9051 2209
rect 9085 2175 9119 2209
rect 9153 2175 9187 2209
rect 9221 2175 9255 2209
rect 9289 2175 9323 2209
rect 9357 2175 9391 2209
rect 9425 2175 9459 2209
rect 9493 2175 9527 2209
rect 9561 2175 9595 2209
rect 9629 2175 9663 2209
rect 9697 2175 9731 2209
rect 9765 2175 9799 2209
rect 9833 2175 9867 2209
rect 9901 2175 9935 2209
rect 9969 2175 10003 2209
rect 10037 2175 10071 2209
rect 10105 2175 10139 2209
rect 10173 2175 10207 2209
rect 10241 2175 10312 2209
rect 10346 2175 10380 2209
rect 10414 2175 10448 2209
rect 10482 2175 10516 2209
rect 10550 2175 10584 2209
rect 10618 2175 10652 2209
rect 10686 2175 10720 2209
rect 10754 2175 10788 2209
rect 10822 2175 10856 2209
rect 10890 2175 10924 2209
rect 10958 2175 10992 2209
rect 11026 2175 11060 2209
rect 11094 2175 11128 2209
rect 11162 2175 11196 2209
rect 11230 2175 11264 2209
rect 11298 2175 11332 2209
rect 11366 2175 11400 2209
rect 11434 2175 11468 2209
rect 11502 2175 11536 2209
rect 11570 2175 11652 2209
rect 11686 2175 11720 2209
rect 11754 2175 11788 2209
rect 11822 2175 11856 2209
rect 11890 2175 11924 2209
rect 11958 2175 11992 2209
rect 12026 2175 12060 2209
rect 12094 2175 12128 2209
rect 12162 2175 12196 2209
rect 12230 2175 12264 2209
rect 12298 2175 12332 2209
rect 12366 2175 12400 2209
rect 12434 2175 12468 2209
rect 12502 2206 13458 2209
rect 12502 2175 12573 2206
rect 8643 2172 12573 2175
rect 12607 2172 12641 2206
rect 12675 2172 12709 2206
rect 12743 2172 12777 2206
rect 12811 2172 12845 2206
rect 12879 2172 12913 2206
rect 12947 2172 12981 2206
rect 13015 2172 13049 2206
rect 13083 2172 13117 2206
rect 13151 2172 13185 2206
rect 13219 2172 13253 2206
rect 13287 2172 13321 2206
rect 13355 2172 13458 2206
rect 8643 2140 13458 2172
rect 8677 2106 8711 2140
rect 8745 2106 8779 2140
rect 8813 2106 8847 2140
rect 8881 2106 8915 2140
rect 8949 2106 8983 2140
rect 9017 2106 9051 2140
rect 9085 2106 9119 2140
rect 9153 2106 9187 2140
rect 9221 2106 9255 2140
rect 9289 2106 9323 2140
rect 9357 2106 9391 2140
rect 9425 2106 9459 2140
rect 9493 2106 9527 2140
rect 9561 2106 9595 2140
rect 9629 2106 9663 2140
rect 9697 2106 9731 2140
rect 9765 2106 9799 2140
rect 9833 2106 9867 2140
rect 9901 2106 9935 2140
rect 9969 2106 10003 2140
rect 10037 2106 10071 2140
rect 10105 2106 10139 2140
rect 10173 2106 10207 2140
rect 10241 2106 10312 2140
rect 10346 2106 10380 2140
rect 10414 2106 10448 2140
rect 10482 2106 10516 2140
rect 10550 2106 10584 2140
rect 10618 2106 10652 2140
rect 10686 2106 10720 2140
rect 10754 2106 10788 2140
rect 10822 2106 10856 2140
rect 10890 2106 10924 2140
rect 10958 2106 10992 2140
rect 11026 2106 11060 2140
rect 11094 2106 11128 2140
rect 11162 2106 11196 2140
rect 11230 2106 11264 2140
rect 11298 2106 11332 2140
rect 11366 2106 11400 2140
rect 11434 2106 11468 2140
rect 11502 2106 11536 2140
rect 11570 2106 11652 2140
rect 11686 2106 11720 2140
rect 11754 2106 11788 2140
rect 11822 2106 11856 2140
rect 11890 2106 11924 2140
rect 11958 2106 11992 2140
rect 12026 2106 12060 2140
rect 12094 2106 12128 2140
rect 12162 2106 12196 2140
rect 12230 2106 12264 2140
rect 12298 2106 12332 2140
rect 12366 2106 12400 2140
rect 12434 2106 12468 2140
rect 12502 2137 13458 2140
rect 12502 2106 12573 2137
rect 8643 2103 12573 2106
rect 12607 2103 12641 2137
rect 12675 2103 12709 2137
rect 12743 2103 12777 2137
rect 12811 2103 12845 2137
rect 12879 2103 12913 2137
rect 12947 2103 12981 2137
rect 13015 2103 13049 2137
rect 13083 2103 13117 2137
rect 13151 2103 13185 2137
rect 13219 2103 13253 2137
rect 13287 2103 13321 2137
rect 13355 2103 13458 2137
rect 8643 2071 13458 2103
rect 8677 2037 8711 2071
rect 8745 2037 8779 2071
rect 8813 2037 8847 2071
rect 8881 2037 8915 2071
rect 8949 2037 8983 2071
rect 9017 2037 9051 2071
rect 9085 2037 9119 2071
rect 9153 2037 9187 2071
rect 9221 2037 9255 2071
rect 9289 2037 9323 2071
rect 9357 2037 9391 2071
rect 9425 2037 9459 2071
rect 9493 2037 9527 2071
rect 9561 2037 9595 2071
rect 9629 2037 9663 2071
rect 9697 2037 9731 2071
rect 9765 2037 9799 2071
rect 9833 2037 9867 2071
rect 9901 2037 9935 2071
rect 9969 2037 10003 2071
rect 10037 2037 10071 2071
rect 10105 2037 10139 2071
rect 10173 2037 10207 2071
rect 10241 2037 10312 2071
rect 10346 2037 10380 2071
rect 10414 2037 10448 2071
rect 10482 2037 10516 2071
rect 10550 2037 10584 2071
rect 10618 2037 10652 2071
rect 10686 2037 10720 2071
rect 10754 2037 10788 2071
rect 10822 2037 10856 2071
rect 10890 2037 10924 2071
rect 10958 2037 10992 2071
rect 11026 2037 11060 2071
rect 11094 2037 11128 2071
rect 11162 2037 11196 2071
rect 11230 2037 11264 2071
rect 11298 2037 11332 2071
rect 11366 2037 11400 2071
rect 11434 2037 11468 2071
rect 11502 2037 11536 2071
rect 11570 2037 11652 2071
rect 11686 2037 11720 2071
rect 11754 2037 11788 2071
rect 11822 2037 11856 2071
rect 11890 2037 11924 2071
rect 11958 2037 11992 2071
rect 12026 2037 12060 2071
rect 12094 2037 12128 2071
rect 12162 2037 12196 2071
rect 12230 2037 12264 2071
rect 12298 2037 12332 2071
rect 12366 2037 12400 2071
rect 12434 2037 12468 2071
rect 12502 2068 13458 2071
rect 12502 2037 12573 2068
rect 8643 2034 12573 2037
rect 12607 2034 12641 2068
rect 12675 2034 12709 2068
rect 12743 2034 12777 2068
rect 12811 2034 12845 2068
rect 12879 2034 12913 2068
rect 12947 2034 12981 2068
rect 13015 2034 13049 2068
rect 13083 2034 13117 2068
rect 13151 2034 13185 2068
rect 13219 2034 13253 2068
rect 13287 2034 13321 2068
rect 13355 2034 13458 2068
rect 8643 2002 13458 2034
rect 8677 1968 8711 2002
rect 8745 1968 8779 2002
rect 8813 1968 8847 2002
rect 8881 1968 8915 2002
rect 8949 1968 8983 2002
rect 9017 1968 9051 2002
rect 9085 1968 9119 2002
rect 9153 1968 9187 2002
rect 9221 1968 9255 2002
rect 9289 1968 9323 2002
rect 9357 1968 9391 2002
rect 9425 1968 9459 2002
rect 9493 1968 9527 2002
rect 9561 1968 9595 2002
rect 9629 1968 9663 2002
rect 9697 1968 9731 2002
rect 9765 1968 9799 2002
rect 9833 1968 9867 2002
rect 9901 1968 9935 2002
rect 9969 1968 10003 2002
rect 10037 1968 10071 2002
rect 10105 1968 10139 2002
rect 10173 1968 10207 2002
rect 10241 1968 10312 2002
rect 10346 1968 10380 2002
rect 10414 1968 10448 2002
rect 10482 1968 10516 2002
rect 10550 1968 10584 2002
rect 10618 1968 10652 2002
rect 10686 1968 10720 2002
rect 10754 1968 10788 2002
rect 10822 1968 10856 2002
rect 10890 1968 10924 2002
rect 10958 1968 10992 2002
rect 11026 1968 11060 2002
rect 11094 1968 11128 2002
rect 11162 1968 11196 2002
rect 11230 1968 11264 2002
rect 11298 1968 11332 2002
rect 11366 1968 11400 2002
rect 11434 1968 11468 2002
rect 11502 1968 11536 2002
rect 11570 1968 11652 2002
rect 11686 1968 11720 2002
rect 11754 1968 11788 2002
rect 11822 1968 11856 2002
rect 11890 1968 11924 2002
rect 11958 1968 11992 2002
rect 12026 1968 12060 2002
rect 12094 1968 12128 2002
rect 12162 1968 12196 2002
rect 12230 1968 12264 2002
rect 12298 1968 12332 2002
rect 12366 1968 12400 2002
rect 12434 1968 12468 2002
rect 12502 1999 13458 2002
rect 12502 1968 12573 1999
rect 8643 1965 12573 1968
rect 12607 1965 12641 1999
rect 12675 1965 12709 1999
rect 12743 1965 12777 1999
rect 12811 1965 12845 1999
rect 12879 1965 12913 1999
rect 12947 1965 12981 1999
rect 13015 1965 13049 1999
rect 13083 1965 13117 1999
rect 13151 1965 13185 1999
rect 13219 1965 13253 1999
rect 13287 1965 13321 1999
rect 13355 1965 13458 1999
rect 8643 1933 13458 1965
rect 8677 1899 8711 1933
rect 8745 1899 8779 1933
rect 8813 1899 8847 1933
rect 8881 1899 8915 1933
rect 8949 1899 8983 1933
rect 9017 1899 9051 1933
rect 9085 1899 9119 1933
rect 9153 1899 9187 1933
rect 9221 1899 9255 1933
rect 9289 1899 9323 1933
rect 9357 1899 9391 1933
rect 9425 1899 9459 1933
rect 9493 1899 9527 1933
rect 9561 1899 9595 1933
rect 9629 1899 9663 1933
rect 9697 1899 9731 1933
rect 9765 1899 9799 1933
rect 9833 1899 9867 1933
rect 9901 1899 9935 1933
rect 9969 1899 10003 1933
rect 10037 1899 10071 1933
rect 10105 1899 10139 1933
rect 10173 1899 10207 1933
rect 10241 1899 10312 1933
rect 10346 1899 10380 1933
rect 10414 1899 10448 1933
rect 10482 1899 10516 1933
rect 10550 1899 10584 1933
rect 10618 1899 10652 1933
rect 10686 1899 10720 1933
rect 10754 1899 10788 1933
rect 10822 1899 10856 1933
rect 10890 1899 10924 1933
rect 10958 1899 10992 1933
rect 11026 1899 11060 1933
rect 11094 1899 11128 1933
rect 11162 1899 11196 1933
rect 11230 1899 11264 1933
rect 11298 1899 11332 1933
rect 11366 1899 11400 1933
rect 11434 1899 11468 1933
rect 11502 1899 11536 1933
rect 11570 1899 11652 1933
rect 11686 1899 11720 1933
rect 11754 1899 11788 1933
rect 11822 1899 11856 1933
rect 11890 1899 11924 1933
rect 11958 1899 11992 1933
rect 12026 1899 12060 1933
rect 12094 1899 12128 1933
rect 12162 1899 12196 1933
rect 12230 1899 12264 1933
rect 12298 1899 12332 1933
rect 12366 1899 12400 1933
rect 12434 1899 12468 1933
rect 12502 1930 13458 1933
rect 12502 1899 12573 1930
rect 8643 1896 12573 1899
rect 12607 1896 12641 1930
rect 12675 1896 12709 1930
rect 12743 1896 12777 1930
rect 12811 1896 12845 1930
rect 12879 1896 12913 1930
rect 12947 1896 12981 1930
rect 13015 1896 13049 1930
rect 13083 1896 13117 1930
rect 13151 1896 13185 1930
rect 13219 1896 13253 1930
rect 13287 1896 13321 1930
rect 13355 1896 13458 1930
rect 8643 1864 13458 1896
rect 8677 1830 8711 1864
rect 8745 1830 8779 1864
rect 8813 1830 8847 1864
rect 8881 1830 8915 1864
rect 8949 1830 8983 1864
rect 9017 1830 9051 1864
rect 9085 1830 9119 1864
rect 9153 1830 9187 1864
rect 9221 1830 9255 1864
rect 9289 1830 9323 1864
rect 9357 1830 9391 1864
rect 9425 1830 9459 1864
rect 9493 1830 9527 1864
rect 9561 1830 9595 1864
rect 9629 1830 9663 1864
rect 9697 1830 9731 1864
rect 9765 1830 9799 1864
rect 9833 1830 9867 1864
rect 9901 1830 9935 1864
rect 9969 1830 10003 1864
rect 10037 1830 10071 1864
rect 10105 1830 10139 1864
rect 10173 1830 10207 1864
rect 10241 1830 10312 1864
rect 10346 1830 10380 1864
rect 10414 1830 10448 1864
rect 10482 1830 10516 1864
rect 10550 1830 10584 1864
rect 10618 1830 10652 1864
rect 10686 1830 10720 1864
rect 10754 1830 10788 1864
rect 10822 1830 10856 1864
rect 10890 1830 10924 1864
rect 10958 1830 10992 1864
rect 11026 1830 11060 1864
rect 11094 1830 11128 1864
rect 11162 1830 11196 1864
rect 11230 1830 11264 1864
rect 11298 1830 11332 1864
rect 11366 1830 11400 1864
rect 11434 1830 11468 1864
rect 11502 1830 11536 1864
rect 11570 1830 11652 1864
rect 11686 1830 11720 1864
rect 11754 1830 11788 1864
rect 11822 1830 11856 1864
rect 11890 1830 11924 1864
rect 11958 1830 11992 1864
rect 12026 1830 12060 1864
rect 12094 1830 12128 1864
rect 12162 1830 12196 1864
rect 12230 1830 12264 1864
rect 12298 1830 12332 1864
rect 12366 1830 12400 1864
rect 12434 1830 12468 1864
rect 12502 1861 13458 1864
rect 12502 1830 12573 1861
rect 8643 1795 12573 1830
rect 8677 1761 8711 1795
rect 8745 1761 8779 1795
rect 8813 1761 8847 1795
rect 8881 1761 8915 1795
rect 8949 1761 8983 1795
rect 9017 1761 9051 1795
rect 9085 1761 9119 1795
rect 9153 1761 9187 1795
rect 9221 1761 9255 1795
rect 9289 1761 9323 1795
rect 9357 1761 9391 1795
rect 9425 1761 9459 1795
rect 9493 1761 9527 1795
rect 9561 1761 9595 1795
rect 9629 1761 9663 1795
rect 9697 1761 9731 1795
rect 9765 1761 9799 1795
rect 9833 1761 9867 1795
rect 9901 1761 9935 1795
rect 9969 1761 10003 1795
rect 10037 1761 10071 1795
rect 10105 1761 10139 1795
rect 10173 1761 10207 1795
rect 10241 1761 10312 1795
rect 10346 1761 10380 1795
rect 10414 1761 10448 1795
rect 10482 1761 10516 1795
rect 10550 1761 10584 1795
rect 10618 1761 10652 1795
rect 10686 1761 10720 1795
rect 10754 1761 10788 1795
rect 10822 1761 10856 1795
rect 10890 1761 10924 1795
rect 10958 1761 10992 1795
rect 11026 1761 11060 1795
rect 11094 1761 11128 1795
rect 11162 1761 11196 1795
rect 11230 1761 11264 1795
rect 11298 1761 11332 1795
rect 11366 1761 11400 1795
rect 11434 1761 11468 1795
rect 11502 1761 11536 1795
rect 11570 1761 11652 1795
rect 11686 1761 11720 1795
rect 11754 1761 11788 1795
rect 11822 1761 11856 1795
rect 11890 1761 11924 1795
rect 11958 1761 11992 1795
rect 12026 1761 12060 1795
rect 12094 1761 12128 1795
rect 12162 1761 12196 1795
rect 12230 1761 12264 1795
rect 12298 1761 12332 1795
rect 12366 1761 12400 1795
rect 12434 1761 12468 1795
rect 12502 1761 12573 1795
rect 8643 1726 12573 1761
rect 8677 1692 8711 1726
rect 8745 1692 8779 1726
rect 8813 1692 8847 1726
rect 8881 1692 8915 1726
rect 8949 1692 8983 1726
rect 9017 1692 9051 1726
rect 9085 1692 9119 1726
rect 9153 1692 9187 1726
rect 9221 1692 9255 1726
rect 9289 1692 9323 1726
rect 9357 1692 9391 1726
rect 9425 1692 9459 1726
rect 9493 1692 9527 1726
rect 9561 1692 9595 1726
rect 9629 1692 9663 1726
rect 9697 1692 9731 1726
rect 9765 1692 9799 1726
rect 9833 1692 9867 1726
rect 9901 1692 9935 1726
rect 9969 1692 10003 1726
rect 10037 1692 10071 1726
rect 10105 1692 10139 1726
rect 10173 1692 10207 1726
rect 10241 1692 10312 1726
rect 10346 1692 10380 1726
rect 10414 1692 10448 1726
rect 10482 1692 10516 1726
rect 10550 1692 10584 1726
rect 10618 1692 10652 1726
rect 10686 1692 10720 1726
rect 10754 1692 10788 1726
rect 10822 1692 10856 1726
rect 10890 1692 10924 1726
rect 10958 1692 10992 1726
rect 11026 1692 11060 1726
rect 11094 1692 11128 1726
rect 11162 1692 11196 1726
rect 11230 1692 11264 1726
rect 11298 1692 11332 1726
rect 11366 1692 11400 1726
rect 11434 1692 11468 1726
rect 11502 1692 11536 1726
rect 11570 1692 11652 1726
rect 11686 1692 11720 1726
rect 11754 1692 11788 1726
rect 11822 1692 11856 1726
rect 11890 1692 11924 1726
rect 11958 1692 11992 1726
rect 12026 1692 12060 1726
rect 12094 1692 12128 1726
rect 12162 1692 12196 1726
rect 12230 1692 12264 1726
rect 12298 1692 12332 1726
rect 12366 1692 12400 1726
rect 12434 1692 12468 1726
rect 12502 1692 12573 1726
rect 8643 1657 12573 1692
rect 8677 1623 8711 1657
rect 8745 1623 8779 1657
rect 8813 1623 8847 1657
rect 8881 1623 8915 1657
rect 8949 1623 8983 1657
rect 9017 1623 9051 1657
rect 9085 1623 9119 1657
rect 9153 1623 9187 1657
rect 9221 1623 9255 1657
rect 9289 1623 9323 1657
rect 9357 1623 9391 1657
rect 9425 1623 9459 1657
rect 9493 1623 9527 1657
rect 9561 1623 9595 1657
rect 9629 1623 9663 1657
rect 9697 1623 9731 1657
rect 9765 1623 9799 1657
rect 9833 1623 9867 1657
rect 9901 1623 9935 1657
rect 9969 1623 10003 1657
rect 10037 1623 10071 1657
rect 10105 1623 10139 1657
rect 10173 1623 10207 1657
rect 10241 1623 10312 1657
rect 10346 1623 10380 1657
rect 10414 1623 10448 1657
rect 10482 1623 10516 1657
rect 10550 1623 10584 1657
rect 10618 1623 10652 1657
rect 10686 1623 10720 1657
rect 10754 1623 10788 1657
rect 10822 1623 10856 1657
rect 10890 1623 10924 1657
rect 10958 1623 10992 1657
rect 11026 1623 11060 1657
rect 11094 1623 11128 1657
rect 11162 1623 11196 1657
rect 11230 1623 11264 1657
rect 11298 1623 11332 1657
rect 11366 1623 11400 1657
rect 11434 1623 11468 1657
rect 11502 1623 11536 1657
rect 11570 1623 11652 1657
rect 11686 1623 11720 1657
rect 11754 1623 11788 1657
rect 11822 1623 11856 1657
rect 11890 1623 11924 1657
rect 11958 1623 11992 1657
rect 12026 1623 12060 1657
rect 12094 1623 12128 1657
rect 12162 1623 12196 1657
rect 12230 1623 12264 1657
rect 12298 1623 12332 1657
rect 12366 1623 12400 1657
rect 12434 1623 12468 1657
rect 12502 1623 12573 1657
rect 13355 1623 13458 1861
rect 8643 1589 13458 1623
rect 1460 1555 1507 1589
rect 1541 1555 1575 1589
rect 1609 1555 1643 1589
rect 1460 1521 1677 1555
rect 8388 1555 8412 1589
rect 8446 1555 8482 1589
rect 8516 1555 8552 1589
rect 8586 1555 8622 1589
rect 8656 1555 8692 1589
rect 8726 1555 8762 1589
rect 8796 1555 8832 1589
rect 8866 1555 8902 1589
rect 8936 1555 8972 1589
rect 9006 1555 9043 1589
rect 9077 1555 9114 1589
rect 9148 1555 9185 1589
rect 9219 1555 9256 1589
rect 9290 1555 9327 1589
rect 9361 1555 9398 1589
rect 9432 1555 9469 1589
rect 9503 1555 9540 1589
rect 9574 1555 9611 1589
rect 9645 1555 9682 1589
rect 9716 1555 9753 1589
rect 9787 1555 9824 1589
rect 9858 1555 9895 1589
rect 9929 1555 9966 1589
rect 10000 1583 13458 1589
rect 10000 1555 10024 1583
rect 8388 1521 10024 1555
rect 1460 1487 1531 1521
rect 1565 1487 1600 1521
rect 1634 1487 1669 1521
rect 1703 1487 1738 1521
rect 1772 1487 1807 1521
rect 1841 1487 1876 1521
rect 1910 1487 1945 1521
rect 1979 1487 2014 1521
rect 2048 1487 2083 1521
rect 2117 1487 2152 1521
rect 2186 1487 2221 1521
rect 2255 1487 2290 1521
rect 2324 1487 2359 1521
rect 2393 1487 2428 1521
rect 2462 1487 2497 1521
rect 2531 1487 2566 1521
rect 2600 1487 2635 1521
rect 2669 1487 2704 1521
rect 2738 1487 2773 1521
rect 2807 1487 2842 1521
rect 2876 1487 2911 1521
rect 2945 1487 2980 1521
rect 3014 1487 3049 1521
rect 3083 1487 3118 1521
rect 3152 1487 3187 1521
rect 3221 1487 3256 1521
rect 3290 1487 3325 1521
rect 3359 1487 3394 1521
rect 3428 1487 3463 1521
rect 3497 1487 3532 1521
rect 3566 1487 3601 1521
rect 3635 1487 3670 1521
rect 3704 1487 3739 1521
rect 3773 1487 3808 1521
rect 3842 1487 3877 1521
rect 3911 1487 3946 1521
rect 3980 1487 4015 1521
rect 4049 1487 4084 1521
rect 4118 1487 4153 1521
rect 4187 1487 4222 1521
rect 4256 1487 4291 1521
rect 4325 1487 4360 1521
rect 4394 1487 4429 1521
rect 4463 1487 4498 1521
rect 4532 1487 4567 1521
rect 4601 1487 4636 1521
rect 4670 1487 4705 1521
rect 4739 1487 4774 1521
rect 4808 1487 4843 1521
rect 4877 1487 4912 1521
rect 4946 1487 4981 1521
rect 5015 1487 5050 1521
rect 5084 1487 5119 1521
rect 5153 1487 5188 1521
rect 5222 1487 5257 1521
rect 5291 1487 5326 1521
rect 5360 1487 5395 1521
rect 5429 1487 5464 1521
rect 5498 1487 5533 1521
rect 5567 1487 5602 1521
rect 5636 1487 5671 1521
rect 5705 1487 5740 1521
rect 5774 1487 5809 1521
rect 5843 1487 5878 1521
rect 5912 1487 5947 1521
rect 5981 1487 6016 1521
rect 6050 1487 6085 1521
rect 6119 1487 6154 1521
rect 1460 1453 6154 1487
rect 1460 1443 1531 1453
rect 1086 1419 1531 1443
rect 1565 1419 1600 1453
rect 1634 1419 1669 1453
rect 1703 1419 1738 1453
rect 1772 1419 1807 1453
rect 1841 1419 1876 1453
rect 1910 1419 1945 1453
rect 1979 1419 2014 1453
rect 2048 1419 2083 1453
rect 2117 1419 2152 1453
rect 2186 1419 2221 1453
rect 2255 1419 2290 1453
rect 2324 1419 2359 1453
rect 2393 1419 2428 1453
rect 2462 1419 2497 1453
rect 2531 1419 2566 1453
rect 2600 1419 2635 1453
rect 2669 1419 2704 1453
rect 2738 1419 2773 1453
rect 2807 1419 2842 1453
rect 2876 1419 2911 1453
rect 2945 1419 2980 1453
rect 3014 1419 3049 1453
rect 3083 1419 3118 1453
rect 3152 1419 3187 1453
rect 3221 1419 3256 1453
rect 3290 1419 3325 1453
rect 3359 1419 3394 1453
rect 3428 1419 3463 1453
rect 3497 1419 3532 1453
rect 3566 1419 3601 1453
rect 3635 1419 3670 1453
rect 3704 1419 3739 1453
rect 3773 1419 3808 1453
rect 3842 1419 3877 1453
rect 3911 1419 3946 1453
rect 3980 1419 4015 1453
rect 4049 1419 4084 1453
rect 4118 1419 4153 1453
rect 4187 1419 4222 1453
rect 4256 1419 4291 1453
rect 4325 1419 4360 1453
rect 4394 1419 4429 1453
rect 4463 1419 4498 1453
rect 4532 1419 4567 1453
rect 4601 1419 4636 1453
rect 4670 1419 4705 1453
rect 4739 1419 4774 1453
rect 4808 1419 4843 1453
rect 4877 1419 4912 1453
rect 4946 1419 4981 1453
rect 5015 1419 5050 1453
rect 5084 1419 5119 1453
rect 5153 1419 5188 1453
rect 5222 1419 5257 1453
rect 5291 1419 5326 1453
rect 5360 1419 5395 1453
rect 5429 1419 5464 1453
rect 5498 1419 5533 1453
rect 5567 1419 5602 1453
rect 5636 1419 5671 1453
rect 5705 1419 5740 1453
rect 5774 1419 5809 1453
rect 5843 1419 5878 1453
rect 5912 1419 5947 1453
rect 5981 1419 6016 1453
rect 6050 1419 6085 1453
rect 6119 1419 6154 1453
rect 8364 1487 8412 1521
rect 8446 1487 8482 1521
rect 8516 1487 8552 1521
rect 8586 1487 8622 1521
rect 8656 1487 8692 1521
rect 8726 1487 8762 1521
rect 8796 1487 8832 1521
rect 8866 1487 8902 1521
rect 8936 1487 8972 1521
rect 9006 1487 9043 1521
rect 9077 1487 9114 1521
rect 9148 1487 9185 1521
rect 9219 1487 9256 1521
rect 9290 1487 9327 1521
rect 9361 1487 9398 1521
rect 9432 1487 9469 1521
rect 9503 1487 9540 1521
rect 9574 1487 9611 1521
rect 9645 1487 9682 1521
rect 9716 1487 9753 1521
rect 9787 1487 9824 1521
rect 9858 1487 9895 1521
rect 9929 1487 9966 1521
rect 10000 1487 10024 1521
rect 8364 1453 10024 1487
rect 8364 1419 8412 1453
rect 8446 1419 8482 1453
rect 8516 1419 8552 1453
rect 8586 1419 8622 1453
rect 8656 1419 8692 1453
rect 8726 1419 8762 1453
rect 8796 1419 8832 1453
rect 8866 1419 8902 1453
rect 8936 1419 8972 1453
rect 9006 1419 9043 1453
rect 9077 1419 9114 1453
rect 9148 1419 9185 1453
rect 9219 1419 9256 1453
rect 9290 1419 9327 1453
rect 9361 1419 9398 1453
rect 9432 1419 9469 1453
rect 9503 1419 9540 1453
rect 9574 1419 9611 1453
rect 9645 1419 9682 1453
rect 9716 1419 9753 1453
rect 9787 1419 9824 1453
rect 9858 1419 9895 1453
rect 9929 1419 9966 1453
rect 10000 1419 10024 1453
rect 24119 5522 24540 5532
rect 24119 5488 24153 5522
rect 24187 5488 24221 5522
rect 24255 5488 24289 5522
rect 24323 5488 24357 5522
rect 24391 5488 24425 5522
rect 24459 5488 24493 5522
rect 24527 5488 24540 5522
rect 24119 5453 24540 5488
rect 24119 5419 24153 5453
rect 24187 5419 24221 5453
rect 24255 5419 24289 5453
rect 24323 5419 24357 5453
rect 24391 5419 24425 5453
rect 24459 5419 24493 5453
rect 24527 5419 24540 5453
rect 24119 5384 24540 5419
rect 24119 5350 24153 5384
rect 24187 5350 24221 5384
rect 24255 5350 24289 5384
rect 24323 5350 24357 5384
rect 24391 5350 24425 5384
rect 24459 5350 24493 5384
rect 24527 5350 24540 5384
rect 24119 5315 24540 5350
rect 24119 5281 24153 5315
rect 24187 5281 24221 5315
rect 24255 5281 24289 5315
rect 24323 5281 24357 5315
rect 24391 5281 24425 5315
rect 24459 5281 24493 5315
rect 24527 5281 24540 5315
rect 24119 5246 24540 5281
rect 24119 5212 24153 5246
rect 24187 5212 24221 5246
rect 24255 5212 24289 5246
rect 24323 5212 24357 5246
rect 24391 5212 24425 5246
rect 24459 5212 24493 5246
rect 24527 5212 24540 5246
rect 24119 5177 24540 5212
rect 24119 5143 24153 5177
rect 24187 5143 24221 5177
rect 24255 5143 24289 5177
rect 24323 5143 24357 5177
rect 24391 5143 24425 5177
rect 24459 5143 24493 5177
rect 24527 5143 24540 5177
rect 24119 5108 24540 5143
rect 24119 5074 24153 5108
rect 24187 5074 24221 5108
rect 24255 5074 24289 5108
rect 24323 5074 24357 5108
rect 24391 5074 24425 5108
rect 24459 5074 24493 5108
rect 24527 5074 24540 5108
rect 24119 5039 24540 5074
rect 24119 5005 24153 5039
rect 24187 5005 24221 5039
rect 24255 5005 24289 5039
rect 24323 5005 24357 5039
rect 24391 5005 24425 5039
rect 24459 5005 24493 5039
rect 24527 5005 24540 5039
rect 24119 4970 24540 5005
rect 24119 4936 24153 4970
rect 24187 4936 24221 4970
rect 24255 4936 24289 4970
rect 24323 4936 24357 4970
rect 24391 4936 24425 4970
rect 24459 4936 24493 4970
rect 24527 4936 24540 4970
rect 24119 4901 24540 4936
rect 24119 4867 24153 4901
rect 24187 4867 24221 4901
rect 24255 4867 24289 4901
rect 24323 4867 24357 4901
rect 24391 4867 24425 4901
rect 24459 4867 24493 4901
rect 24527 4867 24540 4901
rect 24119 4832 24540 4867
rect 24119 4798 24153 4832
rect 24187 4798 24221 4832
rect 24255 4798 24289 4832
rect 24323 4798 24357 4832
rect 24391 4798 24425 4832
rect 24459 4798 24493 4832
rect 24527 4798 24540 4832
rect 24119 4763 24540 4798
rect 24119 4729 24153 4763
rect 24187 4729 24221 4763
rect 24255 4729 24289 4763
rect 24323 4729 24357 4763
rect 24391 4729 24425 4763
rect 24459 4729 24493 4763
rect 24527 4729 24540 4763
rect 24119 4694 24540 4729
rect 24527 2348 24540 4694
rect 24119 2324 24540 2348
rect 20507 942 20558 976
rect 20592 942 20627 976
rect 20661 942 20696 976
rect 20730 942 20765 976
rect 20799 942 20834 976
rect 20868 942 20903 976
rect 20937 942 20972 976
rect 21006 942 21041 976
rect 21075 942 21110 976
rect 21144 942 21179 976
rect 21213 942 21248 976
rect 21282 942 21317 976
rect 21351 942 21386 976
rect 21420 942 21455 976
rect 21489 942 21524 976
rect 21558 942 21593 976
rect 21627 942 21662 976
rect 21696 942 21731 976
rect 21765 942 21800 976
rect 21834 942 21869 976
rect 21903 942 21938 976
rect 21972 942 22007 976
rect 22041 942 22076 976
rect 22110 942 22145 976
rect 22179 942 22214 976
rect 22248 942 22283 976
rect 22317 942 22352 976
rect 22386 942 22421 976
rect 22455 942 22490 976
rect 22524 942 22559 976
rect 22593 942 22628 976
rect 22662 942 22697 976
rect 22731 942 22766 976
rect 22800 942 22835 976
rect 22869 942 22904 976
rect 22938 942 22973 976
rect 20507 908 22973 942
rect 20507 874 20558 908
rect 20592 874 20627 908
rect 20661 874 20696 908
rect 20730 874 20765 908
rect 20799 874 20834 908
rect 20868 874 20903 908
rect 20937 874 20972 908
rect 21006 874 21041 908
rect 21075 874 21110 908
rect 21144 874 21179 908
rect 21213 874 21248 908
rect 21282 874 21317 908
rect 21351 874 21386 908
rect 21420 874 21455 908
rect 21489 874 21524 908
rect 21558 874 21593 908
rect 21627 874 21662 908
rect 21696 874 21731 908
rect 21765 874 21800 908
rect 21834 874 21869 908
rect 21903 874 21938 908
rect 21972 874 22007 908
rect 22041 874 22076 908
rect 22110 874 22145 908
rect 22179 874 22214 908
rect 22248 874 22283 908
rect 22317 874 22352 908
rect 22386 874 22421 908
rect 22455 874 22490 908
rect 22524 874 22559 908
rect 22593 874 22628 908
rect 22662 874 22697 908
rect 22731 874 22766 908
rect 22800 874 22835 908
rect 22869 874 22904 908
rect 22938 874 22973 908
rect 278 822 448 857
rect 312 788 346 822
rect 380 788 414 822
rect 20507 840 22973 874
rect 20507 806 20558 840
rect 20592 806 20627 840
rect 20661 806 20696 840
rect 20730 806 20765 840
rect 20799 806 20834 840
rect 20868 806 20903 840
rect 20937 806 20972 840
rect 21006 806 21041 840
rect 21075 806 21110 840
rect 21144 806 21179 840
rect 21213 806 21248 840
rect 21282 806 21317 840
rect 21351 806 21386 840
rect 21420 806 21455 840
rect 21489 806 21524 840
rect 21558 806 21593 840
rect 21627 806 21662 840
rect 21696 806 21731 840
rect 21765 806 21800 840
rect 21834 806 21869 840
rect 21903 806 21938 840
rect 21972 806 22007 840
rect 22041 806 22076 840
rect 22110 806 22145 840
rect 22179 806 22214 840
rect 22248 806 22283 840
rect 22317 806 22352 840
rect 22386 806 22421 840
rect 22455 806 22490 840
rect 22524 806 22559 840
rect 22593 806 22628 840
rect 22662 806 22697 840
rect 22731 806 22766 840
rect 22800 806 22835 840
rect 22869 806 22904 840
rect 22938 806 22973 840
rect 24095 806 24119 1010
rect 278 753 448 788
rect 312 719 346 753
rect 380 719 414 753
rect 278 684 448 719
rect 312 650 346 684
rect 380 650 414 684
rect 278 615 448 650
rect 312 581 346 615
rect 380 581 414 615
rect 278 546 448 581
rect 312 512 346 546
rect 380 512 414 546
rect 278 477 448 512
rect 312 443 346 477
rect 380 443 414 477
rect 278 408 448 443
rect 312 374 346 408
rect 380 374 414 408
rect 278 339 448 374
rect 312 305 346 339
rect 380 305 414 339
rect 278 270 448 305
rect 312 236 346 270
rect 380 236 414 270
rect 278 201 448 236
rect 312 167 346 201
rect 380 167 414 201
rect 278 133 448 167
<< mvpsubdiffcont >>
rect 22818 9261 22852 9295
rect 22886 9261 22920 9295
rect 22954 9261 22988 9295
rect 23022 9261 23056 9295
rect 23090 9261 23124 9295
rect 23158 9261 23192 9295
rect 23226 9261 23260 9295
rect 23294 9261 23328 9295
rect 23362 9261 23396 9295
rect 23430 9261 23464 9295
rect 23498 9261 23532 9295
rect 23566 9261 23600 9295
rect 23638 9284 23672 9318
rect 23706 9284 23740 9318
rect 23774 9284 23808 9318
rect 23842 9284 23876 9318
rect 23910 9284 23944 9318
rect 23978 9284 24012 9318
rect 24046 9284 24080 9318
rect 24114 9284 24148 9318
rect 22818 9192 22852 9226
rect 22886 9192 22920 9226
rect 22954 9192 22988 9226
rect 23022 9192 23056 9226
rect 23090 9192 23124 9226
rect 23158 9192 23192 9226
rect 23226 9192 23260 9226
rect 23294 9192 23328 9226
rect 23362 9192 23396 9226
rect 23430 9192 23464 9226
rect 23498 9192 23532 9226
rect 23566 9192 23600 9226
rect 23638 9211 23672 9245
rect 23706 9211 23740 9245
rect 23774 9211 23808 9245
rect 23842 9211 23876 9245
rect 23910 9211 23944 9245
rect 23978 9211 24012 9245
rect 24046 9211 24080 9245
rect 24114 9211 24148 9245
rect 22818 9123 22852 9157
rect 22886 9123 22920 9157
rect 22954 9123 22988 9157
rect 23022 9123 23056 9157
rect 23090 9123 23124 9157
rect 23158 9123 23192 9157
rect 23226 9123 23260 9157
rect 23294 9123 23328 9157
rect 23362 9123 23396 9157
rect 23430 9123 23464 9157
rect 23498 9123 23532 9157
rect 23566 9123 23600 9157
rect 23638 9138 23672 9172
rect 23706 9138 23740 9172
rect 23774 9138 23808 9172
rect 23842 9138 23876 9172
rect 23910 9138 23944 9172
rect 23978 9138 24012 9172
rect 24046 9138 24080 9172
rect 24114 9138 24148 9172
rect 22818 9054 22852 9088
rect 22886 9054 22920 9088
rect 22954 9054 22988 9088
rect 23022 9054 23056 9088
rect 23090 9054 23124 9088
rect 23158 9054 23192 9088
rect 23226 9054 23260 9088
rect 23294 9054 23328 9088
rect 23362 9054 23396 9088
rect 23430 9054 23464 9088
rect 23498 9054 23532 9088
rect 23566 9054 23600 9088
rect 23638 9065 23672 9099
rect 23706 9065 23740 9099
rect 23774 9065 23808 9099
rect 23842 9065 23876 9099
rect 23910 9065 23944 9099
rect 23978 9065 24012 9099
rect 24046 9065 24080 9099
rect 24114 9065 24148 9099
rect 22818 8985 22852 9019
rect 22886 8985 22920 9019
rect 22954 8985 22988 9019
rect 23022 8985 23056 9019
rect 23090 8985 23124 9019
rect 23158 8985 23192 9019
rect 23226 8985 23260 9019
rect 23294 8985 23328 9019
rect 23362 8985 23396 9019
rect 23430 8985 23464 9019
rect 23498 8985 23532 9019
rect 23566 8985 23600 9019
rect 23638 8991 23672 9025
rect 23706 8991 23740 9025
rect 23774 8991 23808 9025
rect 23842 8991 23876 9025
rect 23910 8991 23944 9025
rect 23978 8991 24012 9025
rect 24046 8991 24080 9025
rect 24114 8991 24148 9025
rect 22818 8916 22852 8950
rect 22886 8916 22920 8950
rect 22954 8916 22988 8950
rect 23022 8916 23056 8950
rect 23090 8916 23124 8950
rect 23158 8916 23192 8950
rect 23226 8916 23260 8950
rect 23294 8916 23328 8950
rect 23362 8916 23396 8950
rect 23430 8916 23464 8950
rect 23498 8916 23532 8950
rect 23566 8916 23600 8950
rect 23638 8917 23672 8951
rect 23706 8917 23740 8951
rect 23774 8917 23808 8951
rect 23842 8917 23876 8951
rect 23910 8917 23944 8951
rect 23978 8917 24012 8951
rect 24046 8917 24080 8951
rect 24114 8917 24148 8951
rect 22818 8847 22852 8881
rect 22886 8847 22920 8881
rect 22954 8847 22988 8881
rect 23022 8847 23056 8881
rect 23090 8847 23124 8881
rect 23158 8847 23192 8881
rect 23226 8847 23260 8881
rect 23294 8847 23328 8881
rect 23362 8847 23396 8881
rect 23430 8847 23464 8881
rect 23498 8847 23532 8881
rect 23566 8847 23600 8881
rect 23638 8843 23672 8877
rect 23706 8843 23740 8877
rect 23774 8843 23808 8877
rect 23842 8843 23876 8877
rect 23910 8843 23944 8877
rect 23978 8843 24012 8877
rect 24046 8843 24080 8877
rect 24114 8843 24148 8877
rect 22818 8778 22852 8812
rect 22886 8778 22920 8812
rect 22954 8778 22988 8812
rect 23022 8778 23056 8812
rect 23090 8778 23124 8812
rect 23158 8778 23192 8812
rect 23226 8778 23260 8812
rect 23294 8778 23328 8812
rect 23362 8778 23396 8812
rect 23430 8778 23464 8812
rect 23498 8778 23532 8812
rect 23566 8778 23600 8812
rect 23638 8769 23672 8803
rect 23706 8769 23740 8803
rect 23774 8769 23808 8803
rect 23842 8769 23876 8803
rect 23910 8769 23944 8803
rect 23978 8769 24012 8803
rect 24046 8769 24080 8803
rect 24114 8769 24148 8803
rect 22818 8709 22852 8743
rect 22886 8709 22920 8743
rect 22954 8709 22988 8743
rect 23022 8709 23056 8743
rect 23090 8709 23124 8743
rect 23158 8709 23192 8743
rect 23226 8709 23260 8743
rect 23294 8709 23328 8743
rect 23362 8709 23396 8743
rect 23430 8709 23464 8743
rect 23498 8709 23532 8743
rect 23566 8709 23600 8743
rect 22818 8640 22852 8674
rect 22886 8640 22920 8674
rect 22954 8640 22988 8674
rect 23022 8640 23056 8674
rect 23090 8640 23124 8674
rect 23158 8640 23192 8674
rect 23226 8640 23260 8674
rect 23294 8640 23328 8674
rect 23362 8640 23396 8674
rect 23430 8640 23464 8674
rect 23498 8640 23532 8674
rect 23566 8640 23600 8674
rect 22818 8571 22852 8605
rect 22886 8571 22920 8605
rect 22954 8571 22988 8605
rect 23022 8571 23056 8605
rect 23090 8571 23124 8605
rect 23158 8571 23192 8605
rect 23226 8571 23260 8605
rect 23294 8571 23328 8605
rect 23362 8571 23396 8605
rect 23430 8571 23464 8605
rect 23498 8571 23532 8605
rect 23566 8571 23600 8605
rect 22818 8502 22852 8536
rect 22886 8502 22920 8536
rect 22954 8502 22988 8536
rect 23022 8502 23056 8536
rect 23090 8502 23124 8536
rect 23158 8502 23192 8536
rect 23226 8502 23260 8536
rect 23294 8502 23328 8536
rect 23362 8502 23396 8536
rect 23430 8502 23464 8536
rect 23498 8502 23532 8536
rect 23566 8502 23600 8536
rect 22818 8433 22852 8467
rect 22886 8433 22920 8467
rect 22954 8433 22988 8467
rect 23022 8433 23056 8467
rect 23090 8433 23124 8467
rect 23158 8433 23192 8467
rect 23226 8433 23260 8467
rect 23294 8433 23328 8467
rect 23362 8433 23396 8467
rect 23430 8433 23464 8467
rect 23498 8433 23532 8467
rect 23566 8433 23600 8467
rect 22818 8364 22852 8398
rect 22886 8364 22920 8398
rect 22954 8364 22988 8398
rect 23022 8364 23056 8398
rect 23090 8364 23124 8398
rect 23158 8364 23192 8398
rect 23226 8364 23260 8398
rect 23294 8364 23328 8398
rect 23362 8364 23396 8398
rect 23430 8364 23464 8398
rect 23498 8364 23532 8398
rect 23566 8364 23600 8398
rect 22818 8295 22852 8329
rect 22886 8295 22920 8329
rect 22954 8295 22988 8329
rect 23022 8295 23056 8329
rect 23090 8295 23124 8329
rect 23158 8295 23192 8329
rect 23226 8295 23260 8329
rect 23294 8295 23328 8329
rect 23362 8295 23396 8329
rect 23430 8295 23464 8329
rect 23498 8295 23532 8329
rect 23566 8295 23600 8329
rect 22818 8226 22852 8260
rect 22886 8226 22920 8260
rect 22954 8226 22988 8260
rect 23022 8226 23056 8260
rect 23090 8226 23124 8260
rect 23158 8226 23192 8260
rect 23226 8226 23260 8260
rect 23294 8226 23328 8260
rect 23362 8226 23396 8260
rect 23430 8226 23464 8260
rect 23498 8226 23532 8260
rect 23566 8226 23600 8260
rect 22818 8157 22852 8191
rect 22886 8157 22920 8191
rect 22954 8157 22988 8191
rect 23022 8157 23056 8191
rect 23090 8157 23124 8191
rect 23158 8157 23192 8191
rect 23226 8157 23260 8191
rect 23294 8157 23328 8191
rect 23362 8157 23396 8191
rect 23430 8157 23464 8191
rect 23498 8157 23532 8191
rect 23566 8157 23600 8191
rect 22818 8088 22852 8122
rect 22886 8088 22920 8122
rect 22954 8088 22988 8122
rect 23022 8088 23056 8122
rect 23090 8088 23124 8122
rect 23158 8088 23192 8122
rect 23226 8088 23260 8122
rect 23294 8088 23328 8122
rect 23362 8088 23396 8122
rect 23430 8088 23464 8122
rect 23498 8088 23532 8122
rect 23566 8088 23600 8122
rect 22818 8019 22852 8053
rect 22886 8019 22920 8053
rect 22954 8019 22988 8053
rect 23022 8019 23056 8053
rect 23090 8019 23124 8053
rect 23158 8019 23192 8053
rect 23226 8019 23260 8053
rect 23294 8019 23328 8053
rect 23362 8019 23396 8053
rect 23430 8019 23464 8053
rect 23498 8019 23532 8053
rect 23566 8019 23600 8053
rect 22818 7950 22852 7984
rect 22886 7950 22920 7984
rect 22954 7950 22988 7984
rect 23022 7950 23056 7984
rect 23090 7950 23124 7984
rect 23158 7950 23192 7984
rect 23226 7950 23260 7984
rect 23294 7950 23328 7984
rect 23362 7950 23396 7984
rect 23430 7950 23464 7984
rect 23498 7950 23532 7984
rect 23566 7950 23600 7984
rect 22818 7881 22852 7915
rect 22886 7881 22920 7915
rect 22954 7881 22988 7915
rect 23022 7881 23056 7915
rect 23090 7881 23124 7915
rect 23158 7881 23192 7915
rect 23226 7881 23260 7915
rect 23294 7881 23328 7915
rect 23362 7881 23396 7915
rect 23430 7881 23464 7915
rect 23498 7881 23532 7915
rect 23566 7881 23600 7915
rect 22818 7812 22852 7846
rect 22886 7812 22920 7846
rect 22954 7812 22988 7846
rect 23022 7812 23056 7846
rect 23090 7812 23124 7846
rect 23158 7812 23192 7846
rect 23226 7812 23260 7846
rect 23294 7812 23328 7846
rect 23362 7812 23396 7846
rect 23430 7812 23464 7846
rect 23498 7812 23532 7846
rect 23566 7812 23600 7846
rect 22818 7743 22852 7777
rect 22886 7743 22920 7777
rect 22954 7743 22988 7777
rect 23022 7743 23056 7777
rect 23090 7743 23124 7777
rect 23158 7743 23192 7777
rect 23226 7743 23260 7777
rect 23294 7743 23328 7777
rect 23362 7743 23396 7777
rect 23430 7743 23464 7777
rect 23498 7743 23532 7777
rect 23566 7743 23600 7777
rect 22818 7674 22852 7708
rect 22886 7674 22920 7708
rect 22954 7674 22988 7708
rect 23022 7674 23056 7708
rect 23090 7674 23124 7708
rect 23158 7674 23192 7708
rect 23226 7674 23260 7708
rect 23294 7674 23328 7708
rect 23362 7674 23396 7708
rect 23430 7674 23464 7708
rect 23498 7674 23532 7708
rect 23566 7674 23600 7708
rect 22818 7605 22852 7639
rect 22886 7605 22920 7639
rect 22954 7605 22988 7639
rect 23022 7605 23056 7639
rect 23090 7605 23124 7639
rect 23158 7605 23192 7639
rect 23226 7605 23260 7639
rect 23294 7605 23328 7639
rect 23362 7605 23396 7639
rect 23430 7605 23464 7639
rect 23498 7605 23532 7639
rect 23566 7605 23600 7639
rect 22818 7536 22852 7570
rect 22886 7536 22920 7570
rect 22954 7536 22988 7570
rect 23022 7536 23056 7570
rect 23090 7536 23124 7570
rect 23158 7536 23192 7570
rect 23226 7536 23260 7570
rect 23294 7536 23328 7570
rect 23362 7536 23396 7570
rect 23430 7536 23464 7570
rect 23498 7536 23532 7570
rect 23566 7536 23600 7570
rect 22818 7467 22852 7501
rect 22886 7467 22920 7501
rect 22954 7467 22988 7501
rect 23022 7467 23056 7501
rect 23090 7467 23124 7501
rect 23158 7467 23192 7501
rect 23226 7467 23260 7501
rect 23294 7467 23328 7501
rect 23362 7467 23396 7501
rect 23430 7467 23464 7501
rect 23498 7467 23532 7501
rect 23566 7467 23600 7501
rect 22818 7398 22852 7432
rect 22886 7398 22920 7432
rect 22954 7398 22988 7432
rect 23022 7398 23056 7432
rect 23090 7398 23124 7432
rect 23158 7398 23192 7432
rect 23226 7398 23260 7432
rect 23294 7398 23328 7432
rect 23362 7398 23396 7432
rect 23430 7398 23464 7432
rect 23498 7398 23532 7432
rect 23566 7398 23600 7432
rect 22818 7329 22852 7363
rect 22886 7329 22920 7363
rect 22954 7329 22988 7363
rect 23022 7329 23056 7363
rect 23090 7329 23124 7363
rect 23158 7329 23192 7363
rect 23226 7329 23260 7363
rect 23294 7329 23328 7363
rect 23362 7329 23396 7363
rect 23430 7329 23464 7363
rect 23498 7329 23532 7363
rect 23566 7329 23600 7363
rect 22818 7260 22852 7294
rect 22886 7260 22920 7294
rect 22954 7260 22988 7294
rect 23022 7260 23056 7294
rect 23090 7260 23124 7294
rect 23158 7260 23192 7294
rect 23226 7260 23260 7294
rect 23294 7260 23328 7294
rect 23362 7260 23396 7294
rect 23430 7260 23464 7294
rect 23498 7260 23532 7294
rect 23566 7260 23600 7294
rect 22818 7191 22852 7225
rect 22886 7191 22920 7225
rect 22954 7191 22988 7225
rect 23022 7191 23056 7225
rect 23090 7191 23124 7225
rect 23158 7191 23192 7225
rect 23226 7191 23260 7225
rect 23294 7191 23328 7225
rect 23362 7191 23396 7225
rect 23430 7191 23464 7225
rect 23498 7191 23532 7225
rect 23566 7191 23600 7225
rect 22818 7122 22852 7156
rect 22886 7122 22920 7156
rect 22954 7122 22988 7156
rect 23022 7122 23056 7156
rect 23090 7122 23124 7156
rect 23158 7122 23192 7156
rect 23226 7122 23260 7156
rect 23294 7122 23328 7156
rect 23362 7122 23396 7156
rect 23430 7122 23464 7156
rect 23498 7122 23532 7156
rect 23566 7122 23600 7156
rect 22818 7053 22852 7087
rect 22886 7053 22920 7087
rect 22954 7053 22988 7087
rect 23022 7053 23056 7087
rect 23090 7053 23124 7087
rect 23158 7053 23192 7087
rect 23226 7053 23260 7087
rect 23294 7053 23328 7087
rect 23362 7053 23396 7087
rect 23430 7053 23464 7087
rect 23498 7053 23532 7087
rect 23566 7053 23600 7087
rect 22818 6984 22852 7018
rect 22886 6984 22920 7018
rect 22954 6984 22988 7018
rect 23022 6984 23056 7018
rect 23090 6984 23124 7018
rect 23158 6984 23192 7018
rect 23226 6984 23260 7018
rect 23294 6984 23328 7018
rect 23362 6984 23396 7018
rect 23430 6984 23464 7018
rect 23498 6984 23532 7018
rect 23566 6984 23600 7018
rect 22818 6915 22852 6949
rect 22886 6915 22920 6949
rect 22954 6915 22988 6949
rect 23022 6915 23056 6949
rect 23090 6915 23124 6949
rect 23158 6915 23192 6949
rect 23226 6915 23260 6949
rect 23294 6915 23328 6949
rect 23362 6915 23396 6949
rect 23430 6915 23464 6949
rect 23498 6915 23532 6949
rect 23566 6915 23600 6949
rect 22818 6846 22852 6880
rect 22886 6846 22920 6880
rect 22954 6846 22988 6880
rect 23022 6846 23056 6880
rect 23090 6846 23124 6880
rect 23158 6846 23192 6880
rect 23226 6846 23260 6880
rect 23294 6846 23328 6880
rect 23362 6846 23396 6880
rect 23430 6846 23464 6880
rect 23498 6846 23532 6880
rect 23566 6846 23600 6880
rect 22818 5485 23600 6811
rect 22842 4794 22944 5440
rect 22979 5406 23013 5440
rect 23048 5406 23082 5440
rect 23117 5406 23151 5440
rect 23186 5406 23220 5440
rect 23255 5406 23289 5440
rect 23324 5406 23358 5440
rect 23393 5406 23427 5440
rect 23462 5406 23496 5440
rect 23531 5406 23565 5440
rect 23600 5406 23634 5440
rect 23669 5406 23703 5440
rect 23738 5406 23772 5440
rect 22979 5338 23013 5372
rect 23048 5338 23082 5372
rect 23117 5338 23151 5372
rect 23186 5338 23220 5372
rect 23255 5338 23289 5372
rect 23324 5338 23358 5372
rect 23393 5338 23427 5372
rect 23462 5338 23496 5372
rect 23531 5338 23565 5372
rect 23600 5338 23634 5372
rect 23669 5338 23703 5372
rect 23738 5338 23772 5372
rect 22979 5270 23013 5304
rect 23048 5270 23082 5304
rect 23117 5270 23151 5304
rect 23186 5270 23220 5304
rect 23255 5270 23289 5304
rect 23324 5270 23358 5304
rect 23393 5270 23427 5304
rect 23462 5270 23496 5304
rect 23531 5270 23565 5304
rect 23600 5270 23634 5304
rect 23669 5270 23703 5304
rect 23738 5270 23772 5304
rect 22979 5202 23013 5236
rect 23048 5202 23082 5236
rect 23117 5202 23151 5236
rect 23186 5202 23220 5236
rect 23255 5202 23289 5236
rect 23324 5202 23358 5236
rect 23393 5202 23427 5236
rect 23462 5202 23496 5236
rect 23531 5202 23565 5236
rect 23600 5202 23634 5236
rect 23669 5202 23703 5236
rect 23738 5202 23772 5236
rect 22979 5134 23013 5168
rect 23048 5134 23082 5168
rect 23117 5134 23151 5168
rect 23186 5134 23220 5168
rect 23255 5134 23289 5168
rect 23324 5134 23358 5168
rect 23393 5134 23427 5168
rect 23462 5134 23496 5168
rect 23531 5134 23565 5168
rect 23600 5134 23634 5168
rect 23669 5134 23703 5168
rect 23738 5134 23772 5168
rect 22979 5066 23013 5100
rect 23048 5066 23082 5100
rect 23117 5066 23151 5100
rect 23186 5066 23220 5100
rect 23255 5066 23289 5100
rect 23324 5066 23358 5100
rect 23393 5066 23427 5100
rect 23462 5066 23496 5100
rect 23531 5066 23565 5100
rect 23600 5066 23634 5100
rect 23669 5066 23703 5100
rect 23738 5066 23772 5100
rect 22979 4998 23013 5032
rect 23048 4998 23082 5032
rect 23117 4998 23151 5032
rect 23186 4998 23220 5032
rect 23255 4998 23289 5032
rect 23324 4998 23358 5032
rect 23393 4998 23427 5032
rect 23462 4998 23496 5032
rect 23531 4998 23565 5032
rect 23600 4998 23634 5032
rect 23669 4998 23703 5032
rect 23738 4998 23772 5032
rect 22979 4930 23013 4964
rect 23048 4930 23082 4964
rect 23117 4930 23151 4964
rect 23186 4930 23220 4964
rect 23255 4930 23289 4964
rect 23324 4930 23358 4964
rect 23393 4930 23427 4964
rect 23462 4930 23496 4964
rect 23531 4930 23565 4964
rect 23600 4930 23634 4964
rect 23669 4930 23703 4964
rect 23738 4930 23772 4964
rect 22979 4862 23013 4896
rect 23048 4862 23082 4896
rect 23117 4862 23151 4896
rect 23186 4862 23220 4896
rect 23255 4862 23289 4896
rect 23324 4862 23358 4896
rect 23393 4862 23427 4896
rect 23462 4862 23496 4896
rect 23531 4862 23565 4896
rect 23600 4862 23634 4896
rect 23669 4862 23703 4896
rect 23738 4862 23772 4896
rect 22979 4794 23013 4828
rect 23048 4794 23082 4828
rect 23117 4794 23151 4828
rect 23186 4794 23220 4828
rect 23255 4794 23289 4828
rect 23324 4794 23358 4828
rect 23393 4794 23427 4828
rect 23462 4794 23496 4828
rect 23531 4794 23565 4828
rect 23600 4794 23634 4828
rect 23669 4794 23703 4828
rect 23738 4794 23772 4828
rect 696 4703 730 4737
rect 764 4703 798 4737
rect 832 4703 866 4737
rect 696 4631 730 4665
rect 764 4631 798 4665
rect 832 4631 866 4665
rect 696 4559 730 4593
rect 764 4559 798 4593
rect 832 4559 866 4593
rect 23597 4703 23631 4737
rect 23665 4703 23699 4737
rect 23733 4703 23767 4737
rect 23597 4634 23631 4668
rect 23665 4634 23699 4668
rect 23733 4634 23767 4668
rect 696 4487 730 4521
rect 764 4487 798 4521
rect 832 4487 866 4521
rect 696 4415 730 4449
rect 764 4415 798 4449
rect 832 4415 866 4449
rect 696 4343 730 4377
rect 764 4343 798 4377
rect 832 4343 866 4377
rect 696 4271 730 4305
rect 764 4271 798 4305
rect 832 4271 866 4305
rect 696 4199 730 4233
rect 764 4199 798 4233
rect 832 4199 866 4233
rect 696 4127 730 4161
rect 764 4127 798 4161
rect 832 4127 866 4161
rect 696 4055 730 4089
rect 764 4055 798 4089
rect 832 4055 866 4089
rect 696 3983 730 4017
rect 764 3983 798 4017
rect 832 3983 866 4017
rect 696 3912 730 3946
rect 764 3912 798 3946
rect 832 3912 866 3946
rect 696 3841 730 3875
rect 764 3841 798 3875
rect 832 3841 866 3875
rect 696 3770 730 3804
rect 764 3770 798 3804
rect 832 3770 866 3804
rect 696 3699 730 3733
rect 764 3699 798 3733
rect 832 3699 866 3733
rect 696 3628 730 3662
rect 764 3628 798 3662
rect 832 3628 866 3662
rect 696 3557 730 3591
rect 764 3557 798 3591
rect 832 3557 866 3591
rect 696 3486 730 3520
rect 764 3486 798 3520
rect 832 3486 866 3520
rect 696 3415 730 3449
rect 764 3415 798 3449
rect 832 3415 866 3449
rect 696 3344 730 3378
rect 764 3344 798 3378
rect 832 3344 866 3378
rect 696 3252 730 3286
rect 764 3252 798 3286
rect 832 3252 866 3286
rect 696 3182 730 3216
rect 764 3183 798 3217
rect 832 3183 866 3217
rect 696 3112 730 3146
rect 764 3114 798 3148
rect 832 3114 866 3148
rect 696 3042 730 3076
rect 764 3045 798 3079
rect 832 3045 866 3079
rect 696 2972 730 3006
rect 764 2976 798 3010
rect 832 2976 866 3010
rect 696 2903 730 2937
rect 696 2834 730 2868
rect 696 2765 730 2799
rect 696 2696 730 2730
rect 696 2627 730 2661
rect 696 2558 730 2592
rect 696 2489 730 2523
rect 696 2420 730 2454
rect 696 2351 730 2385
rect 696 2282 730 2316
rect 696 2213 730 2247
rect 696 2144 730 2178
rect 696 2075 730 2109
rect 696 2006 730 2040
rect 696 1937 730 1971
rect 696 1868 730 1902
rect 696 1799 730 1833
rect 696 1730 730 1764
rect 696 1661 730 1695
rect 696 1592 730 1626
rect 696 1523 730 1557
rect 696 1454 730 1488
rect 696 1385 730 1419
rect 696 1316 730 1350
rect 696 1247 730 1281
rect 764 1261 866 2941
rect 23597 4565 23631 4599
rect 23665 4565 23699 4599
rect 23733 4565 23767 4599
rect 23597 4496 23631 4530
rect 23665 4496 23699 4530
rect 23733 4496 23767 4530
rect 23597 4427 23631 4461
rect 23665 4427 23699 4461
rect 23733 4427 23767 4461
rect 23597 4358 23631 4392
rect 23665 4358 23699 4392
rect 23733 4358 23767 4392
rect 23597 4289 23631 4323
rect 23665 4289 23699 4323
rect 23733 4289 23767 4323
rect 23597 4220 23631 4254
rect 23665 4220 23699 4254
rect 23733 4220 23767 4254
rect 23597 4151 23631 4185
rect 23665 4151 23699 4185
rect 23733 4151 23767 4185
rect 23597 2110 23767 4116
rect 13751 2018 13785 2052
rect 13819 2018 13853 2052
rect 13887 2018 13921 2052
rect 13955 2018 13989 2052
rect 14023 2018 14057 2052
rect 14091 2018 14125 2052
rect 14159 2018 14193 2052
rect 14227 2018 14261 2052
rect 14295 2018 14329 2052
rect 14363 2018 14397 2052
rect 14489 2042 14523 2076
rect 14567 2042 14601 2076
rect 13751 1946 13785 1980
rect 13819 1946 13853 1980
rect 13887 1946 13921 1980
rect 13955 1946 13989 1980
rect 14023 1946 14057 1980
rect 14091 1946 14125 1980
rect 14159 1946 14193 1980
rect 14227 1946 14261 1980
rect 14295 1946 14329 1980
rect 14363 1946 14397 1980
rect 14545 1974 14579 2008
rect 14455 1934 14489 1968
rect 13751 1874 13785 1908
rect 13819 1874 13853 1908
rect 13887 1874 13921 1908
rect 13955 1874 13989 1908
rect 14023 1874 14057 1908
rect 14091 1874 14125 1908
rect 14159 1874 14193 1908
rect 14227 1874 14261 1908
rect 14295 1874 14329 1908
rect 14363 1874 14397 1908
rect 14523 1905 14557 1939
rect 14455 1863 14489 1897
rect 14591 1882 14625 1916
rect 14523 1836 14557 1870
rect 13751 1802 13785 1836
rect 13819 1802 13853 1836
rect 13887 1802 13921 1836
rect 13955 1802 13989 1836
rect 14023 1802 14057 1836
rect 14091 1802 14125 1836
rect 14159 1802 14193 1836
rect 14227 1802 14261 1836
rect 14295 1802 14329 1836
rect 14363 1802 14397 1836
rect 14455 1792 14489 1826
rect 14591 1812 14625 1846
rect 14523 1767 14557 1801
rect 13751 1730 13785 1764
rect 13819 1730 13853 1764
rect 13887 1730 13921 1764
rect 13955 1730 13989 1764
rect 14023 1730 14057 1764
rect 14091 1730 14125 1764
rect 14159 1730 14193 1764
rect 14227 1730 14261 1764
rect 14295 1730 14329 1764
rect 14363 1730 14397 1764
rect 14455 1721 14489 1755
rect 14591 1742 14625 1776
rect 14523 1698 14557 1732
rect 13751 1658 13785 1692
rect 13819 1658 13853 1692
rect 13887 1658 13921 1692
rect 13955 1658 13989 1692
rect 14023 1658 14057 1692
rect 14091 1658 14125 1692
rect 14159 1658 14193 1692
rect 14227 1658 14261 1692
rect 14295 1658 14329 1692
rect 14363 1658 14397 1692
rect 14455 1650 14489 1684
rect 14591 1672 14625 1706
rect 14523 1629 14557 1663
rect 13751 1586 13785 1620
rect 13819 1586 13853 1620
rect 13887 1586 13921 1620
rect 13955 1586 13989 1620
rect 14023 1586 14057 1620
rect 14091 1586 14125 1620
rect 14159 1586 14193 1620
rect 14227 1586 14261 1620
rect 14295 1586 14329 1620
rect 14363 1586 14397 1620
rect 14455 1579 14489 1613
rect 14591 1602 14625 1636
rect 14523 1560 14557 1594
rect 13751 1514 13785 1548
rect 13819 1514 13853 1548
rect 13887 1514 13921 1548
rect 13955 1514 13989 1548
rect 14023 1514 14057 1548
rect 14091 1514 14125 1548
rect 14159 1514 14193 1548
rect 14227 1514 14261 1548
rect 14295 1514 14329 1548
rect 14363 1514 14397 1548
rect 14455 1507 14489 1541
rect 14591 1532 14625 1566
rect 14523 1491 14557 1525
rect 13751 1441 13785 1475
rect 13819 1441 13853 1475
rect 13887 1441 13921 1475
rect 13955 1441 13989 1475
rect 14023 1441 14057 1475
rect 14091 1441 14125 1475
rect 14159 1441 14193 1475
rect 14227 1441 14261 1475
rect 14295 1441 14329 1475
rect 14363 1441 14397 1475
rect 14455 1435 14489 1469
rect 14591 1462 14625 1496
rect 14523 1422 14557 1456
rect 13751 1368 13785 1402
rect 13819 1368 13853 1402
rect 13887 1368 13921 1402
rect 13955 1368 13989 1402
rect 14023 1368 14057 1402
rect 14091 1368 14125 1402
rect 14159 1368 14193 1402
rect 14227 1368 14261 1402
rect 14295 1368 14329 1402
rect 14363 1368 14397 1402
rect 14455 1363 14489 1397
rect 14591 1392 14625 1426
rect 14523 1353 14557 1387
rect 13751 1261 14397 1329
rect 14455 1291 14489 1325
rect 14591 1322 14625 1356
rect 14523 1284 14557 1318
rect 696 1178 730 1212
rect 696 1109 730 1143
rect 764 1091 934 1261
rect 969 1227 1003 1261
rect 1038 1227 1072 1261
rect 1107 1227 1141 1261
rect 1176 1227 1210 1261
rect 1245 1227 1279 1261
rect 1314 1227 1348 1261
rect 1383 1227 1417 1261
rect 1452 1227 1486 1261
rect 1521 1227 1555 1261
rect 1590 1227 1624 1261
rect 1659 1227 1693 1261
rect 1728 1227 1762 1261
rect 1797 1227 1831 1261
rect 1866 1227 1900 1261
rect 1935 1227 1969 1261
rect 2004 1227 2038 1261
rect 2073 1227 2107 1261
rect 2142 1227 2176 1261
rect 2211 1227 2245 1261
rect 2280 1227 2314 1261
rect 2349 1227 2383 1261
rect 2418 1227 2452 1261
rect 2487 1227 2521 1261
rect 2556 1227 2590 1261
rect 2625 1227 2659 1261
rect 2694 1227 2728 1261
rect 2763 1227 2797 1261
rect 2832 1227 2866 1261
rect 2901 1227 2935 1261
rect 2970 1227 3004 1261
rect 3039 1227 3073 1261
rect 3108 1227 3142 1261
rect 3177 1227 3211 1261
rect 3246 1227 3280 1261
rect 3315 1227 3349 1261
rect 3384 1227 3418 1261
rect 3453 1227 3487 1261
rect 3522 1227 3556 1261
rect 3591 1227 3625 1261
rect 3660 1227 3694 1261
rect 3729 1227 3763 1261
rect 3798 1227 3832 1261
rect 3867 1227 3901 1261
rect 3936 1227 3970 1261
rect 4005 1227 4039 1261
rect 4074 1227 4108 1261
rect 4143 1227 4177 1261
rect 4212 1227 4246 1261
rect 4281 1227 4315 1261
rect 4350 1227 4384 1261
rect 4419 1227 4453 1261
rect 4488 1227 4522 1261
rect 4557 1227 4591 1261
rect 4626 1227 4660 1261
rect 4695 1227 4729 1261
rect 4764 1227 4798 1261
rect 4833 1227 4867 1261
rect 4902 1227 4936 1261
rect 4971 1227 5005 1261
rect 5040 1227 5074 1261
rect 5109 1227 5143 1261
rect 5178 1227 5212 1261
rect 5247 1227 5281 1261
rect 5316 1227 5350 1261
rect 5385 1227 5419 1261
rect 5454 1227 5488 1261
rect 969 1159 1003 1193
rect 1038 1159 1072 1193
rect 1107 1159 1141 1193
rect 1176 1159 1210 1193
rect 1245 1159 1279 1193
rect 1314 1159 1348 1193
rect 1383 1159 1417 1193
rect 1452 1159 1486 1193
rect 1521 1159 1555 1193
rect 1590 1159 1624 1193
rect 1659 1159 1693 1193
rect 1728 1159 1762 1193
rect 1797 1159 1831 1193
rect 1866 1159 1900 1193
rect 1935 1159 1969 1193
rect 2004 1159 2038 1193
rect 2073 1159 2107 1193
rect 2142 1159 2176 1193
rect 2211 1159 2245 1193
rect 2280 1159 2314 1193
rect 2349 1159 2383 1193
rect 2418 1159 2452 1193
rect 2487 1159 2521 1193
rect 2556 1159 2590 1193
rect 2625 1159 2659 1193
rect 2694 1159 2728 1193
rect 2763 1159 2797 1193
rect 2832 1159 2866 1193
rect 2901 1159 2935 1193
rect 2970 1159 3004 1193
rect 3039 1159 3073 1193
rect 3108 1159 3142 1193
rect 3177 1159 3211 1193
rect 3246 1159 3280 1193
rect 3315 1159 3349 1193
rect 3384 1159 3418 1193
rect 3453 1159 3487 1193
rect 3522 1159 3556 1193
rect 3591 1159 3625 1193
rect 3660 1159 3694 1193
rect 3729 1159 3763 1193
rect 3798 1159 3832 1193
rect 3867 1159 3901 1193
rect 3936 1159 3970 1193
rect 4005 1159 4039 1193
rect 4074 1159 4108 1193
rect 4143 1159 4177 1193
rect 4212 1159 4246 1193
rect 4281 1159 4315 1193
rect 4350 1159 4384 1193
rect 4419 1159 4453 1193
rect 4488 1159 4522 1193
rect 4557 1159 4591 1193
rect 4626 1159 4660 1193
rect 4695 1159 4729 1193
rect 4764 1159 4798 1193
rect 4833 1159 4867 1193
rect 4902 1159 4936 1193
rect 4971 1159 5005 1193
rect 5040 1159 5074 1193
rect 5109 1159 5143 1193
rect 5178 1159 5212 1193
rect 5247 1159 5281 1193
rect 5316 1159 5350 1193
rect 5385 1159 5419 1193
rect 5454 1159 5488 1193
rect 969 1091 1003 1125
rect 1038 1091 1072 1125
rect 1107 1091 1141 1125
rect 1176 1091 1210 1125
rect 1245 1091 1279 1125
rect 1314 1091 1348 1125
rect 1383 1091 1417 1125
rect 1452 1091 1486 1125
rect 1521 1091 1555 1125
rect 1590 1091 1624 1125
rect 1659 1091 1693 1125
rect 1728 1091 1762 1125
rect 1797 1091 1831 1125
rect 1866 1091 1900 1125
rect 1935 1091 1969 1125
rect 2004 1091 2038 1125
rect 2073 1091 2107 1125
rect 2142 1091 2176 1125
rect 2211 1091 2245 1125
rect 2280 1091 2314 1125
rect 2349 1091 2383 1125
rect 2418 1091 2452 1125
rect 2487 1091 2521 1125
rect 2556 1091 2590 1125
rect 2625 1091 2659 1125
rect 2694 1091 2728 1125
rect 2763 1091 2797 1125
rect 2832 1091 2866 1125
rect 2901 1091 2935 1125
rect 2970 1091 3004 1125
rect 3039 1091 3073 1125
rect 3108 1091 3142 1125
rect 3177 1091 3211 1125
rect 3246 1091 3280 1125
rect 3315 1091 3349 1125
rect 3384 1091 3418 1125
rect 3453 1091 3487 1125
rect 3522 1091 3556 1125
rect 3591 1091 3625 1125
rect 3660 1091 3694 1125
rect 3729 1091 3763 1125
rect 3798 1091 3832 1125
rect 3867 1091 3901 1125
rect 3936 1091 3970 1125
rect 4005 1091 4039 1125
rect 4074 1091 4108 1125
rect 4143 1091 4177 1125
rect 4212 1091 4246 1125
rect 4281 1091 4315 1125
rect 4350 1091 4384 1125
rect 4419 1091 4453 1125
rect 4488 1091 4522 1125
rect 4557 1091 4591 1125
rect 4626 1091 4660 1125
rect 4695 1091 4729 1125
rect 4764 1091 4798 1125
rect 4833 1091 4867 1125
rect 4902 1091 4936 1125
rect 4971 1091 5005 1125
rect 5040 1091 5074 1125
rect 5109 1091 5143 1125
rect 5178 1091 5212 1125
rect 5247 1091 5281 1125
rect 5316 1091 5350 1125
rect 5385 1091 5419 1125
rect 5454 1091 5488 1125
rect 5523 1091 14397 1261
rect 14455 1219 14489 1253
rect 14591 1252 14625 1286
rect 14523 1215 14557 1249
rect 14591 1182 14625 1216
rect 14455 1147 14489 1181
rect 14523 1145 14557 1179
rect 14591 1112 14625 1146
rect 14701 1143 19563 2061
rect 19598 2027 19632 2061
rect 19667 2027 19701 2061
rect 19736 2027 19770 2061
rect 19805 2027 19839 2061
rect 19874 2027 19908 2061
rect 19943 2027 19977 2061
rect 20012 2027 20046 2061
rect 20081 2027 20115 2061
rect 20150 2027 20184 2061
rect 20219 2027 20253 2061
rect 20288 2027 20322 2061
rect 20357 2027 20391 2061
rect 20426 2027 20460 2061
rect 20495 2027 20529 2061
rect 20564 2027 20598 2061
rect 20633 2027 20667 2061
rect 20702 2027 20736 2061
rect 20771 2027 20805 2061
rect 20840 2027 20874 2061
rect 20909 2027 20943 2061
rect 20978 2027 21012 2061
rect 21047 2027 21081 2061
rect 21116 2027 21150 2061
rect 21185 2027 21219 2061
rect 21254 2027 21288 2061
rect 21323 2027 21357 2061
rect 21392 2027 21426 2061
rect 21461 2027 21495 2061
rect 21530 2027 21564 2061
rect 21599 2027 21633 2061
rect 21668 2027 21702 2061
rect 21737 2027 21771 2061
rect 21806 2027 21840 2061
rect 21875 2027 21909 2061
rect 21944 2027 21978 2061
rect 22013 2027 22047 2061
rect 22082 2027 22116 2061
rect 22151 2027 22185 2061
rect 22220 2027 22254 2061
rect 22289 2027 22323 2061
rect 22358 2027 22392 2061
rect 22427 2027 22461 2061
rect 22496 2027 22530 2061
rect 22565 2027 22599 2061
rect 22634 2027 22668 2061
rect 22703 2027 22737 2061
rect 22772 2027 22806 2061
rect 22841 2027 22875 2061
rect 22910 2027 22944 2061
rect 22979 2027 23013 2061
rect 23048 2027 23082 2061
rect 23117 2027 23151 2061
rect 23186 2027 23220 2061
rect 23255 2027 23289 2061
rect 23324 2027 23358 2061
rect 23393 2027 23427 2061
rect 23462 2027 23496 2061
rect 23531 2027 23565 2061
rect 23600 2027 23634 2061
rect 23669 2027 23703 2061
rect 23738 2027 23772 2061
rect 19598 1959 19632 1993
rect 19667 1959 19701 1993
rect 19736 1959 19770 1993
rect 19805 1959 19839 1993
rect 19874 1959 19908 1993
rect 19943 1959 19977 1993
rect 20012 1959 20046 1993
rect 20081 1959 20115 1993
rect 20150 1959 20184 1993
rect 20219 1959 20253 1993
rect 20288 1959 20322 1993
rect 20357 1959 20391 1993
rect 20426 1959 20460 1993
rect 20495 1959 20529 1993
rect 20564 1959 20598 1993
rect 20633 1959 20667 1993
rect 20702 1959 20736 1993
rect 20771 1959 20805 1993
rect 20840 1959 20874 1993
rect 20909 1959 20943 1993
rect 20978 1959 21012 1993
rect 21047 1959 21081 1993
rect 21116 1959 21150 1993
rect 21185 1959 21219 1993
rect 21254 1959 21288 1993
rect 21323 1959 21357 1993
rect 21392 1959 21426 1993
rect 21461 1959 21495 1993
rect 21530 1959 21564 1993
rect 21599 1959 21633 1993
rect 21668 1959 21702 1993
rect 21737 1959 21771 1993
rect 21806 1959 21840 1993
rect 21875 1959 21909 1993
rect 21944 1959 21978 1993
rect 22013 1959 22047 1993
rect 22082 1959 22116 1993
rect 22151 1959 22185 1993
rect 22220 1959 22254 1993
rect 22289 1959 22323 1993
rect 22358 1959 22392 1993
rect 22427 1959 22461 1993
rect 22496 1959 22530 1993
rect 22565 1959 22599 1993
rect 22634 1959 22668 1993
rect 22703 1959 22737 1993
rect 22772 1959 22806 1993
rect 22841 1959 22875 1993
rect 22910 1959 22944 1993
rect 22979 1959 23013 1993
rect 23048 1959 23082 1993
rect 23117 1959 23151 1993
rect 23186 1959 23220 1993
rect 23255 1959 23289 1993
rect 23324 1959 23358 1993
rect 23393 1959 23427 1993
rect 23462 1959 23496 1993
rect 23531 1959 23565 1993
rect 23600 1959 23634 1993
rect 23669 1959 23703 1993
rect 23738 1959 23772 1993
rect 19598 1891 19632 1925
rect 19667 1891 19701 1925
rect 19736 1891 19770 1925
rect 19805 1891 19839 1925
rect 19874 1891 19908 1925
rect 19943 1891 19977 1925
rect 20012 1891 20046 1925
rect 20081 1891 20115 1925
rect 20150 1891 20184 1925
rect 20219 1891 20253 1925
rect 20288 1891 20322 1925
rect 20357 1891 20391 1925
rect 20426 1891 20460 1925
rect 20495 1891 20529 1925
rect 20564 1891 20598 1925
rect 20633 1891 20667 1925
rect 20702 1891 20736 1925
rect 20771 1891 20805 1925
rect 20840 1891 20874 1925
rect 20909 1891 20943 1925
rect 20978 1891 21012 1925
rect 21047 1891 21081 1925
rect 21116 1891 21150 1925
rect 21185 1891 21219 1925
rect 21254 1891 21288 1925
rect 21323 1891 21357 1925
rect 21392 1891 21426 1925
rect 21461 1891 21495 1925
rect 21530 1891 21564 1925
rect 21599 1891 21633 1925
rect 21668 1891 21702 1925
rect 21737 1891 21771 1925
rect 21806 1891 21840 1925
rect 21875 1891 21909 1925
rect 21944 1891 21978 1925
rect 22013 1891 22047 1925
rect 22082 1891 22116 1925
rect 22151 1891 22185 1925
rect 22220 1891 22254 1925
rect 22289 1891 22323 1925
rect 22358 1891 22392 1925
rect 22427 1891 22461 1925
rect 22496 1891 22530 1925
rect 22565 1891 22599 1925
rect 22634 1891 22668 1925
rect 22703 1891 22737 1925
rect 22772 1891 22806 1925
rect 22841 1891 22875 1925
rect 22910 1891 22944 1925
rect 22979 1891 23013 1925
rect 23048 1891 23082 1925
rect 23117 1891 23151 1925
rect 23186 1891 23220 1925
rect 23255 1891 23289 1925
rect 23324 1891 23358 1925
rect 23393 1891 23427 1925
rect 23462 1891 23496 1925
rect 23531 1891 23565 1925
rect 23600 1891 23634 1925
rect 23669 1891 23703 1925
rect 23738 1891 23772 1925
rect 19598 1823 19632 1857
rect 19667 1823 19701 1857
rect 19736 1823 19770 1857
rect 19805 1823 19839 1857
rect 19874 1823 19908 1857
rect 19943 1823 19977 1857
rect 20012 1823 20046 1857
rect 20081 1823 20115 1857
rect 20150 1823 20184 1857
rect 20219 1823 20253 1857
rect 20288 1823 20322 1857
rect 20357 1823 20391 1857
rect 20426 1823 20460 1857
rect 20495 1823 20529 1857
rect 20564 1823 20598 1857
rect 20633 1823 20667 1857
rect 20702 1823 20736 1857
rect 20771 1823 20805 1857
rect 20840 1823 20874 1857
rect 20909 1823 20943 1857
rect 20978 1823 21012 1857
rect 21047 1823 21081 1857
rect 21116 1823 21150 1857
rect 21185 1823 21219 1857
rect 21254 1823 21288 1857
rect 21323 1823 21357 1857
rect 21392 1823 21426 1857
rect 21461 1823 21495 1857
rect 21530 1823 21564 1857
rect 21599 1823 21633 1857
rect 21668 1823 21702 1857
rect 21737 1823 21771 1857
rect 21806 1823 21840 1857
rect 21875 1823 21909 1857
rect 21944 1823 21978 1857
rect 22013 1823 22047 1857
rect 22082 1823 22116 1857
rect 22151 1823 22185 1857
rect 22220 1823 22254 1857
rect 22289 1823 22323 1857
rect 22358 1823 22392 1857
rect 22427 1823 22461 1857
rect 22496 1823 22530 1857
rect 22565 1823 22599 1857
rect 22634 1823 22668 1857
rect 22703 1823 22737 1857
rect 22772 1823 22806 1857
rect 22841 1823 22875 1857
rect 22910 1823 22944 1857
rect 22979 1823 23013 1857
rect 23048 1823 23082 1857
rect 23117 1823 23151 1857
rect 23186 1823 23220 1857
rect 23255 1823 23289 1857
rect 23324 1823 23358 1857
rect 23393 1823 23427 1857
rect 23462 1823 23496 1857
rect 23531 1823 23565 1857
rect 23600 1823 23634 1857
rect 23669 1823 23703 1857
rect 23738 1823 23772 1857
rect 19598 1755 19632 1789
rect 19667 1755 19701 1789
rect 19736 1755 19770 1789
rect 19805 1755 19839 1789
rect 19874 1755 19908 1789
rect 19943 1755 19977 1789
rect 20012 1755 20046 1789
rect 20081 1755 20115 1789
rect 20150 1755 20184 1789
rect 20219 1755 20253 1789
rect 20288 1755 20322 1789
rect 20357 1755 20391 1789
rect 20426 1755 20460 1789
rect 20495 1755 20529 1789
rect 20564 1755 20598 1789
rect 20633 1755 20667 1789
rect 20702 1755 20736 1789
rect 20771 1755 20805 1789
rect 20840 1755 20874 1789
rect 20909 1755 20943 1789
rect 20978 1755 21012 1789
rect 21047 1755 21081 1789
rect 21116 1755 21150 1789
rect 21185 1755 21219 1789
rect 21254 1755 21288 1789
rect 21323 1755 21357 1789
rect 21392 1755 21426 1789
rect 21461 1755 21495 1789
rect 21530 1755 21564 1789
rect 21599 1755 21633 1789
rect 21668 1755 21702 1789
rect 21737 1755 21771 1789
rect 21806 1755 21840 1789
rect 21875 1755 21909 1789
rect 21944 1755 21978 1789
rect 22013 1755 22047 1789
rect 22082 1755 22116 1789
rect 22151 1755 22185 1789
rect 22220 1755 22254 1789
rect 22289 1755 22323 1789
rect 22358 1755 22392 1789
rect 22427 1755 22461 1789
rect 22496 1755 22530 1789
rect 22565 1755 22599 1789
rect 22634 1755 22668 1789
rect 22703 1755 22737 1789
rect 22772 1755 22806 1789
rect 22841 1755 22875 1789
rect 22910 1755 22944 1789
rect 22979 1755 23013 1789
rect 23048 1755 23082 1789
rect 23117 1755 23151 1789
rect 23186 1755 23220 1789
rect 23255 1755 23289 1789
rect 23324 1755 23358 1789
rect 23393 1755 23427 1789
rect 23462 1755 23496 1789
rect 23531 1755 23565 1789
rect 23600 1755 23634 1789
rect 23669 1755 23703 1789
rect 23738 1755 23772 1789
rect 19598 1687 19632 1721
rect 19667 1687 19701 1721
rect 19736 1687 19770 1721
rect 19805 1687 19839 1721
rect 19874 1687 19908 1721
rect 19943 1687 19977 1721
rect 20012 1687 20046 1721
rect 20081 1687 20115 1721
rect 20150 1687 20184 1721
rect 20219 1687 20253 1721
rect 20288 1687 20322 1721
rect 20357 1687 20391 1721
rect 20426 1687 20460 1721
rect 20495 1687 20529 1721
rect 20564 1687 20598 1721
rect 20633 1687 20667 1721
rect 20702 1687 20736 1721
rect 20771 1687 20805 1721
rect 20840 1687 20874 1721
rect 20909 1687 20943 1721
rect 20978 1687 21012 1721
rect 21047 1687 21081 1721
rect 21116 1687 21150 1721
rect 21185 1687 21219 1721
rect 21254 1687 21288 1721
rect 21323 1687 21357 1721
rect 21392 1687 21426 1721
rect 21461 1687 21495 1721
rect 21530 1687 21564 1721
rect 21599 1687 21633 1721
rect 21668 1687 21702 1721
rect 21737 1687 21771 1721
rect 21806 1687 21840 1721
rect 21875 1687 21909 1721
rect 21944 1687 21978 1721
rect 22013 1687 22047 1721
rect 22082 1687 22116 1721
rect 22151 1687 22185 1721
rect 22220 1687 22254 1721
rect 22289 1687 22323 1721
rect 22358 1687 22392 1721
rect 22427 1687 22461 1721
rect 22496 1687 22530 1721
rect 22565 1687 22599 1721
rect 22634 1687 22668 1721
rect 22703 1687 22737 1721
rect 22772 1687 22806 1721
rect 22841 1687 22875 1721
rect 22910 1687 22944 1721
rect 22979 1687 23013 1721
rect 23048 1687 23082 1721
rect 23117 1687 23151 1721
rect 23186 1687 23220 1721
rect 23255 1687 23289 1721
rect 23324 1687 23358 1721
rect 23393 1687 23427 1721
rect 23462 1687 23496 1721
rect 23531 1687 23565 1721
rect 23600 1687 23634 1721
rect 23669 1687 23703 1721
rect 23738 1687 23772 1721
rect 19598 1619 19632 1653
rect 19667 1619 19701 1653
rect 19736 1619 19770 1653
rect 19805 1619 19839 1653
rect 19874 1619 19908 1653
rect 19943 1619 19977 1653
rect 20012 1619 20046 1653
rect 20081 1619 20115 1653
rect 20150 1619 20184 1653
rect 20219 1619 20253 1653
rect 20288 1619 20322 1653
rect 20357 1619 20391 1653
rect 20426 1619 20460 1653
rect 20495 1619 20529 1653
rect 20564 1619 20598 1653
rect 20633 1619 20667 1653
rect 20702 1619 20736 1653
rect 20771 1619 20805 1653
rect 20840 1619 20874 1653
rect 20909 1619 20943 1653
rect 20978 1619 21012 1653
rect 21047 1619 21081 1653
rect 21116 1619 21150 1653
rect 21185 1619 21219 1653
rect 21254 1619 21288 1653
rect 21323 1619 21357 1653
rect 21392 1619 21426 1653
rect 21461 1619 21495 1653
rect 21530 1619 21564 1653
rect 21599 1619 21633 1653
rect 21668 1619 21702 1653
rect 21737 1619 21771 1653
rect 21806 1619 21840 1653
rect 21875 1619 21909 1653
rect 21944 1619 21978 1653
rect 22013 1619 22047 1653
rect 22082 1619 22116 1653
rect 22151 1619 22185 1653
rect 22220 1619 22254 1653
rect 22289 1619 22323 1653
rect 22358 1619 22392 1653
rect 22427 1619 22461 1653
rect 22496 1619 22530 1653
rect 22565 1619 22599 1653
rect 22634 1619 22668 1653
rect 22703 1619 22737 1653
rect 22772 1619 22806 1653
rect 22841 1619 22875 1653
rect 22910 1619 22944 1653
rect 22979 1619 23013 1653
rect 23048 1619 23082 1653
rect 23117 1619 23151 1653
rect 23186 1619 23220 1653
rect 23255 1619 23289 1653
rect 23324 1619 23358 1653
rect 23393 1619 23427 1653
rect 23462 1619 23496 1653
rect 23531 1619 23565 1653
rect 23600 1619 23634 1653
rect 23669 1619 23703 1653
rect 23738 1619 23772 1653
rect 19598 1551 19632 1585
rect 19667 1551 19701 1585
rect 19736 1551 19770 1585
rect 19805 1551 19839 1585
rect 19874 1551 19908 1585
rect 19943 1551 19977 1585
rect 20012 1551 20046 1585
rect 20081 1551 20115 1585
rect 20150 1551 20184 1585
rect 20219 1551 20253 1585
rect 20288 1551 20322 1585
rect 20357 1551 20391 1585
rect 20426 1551 20460 1585
rect 20495 1551 20529 1585
rect 20564 1551 20598 1585
rect 20633 1551 20667 1585
rect 20702 1551 20736 1585
rect 20771 1551 20805 1585
rect 20840 1551 20874 1585
rect 20909 1551 20943 1585
rect 20978 1551 21012 1585
rect 21047 1551 21081 1585
rect 21116 1551 21150 1585
rect 21185 1551 21219 1585
rect 21254 1551 21288 1585
rect 21323 1551 21357 1585
rect 21392 1551 21426 1585
rect 21461 1551 21495 1585
rect 21530 1551 21564 1585
rect 21599 1551 21633 1585
rect 21668 1551 21702 1585
rect 21737 1551 21771 1585
rect 21806 1551 21840 1585
rect 21875 1551 21909 1585
rect 21944 1551 21978 1585
rect 22013 1551 22047 1585
rect 22082 1551 22116 1585
rect 22151 1551 22185 1585
rect 22220 1551 22254 1585
rect 22289 1551 22323 1585
rect 22358 1551 22392 1585
rect 22427 1551 22461 1585
rect 22496 1551 22530 1585
rect 22565 1551 22599 1585
rect 22634 1551 22668 1585
rect 22703 1551 22737 1585
rect 22772 1551 22806 1585
rect 22841 1551 22875 1585
rect 22910 1551 22944 1585
rect 22979 1551 23013 1585
rect 23048 1551 23082 1585
rect 23117 1551 23151 1585
rect 23186 1551 23220 1585
rect 23255 1551 23289 1585
rect 23324 1551 23358 1585
rect 23393 1551 23427 1585
rect 23462 1551 23496 1585
rect 23531 1551 23565 1585
rect 23600 1551 23634 1585
rect 23669 1551 23703 1585
rect 23738 1551 23772 1585
rect 19598 1483 19632 1517
rect 19667 1483 19701 1517
rect 19736 1483 19770 1517
rect 19805 1483 19839 1517
rect 19874 1483 19908 1517
rect 19943 1483 19977 1517
rect 20012 1483 20046 1517
rect 20081 1483 20115 1517
rect 20150 1483 20184 1517
rect 20219 1483 20253 1517
rect 20288 1483 20322 1517
rect 20357 1483 20391 1517
rect 20426 1483 20460 1517
rect 20495 1483 20529 1517
rect 20564 1483 20598 1517
rect 20633 1483 20667 1517
rect 20702 1483 20736 1517
rect 20771 1483 20805 1517
rect 20840 1483 20874 1517
rect 20909 1483 20943 1517
rect 20978 1483 21012 1517
rect 21047 1483 21081 1517
rect 21116 1483 21150 1517
rect 21185 1483 21219 1517
rect 21254 1483 21288 1517
rect 21323 1483 21357 1517
rect 21392 1483 21426 1517
rect 21461 1483 21495 1517
rect 21530 1483 21564 1517
rect 21599 1483 21633 1517
rect 21668 1483 21702 1517
rect 21737 1483 21771 1517
rect 21806 1483 21840 1517
rect 21875 1483 21909 1517
rect 21944 1483 21978 1517
rect 22013 1483 22047 1517
rect 22082 1483 22116 1517
rect 22151 1483 22185 1517
rect 22220 1483 22254 1517
rect 22289 1483 22323 1517
rect 22358 1483 22392 1517
rect 22427 1483 22461 1517
rect 22496 1483 22530 1517
rect 22565 1483 22599 1517
rect 22634 1483 22668 1517
rect 22703 1483 22737 1517
rect 22772 1483 22806 1517
rect 22841 1483 22875 1517
rect 22910 1483 22944 1517
rect 22979 1483 23013 1517
rect 23048 1483 23082 1517
rect 23117 1483 23151 1517
rect 23186 1483 23220 1517
rect 23255 1483 23289 1517
rect 23324 1483 23358 1517
rect 23393 1483 23427 1517
rect 23462 1483 23496 1517
rect 23531 1483 23565 1517
rect 23600 1483 23634 1517
rect 23669 1483 23703 1517
rect 23738 1483 23772 1517
rect 19598 1415 19632 1449
rect 19667 1415 19701 1449
rect 19736 1415 19770 1449
rect 19805 1415 19839 1449
rect 19874 1415 19908 1449
rect 19943 1415 19977 1449
rect 20012 1415 20046 1449
rect 20081 1415 20115 1449
rect 20150 1415 20184 1449
rect 20219 1415 20253 1449
rect 20288 1415 20322 1449
rect 20357 1415 20391 1449
rect 20426 1415 20460 1449
rect 20495 1415 20529 1449
rect 20564 1415 20598 1449
rect 20633 1415 20667 1449
rect 20702 1415 20736 1449
rect 20771 1415 20805 1449
rect 20840 1415 20874 1449
rect 20909 1415 20943 1449
rect 20978 1415 21012 1449
rect 21047 1415 21081 1449
rect 21116 1415 21150 1449
rect 21185 1415 21219 1449
rect 21254 1415 21288 1449
rect 21323 1415 21357 1449
rect 21392 1415 21426 1449
rect 21461 1415 21495 1449
rect 21530 1415 21564 1449
rect 21599 1415 21633 1449
rect 21668 1415 21702 1449
rect 21737 1415 21771 1449
rect 21806 1415 21840 1449
rect 21875 1415 21909 1449
rect 21944 1415 21978 1449
rect 22013 1415 22047 1449
rect 22082 1415 22116 1449
rect 22151 1415 22185 1449
rect 22220 1415 22254 1449
rect 22289 1415 22323 1449
rect 22358 1415 22392 1449
rect 22427 1415 22461 1449
rect 22496 1415 22530 1449
rect 22565 1415 22599 1449
rect 22634 1415 22668 1449
rect 22703 1415 22737 1449
rect 22772 1415 22806 1449
rect 22841 1415 22875 1449
rect 22910 1415 22944 1449
rect 22979 1415 23013 1449
rect 23048 1415 23082 1449
rect 23117 1415 23151 1449
rect 23186 1415 23220 1449
rect 23255 1415 23289 1449
rect 23324 1415 23358 1449
rect 23393 1415 23427 1449
rect 23462 1415 23496 1449
rect 23531 1415 23565 1449
rect 23600 1415 23634 1449
rect 23669 1415 23703 1449
rect 23738 1415 23772 1449
rect 19598 1347 19632 1381
rect 19667 1347 19701 1381
rect 19736 1347 19770 1381
rect 19805 1347 19839 1381
rect 19874 1347 19908 1381
rect 19943 1347 19977 1381
rect 20012 1347 20046 1381
rect 20081 1347 20115 1381
rect 20150 1347 20184 1381
rect 20219 1347 20253 1381
rect 20288 1347 20322 1381
rect 20357 1347 20391 1381
rect 20426 1347 20460 1381
rect 20495 1347 20529 1381
rect 20564 1347 20598 1381
rect 20633 1347 20667 1381
rect 20702 1347 20736 1381
rect 20771 1347 20805 1381
rect 20840 1347 20874 1381
rect 20909 1347 20943 1381
rect 20978 1347 21012 1381
rect 21047 1347 21081 1381
rect 21116 1347 21150 1381
rect 21185 1347 21219 1381
rect 21254 1347 21288 1381
rect 21323 1347 21357 1381
rect 21392 1347 21426 1381
rect 21461 1347 21495 1381
rect 21530 1347 21564 1381
rect 21599 1347 21633 1381
rect 21668 1347 21702 1381
rect 21737 1347 21771 1381
rect 21806 1347 21840 1381
rect 21875 1347 21909 1381
rect 21944 1347 21978 1381
rect 22013 1347 22047 1381
rect 22082 1347 22116 1381
rect 22151 1347 22185 1381
rect 22220 1347 22254 1381
rect 22289 1347 22323 1381
rect 22358 1347 22392 1381
rect 22427 1347 22461 1381
rect 22496 1347 22530 1381
rect 22565 1347 22599 1381
rect 22634 1347 22668 1381
rect 22703 1347 22737 1381
rect 22772 1347 22806 1381
rect 22841 1347 22875 1381
rect 22910 1347 22944 1381
rect 22979 1347 23013 1381
rect 23048 1347 23082 1381
rect 23117 1347 23151 1381
rect 23186 1347 23220 1381
rect 23255 1347 23289 1381
rect 23324 1347 23358 1381
rect 23393 1347 23427 1381
rect 23462 1347 23496 1381
rect 23531 1347 23565 1381
rect 23600 1347 23634 1381
rect 23669 1347 23703 1381
rect 23738 1347 23772 1381
rect 19598 1279 19632 1313
rect 19667 1279 19701 1313
rect 19736 1279 19770 1313
rect 19805 1279 19839 1313
rect 19874 1279 19908 1313
rect 19943 1279 19977 1313
rect 20012 1279 20046 1313
rect 20081 1279 20115 1313
rect 20150 1279 20184 1313
rect 20219 1279 20253 1313
rect 20288 1279 20322 1313
rect 20357 1279 20391 1313
rect 20426 1279 20460 1313
rect 20495 1279 20529 1313
rect 20564 1279 20598 1313
rect 20633 1279 20667 1313
rect 20702 1279 20736 1313
rect 20771 1279 20805 1313
rect 20840 1279 20874 1313
rect 20909 1279 20943 1313
rect 20978 1279 21012 1313
rect 21047 1279 21081 1313
rect 21116 1279 21150 1313
rect 21185 1279 21219 1313
rect 21254 1279 21288 1313
rect 21323 1279 21357 1313
rect 21392 1279 21426 1313
rect 21461 1279 21495 1313
rect 21530 1279 21564 1313
rect 21599 1279 21633 1313
rect 21668 1279 21702 1313
rect 21737 1279 21771 1313
rect 21806 1279 21840 1313
rect 21875 1279 21909 1313
rect 21944 1279 21978 1313
rect 22013 1279 22047 1313
rect 22082 1279 22116 1313
rect 22151 1279 22185 1313
rect 22220 1279 22254 1313
rect 22289 1279 22323 1313
rect 22358 1279 22392 1313
rect 22427 1279 22461 1313
rect 22496 1279 22530 1313
rect 22565 1279 22599 1313
rect 22634 1279 22668 1313
rect 22703 1279 22737 1313
rect 22772 1279 22806 1313
rect 22841 1279 22875 1313
rect 22910 1279 22944 1313
rect 22979 1279 23013 1313
rect 23048 1279 23082 1313
rect 23117 1279 23151 1313
rect 23186 1279 23220 1313
rect 23255 1279 23289 1313
rect 23324 1279 23358 1313
rect 23393 1279 23427 1313
rect 23462 1279 23496 1313
rect 23531 1279 23565 1313
rect 23600 1279 23634 1313
rect 23669 1279 23703 1313
rect 23738 1279 23772 1313
rect 19598 1211 19632 1245
rect 19667 1211 19701 1245
rect 19736 1211 19770 1245
rect 19805 1211 19839 1245
rect 19874 1211 19908 1245
rect 19943 1211 19977 1245
rect 20012 1211 20046 1245
rect 20081 1211 20115 1245
rect 20150 1211 20184 1245
rect 20219 1211 20253 1245
rect 20288 1211 20322 1245
rect 20357 1211 20391 1245
rect 20426 1211 20460 1245
rect 20495 1211 20529 1245
rect 20564 1211 20598 1245
rect 20633 1211 20667 1245
rect 20702 1211 20736 1245
rect 20771 1211 20805 1245
rect 20840 1211 20874 1245
rect 20909 1211 20943 1245
rect 20978 1211 21012 1245
rect 21047 1211 21081 1245
rect 21116 1211 21150 1245
rect 21185 1211 21219 1245
rect 21254 1211 21288 1245
rect 21323 1211 21357 1245
rect 21392 1211 21426 1245
rect 21461 1211 21495 1245
rect 21530 1211 21564 1245
rect 21599 1211 21633 1245
rect 21668 1211 21702 1245
rect 21737 1211 21771 1245
rect 21806 1211 21840 1245
rect 21875 1211 21909 1245
rect 21944 1211 21978 1245
rect 22013 1211 22047 1245
rect 22082 1211 22116 1245
rect 22151 1211 22185 1245
rect 22220 1211 22254 1245
rect 22289 1211 22323 1245
rect 22358 1211 22392 1245
rect 22427 1211 22461 1245
rect 22496 1211 22530 1245
rect 22565 1211 22599 1245
rect 22634 1211 22668 1245
rect 22703 1211 22737 1245
rect 22772 1211 22806 1245
rect 22841 1211 22875 1245
rect 22910 1211 22944 1245
rect 22979 1211 23013 1245
rect 23048 1211 23082 1245
rect 23117 1211 23151 1245
rect 23186 1211 23220 1245
rect 23255 1211 23289 1245
rect 23324 1211 23358 1245
rect 23393 1211 23427 1245
rect 23462 1211 23496 1245
rect 23531 1211 23565 1245
rect 23600 1211 23634 1245
rect 23669 1211 23703 1245
rect 23738 1211 23772 1245
rect 19598 1143 19632 1177
rect 19667 1143 19701 1177
rect 19736 1143 19770 1177
rect 19805 1143 19839 1177
rect 19874 1143 19908 1177
rect 19943 1143 19977 1177
rect 20012 1143 20046 1177
rect 20081 1143 20115 1177
rect 20150 1143 20184 1177
rect 20219 1143 20253 1177
rect 20288 1143 20322 1177
rect 20357 1143 20391 1177
rect 20426 1143 20460 1177
rect 20495 1143 20529 1177
rect 20564 1143 20598 1177
rect 20633 1143 20667 1177
rect 20702 1143 20736 1177
rect 20771 1143 20805 1177
rect 20840 1143 20874 1177
rect 20909 1143 20943 1177
rect 20978 1143 21012 1177
rect 21047 1143 21081 1177
rect 21116 1143 21150 1177
rect 21185 1143 21219 1177
rect 21254 1143 21288 1177
rect 21323 1143 21357 1177
rect 21392 1143 21426 1177
rect 21461 1143 21495 1177
rect 21530 1143 21564 1177
rect 21599 1143 21633 1177
rect 21668 1143 21702 1177
rect 21737 1143 21771 1177
rect 21806 1143 21840 1177
rect 21875 1143 21909 1177
rect 21944 1143 21978 1177
rect 22013 1143 22047 1177
rect 22082 1143 22116 1177
rect 22151 1143 22185 1177
rect 22220 1143 22254 1177
rect 22289 1143 22323 1177
rect 22358 1143 22392 1177
rect 22427 1143 22461 1177
rect 22496 1143 22530 1177
rect 22565 1143 22599 1177
rect 22634 1143 22668 1177
rect 22703 1143 22737 1177
rect 22772 1143 22806 1177
rect 22841 1143 22875 1177
rect 22910 1143 22944 1177
rect 22979 1143 23013 1177
rect 23048 1143 23082 1177
rect 23117 1143 23151 1177
rect 23186 1143 23220 1177
rect 23255 1143 23289 1177
rect 23324 1143 23358 1177
rect 23393 1143 23427 1177
rect 23462 1143 23496 1177
rect 23531 1143 23565 1177
rect 23600 1143 23634 1177
rect 23669 1143 23703 1177
rect 23738 1143 23772 1177
rect 696 1040 730 1074
rect 696 971 730 1005
rect 764 1003 866 1091
rect 14455 1075 14489 1109
rect 14523 1075 14557 1109
rect 14591 1042 14625 1076
rect 901 1003 935 1037
rect 970 1003 1004 1037
rect 1039 1003 1073 1037
rect 1108 1003 1142 1037
rect 1177 1003 1211 1037
rect 1246 1003 1280 1037
rect 1315 1003 1349 1037
rect 1384 1003 1418 1037
rect 1453 1003 1487 1037
rect 1522 1003 1556 1037
rect 1591 1003 1625 1037
rect 1660 1003 1694 1037
rect 1729 1003 1763 1037
rect 1798 1003 1832 1037
rect 1867 1003 1901 1037
rect 1936 1003 1970 1037
rect 2005 1003 2039 1037
rect 2074 1003 2108 1037
rect 2143 1003 2177 1037
rect 2212 1003 2246 1037
rect 2281 1003 2315 1037
rect 2350 1003 2384 1037
rect 2419 969 14489 1037
rect 14523 1005 14557 1039
rect 14591 972 14625 1006
rect 764 935 798 969
rect 833 935 867 969
rect 902 935 936 969
rect 971 935 1005 969
rect 1040 935 1074 969
rect 1109 935 1143 969
rect 1178 935 1212 969
rect 1247 935 1281 969
rect 1316 935 1350 969
rect 1385 935 1419 969
rect 1454 935 1488 969
rect 1523 935 1557 969
rect 1592 935 1626 969
rect 1661 935 1695 969
rect 1730 935 1764 969
rect 1799 935 1833 969
rect 1868 935 1902 969
rect 1937 935 1971 969
rect 2006 935 2040 969
rect 2075 935 2109 969
rect 2144 935 2178 969
rect 2213 935 2247 969
rect 2282 935 2316 969
rect 2351 935 14557 969
rect 2351 901 14523 935
rect 14591 901 14625 935
rect 730 867 764 901
rect 799 867 833 901
rect 868 867 902 901
rect 937 867 971 901
rect 1006 867 1040 901
rect 1075 867 1109 901
rect 1144 867 1178 901
rect 1213 867 1247 901
rect 1282 867 1316 901
rect 1351 867 1385 901
rect 1420 867 1454 901
rect 1489 867 1523 901
rect 1558 867 1592 901
rect 1627 867 1661 901
rect 1696 867 1730 901
rect 1765 867 1799 901
rect 1834 867 1868 901
rect 1903 867 1937 901
rect 1972 867 2006 901
rect 2041 867 2075 901
rect 2110 867 2144 901
rect 2179 867 2213 901
rect 2248 867 2282 901
rect 2317 867 14523 901
<< mvnsubdiffcont >>
rect 24370 9157 24540 9395
rect 24370 9087 24404 9121
rect 24438 9087 24472 9121
rect 24506 9087 24540 9121
rect 24370 9017 24404 9051
rect 24438 9017 24472 9051
rect 24506 9017 24540 9051
rect 24370 8947 24404 8981
rect 24438 8947 24472 8981
rect 24506 8947 24540 8981
rect 24370 8878 24404 8912
rect 24438 8878 24472 8912
rect 24506 8878 24540 8912
rect 24370 8809 24404 8843
rect 24438 8809 24472 8843
rect 24506 8809 24540 8843
rect 24370 8740 24404 8774
rect 24438 8740 24472 8774
rect 24506 8740 24540 8774
rect 24370 8671 24404 8705
rect 24438 8671 24472 8705
rect 24506 8671 24540 8705
rect 24370 8602 24540 8636
rect 24370 8568 24537 8602
rect 23755 8534 23789 8568
rect 23823 8534 23857 8568
rect 23891 8534 23925 8568
rect 23959 8534 23993 8568
rect 24027 8534 24061 8568
rect 24095 8534 24129 8568
rect 24163 8534 24197 8568
rect 24231 8534 24265 8568
rect 24299 8534 24333 8568
rect 24367 8534 24537 8568
rect 23755 8465 23789 8499
rect 23823 8465 23857 8499
rect 23891 8465 23925 8499
rect 23959 8465 23993 8499
rect 24027 8465 24061 8499
rect 24095 8465 24129 8499
rect 24163 8465 24197 8499
rect 24231 8465 24265 8499
rect 24299 8465 24333 8499
rect 24367 8465 24401 8499
rect 24435 8465 24469 8499
rect 24503 8465 24537 8499
rect 23755 8396 23789 8430
rect 23823 8396 23857 8430
rect 23891 8396 23925 8430
rect 23959 8396 23993 8430
rect 24027 8396 24061 8430
rect 24095 8396 24129 8430
rect 24163 8396 24197 8430
rect 24231 8396 24265 8430
rect 24299 8396 24333 8430
rect 24367 8396 24401 8430
rect 24435 8396 24469 8430
rect 24503 8396 24537 8430
rect 23755 8327 23789 8361
rect 23823 8327 23857 8361
rect 23891 8327 23925 8361
rect 23959 8327 23993 8361
rect 24027 8327 24061 8361
rect 24095 8327 24129 8361
rect 24163 8327 24197 8361
rect 24231 8327 24265 8361
rect 24299 8327 24333 8361
rect 24367 8327 24401 8361
rect 24435 8327 24469 8361
rect 24503 8327 24537 8361
rect 23755 8258 23789 8292
rect 23823 8258 23857 8292
rect 23891 8258 23925 8292
rect 23959 8258 23993 8292
rect 24027 8258 24061 8292
rect 24095 8258 24129 8292
rect 24163 8258 24197 8292
rect 24231 8258 24265 8292
rect 24299 8258 24333 8292
rect 24367 8258 24401 8292
rect 24435 8258 24469 8292
rect 24503 8258 24537 8292
rect 23755 8189 23789 8223
rect 23823 8189 23857 8223
rect 23891 8189 23925 8223
rect 23959 8189 23993 8223
rect 24027 8189 24061 8223
rect 24095 8189 24129 8223
rect 24163 8189 24197 8223
rect 24231 8189 24265 8223
rect 24299 8189 24333 8223
rect 24367 8189 24401 8223
rect 24435 8189 24469 8223
rect 24503 8189 24537 8223
rect 23755 8120 23789 8154
rect 23823 8120 23857 8154
rect 23891 8120 23925 8154
rect 23959 8120 23993 8154
rect 24027 8120 24061 8154
rect 24095 8120 24129 8154
rect 24163 8120 24197 8154
rect 24231 8120 24265 8154
rect 24299 8120 24333 8154
rect 24367 8120 24401 8154
rect 24435 8120 24469 8154
rect 24503 8120 24537 8154
rect 23755 8051 23789 8085
rect 23823 8051 23857 8085
rect 23891 8051 23925 8085
rect 23959 8051 23993 8085
rect 24027 8051 24061 8085
rect 24095 8051 24129 8085
rect 24163 8051 24197 8085
rect 24231 8051 24265 8085
rect 24299 8051 24333 8085
rect 24367 8051 24401 8085
rect 24435 8051 24469 8085
rect 24503 8051 24537 8085
rect 23755 7982 23789 8016
rect 23823 7982 23857 8016
rect 23891 7982 23925 8016
rect 23959 7982 23993 8016
rect 24027 7982 24061 8016
rect 24095 7982 24129 8016
rect 24163 7982 24197 8016
rect 24231 7982 24265 8016
rect 24299 7982 24333 8016
rect 24367 7982 24401 8016
rect 24435 7982 24469 8016
rect 24503 7982 24537 8016
rect 23755 7913 23789 7947
rect 23823 7913 23857 7947
rect 23891 7913 23925 7947
rect 23959 7913 23993 7947
rect 24027 7913 24061 7947
rect 24095 7913 24129 7947
rect 24163 7913 24197 7947
rect 24231 7913 24265 7947
rect 24299 7913 24333 7947
rect 24367 7913 24401 7947
rect 24435 7913 24469 7947
rect 24503 7913 24537 7947
rect 23755 7844 23789 7878
rect 23823 7844 23857 7878
rect 23891 7844 23925 7878
rect 23959 7844 23993 7878
rect 24027 7844 24061 7878
rect 24095 7844 24129 7878
rect 24163 7844 24197 7878
rect 24231 7844 24265 7878
rect 24299 7844 24333 7878
rect 24367 7844 24401 7878
rect 24435 7844 24469 7878
rect 24503 7844 24537 7878
rect 23755 7775 23789 7809
rect 23823 7775 23857 7809
rect 23891 7775 23925 7809
rect 23959 7775 23993 7809
rect 24027 7775 24061 7809
rect 24095 7775 24129 7809
rect 24163 7775 24197 7809
rect 24231 7775 24265 7809
rect 24299 7775 24333 7809
rect 24367 7775 24401 7809
rect 24435 7775 24469 7809
rect 24503 7775 24537 7809
rect 23755 7706 23789 7740
rect 23823 7706 23857 7740
rect 23891 7706 23925 7740
rect 23959 7706 23993 7740
rect 24027 7706 24061 7740
rect 24095 7706 24129 7740
rect 24163 7706 24197 7740
rect 24231 7706 24265 7740
rect 24299 7706 24333 7740
rect 24367 7706 24401 7740
rect 24435 7706 24469 7740
rect 24503 7706 24537 7740
rect 23755 7637 23789 7671
rect 23823 7637 23857 7671
rect 23891 7637 23925 7671
rect 23959 7637 23993 7671
rect 24027 7637 24061 7671
rect 24095 7637 24129 7671
rect 24163 7637 24197 7671
rect 24231 7637 24265 7671
rect 24299 7637 24333 7671
rect 24367 7637 24401 7671
rect 24435 7637 24469 7671
rect 24503 7637 24537 7671
rect 23755 7568 23789 7602
rect 23823 7568 23857 7602
rect 23891 7568 23925 7602
rect 23959 7568 23993 7602
rect 24027 7568 24061 7602
rect 24095 7568 24129 7602
rect 24163 7568 24197 7602
rect 24231 7568 24265 7602
rect 24299 7568 24333 7602
rect 24367 7568 24401 7602
rect 24435 7568 24469 7602
rect 24503 7568 24537 7602
rect 23755 7499 23789 7533
rect 23823 7499 23857 7533
rect 23891 7499 23925 7533
rect 23959 7499 23993 7533
rect 24027 7499 24061 7533
rect 24095 7499 24129 7533
rect 24163 7499 24197 7533
rect 24231 7499 24265 7533
rect 24299 7499 24333 7533
rect 24367 7499 24401 7533
rect 24435 7499 24469 7533
rect 24503 7499 24537 7533
rect 23755 7430 23789 7464
rect 23823 7430 23857 7464
rect 23891 7430 23925 7464
rect 23959 7430 23993 7464
rect 24027 7430 24061 7464
rect 24095 7430 24129 7464
rect 24163 7430 24197 7464
rect 24231 7430 24265 7464
rect 24299 7430 24333 7464
rect 24367 7430 24401 7464
rect 24435 7430 24469 7464
rect 24503 7430 24537 7464
rect 23755 7361 23789 7395
rect 23823 7361 23857 7395
rect 23891 7361 23925 7395
rect 23959 7361 23993 7395
rect 24027 7361 24061 7395
rect 24095 7361 24129 7395
rect 24163 7361 24197 7395
rect 24231 7361 24265 7395
rect 24299 7361 24333 7395
rect 24367 7361 24401 7395
rect 24435 7361 24469 7395
rect 24503 7361 24537 7395
rect 23755 7292 23789 7326
rect 23823 7292 23857 7326
rect 23891 7292 23925 7326
rect 23959 7292 23993 7326
rect 24027 7292 24061 7326
rect 24095 7292 24129 7326
rect 24163 7292 24197 7326
rect 24231 7292 24265 7326
rect 24299 7292 24333 7326
rect 24367 7292 24401 7326
rect 24435 7292 24469 7326
rect 24503 7292 24537 7326
rect 23755 7223 23789 7257
rect 23823 7223 23857 7257
rect 23891 7223 23925 7257
rect 23959 7223 23993 7257
rect 24027 7223 24061 7257
rect 24095 7223 24129 7257
rect 24163 7223 24197 7257
rect 24231 7223 24265 7257
rect 24299 7223 24333 7257
rect 24367 7223 24401 7257
rect 24435 7223 24469 7257
rect 24503 7223 24537 7257
rect 23755 7154 23789 7188
rect 23823 7154 23857 7188
rect 23891 7154 23925 7188
rect 23959 7154 23993 7188
rect 24027 7154 24061 7188
rect 24095 7154 24129 7188
rect 24163 7154 24197 7188
rect 24231 7154 24265 7188
rect 24299 7154 24333 7188
rect 24367 7154 24401 7188
rect 24435 7154 24469 7188
rect 24503 7154 24537 7188
rect 23755 7085 23789 7119
rect 23823 7085 23857 7119
rect 23891 7085 23925 7119
rect 23959 7085 23993 7119
rect 24027 7085 24061 7119
rect 24095 7085 24129 7119
rect 24163 7085 24197 7119
rect 24231 7085 24265 7119
rect 24299 7085 24333 7119
rect 24367 7085 24401 7119
rect 24435 7085 24469 7119
rect 24503 7085 24537 7119
rect 23755 7016 23789 7050
rect 23823 7016 23857 7050
rect 23891 7016 23925 7050
rect 23959 7016 23993 7050
rect 24027 7016 24061 7050
rect 24095 7016 24129 7050
rect 24163 7016 24197 7050
rect 24231 7016 24265 7050
rect 24299 7016 24333 7050
rect 24367 7016 24401 7050
rect 24435 7016 24469 7050
rect 24503 7016 24537 7050
rect 23755 6947 23789 6981
rect 23823 6947 23857 6981
rect 23891 6947 23925 6981
rect 23959 6947 23993 6981
rect 24027 6947 24061 6981
rect 24095 6947 24129 6981
rect 24163 6947 24197 6981
rect 24231 6947 24265 6981
rect 24299 6947 24333 6981
rect 24367 6947 24401 6981
rect 24435 6947 24469 6981
rect 24503 6947 24537 6981
rect 23755 6878 23789 6912
rect 23823 6878 23857 6912
rect 23891 6878 23925 6912
rect 23959 6878 23993 6912
rect 24027 6878 24061 6912
rect 24095 6878 24129 6912
rect 24163 6878 24197 6912
rect 24231 6878 24265 6912
rect 24299 6878 24333 6912
rect 24367 6878 24401 6912
rect 24435 6878 24469 6912
rect 24503 6878 24537 6912
rect 23755 6809 23789 6843
rect 23823 6809 23857 6843
rect 23891 6809 23925 6843
rect 23959 6809 23993 6843
rect 24027 6809 24061 6843
rect 24095 6809 24129 6843
rect 24163 6809 24197 6843
rect 24231 6809 24265 6843
rect 24299 6809 24333 6843
rect 24367 6809 24401 6843
rect 24435 6809 24469 6843
rect 24503 6809 24537 6843
rect 23755 6740 23789 6774
rect 23823 6740 23857 6774
rect 23891 6740 23925 6774
rect 23959 6740 23993 6774
rect 24027 6740 24061 6774
rect 24095 6740 24129 6774
rect 24163 6740 24197 6774
rect 24231 6740 24265 6774
rect 24299 6740 24333 6774
rect 24367 6740 24401 6774
rect 24435 6740 24469 6774
rect 24503 6740 24537 6774
rect 23755 6671 23789 6705
rect 23823 6671 23857 6705
rect 23891 6671 23925 6705
rect 23959 6671 23993 6705
rect 24027 6671 24061 6705
rect 24095 6671 24129 6705
rect 24163 6671 24197 6705
rect 24231 6671 24265 6705
rect 24299 6671 24333 6705
rect 24367 6671 24401 6705
rect 24435 6671 24469 6705
rect 24503 6671 24537 6705
rect 23755 6602 23789 6636
rect 23823 6602 23857 6636
rect 23891 6602 23925 6636
rect 23959 6602 23993 6636
rect 24027 6602 24061 6636
rect 24095 6602 24129 6636
rect 24163 6602 24197 6636
rect 24231 6602 24265 6636
rect 24299 6602 24333 6636
rect 24367 6602 24401 6636
rect 24435 6602 24469 6636
rect 24503 6602 24537 6636
rect 23755 6533 23789 6567
rect 23823 6533 23857 6567
rect 23891 6533 23925 6567
rect 23959 6533 23993 6567
rect 24027 6533 24061 6567
rect 24095 6533 24129 6567
rect 24163 6533 24197 6567
rect 24231 6533 24265 6567
rect 24299 6533 24333 6567
rect 24367 6533 24401 6567
rect 24435 6533 24469 6567
rect 24503 6533 24537 6567
rect 23755 6464 23789 6498
rect 23823 6464 23857 6498
rect 23891 6464 23925 6498
rect 23959 6464 23993 6498
rect 24027 6464 24061 6498
rect 24095 6464 24129 6498
rect 24163 6464 24197 6498
rect 24231 6464 24265 6498
rect 24299 6464 24333 6498
rect 24367 6464 24401 6498
rect 24435 6464 24469 6498
rect 24503 6464 24537 6498
rect 23755 6395 23789 6429
rect 23823 6395 23857 6429
rect 23891 6395 23925 6429
rect 23959 6395 23993 6429
rect 24027 6395 24061 6429
rect 24095 6395 24129 6429
rect 24163 6395 24197 6429
rect 24231 6395 24265 6429
rect 24299 6395 24333 6429
rect 24367 6395 24401 6429
rect 24435 6395 24469 6429
rect 24503 6395 24537 6429
rect 23755 6326 23789 6360
rect 23823 6326 23857 6360
rect 23891 6326 23925 6360
rect 23959 6326 23993 6360
rect 24027 6326 24061 6360
rect 24095 6326 24129 6360
rect 24163 6326 24197 6360
rect 24231 6326 24265 6360
rect 24299 6326 24333 6360
rect 24367 6326 24401 6360
rect 24435 6326 24469 6360
rect 24503 6326 24537 6360
rect 23755 6257 23789 6291
rect 23823 6257 23857 6291
rect 23891 6257 23925 6291
rect 23959 6257 23993 6291
rect 24027 6257 24061 6291
rect 24095 6257 24129 6291
rect 24163 6257 24197 6291
rect 24231 6257 24265 6291
rect 24299 6257 24333 6291
rect 24367 6257 24401 6291
rect 24435 6257 24469 6291
rect 24503 6257 24537 6291
rect 23755 6188 23789 6222
rect 23823 6188 23857 6222
rect 23891 6188 23925 6222
rect 23959 6188 23993 6222
rect 24027 6188 24061 6222
rect 24095 6188 24129 6222
rect 24163 6188 24197 6222
rect 24231 6188 24265 6222
rect 24299 6188 24333 6222
rect 24367 6188 24401 6222
rect 24435 6188 24469 6222
rect 24503 6188 24537 6222
rect 23755 6119 23789 6153
rect 23823 6119 23857 6153
rect 23891 6119 23925 6153
rect 23959 6119 23993 6153
rect 24027 6119 24061 6153
rect 24095 6119 24129 6153
rect 24163 6119 24197 6153
rect 24231 6119 24265 6153
rect 24299 6119 24333 6153
rect 24367 6119 24401 6153
rect 24435 6119 24469 6153
rect 24503 6119 24537 6153
rect 23755 6050 23789 6084
rect 23823 6050 23857 6084
rect 23891 6050 23925 6084
rect 23959 6050 23993 6084
rect 24027 6050 24061 6084
rect 24095 6050 24129 6084
rect 24163 6050 24197 6084
rect 24231 6050 24265 6084
rect 24299 6050 24333 6084
rect 24367 6050 24401 6084
rect 24435 6050 24469 6084
rect 24503 6050 24537 6084
rect 23755 5981 23789 6015
rect 23823 5981 23857 6015
rect 23891 5981 23925 6015
rect 23959 5981 23993 6015
rect 24027 5981 24061 6015
rect 24095 5981 24129 6015
rect 24163 5981 24197 6015
rect 24231 5981 24265 6015
rect 24299 5981 24333 6015
rect 24367 5981 24401 6015
rect 24435 5981 24469 6015
rect 24503 5981 24537 6015
rect 23755 5912 23789 5946
rect 23823 5912 23857 5946
rect 23891 5912 23925 5946
rect 23959 5912 23993 5946
rect 24027 5912 24061 5946
rect 24095 5912 24129 5946
rect 24163 5912 24197 5946
rect 24231 5912 24265 5946
rect 24299 5912 24333 5946
rect 24367 5912 24401 5946
rect 24435 5912 24469 5946
rect 24503 5912 24537 5946
rect 23755 5639 24537 5877
rect 24153 5557 24187 5591
rect 24221 5557 24255 5591
rect 24289 5557 24323 5591
rect 24357 5557 24391 5591
rect 24425 5557 24459 5591
rect 24493 5557 24527 5591
rect 278 4449 312 4483
rect 346 4449 380 4483
rect 414 4449 448 4483
rect 278 4379 312 4413
rect 346 4379 380 4413
rect 414 4379 448 4413
rect 278 4309 312 4343
rect 346 4309 380 4343
rect 414 4309 448 4343
rect 278 4239 312 4273
rect 346 4239 380 4273
rect 414 4239 448 4273
rect 278 4169 312 4203
rect 346 4169 380 4203
rect 414 4169 448 4203
rect 278 4100 312 4134
rect 346 4100 380 4134
rect 414 4100 448 4134
rect 278 4031 312 4065
rect 346 4031 380 4065
rect 414 4031 448 4065
rect 278 3962 312 3996
rect 346 3962 380 3996
rect 414 3962 448 3996
rect 278 3893 312 3927
rect 346 3893 380 3927
rect 414 3893 448 3927
rect 278 3824 312 3858
rect 346 3824 380 3858
rect 414 3824 448 3858
rect 278 3755 312 3789
rect 346 3755 380 3789
rect 414 3755 448 3789
rect 278 3686 312 3720
rect 346 3686 380 3720
rect 414 3686 448 3720
rect 278 3617 312 3651
rect 346 3617 380 3651
rect 414 3617 448 3651
rect 278 3548 312 3582
rect 346 3548 380 3582
rect 414 3548 448 3582
rect 278 3479 312 3513
rect 346 3479 380 3513
rect 414 3479 448 3513
rect 278 3410 312 3444
rect 346 3410 380 3444
rect 414 3410 448 3444
rect 278 3341 312 3375
rect 346 3341 380 3375
rect 414 3341 448 3375
rect 278 3272 312 3306
rect 346 3272 380 3306
rect 414 3272 448 3306
rect 278 3203 312 3237
rect 346 3203 380 3237
rect 414 3203 448 3237
rect 278 3134 312 3168
rect 346 3134 380 3168
rect 414 3134 448 3168
rect 278 3065 312 3099
rect 346 3065 380 3099
rect 414 3065 448 3099
rect 278 2996 312 3030
rect 346 2996 380 3030
rect 414 2996 448 3030
rect 278 2927 312 2961
rect 346 2927 380 2961
rect 414 2927 448 2961
rect 278 2858 312 2892
rect 346 2858 380 2892
rect 414 2858 448 2892
rect 278 2789 312 2823
rect 346 2789 380 2823
rect 414 2789 448 2823
rect 278 2720 312 2754
rect 346 2720 380 2754
rect 414 2720 448 2754
rect 278 2651 312 2685
rect 346 2651 380 2685
rect 414 2651 448 2685
rect 278 2582 312 2616
rect 346 2582 380 2616
rect 414 2582 448 2616
rect 278 2513 312 2547
rect 346 2513 380 2547
rect 414 2513 448 2547
rect 278 2444 312 2478
rect 346 2444 380 2478
rect 414 2444 448 2478
rect 278 2375 312 2409
rect 346 2375 380 2409
rect 414 2375 448 2409
rect 278 2306 312 2340
rect 346 2306 380 2340
rect 414 2306 448 2340
rect 278 2237 312 2271
rect 346 2237 380 2271
rect 414 2237 448 2271
rect 278 2168 312 2202
rect 346 2168 380 2202
rect 414 2168 448 2202
rect 278 2099 312 2133
rect 346 2099 380 2133
rect 414 2099 448 2133
rect 278 2030 312 2064
rect 346 2030 380 2064
rect 414 2030 448 2064
rect 278 1961 312 1995
rect 346 1961 380 1995
rect 414 1961 448 1995
rect 278 1892 312 1926
rect 346 1892 380 1926
rect 414 1892 448 1926
rect 278 1823 312 1857
rect 346 1823 380 1857
rect 414 1823 448 1857
rect 278 1754 312 1788
rect 346 1754 380 1788
rect 414 1754 448 1788
rect 278 1685 312 1719
rect 346 1685 380 1719
rect 414 1685 448 1719
rect 278 1616 312 1650
rect 346 1616 380 1650
rect 414 1616 448 1650
rect 278 1547 312 1581
rect 346 1547 380 1581
rect 414 1547 448 1581
rect 278 1478 312 1512
rect 346 1478 380 1512
rect 414 1478 448 1512
rect 278 1409 312 1443
rect 346 1409 380 1443
rect 414 1409 448 1443
rect 278 1340 312 1374
rect 346 1340 380 1374
rect 414 1340 448 1374
rect 278 1271 312 1305
rect 346 1271 380 1305
rect 414 1271 448 1305
rect 278 1202 312 1236
rect 346 1202 380 1236
rect 414 1202 448 1236
rect 278 1133 312 1167
rect 346 1133 380 1167
rect 414 1133 448 1167
rect 278 1064 312 1098
rect 346 1064 380 1098
rect 414 1064 448 1098
rect 278 995 312 1029
rect 346 995 380 1029
rect 414 995 448 1029
rect 278 926 312 960
rect 346 926 380 960
rect 414 926 448 960
rect 278 857 312 891
rect 346 857 380 891
rect 414 857 448 891
rect 1086 4516 1120 4550
rect 1154 4516 1188 4550
rect 1222 4516 1256 4550
rect 1290 4516 1324 4550
rect 1358 4516 1392 4550
rect 1426 4516 1460 4550
rect 1507 4506 1541 4540
rect 1609 4506 6335 4574
rect 6370 4540 6404 4574
rect 6439 4540 6473 4574
rect 6508 4540 6542 4574
rect 6577 4540 6611 4574
rect 6646 4540 6680 4574
rect 6715 4540 6749 4574
rect 6784 4540 6818 4574
rect 6853 4540 6887 4574
rect 6922 4540 6956 4574
rect 6991 4540 7025 4574
rect 7060 4540 7094 4574
rect 7129 4540 7163 4574
rect 7198 4540 7232 4574
rect 7267 4540 7301 4574
rect 7336 4540 7370 4574
rect 7405 4540 7439 4574
rect 7474 4540 7508 4574
rect 7543 4540 7577 4574
rect 7612 4540 7646 4574
rect 7681 4540 7715 4574
rect 7750 4540 7784 4574
rect 7819 4540 7853 4574
rect 7888 4540 7922 4574
rect 7957 4540 7991 4574
rect 8026 4540 8060 4574
rect 8095 4540 8129 4574
rect 8164 4540 8198 4574
rect 8233 4540 8267 4574
rect 8302 4540 8336 4574
rect 8371 4540 8405 4574
rect 8440 4540 8474 4574
rect 8509 4540 8543 4574
rect 8578 4540 8612 4574
rect 8647 4540 8681 4574
rect 8716 4540 8750 4574
rect 8785 4540 8819 4574
rect 8854 4540 8888 4574
rect 8923 4540 8957 4574
rect 8992 4540 9026 4574
rect 9061 4540 9095 4574
rect 9130 4540 9164 4574
rect 9199 4540 9233 4574
rect 9268 4540 9302 4574
rect 9337 4540 9371 4574
rect 9406 4540 9440 4574
rect 9475 4540 9509 4574
rect 9544 4540 9578 4574
rect 9613 4540 9647 4574
rect 9682 4540 9716 4574
rect 9751 4540 9785 4574
rect 9820 4540 9854 4574
rect 9889 4540 9923 4574
rect 9958 4540 9992 4574
rect 1086 4447 1120 4481
rect 1154 4447 1188 4481
rect 1222 4447 1256 4481
rect 1290 4447 1324 4481
rect 1358 4447 1392 4481
rect 1426 4447 1460 4481
rect 1575 4472 8681 4506
rect 8716 4472 8750 4506
rect 8785 4472 8819 4506
rect 8854 4472 8888 4506
rect 8923 4472 8957 4506
rect 8992 4472 9026 4506
rect 9061 4472 9095 4506
rect 9130 4472 9164 4506
rect 9199 4472 9233 4506
rect 9268 4472 9302 4506
rect 9337 4472 9371 4506
rect 9406 4472 9440 4506
rect 9475 4472 9509 4506
rect 9544 4472 9578 4506
rect 9613 4472 9647 4506
rect 9682 4472 9716 4506
rect 9751 4472 9785 4506
rect 9820 4472 9854 4506
rect 9889 4472 9923 4506
rect 9958 4472 9992 4506
rect 1507 4437 1541 4471
rect 1086 4378 1120 4412
rect 1154 4378 1188 4412
rect 1222 4378 1256 4412
rect 1290 4378 1324 4412
rect 1358 4378 1392 4412
rect 1426 4378 1460 4412
rect 1575 4402 1609 4436
rect 1643 4404 8681 4472
rect 8716 4404 8750 4438
rect 8785 4404 8819 4438
rect 8854 4404 8888 4438
rect 8923 4404 8957 4438
rect 8992 4404 9026 4438
rect 9061 4404 9095 4438
rect 9130 4404 9164 4438
rect 9199 4404 9233 4438
rect 9268 4404 9302 4438
rect 9337 4404 9371 4438
rect 9406 4404 9440 4438
rect 9475 4404 9509 4438
rect 9544 4404 9578 4438
rect 9613 4404 9647 4438
rect 9682 4404 9716 4438
rect 9751 4404 9785 4438
rect 9820 4404 9854 4438
rect 9889 4404 9923 4438
rect 9958 4404 9992 4438
rect 1507 4368 1541 4402
rect 1086 4309 1120 4343
rect 1154 4309 1188 4343
rect 1222 4309 1256 4343
rect 1290 4309 1324 4343
rect 1358 4309 1392 4343
rect 1426 4309 1460 4343
rect 1507 4299 1541 4333
rect 1575 4332 1609 4366
rect 1643 4334 1677 4368
rect 1711 4325 1745 4359
rect 1780 4325 1814 4359
rect 1849 4325 1883 4359
rect 1918 4325 1952 4359
rect 1987 4325 2021 4359
rect 2056 4325 2090 4359
rect 2125 4325 2159 4359
rect 2194 4325 2228 4359
rect 2263 4325 2297 4359
rect 2332 4325 2366 4359
rect 1086 4240 1120 4274
rect 1154 4240 1188 4274
rect 1222 4240 1256 4274
rect 1290 4240 1324 4274
rect 1358 4240 1392 4274
rect 1426 4240 1460 4274
rect 1507 4230 1541 4264
rect 1575 4262 1609 4296
rect 1643 4264 1677 4298
rect 1711 4257 1745 4291
rect 1780 4257 1814 4291
rect 1849 4257 1883 4291
rect 1918 4257 1952 4291
rect 1987 4257 2021 4291
rect 2056 4257 2090 4291
rect 2125 4257 2159 4291
rect 2194 4257 2228 4291
rect 2263 4257 2297 4291
rect 2332 4257 2366 4291
rect 1086 4171 1120 4205
rect 1154 4171 1188 4205
rect 1222 4171 1256 4205
rect 1290 4171 1324 4205
rect 1358 4171 1392 4205
rect 1426 4171 1460 4205
rect 1507 4161 1541 4195
rect 1575 4192 1609 4226
rect 1643 4194 1677 4228
rect 1711 4189 1745 4223
rect 1780 4189 1814 4223
rect 1849 4189 1883 4223
rect 1918 4189 1952 4223
rect 1987 4189 2021 4223
rect 2056 4189 2090 4223
rect 2125 4189 2159 4223
rect 2194 4189 2228 4223
rect 2263 4189 2297 4223
rect 2332 4189 2366 4223
rect 2401 4189 4135 4359
rect 8643 4336 8681 4404
rect 8711 4336 8745 4370
rect 8779 4336 8813 4370
rect 8847 4336 8881 4370
rect 8915 4336 8949 4370
rect 8983 4336 9017 4370
rect 9051 4336 9085 4370
rect 9119 4336 9153 4370
rect 9187 4336 9221 4370
rect 9255 4336 9289 4370
rect 9323 4336 9357 4370
rect 9391 4336 9425 4370
rect 9459 4336 9493 4370
rect 9527 4336 9561 4370
rect 9595 4336 9629 4370
rect 9663 4336 9697 4370
rect 9731 4336 9765 4370
rect 9799 4336 9833 4370
rect 9867 4336 9901 4370
rect 9935 4336 9969 4370
rect 10003 4336 10037 4370
rect 10071 4336 10105 4370
rect 10139 4336 10173 4370
rect 10207 4336 10241 4370
rect 10312 4337 10346 4371
rect 10380 4337 10414 4371
rect 10448 4337 10482 4371
rect 10516 4337 10550 4371
rect 10584 4337 10618 4371
rect 10652 4337 10686 4371
rect 10720 4337 10754 4371
rect 10788 4337 10822 4371
rect 10856 4337 10890 4371
rect 10924 4337 10958 4371
rect 10992 4337 11026 4371
rect 11060 4337 11094 4371
rect 11128 4337 11162 4371
rect 11196 4337 11230 4371
rect 11264 4337 11298 4371
rect 11332 4337 11366 4371
rect 11400 4337 11434 4371
rect 11468 4337 11502 4371
rect 11536 4337 11570 4371
rect 4179 4300 4213 4334
rect 4248 4300 4282 4334
rect 4317 4300 4351 4334
rect 4386 4300 4420 4334
rect 4455 4300 4489 4334
rect 4524 4300 4558 4334
rect 4593 4300 4627 4334
rect 4662 4300 4696 4334
rect 4731 4300 4765 4334
rect 4800 4300 4834 4334
rect 4869 4300 4903 4334
rect 4938 4300 4972 4334
rect 5007 4300 5041 4334
rect 5076 4300 5110 4334
rect 5145 4300 5179 4334
rect 5214 4300 5248 4334
rect 5283 4300 5317 4334
rect 5352 4300 5386 4334
rect 5421 4300 5455 4334
rect 4179 4232 4213 4266
rect 4248 4232 4282 4266
rect 4317 4232 4351 4266
rect 4386 4232 4420 4266
rect 4455 4232 4489 4266
rect 4524 4232 4558 4266
rect 4593 4232 4627 4266
rect 4662 4232 4696 4266
rect 4731 4232 4765 4266
rect 4800 4232 4834 4266
rect 4869 4232 4903 4266
rect 4938 4232 4972 4266
rect 5007 4232 5041 4266
rect 5076 4232 5110 4266
rect 5145 4232 5179 4266
rect 5214 4232 5248 4266
rect 5283 4232 5317 4266
rect 5352 4232 5386 4266
rect 5421 4232 5455 4266
rect 1086 4102 1120 4136
rect 1154 4102 1188 4136
rect 1222 4102 1256 4136
rect 1290 4102 1324 4136
rect 1358 4102 1392 4136
rect 1426 4102 1460 4136
rect 1507 4092 1541 4126
rect 1575 4122 1609 4156
rect 1643 4124 1677 4158
rect 4179 4164 4213 4198
rect 4248 4164 4282 4198
rect 4317 4164 4351 4198
rect 4386 4164 4420 4198
rect 4455 4164 4489 4198
rect 4524 4164 4558 4198
rect 4593 4164 4627 4198
rect 4662 4164 4696 4198
rect 4731 4164 4765 4198
rect 4800 4164 4834 4198
rect 4869 4164 4903 4198
rect 4938 4164 4972 4198
rect 5007 4164 5041 4198
rect 5076 4164 5110 4198
rect 5145 4164 5179 4198
rect 5214 4164 5248 4198
rect 5283 4164 5317 4198
rect 5352 4164 5386 4198
rect 5421 4164 5455 4198
rect 4179 4096 4213 4130
rect 4248 4096 4282 4130
rect 4317 4096 4351 4130
rect 4386 4096 4420 4130
rect 4455 4096 4489 4130
rect 4524 4096 4558 4130
rect 4593 4096 4627 4130
rect 4662 4096 4696 4130
rect 4731 4096 4765 4130
rect 4800 4096 4834 4130
rect 4869 4096 4903 4130
rect 4938 4096 4972 4130
rect 5007 4096 5041 4130
rect 5076 4096 5110 4130
rect 5145 4096 5179 4130
rect 5214 4096 5248 4130
rect 5283 4096 5317 4130
rect 5352 4096 5386 4130
rect 5421 4096 5455 4130
rect 1086 4033 1120 4067
rect 1154 4033 1188 4067
rect 1222 4033 1256 4067
rect 1290 4033 1324 4067
rect 1358 4033 1392 4067
rect 1426 4033 1460 4067
rect 1507 4023 1541 4057
rect 1575 4052 1609 4086
rect 1643 4054 1677 4088
rect 1086 3964 1120 3998
rect 1154 3964 1188 3998
rect 1222 3964 1256 3998
rect 1290 3964 1324 3998
rect 1358 3964 1392 3998
rect 1426 3964 1460 3998
rect 1507 3954 1541 3988
rect 1575 3982 1609 4016
rect 1643 3984 1677 4018
rect 4179 4028 4213 4062
rect 4248 4028 4282 4062
rect 4317 4028 4351 4062
rect 4386 4028 4420 4062
rect 4455 4028 4489 4062
rect 4524 4028 4558 4062
rect 4593 4028 4627 4062
rect 4662 4028 4696 4062
rect 4731 4028 4765 4062
rect 4800 4028 4834 4062
rect 4869 4028 4903 4062
rect 4938 4028 4972 4062
rect 5007 4028 5041 4062
rect 5076 4028 5110 4062
rect 5145 4028 5179 4062
rect 5214 4028 5248 4062
rect 5283 4028 5317 4062
rect 5352 4028 5386 4062
rect 5421 4028 5455 4062
rect 1086 3895 1120 3929
rect 1154 3895 1188 3929
rect 1222 3895 1256 3929
rect 1290 3895 1324 3929
rect 1358 3895 1392 3929
rect 1426 3895 1460 3929
rect 1507 3885 1541 3919
rect 1575 3912 1609 3946
rect 1643 3914 1677 3948
rect 1086 3826 1120 3860
rect 1154 3826 1188 3860
rect 1222 3826 1256 3860
rect 1290 3826 1324 3860
rect 1358 3826 1392 3860
rect 1426 3826 1460 3860
rect 1507 3816 1541 3850
rect 1575 3842 1609 3876
rect 1643 3844 1677 3878
rect 4179 3960 4213 3994
rect 4248 3960 4282 3994
rect 4317 3960 4351 3994
rect 4386 3960 4420 3994
rect 4455 3960 4489 3994
rect 4524 3960 4558 3994
rect 4593 3960 4627 3994
rect 4662 3960 4696 3994
rect 4731 3960 4765 3994
rect 4800 3960 4834 3994
rect 4869 3960 4903 3994
rect 4938 3960 4972 3994
rect 5007 3960 5041 3994
rect 5076 3960 5110 3994
rect 5145 3960 5179 3994
rect 5214 3960 5248 3994
rect 5283 3960 5317 3994
rect 5352 3960 5386 3994
rect 5421 3960 5455 3994
rect 4179 3892 4213 3926
rect 4248 3892 4282 3926
rect 4317 3892 4351 3926
rect 4386 3892 4420 3926
rect 4455 3892 4489 3926
rect 4524 3892 4558 3926
rect 4593 3892 4627 3926
rect 4662 3892 4696 3926
rect 4731 3892 4765 3926
rect 4800 3892 4834 3926
rect 4869 3892 4903 3926
rect 4938 3892 4972 3926
rect 5007 3892 5041 3926
rect 5076 3892 5110 3926
rect 5145 3892 5179 3926
rect 5214 3892 5248 3926
rect 5283 3892 5317 3926
rect 5352 3892 5386 3926
rect 5421 3892 5455 3926
rect 5490 3892 8584 4334
rect 8643 4266 8677 4300
rect 8711 4266 8745 4300
rect 8779 4266 8813 4300
rect 8847 4266 8881 4300
rect 8915 4266 8949 4300
rect 8983 4266 9017 4300
rect 9051 4266 9085 4300
rect 9119 4266 9153 4300
rect 9187 4266 9221 4300
rect 9255 4266 9289 4300
rect 9323 4266 9357 4300
rect 9391 4266 9425 4300
rect 9459 4266 9493 4300
rect 9527 4266 9561 4300
rect 9595 4266 9629 4300
rect 9663 4266 9697 4300
rect 9731 4266 9765 4300
rect 9799 4266 9833 4300
rect 9867 4266 9901 4300
rect 9935 4266 9969 4300
rect 10003 4266 10037 4300
rect 10071 4266 10105 4300
rect 10139 4266 10173 4300
rect 10207 4266 10241 4300
rect 10312 4267 10346 4301
rect 10380 4267 10414 4301
rect 10448 4267 10482 4301
rect 10516 4267 10550 4301
rect 10584 4267 10618 4301
rect 10652 4267 10686 4301
rect 10720 4267 10754 4301
rect 10788 4267 10822 4301
rect 10856 4267 10890 4301
rect 10924 4267 10958 4301
rect 10992 4267 11026 4301
rect 11060 4267 11094 4301
rect 11128 4267 11162 4301
rect 11196 4267 11230 4301
rect 11264 4267 11298 4301
rect 11332 4267 11366 4301
rect 11400 4267 11434 4301
rect 11468 4267 11502 4301
rect 11536 4267 11570 4301
rect 8643 4196 8677 4230
rect 8711 4196 8745 4230
rect 8779 4196 8813 4230
rect 8847 4196 8881 4230
rect 8915 4196 8949 4230
rect 8983 4196 9017 4230
rect 9051 4196 9085 4230
rect 9119 4196 9153 4230
rect 9187 4196 9221 4230
rect 9255 4196 9289 4230
rect 9323 4196 9357 4230
rect 9391 4196 9425 4230
rect 9459 4196 9493 4230
rect 9527 4196 9561 4230
rect 9595 4196 9629 4230
rect 9663 4196 9697 4230
rect 9731 4196 9765 4230
rect 9799 4196 9833 4230
rect 9867 4196 9901 4230
rect 9935 4196 9969 4230
rect 10003 4196 10037 4230
rect 10071 4196 10105 4230
rect 10139 4196 10173 4230
rect 10207 4196 10241 4230
rect 10312 4197 10346 4231
rect 10380 4197 10414 4231
rect 10448 4197 10482 4231
rect 10516 4197 10550 4231
rect 10584 4197 10618 4231
rect 10652 4197 10686 4231
rect 10720 4197 10754 4231
rect 10788 4197 10822 4231
rect 10856 4197 10890 4231
rect 10924 4197 10958 4231
rect 10992 4197 11026 4231
rect 11060 4197 11094 4231
rect 11128 4197 11162 4231
rect 11196 4197 11230 4231
rect 11264 4197 11298 4231
rect 11332 4197 11366 4231
rect 11400 4197 11434 4231
rect 11468 4197 11502 4231
rect 11536 4197 11570 4231
rect 8643 4126 8677 4160
rect 8711 4126 8745 4160
rect 8779 4126 8813 4160
rect 8847 4126 8881 4160
rect 8915 4126 8949 4160
rect 8983 4126 9017 4160
rect 9051 4126 9085 4160
rect 9119 4126 9153 4160
rect 9187 4126 9221 4160
rect 9255 4126 9289 4160
rect 9323 4126 9357 4160
rect 9391 4126 9425 4160
rect 9459 4126 9493 4160
rect 9527 4126 9561 4160
rect 9595 4126 9629 4160
rect 9663 4126 9697 4160
rect 9731 4126 9765 4160
rect 9799 4126 9833 4160
rect 9867 4126 9901 4160
rect 9935 4126 9969 4160
rect 10003 4126 10037 4160
rect 10071 4126 10105 4160
rect 10139 4126 10173 4160
rect 10207 4126 10241 4160
rect 10312 4127 10346 4161
rect 10380 4127 10414 4161
rect 10448 4127 10482 4161
rect 10516 4127 10550 4161
rect 10584 4127 10618 4161
rect 10652 4127 10686 4161
rect 10720 4127 10754 4161
rect 10788 4127 10822 4161
rect 10856 4127 10890 4161
rect 10924 4127 10958 4161
rect 10992 4127 11026 4161
rect 11060 4127 11094 4161
rect 11128 4127 11162 4161
rect 11196 4127 11230 4161
rect 11264 4127 11298 4161
rect 11332 4127 11366 4161
rect 11400 4127 11434 4161
rect 11468 4127 11502 4161
rect 11536 4127 11570 4161
rect 8643 4056 8677 4090
rect 8711 4056 8745 4090
rect 8779 4056 8813 4090
rect 8847 4056 8881 4090
rect 8915 4056 8949 4090
rect 8983 4056 9017 4090
rect 9051 4056 9085 4090
rect 9119 4056 9153 4090
rect 9187 4056 9221 4090
rect 9255 4056 9289 4090
rect 9323 4056 9357 4090
rect 9391 4056 9425 4090
rect 9459 4056 9493 4090
rect 9527 4056 9561 4090
rect 9595 4056 9629 4090
rect 9663 4056 9697 4090
rect 9731 4056 9765 4090
rect 9799 4056 9833 4090
rect 9867 4056 9901 4090
rect 9935 4056 9969 4090
rect 10003 4056 10037 4090
rect 10071 4056 10105 4090
rect 10139 4056 10173 4090
rect 10207 4056 10241 4090
rect 10312 4057 10346 4091
rect 10380 4057 10414 4091
rect 10448 4057 10482 4091
rect 10516 4057 10550 4091
rect 10584 4057 10618 4091
rect 10652 4057 10686 4091
rect 10720 4057 10754 4091
rect 10788 4057 10822 4091
rect 10856 4057 10890 4091
rect 10924 4057 10958 4091
rect 10992 4057 11026 4091
rect 11060 4057 11094 4091
rect 11128 4057 11162 4091
rect 11196 4057 11230 4091
rect 11264 4057 11298 4091
rect 11332 4057 11366 4091
rect 11400 4057 11434 4091
rect 11468 4057 11502 4091
rect 11536 4057 11570 4091
rect 8643 3986 8677 4020
rect 8711 3986 8745 4020
rect 8779 3986 8813 4020
rect 8847 3986 8881 4020
rect 8915 3986 8949 4020
rect 8983 3986 9017 4020
rect 9051 3986 9085 4020
rect 9119 3986 9153 4020
rect 9187 3986 9221 4020
rect 9255 3986 9289 4020
rect 9323 3986 9357 4020
rect 9391 3986 9425 4020
rect 9459 3986 9493 4020
rect 9527 3986 9561 4020
rect 9595 3986 9629 4020
rect 9663 3986 9697 4020
rect 9731 3986 9765 4020
rect 9799 3986 9833 4020
rect 9867 3986 9901 4020
rect 9935 3986 9969 4020
rect 10003 3986 10037 4020
rect 10071 3986 10105 4020
rect 10139 3986 10173 4020
rect 10207 3986 10241 4020
rect 10312 3987 10346 4021
rect 10380 3987 10414 4021
rect 10448 3987 10482 4021
rect 10516 3987 10550 4021
rect 10584 3987 10618 4021
rect 10652 3987 10686 4021
rect 10720 3987 10754 4021
rect 10788 3987 10822 4021
rect 10856 3987 10890 4021
rect 10924 3987 10958 4021
rect 10992 3987 11026 4021
rect 11060 3987 11094 4021
rect 11128 3987 11162 4021
rect 11196 3987 11230 4021
rect 11264 3987 11298 4021
rect 11332 3987 11366 4021
rect 11400 3987 11434 4021
rect 11468 3987 11502 4021
rect 11536 3987 11570 4021
rect 8643 3916 8677 3950
rect 8711 3916 8745 3950
rect 8779 3916 8813 3950
rect 8847 3916 8881 3950
rect 8915 3916 8949 3950
rect 8983 3916 9017 3950
rect 9051 3916 9085 3950
rect 9119 3916 9153 3950
rect 9187 3916 9221 3950
rect 9255 3916 9289 3950
rect 9323 3916 9357 3950
rect 9391 3916 9425 3950
rect 9459 3916 9493 3950
rect 9527 3916 9561 3950
rect 9595 3916 9629 3950
rect 9663 3916 9697 3950
rect 9731 3916 9765 3950
rect 9799 3916 9833 3950
rect 9867 3916 9901 3950
rect 9935 3916 9969 3950
rect 10003 3916 10037 3950
rect 10071 3916 10105 3950
rect 10139 3916 10173 3950
rect 10207 3916 10241 3950
rect 10312 3917 10346 3951
rect 10380 3917 10414 3951
rect 10448 3917 10482 3951
rect 10516 3917 10550 3951
rect 10584 3917 10618 3951
rect 10652 3917 10686 3951
rect 10720 3917 10754 3951
rect 10788 3917 10822 3951
rect 10856 3917 10890 3951
rect 10924 3917 10958 3951
rect 10992 3917 11026 3951
rect 11060 3917 11094 3951
rect 11128 3917 11162 3951
rect 11196 3917 11230 3951
rect 11264 3917 11298 3951
rect 11332 3917 11366 3951
rect 11400 3917 11434 3951
rect 11468 3917 11502 3951
rect 11536 3917 11570 3951
rect 1086 3757 1120 3791
rect 1154 3757 1188 3791
rect 1222 3757 1256 3791
rect 1290 3757 1324 3791
rect 1358 3757 1392 3791
rect 1426 3757 1460 3791
rect 1507 3747 1541 3781
rect 1575 3772 1609 3806
rect 1643 3774 1677 3808
rect 1086 3688 1120 3722
rect 1154 3688 1188 3722
rect 1222 3688 1256 3722
rect 1290 3688 1324 3722
rect 1358 3688 1392 3722
rect 1426 3688 1460 3722
rect 1507 3678 1541 3712
rect 1575 3702 1609 3736
rect 1643 3704 1677 3738
rect 1086 1443 1460 3653
rect 1507 3609 1541 3643
rect 1575 3632 1609 3666
rect 1643 3634 1677 3668
rect 1507 3540 1541 3574
rect 1575 3562 1609 3596
rect 1643 3564 1677 3598
rect 1507 3471 1541 3505
rect 1575 3492 1609 3526
rect 1643 3494 1677 3528
rect 1507 3402 1541 3436
rect 1575 3422 1609 3456
rect 1643 3424 1677 3458
rect 1507 3333 1541 3367
rect 1575 3352 1609 3386
rect 1643 3354 1677 3388
rect 1507 3264 1541 3298
rect 1575 3282 1609 3316
rect 1643 3284 1677 3318
rect 8643 3846 8677 3880
rect 8711 3846 8745 3880
rect 8779 3846 8813 3880
rect 8847 3846 8881 3880
rect 8915 3846 8949 3880
rect 8983 3846 9017 3880
rect 9051 3846 9085 3880
rect 9119 3846 9153 3880
rect 9187 3846 9221 3880
rect 9255 3846 9289 3880
rect 9323 3846 9357 3880
rect 9391 3846 9425 3880
rect 9459 3846 9493 3880
rect 9527 3846 9561 3880
rect 9595 3846 9629 3880
rect 9663 3846 9697 3880
rect 9731 3846 9765 3880
rect 9799 3846 9833 3880
rect 9867 3846 9901 3880
rect 9935 3846 9969 3880
rect 10003 3846 10037 3880
rect 10071 3846 10105 3880
rect 10139 3846 10173 3880
rect 10207 3846 10241 3880
rect 10312 3847 10346 3881
rect 10380 3847 10414 3881
rect 10448 3847 10482 3881
rect 10516 3847 10550 3881
rect 10584 3847 10618 3881
rect 10652 3847 10686 3881
rect 10720 3847 10754 3881
rect 10788 3847 10822 3881
rect 10856 3847 10890 3881
rect 10924 3847 10958 3881
rect 10992 3847 11026 3881
rect 11060 3847 11094 3881
rect 11128 3847 11162 3881
rect 11196 3847 11230 3881
rect 11264 3847 11298 3881
rect 11332 3847 11366 3881
rect 11400 3847 11434 3881
rect 11468 3847 11502 3881
rect 11536 3847 11570 3881
rect 8643 3776 8677 3810
rect 8711 3776 8745 3810
rect 8779 3776 8813 3810
rect 8847 3776 8881 3810
rect 8915 3776 8949 3810
rect 8983 3776 9017 3810
rect 9051 3776 9085 3810
rect 9119 3776 9153 3810
rect 9187 3776 9221 3810
rect 9255 3776 9289 3810
rect 9323 3776 9357 3810
rect 9391 3776 9425 3810
rect 9459 3776 9493 3810
rect 9527 3776 9561 3810
rect 9595 3776 9629 3810
rect 9663 3776 9697 3810
rect 9731 3776 9765 3810
rect 9799 3776 9833 3810
rect 9867 3776 9901 3810
rect 9935 3776 9969 3810
rect 10003 3776 10037 3810
rect 10071 3776 10105 3810
rect 10139 3776 10173 3810
rect 10207 3776 10241 3810
rect 10312 3777 10346 3811
rect 10380 3777 10414 3811
rect 10448 3777 10482 3811
rect 10516 3777 10550 3811
rect 10584 3777 10618 3811
rect 10652 3777 10686 3811
rect 10720 3777 10754 3811
rect 10788 3777 10822 3811
rect 10856 3777 10890 3811
rect 10924 3777 10958 3811
rect 10992 3777 11026 3811
rect 11060 3777 11094 3811
rect 11128 3777 11162 3811
rect 11196 3777 11230 3811
rect 11264 3777 11298 3811
rect 11332 3777 11366 3811
rect 11400 3777 11434 3811
rect 11468 3777 11502 3811
rect 11536 3777 11570 3811
rect 8643 3706 8677 3740
rect 8711 3706 8745 3740
rect 8779 3706 8813 3740
rect 8847 3706 8881 3740
rect 8915 3706 8949 3740
rect 8983 3706 9017 3740
rect 9051 3706 9085 3740
rect 9119 3706 9153 3740
rect 9187 3706 9221 3740
rect 9255 3706 9289 3740
rect 9323 3706 9357 3740
rect 9391 3706 9425 3740
rect 9459 3706 9493 3740
rect 9527 3706 9561 3740
rect 9595 3706 9629 3740
rect 9663 3706 9697 3740
rect 9731 3706 9765 3740
rect 9799 3706 9833 3740
rect 9867 3706 9901 3740
rect 9935 3706 9969 3740
rect 10003 3706 10037 3740
rect 10071 3706 10105 3740
rect 10139 3706 10173 3740
rect 10207 3706 10241 3740
rect 10312 3707 10346 3741
rect 10380 3707 10414 3741
rect 10448 3707 10482 3741
rect 10516 3707 10550 3741
rect 10584 3707 10618 3741
rect 10652 3707 10686 3741
rect 10720 3707 10754 3741
rect 10788 3707 10822 3741
rect 10856 3707 10890 3741
rect 10924 3707 10958 3741
rect 10992 3707 11026 3741
rect 11060 3707 11094 3741
rect 11128 3707 11162 3741
rect 11196 3707 11230 3741
rect 11264 3707 11298 3741
rect 11332 3707 11366 3741
rect 11400 3707 11434 3741
rect 11468 3707 11502 3741
rect 11536 3707 11570 3741
rect 8643 3636 8677 3670
rect 8711 3636 8745 3670
rect 8779 3636 8813 3670
rect 8847 3636 8881 3670
rect 8915 3636 8949 3670
rect 8983 3636 9017 3670
rect 9051 3636 9085 3670
rect 9119 3636 9153 3670
rect 9187 3636 9221 3670
rect 9255 3636 9289 3670
rect 9323 3636 9357 3670
rect 9391 3636 9425 3670
rect 9459 3636 9493 3670
rect 9527 3636 9561 3670
rect 9595 3636 9629 3670
rect 9663 3636 9697 3670
rect 9731 3636 9765 3670
rect 9799 3636 9833 3670
rect 9867 3636 9901 3670
rect 9935 3636 9969 3670
rect 10003 3636 10037 3670
rect 10071 3636 10105 3670
rect 10139 3636 10173 3670
rect 10207 3636 10241 3670
rect 10312 3637 10346 3671
rect 10380 3637 10414 3671
rect 10448 3637 10482 3671
rect 10516 3637 10550 3671
rect 10584 3637 10618 3671
rect 10652 3637 10686 3671
rect 10720 3637 10754 3671
rect 10788 3637 10822 3671
rect 10856 3637 10890 3671
rect 10924 3637 10958 3671
rect 10992 3637 11026 3671
rect 11060 3637 11094 3671
rect 11128 3637 11162 3671
rect 11196 3637 11230 3671
rect 11264 3637 11298 3671
rect 11332 3637 11366 3671
rect 11400 3637 11434 3671
rect 11468 3637 11502 3671
rect 11536 3637 11570 3671
rect 8643 3566 8677 3600
rect 8711 3566 8745 3600
rect 8779 3566 8813 3600
rect 8847 3566 8881 3600
rect 8915 3566 8949 3600
rect 8983 3566 9017 3600
rect 9051 3566 9085 3600
rect 9119 3566 9153 3600
rect 9187 3566 9221 3600
rect 9255 3566 9289 3600
rect 9323 3566 9357 3600
rect 9391 3566 9425 3600
rect 9459 3566 9493 3600
rect 9527 3566 9561 3600
rect 9595 3566 9629 3600
rect 9663 3566 9697 3600
rect 9731 3566 9765 3600
rect 9799 3566 9833 3600
rect 9867 3566 9901 3600
rect 9935 3566 9969 3600
rect 10003 3566 10037 3600
rect 10071 3566 10105 3600
rect 10139 3566 10173 3600
rect 10207 3566 10241 3600
rect 10312 3567 10346 3601
rect 10380 3567 10414 3601
rect 10448 3567 10482 3601
rect 10516 3567 10550 3601
rect 10584 3567 10618 3601
rect 10652 3567 10686 3601
rect 10720 3567 10754 3601
rect 10788 3567 10822 3601
rect 10856 3567 10890 3601
rect 10924 3567 10958 3601
rect 10992 3567 11026 3601
rect 11060 3567 11094 3601
rect 11128 3567 11162 3601
rect 11196 3567 11230 3601
rect 11264 3567 11298 3601
rect 11332 3567 11366 3601
rect 11400 3567 11434 3601
rect 11468 3567 11502 3601
rect 11536 3567 11570 3601
rect 8643 3496 8677 3530
rect 8711 3496 8745 3530
rect 8779 3496 8813 3530
rect 8847 3496 8881 3530
rect 8915 3496 8949 3530
rect 8983 3496 9017 3530
rect 9051 3496 9085 3530
rect 9119 3496 9153 3530
rect 9187 3496 9221 3530
rect 9255 3496 9289 3530
rect 9323 3496 9357 3530
rect 9391 3496 9425 3530
rect 9459 3496 9493 3530
rect 9527 3496 9561 3530
rect 9595 3496 9629 3530
rect 9663 3496 9697 3530
rect 9731 3496 9765 3530
rect 9799 3496 9833 3530
rect 9867 3496 9901 3530
rect 9935 3496 9969 3530
rect 10003 3496 10037 3530
rect 10071 3496 10105 3530
rect 10139 3496 10173 3530
rect 10207 3496 10241 3530
rect 10312 3497 10346 3531
rect 10380 3497 10414 3531
rect 10448 3497 10482 3531
rect 10516 3497 10550 3531
rect 10584 3497 10618 3531
rect 10652 3497 10686 3531
rect 10720 3497 10754 3531
rect 10788 3497 10822 3531
rect 10856 3497 10890 3531
rect 10924 3497 10958 3531
rect 10992 3497 11026 3531
rect 11060 3497 11094 3531
rect 11128 3497 11162 3531
rect 11196 3497 11230 3531
rect 11264 3497 11298 3531
rect 11332 3497 11366 3531
rect 11400 3497 11434 3531
rect 11468 3497 11502 3531
rect 11536 3497 11570 3531
rect 8643 3426 8677 3460
rect 8711 3426 8745 3460
rect 8779 3426 8813 3460
rect 8847 3426 8881 3460
rect 8915 3426 8949 3460
rect 8983 3426 9017 3460
rect 9051 3426 9085 3460
rect 9119 3426 9153 3460
rect 9187 3426 9221 3460
rect 9255 3426 9289 3460
rect 9323 3426 9357 3460
rect 9391 3426 9425 3460
rect 9459 3426 9493 3460
rect 9527 3426 9561 3460
rect 9595 3426 9629 3460
rect 9663 3426 9697 3460
rect 9731 3426 9765 3460
rect 9799 3426 9833 3460
rect 9867 3426 9901 3460
rect 9935 3426 9969 3460
rect 10003 3426 10037 3460
rect 10071 3426 10105 3460
rect 10139 3426 10173 3460
rect 10207 3426 10241 3460
rect 10312 3427 10346 3461
rect 10380 3427 10414 3461
rect 10448 3427 10482 3461
rect 10516 3427 10550 3461
rect 10584 3427 10618 3461
rect 10652 3427 10686 3461
rect 10720 3427 10754 3461
rect 10788 3427 10822 3461
rect 10856 3427 10890 3461
rect 10924 3427 10958 3461
rect 10992 3427 11026 3461
rect 11060 3427 11094 3461
rect 11128 3427 11162 3461
rect 11196 3427 11230 3461
rect 11264 3427 11298 3461
rect 11332 3427 11366 3461
rect 11400 3427 11434 3461
rect 11468 3427 11502 3461
rect 11536 3427 11570 3461
rect 8643 3356 8677 3390
rect 8711 3356 8745 3390
rect 8779 3356 8813 3390
rect 8847 3356 8881 3390
rect 8915 3356 8949 3390
rect 8983 3356 9017 3390
rect 9051 3356 9085 3390
rect 9119 3356 9153 3390
rect 9187 3356 9221 3390
rect 9255 3356 9289 3390
rect 9323 3356 9357 3390
rect 9391 3356 9425 3390
rect 9459 3356 9493 3390
rect 9527 3356 9561 3390
rect 9595 3356 9629 3390
rect 9663 3356 9697 3390
rect 9731 3356 9765 3390
rect 9799 3356 9833 3390
rect 9867 3356 9901 3390
rect 9935 3356 9969 3390
rect 10003 3356 10037 3390
rect 10071 3356 10105 3390
rect 10139 3356 10173 3390
rect 10207 3356 10241 3390
rect 10312 3357 10346 3391
rect 10380 3357 10414 3391
rect 10448 3357 10482 3391
rect 10516 3357 10550 3391
rect 10584 3357 10618 3391
rect 10652 3357 10686 3391
rect 10720 3357 10754 3391
rect 10788 3357 10822 3391
rect 10856 3357 10890 3391
rect 10924 3357 10958 3391
rect 10992 3357 11026 3391
rect 11060 3357 11094 3391
rect 11128 3357 11162 3391
rect 11196 3357 11230 3391
rect 11264 3357 11298 3391
rect 11332 3357 11366 3391
rect 11400 3357 11434 3391
rect 11468 3357 11502 3391
rect 11536 3357 11570 3391
rect 8643 3286 8677 3320
rect 8711 3286 8745 3320
rect 8779 3286 8813 3320
rect 8847 3286 8881 3320
rect 8915 3286 8949 3320
rect 8983 3286 9017 3320
rect 9051 3286 9085 3320
rect 9119 3286 9153 3320
rect 9187 3286 9221 3320
rect 9255 3286 9289 3320
rect 9323 3286 9357 3320
rect 9391 3286 9425 3320
rect 9459 3286 9493 3320
rect 9527 3286 9561 3320
rect 9595 3286 9629 3320
rect 9663 3286 9697 3320
rect 9731 3286 9765 3320
rect 9799 3286 9833 3320
rect 9867 3286 9901 3320
rect 9935 3286 9969 3320
rect 10003 3286 10037 3320
rect 10071 3286 10105 3320
rect 10139 3286 10173 3320
rect 10207 3286 10241 3320
rect 10312 3287 10346 3321
rect 10380 3287 10414 3321
rect 10448 3287 10482 3321
rect 10516 3287 10550 3321
rect 10584 3287 10618 3321
rect 10652 3287 10686 3321
rect 10720 3287 10754 3321
rect 10788 3287 10822 3321
rect 10856 3287 10890 3321
rect 10924 3287 10958 3321
rect 10992 3287 11026 3321
rect 11060 3287 11094 3321
rect 11128 3287 11162 3321
rect 11196 3287 11230 3321
rect 11264 3287 11298 3321
rect 11332 3287 11366 3321
rect 11400 3287 11434 3321
rect 11468 3287 11502 3321
rect 11536 3287 11570 3321
rect 1507 3195 1541 3229
rect 1575 3212 1609 3246
rect 1643 3214 1677 3248
rect 1740 3224 1774 3258
rect 1809 3224 1843 3258
rect 1878 3224 1912 3258
rect 1947 3224 1981 3258
rect 2016 3224 2050 3258
rect 2085 3224 2119 3258
rect 2154 3224 2188 3258
rect 2223 3224 2257 3258
rect 2292 3224 2326 3258
rect 2361 3224 2395 3258
rect 2430 3224 2464 3258
rect 2499 3224 2533 3258
rect 2568 3224 2602 3258
rect 2637 3224 2671 3258
rect 2706 3224 2740 3258
rect 2775 3224 2809 3258
rect 1507 3126 1541 3160
rect 1575 3142 1609 3176
rect 1643 3144 1677 3178
rect 1740 3156 1774 3190
rect 1809 3156 1843 3190
rect 1878 3156 1912 3190
rect 1947 3156 1981 3190
rect 2016 3156 2050 3190
rect 2085 3156 2119 3190
rect 2154 3156 2188 3190
rect 2223 3156 2257 3190
rect 2292 3156 2326 3190
rect 2361 3156 2395 3190
rect 2430 3156 2464 3190
rect 2499 3156 2533 3190
rect 2568 3156 2602 3190
rect 2637 3156 2671 3190
rect 2706 3156 2740 3190
rect 2775 3156 2809 3190
rect 1507 3057 1541 3091
rect 1575 3073 1609 3107
rect 1643 3074 1677 3108
rect 1740 3088 1774 3122
rect 1809 3088 1843 3122
rect 1878 3088 1912 3122
rect 1947 3088 1981 3122
rect 2016 3088 2050 3122
rect 2085 3088 2119 3122
rect 2154 3088 2188 3122
rect 2223 3088 2257 3122
rect 2292 3088 2326 3122
rect 2361 3088 2395 3122
rect 2430 3088 2464 3122
rect 2499 3088 2533 3122
rect 2568 3088 2602 3122
rect 2637 3088 2671 3122
rect 2706 3088 2740 3122
rect 2775 3088 2809 3122
rect 2844 3088 4782 3258
rect 8643 3216 8677 3250
rect 8711 3216 8745 3250
rect 8779 3216 8813 3250
rect 8847 3216 8881 3250
rect 8915 3216 8949 3250
rect 8983 3216 9017 3250
rect 9051 3216 9085 3250
rect 9119 3216 9153 3250
rect 9187 3216 9221 3250
rect 9255 3216 9289 3250
rect 9323 3216 9357 3250
rect 9391 3216 9425 3250
rect 9459 3216 9493 3250
rect 9527 3216 9561 3250
rect 9595 3216 9629 3250
rect 9663 3216 9697 3250
rect 9731 3216 9765 3250
rect 9799 3216 9833 3250
rect 9867 3216 9901 3250
rect 9935 3216 9969 3250
rect 10003 3216 10037 3250
rect 10071 3216 10105 3250
rect 10139 3216 10173 3250
rect 10207 3216 10241 3250
rect 10312 3217 10346 3251
rect 10380 3217 10414 3251
rect 10448 3217 10482 3251
rect 10516 3217 10550 3251
rect 10584 3217 10618 3251
rect 10652 3217 10686 3251
rect 10720 3217 10754 3251
rect 10788 3217 10822 3251
rect 10856 3217 10890 3251
rect 10924 3217 10958 3251
rect 10992 3217 11026 3251
rect 11060 3217 11094 3251
rect 11128 3217 11162 3251
rect 11196 3217 11230 3251
rect 11264 3217 11298 3251
rect 11332 3217 11366 3251
rect 11400 3217 11434 3251
rect 11468 3217 11502 3251
rect 11536 3217 11570 3251
rect 8643 3146 8677 3180
rect 8711 3146 8745 3180
rect 8779 3146 8813 3180
rect 8847 3146 8881 3180
rect 8915 3146 8949 3180
rect 8983 3146 9017 3180
rect 9051 3146 9085 3180
rect 9119 3146 9153 3180
rect 9187 3146 9221 3180
rect 9255 3146 9289 3180
rect 9323 3146 9357 3180
rect 9391 3146 9425 3180
rect 9459 3146 9493 3180
rect 9527 3146 9561 3180
rect 9595 3146 9629 3180
rect 9663 3146 9697 3180
rect 9731 3146 9765 3180
rect 9799 3146 9833 3180
rect 9867 3146 9901 3180
rect 9935 3146 9969 3180
rect 10003 3146 10037 3180
rect 10071 3146 10105 3180
rect 10139 3146 10173 3180
rect 10207 3146 10241 3180
rect 10312 3147 10346 3181
rect 10380 3147 10414 3181
rect 10448 3147 10482 3181
rect 10516 3147 10550 3181
rect 10584 3147 10618 3181
rect 10652 3147 10686 3181
rect 10720 3147 10754 3181
rect 10788 3147 10822 3181
rect 10856 3147 10890 3181
rect 10924 3147 10958 3181
rect 10992 3147 11026 3181
rect 11060 3147 11094 3181
rect 11128 3147 11162 3181
rect 11196 3147 11230 3181
rect 11264 3147 11298 3181
rect 11332 3147 11366 3181
rect 11400 3147 11434 3181
rect 11468 3147 11502 3181
rect 11536 3147 11570 3181
rect 1507 2988 1541 3022
rect 1575 3004 1609 3038
rect 1643 3004 1677 3038
rect 1507 2919 1541 2953
rect 1575 2935 1609 2969
rect 1643 2935 1677 2969
rect 1507 2850 1541 2884
rect 1575 2866 1609 2900
rect 1643 2866 1677 2900
rect 1507 2781 1541 2815
rect 1575 2797 1609 2831
rect 1643 2797 1677 2831
rect 1507 2712 1541 2746
rect 1575 2728 1609 2762
rect 1643 2728 1677 2762
rect 1507 2643 1541 2677
rect 1575 2659 1609 2693
rect 1643 2659 1677 2693
rect 1507 2575 1541 2609
rect 1575 2590 1609 2624
rect 1643 2590 1677 2624
rect 1507 2507 1541 2541
rect 1575 2521 1609 2555
rect 1643 2521 1677 2555
rect 1507 2439 1541 2473
rect 1575 2452 1609 2486
rect 1643 2452 1677 2486
rect 1507 2371 1541 2405
rect 1575 2383 1609 2417
rect 1643 2383 1677 2417
rect 8643 3076 8677 3110
rect 8711 3076 8745 3110
rect 8779 3076 8813 3110
rect 8847 3076 8881 3110
rect 8915 3076 8949 3110
rect 8983 3076 9017 3110
rect 9051 3076 9085 3110
rect 9119 3076 9153 3110
rect 9187 3076 9221 3110
rect 9255 3076 9289 3110
rect 9323 3076 9357 3110
rect 9391 3076 9425 3110
rect 9459 3076 9493 3110
rect 9527 3076 9561 3110
rect 9595 3076 9629 3110
rect 9663 3076 9697 3110
rect 9731 3076 9765 3110
rect 9799 3076 9833 3110
rect 9867 3076 9901 3110
rect 9935 3076 9969 3110
rect 10003 3076 10037 3110
rect 10071 3076 10105 3110
rect 10139 3076 10173 3110
rect 10207 3076 10241 3110
rect 10312 3077 10346 3111
rect 10380 3077 10414 3111
rect 10448 3077 10482 3111
rect 10516 3077 10550 3111
rect 10584 3077 10618 3111
rect 10652 3077 10686 3111
rect 10720 3077 10754 3111
rect 10788 3077 10822 3111
rect 10856 3077 10890 3111
rect 10924 3077 10958 3111
rect 10992 3077 11026 3111
rect 11060 3077 11094 3111
rect 11128 3077 11162 3111
rect 11196 3077 11230 3111
rect 11264 3077 11298 3111
rect 11332 3077 11366 3111
rect 11400 3077 11434 3111
rect 11468 3077 11502 3111
rect 11536 3077 11570 3111
rect 8643 3006 8677 3040
rect 8711 3006 8745 3040
rect 8779 3006 8813 3040
rect 8847 3006 8881 3040
rect 8915 3006 8949 3040
rect 8983 3006 9017 3040
rect 9051 3006 9085 3040
rect 9119 3006 9153 3040
rect 9187 3006 9221 3040
rect 9255 3006 9289 3040
rect 9323 3006 9357 3040
rect 9391 3006 9425 3040
rect 9459 3006 9493 3040
rect 9527 3006 9561 3040
rect 9595 3006 9629 3040
rect 9663 3006 9697 3040
rect 9731 3006 9765 3040
rect 9799 3006 9833 3040
rect 9867 3006 9901 3040
rect 9935 3006 9969 3040
rect 10003 3006 10037 3040
rect 10071 3006 10105 3040
rect 10139 3006 10173 3040
rect 10207 3006 10241 3040
rect 10312 3007 10346 3041
rect 10380 3007 10414 3041
rect 10448 3007 10482 3041
rect 10516 3007 10550 3041
rect 10584 3007 10618 3041
rect 10652 3007 10686 3041
rect 10720 3007 10754 3041
rect 10788 3007 10822 3041
rect 10856 3007 10890 3041
rect 10924 3007 10958 3041
rect 10992 3007 11026 3041
rect 11060 3007 11094 3041
rect 11128 3007 11162 3041
rect 11196 3007 11230 3041
rect 11264 3007 11298 3041
rect 11332 3007 11366 3041
rect 11400 3007 11434 3041
rect 11468 3007 11502 3041
rect 11536 3007 11570 3041
rect 8643 2936 8677 2970
rect 8711 2936 8745 2970
rect 8779 2936 8813 2970
rect 8847 2936 8881 2970
rect 8915 2936 8949 2970
rect 8983 2936 9017 2970
rect 9051 2936 9085 2970
rect 9119 2936 9153 2970
rect 9187 2936 9221 2970
rect 9255 2936 9289 2970
rect 9323 2936 9357 2970
rect 9391 2936 9425 2970
rect 9459 2936 9493 2970
rect 9527 2936 9561 2970
rect 9595 2936 9629 2970
rect 9663 2936 9697 2970
rect 9731 2936 9765 2970
rect 9799 2936 9833 2970
rect 9867 2936 9901 2970
rect 9935 2936 9969 2970
rect 10003 2936 10037 2970
rect 10071 2936 10105 2970
rect 10139 2936 10173 2970
rect 10207 2936 10241 2970
rect 10312 2937 10346 2971
rect 10380 2937 10414 2971
rect 10448 2937 10482 2971
rect 10516 2937 10550 2971
rect 10584 2937 10618 2971
rect 10652 2937 10686 2971
rect 10720 2937 10754 2971
rect 10788 2937 10822 2971
rect 10856 2937 10890 2971
rect 10924 2937 10958 2971
rect 10992 2937 11026 2971
rect 11060 2937 11094 2971
rect 11128 2937 11162 2971
rect 11196 2937 11230 2971
rect 11264 2937 11298 2971
rect 11332 2937 11366 2971
rect 11400 2937 11434 2971
rect 11468 2937 11502 2971
rect 11536 2937 11570 2971
rect 8643 2866 8677 2900
rect 8711 2866 8745 2900
rect 8779 2866 8813 2900
rect 8847 2866 8881 2900
rect 8915 2866 8949 2900
rect 8983 2866 9017 2900
rect 9051 2866 9085 2900
rect 9119 2866 9153 2900
rect 9187 2866 9221 2900
rect 9255 2866 9289 2900
rect 9323 2866 9357 2900
rect 9391 2866 9425 2900
rect 9459 2866 9493 2900
rect 9527 2866 9561 2900
rect 9595 2866 9629 2900
rect 9663 2866 9697 2900
rect 9731 2866 9765 2900
rect 9799 2866 9833 2900
rect 9867 2866 9901 2900
rect 9935 2866 9969 2900
rect 10003 2866 10037 2900
rect 10071 2866 10105 2900
rect 10139 2866 10173 2900
rect 10207 2866 10241 2900
rect 10312 2867 10346 2901
rect 10380 2867 10414 2901
rect 10448 2867 10482 2901
rect 10516 2867 10550 2901
rect 10584 2867 10618 2901
rect 10652 2867 10686 2901
rect 10720 2867 10754 2901
rect 10788 2867 10822 2901
rect 10856 2867 10890 2901
rect 10924 2867 10958 2901
rect 10992 2867 11026 2901
rect 11060 2867 11094 2901
rect 11128 2867 11162 2901
rect 11196 2867 11230 2901
rect 11264 2867 11298 2901
rect 11332 2867 11366 2901
rect 11400 2867 11434 2901
rect 11468 2867 11502 2901
rect 11536 2867 11570 2901
rect 8643 2796 8677 2830
rect 8711 2796 8745 2830
rect 8779 2796 8813 2830
rect 8847 2796 8881 2830
rect 8915 2796 8949 2830
rect 8983 2796 9017 2830
rect 9051 2796 9085 2830
rect 9119 2796 9153 2830
rect 9187 2796 9221 2830
rect 9255 2796 9289 2830
rect 9323 2796 9357 2830
rect 9391 2796 9425 2830
rect 9459 2796 9493 2830
rect 9527 2796 9561 2830
rect 9595 2796 9629 2830
rect 9663 2796 9697 2830
rect 9731 2796 9765 2830
rect 9799 2796 9833 2830
rect 9867 2796 9901 2830
rect 9935 2796 9969 2830
rect 10003 2796 10037 2830
rect 10071 2796 10105 2830
rect 10139 2796 10173 2830
rect 10207 2796 10241 2830
rect 10312 2797 10346 2831
rect 10380 2797 10414 2831
rect 10448 2797 10482 2831
rect 10516 2797 10550 2831
rect 10584 2797 10618 2831
rect 10652 2797 10686 2831
rect 10720 2797 10754 2831
rect 10788 2797 10822 2831
rect 10856 2797 10890 2831
rect 10924 2797 10958 2831
rect 10992 2797 11026 2831
rect 11060 2797 11094 2831
rect 11128 2797 11162 2831
rect 11196 2797 11230 2831
rect 11264 2797 11298 2831
rect 11332 2797 11366 2831
rect 11400 2797 11434 2831
rect 11468 2797 11502 2831
rect 11536 2797 11570 2831
rect 8643 2727 8677 2761
rect 8711 2727 8745 2761
rect 8779 2727 8813 2761
rect 8847 2727 8881 2761
rect 8915 2727 8949 2761
rect 8983 2727 9017 2761
rect 9051 2727 9085 2761
rect 9119 2727 9153 2761
rect 9187 2727 9221 2761
rect 9255 2727 9289 2761
rect 9323 2727 9357 2761
rect 9391 2727 9425 2761
rect 9459 2727 9493 2761
rect 9527 2727 9561 2761
rect 9595 2727 9629 2761
rect 9663 2727 9697 2761
rect 9731 2727 9765 2761
rect 9799 2727 9833 2761
rect 9867 2727 9901 2761
rect 9935 2727 9969 2761
rect 10003 2727 10037 2761
rect 10071 2727 10105 2761
rect 10139 2727 10173 2761
rect 10207 2727 10241 2761
rect 10312 2727 10346 2761
rect 10380 2727 10414 2761
rect 10448 2727 10482 2761
rect 10516 2727 10550 2761
rect 10584 2727 10618 2761
rect 10652 2727 10686 2761
rect 10720 2727 10754 2761
rect 10788 2727 10822 2761
rect 10856 2727 10890 2761
rect 10924 2727 10958 2761
rect 10992 2727 11026 2761
rect 11060 2727 11094 2761
rect 11128 2727 11162 2761
rect 11196 2727 11230 2761
rect 11264 2727 11298 2761
rect 11332 2727 11366 2761
rect 11400 2727 11434 2761
rect 11468 2727 11502 2761
rect 11536 2727 11570 2761
rect 12595 4329 12629 4363
rect 12663 4329 12697 4363
rect 12731 4329 12765 4363
rect 12799 4329 12833 4363
rect 12867 4329 12901 4363
rect 12935 4329 12969 4363
rect 13003 4329 13037 4363
rect 13071 4329 13105 4363
rect 13139 4329 13173 4363
rect 13207 4329 13241 4363
rect 13275 4329 13309 4363
rect 13343 4329 13377 4363
rect 12595 4259 12629 4293
rect 12663 4259 12697 4293
rect 12731 4259 12765 4293
rect 12799 4259 12833 4293
rect 12867 4259 12901 4293
rect 12935 4259 12969 4293
rect 13003 4259 13037 4293
rect 13071 4259 13105 4293
rect 13139 4259 13173 4293
rect 13207 4259 13241 4293
rect 13275 4259 13309 4293
rect 13343 4259 13377 4293
rect 12595 4189 12629 4223
rect 12663 4189 12697 4223
rect 12731 4189 12765 4223
rect 12799 4189 12833 4223
rect 12867 4189 12901 4223
rect 12935 4189 12969 4223
rect 13003 4189 13037 4223
rect 13071 4189 13105 4223
rect 13139 4189 13173 4223
rect 13207 4189 13241 4223
rect 13275 4189 13309 4223
rect 13343 4189 13377 4223
rect 12595 4119 12629 4153
rect 12663 4119 12697 4153
rect 12731 4119 12765 4153
rect 12799 4119 12833 4153
rect 12867 4119 12901 4153
rect 12935 4119 12969 4153
rect 13003 4119 13037 4153
rect 13071 4119 13105 4153
rect 13139 4119 13173 4153
rect 13207 4119 13241 4153
rect 13275 4119 13309 4153
rect 13343 4119 13377 4153
rect 12595 4049 12629 4083
rect 12663 4049 12697 4083
rect 12731 4049 12765 4083
rect 12799 4049 12833 4083
rect 12867 4049 12901 4083
rect 12935 4049 12969 4083
rect 13003 4049 13037 4083
rect 13071 4049 13105 4083
rect 13139 4049 13173 4083
rect 13207 4049 13241 4083
rect 13275 4049 13309 4083
rect 13343 4049 13377 4083
rect 12595 3979 12629 4013
rect 12663 3979 12697 4013
rect 12731 3979 12765 4013
rect 12799 3979 12833 4013
rect 12867 3979 12901 4013
rect 12935 3979 12969 4013
rect 13003 3979 13037 4013
rect 13071 3979 13105 4013
rect 13139 3979 13173 4013
rect 13207 3979 13241 4013
rect 13275 3979 13309 4013
rect 13343 3979 13377 4013
rect 12595 3909 12629 3943
rect 12663 3909 12697 3943
rect 12731 3909 12765 3943
rect 12799 3909 12833 3943
rect 12867 3909 12901 3943
rect 12935 3909 12969 3943
rect 13003 3909 13037 3943
rect 13071 3909 13105 3943
rect 13139 3909 13173 3943
rect 13207 3909 13241 3943
rect 13275 3909 13309 3943
rect 13343 3909 13377 3943
rect 12595 3839 12629 3873
rect 12663 3839 12697 3873
rect 12731 3839 12765 3873
rect 12799 3839 12833 3873
rect 12867 3839 12901 3873
rect 12935 3839 12969 3873
rect 13003 3839 13037 3873
rect 13071 3839 13105 3873
rect 13139 3839 13173 3873
rect 13207 3839 13241 3873
rect 13275 3839 13309 3873
rect 13343 3839 13377 3873
rect 12595 3769 12629 3803
rect 12663 3769 12697 3803
rect 12731 3769 12765 3803
rect 12799 3769 12833 3803
rect 12867 3769 12901 3803
rect 12935 3769 12969 3803
rect 13003 3769 13037 3803
rect 13071 3769 13105 3803
rect 13139 3769 13173 3803
rect 13207 3769 13241 3803
rect 13275 3769 13309 3803
rect 13343 3769 13377 3803
rect 12595 3699 12629 3733
rect 12663 3699 12697 3733
rect 12731 3699 12765 3733
rect 12799 3699 12833 3733
rect 12867 3699 12901 3733
rect 12935 3699 12969 3733
rect 13003 3699 13037 3733
rect 13071 3699 13105 3733
rect 13139 3699 13173 3733
rect 13207 3699 13241 3733
rect 13275 3699 13309 3733
rect 13343 3699 13377 3733
rect 12595 3629 12629 3663
rect 12663 3629 12697 3663
rect 12731 3629 12765 3663
rect 12799 3629 12833 3663
rect 12867 3629 12901 3663
rect 12935 3629 12969 3663
rect 13003 3629 13037 3663
rect 13071 3629 13105 3663
rect 13139 3629 13173 3663
rect 13207 3629 13241 3663
rect 13275 3629 13309 3663
rect 13343 3629 13377 3663
rect 12595 3559 12629 3593
rect 12663 3559 12697 3593
rect 12731 3559 12765 3593
rect 12799 3559 12833 3593
rect 12867 3559 12901 3593
rect 12935 3559 12969 3593
rect 13003 3559 13037 3593
rect 13071 3559 13105 3593
rect 13139 3559 13173 3593
rect 13207 3559 13241 3593
rect 13275 3559 13309 3593
rect 13343 3559 13377 3593
rect 12595 3489 12629 3523
rect 12663 3489 12697 3523
rect 12731 3489 12765 3523
rect 12799 3489 12833 3523
rect 12867 3489 12901 3523
rect 12935 3489 12969 3523
rect 13003 3489 13037 3523
rect 13071 3489 13105 3523
rect 13139 3489 13173 3523
rect 13207 3489 13241 3523
rect 13275 3489 13309 3523
rect 13343 3489 13377 3523
rect 12595 3419 12629 3453
rect 12663 3419 12697 3453
rect 12731 3419 12765 3453
rect 12799 3419 12833 3453
rect 12867 3419 12901 3453
rect 12935 3419 12969 3453
rect 13003 3419 13037 3453
rect 13071 3419 13105 3453
rect 13139 3419 13173 3453
rect 13207 3419 13241 3453
rect 13275 3419 13309 3453
rect 13343 3419 13377 3453
rect 12595 3349 12629 3383
rect 12663 3349 12697 3383
rect 12731 3349 12765 3383
rect 12799 3349 12833 3383
rect 12867 3349 12901 3383
rect 12935 3349 12969 3383
rect 13003 3349 13037 3383
rect 13071 3349 13105 3383
rect 13139 3349 13173 3383
rect 13207 3349 13241 3383
rect 13275 3349 13309 3383
rect 13343 3349 13377 3383
rect 12595 3279 12629 3313
rect 12663 3279 12697 3313
rect 12731 3279 12765 3313
rect 12799 3279 12833 3313
rect 12867 3279 12901 3313
rect 12935 3279 12969 3313
rect 13003 3279 13037 3313
rect 13071 3279 13105 3313
rect 13139 3279 13173 3313
rect 13207 3279 13241 3313
rect 13275 3279 13309 3313
rect 13343 3279 13377 3313
rect 12595 3209 12629 3243
rect 12663 3209 12697 3243
rect 12731 3209 12765 3243
rect 12799 3209 12833 3243
rect 12867 3209 12901 3243
rect 12935 3209 12969 3243
rect 13003 3209 13037 3243
rect 13071 3209 13105 3243
rect 13139 3209 13173 3243
rect 13207 3209 13241 3243
rect 13275 3209 13309 3243
rect 13343 3209 13377 3243
rect 12595 3139 12629 3173
rect 12663 3139 12697 3173
rect 12731 3139 12765 3173
rect 12799 3139 12833 3173
rect 12867 3139 12901 3173
rect 12935 3139 12969 3173
rect 13003 3139 13037 3173
rect 13071 3139 13105 3173
rect 13139 3139 13173 3173
rect 13207 3139 13241 3173
rect 13275 3139 13309 3173
rect 13343 3139 13377 3173
rect 12595 3069 12629 3103
rect 12663 3069 12697 3103
rect 12731 3069 12765 3103
rect 12799 3069 12833 3103
rect 12867 3069 12901 3103
rect 12935 3069 12969 3103
rect 13003 3069 13037 3103
rect 13071 3069 13105 3103
rect 13139 3069 13173 3103
rect 13207 3069 13241 3103
rect 13275 3069 13309 3103
rect 13343 3069 13377 3103
rect 12595 2999 12629 3033
rect 12663 2999 12697 3033
rect 12731 2999 12765 3033
rect 12799 2999 12833 3033
rect 12867 2999 12901 3033
rect 12935 2999 12969 3033
rect 13003 2999 13037 3033
rect 13071 2999 13105 3033
rect 13139 2999 13173 3033
rect 13207 2999 13241 3033
rect 13275 2999 13309 3033
rect 13343 2999 13377 3033
rect 12595 2930 12629 2964
rect 12663 2930 12697 2964
rect 12731 2930 12765 2964
rect 12799 2930 12833 2964
rect 12867 2930 12901 2964
rect 12935 2930 12969 2964
rect 13003 2930 13037 2964
rect 13071 2930 13105 2964
rect 13139 2930 13173 2964
rect 13207 2930 13241 2964
rect 13275 2930 13309 2964
rect 13343 2930 13377 2964
rect 12595 2861 12629 2895
rect 12663 2861 12697 2895
rect 12731 2861 12765 2895
rect 12799 2861 12833 2895
rect 12867 2861 12901 2895
rect 12935 2861 12969 2895
rect 13003 2861 13037 2895
rect 13071 2861 13105 2895
rect 13139 2861 13173 2895
rect 13207 2861 13241 2895
rect 13275 2861 13309 2895
rect 13343 2861 13377 2895
rect 12595 2792 12629 2826
rect 12663 2792 12697 2826
rect 12731 2792 12765 2826
rect 12799 2792 12833 2826
rect 12867 2792 12901 2826
rect 12935 2792 12969 2826
rect 13003 2792 13037 2826
rect 13071 2792 13105 2826
rect 13139 2792 13173 2826
rect 13207 2792 13241 2826
rect 13275 2792 13309 2826
rect 13343 2792 13377 2826
rect 12595 2723 13377 2757
rect 8643 2658 8677 2692
rect 8711 2658 8745 2692
rect 8779 2658 8813 2692
rect 8847 2658 8881 2692
rect 8915 2658 8949 2692
rect 8983 2658 9017 2692
rect 9051 2658 9085 2692
rect 9119 2658 9153 2692
rect 9187 2658 9221 2692
rect 9255 2658 9289 2692
rect 9323 2658 9357 2692
rect 9391 2658 9425 2692
rect 9459 2658 9493 2692
rect 9527 2658 9561 2692
rect 9595 2658 9629 2692
rect 9663 2658 9697 2692
rect 9731 2658 9765 2692
rect 9799 2658 9833 2692
rect 9867 2658 9901 2692
rect 9935 2658 9969 2692
rect 10003 2658 10037 2692
rect 10071 2658 10105 2692
rect 10139 2658 10173 2692
rect 10207 2658 10241 2692
rect 10312 2658 10346 2692
rect 10380 2658 10414 2692
rect 10448 2658 10482 2692
rect 10516 2658 10550 2692
rect 10584 2658 10618 2692
rect 10652 2658 10686 2692
rect 10720 2658 10754 2692
rect 10788 2658 10822 2692
rect 10856 2658 10890 2692
rect 10924 2658 10958 2692
rect 10992 2658 11026 2692
rect 11060 2658 11094 2692
rect 11128 2658 11162 2692
rect 11196 2658 11230 2692
rect 11264 2658 11298 2692
rect 11332 2658 11366 2692
rect 11400 2658 11434 2692
rect 11468 2658 11502 2692
rect 11536 2658 11570 2692
rect 11652 2665 11686 2699
rect 11720 2665 11754 2699
rect 11788 2665 11822 2699
rect 11856 2665 11890 2699
rect 11924 2665 11958 2699
rect 11992 2665 12026 2699
rect 12060 2665 12094 2699
rect 12128 2665 12162 2699
rect 12196 2665 12230 2699
rect 12264 2665 12298 2699
rect 12332 2665 12366 2699
rect 12400 2665 12434 2699
rect 12468 2665 12502 2699
rect 12595 2689 13355 2723
rect 12573 2655 13355 2689
rect 8643 2589 8677 2623
rect 8711 2589 8745 2623
rect 8779 2589 8813 2623
rect 8847 2589 8881 2623
rect 8915 2589 8949 2623
rect 8983 2589 9017 2623
rect 9051 2589 9085 2623
rect 9119 2589 9153 2623
rect 9187 2589 9221 2623
rect 9255 2589 9289 2623
rect 9323 2589 9357 2623
rect 9391 2589 9425 2623
rect 9459 2589 9493 2623
rect 9527 2589 9561 2623
rect 9595 2589 9629 2623
rect 9663 2589 9697 2623
rect 9731 2589 9765 2623
rect 9799 2589 9833 2623
rect 9867 2589 9901 2623
rect 9935 2589 9969 2623
rect 10003 2589 10037 2623
rect 10071 2589 10105 2623
rect 10139 2589 10173 2623
rect 10207 2589 10241 2623
rect 10312 2589 10346 2623
rect 10380 2589 10414 2623
rect 10448 2589 10482 2623
rect 10516 2589 10550 2623
rect 10584 2589 10618 2623
rect 10652 2589 10686 2623
rect 10720 2589 10754 2623
rect 10788 2589 10822 2623
rect 10856 2589 10890 2623
rect 10924 2589 10958 2623
rect 10992 2589 11026 2623
rect 11060 2589 11094 2623
rect 11128 2589 11162 2623
rect 11196 2589 11230 2623
rect 11264 2589 11298 2623
rect 11332 2589 11366 2623
rect 11400 2589 11434 2623
rect 11468 2589 11502 2623
rect 11536 2589 11570 2623
rect 11652 2595 11686 2629
rect 11720 2595 11754 2629
rect 11788 2595 11822 2629
rect 11856 2595 11890 2629
rect 11924 2595 11958 2629
rect 11992 2595 12026 2629
rect 12060 2595 12094 2629
rect 12128 2595 12162 2629
rect 12196 2595 12230 2629
rect 12264 2595 12298 2629
rect 12332 2595 12366 2629
rect 12400 2595 12434 2629
rect 12468 2595 12502 2629
rect 12573 2586 12607 2620
rect 12641 2586 12675 2620
rect 12709 2586 12743 2620
rect 12777 2586 12811 2620
rect 12845 2586 12879 2620
rect 12913 2586 12947 2620
rect 12981 2586 13015 2620
rect 13049 2586 13083 2620
rect 13117 2586 13151 2620
rect 13185 2586 13219 2620
rect 13253 2586 13287 2620
rect 13321 2586 13355 2620
rect 8643 2520 8677 2554
rect 8711 2520 8745 2554
rect 8779 2520 8813 2554
rect 8847 2520 8881 2554
rect 8915 2520 8949 2554
rect 8983 2520 9017 2554
rect 9051 2520 9085 2554
rect 9119 2520 9153 2554
rect 9187 2520 9221 2554
rect 9255 2520 9289 2554
rect 9323 2520 9357 2554
rect 9391 2520 9425 2554
rect 9459 2520 9493 2554
rect 9527 2520 9561 2554
rect 9595 2520 9629 2554
rect 9663 2520 9697 2554
rect 9731 2520 9765 2554
rect 9799 2520 9833 2554
rect 9867 2520 9901 2554
rect 9935 2520 9969 2554
rect 10003 2520 10037 2554
rect 10071 2520 10105 2554
rect 10139 2520 10173 2554
rect 10207 2520 10241 2554
rect 10312 2520 10346 2554
rect 10380 2520 10414 2554
rect 10448 2520 10482 2554
rect 10516 2520 10550 2554
rect 10584 2520 10618 2554
rect 10652 2520 10686 2554
rect 10720 2520 10754 2554
rect 10788 2520 10822 2554
rect 10856 2520 10890 2554
rect 10924 2520 10958 2554
rect 10992 2520 11026 2554
rect 11060 2520 11094 2554
rect 11128 2520 11162 2554
rect 11196 2520 11230 2554
rect 11264 2520 11298 2554
rect 11332 2520 11366 2554
rect 11400 2520 11434 2554
rect 11468 2520 11502 2554
rect 11536 2520 11570 2554
rect 11652 2525 11686 2559
rect 11720 2525 11754 2559
rect 11788 2525 11822 2559
rect 11856 2525 11890 2559
rect 11924 2525 11958 2559
rect 11992 2525 12026 2559
rect 12060 2525 12094 2559
rect 12128 2525 12162 2559
rect 12196 2525 12230 2559
rect 12264 2525 12298 2559
rect 12332 2525 12366 2559
rect 12400 2525 12434 2559
rect 12468 2525 12502 2559
rect 12573 2517 12607 2551
rect 12641 2517 12675 2551
rect 12709 2517 12743 2551
rect 12777 2517 12811 2551
rect 12845 2517 12879 2551
rect 12913 2517 12947 2551
rect 12981 2517 13015 2551
rect 13049 2517 13083 2551
rect 13117 2517 13151 2551
rect 13185 2517 13219 2551
rect 13253 2517 13287 2551
rect 13321 2517 13355 2551
rect 8643 2451 8677 2485
rect 8711 2451 8745 2485
rect 8779 2451 8813 2485
rect 8847 2451 8881 2485
rect 8915 2451 8949 2485
rect 8983 2451 9017 2485
rect 9051 2451 9085 2485
rect 9119 2451 9153 2485
rect 9187 2451 9221 2485
rect 9255 2451 9289 2485
rect 9323 2451 9357 2485
rect 9391 2451 9425 2485
rect 9459 2451 9493 2485
rect 9527 2451 9561 2485
rect 9595 2451 9629 2485
rect 9663 2451 9697 2485
rect 9731 2451 9765 2485
rect 9799 2451 9833 2485
rect 9867 2451 9901 2485
rect 9935 2451 9969 2485
rect 10003 2451 10037 2485
rect 10071 2451 10105 2485
rect 10139 2451 10173 2485
rect 10207 2451 10241 2485
rect 10312 2451 10346 2485
rect 10380 2451 10414 2485
rect 10448 2451 10482 2485
rect 10516 2451 10550 2485
rect 10584 2451 10618 2485
rect 10652 2451 10686 2485
rect 10720 2451 10754 2485
rect 10788 2451 10822 2485
rect 10856 2451 10890 2485
rect 10924 2451 10958 2485
rect 10992 2451 11026 2485
rect 11060 2451 11094 2485
rect 11128 2451 11162 2485
rect 11196 2451 11230 2485
rect 11264 2451 11298 2485
rect 11332 2451 11366 2485
rect 11400 2451 11434 2485
rect 11468 2451 11502 2485
rect 11536 2451 11570 2485
rect 11652 2455 11686 2489
rect 11720 2455 11754 2489
rect 11788 2455 11822 2489
rect 11856 2455 11890 2489
rect 11924 2455 11958 2489
rect 11992 2455 12026 2489
rect 12060 2455 12094 2489
rect 12128 2455 12162 2489
rect 12196 2455 12230 2489
rect 12264 2455 12298 2489
rect 12332 2455 12366 2489
rect 12400 2455 12434 2489
rect 12468 2455 12502 2489
rect 12573 2448 12607 2482
rect 12641 2448 12675 2482
rect 12709 2448 12743 2482
rect 12777 2448 12811 2482
rect 12845 2448 12879 2482
rect 12913 2448 12947 2482
rect 12981 2448 13015 2482
rect 13049 2448 13083 2482
rect 13117 2448 13151 2482
rect 13185 2448 13219 2482
rect 13253 2448 13287 2482
rect 13321 2448 13355 2482
rect 8643 2382 8677 2416
rect 8711 2382 8745 2416
rect 8779 2382 8813 2416
rect 8847 2382 8881 2416
rect 8915 2382 8949 2416
rect 8983 2382 9017 2416
rect 9051 2382 9085 2416
rect 9119 2382 9153 2416
rect 9187 2382 9221 2416
rect 9255 2382 9289 2416
rect 9323 2382 9357 2416
rect 9391 2382 9425 2416
rect 9459 2382 9493 2416
rect 9527 2382 9561 2416
rect 9595 2382 9629 2416
rect 9663 2382 9697 2416
rect 9731 2382 9765 2416
rect 9799 2382 9833 2416
rect 9867 2382 9901 2416
rect 9935 2382 9969 2416
rect 10003 2382 10037 2416
rect 10071 2382 10105 2416
rect 10139 2382 10173 2416
rect 10207 2382 10241 2416
rect 10312 2382 10346 2416
rect 10380 2382 10414 2416
rect 10448 2382 10482 2416
rect 10516 2382 10550 2416
rect 10584 2382 10618 2416
rect 10652 2382 10686 2416
rect 10720 2382 10754 2416
rect 10788 2382 10822 2416
rect 10856 2382 10890 2416
rect 10924 2382 10958 2416
rect 10992 2382 11026 2416
rect 11060 2382 11094 2416
rect 11128 2382 11162 2416
rect 11196 2382 11230 2416
rect 11264 2382 11298 2416
rect 11332 2382 11366 2416
rect 11400 2382 11434 2416
rect 11468 2382 11502 2416
rect 11536 2382 11570 2416
rect 11652 2385 11686 2419
rect 11720 2385 11754 2419
rect 11788 2385 11822 2419
rect 11856 2385 11890 2419
rect 11924 2385 11958 2419
rect 11992 2385 12026 2419
rect 12060 2385 12094 2419
rect 12128 2385 12162 2419
rect 12196 2385 12230 2419
rect 12264 2385 12298 2419
rect 12332 2385 12366 2419
rect 12400 2385 12434 2419
rect 12468 2385 12502 2419
rect 12573 2379 12607 2413
rect 12641 2379 12675 2413
rect 12709 2379 12743 2413
rect 12777 2379 12811 2413
rect 12845 2379 12879 2413
rect 12913 2379 12947 2413
rect 12981 2379 13015 2413
rect 13049 2379 13083 2413
rect 13117 2379 13151 2413
rect 13185 2379 13219 2413
rect 13253 2379 13287 2413
rect 13321 2379 13355 2413
rect 1507 2303 1541 2337
rect 1575 2314 1609 2348
rect 1643 2314 1677 2348
rect 1740 2327 1774 2361
rect 1809 2327 1843 2361
rect 1878 2327 1912 2361
rect 1947 2327 1981 2361
rect 2016 2327 2050 2361
rect 2085 2327 2119 2361
rect 2154 2327 2188 2361
rect 2223 2327 2257 2361
rect 2292 2327 2326 2361
rect 2361 2327 2395 2361
rect 2430 2327 2464 2361
rect 2499 2327 2533 2361
rect 2568 2327 2602 2361
rect 2637 2327 2671 2361
rect 2706 2327 2740 2361
rect 2775 2327 2809 2361
rect 1507 2235 1541 2269
rect 1575 2245 1609 2279
rect 1643 2245 1677 2279
rect 1740 2259 1774 2293
rect 1809 2259 1843 2293
rect 1878 2259 1912 2293
rect 1947 2259 1981 2293
rect 2016 2259 2050 2293
rect 2085 2259 2119 2293
rect 2154 2259 2188 2293
rect 2223 2259 2257 2293
rect 2292 2259 2326 2293
rect 2361 2259 2395 2293
rect 2430 2259 2464 2293
rect 2499 2259 2533 2293
rect 2568 2259 2602 2293
rect 2637 2259 2671 2293
rect 2706 2259 2740 2293
rect 2775 2259 2809 2293
rect 1507 2167 1541 2201
rect 1575 2176 1609 2210
rect 1643 2176 1677 2210
rect 1740 2191 1774 2225
rect 1809 2191 1843 2225
rect 1878 2191 1912 2225
rect 1947 2191 1981 2225
rect 2016 2191 2050 2225
rect 2085 2191 2119 2225
rect 2154 2191 2188 2225
rect 2223 2191 2257 2225
rect 2292 2191 2326 2225
rect 2361 2191 2395 2225
rect 2430 2191 2464 2225
rect 2499 2191 2533 2225
rect 2568 2191 2602 2225
rect 2637 2191 2671 2225
rect 2706 2191 2740 2225
rect 2775 2191 2809 2225
rect 2844 2191 4782 2361
rect 8643 2313 8677 2347
rect 8711 2313 8745 2347
rect 8779 2313 8813 2347
rect 8847 2313 8881 2347
rect 8915 2313 8949 2347
rect 8983 2313 9017 2347
rect 9051 2313 9085 2347
rect 9119 2313 9153 2347
rect 9187 2313 9221 2347
rect 9255 2313 9289 2347
rect 9323 2313 9357 2347
rect 9391 2313 9425 2347
rect 9459 2313 9493 2347
rect 9527 2313 9561 2347
rect 9595 2313 9629 2347
rect 9663 2313 9697 2347
rect 9731 2313 9765 2347
rect 9799 2313 9833 2347
rect 9867 2313 9901 2347
rect 9935 2313 9969 2347
rect 10003 2313 10037 2347
rect 10071 2313 10105 2347
rect 10139 2313 10173 2347
rect 10207 2313 10241 2347
rect 10312 2313 10346 2347
rect 10380 2313 10414 2347
rect 10448 2313 10482 2347
rect 10516 2313 10550 2347
rect 10584 2313 10618 2347
rect 10652 2313 10686 2347
rect 10720 2313 10754 2347
rect 10788 2313 10822 2347
rect 10856 2313 10890 2347
rect 10924 2313 10958 2347
rect 10992 2313 11026 2347
rect 11060 2313 11094 2347
rect 11128 2313 11162 2347
rect 11196 2313 11230 2347
rect 11264 2313 11298 2347
rect 11332 2313 11366 2347
rect 11400 2313 11434 2347
rect 11468 2313 11502 2347
rect 11536 2313 11570 2347
rect 11652 2315 11686 2349
rect 11720 2315 11754 2349
rect 11788 2315 11822 2349
rect 11856 2315 11890 2349
rect 11924 2315 11958 2349
rect 11992 2315 12026 2349
rect 12060 2315 12094 2349
rect 12128 2315 12162 2349
rect 12196 2315 12230 2349
rect 12264 2315 12298 2349
rect 12332 2315 12366 2349
rect 12400 2315 12434 2349
rect 12468 2315 12502 2349
rect 12573 2310 12607 2344
rect 12641 2310 12675 2344
rect 12709 2310 12743 2344
rect 12777 2310 12811 2344
rect 12845 2310 12879 2344
rect 12913 2310 12947 2344
rect 12981 2310 13015 2344
rect 13049 2310 13083 2344
rect 13117 2310 13151 2344
rect 13185 2310 13219 2344
rect 13253 2310 13287 2344
rect 13321 2310 13355 2344
rect 8643 2244 8677 2278
rect 8711 2244 8745 2278
rect 8779 2244 8813 2278
rect 8847 2244 8881 2278
rect 8915 2244 8949 2278
rect 8983 2244 9017 2278
rect 9051 2244 9085 2278
rect 9119 2244 9153 2278
rect 9187 2244 9221 2278
rect 9255 2244 9289 2278
rect 9323 2244 9357 2278
rect 9391 2244 9425 2278
rect 9459 2244 9493 2278
rect 9527 2244 9561 2278
rect 9595 2244 9629 2278
rect 9663 2244 9697 2278
rect 9731 2244 9765 2278
rect 9799 2244 9833 2278
rect 9867 2244 9901 2278
rect 9935 2244 9969 2278
rect 10003 2244 10037 2278
rect 10071 2244 10105 2278
rect 10139 2244 10173 2278
rect 10207 2244 10241 2278
rect 10312 2244 10346 2278
rect 10380 2244 10414 2278
rect 10448 2244 10482 2278
rect 10516 2244 10550 2278
rect 10584 2244 10618 2278
rect 10652 2244 10686 2278
rect 10720 2244 10754 2278
rect 10788 2244 10822 2278
rect 10856 2244 10890 2278
rect 10924 2244 10958 2278
rect 10992 2244 11026 2278
rect 11060 2244 11094 2278
rect 11128 2244 11162 2278
rect 11196 2244 11230 2278
rect 11264 2244 11298 2278
rect 11332 2244 11366 2278
rect 11400 2244 11434 2278
rect 11468 2244 11502 2278
rect 11536 2244 11570 2278
rect 11652 2245 11686 2279
rect 11720 2245 11754 2279
rect 11788 2245 11822 2279
rect 11856 2245 11890 2279
rect 11924 2245 11958 2279
rect 11992 2245 12026 2279
rect 12060 2245 12094 2279
rect 12128 2245 12162 2279
rect 12196 2245 12230 2279
rect 12264 2245 12298 2279
rect 12332 2245 12366 2279
rect 12400 2245 12434 2279
rect 12468 2245 12502 2279
rect 12573 2241 12607 2275
rect 12641 2241 12675 2275
rect 12709 2241 12743 2275
rect 12777 2241 12811 2275
rect 12845 2241 12879 2275
rect 12913 2241 12947 2275
rect 12981 2241 13015 2275
rect 13049 2241 13083 2275
rect 13117 2241 13151 2275
rect 13185 2241 13219 2275
rect 13253 2241 13287 2275
rect 13321 2241 13355 2275
rect 1507 2099 1541 2133
rect 1575 2107 1609 2141
rect 1643 2107 1677 2141
rect 1507 2031 1541 2065
rect 1575 2038 1609 2072
rect 1643 2038 1677 2072
rect 1507 1963 1541 1997
rect 1575 1969 1609 2003
rect 1643 1969 1677 2003
rect 1507 1895 1541 1929
rect 1575 1900 1609 1934
rect 1643 1900 1677 1934
rect 1507 1827 1541 1861
rect 1575 1831 1609 1865
rect 1643 1831 1677 1865
rect 1507 1759 1541 1793
rect 1575 1762 1609 1796
rect 1643 1762 1677 1796
rect 1507 1691 1541 1725
rect 1575 1693 1609 1727
rect 1643 1693 1677 1727
rect 1507 1623 1541 1657
rect 1575 1624 1609 1658
rect 1643 1624 1677 1658
rect 8643 2175 8677 2209
rect 8711 2175 8745 2209
rect 8779 2175 8813 2209
rect 8847 2175 8881 2209
rect 8915 2175 8949 2209
rect 8983 2175 9017 2209
rect 9051 2175 9085 2209
rect 9119 2175 9153 2209
rect 9187 2175 9221 2209
rect 9255 2175 9289 2209
rect 9323 2175 9357 2209
rect 9391 2175 9425 2209
rect 9459 2175 9493 2209
rect 9527 2175 9561 2209
rect 9595 2175 9629 2209
rect 9663 2175 9697 2209
rect 9731 2175 9765 2209
rect 9799 2175 9833 2209
rect 9867 2175 9901 2209
rect 9935 2175 9969 2209
rect 10003 2175 10037 2209
rect 10071 2175 10105 2209
rect 10139 2175 10173 2209
rect 10207 2175 10241 2209
rect 10312 2175 10346 2209
rect 10380 2175 10414 2209
rect 10448 2175 10482 2209
rect 10516 2175 10550 2209
rect 10584 2175 10618 2209
rect 10652 2175 10686 2209
rect 10720 2175 10754 2209
rect 10788 2175 10822 2209
rect 10856 2175 10890 2209
rect 10924 2175 10958 2209
rect 10992 2175 11026 2209
rect 11060 2175 11094 2209
rect 11128 2175 11162 2209
rect 11196 2175 11230 2209
rect 11264 2175 11298 2209
rect 11332 2175 11366 2209
rect 11400 2175 11434 2209
rect 11468 2175 11502 2209
rect 11536 2175 11570 2209
rect 11652 2175 11686 2209
rect 11720 2175 11754 2209
rect 11788 2175 11822 2209
rect 11856 2175 11890 2209
rect 11924 2175 11958 2209
rect 11992 2175 12026 2209
rect 12060 2175 12094 2209
rect 12128 2175 12162 2209
rect 12196 2175 12230 2209
rect 12264 2175 12298 2209
rect 12332 2175 12366 2209
rect 12400 2175 12434 2209
rect 12468 2175 12502 2209
rect 12573 2172 12607 2206
rect 12641 2172 12675 2206
rect 12709 2172 12743 2206
rect 12777 2172 12811 2206
rect 12845 2172 12879 2206
rect 12913 2172 12947 2206
rect 12981 2172 13015 2206
rect 13049 2172 13083 2206
rect 13117 2172 13151 2206
rect 13185 2172 13219 2206
rect 13253 2172 13287 2206
rect 13321 2172 13355 2206
rect 8643 2106 8677 2140
rect 8711 2106 8745 2140
rect 8779 2106 8813 2140
rect 8847 2106 8881 2140
rect 8915 2106 8949 2140
rect 8983 2106 9017 2140
rect 9051 2106 9085 2140
rect 9119 2106 9153 2140
rect 9187 2106 9221 2140
rect 9255 2106 9289 2140
rect 9323 2106 9357 2140
rect 9391 2106 9425 2140
rect 9459 2106 9493 2140
rect 9527 2106 9561 2140
rect 9595 2106 9629 2140
rect 9663 2106 9697 2140
rect 9731 2106 9765 2140
rect 9799 2106 9833 2140
rect 9867 2106 9901 2140
rect 9935 2106 9969 2140
rect 10003 2106 10037 2140
rect 10071 2106 10105 2140
rect 10139 2106 10173 2140
rect 10207 2106 10241 2140
rect 10312 2106 10346 2140
rect 10380 2106 10414 2140
rect 10448 2106 10482 2140
rect 10516 2106 10550 2140
rect 10584 2106 10618 2140
rect 10652 2106 10686 2140
rect 10720 2106 10754 2140
rect 10788 2106 10822 2140
rect 10856 2106 10890 2140
rect 10924 2106 10958 2140
rect 10992 2106 11026 2140
rect 11060 2106 11094 2140
rect 11128 2106 11162 2140
rect 11196 2106 11230 2140
rect 11264 2106 11298 2140
rect 11332 2106 11366 2140
rect 11400 2106 11434 2140
rect 11468 2106 11502 2140
rect 11536 2106 11570 2140
rect 11652 2106 11686 2140
rect 11720 2106 11754 2140
rect 11788 2106 11822 2140
rect 11856 2106 11890 2140
rect 11924 2106 11958 2140
rect 11992 2106 12026 2140
rect 12060 2106 12094 2140
rect 12128 2106 12162 2140
rect 12196 2106 12230 2140
rect 12264 2106 12298 2140
rect 12332 2106 12366 2140
rect 12400 2106 12434 2140
rect 12468 2106 12502 2140
rect 12573 2103 12607 2137
rect 12641 2103 12675 2137
rect 12709 2103 12743 2137
rect 12777 2103 12811 2137
rect 12845 2103 12879 2137
rect 12913 2103 12947 2137
rect 12981 2103 13015 2137
rect 13049 2103 13083 2137
rect 13117 2103 13151 2137
rect 13185 2103 13219 2137
rect 13253 2103 13287 2137
rect 13321 2103 13355 2137
rect 8643 2037 8677 2071
rect 8711 2037 8745 2071
rect 8779 2037 8813 2071
rect 8847 2037 8881 2071
rect 8915 2037 8949 2071
rect 8983 2037 9017 2071
rect 9051 2037 9085 2071
rect 9119 2037 9153 2071
rect 9187 2037 9221 2071
rect 9255 2037 9289 2071
rect 9323 2037 9357 2071
rect 9391 2037 9425 2071
rect 9459 2037 9493 2071
rect 9527 2037 9561 2071
rect 9595 2037 9629 2071
rect 9663 2037 9697 2071
rect 9731 2037 9765 2071
rect 9799 2037 9833 2071
rect 9867 2037 9901 2071
rect 9935 2037 9969 2071
rect 10003 2037 10037 2071
rect 10071 2037 10105 2071
rect 10139 2037 10173 2071
rect 10207 2037 10241 2071
rect 10312 2037 10346 2071
rect 10380 2037 10414 2071
rect 10448 2037 10482 2071
rect 10516 2037 10550 2071
rect 10584 2037 10618 2071
rect 10652 2037 10686 2071
rect 10720 2037 10754 2071
rect 10788 2037 10822 2071
rect 10856 2037 10890 2071
rect 10924 2037 10958 2071
rect 10992 2037 11026 2071
rect 11060 2037 11094 2071
rect 11128 2037 11162 2071
rect 11196 2037 11230 2071
rect 11264 2037 11298 2071
rect 11332 2037 11366 2071
rect 11400 2037 11434 2071
rect 11468 2037 11502 2071
rect 11536 2037 11570 2071
rect 11652 2037 11686 2071
rect 11720 2037 11754 2071
rect 11788 2037 11822 2071
rect 11856 2037 11890 2071
rect 11924 2037 11958 2071
rect 11992 2037 12026 2071
rect 12060 2037 12094 2071
rect 12128 2037 12162 2071
rect 12196 2037 12230 2071
rect 12264 2037 12298 2071
rect 12332 2037 12366 2071
rect 12400 2037 12434 2071
rect 12468 2037 12502 2071
rect 12573 2034 12607 2068
rect 12641 2034 12675 2068
rect 12709 2034 12743 2068
rect 12777 2034 12811 2068
rect 12845 2034 12879 2068
rect 12913 2034 12947 2068
rect 12981 2034 13015 2068
rect 13049 2034 13083 2068
rect 13117 2034 13151 2068
rect 13185 2034 13219 2068
rect 13253 2034 13287 2068
rect 13321 2034 13355 2068
rect 8643 1968 8677 2002
rect 8711 1968 8745 2002
rect 8779 1968 8813 2002
rect 8847 1968 8881 2002
rect 8915 1968 8949 2002
rect 8983 1968 9017 2002
rect 9051 1968 9085 2002
rect 9119 1968 9153 2002
rect 9187 1968 9221 2002
rect 9255 1968 9289 2002
rect 9323 1968 9357 2002
rect 9391 1968 9425 2002
rect 9459 1968 9493 2002
rect 9527 1968 9561 2002
rect 9595 1968 9629 2002
rect 9663 1968 9697 2002
rect 9731 1968 9765 2002
rect 9799 1968 9833 2002
rect 9867 1968 9901 2002
rect 9935 1968 9969 2002
rect 10003 1968 10037 2002
rect 10071 1968 10105 2002
rect 10139 1968 10173 2002
rect 10207 1968 10241 2002
rect 10312 1968 10346 2002
rect 10380 1968 10414 2002
rect 10448 1968 10482 2002
rect 10516 1968 10550 2002
rect 10584 1968 10618 2002
rect 10652 1968 10686 2002
rect 10720 1968 10754 2002
rect 10788 1968 10822 2002
rect 10856 1968 10890 2002
rect 10924 1968 10958 2002
rect 10992 1968 11026 2002
rect 11060 1968 11094 2002
rect 11128 1968 11162 2002
rect 11196 1968 11230 2002
rect 11264 1968 11298 2002
rect 11332 1968 11366 2002
rect 11400 1968 11434 2002
rect 11468 1968 11502 2002
rect 11536 1968 11570 2002
rect 11652 1968 11686 2002
rect 11720 1968 11754 2002
rect 11788 1968 11822 2002
rect 11856 1968 11890 2002
rect 11924 1968 11958 2002
rect 11992 1968 12026 2002
rect 12060 1968 12094 2002
rect 12128 1968 12162 2002
rect 12196 1968 12230 2002
rect 12264 1968 12298 2002
rect 12332 1968 12366 2002
rect 12400 1968 12434 2002
rect 12468 1968 12502 2002
rect 12573 1965 12607 1999
rect 12641 1965 12675 1999
rect 12709 1965 12743 1999
rect 12777 1965 12811 1999
rect 12845 1965 12879 1999
rect 12913 1965 12947 1999
rect 12981 1965 13015 1999
rect 13049 1965 13083 1999
rect 13117 1965 13151 1999
rect 13185 1965 13219 1999
rect 13253 1965 13287 1999
rect 13321 1965 13355 1999
rect 8643 1899 8677 1933
rect 8711 1899 8745 1933
rect 8779 1899 8813 1933
rect 8847 1899 8881 1933
rect 8915 1899 8949 1933
rect 8983 1899 9017 1933
rect 9051 1899 9085 1933
rect 9119 1899 9153 1933
rect 9187 1899 9221 1933
rect 9255 1899 9289 1933
rect 9323 1899 9357 1933
rect 9391 1899 9425 1933
rect 9459 1899 9493 1933
rect 9527 1899 9561 1933
rect 9595 1899 9629 1933
rect 9663 1899 9697 1933
rect 9731 1899 9765 1933
rect 9799 1899 9833 1933
rect 9867 1899 9901 1933
rect 9935 1899 9969 1933
rect 10003 1899 10037 1933
rect 10071 1899 10105 1933
rect 10139 1899 10173 1933
rect 10207 1899 10241 1933
rect 10312 1899 10346 1933
rect 10380 1899 10414 1933
rect 10448 1899 10482 1933
rect 10516 1899 10550 1933
rect 10584 1899 10618 1933
rect 10652 1899 10686 1933
rect 10720 1899 10754 1933
rect 10788 1899 10822 1933
rect 10856 1899 10890 1933
rect 10924 1899 10958 1933
rect 10992 1899 11026 1933
rect 11060 1899 11094 1933
rect 11128 1899 11162 1933
rect 11196 1899 11230 1933
rect 11264 1899 11298 1933
rect 11332 1899 11366 1933
rect 11400 1899 11434 1933
rect 11468 1899 11502 1933
rect 11536 1899 11570 1933
rect 11652 1899 11686 1933
rect 11720 1899 11754 1933
rect 11788 1899 11822 1933
rect 11856 1899 11890 1933
rect 11924 1899 11958 1933
rect 11992 1899 12026 1933
rect 12060 1899 12094 1933
rect 12128 1899 12162 1933
rect 12196 1899 12230 1933
rect 12264 1899 12298 1933
rect 12332 1899 12366 1933
rect 12400 1899 12434 1933
rect 12468 1899 12502 1933
rect 12573 1896 12607 1930
rect 12641 1896 12675 1930
rect 12709 1896 12743 1930
rect 12777 1896 12811 1930
rect 12845 1896 12879 1930
rect 12913 1896 12947 1930
rect 12981 1896 13015 1930
rect 13049 1896 13083 1930
rect 13117 1896 13151 1930
rect 13185 1896 13219 1930
rect 13253 1896 13287 1930
rect 13321 1896 13355 1930
rect 8643 1830 8677 1864
rect 8711 1830 8745 1864
rect 8779 1830 8813 1864
rect 8847 1830 8881 1864
rect 8915 1830 8949 1864
rect 8983 1830 9017 1864
rect 9051 1830 9085 1864
rect 9119 1830 9153 1864
rect 9187 1830 9221 1864
rect 9255 1830 9289 1864
rect 9323 1830 9357 1864
rect 9391 1830 9425 1864
rect 9459 1830 9493 1864
rect 9527 1830 9561 1864
rect 9595 1830 9629 1864
rect 9663 1830 9697 1864
rect 9731 1830 9765 1864
rect 9799 1830 9833 1864
rect 9867 1830 9901 1864
rect 9935 1830 9969 1864
rect 10003 1830 10037 1864
rect 10071 1830 10105 1864
rect 10139 1830 10173 1864
rect 10207 1830 10241 1864
rect 10312 1830 10346 1864
rect 10380 1830 10414 1864
rect 10448 1830 10482 1864
rect 10516 1830 10550 1864
rect 10584 1830 10618 1864
rect 10652 1830 10686 1864
rect 10720 1830 10754 1864
rect 10788 1830 10822 1864
rect 10856 1830 10890 1864
rect 10924 1830 10958 1864
rect 10992 1830 11026 1864
rect 11060 1830 11094 1864
rect 11128 1830 11162 1864
rect 11196 1830 11230 1864
rect 11264 1830 11298 1864
rect 11332 1830 11366 1864
rect 11400 1830 11434 1864
rect 11468 1830 11502 1864
rect 11536 1830 11570 1864
rect 11652 1830 11686 1864
rect 11720 1830 11754 1864
rect 11788 1830 11822 1864
rect 11856 1830 11890 1864
rect 11924 1830 11958 1864
rect 11992 1830 12026 1864
rect 12060 1830 12094 1864
rect 12128 1830 12162 1864
rect 12196 1830 12230 1864
rect 12264 1830 12298 1864
rect 12332 1830 12366 1864
rect 12400 1830 12434 1864
rect 12468 1830 12502 1864
rect 8643 1761 8677 1795
rect 8711 1761 8745 1795
rect 8779 1761 8813 1795
rect 8847 1761 8881 1795
rect 8915 1761 8949 1795
rect 8983 1761 9017 1795
rect 9051 1761 9085 1795
rect 9119 1761 9153 1795
rect 9187 1761 9221 1795
rect 9255 1761 9289 1795
rect 9323 1761 9357 1795
rect 9391 1761 9425 1795
rect 9459 1761 9493 1795
rect 9527 1761 9561 1795
rect 9595 1761 9629 1795
rect 9663 1761 9697 1795
rect 9731 1761 9765 1795
rect 9799 1761 9833 1795
rect 9867 1761 9901 1795
rect 9935 1761 9969 1795
rect 10003 1761 10037 1795
rect 10071 1761 10105 1795
rect 10139 1761 10173 1795
rect 10207 1761 10241 1795
rect 10312 1761 10346 1795
rect 10380 1761 10414 1795
rect 10448 1761 10482 1795
rect 10516 1761 10550 1795
rect 10584 1761 10618 1795
rect 10652 1761 10686 1795
rect 10720 1761 10754 1795
rect 10788 1761 10822 1795
rect 10856 1761 10890 1795
rect 10924 1761 10958 1795
rect 10992 1761 11026 1795
rect 11060 1761 11094 1795
rect 11128 1761 11162 1795
rect 11196 1761 11230 1795
rect 11264 1761 11298 1795
rect 11332 1761 11366 1795
rect 11400 1761 11434 1795
rect 11468 1761 11502 1795
rect 11536 1761 11570 1795
rect 11652 1761 11686 1795
rect 11720 1761 11754 1795
rect 11788 1761 11822 1795
rect 11856 1761 11890 1795
rect 11924 1761 11958 1795
rect 11992 1761 12026 1795
rect 12060 1761 12094 1795
rect 12128 1761 12162 1795
rect 12196 1761 12230 1795
rect 12264 1761 12298 1795
rect 12332 1761 12366 1795
rect 12400 1761 12434 1795
rect 12468 1761 12502 1795
rect 8643 1692 8677 1726
rect 8711 1692 8745 1726
rect 8779 1692 8813 1726
rect 8847 1692 8881 1726
rect 8915 1692 8949 1726
rect 8983 1692 9017 1726
rect 9051 1692 9085 1726
rect 9119 1692 9153 1726
rect 9187 1692 9221 1726
rect 9255 1692 9289 1726
rect 9323 1692 9357 1726
rect 9391 1692 9425 1726
rect 9459 1692 9493 1726
rect 9527 1692 9561 1726
rect 9595 1692 9629 1726
rect 9663 1692 9697 1726
rect 9731 1692 9765 1726
rect 9799 1692 9833 1726
rect 9867 1692 9901 1726
rect 9935 1692 9969 1726
rect 10003 1692 10037 1726
rect 10071 1692 10105 1726
rect 10139 1692 10173 1726
rect 10207 1692 10241 1726
rect 10312 1692 10346 1726
rect 10380 1692 10414 1726
rect 10448 1692 10482 1726
rect 10516 1692 10550 1726
rect 10584 1692 10618 1726
rect 10652 1692 10686 1726
rect 10720 1692 10754 1726
rect 10788 1692 10822 1726
rect 10856 1692 10890 1726
rect 10924 1692 10958 1726
rect 10992 1692 11026 1726
rect 11060 1692 11094 1726
rect 11128 1692 11162 1726
rect 11196 1692 11230 1726
rect 11264 1692 11298 1726
rect 11332 1692 11366 1726
rect 11400 1692 11434 1726
rect 11468 1692 11502 1726
rect 11536 1692 11570 1726
rect 11652 1692 11686 1726
rect 11720 1692 11754 1726
rect 11788 1692 11822 1726
rect 11856 1692 11890 1726
rect 11924 1692 11958 1726
rect 11992 1692 12026 1726
rect 12060 1692 12094 1726
rect 12128 1692 12162 1726
rect 12196 1692 12230 1726
rect 12264 1692 12298 1726
rect 12332 1692 12366 1726
rect 12400 1692 12434 1726
rect 12468 1692 12502 1726
rect 8643 1623 8677 1657
rect 8711 1623 8745 1657
rect 8779 1623 8813 1657
rect 8847 1623 8881 1657
rect 8915 1623 8949 1657
rect 8983 1623 9017 1657
rect 9051 1623 9085 1657
rect 9119 1623 9153 1657
rect 9187 1623 9221 1657
rect 9255 1623 9289 1657
rect 9323 1623 9357 1657
rect 9391 1623 9425 1657
rect 9459 1623 9493 1657
rect 9527 1623 9561 1657
rect 9595 1623 9629 1657
rect 9663 1623 9697 1657
rect 9731 1623 9765 1657
rect 9799 1623 9833 1657
rect 9867 1623 9901 1657
rect 9935 1623 9969 1657
rect 10003 1623 10037 1657
rect 10071 1623 10105 1657
rect 10139 1623 10173 1657
rect 10207 1623 10241 1657
rect 10312 1623 10346 1657
rect 10380 1623 10414 1657
rect 10448 1623 10482 1657
rect 10516 1623 10550 1657
rect 10584 1623 10618 1657
rect 10652 1623 10686 1657
rect 10720 1623 10754 1657
rect 10788 1623 10822 1657
rect 10856 1623 10890 1657
rect 10924 1623 10958 1657
rect 10992 1623 11026 1657
rect 11060 1623 11094 1657
rect 11128 1623 11162 1657
rect 11196 1623 11230 1657
rect 11264 1623 11298 1657
rect 11332 1623 11366 1657
rect 11400 1623 11434 1657
rect 11468 1623 11502 1657
rect 11536 1623 11570 1657
rect 11652 1623 11686 1657
rect 11720 1623 11754 1657
rect 11788 1623 11822 1657
rect 11856 1623 11890 1657
rect 11924 1623 11958 1657
rect 11992 1623 12026 1657
rect 12060 1623 12094 1657
rect 12128 1623 12162 1657
rect 12196 1623 12230 1657
rect 12264 1623 12298 1657
rect 12332 1623 12366 1657
rect 12400 1623 12434 1657
rect 12468 1623 12502 1657
rect 12573 1623 13355 1861
rect 1507 1555 1541 1589
rect 1575 1555 1609 1589
rect 1643 1555 1677 1589
rect 8412 1555 8446 1589
rect 8482 1555 8516 1589
rect 8552 1555 8586 1589
rect 8622 1555 8656 1589
rect 8692 1555 8726 1589
rect 8762 1555 8796 1589
rect 8832 1555 8866 1589
rect 8902 1555 8936 1589
rect 8972 1555 9006 1589
rect 9043 1555 9077 1589
rect 9114 1555 9148 1589
rect 9185 1555 9219 1589
rect 9256 1555 9290 1589
rect 9327 1555 9361 1589
rect 9398 1555 9432 1589
rect 9469 1555 9503 1589
rect 9540 1555 9574 1589
rect 9611 1555 9645 1589
rect 9682 1555 9716 1589
rect 9753 1555 9787 1589
rect 9824 1555 9858 1589
rect 9895 1555 9929 1589
rect 9966 1555 10000 1589
rect 1531 1487 1565 1521
rect 1600 1487 1634 1521
rect 1669 1487 1703 1521
rect 1738 1487 1772 1521
rect 1807 1487 1841 1521
rect 1876 1487 1910 1521
rect 1945 1487 1979 1521
rect 2014 1487 2048 1521
rect 2083 1487 2117 1521
rect 2152 1487 2186 1521
rect 2221 1487 2255 1521
rect 2290 1487 2324 1521
rect 2359 1487 2393 1521
rect 2428 1487 2462 1521
rect 2497 1487 2531 1521
rect 2566 1487 2600 1521
rect 2635 1487 2669 1521
rect 2704 1487 2738 1521
rect 2773 1487 2807 1521
rect 2842 1487 2876 1521
rect 2911 1487 2945 1521
rect 2980 1487 3014 1521
rect 3049 1487 3083 1521
rect 3118 1487 3152 1521
rect 3187 1487 3221 1521
rect 3256 1487 3290 1521
rect 3325 1487 3359 1521
rect 3394 1487 3428 1521
rect 3463 1487 3497 1521
rect 3532 1487 3566 1521
rect 3601 1487 3635 1521
rect 3670 1487 3704 1521
rect 3739 1487 3773 1521
rect 3808 1487 3842 1521
rect 3877 1487 3911 1521
rect 3946 1487 3980 1521
rect 4015 1487 4049 1521
rect 4084 1487 4118 1521
rect 4153 1487 4187 1521
rect 4222 1487 4256 1521
rect 4291 1487 4325 1521
rect 4360 1487 4394 1521
rect 4429 1487 4463 1521
rect 4498 1487 4532 1521
rect 4567 1487 4601 1521
rect 4636 1487 4670 1521
rect 4705 1487 4739 1521
rect 4774 1487 4808 1521
rect 4843 1487 4877 1521
rect 4912 1487 4946 1521
rect 4981 1487 5015 1521
rect 5050 1487 5084 1521
rect 5119 1487 5153 1521
rect 5188 1487 5222 1521
rect 5257 1487 5291 1521
rect 5326 1487 5360 1521
rect 5395 1487 5429 1521
rect 5464 1487 5498 1521
rect 5533 1487 5567 1521
rect 5602 1487 5636 1521
rect 5671 1487 5705 1521
rect 5740 1487 5774 1521
rect 5809 1487 5843 1521
rect 5878 1487 5912 1521
rect 5947 1487 5981 1521
rect 6016 1487 6050 1521
rect 6085 1487 6119 1521
rect 1531 1419 1565 1453
rect 1600 1419 1634 1453
rect 1669 1419 1703 1453
rect 1738 1419 1772 1453
rect 1807 1419 1841 1453
rect 1876 1419 1910 1453
rect 1945 1419 1979 1453
rect 2014 1419 2048 1453
rect 2083 1419 2117 1453
rect 2152 1419 2186 1453
rect 2221 1419 2255 1453
rect 2290 1419 2324 1453
rect 2359 1419 2393 1453
rect 2428 1419 2462 1453
rect 2497 1419 2531 1453
rect 2566 1419 2600 1453
rect 2635 1419 2669 1453
rect 2704 1419 2738 1453
rect 2773 1419 2807 1453
rect 2842 1419 2876 1453
rect 2911 1419 2945 1453
rect 2980 1419 3014 1453
rect 3049 1419 3083 1453
rect 3118 1419 3152 1453
rect 3187 1419 3221 1453
rect 3256 1419 3290 1453
rect 3325 1419 3359 1453
rect 3394 1419 3428 1453
rect 3463 1419 3497 1453
rect 3532 1419 3566 1453
rect 3601 1419 3635 1453
rect 3670 1419 3704 1453
rect 3739 1419 3773 1453
rect 3808 1419 3842 1453
rect 3877 1419 3911 1453
rect 3946 1419 3980 1453
rect 4015 1419 4049 1453
rect 4084 1419 4118 1453
rect 4153 1419 4187 1453
rect 4222 1419 4256 1453
rect 4291 1419 4325 1453
rect 4360 1419 4394 1453
rect 4429 1419 4463 1453
rect 4498 1419 4532 1453
rect 4567 1419 4601 1453
rect 4636 1419 4670 1453
rect 4705 1419 4739 1453
rect 4774 1419 4808 1453
rect 4843 1419 4877 1453
rect 4912 1419 4946 1453
rect 4981 1419 5015 1453
rect 5050 1419 5084 1453
rect 5119 1419 5153 1453
rect 5188 1419 5222 1453
rect 5257 1419 5291 1453
rect 5326 1419 5360 1453
rect 5395 1419 5429 1453
rect 5464 1419 5498 1453
rect 5533 1419 5567 1453
rect 5602 1419 5636 1453
rect 5671 1419 5705 1453
rect 5740 1419 5774 1453
rect 5809 1419 5843 1453
rect 5878 1419 5912 1453
rect 5947 1419 5981 1453
rect 6016 1419 6050 1453
rect 6085 1419 6119 1453
rect 6154 1419 8364 1521
rect 8412 1487 8446 1521
rect 8482 1487 8516 1521
rect 8552 1487 8586 1521
rect 8622 1487 8656 1521
rect 8692 1487 8726 1521
rect 8762 1487 8796 1521
rect 8832 1487 8866 1521
rect 8902 1487 8936 1521
rect 8972 1487 9006 1521
rect 9043 1487 9077 1521
rect 9114 1487 9148 1521
rect 9185 1487 9219 1521
rect 9256 1487 9290 1521
rect 9327 1487 9361 1521
rect 9398 1487 9432 1521
rect 9469 1487 9503 1521
rect 9540 1487 9574 1521
rect 9611 1487 9645 1521
rect 9682 1487 9716 1521
rect 9753 1487 9787 1521
rect 9824 1487 9858 1521
rect 9895 1487 9929 1521
rect 9966 1487 10000 1521
rect 8412 1419 8446 1453
rect 8482 1419 8516 1453
rect 8552 1419 8586 1453
rect 8622 1419 8656 1453
rect 8692 1419 8726 1453
rect 8762 1419 8796 1453
rect 8832 1419 8866 1453
rect 8902 1419 8936 1453
rect 8972 1419 9006 1453
rect 9043 1419 9077 1453
rect 9114 1419 9148 1453
rect 9185 1419 9219 1453
rect 9256 1419 9290 1453
rect 9327 1419 9361 1453
rect 9398 1419 9432 1453
rect 9469 1419 9503 1453
rect 9540 1419 9574 1453
rect 9611 1419 9645 1453
rect 9682 1419 9716 1453
rect 9753 1419 9787 1453
rect 9824 1419 9858 1453
rect 9895 1419 9929 1453
rect 9966 1419 10000 1453
rect 23949 4694 24119 5532
rect 24153 5488 24187 5522
rect 24221 5488 24255 5522
rect 24289 5488 24323 5522
rect 24357 5488 24391 5522
rect 24425 5488 24459 5522
rect 24493 5488 24527 5522
rect 24153 5419 24187 5453
rect 24221 5419 24255 5453
rect 24289 5419 24323 5453
rect 24357 5419 24391 5453
rect 24425 5419 24459 5453
rect 24493 5419 24527 5453
rect 24153 5350 24187 5384
rect 24221 5350 24255 5384
rect 24289 5350 24323 5384
rect 24357 5350 24391 5384
rect 24425 5350 24459 5384
rect 24493 5350 24527 5384
rect 24153 5281 24187 5315
rect 24221 5281 24255 5315
rect 24289 5281 24323 5315
rect 24357 5281 24391 5315
rect 24425 5281 24459 5315
rect 24493 5281 24527 5315
rect 24153 5212 24187 5246
rect 24221 5212 24255 5246
rect 24289 5212 24323 5246
rect 24357 5212 24391 5246
rect 24425 5212 24459 5246
rect 24493 5212 24527 5246
rect 24153 5143 24187 5177
rect 24221 5143 24255 5177
rect 24289 5143 24323 5177
rect 24357 5143 24391 5177
rect 24425 5143 24459 5177
rect 24493 5143 24527 5177
rect 24153 5074 24187 5108
rect 24221 5074 24255 5108
rect 24289 5074 24323 5108
rect 24357 5074 24391 5108
rect 24425 5074 24459 5108
rect 24493 5074 24527 5108
rect 24153 5005 24187 5039
rect 24221 5005 24255 5039
rect 24289 5005 24323 5039
rect 24357 5005 24391 5039
rect 24425 5005 24459 5039
rect 24493 5005 24527 5039
rect 24153 4936 24187 4970
rect 24221 4936 24255 4970
rect 24289 4936 24323 4970
rect 24357 4936 24391 4970
rect 24425 4936 24459 4970
rect 24493 4936 24527 4970
rect 24153 4867 24187 4901
rect 24221 4867 24255 4901
rect 24289 4867 24323 4901
rect 24357 4867 24391 4901
rect 24425 4867 24459 4901
rect 24493 4867 24527 4901
rect 24153 4798 24187 4832
rect 24221 4798 24255 4832
rect 24289 4798 24323 4832
rect 24357 4798 24391 4832
rect 24425 4798 24459 4832
rect 24493 4798 24527 4832
rect 24153 4729 24187 4763
rect 24221 4729 24255 4763
rect 24289 4729 24323 4763
rect 24357 4729 24391 4763
rect 24425 4729 24459 4763
rect 24493 4729 24527 4763
rect 23949 2348 24527 4694
rect 23949 1010 24119 2348
rect 23949 976 24095 1010
rect 20558 942 20592 976
rect 20627 942 20661 976
rect 20696 942 20730 976
rect 20765 942 20799 976
rect 20834 942 20868 976
rect 20903 942 20937 976
rect 20972 942 21006 976
rect 21041 942 21075 976
rect 21110 942 21144 976
rect 21179 942 21213 976
rect 21248 942 21282 976
rect 21317 942 21351 976
rect 21386 942 21420 976
rect 21455 942 21489 976
rect 21524 942 21558 976
rect 21593 942 21627 976
rect 21662 942 21696 976
rect 21731 942 21765 976
rect 21800 942 21834 976
rect 21869 942 21903 976
rect 21938 942 21972 976
rect 22007 942 22041 976
rect 22076 942 22110 976
rect 22145 942 22179 976
rect 22214 942 22248 976
rect 22283 942 22317 976
rect 22352 942 22386 976
rect 22421 942 22455 976
rect 22490 942 22524 976
rect 22559 942 22593 976
rect 22628 942 22662 976
rect 22697 942 22731 976
rect 22766 942 22800 976
rect 22835 942 22869 976
rect 22904 942 22938 976
rect 20558 874 20592 908
rect 20627 874 20661 908
rect 20696 874 20730 908
rect 20765 874 20799 908
rect 20834 874 20868 908
rect 20903 874 20937 908
rect 20972 874 21006 908
rect 21041 874 21075 908
rect 21110 874 21144 908
rect 21179 874 21213 908
rect 21248 874 21282 908
rect 21317 874 21351 908
rect 21386 874 21420 908
rect 21455 874 21489 908
rect 21524 874 21558 908
rect 21593 874 21627 908
rect 21662 874 21696 908
rect 21731 874 21765 908
rect 21800 874 21834 908
rect 21869 874 21903 908
rect 21938 874 21972 908
rect 22007 874 22041 908
rect 22076 874 22110 908
rect 22145 874 22179 908
rect 22214 874 22248 908
rect 22283 874 22317 908
rect 22352 874 22386 908
rect 22421 874 22455 908
rect 22490 874 22524 908
rect 22559 874 22593 908
rect 22628 874 22662 908
rect 22697 874 22731 908
rect 22766 874 22800 908
rect 22835 874 22869 908
rect 22904 874 22938 908
rect 278 788 312 822
rect 346 788 380 822
rect 414 788 448 822
rect 20558 806 20592 840
rect 20627 806 20661 840
rect 20696 806 20730 840
rect 20765 806 20799 840
rect 20834 806 20868 840
rect 20903 806 20937 840
rect 20972 806 21006 840
rect 21041 806 21075 840
rect 21110 806 21144 840
rect 21179 806 21213 840
rect 21248 806 21282 840
rect 21317 806 21351 840
rect 21386 806 21420 840
rect 21455 806 21489 840
rect 21524 806 21558 840
rect 21593 806 21627 840
rect 21662 806 21696 840
rect 21731 806 21765 840
rect 21800 806 21834 840
rect 21869 806 21903 840
rect 21938 806 21972 840
rect 22007 806 22041 840
rect 22076 806 22110 840
rect 22145 806 22179 840
rect 22214 806 22248 840
rect 22283 806 22317 840
rect 22352 806 22386 840
rect 22421 806 22455 840
rect 22490 806 22524 840
rect 22559 806 22593 840
rect 22628 806 22662 840
rect 22697 806 22731 840
rect 22766 806 22800 840
rect 22835 806 22869 840
rect 22904 806 22938 840
rect 22973 806 24095 976
rect 278 719 312 753
rect 346 719 380 753
rect 414 719 448 753
rect 278 650 312 684
rect 346 650 380 684
rect 414 650 448 684
rect 278 581 312 615
rect 346 581 380 615
rect 414 581 448 615
rect 278 512 312 546
rect 346 512 380 546
rect 414 512 448 546
rect 278 443 312 477
rect 346 443 380 477
rect 414 443 448 477
rect 278 374 312 408
rect 346 374 380 408
rect 414 374 448 408
rect 278 305 312 339
rect 346 305 380 339
rect 414 305 448 339
rect 278 236 312 270
rect 346 236 380 270
rect 414 236 448 270
rect 278 167 312 201
rect 346 167 380 201
rect 414 167 448 201
<< poly >>
rect 3994 4076 4062 4093
rect 1786 4060 1920 4076
rect 1786 4026 1802 4060
rect 1836 4026 1870 4060
rect 1904 4026 1920 4060
rect 1786 4010 1920 4026
rect 3928 4060 4062 4076
rect 3928 4026 3944 4060
rect 3978 4026 4012 4060
rect 4046 4026 4062 4060
rect 3928 4010 4062 4026
rect 3994 3993 4062 4010
rect 16960 4273 17028 4290
rect 19168 4273 19236 4290
rect 16960 4257 17094 4273
rect 16960 4223 16976 4257
rect 17010 4223 17044 4257
rect 17078 4223 17094 4257
rect 16960 4207 17094 4223
rect 19102 4257 19236 4273
rect 19102 4223 19118 4257
rect 19152 4223 19186 4257
rect 19220 4223 19236 4257
rect 19102 4207 19236 4223
rect 16960 4190 17028 4207
rect 19168 4190 19236 4207
<< polycont >>
rect 1802 4026 1836 4060
rect 1870 4026 1904 4060
rect 3944 4026 3978 4060
rect 4012 4026 4046 4060
rect 16976 4223 17010 4257
rect 17044 4223 17078 4257
rect 19118 4223 19152 4257
rect 19186 4223 19220 4257
<< locali >>
rect 24370 9395 24540 9419
rect 22766 9342 23600 9372
rect 22766 9318 24159 9342
rect 22766 9295 23638 9318
rect 22766 9261 22818 9295
rect 22852 9261 22886 9295
rect 22920 9261 22954 9295
rect 22988 9261 23022 9295
rect 23056 9261 23090 9295
rect 23124 9261 23158 9295
rect 23192 9261 23226 9295
rect 23260 9261 23294 9295
rect 23328 9261 23362 9295
rect 23396 9261 23430 9295
rect 23464 9261 23498 9295
rect 23532 9261 23566 9295
rect 23600 9284 23638 9295
rect 23672 9284 23706 9318
rect 23740 9284 23774 9318
rect 23808 9284 23842 9318
rect 23876 9284 23910 9318
rect 23944 9284 23978 9318
rect 24012 9284 24046 9318
rect 24080 9284 24114 9318
rect 24148 9284 24159 9318
rect 23600 9261 24159 9284
rect 22766 9245 24159 9261
rect 22766 9226 23638 9245
rect 22766 9192 22818 9226
rect 22852 9192 22886 9226
rect 22920 9192 22954 9226
rect 22988 9192 23022 9226
rect 23056 9192 23090 9226
rect 23124 9192 23158 9226
rect 23192 9192 23226 9226
rect 23260 9192 23294 9226
rect 23328 9192 23362 9226
rect 23396 9192 23430 9226
rect 23464 9192 23498 9226
rect 23532 9192 23566 9226
rect 23600 9211 23638 9226
rect 23672 9211 23706 9245
rect 23740 9211 23774 9245
rect 23808 9211 23842 9245
rect 23876 9211 23910 9245
rect 23944 9211 23978 9245
rect 24012 9211 24046 9245
rect 24080 9211 24114 9245
rect 24148 9211 24159 9245
rect 23600 9192 24159 9211
rect 22766 9172 24159 9192
rect 22766 9157 23638 9172
rect 22766 9123 22818 9157
rect 22852 9123 22886 9157
rect 22920 9123 22954 9157
rect 22988 9123 23022 9157
rect 23056 9123 23090 9157
rect 23124 9123 23158 9157
rect 23192 9123 23226 9157
rect 23260 9123 23294 9157
rect 23328 9123 23362 9157
rect 23396 9123 23430 9157
rect 23464 9123 23498 9157
rect 23532 9123 23566 9157
rect 23600 9138 23638 9157
rect 23672 9138 23706 9172
rect 23740 9138 23774 9172
rect 23808 9138 23842 9172
rect 23876 9138 23910 9172
rect 23944 9138 23978 9172
rect 24012 9138 24046 9172
rect 24080 9138 24114 9172
rect 24148 9138 24159 9172
rect 23600 9123 24159 9138
rect 22766 9099 24159 9123
rect 22766 9088 23638 9099
rect 22766 9054 22818 9088
rect 22852 9054 22886 9088
rect 22920 9054 22954 9088
rect 22988 9054 23022 9088
rect 23056 9054 23090 9088
rect 23124 9054 23158 9088
rect 23192 9054 23226 9088
rect 23260 9054 23294 9088
rect 23328 9054 23362 9088
rect 23396 9054 23430 9088
rect 23464 9054 23498 9088
rect 23532 9054 23566 9088
rect 23600 9065 23638 9088
rect 23672 9065 23706 9099
rect 23740 9065 23774 9099
rect 23808 9065 23842 9099
rect 23876 9065 23910 9099
rect 23944 9065 23978 9099
rect 24012 9065 24046 9099
rect 24080 9065 24114 9099
rect 24148 9065 24159 9099
rect 23600 9054 24159 9065
rect 22766 9025 24159 9054
rect 22766 9019 23638 9025
rect 22766 8997 22818 9019
rect 22852 8997 22886 9019
rect 22920 8997 22954 9019
rect 22988 8997 23022 9019
rect 23056 8997 23090 9019
rect 23124 8997 23158 9019
rect 23192 8997 23226 9019
rect 23260 8997 23294 9019
rect 23328 8997 23362 9019
rect 23396 8997 23430 9019
rect 23464 8997 23498 9019
rect 22766 8603 22798 8997
rect 23480 8985 23498 8997
rect 23532 8985 23566 9019
rect 23600 8991 23638 9019
rect 23672 8991 23706 9025
rect 23740 8991 23774 9025
rect 23808 8991 23842 9025
rect 23876 8991 23910 9025
rect 23944 8991 23978 9025
rect 24012 8991 24046 9025
rect 24080 8991 24114 9025
rect 24148 8991 24159 9025
rect 23600 8985 24159 8991
rect 23480 8951 24159 8985
rect 23480 8950 23638 8951
rect 23480 8916 23498 8950
rect 23532 8916 23566 8950
rect 23600 8917 23638 8950
rect 23672 8917 23706 8951
rect 23740 8917 23774 8951
rect 23808 8917 23842 8951
rect 23876 8917 23910 8951
rect 23944 8917 23978 8951
rect 24012 8917 24046 8951
rect 24080 8917 24114 8951
rect 24148 8917 24159 8951
rect 23600 8916 24159 8917
rect 23480 8881 24159 8916
rect 23480 8847 23498 8881
rect 23532 8847 23566 8881
rect 23600 8877 24159 8881
rect 23600 8847 23638 8877
rect 23480 8843 23638 8847
rect 23672 8843 23706 8877
rect 23740 8843 23774 8877
rect 23808 8843 23842 8877
rect 23876 8843 23910 8877
rect 23944 8843 23978 8877
rect 24012 8843 24046 8877
rect 24080 8843 24114 8877
rect 24148 8843 24159 8877
rect 23480 8812 24159 8843
rect 23480 8778 23498 8812
rect 23532 8778 23566 8812
rect 23600 8803 24159 8812
rect 23600 8778 23638 8803
rect 23480 8769 23638 8778
rect 23672 8769 23706 8803
rect 23740 8769 23774 8803
rect 23808 8769 23842 8803
rect 23876 8769 23910 8803
rect 23944 8769 23978 8803
rect 24012 8769 24046 8803
rect 24080 8769 24114 8803
rect 24148 8769 24159 8803
rect 23480 8745 24159 8769
rect 24370 9121 24540 9157
rect 24404 9087 24438 9121
rect 24472 9087 24506 9121
rect 24370 9051 24540 9087
rect 24404 9017 24438 9051
rect 24472 9017 24506 9051
rect 24370 8981 24540 9017
rect 24404 8947 24438 8981
rect 24472 8947 24506 8981
rect 24370 8912 24540 8947
rect 24404 8878 24438 8912
rect 24472 8878 24506 8912
rect 24370 8843 24540 8878
rect 24404 8809 24438 8843
rect 24472 8809 24506 8843
rect 24370 8774 24540 8809
rect 23480 8743 23600 8745
rect 23480 8709 23498 8743
rect 23532 8709 23566 8743
rect 23480 8674 23600 8709
rect 24404 8740 24438 8774
rect 24472 8740 24506 8774
rect 24370 8705 24540 8740
rect 24404 8680 24438 8705
rect 24472 8680 24506 8705
rect 23480 8640 23498 8674
rect 23532 8640 23566 8674
rect 23480 8605 23600 8640
rect 23480 8603 23498 8605
rect 22766 8571 22818 8603
rect 22852 8571 22886 8603
rect 22920 8571 22954 8603
rect 22988 8571 23022 8603
rect 23056 8571 23090 8603
rect 23124 8571 23158 8603
rect 23192 8571 23226 8603
rect 23260 8571 23294 8603
rect 23328 8571 23362 8603
rect 23396 8571 23430 8603
rect 23464 8571 23498 8603
rect 23532 8571 23566 8605
rect 24535 8636 24540 8671
rect 22766 8564 23600 8571
rect 22766 8530 22798 8564
rect 22832 8536 22870 8564
rect 22904 8536 22942 8564
rect 22976 8536 23014 8564
rect 23048 8536 23086 8564
rect 23120 8536 23158 8564
rect 23192 8536 23230 8564
rect 23264 8536 23302 8564
rect 23336 8536 23374 8564
rect 23408 8536 23446 8564
rect 23480 8536 23600 8564
rect 22852 8530 22870 8536
rect 22920 8530 22942 8536
rect 22988 8530 23014 8536
rect 23056 8530 23086 8536
rect 22766 8502 22818 8530
rect 22852 8502 22886 8530
rect 22920 8502 22954 8530
rect 22988 8502 23022 8530
rect 23056 8502 23090 8530
rect 23124 8502 23158 8536
rect 23192 8502 23226 8536
rect 23264 8530 23294 8536
rect 23336 8530 23362 8536
rect 23408 8530 23430 8536
rect 23480 8530 23498 8536
rect 23260 8502 23294 8530
rect 23328 8502 23362 8530
rect 23396 8502 23430 8530
rect 23464 8502 23498 8530
rect 23532 8502 23566 8536
rect 22766 8491 23600 8502
rect 22766 8457 22798 8491
rect 22832 8467 22870 8491
rect 22904 8467 22942 8491
rect 22976 8467 23014 8491
rect 23048 8467 23086 8491
rect 23120 8467 23158 8491
rect 23192 8467 23230 8491
rect 23264 8467 23302 8491
rect 23336 8467 23374 8491
rect 23408 8467 23446 8491
rect 23480 8467 23600 8491
rect 22852 8457 22870 8467
rect 22920 8457 22942 8467
rect 22988 8457 23014 8467
rect 23056 8457 23086 8467
rect 22766 8433 22818 8457
rect 22852 8433 22886 8457
rect 22920 8433 22954 8457
rect 22988 8433 23022 8457
rect 23056 8433 23090 8457
rect 23124 8433 23158 8467
rect 23192 8433 23226 8467
rect 23264 8457 23294 8467
rect 23336 8457 23362 8467
rect 23408 8457 23430 8467
rect 23480 8457 23498 8467
rect 23260 8433 23294 8457
rect 23328 8433 23362 8457
rect 23396 8433 23430 8457
rect 23464 8433 23498 8457
rect 23532 8433 23566 8467
rect 22766 8418 23600 8433
rect 22766 8384 22798 8418
rect 22832 8398 22870 8418
rect 22904 8398 22942 8418
rect 22976 8398 23014 8418
rect 23048 8398 23086 8418
rect 23120 8398 23158 8418
rect 23192 8398 23230 8418
rect 23264 8398 23302 8418
rect 23336 8398 23374 8418
rect 23408 8398 23446 8418
rect 23480 8398 23600 8418
rect 22852 8384 22870 8398
rect 22920 8384 22942 8398
rect 22988 8384 23014 8398
rect 23056 8384 23086 8398
rect 22766 8364 22818 8384
rect 22852 8364 22886 8384
rect 22920 8364 22954 8384
rect 22988 8364 23022 8384
rect 23056 8364 23090 8384
rect 23124 8364 23158 8398
rect 23192 8364 23226 8398
rect 23264 8384 23294 8398
rect 23336 8384 23362 8398
rect 23408 8384 23430 8398
rect 23480 8384 23498 8398
rect 23260 8364 23294 8384
rect 23328 8364 23362 8384
rect 23396 8364 23430 8384
rect 23464 8364 23498 8384
rect 23532 8364 23566 8398
rect 22766 8345 23600 8364
rect 22766 8311 22798 8345
rect 22832 8329 22870 8345
rect 22904 8329 22942 8345
rect 22976 8329 23014 8345
rect 23048 8329 23086 8345
rect 23120 8329 23158 8345
rect 23192 8329 23230 8345
rect 23264 8329 23302 8345
rect 23336 8329 23374 8345
rect 23408 8329 23446 8345
rect 23480 8329 23600 8345
rect 22852 8311 22870 8329
rect 22920 8311 22942 8329
rect 22988 8311 23014 8329
rect 23056 8311 23086 8329
rect 22766 8295 22818 8311
rect 22852 8295 22886 8311
rect 22920 8295 22954 8311
rect 22988 8295 23022 8311
rect 23056 8295 23090 8311
rect 23124 8295 23158 8329
rect 23192 8295 23226 8329
rect 23264 8311 23294 8329
rect 23336 8311 23362 8329
rect 23408 8311 23430 8329
rect 23480 8311 23498 8329
rect 23260 8295 23294 8311
rect 23328 8295 23362 8311
rect 23396 8295 23430 8311
rect 23464 8295 23498 8311
rect 23532 8295 23566 8329
rect 22766 8272 23600 8295
rect 22766 8238 22798 8272
rect 22832 8260 22870 8272
rect 22904 8260 22942 8272
rect 22976 8260 23014 8272
rect 23048 8260 23086 8272
rect 23120 8260 23158 8272
rect 23192 8260 23230 8272
rect 23264 8260 23302 8272
rect 23336 8260 23374 8272
rect 23408 8260 23446 8272
rect 23480 8260 23600 8272
rect 22852 8238 22870 8260
rect 22920 8238 22942 8260
rect 22988 8238 23014 8260
rect 23056 8238 23086 8260
rect 22766 8226 22818 8238
rect 22852 8226 22886 8238
rect 22920 8226 22954 8238
rect 22988 8226 23022 8238
rect 23056 8226 23090 8238
rect 23124 8226 23158 8260
rect 23192 8226 23226 8260
rect 23264 8238 23294 8260
rect 23336 8238 23362 8260
rect 23408 8238 23430 8260
rect 23480 8238 23498 8260
rect 23260 8226 23294 8238
rect 23328 8226 23362 8238
rect 23396 8226 23430 8238
rect 23464 8226 23498 8238
rect 23532 8226 23566 8260
rect 22766 8199 23600 8226
rect 22766 8165 22798 8199
rect 22832 8191 22870 8199
rect 22904 8191 22942 8199
rect 22976 8191 23014 8199
rect 23048 8191 23086 8199
rect 23120 8191 23158 8199
rect 23192 8191 23230 8199
rect 23264 8191 23302 8199
rect 23336 8191 23374 8199
rect 23408 8191 23446 8199
rect 23480 8191 23600 8199
rect 22852 8165 22870 8191
rect 22920 8165 22942 8191
rect 22988 8165 23014 8191
rect 23056 8165 23086 8191
rect 22766 8157 22818 8165
rect 22852 8157 22886 8165
rect 22920 8157 22954 8165
rect 22988 8157 23022 8165
rect 23056 8157 23090 8165
rect 23124 8157 23158 8191
rect 23192 8157 23226 8191
rect 23264 8165 23294 8191
rect 23336 8165 23362 8191
rect 23408 8165 23430 8191
rect 23480 8165 23498 8191
rect 23260 8157 23294 8165
rect 23328 8157 23362 8165
rect 23396 8157 23430 8165
rect 23464 8157 23498 8165
rect 23532 8157 23566 8191
rect 22766 8126 23600 8157
rect 22766 8092 22798 8126
rect 22832 8122 22870 8126
rect 22904 8122 22942 8126
rect 22976 8122 23014 8126
rect 23048 8122 23086 8126
rect 23120 8122 23158 8126
rect 23192 8122 23230 8126
rect 23264 8122 23302 8126
rect 23336 8122 23374 8126
rect 23408 8122 23446 8126
rect 23480 8122 23600 8126
rect 22852 8092 22870 8122
rect 22920 8092 22942 8122
rect 22988 8092 23014 8122
rect 23056 8092 23086 8122
rect 22766 8088 22818 8092
rect 22852 8088 22886 8092
rect 22920 8088 22954 8092
rect 22988 8088 23022 8092
rect 23056 8088 23090 8092
rect 23124 8088 23158 8122
rect 23192 8088 23226 8122
rect 23264 8092 23294 8122
rect 23336 8092 23362 8122
rect 23408 8092 23430 8122
rect 23480 8092 23498 8122
rect 23260 8088 23294 8092
rect 23328 8088 23362 8092
rect 23396 8088 23430 8092
rect 23464 8088 23498 8092
rect 23532 8088 23566 8122
rect 22766 8053 23600 8088
rect 22766 8019 22798 8053
rect 22852 8019 22870 8053
rect 22920 8019 22942 8053
rect 22988 8019 23014 8053
rect 23056 8019 23086 8053
rect 23124 8019 23158 8053
rect 23192 8019 23226 8053
rect 23264 8019 23294 8053
rect 23336 8019 23362 8053
rect 23408 8019 23430 8053
rect 23480 8019 23498 8053
rect 23532 8019 23566 8053
rect 22766 7984 23600 8019
rect 22766 7980 22818 7984
rect 22852 7980 22886 7984
rect 22920 7980 22954 7984
rect 22988 7980 23022 7984
rect 23056 7980 23090 7984
rect 22766 7946 22798 7980
rect 22852 7950 22870 7980
rect 22920 7950 22942 7980
rect 22988 7950 23014 7980
rect 23056 7950 23086 7980
rect 23124 7950 23158 7984
rect 23192 7950 23226 7984
rect 23260 7980 23294 7984
rect 23328 7980 23362 7984
rect 23396 7980 23430 7984
rect 23464 7980 23498 7984
rect 23264 7950 23294 7980
rect 23336 7950 23362 7980
rect 23408 7950 23430 7980
rect 23480 7950 23498 7980
rect 23532 7950 23566 7984
rect 22832 7946 22870 7950
rect 22904 7946 22942 7950
rect 22976 7946 23014 7950
rect 23048 7946 23086 7950
rect 23120 7946 23158 7950
rect 23192 7946 23230 7950
rect 23264 7946 23302 7950
rect 23336 7946 23374 7950
rect 23408 7946 23446 7950
rect 23480 7946 23600 7950
rect 22766 7915 23600 7946
rect 22766 7907 22818 7915
rect 22852 7907 22886 7915
rect 22920 7907 22954 7915
rect 22988 7907 23022 7915
rect 23056 7907 23090 7915
rect 22766 7873 22798 7907
rect 22852 7881 22870 7907
rect 22920 7881 22942 7907
rect 22988 7881 23014 7907
rect 23056 7881 23086 7907
rect 23124 7881 23158 7915
rect 23192 7881 23226 7915
rect 23260 7907 23294 7915
rect 23328 7907 23362 7915
rect 23396 7907 23430 7915
rect 23464 7907 23498 7915
rect 23264 7881 23294 7907
rect 23336 7881 23362 7907
rect 23408 7881 23430 7907
rect 23480 7881 23498 7907
rect 23532 7881 23566 7915
rect 22832 7873 22870 7881
rect 22904 7873 22942 7881
rect 22976 7873 23014 7881
rect 23048 7873 23086 7881
rect 23120 7873 23158 7881
rect 23192 7873 23230 7881
rect 23264 7873 23302 7881
rect 23336 7873 23374 7881
rect 23408 7873 23446 7881
rect 23480 7873 23600 7881
rect 22766 7846 23600 7873
rect 22766 7834 22818 7846
rect 22852 7834 22886 7846
rect 22920 7834 22954 7846
rect 22988 7834 23022 7846
rect 23056 7834 23090 7846
rect 22766 7800 22798 7834
rect 22852 7812 22870 7834
rect 22920 7812 22942 7834
rect 22988 7812 23014 7834
rect 23056 7812 23086 7834
rect 23124 7812 23158 7846
rect 23192 7812 23226 7846
rect 23260 7834 23294 7846
rect 23328 7834 23362 7846
rect 23396 7834 23430 7846
rect 23464 7834 23498 7846
rect 23264 7812 23294 7834
rect 23336 7812 23362 7834
rect 23408 7812 23430 7834
rect 23480 7812 23498 7834
rect 23532 7812 23566 7846
rect 22832 7800 22870 7812
rect 22904 7800 22942 7812
rect 22976 7800 23014 7812
rect 23048 7800 23086 7812
rect 23120 7800 23158 7812
rect 23192 7800 23230 7812
rect 23264 7800 23302 7812
rect 23336 7800 23374 7812
rect 23408 7800 23446 7812
rect 23480 7800 23600 7812
rect 22766 7777 23600 7800
rect 22766 7761 22818 7777
rect 22852 7761 22886 7777
rect 22920 7761 22954 7777
rect 22988 7761 23022 7777
rect 23056 7761 23090 7777
rect 22766 7727 22798 7761
rect 22852 7743 22870 7761
rect 22920 7743 22942 7761
rect 22988 7743 23014 7761
rect 23056 7743 23086 7761
rect 23124 7743 23158 7777
rect 23192 7743 23226 7777
rect 23260 7761 23294 7777
rect 23328 7761 23362 7777
rect 23396 7761 23430 7777
rect 23464 7761 23498 7777
rect 23264 7743 23294 7761
rect 23336 7743 23362 7761
rect 23408 7743 23430 7761
rect 23480 7743 23498 7761
rect 23532 7743 23566 7777
rect 22832 7727 22870 7743
rect 22904 7727 22942 7743
rect 22976 7727 23014 7743
rect 23048 7727 23086 7743
rect 23120 7727 23158 7743
rect 23192 7727 23230 7743
rect 23264 7727 23302 7743
rect 23336 7727 23374 7743
rect 23408 7727 23446 7743
rect 23480 7727 23600 7743
rect 22766 7708 23600 7727
rect 22766 7688 22818 7708
rect 22852 7688 22886 7708
rect 22920 7688 22954 7708
rect 22988 7688 23022 7708
rect 23056 7688 23090 7708
rect 22766 7654 22798 7688
rect 22852 7674 22870 7688
rect 22920 7674 22942 7688
rect 22988 7674 23014 7688
rect 23056 7674 23086 7688
rect 23124 7674 23158 7708
rect 23192 7674 23226 7708
rect 23260 7688 23294 7708
rect 23328 7688 23362 7708
rect 23396 7688 23430 7708
rect 23464 7688 23498 7708
rect 23264 7674 23294 7688
rect 23336 7674 23362 7688
rect 23408 7674 23430 7688
rect 23480 7674 23498 7688
rect 23532 7674 23566 7708
rect 22832 7654 22870 7674
rect 22904 7654 22942 7674
rect 22976 7654 23014 7674
rect 23048 7654 23086 7674
rect 23120 7654 23158 7674
rect 23192 7654 23230 7674
rect 23264 7654 23302 7674
rect 23336 7654 23374 7674
rect 23408 7654 23446 7674
rect 23480 7654 23600 7674
rect 22766 7639 23600 7654
rect 22766 7615 22818 7639
rect 22852 7615 22886 7639
rect 22920 7615 22954 7639
rect 22988 7615 23022 7639
rect 23056 7615 23090 7639
rect 22766 7581 22798 7615
rect 22852 7605 22870 7615
rect 22920 7605 22942 7615
rect 22988 7605 23014 7615
rect 23056 7605 23086 7615
rect 23124 7605 23158 7639
rect 23192 7605 23226 7639
rect 23260 7615 23294 7639
rect 23328 7615 23362 7639
rect 23396 7615 23430 7639
rect 23464 7615 23498 7639
rect 23264 7605 23294 7615
rect 23336 7605 23362 7615
rect 23408 7605 23430 7615
rect 23480 7605 23498 7615
rect 23532 7605 23566 7639
rect 22832 7581 22870 7605
rect 22904 7581 22942 7605
rect 22976 7581 23014 7605
rect 23048 7581 23086 7605
rect 23120 7581 23158 7605
rect 23192 7581 23230 7605
rect 23264 7581 23302 7605
rect 23336 7581 23374 7605
rect 23408 7581 23446 7605
rect 23480 7581 23600 7605
rect 22766 7570 23600 7581
rect 22766 7542 22818 7570
rect 22852 7542 22886 7570
rect 22920 7542 22954 7570
rect 22988 7542 23022 7570
rect 23056 7542 23090 7570
rect 22766 7508 22798 7542
rect 22852 7536 22870 7542
rect 22920 7536 22942 7542
rect 22988 7536 23014 7542
rect 23056 7536 23086 7542
rect 23124 7536 23158 7570
rect 23192 7536 23226 7570
rect 23260 7542 23294 7570
rect 23328 7542 23362 7570
rect 23396 7542 23430 7570
rect 23464 7542 23498 7570
rect 23264 7536 23294 7542
rect 23336 7536 23362 7542
rect 23408 7536 23430 7542
rect 23480 7536 23498 7542
rect 23532 7536 23566 7570
rect 22832 7508 22870 7536
rect 22904 7508 22942 7536
rect 22976 7508 23014 7536
rect 23048 7508 23086 7536
rect 23120 7508 23158 7536
rect 23192 7508 23230 7536
rect 23264 7508 23302 7536
rect 23336 7508 23374 7536
rect 23408 7508 23446 7536
rect 23480 7508 23600 7536
rect 22766 7501 23600 7508
rect 22766 7469 22818 7501
rect 22852 7469 22886 7501
rect 22920 7469 22954 7501
rect 22988 7469 23022 7501
rect 23056 7469 23090 7501
rect 22766 7435 22798 7469
rect 22852 7467 22870 7469
rect 22920 7467 22942 7469
rect 22988 7467 23014 7469
rect 23056 7467 23086 7469
rect 23124 7467 23158 7501
rect 23192 7467 23226 7501
rect 23260 7469 23294 7501
rect 23328 7469 23362 7501
rect 23396 7469 23430 7501
rect 23464 7469 23498 7501
rect 23264 7467 23294 7469
rect 23336 7467 23362 7469
rect 23408 7467 23430 7469
rect 23480 7467 23498 7469
rect 23532 7467 23566 7501
rect 22832 7435 22870 7467
rect 22904 7435 22942 7467
rect 22976 7435 23014 7467
rect 23048 7435 23086 7467
rect 23120 7435 23158 7467
rect 23192 7435 23230 7467
rect 23264 7435 23302 7467
rect 23336 7435 23374 7467
rect 23408 7435 23446 7467
rect 23480 7435 23600 7467
rect 22766 7432 23600 7435
rect 22766 7398 22818 7432
rect 22852 7398 22886 7432
rect 22920 7398 22954 7432
rect 22988 7398 23022 7432
rect 23056 7398 23090 7432
rect 23124 7398 23158 7432
rect 23192 7398 23226 7432
rect 23260 7398 23294 7432
rect 23328 7398 23362 7432
rect 23396 7398 23430 7432
rect 23464 7398 23498 7432
rect 23532 7398 23566 7432
rect 22766 7396 23600 7398
rect 22766 7362 22798 7396
rect 22832 7363 22870 7396
rect 22904 7363 22942 7396
rect 22976 7363 23014 7396
rect 23048 7363 23086 7396
rect 23120 7363 23158 7396
rect 23192 7363 23230 7396
rect 23264 7363 23302 7396
rect 23336 7363 23374 7396
rect 23408 7363 23446 7396
rect 23480 7363 23600 7396
rect 22852 7362 22870 7363
rect 22920 7362 22942 7363
rect 22988 7362 23014 7363
rect 23056 7362 23086 7363
rect 22766 7329 22818 7362
rect 22852 7329 22886 7362
rect 22920 7329 22954 7362
rect 22988 7329 23022 7362
rect 23056 7329 23090 7362
rect 23124 7329 23158 7363
rect 23192 7329 23226 7363
rect 23264 7362 23294 7363
rect 23336 7362 23362 7363
rect 23408 7362 23430 7363
rect 23480 7362 23498 7363
rect 23260 7329 23294 7362
rect 23328 7329 23362 7362
rect 23396 7329 23430 7362
rect 23464 7329 23498 7362
rect 23532 7329 23566 7363
rect 22766 7323 23600 7329
rect 22766 7289 22798 7323
rect 22832 7294 22870 7323
rect 22904 7294 22942 7323
rect 22976 7294 23014 7323
rect 23048 7294 23086 7323
rect 23120 7294 23158 7323
rect 23192 7294 23230 7323
rect 23264 7294 23302 7323
rect 23336 7294 23374 7323
rect 23408 7294 23446 7323
rect 23480 7294 23600 7323
rect 22852 7289 22870 7294
rect 22920 7289 22942 7294
rect 22988 7289 23014 7294
rect 23056 7289 23086 7294
rect 22766 7260 22818 7289
rect 22852 7260 22886 7289
rect 22920 7260 22954 7289
rect 22988 7260 23022 7289
rect 23056 7260 23090 7289
rect 23124 7260 23158 7294
rect 23192 7260 23226 7294
rect 23264 7289 23294 7294
rect 23336 7289 23362 7294
rect 23408 7289 23430 7294
rect 23480 7289 23498 7294
rect 23260 7260 23294 7289
rect 23328 7260 23362 7289
rect 23396 7260 23430 7289
rect 23464 7260 23498 7289
rect 23532 7260 23566 7294
rect 22766 7250 23600 7260
rect 22766 7216 22798 7250
rect 22832 7225 22870 7250
rect 22904 7225 22942 7250
rect 22976 7225 23014 7250
rect 23048 7225 23086 7250
rect 23120 7225 23158 7250
rect 23192 7225 23230 7250
rect 23264 7225 23302 7250
rect 23336 7225 23374 7250
rect 23408 7225 23446 7250
rect 23480 7225 23600 7250
rect 22852 7216 22870 7225
rect 22920 7216 22942 7225
rect 22988 7216 23014 7225
rect 23056 7216 23086 7225
rect 22766 7191 22818 7216
rect 22852 7191 22886 7216
rect 22920 7191 22954 7216
rect 22988 7191 23022 7216
rect 23056 7191 23090 7216
rect 23124 7191 23158 7225
rect 23192 7191 23226 7225
rect 23264 7216 23294 7225
rect 23336 7216 23362 7225
rect 23408 7216 23430 7225
rect 23480 7216 23498 7225
rect 23260 7191 23294 7216
rect 23328 7191 23362 7216
rect 23396 7191 23430 7216
rect 23464 7191 23498 7216
rect 23532 7191 23566 7225
rect 22766 7177 23600 7191
rect 22766 7143 22798 7177
rect 22832 7156 22870 7177
rect 22904 7156 22942 7177
rect 22976 7156 23014 7177
rect 23048 7156 23086 7177
rect 23120 7156 23158 7177
rect 23192 7156 23230 7177
rect 23264 7156 23302 7177
rect 23336 7156 23374 7177
rect 23408 7156 23446 7177
rect 23480 7156 23600 7177
rect 22852 7143 22870 7156
rect 22920 7143 22942 7156
rect 22988 7143 23014 7156
rect 23056 7143 23086 7156
rect 22766 7122 22818 7143
rect 22852 7122 22886 7143
rect 22920 7122 22954 7143
rect 22988 7122 23022 7143
rect 23056 7122 23090 7143
rect 23124 7122 23158 7156
rect 23192 7122 23226 7156
rect 23264 7143 23294 7156
rect 23336 7143 23362 7156
rect 23408 7143 23430 7156
rect 23480 7143 23498 7156
rect 23260 7122 23294 7143
rect 23328 7122 23362 7143
rect 23396 7122 23430 7143
rect 23464 7122 23498 7143
rect 23532 7122 23566 7156
rect 22766 7104 23600 7122
rect 22766 7070 22798 7104
rect 22832 7087 22870 7104
rect 22904 7087 22942 7104
rect 22976 7087 23014 7104
rect 23048 7087 23086 7104
rect 23120 7087 23158 7104
rect 23192 7087 23230 7104
rect 23264 7087 23302 7104
rect 23336 7087 23374 7104
rect 23408 7087 23446 7104
rect 23480 7087 23600 7104
rect 22852 7070 22870 7087
rect 22920 7070 22942 7087
rect 22988 7070 23014 7087
rect 23056 7070 23086 7087
rect 22766 7053 22818 7070
rect 22852 7053 22886 7070
rect 22920 7053 22954 7070
rect 22988 7053 23022 7070
rect 23056 7053 23090 7070
rect 23124 7053 23158 7087
rect 23192 7053 23226 7087
rect 23264 7070 23294 7087
rect 23336 7070 23362 7087
rect 23408 7070 23430 7087
rect 23480 7070 23498 7087
rect 23260 7053 23294 7070
rect 23328 7053 23362 7070
rect 23396 7053 23430 7070
rect 23464 7053 23498 7070
rect 23532 7053 23566 7087
rect 22766 7031 23600 7053
rect 22766 6997 22798 7031
rect 22832 7018 22870 7031
rect 22904 7018 22942 7031
rect 22976 7018 23014 7031
rect 23048 7018 23086 7031
rect 23120 7018 23158 7031
rect 23192 7018 23230 7031
rect 23264 7018 23302 7031
rect 23336 7018 23374 7031
rect 23408 7018 23446 7031
rect 23480 7018 23600 7031
rect 22852 6997 22870 7018
rect 22920 6997 22942 7018
rect 22988 6997 23014 7018
rect 23056 6997 23086 7018
rect 22766 6984 22818 6997
rect 22852 6984 22886 6997
rect 22920 6984 22954 6997
rect 22988 6984 23022 6997
rect 23056 6984 23090 6997
rect 23124 6984 23158 7018
rect 23192 6984 23226 7018
rect 23264 6997 23294 7018
rect 23336 6997 23362 7018
rect 23408 6997 23430 7018
rect 23480 6997 23498 7018
rect 23260 6984 23294 6997
rect 23328 6984 23362 6997
rect 23396 6984 23430 6997
rect 23464 6984 23498 6997
rect 23532 6984 23566 7018
rect 22766 6958 23600 6984
rect 22766 6924 22798 6958
rect 22832 6949 22870 6958
rect 22904 6949 22942 6958
rect 22976 6949 23014 6958
rect 23048 6949 23086 6958
rect 23120 6949 23158 6958
rect 23192 6949 23230 6958
rect 23264 6949 23302 6958
rect 23336 6949 23374 6958
rect 23408 6949 23446 6958
rect 23480 6949 23600 6958
rect 22852 6924 22870 6949
rect 22920 6924 22942 6949
rect 22988 6924 23014 6949
rect 23056 6924 23086 6949
rect 22766 6915 22818 6924
rect 22852 6915 22886 6924
rect 22920 6915 22954 6924
rect 22988 6915 23022 6924
rect 23056 6915 23090 6924
rect 23124 6915 23158 6949
rect 23192 6915 23226 6949
rect 23264 6924 23294 6949
rect 23336 6924 23362 6949
rect 23408 6924 23430 6949
rect 23480 6924 23498 6949
rect 23260 6915 23294 6924
rect 23328 6915 23362 6924
rect 23396 6915 23430 6924
rect 23464 6915 23498 6924
rect 23532 6915 23566 6949
rect 22766 6885 23600 6915
rect 22766 6851 22798 6885
rect 22832 6880 22870 6885
rect 22904 6880 22942 6885
rect 22976 6880 23014 6885
rect 23048 6880 23086 6885
rect 23120 6880 23158 6885
rect 23192 6880 23230 6885
rect 23264 6880 23302 6885
rect 23336 6880 23374 6885
rect 23408 6880 23446 6885
rect 23480 6880 23600 6885
rect 22852 6851 22870 6880
rect 22920 6851 22942 6880
rect 22988 6851 23014 6880
rect 23056 6851 23086 6880
rect 22766 6846 22818 6851
rect 22852 6846 22886 6851
rect 22920 6846 22954 6851
rect 22988 6846 23022 6851
rect 23056 6846 23090 6851
rect 23124 6846 23158 6880
rect 23192 6846 23226 6880
rect 23264 6851 23294 6880
rect 23336 6851 23362 6880
rect 23408 6851 23430 6880
rect 23480 6851 23498 6880
rect 23260 6846 23294 6851
rect 23328 6846 23362 6851
rect 23396 6846 23430 6851
rect 23464 6846 23498 6851
rect 23532 6846 23566 6880
rect 22766 6812 23600 6846
rect 22766 6778 22798 6812
rect 22832 6811 22870 6812
rect 22904 6811 22942 6812
rect 22976 6811 23014 6812
rect 23048 6811 23086 6812
rect 23120 6811 23158 6812
rect 23192 6811 23230 6812
rect 23264 6811 23302 6812
rect 23336 6811 23374 6812
rect 23408 6811 23446 6812
rect 23480 6811 23600 6812
rect 22766 6739 22818 6778
rect 22766 6705 22798 6739
rect 22766 6666 22818 6705
rect 22766 6632 22798 6666
rect 22766 6593 22818 6632
rect 22766 6559 22798 6593
rect 22766 6520 22818 6559
rect 22766 6486 22798 6520
rect 22766 6447 22818 6486
rect 22766 6413 22798 6447
rect 22766 6374 22818 6413
rect 22766 6340 22798 6374
rect 22766 6301 22818 6340
rect 22766 6267 22798 6301
rect 22766 6228 22818 6267
rect 22766 6194 22798 6228
rect 22766 6155 22818 6194
rect 22766 6121 22798 6155
rect 22766 6082 22818 6121
rect 22766 6048 22798 6082
rect 22766 6009 22818 6048
rect 22766 5975 22798 6009
rect 22766 5936 22818 5975
rect 22766 5902 22798 5936
rect 22766 5863 22818 5902
rect 22766 5829 22798 5863
rect 22766 5790 22818 5829
rect 22766 5756 22798 5790
rect 22766 5717 22818 5756
rect 22766 5683 22798 5717
rect 22766 5644 22818 5683
rect 22766 5610 22798 5644
rect 23752 8568 23781 8592
rect 23752 8534 23755 8568
rect 24537 8534 24540 8602
rect 23752 8499 23781 8534
rect 24535 8499 24540 8534
rect 23752 8465 23755 8499
rect 24537 8465 24540 8499
rect 23752 8430 23781 8465
rect 24535 8430 24540 8465
rect 23752 8396 23755 8430
rect 24537 8396 24540 8430
rect 23752 8361 23781 8396
rect 24535 8361 24540 8396
rect 23752 8327 23755 8361
rect 24537 8327 24540 8361
rect 23752 8292 23781 8327
rect 24535 8292 24540 8327
rect 23752 8258 23755 8292
rect 24537 8258 24540 8292
rect 23752 8223 23781 8258
rect 24535 8223 24540 8258
rect 23752 8189 23755 8223
rect 24537 8189 24540 8223
rect 23752 8154 23781 8189
rect 24535 8154 24540 8189
rect 23752 8120 23755 8154
rect 24537 8120 24540 8154
rect 23752 8085 23781 8120
rect 24535 8085 24540 8120
rect 23752 8051 23755 8085
rect 24537 8051 24540 8085
rect 23752 8016 23781 8051
rect 24535 8016 24540 8051
rect 23752 7982 23755 8016
rect 24537 7982 24540 8016
rect 23752 7947 23781 7982
rect 24535 7947 24540 7982
rect 23752 7913 23755 7947
rect 24537 7913 24540 7947
rect 23752 7878 23781 7913
rect 24535 7878 24540 7913
rect 23752 7844 23755 7878
rect 23789 7844 23823 7854
rect 23857 7844 23891 7854
rect 23925 7844 23959 7854
rect 23993 7844 24027 7854
rect 24061 7844 24095 7854
rect 24129 7844 24163 7854
rect 24197 7844 24231 7854
rect 24265 7844 24299 7854
rect 24333 7844 24367 7854
rect 24401 7844 24435 7854
rect 24469 7844 24503 7854
rect 24537 7844 24540 7878
rect 23752 7815 24540 7844
rect 23752 7809 23781 7815
rect 23815 7809 23853 7815
rect 23887 7809 23925 7815
rect 23752 7775 23755 7809
rect 23815 7781 23823 7809
rect 23887 7781 23891 7809
rect 23789 7775 23823 7781
rect 23857 7775 23891 7781
rect 23959 7809 23997 7815
rect 24031 7809 24069 7815
rect 24103 7809 24141 7815
rect 24175 7809 24213 7815
rect 24247 7809 24285 7815
rect 24319 7809 24357 7815
rect 24391 7809 24429 7815
rect 24463 7809 24501 7815
rect 24535 7809 24540 7815
rect 23925 7775 23959 7781
rect 23993 7781 23997 7809
rect 24061 7781 24069 7809
rect 24129 7781 24141 7809
rect 24197 7781 24213 7809
rect 24265 7781 24285 7809
rect 24333 7781 24357 7809
rect 24401 7781 24429 7809
rect 24469 7781 24501 7809
rect 23993 7775 24027 7781
rect 24061 7775 24095 7781
rect 24129 7775 24163 7781
rect 24197 7775 24231 7781
rect 24265 7775 24299 7781
rect 24333 7775 24367 7781
rect 24401 7775 24435 7781
rect 24469 7775 24503 7781
rect 24537 7775 24540 7809
rect 23752 7742 24540 7775
rect 23752 7740 23781 7742
rect 23815 7740 23853 7742
rect 23887 7740 23925 7742
rect 23752 7706 23755 7740
rect 23815 7708 23823 7740
rect 23887 7708 23891 7740
rect 23789 7706 23823 7708
rect 23857 7706 23891 7708
rect 23959 7740 23997 7742
rect 24031 7740 24069 7742
rect 24103 7740 24141 7742
rect 24175 7740 24213 7742
rect 24247 7740 24285 7742
rect 24319 7740 24357 7742
rect 24391 7740 24429 7742
rect 24463 7740 24501 7742
rect 24535 7740 24540 7742
rect 23925 7706 23959 7708
rect 23993 7708 23997 7740
rect 24061 7708 24069 7740
rect 24129 7708 24141 7740
rect 24197 7708 24213 7740
rect 24265 7708 24285 7740
rect 24333 7708 24357 7740
rect 24401 7708 24429 7740
rect 24469 7708 24501 7740
rect 23993 7706 24027 7708
rect 24061 7706 24095 7708
rect 24129 7706 24163 7708
rect 24197 7706 24231 7708
rect 24265 7706 24299 7708
rect 24333 7706 24367 7708
rect 24401 7706 24435 7708
rect 24469 7706 24503 7708
rect 24537 7706 24540 7740
rect 23752 7671 24540 7706
rect 23752 7637 23755 7671
rect 23789 7669 23823 7671
rect 23857 7669 23891 7671
rect 23815 7637 23823 7669
rect 23887 7637 23891 7669
rect 23925 7669 23959 7671
rect 23752 7635 23781 7637
rect 23815 7635 23853 7637
rect 23887 7635 23925 7637
rect 23993 7669 24027 7671
rect 24061 7669 24095 7671
rect 24129 7669 24163 7671
rect 24197 7669 24231 7671
rect 24265 7669 24299 7671
rect 24333 7669 24367 7671
rect 24401 7669 24435 7671
rect 24469 7669 24503 7671
rect 23993 7637 23997 7669
rect 24061 7637 24069 7669
rect 24129 7637 24141 7669
rect 24197 7637 24213 7669
rect 24265 7637 24285 7669
rect 24333 7637 24357 7669
rect 24401 7637 24429 7669
rect 24469 7637 24501 7669
rect 24537 7637 24540 7671
rect 23959 7635 23997 7637
rect 24031 7635 24069 7637
rect 24103 7635 24141 7637
rect 24175 7635 24213 7637
rect 24247 7635 24285 7637
rect 24319 7635 24357 7637
rect 24391 7635 24429 7637
rect 24463 7635 24501 7637
rect 24535 7635 24540 7637
rect 23752 7602 24540 7635
rect 23752 7568 23755 7602
rect 23789 7596 23823 7602
rect 23857 7596 23891 7602
rect 23815 7568 23823 7596
rect 23887 7568 23891 7596
rect 23925 7596 23959 7602
rect 23752 7562 23781 7568
rect 23815 7562 23853 7568
rect 23887 7562 23925 7568
rect 23993 7596 24027 7602
rect 24061 7596 24095 7602
rect 24129 7596 24163 7602
rect 24197 7596 24231 7602
rect 24265 7596 24299 7602
rect 24333 7596 24367 7602
rect 24401 7596 24435 7602
rect 24469 7596 24503 7602
rect 23993 7568 23997 7596
rect 24061 7568 24069 7596
rect 24129 7568 24141 7596
rect 24197 7568 24213 7596
rect 24265 7568 24285 7596
rect 24333 7568 24357 7596
rect 24401 7568 24429 7596
rect 24469 7568 24501 7596
rect 24537 7568 24540 7602
rect 23959 7562 23997 7568
rect 24031 7562 24069 7568
rect 24103 7562 24141 7568
rect 24175 7562 24213 7568
rect 24247 7562 24285 7568
rect 24319 7562 24357 7568
rect 24391 7562 24429 7568
rect 24463 7562 24501 7568
rect 24535 7562 24540 7568
rect 23752 7533 24540 7562
rect 23752 7499 23755 7533
rect 23789 7523 23823 7533
rect 23857 7523 23891 7533
rect 23815 7499 23823 7523
rect 23887 7499 23891 7523
rect 23925 7523 23959 7533
rect 23752 7489 23781 7499
rect 23815 7489 23853 7499
rect 23887 7489 23925 7499
rect 23993 7523 24027 7533
rect 24061 7523 24095 7533
rect 24129 7523 24163 7533
rect 24197 7523 24231 7533
rect 24265 7523 24299 7533
rect 24333 7523 24367 7533
rect 24401 7523 24435 7533
rect 24469 7523 24503 7533
rect 23993 7499 23997 7523
rect 24061 7499 24069 7523
rect 24129 7499 24141 7523
rect 24197 7499 24213 7523
rect 24265 7499 24285 7523
rect 24333 7499 24357 7523
rect 24401 7499 24429 7523
rect 24469 7499 24501 7523
rect 24537 7499 24540 7533
rect 23959 7489 23997 7499
rect 24031 7489 24069 7499
rect 24103 7489 24141 7499
rect 24175 7489 24213 7499
rect 24247 7489 24285 7499
rect 24319 7489 24357 7499
rect 24391 7489 24429 7499
rect 24463 7489 24501 7499
rect 24535 7489 24540 7499
rect 23752 7464 24540 7489
rect 23752 7430 23755 7464
rect 23789 7450 23823 7464
rect 23857 7450 23891 7464
rect 23815 7430 23823 7450
rect 23887 7430 23891 7450
rect 23925 7450 23959 7464
rect 23752 7416 23781 7430
rect 23815 7416 23853 7430
rect 23887 7416 23925 7430
rect 23993 7450 24027 7464
rect 24061 7450 24095 7464
rect 24129 7450 24163 7464
rect 24197 7450 24231 7464
rect 24265 7450 24299 7464
rect 24333 7450 24367 7464
rect 24401 7450 24435 7464
rect 24469 7450 24503 7464
rect 23993 7430 23997 7450
rect 24061 7430 24069 7450
rect 24129 7430 24141 7450
rect 24197 7430 24213 7450
rect 24265 7430 24285 7450
rect 24333 7430 24357 7450
rect 24401 7430 24429 7450
rect 24469 7430 24501 7450
rect 24537 7430 24540 7464
rect 23959 7416 23997 7430
rect 24031 7416 24069 7430
rect 24103 7416 24141 7430
rect 24175 7416 24213 7430
rect 24247 7416 24285 7430
rect 24319 7416 24357 7430
rect 24391 7416 24429 7430
rect 24463 7416 24501 7430
rect 24535 7416 24540 7430
rect 23752 7395 24540 7416
rect 23752 7361 23755 7395
rect 23789 7377 23823 7395
rect 23857 7377 23891 7395
rect 23815 7361 23823 7377
rect 23887 7361 23891 7377
rect 23925 7377 23959 7395
rect 23752 7343 23781 7361
rect 23815 7343 23853 7361
rect 23887 7343 23925 7361
rect 23993 7377 24027 7395
rect 24061 7377 24095 7395
rect 24129 7377 24163 7395
rect 24197 7377 24231 7395
rect 24265 7377 24299 7395
rect 24333 7377 24367 7395
rect 24401 7377 24435 7395
rect 24469 7377 24503 7395
rect 23993 7361 23997 7377
rect 24061 7361 24069 7377
rect 24129 7361 24141 7377
rect 24197 7361 24213 7377
rect 24265 7361 24285 7377
rect 24333 7361 24357 7377
rect 24401 7361 24429 7377
rect 24469 7361 24501 7377
rect 24537 7361 24540 7395
rect 23959 7343 23997 7361
rect 24031 7343 24069 7361
rect 24103 7343 24141 7361
rect 24175 7343 24213 7361
rect 24247 7343 24285 7361
rect 24319 7343 24357 7361
rect 24391 7343 24429 7361
rect 24463 7343 24501 7361
rect 24535 7343 24540 7361
rect 23752 7326 24540 7343
rect 23752 7292 23755 7326
rect 23789 7304 23823 7326
rect 23857 7304 23891 7326
rect 23815 7292 23823 7304
rect 23887 7292 23891 7304
rect 23925 7304 23959 7326
rect 23752 7270 23781 7292
rect 23815 7270 23853 7292
rect 23887 7270 23925 7292
rect 23993 7304 24027 7326
rect 24061 7304 24095 7326
rect 24129 7304 24163 7326
rect 24197 7304 24231 7326
rect 24265 7304 24299 7326
rect 24333 7304 24367 7326
rect 24401 7304 24435 7326
rect 24469 7304 24503 7326
rect 23993 7292 23997 7304
rect 24061 7292 24069 7304
rect 24129 7292 24141 7304
rect 24197 7292 24213 7304
rect 24265 7292 24285 7304
rect 24333 7292 24357 7304
rect 24401 7292 24429 7304
rect 24469 7292 24501 7304
rect 24537 7292 24540 7326
rect 23959 7270 23997 7292
rect 24031 7270 24069 7292
rect 24103 7270 24141 7292
rect 24175 7270 24213 7292
rect 24247 7270 24285 7292
rect 24319 7270 24357 7292
rect 24391 7270 24429 7292
rect 24463 7270 24501 7292
rect 24535 7270 24540 7292
rect 23752 7257 24540 7270
rect 23752 7223 23755 7257
rect 23789 7231 23823 7257
rect 23857 7231 23891 7257
rect 23815 7223 23823 7231
rect 23887 7223 23891 7231
rect 23925 7231 23959 7257
rect 23752 7197 23781 7223
rect 23815 7197 23853 7223
rect 23887 7197 23925 7223
rect 23993 7231 24027 7257
rect 24061 7231 24095 7257
rect 24129 7231 24163 7257
rect 24197 7231 24231 7257
rect 24265 7231 24299 7257
rect 24333 7231 24367 7257
rect 24401 7231 24435 7257
rect 24469 7231 24503 7257
rect 23993 7223 23997 7231
rect 24061 7223 24069 7231
rect 24129 7223 24141 7231
rect 24197 7223 24213 7231
rect 24265 7223 24285 7231
rect 24333 7223 24357 7231
rect 24401 7223 24429 7231
rect 24469 7223 24501 7231
rect 24537 7223 24540 7257
rect 23959 7197 23997 7223
rect 24031 7197 24069 7223
rect 24103 7197 24141 7223
rect 24175 7197 24213 7223
rect 24247 7197 24285 7223
rect 24319 7197 24357 7223
rect 24391 7197 24429 7223
rect 24463 7197 24501 7223
rect 24535 7197 24540 7223
rect 23752 7188 24540 7197
rect 23752 7154 23755 7188
rect 23789 7158 23823 7188
rect 23857 7158 23891 7188
rect 23815 7154 23823 7158
rect 23887 7154 23891 7158
rect 23925 7158 23959 7188
rect 23752 7124 23781 7154
rect 23815 7124 23853 7154
rect 23887 7124 23925 7154
rect 23993 7158 24027 7188
rect 24061 7158 24095 7188
rect 24129 7158 24163 7188
rect 24197 7158 24231 7188
rect 24265 7158 24299 7188
rect 24333 7158 24367 7188
rect 24401 7158 24435 7188
rect 24469 7158 24503 7188
rect 23993 7154 23997 7158
rect 24061 7154 24069 7158
rect 24129 7154 24141 7158
rect 24197 7154 24213 7158
rect 24265 7154 24285 7158
rect 24333 7154 24357 7158
rect 24401 7154 24429 7158
rect 24469 7154 24501 7158
rect 24537 7154 24540 7188
rect 23959 7124 23997 7154
rect 24031 7124 24069 7154
rect 24103 7124 24141 7154
rect 24175 7124 24213 7154
rect 24247 7124 24285 7154
rect 24319 7124 24357 7154
rect 24391 7124 24429 7154
rect 24463 7124 24501 7154
rect 24535 7124 24540 7154
rect 23752 7119 24540 7124
rect 23752 7085 23755 7119
rect 23789 7085 23823 7119
rect 23857 7085 23891 7119
rect 23925 7085 23959 7119
rect 23993 7085 24027 7119
rect 24061 7085 24095 7119
rect 24129 7085 24163 7119
rect 24197 7085 24231 7119
rect 24265 7085 24299 7119
rect 24333 7085 24367 7119
rect 24401 7085 24435 7119
rect 24469 7085 24503 7119
rect 24537 7085 24540 7119
rect 23752 7051 23781 7085
rect 23815 7051 23853 7085
rect 23887 7051 23925 7085
rect 23959 7051 23997 7085
rect 24031 7051 24069 7085
rect 24103 7051 24141 7085
rect 24175 7051 24213 7085
rect 24247 7051 24285 7085
rect 24319 7051 24357 7085
rect 24391 7051 24429 7085
rect 24463 7051 24501 7085
rect 24535 7051 24540 7085
rect 23752 7050 24540 7051
rect 23752 7016 23755 7050
rect 23789 7016 23823 7050
rect 23857 7016 23891 7050
rect 23925 7016 23959 7050
rect 23993 7016 24027 7050
rect 24061 7016 24095 7050
rect 24129 7016 24163 7050
rect 24197 7016 24231 7050
rect 24265 7016 24299 7050
rect 24333 7016 24367 7050
rect 24401 7016 24435 7050
rect 24469 7016 24503 7050
rect 24537 7016 24540 7050
rect 23752 7012 24540 7016
rect 23752 6981 23781 7012
rect 23815 6981 23853 7012
rect 23887 6981 23925 7012
rect 23752 6947 23755 6981
rect 23815 6978 23823 6981
rect 23887 6978 23891 6981
rect 23789 6947 23823 6978
rect 23857 6947 23891 6978
rect 23959 6981 23997 7012
rect 24031 6981 24069 7012
rect 24103 6981 24141 7012
rect 24175 6981 24213 7012
rect 24247 6981 24285 7012
rect 24319 6981 24357 7012
rect 24391 6981 24429 7012
rect 24463 6981 24501 7012
rect 24535 6981 24540 7012
rect 23925 6947 23959 6978
rect 23993 6978 23997 6981
rect 24061 6978 24069 6981
rect 24129 6978 24141 6981
rect 24197 6978 24213 6981
rect 24265 6978 24285 6981
rect 24333 6978 24357 6981
rect 24401 6978 24429 6981
rect 24469 6978 24501 6981
rect 23993 6947 24027 6978
rect 24061 6947 24095 6978
rect 24129 6947 24163 6978
rect 24197 6947 24231 6978
rect 24265 6947 24299 6978
rect 24333 6947 24367 6978
rect 24401 6947 24435 6978
rect 24469 6947 24503 6978
rect 24537 6947 24540 6981
rect 23752 6939 24540 6947
rect 23752 6912 23781 6939
rect 23815 6912 23853 6939
rect 23887 6912 23925 6939
rect 23752 6878 23755 6912
rect 23815 6905 23823 6912
rect 23887 6905 23891 6912
rect 23789 6878 23823 6905
rect 23857 6878 23891 6905
rect 23959 6912 23997 6939
rect 24031 6912 24069 6939
rect 24103 6912 24141 6939
rect 24175 6912 24213 6939
rect 24247 6912 24285 6939
rect 24319 6912 24357 6939
rect 24391 6912 24429 6939
rect 24463 6912 24501 6939
rect 24535 6912 24540 6939
rect 23925 6878 23959 6905
rect 23993 6905 23997 6912
rect 24061 6905 24069 6912
rect 24129 6905 24141 6912
rect 24197 6905 24213 6912
rect 24265 6905 24285 6912
rect 24333 6905 24357 6912
rect 24401 6905 24429 6912
rect 24469 6905 24501 6912
rect 23993 6878 24027 6905
rect 24061 6878 24095 6905
rect 24129 6878 24163 6905
rect 24197 6878 24231 6905
rect 24265 6878 24299 6905
rect 24333 6878 24367 6905
rect 24401 6878 24435 6905
rect 24469 6878 24503 6905
rect 24537 6878 24540 6912
rect 23752 6866 24540 6878
rect 23752 6843 23781 6866
rect 23815 6843 23853 6866
rect 23887 6843 23925 6866
rect 23752 6809 23755 6843
rect 23815 6832 23823 6843
rect 23887 6832 23891 6843
rect 23789 6809 23823 6832
rect 23857 6809 23891 6832
rect 23959 6843 23997 6866
rect 24031 6843 24069 6866
rect 24103 6843 24141 6866
rect 24175 6843 24213 6866
rect 24247 6843 24285 6866
rect 24319 6843 24357 6866
rect 24391 6843 24429 6866
rect 24463 6843 24501 6866
rect 24535 6843 24540 6866
rect 23925 6809 23959 6832
rect 23993 6832 23997 6843
rect 24061 6832 24069 6843
rect 24129 6832 24141 6843
rect 24197 6832 24213 6843
rect 24265 6832 24285 6843
rect 24333 6832 24357 6843
rect 24401 6832 24429 6843
rect 24469 6832 24501 6843
rect 23993 6809 24027 6832
rect 24061 6809 24095 6832
rect 24129 6809 24163 6832
rect 24197 6809 24231 6832
rect 24265 6809 24299 6832
rect 24333 6809 24367 6832
rect 24401 6809 24435 6832
rect 24469 6809 24503 6832
rect 24537 6809 24540 6843
rect 23752 6793 24540 6809
rect 23752 6774 23781 6793
rect 23815 6774 23853 6793
rect 23887 6774 23925 6793
rect 23752 6740 23755 6774
rect 23815 6759 23823 6774
rect 23887 6759 23891 6774
rect 23789 6740 23823 6759
rect 23857 6740 23891 6759
rect 23959 6774 23997 6793
rect 24031 6774 24069 6793
rect 24103 6774 24141 6793
rect 24175 6774 24213 6793
rect 24247 6774 24285 6793
rect 24319 6774 24357 6793
rect 24391 6774 24429 6793
rect 24463 6774 24501 6793
rect 24535 6774 24540 6793
rect 23925 6740 23959 6759
rect 23993 6759 23997 6774
rect 24061 6759 24069 6774
rect 24129 6759 24141 6774
rect 24197 6759 24213 6774
rect 24265 6759 24285 6774
rect 24333 6759 24357 6774
rect 24401 6759 24429 6774
rect 24469 6759 24501 6774
rect 23993 6740 24027 6759
rect 24061 6740 24095 6759
rect 24129 6740 24163 6759
rect 24197 6740 24231 6759
rect 24265 6740 24299 6759
rect 24333 6740 24367 6759
rect 24401 6740 24435 6759
rect 24469 6740 24503 6759
rect 24537 6740 24540 6774
rect 23752 6720 24540 6740
rect 23752 6705 23781 6720
rect 23815 6705 23853 6720
rect 23887 6705 23925 6720
rect 23752 6671 23755 6705
rect 23815 6686 23823 6705
rect 23887 6686 23891 6705
rect 23789 6671 23823 6686
rect 23857 6671 23891 6686
rect 23959 6705 23997 6720
rect 24031 6705 24069 6720
rect 24103 6705 24141 6720
rect 24175 6705 24213 6720
rect 24247 6705 24285 6720
rect 24319 6705 24357 6720
rect 24391 6705 24429 6720
rect 24463 6705 24501 6720
rect 24535 6705 24540 6720
rect 23925 6671 23959 6686
rect 23993 6686 23997 6705
rect 24061 6686 24069 6705
rect 24129 6686 24141 6705
rect 24197 6686 24213 6705
rect 24265 6686 24285 6705
rect 24333 6686 24357 6705
rect 24401 6686 24429 6705
rect 24469 6686 24501 6705
rect 23993 6671 24027 6686
rect 24061 6671 24095 6686
rect 24129 6671 24163 6686
rect 24197 6671 24231 6686
rect 24265 6671 24299 6686
rect 24333 6671 24367 6686
rect 24401 6671 24435 6686
rect 24469 6671 24503 6686
rect 24537 6671 24540 6705
rect 23752 6647 24540 6671
rect 23752 6636 23781 6647
rect 23815 6636 23853 6647
rect 23887 6636 23925 6647
rect 23752 6602 23755 6636
rect 23815 6613 23823 6636
rect 23887 6613 23891 6636
rect 23789 6602 23823 6613
rect 23857 6602 23891 6613
rect 23959 6636 23997 6647
rect 24031 6636 24069 6647
rect 24103 6636 24141 6647
rect 24175 6636 24213 6647
rect 24247 6636 24285 6647
rect 24319 6636 24357 6647
rect 24391 6636 24429 6647
rect 24463 6636 24501 6647
rect 24535 6636 24540 6647
rect 23925 6602 23959 6613
rect 23993 6613 23997 6636
rect 24061 6613 24069 6636
rect 24129 6613 24141 6636
rect 24197 6613 24213 6636
rect 24265 6613 24285 6636
rect 24333 6613 24357 6636
rect 24401 6613 24429 6636
rect 24469 6613 24501 6636
rect 23993 6602 24027 6613
rect 24061 6602 24095 6613
rect 24129 6602 24163 6613
rect 24197 6602 24231 6613
rect 24265 6602 24299 6613
rect 24333 6602 24367 6613
rect 24401 6602 24435 6613
rect 24469 6602 24503 6613
rect 24537 6602 24540 6636
rect 23752 6574 24540 6602
rect 23752 6567 23781 6574
rect 23815 6567 23853 6574
rect 23887 6567 23925 6574
rect 23752 6533 23755 6567
rect 23815 6540 23823 6567
rect 23887 6540 23891 6567
rect 23789 6533 23823 6540
rect 23857 6533 23891 6540
rect 23959 6567 23997 6574
rect 24031 6567 24069 6574
rect 24103 6567 24141 6574
rect 24175 6567 24213 6574
rect 24247 6567 24285 6574
rect 24319 6567 24357 6574
rect 24391 6567 24429 6574
rect 24463 6567 24501 6574
rect 24535 6567 24540 6574
rect 23925 6533 23959 6540
rect 23993 6540 23997 6567
rect 24061 6540 24069 6567
rect 24129 6540 24141 6567
rect 24197 6540 24213 6567
rect 24265 6540 24285 6567
rect 24333 6540 24357 6567
rect 24401 6540 24429 6567
rect 24469 6540 24501 6567
rect 23993 6533 24027 6540
rect 24061 6533 24095 6540
rect 24129 6533 24163 6540
rect 24197 6533 24231 6540
rect 24265 6533 24299 6540
rect 24333 6533 24367 6540
rect 24401 6533 24435 6540
rect 24469 6533 24503 6540
rect 24537 6533 24540 6567
rect 23752 6501 24540 6533
rect 23752 6498 23781 6501
rect 23815 6498 23853 6501
rect 23887 6498 23925 6501
rect 23752 6464 23755 6498
rect 23815 6467 23823 6498
rect 23887 6467 23891 6498
rect 23789 6464 23823 6467
rect 23857 6464 23891 6467
rect 23959 6498 23997 6501
rect 24031 6498 24069 6501
rect 24103 6498 24141 6501
rect 24175 6498 24213 6501
rect 24247 6498 24285 6501
rect 24319 6498 24357 6501
rect 24391 6498 24429 6501
rect 24463 6498 24501 6501
rect 24535 6498 24540 6501
rect 23925 6464 23959 6467
rect 23993 6467 23997 6498
rect 24061 6467 24069 6498
rect 24129 6467 24141 6498
rect 24197 6467 24213 6498
rect 24265 6467 24285 6498
rect 24333 6467 24357 6498
rect 24401 6467 24429 6498
rect 24469 6467 24501 6498
rect 23993 6464 24027 6467
rect 24061 6464 24095 6467
rect 24129 6464 24163 6467
rect 24197 6464 24231 6467
rect 24265 6464 24299 6467
rect 24333 6464 24367 6467
rect 24401 6464 24435 6467
rect 24469 6464 24503 6467
rect 24537 6464 24540 6498
rect 23752 6429 24540 6464
rect 23752 6395 23755 6429
rect 23789 6428 23823 6429
rect 23857 6428 23891 6429
rect 23815 6395 23823 6428
rect 23887 6395 23891 6428
rect 23925 6428 23959 6429
rect 23752 6394 23781 6395
rect 23815 6394 23853 6395
rect 23887 6394 23925 6395
rect 23993 6428 24027 6429
rect 24061 6428 24095 6429
rect 24129 6428 24163 6429
rect 24197 6428 24231 6429
rect 24265 6428 24299 6429
rect 24333 6428 24367 6429
rect 24401 6428 24435 6429
rect 24469 6428 24503 6429
rect 23993 6395 23997 6428
rect 24061 6395 24069 6428
rect 24129 6395 24141 6428
rect 24197 6395 24213 6428
rect 24265 6395 24285 6428
rect 24333 6395 24357 6428
rect 24401 6395 24429 6428
rect 24469 6395 24501 6428
rect 24537 6395 24540 6429
rect 23959 6394 23997 6395
rect 24031 6394 24069 6395
rect 24103 6394 24141 6395
rect 24175 6394 24213 6395
rect 24247 6394 24285 6395
rect 24319 6394 24357 6395
rect 24391 6394 24429 6395
rect 24463 6394 24501 6395
rect 24535 6394 24540 6395
rect 23752 6360 24540 6394
rect 23752 6326 23755 6360
rect 23789 6355 23823 6360
rect 23857 6355 23891 6360
rect 23815 6326 23823 6355
rect 23887 6326 23891 6355
rect 23925 6355 23959 6360
rect 23752 6321 23781 6326
rect 23815 6321 23853 6326
rect 23887 6321 23925 6326
rect 23993 6355 24027 6360
rect 24061 6355 24095 6360
rect 24129 6355 24163 6360
rect 24197 6355 24231 6360
rect 24265 6355 24299 6360
rect 24333 6355 24367 6360
rect 24401 6355 24435 6360
rect 24469 6355 24503 6360
rect 23993 6326 23997 6355
rect 24061 6326 24069 6355
rect 24129 6326 24141 6355
rect 24197 6326 24213 6355
rect 24265 6326 24285 6355
rect 24333 6326 24357 6355
rect 24401 6326 24429 6355
rect 24469 6326 24501 6355
rect 24537 6326 24540 6360
rect 23959 6321 23997 6326
rect 24031 6321 24069 6326
rect 24103 6321 24141 6326
rect 24175 6321 24213 6326
rect 24247 6321 24285 6326
rect 24319 6321 24357 6326
rect 24391 6321 24429 6326
rect 24463 6321 24501 6326
rect 24535 6321 24540 6326
rect 23752 6291 24540 6321
rect 23752 6257 23755 6291
rect 23789 6282 23823 6291
rect 23857 6282 23891 6291
rect 23815 6257 23823 6282
rect 23887 6257 23891 6282
rect 23925 6282 23959 6291
rect 23752 6248 23781 6257
rect 23815 6248 23853 6257
rect 23887 6248 23925 6257
rect 23993 6282 24027 6291
rect 24061 6282 24095 6291
rect 24129 6282 24163 6291
rect 24197 6282 24231 6291
rect 24265 6282 24299 6291
rect 24333 6282 24367 6291
rect 24401 6282 24435 6291
rect 24469 6282 24503 6291
rect 23993 6257 23997 6282
rect 24061 6257 24069 6282
rect 24129 6257 24141 6282
rect 24197 6257 24213 6282
rect 24265 6257 24285 6282
rect 24333 6257 24357 6282
rect 24401 6257 24429 6282
rect 24469 6257 24501 6282
rect 24537 6257 24540 6291
rect 23959 6248 23997 6257
rect 24031 6248 24069 6257
rect 24103 6248 24141 6257
rect 24175 6248 24213 6257
rect 24247 6248 24285 6257
rect 24319 6248 24357 6257
rect 24391 6248 24429 6257
rect 24463 6248 24501 6257
rect 24535 6248 24540 6257
rect 23752 6222 24540 6248
rect 23752 6188 23755 6222
rect 23789 6209 23823 6222
rect 23857 6209 23891 6222
rect 23815 6188 23823 6209
rect 23887 6188 23891 6209
rect 23925 6209 23959 6222
rect 23752 6175 23781 6188
rect 23815 6175 23853 6188
rect 23887 6175 23925 6188
rect 23993 6209 24027 6222
rect 24061 6209 24095 6222
rect 24129 6209 24163 6222
rect 24197 6209 24231 6222
rect 24265 6209 24299 6222
rect 24333 6209 24367 6222
rect 24401 6209 24435 6222
rect 24469 6209 24503 6222
rect 23993 6188 23997 6209
rect 24061 6188 24069 6209
rect 24129 6188 24141 6209
rect 24197 6188 24213 6209
rect 24265 6188 24285 6209
rect 24333 6188 24357 6209
rect 24401 6188 24429 6209
rect 24469 6188 24501 6209
rect 24537 6188 24540 6222
rect 23959 6175 23997 6188
rect 24031 6175 24069 6188
rect 24103 6175 24141 6188
rect 24175 6175 24213 6188
rect 24247 6175 24285 6188
rect 24319 6175 24357 6188
rect 24391 6175 24429 6188
rect 24463 6175 24501 6188
rect 24535 6175 24540 6188
rect 23752 6153 24540 6175
rect 23752 6119 23755 6153
rect 23789 6136 23823 6153
rect 23857 6136 23891 6153
rect 23815 6119 23823 6136
rect 23887 6119 23891 6136
rect 23925 6136 23959 6153
rect 23752 6102 23781 6119
rect 23815 6102 23853 6119
rect 23887 6102 23925 6119
rect 23993 6136 24027 6153
rect 24061 6136 24095 6153
rect 24129 6136 24163 6153
rect 24197 6136 24231 6153
rect 24265 6136 24299 6153
rect 24333 6136 24367 6153
rect 24401 6136 24435 6153
rect 24469 6136 24503 6153
rect 23993 6119 23997 6136
rect 24061 6119 24069 6136
rect 24129 6119 24141 6136
rect 24197 6119 24213 6136
rect 24265 6119 24285 6136
rect 24333 6119 24357 6136
rect 24401 6119 24429 6136
rect 24469 6119 24501 6136
rect 24537 6119 24540 6153
rect 23959 6102 23997 6119
rect 24031 6102 24069 6119
rect 24103 6102 24141 6119
rect 24175 6102 24213 6119
rect 24247 6102 24285 6119
rect 24319 6102 24357 6119
rect 24391 6102 24429 6119
rect 24463 6102 24501 6119
rect 24535 6102 24540 6119
rect 23752 6084 24540 6102
rect 23752 6050 23755 6084
rect 23789 6063 23823 6084
rect 23857 6063 23891 6084
rect 23815 6050 23823 6063
rect 23887 6050 23891 6063
rect 23925 6063 23959 6084
rect 23752 6029 23781 6050
rect 23815 6029 23853 6050
rect 23887 6029 23925 6050
rect 23993 6063 24027 6084
rect 24061 6063 24095 6084
rect 24129 6063 24163 6084
rect 24197 6063 24231 6084
rect 24265 6063 24299 6084
rect 24333 6063 24367 6084
rect 24401 6063 24435 6084
rect 24469 6063 24503 6084
rect 23993 6050 23997 6063
rect 24061 6050 24069 6063
rect 24129 6050 24141 6063
rect 24197 6050 24213 6063
rect 24265 6050 24285 6063
rect 24333 6050 24357 6063
rect 24401 6050 24429 6063
rect 24469 6050 24501 6063
rect 24537 6050 24540 6084
rect 23959 6029 23997 6050
rect 24031 6029 24069 6050
rect 24103 6029 24141 6050
rect 24175 6029 24213 6050
rect 24247 6029 24285 6050
rect 24319 6029 24357 6050
rect 24391 6029 24429 6050
rect 24463 6029 24501 6050
rect 24535 6029 24540 6050
rect 23752 6015 24540 6029
rect 23752 5981 23755 6015
rect 23789 5990 23823 6015
rect 23857 5990 23891 6015
rect 23815 5981 23823 5990
rect 23887 5981 23891 5990
rect 23925 5990 23959 6015
rect 23752 5956 23781 5981
rect 23815 5956 23853 5981
rect 23887 5956 23925 5981
rect 23993 5990 24027 6015
rect 24061 5990 24095 6015
rect 24129 5990 24163 6015
rect 24197 5990 24231 6015
rect 24265 5990 24299 6015
rect 24333 5990 24367 6015
rect 24401 5990 24435 6015
rect 24469 5990 24503 6015
rect 23993 5981 23997 5990
rect 24061 5981 24069 5990
rect 24129 5981 24141 5990
rect 24197 5981 24213 5990
rect 24265 5981 24285 5990
rect 24333 5981 24357 5990
rect 24401 5981 24429 5990
rect 24469 5981 24501 5990
rect 24537 5981 24540 6015
rect 23959 5956 23997 5981
rect 24031 5956 24069 5981
rect 24103 5956 24141 5981
rect 24175 5956 24213 5981
rect 24247 5956 24285 5981
rect 24319 5956 24357 5981
rect 24391 5956 24429 5981
rect 24463 5956 24501 5981
rect 24535 5956 24540 5981
rect 23752 5946 24540 5956
rect 23752 5912 23755 5946
rect 23789 5917 23823 5946
rect 23857 5917 23891 5946
rect 23815 5912 23823 5917
rect 23887 5912 23891 5917
rect 23925 5917 23959 5946
rect 23752 5883 23781 5912
rect 23815 5883 23853 5912
rect 23887 5883 23925 5912
rect 23993 5917 24027 5946
rect 24061 5917 24095 5946
rect 24129 5917 24163 5946
rect 24197 5917 24231 5946
rect 24265 5917 24299 5946
rect 24333 5917 24367 5946
rect 24401 5917 24435 5946
rect 24469 5917 24503 5946
rect 23993 5912 23997 5917
rect 24061 5912 24069 5917
rect 24129 5912 24141 5917
rect 24197 5912 24213 5917
rect 24265 5912 24285 5917
rect 24333 5912 24357 5917
rect 24401 5912 24429 5917
rect 24469 5912 24501 5917
rect 24537 5912 24540 5946
rect 23959 5883 23997 5912
rect 24031 5883 24069 5912
rect 24103 5883 24141 5912
rect 24175 5883 24213 5912
rect 24247 5883 24285 5912
rect 24319 5883 24357 5912
rect 24391 5883 24429 5912
rect 24463 5883 24501 5912
rect 24535 5883 24540 5912
rect 23752 5877 24540 5883
rect 23752 5639 23755 5877
rect 24537 5639 24540 5877
rect 23752 5615 23981 5639
rect 22766 5571 22818 5610
rect 22766 5537 22798 5571
rect 22766 5498 22818 5537
rect 22766 5464 22798 5498
rect 22832 5464 22870 5485
rect 22904 5464 22942 5485
rect 22976 5464 23014 5485
rect 23048 5464 23086 5485
rect 23120 5464 23158 5485
rect 23192 5464 23230 5485
rect 23264 5464 23302 5485
rect 23336 5464 23374 5485
rect 23408 5464 23446 5485
rect 23480 5464 23600 5485
rect 22766 5463 23600 5464
rect 23949 5532 23981 5615
rect 24087 5591 24540 5639
rect 24087 5557 24153 5591
rect 24187 5557 24221 5591
rect 24255 5557 24289 5591
rect 24323 5557 24357 5591
rect 24391 5557 24425 5591
rect 24459 5557 24493 5591
rect 24527 5557 24540 5591
rect 24087 5532 24540 5557
rect 22766 5440 23796 5463
rect 22766 5425 22842 5440
rect 22944 5425 22979 5440
rect 22766 5391 22798 5425
rect 22832 5391 22842 5425
rect 22976 5406 22979 5425
rect 23013 5425 23048 5440
rect 23013 5406 23014 5425
rect 22976 5391 23014 5406
rect 23082 5425 23117 5440
rect 23151 5425 23186 5440
rect 23220 5425 23255 5440
rect 23289 5425 23324 5440
rect 23358 5425 23393 5440
rect 23427 5425 23462 5440
rect 23082 5406 23086 5425
rect 23151 5406 23158 5425
rect 23220 5406 23230 5425
rect 23289 5406 23302 5425
rect 23358 5406 23374 5425
rect 23427 5406 23446 5425
rect 23496 5406 23531 5440
rect 23565 5406 23600 5440
rect 23634 5406 23669 5440
rect 23703 5406 23738 5440
rect 23772 5406 23796 5440
rect 23048 5391 23086 5406
rect 23120 5391 23158 5406
rect 23192 5391 23230 5406
rect 23264 5391 23302 5406
rect 23336 5391 23374 5406
rect 23408 5391 23446 5406
rect 23480 5391 23796 5406
rect 22766 5352 22842 5391
rect 22944 5372 23796 5391
rect 22944 5352 22979 5372
rect 22766 5318 22798 5352
rect 22832 5318 22842 5352
rect 22976 5338 22979 5352
rect 23013 5352 23048 5372
rect 23013 5338 23014 5352
rect 22976 5318 23014 5338
rect 23082 5352 23117 5372
rect 23151 5352 23186 5372
rect 23220 5352 23255 5372
rect 23289 5352 23324 5372
rect 23358 5352 23393 5372
rect 23427 5352 23462 5372
rect 23082 5338 23086 5352
rect 23151 5338 23158 5352
rect 23220 5338 23230 5352
rect 23289 5338 23302 5352
rect 23358 5338 23374 5352
rect 23427 5338 23446 5352
rect 23496 5338 23531 5372
rect 23565 5338 23600 5372
rect 23634 5338 23669 5372
rect 23703 5338 23738 5372
rect 23772 5338 23796 5372
rect 23048 5318 23086 5338
rect 23120 5318 23158 5338
rect 23192 5318 23230 5338
rect 23264 5318 23302 5338
rect 23336 5318 23374 5338
rect 23408 5318 23446 5338
rect 23480 5318 23796 5338
rect 22766 5280 22842 5318
rect 22944 5304 23796 5318
rect 22944 5280 22979 5304
rect 23013 5280 23048 5304
rect 23082 5280 23117 5304
rect 23151 5280 23186 5304
rect 22766 5246 22782 5280
rect 22816 5246 22842 5280
rect 22962 5270 22979 5280
rect 23035 5270 23048 5280
rect 23108 5270 23117 5280
rect 23181 5270 23186 5280
rect 23220 5280 23255 5304
rect 22962 5246 23001 5270
rect 23035 5246 23074 5270
rect 23108 5246 23147 5270
rect 23181 5246 23220 5270
rect 23254 5270 23255 5280
rect 23289 5280 23324 5304
rect 23358 5280 23393 5304
rect 23427 5280 23462 5304
rect 23496 5280 23531 5304
rect 23289 5270 23294 5280
rect 23358 5270 23368 5280
rect 23427 5270 23442 5280
rect 23496 5270 23516 5280
rect 23565 5274 23600 5304
rect 23634 5274 23669 5304
rect 23703 5274 23738 5304
rect 23565 5270 23593 5274
rect 23634 5270 23665 5274
rect 23703 5270 23737 5274
rect 23772 5270 23796 5304
rect 23254 5246 23294 5270
rect 23328 5246 23368 5270
rect 23402 5246 23442 5270
rect 23476 5246 23516 5270
rect 23550 5246 23593 5270
rect 22766 5208 22842 5246
rect 22944 5240 23593 5246
rect 23627 5240 23665 5270
rect 23699 5240 23737 5270
rect 23771 5240 23796 5270
rect 22944 5236 23796 5240
rect 22944 5208 22979 5236
rect 23013 5208 23048 5236
rect 23082 5208 23117 5236
rect 23151 5208 23186 5236
rect 22766 5174 22782 5208
rect 22816 5174 22842 5208
rect 22962 5202 22979 5208
rect 23035 5202 23048 5208
rect 23108 5202 23117 5208
rect 23181 5202 23186 5208
rect 23220 5208 23255 5236
rect 22962 5174 23001 5202
rect 23035 5174 23074 5202
rect 23108 5174 23147 5202
rect 23181 5174 23220 5202
rect 23254 5202 23255 5208
rect 23289 5208 23324 5236
rect 23358 5208 23393 5236
rect 23427 5208 23462 5236
rect 23496 5208 23531 5236
rect 23289 5202 23294 5208
rect 23358 5202 23368 5208
rect 23427 5202 23442 5208
rect 23496 5202 23516 5208
rect 23565 5202 23600 5236
rect 23634 5202 23669 5236
rect 23703 5202 23738 5236
rect 23772 5202 23796 5236
rect 23254 5174 23294 5202
rect 23328 5174 23368 5202
rect 23402 5174 23442 5202
rect 23476 5174 23516 5202
rect 23550 5201 23796 5202
rect 23550 5174 23593 5201
rect 22766 5136 22842 5174
rect 22944 5168 23593 5174
rect 23627 5168 23665 5201
rect 23699 5168 23737 5201
rect 23771 5168 23796 5201
rect 22944 5136 22979 5168
rect 23013 5136 23048 5168
rect 23082 5136 23117 5168
rect 23151 5136 23186 5168
rect 22766 5102 22782 5136
rect 22816 5102 22842 5136
rect 22962 5134 22979 5136
rect 23035 5134 23048 5136
rect 23108 5134 23117 5136
rect 23181 5134 23186 5136
rect 23220 5136 23255 5168
rect 22962 5102 23001 5134
rect 23035 5102 23074 5134
rect 23108 5102 23147 5134
rect 23181 5102 23220 5134
rect 23254 5134 23255 5136
rect 23289 5136 23324 5168
rect 23358 5136 23393 5168
rect 23427 5136 23462 5168
rect 23496 5136 23531 5168
rect 23565 5167 23593 5168
rect 23634 5167 23665 5168
rect 23703 5167 23737 5168
rect 23289 5134 23294 5136
rect 23358 5134 23368 5136
rect 23427 5134 23442 5136
rect 23496 5134 23516 5136
rect 23565 5134 23600 5167
rect 23634 5134 23669 5167
rect 23703 5134 23738 5167
rect 23772 5134 23796 5168
rect 23254 5102 23294 5134
rect 23328 5102 23368 5134
rect 23402 5102 23442 5134
rect 23476 5102 23516 5134
rect 23550 5128 23796 5134
rect 23550 5102 23593 5128
rect 22766 5064 22842 5102
rect 22944 5100 23593 5102
rect 23627 5100 23665 5128
rect 23699 5100 23737 5128
rect 23771 5100 23796 5128
rect 22944 5066 22979 5100
rect 23013 5066 23048 5100
rect 23082 5066 23117 5100
rect 23151 5066 23186 5100
rect 23220 5066 23255 5100
rect 23289 5066 23324 5100
rect 23358 5066 23393 5100
rect 23427 5066 23462 5100
rect 23496 5066 23531 5100
rect 23565 5094 23593 5100
rect 23634 5094 23665 5100
rect 23703 5094 23737 5100
rect 23565 5066 23600 5094
rect 23634 5066 23669 5094
rect 23703 5066 23738 5094
rect 23772 5066 23796 5100
rect 22944 5064 23796 5066
rect 22766 5030 22782 5064
rect 22816 5030 22842 5064
rect 22962 5032 23001 5064
rect 23035 5032 23074 5064
rect 23108 5032 23147 5064
rect 23181 5032 23220 5064
rect 22962 5030 22979 5032
rect 23035 5030 23048 5032
rect 23108 5030 23117 5032
rect 23181 5030 23186 5032
rect 22766 4992 22842 5030
rect 22944 4998 22979 5030
rect 23013 4998 23048 5030
rect 23082 4998 23117 5030
rect 23151 4998 23186 5030
rect 23254 5032 23294 5064
rect 23328 5032 23368 5064
rect 23402 5032 23442 5064
rect 23476 5032 23516 5064
rect 23550 5055 23796 5064
rect 23550 5032 23593 5055
rect 23627 5032 23665 5055
rect 23699 5032 23737 5055
rect 23771 5032 23796 5055
rect 23254 5030 23255 5032
rect 23220 4998 23255 5030
rect 23289 5030 23294 5032
rect 23358 5030 23368 5032
rect 23427 5030 23442 5032
rect 23496 5030 23516 5032
rect 23289 4998 23324 5030
rect 23358 4998 23393 5030
rect 23427 4998 23462 5030
rect 23496 4998 23531 5030
rect 23565 5021 23593 5032
rect 23634 5021 23665 5032
rect 23703 5021 23737 5032
rect 23565 4998 23600 5021
rect 23634 4998 23669 5021
rect 23703 4998 23738 5021
rect 23772 4998 23796 5032
rect 22944 4992 23796 4998
rect 22766 4958 22782 4992
rect 22816 4958 22842 4992
rect 22962 4964 23001 4992
rect 23035 4964 23074 4992
rect 23108 4964 23147 4992
rect 23181 4964 23220 4992
rect 22962 4958 22979 4964
rect 23035 4958 23048 4964
rect 23108 4958 23117 4964
rect 23181 4958 23186 4964
rect 22766 4794 22842 4958
rect 22944 4930 22979 4958
rect 23013 4930 23048 4958
rect 23082 4930 23117 4958
rect 23151 4930 23186 4958
rect 23254 4964 23294 4992
rect 23328 4964 23368 4992
rect 23402 4964 23442 4992
rect 23476 4964 23516 4992
rect 23550 4982 23796 4992
rect 23550 4964 23593 4982
rect 23627 4964 23665 4982
rect 23699 4964 23737 4982
rect 23771 4964 23796 4982
rect 23254 4958 23255 4964
rect 23220 4930 23255 4958
rect 23289 4958 23294 4964
rect 23358 4958 23368 4964
rect 23427 4958 23442 4964
rect 23496 4958 23516 4964
rect 23289 4930 23324 4958
rect 23358 4930 23393 4958
rect 23427 4930 23462 4958
rect 23496 4930 23531 4958
rect 23565 4948 23593 4964
rect 23634 4948 23665 4964
rect 23703 4948 23737 4964
rect 23565 4930 23600 4948
rect 23634 4930 23669 4948
rect 23703 4930 23738 4948
rect 23772 4930 23796 4964
rect 22944 4909 23796 4930
rect 22944 4896 23593 4909
rect 23627 4896 23665 4909
rect 23699 4896 23737 4909
rect 23771 4896 23796 4909
rect 22944 4862 22979 4896
rect 23013 4862 23048 4896
rect 23082 4862 23117 4896
rect 23151 4862 23186 4896
rect 23220 4862 23255 4896
rect 23289 4862 23324 4896
rect 23358 4862 23393 4896
rect 23427 4862 23462 4896
rect 23496 4862 23531 4896
rect 23565 4875 23593 4896
rect 23634 4875 23665 4896
rect 23703 4875 23737 4896
rect 23565 4862 23600 4875
rect 23634 4862 23669 4875
rect 23703 4862 23738 4875
rect 23772 4862 23796 4896
rect 22944 4836 23796 4862
rect 22944 4828 23593 4836
rect 23627 4828 23665 4836
rect 23699 4828 23737 4836
rect 23771 4828 23796 4836
rect 22944 4794 22979 4828
rect 23013 4794 23048 4828
rect 23082 4794 23117 4828
rect 23151 4794 23186 4828
rect 23220 4794 23255 4828
rect 23289 4794 23324 4828
rect 23358 4794 23393 4828
rect 23427 4794 23462 4828
rect 23496 4794 23531 4828
rect 23565 4802 23593 4828
rect 23634 4802 23665 4828
rect 23703 4802 23737 4828
rect 23565 4794 23600 4802
rect 23634 4794 23669 4802
rect 23703 4794 23738 4802
rect 23772 4794 23796 4828
rect 22766 4771 23796 4794
rect 696 4746 866 4771
rect 696 4737 728 4746
rect 762 4737 800 4746
rect 834 4737 866 4746
rect 762 4712 764 4737
rect 730 4703 764 4712
rect 798 4712 800 4737
rect 798 4703 832 4712
rect 696 4673 866 4703
rect 696 4665 728 4673
rect 762 4672 866 4673
rect 762 4665 800 4672
rect 834 4665 866 4672
rect 762 4639 764 4665
rect 730 4631 764 4639
rect 798 4638 800 4665
rect 798 4631 832 4638
rect 696 4600 866 4631
rect 696 4593 728 4600
rect 762 4598 866 4600
rect 762 4593 800 4598
rect 834 4593 866 4598
rect 762 4566 764 4593
rect 730 4559 764 4566
rect 798 4564 800 4593
rect 23568 4763 23796 4771
rect 23568 4729 23593 4763
rect 23627 4737 23665 4763
rect 23699 4737 23737 4763
rect 23568 4703 23597 4729
rect 23631 4703 23665 4737
rect 23699 4703 23733 4737
rect 23771 4729 23796 4763
rect 23767 4703 23796 4729
rect 23568 4690 23796 4703
rect 23568 4656 23593 4690
rect 23627 4668 23665 4690
rect 23699 4668 23737 4690
rect 23568 4634 23597 4656
rect 23631 4634 23665 4668
rect 23699 4634 23733 4668
rect 23771 4656 23796 4690
rect 23767 4634 23796 4656
rect 23568 4617 23796 4634
rect 23568 4583 23593 4617
rect 23627 4599 23665 4617
rect 23699 4599 23737 4617
rect 798 4559 832 4564
rect 696 4527 866 4559
rect 696 4521 728 4527
rect 762 4524 866 4527
rect 762 4521 800 4524
rect 834 4521 866 4524
rect 278 4483 448 4517
rect 312 4479 346 4483
rect 380 4479 414 4483
rect 278 4413 310 4449
rect 416 4413 448 4449
rect 278 4343 310 4379
rect 416 4343 448 4379
rect 278 4273 310 4309
rect 416 4273 448 4309
rect 278 4203 310 4239
rect 416 4203 448 4239
rect 278 4134 310 4169
rect 416 4134 448 4169
rect 278 4065 310 4100
rect 416 4065 448 4100
rect 278 3996 310 4031
rect 416 3996 448 4031
rect 278 3927 310 3962
rect 416 3927 448 3962
rect 278 3858 310 3893
rect 416 3858 448 3893
rect 278 3789 310 3824
rect 416 3789 448 3824
rect 278 3720 310 3755
rect 416 3720 448 3755
rect 278 3651 310 3686
rect 416 3651 448 3686
rect 278 3582 310 3617
rect 416 3582 448 3617
rect 278 3513 310 3548
rect 416 3513 448 3548
rect 278 3444 310 3479
rect 416 3444 448 3479
rect 278 3375 310 3410
rect 416 3375 448 3410
rect 278 3306 310 3341
rect 416 3306 448 3341
rect 278 3237 310 3272
rect 416 3237 448 3272
rect 278 3168 310 3203
rect 416 3168 448 3203
rect 278 3099 310 3134
rect 416 3099 448 3134
rect 278 3030 310 3065
rect 416 3030 448 3065
rect 278 2961 310 2996
rect 416 2961 448 2996
rect 278 2892 310 2927
rect 416 2892 448 2927
rect 278 2823 310 2858
rect 416 2823 448 2858
rect 278 2754 310 2789
rect 416 2754 448 2789
rect 278 2685 310 2720
rect 416 2685 448 2720
rect 278 2616 310 2651
rect 416 2616 448 2651
rect 278 2573 310 2582
rect 416 2573 448 2582
rect 278 2547 448 2573
rect 312 2534 346 2547
rect 344 2513 346 2534
rect 380 2534 414 2547
rect 380 2513 382 2534
rect 278 2500 310 2513
rect 344 2500 382 2513
rect 416 2500 448 2513
rect 278 2478 448 2500
rect 312 2461 346 2478
rect 344 2444 346 2461
rect 380 2461 414 2478
rect 380 2444 382 2461
rect 278 2427 310 2444
rect 344 2427 382 2444
rect 416 2427 448 2444
rect 278 2409 448 2427
rect 312 2388 346 2409
rect 344 2375 346 2388
rect 380 2388 414 2409
rect 380 2375 382 2388
rect 278 2354 310 2375
rect 344 2354 382 2375
rect 416 2354 448 2375
rect 278 2340 448 2354
rect 312 2315 346 2340
rect 344 2306 346 2315
rect 380 2315 414 2340
rect 380 2306 382 2315
rect 278 2281 310 2306
rect 344 2281 382 2306
rect 416 2281 448 2306
rect 278 2271 448 2281
rect 312 2242 346 2271
rect 344 2237 346 2242
rect 380 2242 414 2271
rect 380 2237 382 2242
rect 278 2208 310 2237
rect 344 2208 382 2237
rect 416 2208 448 2237
rect 278 2202 448 2208
rect 312 2169 346 2202
rect 344 2168 346 2169
rect 380 2169 414 2202
rect 380 2168 382 2169
rect 278 2135 310 2168
rect 344 2135 382 2168
rect 416 2135 448 2168
rect 278 2133 448 2135
rect 312 2099 346 2133
rect 380 2099 414 2133
rect 278 2096 448 2099
rect 278 2064 310 2096
rect 344 2064 382 2096
rect 416 2064 448 2096
rect 344 2062 346 2064
rect 312 2030 346 2062
rect 380 2062 382 2064
rect 380 2030 414 2062
rect 278 2023 448 2030
rect 278 1995 310 2023
rect 344 1995 382 2023
rect 416 1995 448 2023
rect 344 1989 346 1995
rect 312 1961 346 1989
rect 380 1989 382 1995
rect 380 1961 414 1989
rect 278 1950 448 1961
rect 278 1926 310 1950
rect 344 1926 382 1950
rect 416 1926 448 1950
rect 344 1916 346 1926
rect 312 1892 346 1916
rect 380 1916 382 1926
rect 380 1892 414 1916
rect 278 1877 448 1892
rect 278 1857 310 1877
rect 344 1857 382 1877
rect 416 1857 448 1877
rect 344 1843 346 1857
rect 312 1823 346 1843
rect 380 1843 382 1857
rect 380 1823 414 1843
rect 278 1804 448 1823
rect 278 1788 310 1804
rect 344 1788 382 1804
rect 416 1788 448 1804
rect 344 1770 346 1788
rect 312 1754 346 1770
rect 380 1770 382 1788
rect 380 1754 414 1770
rect 278 1731 448 1754
rect 278 1719 310 1731
rect 344 1719 382 1731
rect 416 1719 448 1731
rect 344 1697 346 1719
rect 312 1685 346 1697
rect 380 1697 382 1719
rect 380 1685 414 1697
rect 278 1658 448 1685
rect 278 1650 310 1658
rect 344 1650 382 1658
rect 416 1650 448 1658
rect 344 1624 346 1650
rect 312 1616 346 1624
rect 380 1624 382 1650
rect 380 1616 414 1624
rect 278 1585 448 1616
rect 278 1581 310 1585
rect 344 1581 382 1585
rect 416 1581 448 1585
rect 344 1551 346 1581
rect 312 1547 346 1551
rect 380 1551 382 1581
rect 380 1547 414 1551
rect 278 1512 448 1547
rect 344 1478 346 1512
rect 380 1478 382 1512
rect 278 1443 448 1478
rect 312 1439 346 1443
rect 344 1409 346 1439
rect 380 1439 414 1443
rect 380 1409 382 1439
rect 278 1405 310 1409
rect 344 1405 382 1409
rect 416 1405 448 1409
rect 278 1374 448 1405
rect 312 1366 346 1374
rect 344 1340 346 1366
rect 380 1366 414 1374
rect 380 1340 382 1366
rect 278 1332 310 1340
rect 344 1332 382 1340
rect 416 1332 448 1340
rect 278 1305 448 1332
rect 312 1293 346 1305
rect 344 1271 346 1293
rect 380 1293 414 1305
rect 380 1271 382 1293
rect 278 1259 310 1271
rect 344 1259 382 1271
rect 416 1259 448 1271
rect 278 1236 448 1259
rect 312 1220 346 1236
rect 344 1202 346 1220
rect 380 1220 414 1236
rect 380 1202 382 1220
rect 278 1186 310 1202
rect 344 1186 382 1202
rect 416 1186 448 1202
rect 278 1167 448 1186
rect 312 1147 346 1167
rect 344 1133 346 1147
rect 380 1147 414 1167
rect 380 1133 382 1147
rect 278 1113 310 1133
rect 344 1113 382 1133
rect 416 1113 448 1133
rect 278 1098 448 1113
rect 312 1074 346 1098
rect 344 1064 346 1074
rect 380 1074 414 1098
rect 380 1064 382 1074
rect 278 1040 310 1064
rect 344 1040 382 1064
rect 416 1040 448 1064
rect 278 1029 448 1040
rect 312 1001 346 1029
rect 344 995 346 1001
rect 380 1001 414 1029
rect 380 995 382 1001
rect 278 967 310 995
rect 344 967 382 995
rect 416 967 448 995
rect 278 960 448 967
rect 312 928 346 960
rect 344 926 346 928
rect 380 928 414 960
rect 380 926 382 928
rect 278 894 310 926
rect 344 894 382 926
rect 416 894 448 926
rect 278 891 448 894
rect 312 857 346 891
rect 380 857 414 891
rect 762 4493 764 4521
rect 730 4487 764 4493
rect 798 4490 800 4521
rect 798 4487 832 4490
rect 696 4454 866 4487
rect 696 4449 728 4454
rect 762 4450 866 4454
rect 762 4449 800 4450
rect 834 4449 866 4450
rect 762 4420 764 4449
rect 730 4415 764 4420
rect 798 4416 800 4449
rect 798 4415 832 4416
rect 696 4381 866 4415
rect 696 4377 728 4381
rect 762 4377 866 4381
rect 762 4347 764 4377
rect 730 4343 764 4347
rect 798 4376 832 4377
rect 798 4343 800 4376
rect 696 4342 800 4343
rect 834 4342 866 4343
rect 696 4308 866 4342
rect 696 4305 728 4308
rect 762 4305 866 4308
rect 762 4274 764 4305
rect 730 4271 764 4274
rect 798 4302 832 4305
rect 798 4271 800 4302
rect 696 4268 800 4271
rect 834 4268 866 4271
rect 696 4235 866 4268
rect 696 4233 728 4235
rect 762 4233 866 4235
rect 762 4201 764 4233
rect 730 4199 764 4201
rect 798 4228 832 4233
rect 798 4199 800 4228
rect 696 4194 800 4199
rect 834 4194 866 4199
rect 696 4162 866 4194
rect 696 4161 728 4162
rect 762 4161 866 4162
rect 762 4128 764 4161
rect 730 4127 764 4128
rect 798 4154 832 4161
rect 798 4127 800 4154
rect 696 4120 800 4127
rect 834 4120 866 4127
rect 696 4089 866 4120
rect 762 4055 764 4089
rect 798 4080 832 4089
rect 798 4055 800 4080
rect 696 4046 800 4055
rect 834 4046 866 4055
rect 696 4017 866 4046
rect 730 4016 764 4017
rect 762 3983 764 4016
rect 798 4006 832 4017
rect 798 3983 800 4006
rect 696 3982 728 3983
rect 762 3982 800 3983
rect 696 3972 800 3982
rect 834 3972 866 3983
rect 696 3946 866 3972
rect 730 3943 764 3946
rect 762 3912 764 3943
rect 798 3932 832 3946
rect 798 3912 800 3932
rect 696 3909 728 3912
rect 762 3909 800 3912
rect 696 3898 800 3909
rect 834 3898 866 3912
rect 696 3875 866 3898
rect 730 3870 764 3875
rect 762 3841 764 3870
rect 798 3858 832 3875
rect 798 3841 800 3858
rect 696 3836 728 3841
rect 762 3836 800 3841
rect 696 3824 800 3836
rect 834 3824 866 3841
rect 696 3804 866 3824
rect 730 3797 764 3804
rect 762 3770 764 3797
rect 798 3784 832 3804
rect 798 3770 800 3784
rect 696 3763 728 3770
rect 762 3763 800 3770
rect 696 3750 800 3763
rect 834 3750 866 3770
rect 696 3733 866 3750
rect 730 3724 764 3733
rect 762 3699 764 3724
rect 798 3710 832 3733
rect 798 3699 800 3710
rect 696 3690 728 3699
rect 762 3690 800 3699
rect 696 3676 800 3690
rect 834 3676 866 3699
rect 696 3662 866 3676
rect 730 3651 764 3662
rect 762 3628 764 3651
rect 798 3636 832 3662
rect 798 3628 800 3636
rect 696 3617 728 3628
rect 762 3617 800 3628
rect 696 3602 800 3617
rect 834 3602 866 3628
rect 696 3591 866 3602
rect 730 3578 764 3591
rect 762 3557 764 3578
rect 798 3562 832 3591
rect 798 3557 800 3562
rect 696 3544 728 3557
rect 762 3544 800 3557
rect 696 3528 800 3544
rect 834 3528 866 3557
rect 696 3520 866 3528
rect 730 3505 764 3520
rect 762 3486 764 3505
rect 798 3488 832 3520
rect 798 3486 800 3488
rect 696 3471 728 3486
rect 762 3471 800 3486
rect 696 3454 800 3471
rect 834 3454 866 3486
rect 696 3449 866 3454
rect 730 3432 764 3449
rect 762 3415 764 3432
rect 798 3415 832 3449
rect 696 3398 728 3415
rect 762 3414 866 3415
rect 762 3398 800 3414
rect 696 3380 800 3398
rect 834 3380 866 3414
rect 696 3378 866 3380
rect 730 3359 764 3378
rect 762 3344 764 3359
rect 798 3344 832 3378
rect 696 3325 728 3344
rect 762 3341 866 3344
rect 762 3325 800 3341
rect 696 3307 800 3325
rect 834 3307 866 3341
rect 696 3286 866 3307
rect 762 3252 764 3286
rect 798 3268 832 3286
rect 798 3252 800 3268
rect 696 3234 800 3252
rect 834 3234 866 3252
rect 696 3217 866 3234
rect 696 3216 764 3217
rect 730 3213 764 3216
rect 762 3183 764 3213
rect 798 3195 832 3217
rect 798 3183 800 3195
rect 696 3179 728 3182
rect 762 3179 800 3183
rect 696 3161 800 3179
rect 834 3161 866 3183
rect 696 3148 866 3161
rect 696 3146 764 3148
rect 730 3140 764 3146
rect 762 3114 764 3140
rect 798 3122 832 3148
rect 798 3114 800 3122
rect 696 3106 728 3112
rect 762 3106 800 3114
rect 696 3088 800 3106
rect 834 3088 866 3114
rect 696 3079 866 3088
rect 696 3076 764 3079
rect 730 3067 764 3076
rect 762 3045 764 3067
rect 798 3049 832 3079
rect 798 3045 800 3049
rect 696 3033 728 3042
rect 762 3033 800 3045
rect 696 3015 800 3033
rect 834 3015 866 3045
rect 696 3010 866 3015
rect 696 3006 764 3010
rect 730 2994 764 3006
rect 762 2976 764 2994
rect 798 2976 832 3010
rect 696 2960 728 2972
rect 762 2960 800 2976
rect 696 2942 800 2960
rect 834 2942 866 2976
rect 696 2941 866 2942
rect 696 2937 764 2941
rect 730 2921 764 2937
rect 696 2887 728 2903
rect 762 2887 764 2921
rect 696 2868 764 2887
rect 730 2848 764 2868
rect 696 2814 728 2834
rect 762 2814 764 2848
rect 696 2799 764 2814
rect 730 2775 764 2799
rect 696 2741 728 2765
rect 762 2741 764 2775
rect 696 2730 764 2741
rect 730 2702 764 2730
rect 696 2668 728 2696
rect 762 2668 764 2702
rect 696 2661 764 2668
rect 730 2629 764 2661
rect 696 2595 728 2627
rect 762 2595 764 2629
rect 696 2592 764 2595
rect 730 2558 764 2592
rect 696 2556 764 2558
rect 696 2523 728 2556
rect 762 2522 764 2556
rect 730 2489 764 2522
rect 696 2483 764 2489
rect 696 2454 728 2483
rect 762 2449 764 2483
rect 730 2420 764 2449
rect 696 2411 764 2420
rect 696 2385 728 2411
rect 762 2377 764 2411
rect 730 2351 764 2377
rect 696 2339 764 2351
rect 696 2316 728 2339
rect 762 2305 764 2339
rect 730 2282 764 2305
rect 696 2267 764 2282
rect 696 2247 728 2267
rect 762 2233 764 2267
rect 730 2213 764 2233
rect 696 2195 764 2213
rect 696 2178 728 2195
rect 762 2161 764 2195
rect 730 2144 764 2161
rect 696 2123 764 2144
rect 696 2109 728 2123
rect 762 2089 764 2123
rect 730 2075 764 2089
rect 696 2051 764 2075
rect 696 2040 728 2051
rect 762 2017 764 2051
rect 730 2006 764 2017
rect 696 1979 764 2006
rect 696 1971 728 1979
rect 762 1945 764 1979
rect 730 1937 764 1945
rect 696 1907 764 1937
rect 696 1902 728 1907
rect 762 1873 764 1907
rect 730 1868 764 1873
rect 696 1835 764 1868
rect 696 1833 728 1835
rect 762 1801 764 1835
rect 730 1799 764 1801
rect 696 1764 764 1799
rect 730 1763 764 1764
rect 696 1729 728 1730
rect 762 1729 764 1763
rect 696 1695 764 1729
rect 730 1691 764 1695
rect 696 1657 728 1661
rect 762 1657 764 1691
rect 696 1626 764 1657
rect 730 1619 764 1626
rect 696 1585 728 1592
rect 762 1585 764 1619
rect 696 1557 764 1585
rect 730 1547 764 1557
rect 696 1513 728 1523
rect 762 1513 764 1547
rect 696 1488 764 1513
rect 730 1475 764 1488
rect 696 1441 728 1454
rect 762 1441 764 1475
rect 696 1419 764 1441
rect 730 1403 764 1419
rect 696 1369 728 1385
rect 762 1369 764 1403
rect 696 1350 764 1369
rect 730 1331 764 1350
rect 696 1297 728 1316
rect 762 1297 764 1331
rect 1086 4550 1609 4574
rect 1120 4516 1154 4550
rect 1188 4516 1222 4550
rect 1256 4516 1290 4550
rect 1324 4516 1358 4550
rect 1392 4516 1426 4550
rect 1460 4540 1609 4550
rect 1460 4516 1507 4540
rect 1086 4506 1507 4516
rect 1541 4506 1609 4540
rect 6335 4540 6370 4574
rect 6404 4540 6439 4574
rect 6473 4540 6508 4574
rect 6542 4540 6577 4574
rect 6611 4540 6646 4574
rect 6680 4540 6715 4574
rect 6749 4540 6784 4574
rect 6818 4540 6853 4574
rect 6887 4540 6922 4574
rect 6956 4540 6991 4574
rect 7025 4540 7060 4574
rect 7094 4540 7129 4574
rect 7163 4540 7198 4574
rect 7232 4540 7267 4574
rect 7301 4540 7336 4574
rect 7370 4540 7405 4574
rect 7439 4540 7474 4574
rect 7508 4540 7543 4574
rect 7577 4540 7612 4574
rect 7646 4540 7681 4574
rect 7715 4540 7750 4574
rect 7784 4540 7819 4574
rect 7853 4540 7888 4574
rect 7922 4540 7957 4574
rect 7991 4540 8026 4574
rect 8060 4540 8095 4574
rect 8129 4540 8164 4574
rect 8198 4540 8233 4574
rect 8267 4540 8302 4574
rect 8336 4540 8371 4574
rect 8405 4540 8440 4574
rect 8474 4540 8509 4574
rect 8543 4540 8578 4574
rect 8612 4540 8647 4574
rect 8681 4540 8716 4574
rect 8750 4540 8785 4574
rect 8819 4540 8854 4574
rect 8888 4540 8923 4574
rect 8957 4540 8992 4574
rect 9026 4540 9061 4574
rect 9095 4540 9130 4574
rect 9164 4540 9199 4574
rect 9233 4540 9268 4574
rect 9302 4540 9337 4574
rect 9371 4540 9406 4574
rect 9440 4540 9475 4574
rect 9509 4540 9544 4574
rect 9578 4540 9613 4574
rect 9647 4540 9682 4574
rect 9716 4540 9751 4574
rect 9785 4540 9820 4574
rect 9854 4540 9889 4574
rect 9923 4540 9958 4574
rect 9992 4540 10026 4574
rect 6335 4506 10026 4540
rect 1086 4481 1575 4506
rect 8681 4485 8716 4506
rect 1120 4447 1154 4481
rect 1188 4479 1222 4481
rect 1256 4479 1290 4481
rect 1324 4479 1358 4481
rect 1392 4479 1426 4481
rect 1460 4479 1575 4481
rect 1203 4447 1222 4479
rect 1275 4447 1290 4479
rect 1347 4447 1358 4479
rect 1419 4447 1426 4479
rect 1491 4471 1529 4479
rect 1563 4472 1575 4479
rect 1086 4445 1169 4447
rect 1203 4445 1241 4447
rect 1275 4445 1313 4447
rect 1347 4445 1385 4447
rect 1419 4445 1457 4447
rect 1491 4445 1507 4471
rect 1563 4445 1601 4472
rect 1635 4445 1643 4472
rect 8681 4451 8682 4485
rect 8750 4485 8785 4506
rect 8819 4485 8854 4506
rect 8888 4485 8923 4506
rect 8957 4485 8992 4506
rect 9026 4485 9061 4506
rect 9095 4485 9130 4506
rect 9164 4485 9199 4506
rect 9233 4485 9268 4506
rect 9302 4485 9337 4506
rect 9371 4485 9406 4506
rect 9440 4485 9475 4506
rect 8750 4472 8754 4485
rect 8819 4472 8826 4485
rect 8888 4472 8898 4485
rect 8957 4472 8970 4485
rect 9026 4472 9042 4485
rect 9095 4472 9114 4485
rect 9164 4472 9186 4485
rect 9233 4472 9258 4485
rect 9302 4472 9330 4485
rect 9371 4472 9402 4485
rect 9440 4472 9474 4485
rect 9509 4472 9544 4506
rect 9578 4485 9613 4506
rect 9647 4485 9682 4506
rect 9716 4485 9751 4506
rect 9785 4485 9820 4506
rect 9854 4485 9889 4506
rect 9923 4485 9958 4506
rect 9992 4485 10026 4506
rect 23568 4565 23597 4583
rect 23631 4565 23665 4599
rect 23699 4565 23733 4599
rect 23771 4583 23796 4617
rect 23767 4565 23796 4583
rect 23568 4544 23796 4565
rect 23568 4510 23593 4544
rect 23627 4530 23665 4544
rect 23699 4530 23737 4544
rect 23568 4496 23597 4510
rect 23631 4496 23665 4530
rect 23699 4496 23733 4530
rect 23771 4510 23796 4544
rect 23767 4496 23796 4510
rect 9580 4472 9613 4485
rect 9652 4472 9682 4485
rect 9724 4472 9751 4485
rect 9796 4472 9820 4485
rect 9868 4472 9889 4485
rect 9940 4472 9958 4485
rect 8716 4451 8754 4472
rect 8788 4451 8826 4472
rect 8860 4451 8898 4472
rect 8932 4451 8970 4472
rect 9004 4451 9042 4472
rect 9076 4451 9114 4472
rect 9148 4451 9186 4472
rect 9220 4451 9258 4472
rect 9292 4451 9330 4472
rect 9364 4451 9402 4472
rect 9436 4451 9474 4472
rect 9508 4451 9546 4472
rect 9580 4451 9618 4472
rect 9652 4451 9690 4472
rect 9724 4451 9762 4472
rect 9796 4451 9834 4472
rect 9868 4451 9906 4472
rect 9940 4451 9978 4472
rect 10012 4451 10050 4485
rect 10084 4451 10122 4485
rect 10156 4451 10194 4485
rect 10228 4451 10266 4485
rect 10300 4451 10338 4485
rect 10372 4451 10410 4485
rect 10444 4451 10482 4485
rect 10516 4451 10554 4485
rect 10588 4451 10626 4485
rect 10660 4451 10698 4485
rect 10732 4451 10770 4485
rect 10804 4451 10842 4485
rect 23568 4471 23796 4496
rect 1086 4437 1507 4445
rect 1541 4437 1643 4445
rect 1086 4436 1643 4437
rect 1086 4412 1575 4436
rect 1120 4378 1154 4412
rect 1188 4405 1222 4412
rect 1256 4405 1290 4412
rect 1324 4405 1358 4412
rect 1392 4405 1426 4412
rect 1460 4405 1575 4412
rect 1609 4405 1643 4436
rect 1203 4378 1222 4405
rect 1275 4378 1290 4405
rect 1347 4378 1358 4405
rect 1419 4378 1426 4405
rect 1491 4402 1529 4405
rect 1563 4402 1575 4405
rect 1635 4404 1643 4405
rect 8681 4438 10026 4451
rect 8681 4404 8716 4438
rect 8750 4404 8785 4438
rect 8819 4404 8854 4438
rect 8888 4404 8923 4438
rect 8957 4404 8992 4438
rect 9026 4404 9061 4438
rect 9095 4404 9130 4438
rect 9164 4404 9199 4438
rect 9233 4404 9268 4438
rect 9302 4404 9337 4438
rect 9371 4404 9406 4438
rect 9440 4404 9475 4438
rect 9509 4404 9544 4438
rect 9578 4404 9613 4438
rect 9647 4404 9682 4438
rect 9716 4404 9751 4438
rect 9785 4404 9820 4438
rect 9854 4404 9889 4438
rect 9923 4404 9958 4438
rect 9992 4405 10026 4438
rect 23568 4437 23593 4471
rect 23627 4461 23665 4471
rect 23699 4461 23737 4471
rect 23568 4427 23597 4437
rect 23631 4427 23665 4461
rect 23699 4427 23733 4461
rect 23771 4437 23796 4471
rect 23767 4427 23796 4437
rect 9992 4404 11589 4405
rect 1086 4371 1169 4378
rect 1203 4371 1241 4378
rect 1275 4371 1313 4378
rect 1347 4371 1385 4378
rect 1419 4371 1457 4378
rect 1491 4371 1507 4402
rect 1563 4371 1601 4402
rect 1635 4371 8643 4404
rect 1086 4368 1507 4371
rect 1541 4368 8643 4371
rect 1086 4366 1643 4368
rect 1086 4343 1575 4366
rect 1120 4309 1154 4343
rect 1188 4331 1222 4343
rect 1256 4331 1290 4343
rect 1324 4331 1358 4343
rect 1392 4331 1426 4343
rect 1460 4333 1575 4343
rect 1460 4331 1507 4333
rect 1541 4332 1575 4333
rect 1609 4334 1643 4366
rect 1677 4359 8643 4368
rect 1677 4334 1711 4359
rect 1609 4332 1711 4334
rect 1541 4331 1711 4332
rect 1203 4309 1222 4331
rect 1275 4309 1290 4331
rect 1347 4309 1358 4331
rect 1419 4309 1426 4331
rect 1086 4297 1169 4309
rect 1203 4297 1241 4309
rect 1275 4297 1313 4309
rect 1347 4297 1385 4309
rect 1419 4297 1457 4309
rect 1491 4299 1507 4331
rect 1491 4297 1529 4299
rect 1563 4297 1601 4331
rect 1635 4325 1711 4331
rect 1745 4325 1780 4359
rect 1814 4325 1849 4359
rect 1883 4325 1918 4359
rect 1952 4325 1987 4359
rect 2021 4325 2056 4359
rect 2090 4325 2125 4359
rect 2159 4325 2194 4359
rect 2228 4325 2263 4359
rect 2297 4325 2332 4359
rect 2366 4325 2401 4359
rect 1635 4298 2401 4325
rect 1635 4297 1643 4298
rect 1086 4296 1643 4297
rect 1086 4274 1575 4296
rect 1120 4240 1154 4274
rect 1188 4257 1222 4274
rect 1256 4257 1290 4274
rect 1324 4257 1358 4274
rect 1392 4257 1426 4274
rect 1460 4264 1575 4274
rect 1460 4257 1507 4264
rect 1541 4262 1575 4264
rect 1609 4264 1643 4296
rect 1677 4291 2401 4298
rect 1677 4264 1711 4291
rect 1609 4262 1711 4264
rect 1541 4257 1711 4262
rect 1745 4257 1780 4291
rect 1814 4257 1849 4291
rect 1883 4257 1918 4291
rect 1952 4257 1987 4291
rect 2021 4257 2056 4291
rect 2090 4257 2125 4291
rect 2159 4257 2194 4291
rect 2228 4257 2263 4291
rect 2297 4257 2332 4291
rect 2366 4257 2401 4291
rect 1203 4240 1222 4257
rect 1275 4240 1290 4257
rect 1347 4240 1358 4257
rect 1419 4240 1426 4257
rect 1086 4223 1169 4240
rect 1203 4223 1241 4240
rect 1275 4223 1313 4240
rect 1347 4223 1385 4240
rect 1419 4223 1457 4240
rect 1491 4230 1507 4257
rect 1491 4223 1529 4230
rect 1563 4226 1601 4257
rect 1635 4228 2401 4257
rect 1563 4223 1575 4226
rect 1635 4223 1643 4228
rect 1086 4205 1575 4223
rect 1120 4171 1154 4205
rect 1188 4183 1222 4205
rect 1256 4183 1290 4205
rect 1324 4183 1358 4205
rect 1392 4183 1426 4205
rect 1460 4195 1575 4205
rect 1460 4183 1507 4195
rect 1541 4192 1575 4195
rect 1609 4194 1643 4223
rect 1677 4223 2401 4228
rect 1677 4194 1711 4223
rect 1609 4192 1711 4194
rect 1541 4189 1711 4192
rect 1745 4189 1780 4223
rect 1814 4189 1849 4223
rect 1883 4189 1918 4223
rect 1952 4189 1987 4223
rect 2021 4189 2056 4223
rect 2090 4189 2125 4223
rect 2159 4189 2194 4223
rect 2228 4189 2263 4223
rect 2297 4189 2332 4223
rect 2366 4189 2401 4223
rect 4135 4336 8643 4359
rect 8681 4371 11589 4404
rect 23568 4398 23796 4427
rect 8681 4370 10312 4371
rect 8681 4336 8711 4370
rect 8745 4336 8779 4370
rect 8813 4336 8847 4370
rect 8881 4336 8915 4370
rect 8949 4336 8983 4370
rect 9017 4336 9051 4370
rect 9085 4336 9119 4370
rect 9153 4336 9187 4370
rect 9221 4336 9255 4370
rect 9289 4336 9323 4370
rect 9357 4336 9391 4370
rect 9425 4336 9459 4370
rect 9493 4336 9527 4370
rect 9561 4336 9595 4370
rect 9629 4336 9663 4370
rect 9697 4336 9731 4370
rect 9765 4336 9799 4370
rect 9833 4336 9867 4370
rect 9901 4336 9935 4370
rect 9969 4336 10003 4370
rect 10037 4336 10071 4370
rect 10105 4336 10139 4370
rect 10173 4336 10207 4370
rect 10241 4337 10312 4370
rect 10346 4337 10380 4371
rect 10414 4337 10448 4371
rect 10482 4337 10516 4371
rect 10550 4337 10584 4371
rect 10618 4337 10652 4371
rect 10686 4337 10720 4371
rect 10754 4337 10788 4371
rect 10822 4337 10856 4371
rect 10890 4337 10924 4371
rect 10958 4337 10992 4371
rect 11026 4337 11060 4371
rect 11094 4337 11128 4371
rect 11162 4337 11196 4371
rect 11230 4337 11264 4371
rect 11298 4337 11332 4371
rect 11366 4337 11400 4371
rect 11434 4337 11468 4371
rect 11502 4337 11536 4371
rect 11570 4337 11589 4371
rect 10241 4336 11589 4337
rect 4135 4334 11589 4336
rect 4135 4300 4179 4334
rect 4213 4300 4248 4334
rect 4282 4300 4317 4334
rect 4351 4300 4386 4334
rect 4420 4300 4455 4334
rect 4489 4300 4524 4334
rect 4558 4300 4593 4334
rect 4627 4300 4662 4334
rect 4696 4300 4731 4334
rect 4765 4300 4800 4334
rect 4834 4300 4869 4334
rect 4903 4300 4938 4334
rect 4972 4300 5007 4334
rect 5041 4300 5076 4334
rect 5110 4300 5145 4334
rect 5179 4300 5214 4334
rect 5248 4300 5283 4334
rect 5317 4300 5352 4334
rect 5386 4300 5421 4334
rect 5455 4300 5490 4334
rect 4135 4266 5490 4300
rect 4135 4232 4179 4266
rect 4213 4232 4248 4266
rect 4282 4232 4317 4266
rect 4351 4232 4386 4266
rect 4420 4232 4455 4266
rect 4489 4232 4524 4266
rect 4558 4232 4593 4266
rect 4627 4232 4662 4266
rect 4696 4232 4731 4266
rect 4765 4232 4800 4266
rect 4834 4232 4869 4266
rect 4903 4232 4938 4266
rect 4972 4232 5007 4266
rect 5041 4232 5076 4266
rect 5110 4232 5145 4266
rect 5179 4232 5214 4266
rect 5248 4232 5283 4266
rect 5317 4232 5352 4266
rect 5386 4232 5421 4266
rect 5455 4232 5490 4266
rect 4135 4198 5490 4232
rect 4135 4189 4179 4198
rect 1541 4183 1677 4189
rect 1203 4171 1222 4183
rect 1275 4171 1290 4183
rect 1347 4171 1358 4183
rect 1419 4171 1426 4183
rect 1086 4149 1169 4171
rect 1203 4149 1241 4171
rect 1275 4149 1313 4171
rect 1347 4149 1385 4171
rect 1419 4149 1457 4171
rect 1491 4161 1507 4183
rect 1491 4149 1529 4161
rect 1563 4156 1601 4183
rect 1635 4158 1677 4183
rect 1563 4149 1575 4156
rect 1635 4149 1643 4158
rect 1086 4136 1575 4149
rect 1120 4102 1154 4136
rect 1188 4109 1222 4136
rect 1256 4109 1290 4136
rect 1324 4109 1358 4136
rect 1392 4109 1426 4136
rect 1460 4126 1575 4136
rect 1460 4109 1507 4126
rect 1541 4122 1575 4126
rect 1609 4124 1643 4149
rect 1609 4122 1677 4124
rect 1541 4109 1677 4122
rect 1203 4102 1222 4109
rect 1275 4102 1290 4109
rect 1347 4102 1358 4109
rect 1419 4102 1426 4109
rect 1086 4075 1169 4102
rect 1203 4075 1241 4102
rect 1275 4075 1313 4102
rect 1347 4075 1385 4102
rect 1419 4075 1457 4102
rect 1491 4092 1507 4109
rect 1491 4075 1529 4092
rect 1563 4086 1601 4109
rect 1635 4088 1677 4109
rect 1563 4075 1575 4086
rect 1635 4075 1643 4088
rect 1086 4067 1575 4075
rect 1120 4033 1154 4067
rect 1188 4035 1222 4067
rect 1256 4035 1290 4067
rect 1324 4035 1358 4067
rect 1392 4035 1426 4067
rect 1460 4057 1575 4067
rect 1460 4035 1507 4057
rect 1541 4052 1575 4057
rect 1609 4054 1643 4075
rect 4155 4164 4179 4189
rect 4213 4164 4248 4198
rect 4282 4164 4317 4198
rect 4351 4164 4386 4198
rect 4420 4164 4455 4198
rect 4489 4164 4524 4198
rect 4558 4164 4593 4198
rect 4627 4164 4662 4198
rect 4696 4164 4731 4198
rect 4765 4164 4800 4198
rect 4834 4164 4869 4198
rect 4903 4164 4938 4198
rect 4972 4164 5007 4198
rect 5041 4164 5076 4198
rect 5110 4164 5145 4198
rect 5179 4164 5214 4198
rect 5248 4164 5283 4198
rect 5317 4164 5352 4198
rect 5386 4164 5421 4198
rect 5455 4164 5490 4198
rect 4155 4130 5490 4164
rect 4155 4096 4179 4130
rect 4213 4096 4248 4130
rect 4282 4096 4317 4130
rect 4351 4096 4386 4130
rect 4420 4096 4455 4130
rect 4489 4096 4524 4130
rect 4558 4096 4593 4130
rect 4627 4096 4662 4130
rect 4696 4096 4731 4130
rect 4765 4096 4800 4130
rect 4834 4096 4869 4130
rect 4903 4096 4938 4130
rect 4972 4096 5007 4130
rect 5041 4096 5076 4130
rect 5110 4096 5145 4130
rect 5179 4096 5214 4130
rect 5248 4096 5283 4130
rect 5317 4096 5352 4130
rect 5386 4096 5421 4130
rect 5455 4096 5490 4130
rect 1677 4060 1904 4076
rect 1677 4054 1802 4060
rect 1609 4052 1802 4054
rect 1541 4035 1802 4052
rect 1203 4033 1222 4035
rect 1275 4033 1290 4035
rect 1347 4033 1358 4035
rect 1419 4033 1426 4035
rect 1086 4001 1169 4033
rect 1203 4001 1241 4033
rect 1275 4001 1313 4033
rect 1347 4001 1385 4033
rect 1419 4001 1457 4033
rect 1491 4023 1507 4035
rect 1491 4001 1529 4023
rect 1563 4016 1601 4035
rect 1635 4026 1802 4035
rect 1836 4026 1870 4060
rect 1635 4018 1904 4026
rect 1563 4001 1575 4016
rect 1635 4001 1643 4018
rect 1086 3998 1575 4001
rect 1120 3964 1154 3998
rect 1188 3964 1222 3998
rect 1256 3964 1290 3998
rect 1324 3964 1358 3998
rect 1392 3964 1426 3998
rect 1460 3988 1575 3998
rect 1460 3964 1507 3988
rect 1086 3962 1507 3964
rect 1541 3982 1575 3988
rect 1609 3984 1643 4001
rect 1677 4010 1904 4018
rect 3944 4060 4046 4076
rect 4155 4062 5490 4096
rect 3980 4026 4012 4060
rect 4155 4028 4179 4062
rect 4213 4028 4248 4062
rect 4282 4028 4317 4062
rect 4351 4028 4386 4062
rect 4420 4028 4455 4062
rect 4489 4028 4524 4062
rect 4558 4028 4593 4062
rect 4627 4028 4662 4062
rect 4696 4028 4731 4062
rect 4765 4028 4800 4062
rect 4834 4028 4869 4062
rect 4903 4028 4938 4062
rect 4972 4028 5007 4062
rect 5041 4028 5076 4062
rect 5110 4028 5145 4062
rect 5179 4028 5214 4062
rect 5248 4028 5283 4062
rect 5317 4028 5352 4062
rect 5386 4028 5421 4062
rect 5455 4028 5490 4062
rect 3944 4010 4046 4026
rect 1609 3982 1677 3984
rect 1541 3962 1677 3982
rect 1086 3929 1169 3962
rect 1203 3929 1241 3962
rect 1275 3929 1313 3962
rect 1347 3929 1385 3962
rect 1419 3929 1457 3962
rect 1491 3954 1507 3962
rect 1120 3895 1154 3929
rect 1203 3928 1222 3929
rect 1275 3928 1290 3929
rect 1347 3928 1358 3929
rect 1419 3928 1426 3929
rect 1491 3928 1529 3954
rect 1563 3946 1601 3962
rect 1635 3948 1677 3962
rect 1563 3928 1575 3946
rect 1635 3928 1643 3948
rect 1188 3895 1222 3928
rect 1256 3895 1290 3928
rect 1324 3895 1358 3928
rect 1392 3895 1426 3928
rect 1460 3919 1575 3928
rect 1460 3895 1507 3919
rect 1086 3889 1507 3895
rect 1541 3912 1575 3919
rect 1609 3914 1643 3928
rect 1609 3912 1677 3914
rect 1541 3889 1677 3912
rect 1086 3860 1169 3889
rect 1203 3860 1241 3889
rect 1275 3860 1313 3889
rect 1347 3860 1385 3889
rect 1419 3860 1457 3889
rect 1491 3885 1507 3889
rect 1120 3826 1154 3860
rect 1203 3855 1222 3860
rect 1275 3855 1290 3860
rect 1347 3855 1358 3860
rect 1419 3855 1426 3860
rect 1491 3855 1529 3885
rect 1563 3876 1601 3889
rect 1635 3878 1677 3889
rect 1563 3855 1575 3876
rect 1635 3855 1643 3878
rect 1188 3826 1222 3855
rect 1256 3826 1290 3855
rect 1324 3826 1358 3855
rect 1392 3826 1426 3855
rect 1460 3850 1575 3855
rect 1460 3826 1507 3850
rect 1086 3816 1507 3826
rect 1541 3842 1575 3850
rect 1609 3844 1643 3855
rect 4155 3994 5490 4028
rect 4155 3960 4179 3994
rect 4213 3960 4248 3994
rect 4282 3960 4317 3994
rect 4351 3960 4386 3994
rect 4420 3960 4455 3994
rect 4489 3960 4524 3994
rect 4558 3960 4593 3994
rect 4627 3960 4662 3994
rect 4696 3960 4731 3994
rect 4765 3960 4800 3994
rect 4834 3960 4869 3994
rect 4903 3960 4938 3994
rect 4972 3960 5007 3994
rect 5041 3960 5076 3994
rect 5110 3960 5145 3994
rect 5179 3960 5214 3994
rect 5248 3960 5283 3994
rect 5317 3960 5352 3994
rect 5386 3960 5421 3994
rect 5455 3960 5490 3994
rect 4155 3926 5490 3960
rect 4155 3892 4179 3926
rect 4213 3892 4248 3926
rect 4282 3892 4317 3926
rect 4351 3892 4386 3926
rect 4420 3892 4455 3926
rect 4489 3892 4524 3926
rect 4558 3892 4593 3926
rect 4627 3892 4662 3926
rect 4696 3892 4731 3926
rect 4765 3892 4800 3926
rect 4834 3892 4869 3926
rect 4903 3892 4938 3926
rect 4972 3892 5007 3926
rect 5041 3892 5076 3926
rect 5110 3892 5145 3926
rect 5179 3892 5214 3926
rect 5248 3892 5283 3926
rect 5317 3892 5352 3926
rect 5386 3892 5421 3926
rect 5455 3892 5490 3926
rect 8584 4301 11589 4334
rect 8584 4300 10312 4301
rect 8584 4266 8643 4300
rect 8677 4266 8711 4300
rect 8745 4266 8779 4300
rect 8813 4266 8847 4300
rect 8881 4266 8915 4300
rect 8949 4266 8983 4300
rect 9017 4266 9051 4300
rect 9085 4266 9119 4300
rect 9153 4266 9187 4300
rect 9221 4266 9255 4300
rect 9289 4266 9323 4300
rect 9357 4266 9391 4300
rect 9425 4266 9459 4300
rect 9493 4266 9527 4300
rect 9561 4266 9595 4300
rect 9629 4266 9663 4300
rect 9697 4266 9731 4300
rect 9765 4266 9799 4300
rect 9833 4266 9867 4300
rect 9901 4266 9935 4300
rect 9969 4266 10003 4300
rect 10037 4266 10071 4300
rect 10105 4266 10139 4300
rect 10173 4266 10207 4300
rect 10241 4267 10312 4300
rect 10346 4267 10380 4301
rect 10414 4267 10448 4301
rect 10482 4267 10516 4301
rect 10550 4267 10584 4301
rect 10618 4267 10652 4301
rect 10686 4267 10720 4301
rect 10754 4267 10788 4301
rect 10822 4267 10856 4301
rect 10890 4267 10924 4301
rect 10958 4267 10992 4301
rect 11026 4267 11060 4301
rect 11094 4267 11128 4301
rect 11162 4267 11196 4301
rect 11230 4267 11264 4301
rect 11298 4267 11332 4301
rect 11366 4267 11400 4301
rect 11434 4267 11468 4301
rect 11502 4267 11536 4301
rect 11570 4267 11589 4301
rect 10241 4266 11589 4267
rect 8584 4231 11589 4266
rect 8584 4230 10312 4231
rect 8584 4196 8643 4230
rect 8677 4196 8711 4230
rect 8745 4196 8779 4230
rect 8813 4196 8847 4230
rect 8881 4196 8915 4230
rect 8949 4196 8983 4230
rect 9017 4196 9051 4230
rect 9085 4196 9119 4230
rect 9153 4196 9187 4230
rect 9221 4196 9255 4230
rect 9289 4196 9323 4230
rect 9357 4196 9391 4230
rect 9425 4196 9459 4230
rect 9493 4196 9527 4230
rect 9561 4196 9595 4230
rect 9629 4196 9663 4230
rect 9697 4196 9731 4230
rect 9765 4196 9799 4230
rect 9833 4196 9867 4230
rect 9901 4196 9935 4230
rect 9969 4196 10003 4230
rect 10037 4196 10071 4230
rect 10105 4196 10139 4230
rect 10173 4196 10207 4230
rect 10241 4197 10312 4230
rect 10346 4197 10380 4231
rect 10414 4197 10448 4231
rect 10482 4197 10516 4231
rect 10550 4197 10584 4231
rect 10618 4197 10652 4231
rect 10686 4197 10720 4231
rect 10754 4197 10788 4231
rect 10822 4197 10856 4231
rect 10890 4197 10924 4231
rect 10958 4197 10992 4231
rect 11026 4197 11060 4231
rect 11094 4197 11128 4231
rect 11162 4197 11196 4231
rect 11230 4197 11264 4231
rect 11298 4197 11332 4231
rect 11366 4197 11400 4231
rect 11434 4197 11468 4231
rect 11502 4197 11536 4231
rect 11570 4197 11589 4231
rect 10241 4196 11589 4197
rect 8584 4161 11589 4196
rect 8584 4160 10312 4161
rect 8584 4126 8643 4160
rect 8677 4126 8711 4160
rect 8745 4126 8779 4160
rect 8813 4126 8847 4160
rect 8881 4126 8915 4160
rect 8949 4126 8983 4160
rect 9017 4126 9051 4160
rect 9085 4126 9119 4160
rect 9153 4126 9187 4160
rect 9221 4126 9255 4160
rect 9289 4126 9323 4160
rect 9357 4126 9391 4160
rect 9425 4126 9459 4160
rect 9493 4126 9527 4160
rect 9561 4126 9595 4160
rect 9629 4126 9663 4160
rect 9697 4126 9731 4160
rect 9765 4126 9799 4160
rect 9833 4126 9867 4160
rect 9901 4126 9935 4160
rect 9969 4126 10003 4160
rect 10037 4126 10071 4160
rect 10105 4126 10139 4160
rect 10173 4126 10207 4160
rect 10241 4127 10312 4160
rect 10346 4127 10380 4161
rect 10414 4127 10448 4161
rect 10482 4127 10516 4161
rect 10550 4127 10584 4161
rect 10618 4127 10652 4161
rect 10686 4127 10720 4161
rect 10754 4127 10788 4161
rect 10822 4127 10856 4161
rect 10890 4127 10924 4161
rect 10958 4127 10992 4161
rect 11026 4127 11060 4161
rect 11094 4127 11128 4161
rect 11162 4127 11196 4161
rect 11230 4127 11264 4161
rect 11298 4127 11332 4161
rect 11366 4127 11400 4161
rect 11434 4127 11468 4161
rect 11502 4127 11536 4161
rect 11570 4127 11589 4161
rect 10241 4126 11589 4127
rect 8584 4091 11589 4126
rect 8584 4090 10312 4091
rect 8584 4056 8643 4090
rect 8677 4056 8711 4090
rect 8745 4056 8779 4090
rect 8813 4056 8847 4090
rect 8881 4056 8915 4090
rect 8949 4056 8983 4090
rect 9017 4056 9051 4090
rect 9085 4056 9119 4090
rect 9153 4056 9187 4090
rect 9221 4056 9255 4090
rect 9289 4056 9323 4090
rect 9357 4056 9391 4090
rect 9425 4056 9459 4090
rect 9493 4056 9527 4090
rect 9561 4056 9595 4090
rect 9629 4056 9663 4090
rect 9697 4056 9731 4090
rect 9765 4056 9799 4090
rect 9833 4056 9867 4090
rect 9901 4056 9935 4090
rect 9969 4056 10003 4090
rect 10037 4056 10071 4090
rect 10105 4056 10139 4090
rect 10173 4056 10207 4090
rect 10241 4057 10312 4090
rect 10346 4057 10380 4091
rect 10414 4057 10448 4091
rect 10482 4057 10516 4091
rect 10550 4057 10584 4091
rect 10618 4057 10652 4091
rect 10686 4057 10720 4091
rect 10754 4057 10788 4091
rect 10822 4057 10856 4091
rect 10890 4057 10924 4091
rect 10958 4057 10992 4091
rect 11026 4057 11060 4091
rect 11094 4057 11128 4091
rect 11162 4057 11196 4091
rect 11230 4057 11264 4091
rect 11298 4057 11332 4091
rect 11366 4057 11400 4091
rect 11434 4057 11468 4091
rect 11502 4057 11536 4091
rect 11570 4057 11589 4091
rect 10241 4056 11589 4057
rect 8584 4021 11589 4056
rect 8584 4020 10312 4021
rect 8584 3986 8643 4020
rect 8677 3986 8711 4020
rect 8745 3986 8779 4020
rect 8813 3986 8847 4020
rect 8881 3986 8915 4020
rect 8949 3986 8983 4020
rect 9017 3986 9051 4020
rect 9085 3986 9119 4020
rect 9153 3986 9187 4020
rect 9221 3986 9255 4020
rect 9289 3986 9323 4020
rect 9357 3986 9391 4020
rect 9425 3986 9459 4020
rect 9493 3986 9527 4020
rect 9561 3986 9595 4020
rect 9629 3986 9663 4020
rect 9697 3986 9731 4020
rect 9765 3986 9799 4020
rect 9833 3986 9867 4020
rect 9901 3986 9935 4020
rect 9969 3986 10003 4020
rect 10037 3986 10071 4020
rect 10105 3986 10139 4020
rect 10173 3986 10207 4020
rect 10241 3987 10312 4020
rect 10346 3987 10380 4021
rect 10414 3987 10448 4021
rect 10482 3987 10516 4021
rect 10550 3987 10584 4021
rect 10618 3987 10652 4021
rect 10686 3987 10720 4021
rect 10754 3987 10788 4021
rect 10822 3987 10856 4021
rect 10890 3987 10924 4021
rect 10958 3987 10992 4021
rect 11026 3987 11060 4021
rect 11094 3987 11128 4021
rect 11162 3987 11196 4021
rect 11230 3987 11264 4021
rect 11298 3987 11332 4021
rect 11366 3987 11400 4021
rect 11434 3987 11468 4021
rect 11502 3987 11536 4021
rect 11570 3987 11589 4021
rect 10241 3986 11589 3987
rect 8584 3951 11589 3986
rect 8584 3950 10312 3951
rect 8584 3916 8643 3950
rect 8677 3916 8711 3950
rect 8745 3916 8779 3950
rect 8813 3916 8847 3950
rect 8881 3916 8915 3950
rect 8949 3916 8983 3950
rect 9017 3916 9051 3950
rect 9085 3916 9119 3950
rect 9153 3916 9187 3950
rect 9221 3916 9255 3950
rect 9289 3916 9323 3950
rect 9357 3916 9391 3950
rect 9425 3916 9459 3950
rect 9493 3916 9527 3950
rect 9561 3916 9595 3950
rect 9629 3916 9663 3950
rect 9697 3916 9731 3950
rect 9765 3916 9799 3950
rect 9833 3916 9867 3950
rect 9901 3916 9935 3950
rect 9969 3916 10003 3950
rect 10037 3916 10071 3950
rect 10105 3916 10139 3950
rect 10173 3916 10207 3950
rect 10241 3917 10312 3950
rect 10346 3917 10380 3951
rect 10414 3917 10448 3951
rect 10482 3917 10516 3951
rect 10550 3917 10584 3951
rect 10618 3917 10652 3951
rect 10686 3917 10720 3951
rect 10754 3917 10788 3951
rect 10822 3917 10856 3951
rect 10890 3917 10924 3951
rect 10958 3917 10992 3951
rect 11026 3917 11060 3951
rect 11094 3917 11128 3951
rect 11162 3917 11196 3951
rect 11230 3917 11264 3951
rect 11298 3917 11332 3951
rect 11366 3917 11400 3951
rect 11434 3917 11468 3951
rect 11502 3917 11536 3951
rect 11570 3917 11589 3951
rect 10241 3916 11589 3917
rect 8584 3892 11589 3916
rect 4155 3881 11589 3892
rect 4155 3880 10312 3881
rect 4155 3867 8643 3880
rect 1609 3842 1677 3844
rect 1541 3816 1677 3842
rect 1086 3791 1169 3816
rect 1203 3791 1241 3816
rect 1275 3791 1313 3816
rect 1347 3791 1385 3816
rect 1419 3791 1457 3816
rect 1120 3757 1154 3791
rect 1203 3782 1222 3791
rect 1275 3782 1290 3791
rect 1347 3782 1358 3791
rect 1419 3782 1426 3791
rect 1491 3782 1529 3816
rect 1563 3806 1601 3816
rect 1635 3808 1677 3816
rect 1563 3782 1575 3806
rect 1635 3782 1643 3808
rect 1188 3757 1222 3782
rect 1256 3757 1290 3782
rect 1324 3757 1358 3782
rect 1392 3757 1426 3782
rect 1460 3781 1575 3782
rect 1460 3757 1507 3781
rect 1086 3747 1507 3757
rect 1541 3772 1575 3781
rect 1609 3774 1643 3782
rect 1609 3772 1677 3774
rect 1541 3747 1677 3772
rect 1086 3743 1677 3747
rect 1086 3722 1169 3743
rect 1203 3722 1241 3743
rect 1275 3722 1313 3743
rect 1347 3722 1385 3743
rect 1419 3722 1457 3743
rect 1120 3688 1154 3722
rect 1203 3709 1222 3722
rect 1275 3709 1290 3722
rect 1347 3709 1358 3722
rect 1419 3709 1426 3722
rect 1491 3712 1529 3743
rect 1563 3736 1601 3743
rect 1635 3738 1677 3743
rect 1491 3709 1507 3712
rect 1563 3709 1575 3736
rect 1635 3709 1643 3738
rect 1188 3688 1222 3709
rect 1256 3688 1290 3709
rect 1324 3688 1358 3709
rect 1392 3688 1426 3709
rect 1460 3688 1507 3709
rect 1086 3678 1507 3688
rect 1541 3702 1575 3709
rect 1609 3704 1643 3709
rect 1609 3702 1677 3704
rect 1541 3678 1677 3702
rect 1086 3670 1677 3678
rect 1086 3653 1169 3670
rect 1203 3653 1241 3670
rect 1275 3653 1313 3670
rect 1347 3653 1385 3670
rect 1419 3653 1457 3670
rect 1491 3643 1529 3670
rect 1563 3666 1601 3670
rect 1635 3668 1677 3670
rect 1491 3636 1507 3643
rect 1563 3636 1575 3666
rect 1635 3636 1643 3668
rect 1460 3609 1507 3636
rect 1541 3632 1575 3636
rect 1609 3634 1643 3636
rect 8677 3846 8711 3880
rect 8745 3846 8779 3880
rect 8813 3846 8847 3880
rect 8881 3846 8915 3880
rect 8949 3846 8983 3880
rect 9017 3846 9051 3880
rect 9085 3846 9119 3880
rect 9153 3846 9187 3880
rect 9221 3846 9255 3880
rect 9289 3846 9323 3880
rect 9357 3846 9391 3880
rect 9425 3846 9459 3880
rect 9493 3846 9527 3880
rect 9561 3846 9595 3880
rect 9629 3846 9663 3880
rect 9697 3846 9731 3880
rect 9765 3846 9799 3880
rect 9833 3846 9867 3880
rect 9901 3846 9935 3880
rect 9969 3846 10003 3880
rect 10037 3846 10071 3880
rect 10105 3846 10139 3880
rect 10173 3846 10207 3880
rect 10241 3847 10312 3880
rect 10346 3847 10380 3881
rect 10414 3847 10448 3881
rect 10482 3847 10516 3881
rect 10550 3847 10584 3881
rect 10618 3847 10652 3881
rect 10686 3847 10720 3881
rect 10754 3847 10788 3881
rect 10822 3847 10856 3881
rect 10890 3847 10924 3881
rect 10958 3847 10992 3881
rect 11026 3847 11060 3881
rect 11094 3847 11128 3881
rect 11162 3847 11196 3881
rect 11230 3847 11264 3881
rect 11298 3847 11332 3881
rect 11366 3847 11400 3881
rect 11434 3847 11468 3881
rect 11502 3847 11536 3881
rect 11570 3847 11589 3881
rect 10241 3846 11589 3847
rect 8643 3811 11589 3846
rect 8643 3810 10312 3811
rect 8677 3776 8711 3810
rect 8745 3776 8779 3810
rect 8813 3776 8847 3810
rect 8881 3776 8915 3810
rect 8949 3776 8983 3810
rect 9017 3776 9051 3810
rect 9085 3776 9119 3810
rect 9153 3776 9187 3810
rect 9221 3776 9255 3810
rect 9289 3776 9323 3810
rect 9357 3776 9391 3810
rect 9425 3776 9459 3810
rect 9493 3776 9527 3810
rect 9561 3776 9595 3810
rect 9629 3776 9663 3810
rect 9697 3776 9731 3810
rect 9765 3776 9799 3810
rect 9833 3776 9867 3810
rect 9901 3776 9935 3810
rect 9969 3776 10003 3810
rect 10037 3776 10071 3810
rect 10105 3776 10139 3810
rect 10173 3776 10207 3810
rect 10241 3777 10312 3810
rect 10346 3777 10380 3811
rect 10414 3777 10448 3811
rect 10482 3777 10516 3811
rect 10550 3777 10584 3811
rect 10618 3777 10652 3811
rect 10686 3777 10720 3811
rect 10754 3777 10788 3811
rect 10822 3777 10856 3811
rect 10890 3777 10924 3811
rect 10958 3777 10992 3811
rect 11026 3777 11060 3811
rect 11094 3777 11128 3811
rect 11162 3777 11196 3811
rect 11230 3777 11264 3811
rect 11298 3777 11332 3811
rect 11366 3777 11400 3811
rect 11434 3777 11468 3811
rect 11502 3777 11536 3811
rect 11570 3777 11589 3811
rect 10241 3776 11589 3777
rect 8643 3741 11589 3776
rect 8643 3740 10312 3741
rect 8677 3706 8711 3740
rect 8745 3706 8779 3740
rect 8813 3706 8847 3740
rect 8881 3706 8915 3740
rect 8949 3706 8983 3740
rect 9017 3706 9051 3740
rect 9085 3706 9119 3740
rect 9153 3706 9187 3740
rect 9221 3706 9255 3740
rect 9289 3706 9323 3740
rect 9357 3706 9391 3740
rect 9425 3706 9459 3740
rect 9493 3706 9527 3740
rect 9561 3706 9595 3740
rect 9629 3706 9663 3740
rect 9697 3706 9731 3740
rect 9765 3706 9799 3740
rect 9833 3706 9867 3740
rect 9901 3706 9935 3740
rect 9969 3706 10003 3740
rect 10037 3706 10071 3740
rect 10105 3706 10139 3740
rect 10173 3706 10207 3740
rect 10241 3707 10312 3740
rect 10346 3707 10380 3741
rect 10414 3707 10448 3741
rect 10482 3707 10516 3741
rect 10550 3707 10584 3741
rect 10618 3707 10652 3741
rect 10686 3707 10720 3741
rect 10754 3707 10788 3741
rect 10822 3707 10856 3741
rect 10890 3707 10924 3741
rect 10958 3707 10992 3741
rect 11026 3707 11060 3741
rect 11094 3707 11128 3741
rect 11162 3707 11196 3741
rect 11230 3707 11264 3741
rect 11298 3707 11332 3741
rect 11366 3707 11400 3741
rect 11434 3707 11468 3741
rect 11502 3707 11536 3741
rect 11570 3707 11589 3741
rect 10241 3706 11589 3707
rect 8643 3671 11589 3706
rect 8643 3670 10312 3671
rect 1609 3632 1677 3634
rect 1541 3609 1677 3632
rect 1460 3598 1677 3609
rect 1460 3597 1643 3598
rect 1491 3574 1529 3597
rect 1563 3596 1601 3597
rect 1491 3563 1507 3574
rect 1563 3563 1575 3596
rect 1635 3564 1643 3597
rect 1635 3563 1677 3564
rect 1460 3540 1507 3563
rect 1541 3562 1575 3563
rect 1609 3562 1677 3563
rect 1541 3540 1677 3562
rect 1460 3528 1677 3540
rect 1460 3526 1643 3528
rect 1460 3524 1575 3526
rect 1609 3524 1643 3526
rect 1491 3505 1529 3524
rect 1491 3490 1507 3505
rect 1563 3492 1575 3524
rect 1635 3494 1643 3524
rect 1563 3490 1601 3492
rect 1635 3490 1677 3494
rect 1460 3471 1507 3490
rect 1541 3471 1677 3490
rect 1460 3458 1677 3471
rect 1460 3456 1643 3458
rect 1460 3451 1575 3456
rect 1609 3451 1643 3456
rect 1491 3436 1529 3451
rect 1491 3417 1507 3436
rect 1563 3422 1575 3451
rect 1635 3424 1643 3451
rect 1563 3417 1601 3422
rect 1635 3417 1677 3424
rect 1460 3402 1507 3417
rect 1541 3402 1677 3417
rect 1460 3388 1677 3402
rect 1460 3386 1643 3388
rect 1460 3378 1575 3386
rect 1609 3378 1643 3386
rect 1491 3367 1529 3378
rect 1491 3344 1507 3367
rect 1563 3352 1575 3378
rect 1635 3354 1643 3378
rect 1563 3344 1601 3352
rect 1635 3344 1677 3354
rect 1460 3333 1507 3344
rect 1541 3333 1677 3344
rect 1460 3318 1677 3333
rect 1460 3316 1643 3318
rect 1460 3305 1575 3316
rect 1609 3305 1643 3316
rect 1491 3298 1529 3305
rect 1491 3271 1507 3298
rect 1563 3282 1575 3305
rect 1635 3284 1643 3305
rect 1563 3271 1601 3282
rect 1635 3271 1677 3284
rect 1460 3264 1507 3271
rect 1541 3264 1677 3271
rect 1460 3258 1677 3264
rect 4998 3413 5104 3647
rect 8472 3413 8609 3647
rect 1460 3248 1740 3258
rect 1460 3246 1643 3248
rect 1460 3232 1575 3246
rect 1609 3232 1643 3246
rect 1491 3229 1529 3232
rect 1491 3198 1507 3229
rect 1563 3212 1575 3232
rect 1635 3214 1643 3232
rect 1677 3228 1740 3248
rect 1774 3228 1809 3258
rect 1843 3228 1878 3258
rect 1912 3228 1947 3258
rect 1981 3228 2016 3258
rect 2050 3228 2085 3258
rect 2119 3228 2154 3258
rect 1677 3214 1712 3228
rect 1774 3224 1785 3228
rect 1843 3224 1858 3228
rect 1912 3224 1931 3228
rect 1981 3224 2004 3228
rect 2050 3224 2077 3228
rect 2119 3224 2150 3228
rect 2188 3224 2223 3258
rect 2257 3224 2292 3258
rect 2326 3228 2361 3258
rect 2395 3228 2430 3258
rect 2464 3228 2499 3258
rect 2533 3228 2568 3258
rect 2602 3228 2637 3258
rect 2671 3228 2706 3258
rect 2740 3228 2775 3258
rect 2809 3228 2844 3258
rect 2330 3224 2361 3228
rect 2403 3224 2430 3228
rect 2476 3224 2499 3228
rect 2549 3224 2568 3228
rect 2622 3224 2637 3228
rect 2695 3224 2706 3228
rect 2768 3224 2775 3228
rect 1563 3198 1601 3212
rect 1635 3198 1712 3214
rect 1460 3195 1507 3198
rect 1541 3195 1712 3198
rect 1460 3194 1712 3195
rect 1746 3194 1785 3224
rect 1819 3194 1858 3224
rect 1892 3194 1931 3224
rect 1965 3194 2004 3224
rect 2038 3194 2077 3224
rect 2111 3194 2150 3224
rect 2184 3194 2223 3224
rect 2257 3194 2296 3224
rect 2330 3194 2369 3224
rect 2403 3194 2442 3224
rect 2476 3194 2515 3224
rect 2549 3194 2588 3224
rect 2622 3194 2661 3224
rect 2695 3194 2734 3224
rect 2768 3194 2807 3224
rect 1460 3190 2807 3194
rect 1460 3178 1740 3190
rect 1460 3176 1643 3178
rect 1460 3160 1575 3176
rect 1460 3159 1507 3160
rect 1541 3159 1575 3160
rect 1609 3159 1643 3176
rect 1491 3126 1507 3159
rect 1563 3142 1575 3159
rect 1635 3144 1643 3159
rect 1677 3156 1740 3178
rect 1774 3156 1809 3190
rect 1843 3156 1878 3190
rect 1912 3156 1947 3190
rect 1981 3156 2016 3190
rect 2050 3156 2085 3190
rect 2119 3156 2154 3190
rect 2188 3156 2223 3190
rect 2257 3156 2292 3190
rect 2326 3156 2361 3190
rect 2395 3156 2430 3190
rect 2464 3156 2499 3190
rect 2533 3156 2568 3190
rect 2602 3156 2637 3190
rect 2671 3156 2706 3190
rect 2740 3156 2775 3190
rect 1677 3144 1712 3156
rect 1491 3125 1529 3126
rect 1563 3125 1601 3142
rect 1635 3125 1712 3144
rect 1460 3122 1712 3125
rect 1746 3122 1785 3156
rect 1819 3122 1858 3156
rect 1892 3122 1931 3156
rect 1965 3122 2004 3156
rect 2038 3122 2077 3156
rect 2111 3122 2150 3156
rect 2184 3122 2223 3156
rect 2257 3122 2296 3156
rect 2330 3122 2369 3156
rect 2403 3122 2442 3156
rect 2476 3122 2515 3156
rect 2549 3122 2588 3156
rect 2622 3122 2661 3156
rect 2695 3122 2734 3156
rect 2768 3122 2807 3156
rect 1460 3108 1740 3122
rect 1460 3107 1643 3108
rect 1460 3091 1575 3107
rect 1460 3086 1507 3091
rect 1541 3086 1575 3091
rect 1609 3086 1643 3107
rect 1491 3057 1507 3086
rect 1563 3073 1575 3086
rect 1635 3074 1643 3086
rect 1677 3088 1740 3108
rect 1774 3088 1809 3122
rect 1843 3088 1878 3122
rect 1912 3088 1947 3122
rect 1981 3088 2016 3122
rect 2050 3088 2085 3122
rect 2119 3088 2154 3122
rect 2188 3088 2223 3122
rect 2257 3088 2292 3122
rect 2326 3088 2361 3122
rect 2395 3088 2430 3122
rect 2464 3088 2499 3122
rect 2533 3088 2568 3122
rect 2602 3088 2637 3122
rect 2671 3088 2706 3122
rect 2740 3088 2775 3122
rect 2809 3088 2844 3122
rect 4782 3088 4806 3258
rect 1491 3052 1529 3057
rect 1563 3052 1601 3073
rect 1635 3052 1677 3074
rect 1460 3038 1677 3052
rect 1460 3022 1575 3038
rect 1460 3013 1507 3022
rect 1541 3013 1575 3022
rect 1609 3013 1643 3038
rect 1491 2988 1507 3013
rect 1563 3004 1575 3013
rect 1635 3004 1643 3013
rect 1491 2979 1529 2988
rect 1563 2979 1601 3004
rect 1635 2979 1677 3004
rect 1460 2969 1677 2979
rect 1460 2953 1575 2969
rect 1460 2940 1507 2953
rect 1541 2940 1575 2953
rect 1609 2940 1643 2969
rect 1491 2919 1507 2940
rect 1563 2935 1575 2940
rect 1635 2935 1643 2940
rect 1491 2906 1529 2919
rect 1563 2906 1601 2935
rect 1635 2906 1677 2935
rect 1460 2900 1677 2906
rect 1460 2884 1575 2900
rect 1460 2867 1507 2884
rect 1541 2867 1575 2884
rect 1609 2867 1643 2900
rect 1491 2850 1507 2867
rect 1563 2866 1575 2867
rect 1635 2866 1643 2867
rect 1491 2833 1529 2850
rect 1563 2833 1601 2866
rect 1635 2833 1677 2866
rect 1460 2831 1677 2833
rect 1460 2815 1575 2831
rect 1460 2794 1507 2815
rect 1541 2797 1575 2815
rect 1609 2797 1643 2831
rect 1541 2794 1677 2797
rect 1491 2781 1507 2794
rect 1491 2760 1529 2781
rect 1563 2762 1601 2794
rect 1635 2762 1677 2794
rect 1563 2760 1575 2762
rect 1635 2760 1643 2762
rect 1460 2746 1575 2760
rect 1460 2721 1507 2746
rect 1541 2728 1575 2746
rect 1609 2728 1643 2760
rect 1541 2721 1677 2728
rect 1491 2712 1507 2721
rect 1491 2687 1529 2712
rect 1563 2693 1601 2721
rect 1635 2693 1677 2721
rect 1563 2687 1575 2693
rect 1635 2687 1643 2693
rect 1460 2677 1575 2687
rect 1460 2648 1507 2677
rect 1541 2659 1575 2677
rect 1609 2659 1643 2687
rect 1541 2648 1677 2659
rect 1491 2643 1507 2648
rect 1491 2614 1529 2643
rect 1563 2624 1601 2648
rect 1635 2624 1677 2648
rect 1563 2614 1575 2624
rect 1635 2614 1643 2624
rect 1460 2609 1575 2614
rect 1460 2575 1507 2609
rect 1541 2590 1575 2609
rect 1609 2590 1643 2614
rect 1541 2575 1677 2590
rect 1491 2541 1529 2575
rect 1563 2555 1601 2575
rect 1635 2555 1677 2575
rect 1563 2541 1575 2555
rect 1635 2541 1643 2555
rect 1460 2507 1507 2541
rect 1541 2521 1575 2541
rect 1609 2521 1643 2541
rect 1541 2507 1677 2521
rect 1460 2502 1677 2507
rect 1491 2473 1529 2502
rect 1563 2486 1601 2502
rect 1635 2486 1677 2502
rect 1491 2468 1507 2473
rect 1563 2468 1575 2486
rect 1635 2468 1643 2486
rect 1460 2439 1507 2468
rect 1541 2452 1575 2468
rect 1609 2452 1643 2468
rect 1541 2439 1677 2452
rect 1460 2429 1677 2439
rect 1491 2405 1529 2429
rect 1563 2417 1601 2429
rect 1635 2417 1677 2429
rect 1491 2395 1507 2405
rect 1563 2395 1575 2417
rect 1635 2395 1643 2417
rect 1460 2371 1507 2395
rect 1541 2383 1575 2395
rect 1609 2383 1643 2395
rect 1541 2371 1677 2383
rect 1460 2361 1677 2371
rect 4998 2945 8609 3413
rect 4998 2500 5104 2945
rect 8351 2500 8609 2945
rect 4998 2409 8609 2500
rect 4998 2375 7104 2409
rect 7138 2375 7179 2409
rect 7213 2375 7254 2409
rect 7288 2375 7329 2409
rect 7363 2375 7403 2409
rect 7437 2375 7477 2409
rect 7511 2375 7551 2409
rect 7585 2375 7625 2409
rect 7659 2375 7699 2409
rect 7733 2375 7773 2409
rect 7807 2375 7847 2409
rect 7881 2375 7921 2409
rect 7955 2375 7995 2409
rect 8029 2375 8069 2409
rect 8103 2375 8143 2409
rect 8177 2375 8217 2409
rect 8251 2375 8291 2409
rect 8325 2375 8365 2409
rect 8399 2375 8439 2409
rect 8473 2375 8513 2409
rect 8547 2375 8609 2409
rect 1460 2356 1740 2361
rect 1491 2337 1529 2356
rect 1563 2348 1601 2356
rect 1635 2348 1740 2356
rect 1491 2322 1507 2337
rect 1563 2322 1575 2348
rect 1635 2322 1643 2348
rect 1460 2303 1507 2322
rect 1541 2314 1575 2322
rect 1609 2314 1643 2322
rect 1677 2330 1740 2348
rect 1774 2330 1809 2361
rect 1843 2330 1878 2361
rect 1912 2330 1947 2361
rect 1981 2330 2016 2361
rect 2050 2330 2085 2361
rect 1677 2314 1712 2330
rect 1774 2327 1786 2330
rect 1843 2327 1860 2330
rect 1912 2327 1934 2330
rect 1981 2327 2008 2330
rect 2050 2327 2082 2330
rect 2119 2327 2154 2361
rect 2188 2330 2223 2361
rect 2257 2330 2292 2361
rect 2326 2330 2361 2361
rect 2395 2330 2430 2361
rect 2464 2330 2499 2361
rect 2533 2330 2568 2361
rect 2602 2330 2637 2361
rect 2190 2327 2223 2330
rect 2264 2327 2292 2330
rect 2338 2327 2361 2330
rect 2412 2327 2430 2330
rect 2486 2327 2499 2330
rect 2560 2327 2568 2330
rect 2633 2327 2637 2330
rect 2671 2330 2706 2361
rect 2671 2327 2672 2330
rect 1541 2303 1712 2314
rect 1460 2296 1712 2303
rect 1746 2296 1786 2327
rect 1820 2296 1860 2327
rect 1894 2296 1934 2327
rect 1968 2296 2008 2327
rect 2042 2296 2082 2327
rect 2116 2296 2156 2327
rect 2190 2296 2230 2327
rect 2264 2296 2304 2327
rect 2338 2296 2378 2327
rect 2412 2296 2452 2327
rect 2486 2296 2526 2327
rect 2560 2296 2599 2327
rect 2633 2296 2672 2327
rect 2740 2330 2775 2361
rect 2809 2330 2844 2361
rect 2740 2327 2745 2330
rect 2809 2327 2818 2330
rect 2706 2296 2745 2327
rect 2779 2296 2818 2327
rect 1460 2293 2844 2296
rect 1460 2283 1740 2293
rect 1491 2269 1529 2283
rect 1563 2279 1601 2283
rect 1635 2279 1740 2283
rect 1491 2249 1507 2269
rect 1563 2249 1575 2279
rect 1635 2249 1643 2279
rect 1460 2235 1507 2249
rect 1541 2245 1575 2249
rect 1609 2245 1643 2249
rect 1677 2259 1740 2279
rect 1774 2259 1809 2293
rect 1843 2259 1878 2293
rect 1912 2259 1947 2293
rect 1981 2259 2016 2293
rect 2050 2259 2085 2293
rect 2119 2259 2154 2293
rect 2188 2259 2223 2293
rect 2257 2259 2292 2293
rect 2326 2259 2361 2293
rect 2395 2259 2430 2293
rect 2464 2259 2499 2293
rect 2533 2259 2568 2293
rect 2602 2259 2637 2293
rect 2671 2259 2706 2293
rect 2740 2259 2775 2293
rect 2809 2259 2844 2293
rect 1677 2258 2844 2259
rect 1677 2245 1712 2258
rect 1541 2235 1712 2245
rect 1460 2224 1712 2235
rect 1746 2225 1786 2258
rect 1820 2225 1860 2258
rect 1894 2225 1934 2258
rect 1968 2225 2008 2258
rect 2042 2225 2082 2258
rect 2116 2225 2156 2258
rect 2190 2225 2230 2258
rect 2264 2225 2304 2258
rect 2338 2225 2378 2258
rect 2412 2225 2452 2258
rect 2486 2225 2526 2258
rect 2560 2225 2599 2258
rect 2633 2225 2672 2258
rect 1774 2224 1786 2225
rect 1843 2224 1860 2225
rect 1912 2224 1934 2225
rect 1981 2224 2008 2225
rect 2050 2224 2082 2225
rect 1460 2210 1740 2224
rect 1491 2201 1529 2210
rect 1491 2176 1507 2201
rect 1563 2176 1575 2210
rect 1635 2176 1643 2210
rect 1677 2191 1740 2210
rect 1774 2191 1809 2224
rect 1843 2191 1878 2224
rect 1912 2191 1947 2224
rect 1981 2191 2016 2224
rect 2050 2191 2085 2224
rect 2119 2191 2154 2225
rect 2190 2224 2223 2225
rect 2264 2224 2292 2225
rect 2338 2224 2361 2225
rect 2412 2224 2430 2225
rect 2486 2224 2499 2225
rect 2560 2224 2568 2225
rect 2633 2224 2637 2225
rect 2188 2191 2223 2224
rect 2257 2191 2292 2224
rect 2326 2191 2361 2224
rect 2395 2191 2430 2224
rect 2464 2191 2499 2224
rect 2533 2191 2568 2224
rect 2602 2191 2637 2224
rect 2671 2224 2672 2225
rect 2706 2225 2745 2258
rect 2779 2225 2818 2258
rect 2671 2191 2706 2224
rect 2740 2224 2745 2225
rect 2809 2224 2818 2225
rect 2740 2191 2775 2224
rect 2809 2191 2844 2224
rect 4782 2191 4806 2361
rect 4998 2337 8609 2375
rect 4998 2303 7104 2337
rect 7138 2303 7179 2337
rect 7213 2303 7254 2337
rect 7288 2303 7329 2337
rect 7363 2303 7403 2337
rect 7437 2303 7477 2337
rect 7511 2303 7551 2337
rect 7585 2303 7625 2337
rect 7659 2303 7699 2337
rect 7733 2303 7773 2337
rect 7807 2303 7847 2337
rect 7881 2303 7921 2337
rect 7955 2303 7995 2337
rect 8029 2303 8069 2337
rect 8103 2303 8143 2337
rect 8177 2303 8217 2337
rect 8251 2303 8291 2337
rect 8325 2303 8365 2337
rect 8399 2303 8439 2337
rect 8473 2303 8513 2337
rect 8547 2303 8609 2337
rect 4998 2265 8609 2303
rect 4998 2231 7104 2265
rect 7138 2231 7179 2265
rect 7213 2231 7254 2265
rect 7288 2231 7329 2265
rect 7363 2231 7403 2265
rect 7437 2231 7477 2265
rect 7511 2231 7551 2265
rect 7585 2231 7625 2265
rect 7659 2231 7699 2265
rect 7733 2231 7773 2265
rect 7807 2231 7847 2265
rect 7881 2231 7921 2265
rect 7955 2231 7995 2265
rect 8029 2231 8069 2265
rect 8103 2231 8143 2265
rect 8177 2231 8217 2265
rect 8251 2231 8291 2265
rect 8325 2231 8365 2265
rect 8399 2231 8439 2265
rect 8473 2231 8513 2265
rect 8547 2231 8609 2265
rect 1460 2167 1507 2176
rect 1541 2167 1677 2176
rect 1460 2141 1677 2167
rect 1460 2137 1575 2141
rect 1609 2137 1643 2141
rect 1491 2133 1529 2137
rect 1491 2103 1507 2133
rect 1563 2107 1575 2137
rect 1635 2107 1643 2137
rect 1563 2103 1601 2107
rect 1635 2103 1677 2107
rect 1460 2099 1507 2103
rect 1541 2099 1677 2103
rect 1460 2072 1677 2099
rect 1460 2065 1575 2072
rect 1460 2064 1507 2065
rect 1541 2064 1575 2065
rect 1609 2064 1643 2072
rect 1491 2031 1507 2064
rect 1563 2038 1575 2064
rect 1635 2038 1643 2064
rect 1491 2030 1529 2031
rect 1563 2030 1601 2038
rect 1635 2030 1677 2038
rect 1460 2003 1677 2030
rect 1460 1997 1575 2003
rect 1460 1991 1507 1997
rect 1541 1991 1575 1997
rect 1609 1991 1643 2003
rect 1491 1963 1507 1991
rect 1563 1969 1575 1991
rect 1635 1969 1643 1991
rect 1491 1957 1529 1963
rect 1563 1957 1601 1969
rect 1635 1957 1677 1969
rect 1460 1934 1677 1957
rect 1460 1929 1575 1934
rect 1460 1918 1507 1929
rect 1541 1918 1575 1929
rect 1609 1918 1643 1934
rect 1491 1895 1507 1918
rect 1563 1900 1575 1918
rect 1635 1900 1643 1918
rect 1491 1884 1529 1895
rect 1563 1884 1601 1900
rect 1635 1884 1677 1900
rect 1460 1865 1677 1884
rect 1460 1861 1575 1865
rect 1460 1845 1507 1861
rect 1541 1845 1575 1861
rect 1609 1845 1643 1865
rect 1491 1827 1507 1845
rect 1563 1831 1575 1845
rect 1635 1831 1643 1845
rect 1491 1811 1529 1827
rect 1563 1811 1601 1831
rect 1635 1811 1677 1831
rect 1460 1796 1677 1811
rect 4998 2032 8609 2231
rect 8677 3636 8711 3670
rect 8745 3636 8779 3670
rect 8813 3663 8847 3670
rect 8881 3663 8915 3670
rect 8949 3663 8983 3670
rect 9017 3663 9051 3670
rect 8813 3636 8824 3663
rect 8881 3636 8898 3663
rect 8949 3636 8972 3663
rect 9017 3636 9046 3663
rect 9085 3636 9119 3670
rect 9153 3663 9187 3670
rect 9221 3663 9255 3670
rect 9289 3663 9323 3670
rect 9357 3663 9391 3670
rect 9425 3663 9459 3670
rect 9493 3663 9527 3670
rect 9154 3636 9187 3663
rect 9228 3636 9255 3663
rect 9302 3636 9323 3663
rect 9376 3636 9391 3663
rect 9450 3636 9459 3663
rect 9524 3636 9527 3663
rect 9561 3663 9595 3670
rect 9629 3663 9663 3670
rect 9697 3663 9731 3670
rect 9765 3663 9799 3670
rect 9833 3663 9867 3670
rect 9901 3663 9935 3670
rect 9561 3636 9564 3663
rect 9629 3636 9638 3663
rect 9697 3636 9712 3663
rect 9765 3636 9786 3663
rect 9833 3636 9860 3663
rect 9901 3636 9934 3663
rect 9969 3636 10003 3670
rect 10037 3663 10071 3670
rect 10105 3663 10139 3670
rect 10173 3663 10207 3670
rect 10241 3663 10312 3670
rect 10346 3663 10380 3671
rect 10042 3636 10071 3663
rect 10116 3636 10139 3663
rect 10190 3636 10207 3663
rect 8643 3629 8824 3636
rect 8858 3629 8898 3636
rect 8932 3629 8972 3636
rect 9006 3629 9046 3636
rect 9080 3629 9120 3636
rect 9154 3629 9194 3636
rect 9228 3629 9268 3636
rect 9302 3629 9342 3636
rect 9376 3629 9416 3636
rect 9450 3629 9490 3636
rect 9524 3629 9564 3636
rect 9598 3629 9638 3636
rect 9672 3629 9712 3636
rect 9746 3629 9786 3636
rect 9820 3629 9860 3636
rect 9894 3629 9934 3636
rect 9968 3629 10008 3636
rect 10042 3629 10082 3636
rect 10116 3629 10156 3636
rect 10190 3629 10230 3636
rect 10264 3629 10304 3663
rect 10346 3637 10378 3663
rect 10414 3637 10448 3671
rect 10482 3663 10516 3671
rect 10550 3663 10584 3671
rect 10618 3663 10652 3671
rect 10686 3663 10720 3671
rect 10754 3663 10788 3671
rect 10486 3637 10516 3663
rect 10560 3637 10584 3663
rect 10634 3637 10652 3663
rect 10708 3637 10720 3663
rect 10782 3637 10788 3663
rect 10822 3663 10856 3671
rect 10338 3629 10378 3637
rect 10412 3629 10452 3637
rect 10486 3629 10526 3637
rect 10560 3629 10600 3637
rect 10634 3629 10674 3637
rect 10708 3629 10748 3637
rect 10782 3629 10822 3637
rect 10890 3663 10924 3671
rect 10958 3663 10992 3671
rect 11026 3663 11060 3671
rect 11094 3663 11128 3671
rect 11162 3663 11196 3671
rect 11230 3663 11264 3671
rect 10890 3637 10896 3663
rect 10958 3637 10970 3663
rect 11026 3637 11043 3663
rect 11094 3637 11116 3663
rect 11162 3637 11189 3663
rect 11230 3637 11262 3663
rect 11298 3637 11332 3671
rect 11366 3663 11400 3671
rect 11434 3663 11468 3671
rect 11502 3663 11536 3671
rect 11369 3637 11400 3663
rect 11442 3637 11468 3663
rect 11515 3637 11536 3663
rect 11570 3637 11589 3671
rect 10856 3629 10896 3637
rect 10930 3629 10970 3637
rect 11004 3629 11043 3637
rect 11077 3629 11116 3637
rect 11150 3629 11189 3637
rect 11223 3629 11262 3637
rect 11296 3629 11335 3637
rect 11369 3629 11408 3637
rect 11442 3629 11481 3637
rect 11515 3629 11589 3637
rect 8643 3601 11589 3629
rect 8643 3600 10312 3601
rect 8677 3566 8711 3600
rect 8745 3566 8779 3600
rect 8813 3591 8847 3600
rect 8881 3591 8915 3600
rect 8949 3591 8983 3600
rect 9017 3591 9051 3600
rect 8813 3566 8824 3591
rect 8881 3566 8898 3591
rect 8949 3566 8972 3591
rect 9017 3566 9046 3591
rect 9085 3566 9119 3600
rect 9153 3591 9187 3600
rect 9221 3591 9255 3600
rect 9289 3591 9323 3600
rect 9357 3591 9391 3600
rect 9425 3591 9459 3600
rect 9493 3591 9527 3600
rect 9154 3566 9187 3591
rect 9228 3566 9255 3591
rect 9302 3566 9323 3591
rect 9376 3566 9391 3591
rect 9450 3566 9459 3591
rect 9524 3566 9527 3591
rect 9561 3591 9595 3600
rect 9629 3591 9663 3600
rect 9697 3591 9731 3600
rect 9765 3591 9799 3600
rect 9833 3591 9867 3600
rect 9901 3591 9935 3600
rect 9561 3566 9564 3591
rect 9629 3566 9638 3591
rect 9697 3566 9712 3591
rect 9765 3566 9786 3591
rect 9833 3566 9860 3591
rect 9901 3566 9934 3591
rect 9969 3566 10003 3600
rect 10037 3591 10071 3600
rect 10105 3591 10139 3600
rect 10173 3591 10207 3600
rect 10241 3591 10312 3600
rect 10346 3591 10380 3601
rect 10042 3566 10071 3591
rect 10116 3566 10139 3591
rect 10190 3566 10207 3591
rect 8643 3557 8824 3566
rect 8858 3557 8898 3566
rect 8932 3557 8972 3566
rect 9006 3557 9046 3566
rect 9080 3557 9120 3566
rect 9154 3557 9194 3566
rect 9228 3557 9268 3566
rect 9302 3557 9342 3566
rect 9376 3557 9416 3566
rect 9450 3557 9490 3566
rect 9524 3557 9564 3566
rect 9598 3557 9638 3566
rect 9672 3557 9712 3566
rect 9746 3557 9786 3566
rect 9820 3557 9860 3566
rect 9894 3557 9934 3566
rect 9968 3557 10008 3566
rect 10042 3557 10082 3566
rect 10116 3557 10156 3566
rect 10190 3557 10230 3566
rect 10264 3557 10304 3591
rect 10346 3567 10378 3591
rect 10414 3567 10448 3601
rect 10482 3591 10516 3601
rect 10550 3591 10584 3601
rect 10618 3591 10652 3601
rect 10686 3591 10720 3601
rect 10754 3591 10788 3601
rect 10486 3567 10516 3591
rect 10560 3567 10584 3591
rect 10634 3567 10652 3591
rect 10708 3567 10720 3591
rect 10782 3567 10788 3591
rect 10822 3591 10856 3601
rect 10338 3557 10378 3567
rect 10412 3557 10452 3567
rect 10486 3557 10526 3567
rect 10560 3557 10600 3567
rect 10634 3557 10674 3567
rect 10708 3557 10748 3567
rect 10782 3557 10822 3567
rect 10890 3591 10924 3601
rect 10958 3591 10992 3601
rect 11026 3591 11060 3601
rect 11094 3591 11128 3601
rect 11162 3591 11196 3601
rect 11230 3591 11264 3601
rect 10890 3567 10896 3591
rect 10958 3567 10970 3591
rect 11026 3567 11043 3591
rect 11094 3567 11116 3591
rect 11162 3567 11189 3591
rect 11230 3567 11262 3591
rect 11298 3567 11332 3601
rect 11366 3591 11400 3601
rect 11434 3591 11468 3601
rect 11502 3591 11536 3601
rect 11369 3567 11400 3591
rect 11442 3567 11468 3591
rect 11515 3567 11536 3591
rect 11570 3567 11589 3601
rect 10856 3557 10896 3567
rect 10930 3557 10970 3567
rect 11004 3557 11043 3567
rect 11077 3557 11116 3567
rect 11150 3557 11189 3567
rect 11223 3557 11262 3567
rect 11296 3557 11335 3567
rect 11369 3557 11408 3567
rect 11442 3557 11481 3567
rect 11515 3557 11589 3567
rect 8643 3531 11589 3557
rect 8643 3530 10312 3531
rect 8677 3496 8711 3530
rect 8745 3496 8779 3530
rect 8813 3519 8847 3530
rect 8881 3519 8915 3530
rect 8949 3519 8983 3530
rect 9017 3519 9051 3530
rect 8813 3496 8824 3519
rect 8881 3496 8898 3519
rect 8949 3496 8972 3519
rect 9017 3496 9046 3519
rect 9085 3496 9119 3530
rect 9153 3519 9187 3530
rect 9221 3519 9255 3530
rect 9289 3519 9323 3530
rect 9357 3519 9391 3530
rect 9425 3519 9459 3530
rect 9493 3519 9527 3530
rect 9154 3496 9187 3519
rect 9228 3496 9255 3519
rect 9302 3496 9323 3519
rect 9376 3496 9391 3519
rect 9450 3496 9459 3519
rect 9524 3496 9527 3519
rect 9561 3519 9595 3530
rect 9629 3519 9663 3530
rect 9697 3519 9731 3530
rect 9765 3519 9799 3530
rect 9833 3519 9867 3530
rect 9901 3519 9935 3530
rect 9561 3496 9564 3519
rect 9629 3496 9638 3519
rect 9697 3496 9712 3519
rect 9765 3496 9786 3519
rect 9833 3496 9860 3519
rect 9901 3496 9934 3519
rect 9969 3496 10003 3530
rect 10037 3519 10071 3530
rect 10105 3519 10139 3530
rect 10173 3519 10207 3530
rect 10241 3519 10312 3530
rect 10346 3519 10380 3531
rect 10042 3496 10071 3519
rect 10116 3496 10139 3519
rect 10190 3496 10207 3519
rect 8643 3485 8824 3496
rect 8858 3485 8898 3496
rect 8932 3485 8972 3496
rect 9006 3485 9046 3496
rect 9080 3485 9120 3496
rect 9154 3485 9194 3496
rect 9228 3485 9268 3496
rect 9302 3485 9342 3496
rect 9376 3485 9416 3496
rect 9450 3485 9490 3496
rect 9524 3485 9564 3496
rect 9598 3485 9638 3496
rect 9672 3485 9712 3496
rect 9746 3485 9786 3496
rect 9820 3485 9860 3496
rect 9894 3485 9934 3496
rect 9968 3485 10008 3496
rect 10042 3485 10082 3496
rect 10116 3485 10156 3496
rect 10190 3485 10230 3496
rect 10264 3485 10304 3519
rect 10346 3497 10378 3519
rect 10414 3497 10448 3531
rect 10482 3519 10516 3531
rect 10550 3519 10584 3531
rect 10618 3519 10652 3531
rect 10686 3519 10720 3531
rect 10754 3519 10788 3531
rect 10486 3497 10516 3519
rect 10560 3497 10584 3519
rect 10634 3497 10652 3519
rect 10708 3497 10720 3519
rect 10782 3497 10788 3519
rect 10822 3519 10856 3531
rect 10338 3485 10378 3497
rect 10412 3485 10452 3497
rect 10486 3485 10526 3497
rect 10560 3485 10600 3497
rect 10634 3485 10674 3497
rect 10708 3485 10748 3497
rect 10782 3485 10822 3497
rect 10890 3519 10924 3531
rect 10958 3519 10992 3531
rect 11026 3519 11060 3531
rect 11094 3519 11128 3531
rect 11162 3519 11196 3531
rect 11230 3519 11264 3531
rect 10890 3497 10896 3519
rect 10958 3497 10970 3519
rect 11026 3497 11043 3519
rect 11094 3497 11116 3519
rect 11162 3497 11189 3519
rect 11230 3497 11262 3519
rect 11298 3497 11332 3531
rect 11366 3519 11400 3531
rect 11434 3519 11468 3531
rect 11502 3519 11536 3531
rect 11369 3497 11400 3519
rect 11442 3497 11468 3519
rect 11515 3497 11536 3519
rect 11570 3497 11589 3531
rect 10856 3485 10896 3497
rect 10930 3485 10970 3497
rect 11004 3485 11043 3497
rect 11077 3485 11116 3497
rect 11150 3485 11189 3497
rect 11223 3485 11262 3497
rect 11296 3485 11335 3497
rect 11369 3485 11408 3497
rect 11442 3485 11481 3497
rect 11515 3485 11589 3497
rect 8643 3475 11589 3485
rect 12582 4363 13390 4387
rect 12582 4329 12595 4363
rect 12629 4329 12663 4363
rect 12697 4329 12731 4363
rect 12765 4329 12799 4363
rect 12833 4329 12867 4363
rect 12901 4329 12935 4363
rect 12969 4329 13003 4363
rect 13037 4329 13071 4363
rect 13105 4329 13139 4363
rect 13173 4329 13207 4363
rect 13241 4329 13275 4363
rect 13309 4329 13343 4363
rect 13377 4329 13390 4363
rect 12582 4293 13390 4329
rect 12582 4259 12595 4293
rect 12629 4259 12663 4293
rect 12697 4259 12731 4293
rect 12765 4259 12799 4293
rect 12833 4259 12867 4293
rect 12901 4259 12935 4293
rect 12969 4259 13003 4293
rect 13037 4259 13071 4293
rect 13105 4259 13139 4293
rect 13173 4259 13207 4293
rect 13241 4259 13275 4293
rect 13309 4259 13343 4293
rect 13377 4259 13390 4293
rect 23568 4364 23593 4398
rect 23627 4392 23665 4398
rect 23699 4392 23737 4398
rect 23568 4358 23597 4364
rect 23631 4358 23665 4392
rect 23699 4358 23733 4392
rect 23771 4364 23796 4398
rect 23767 4358 23796 4364
rect 23568 4325 23796 4358
rect 23568 4291 23593 4325
rect 23627 4323 23665 4325
rect 23699 4323 23737 4325
rect 23568 4289 23597 4291
rect 23631 4289 23665 4323
rect 23699 4289 23733 4323
rect 23771 4291 23796 4325
rect 23767 4289 23796 4291
rect 12582 4223 13390 4259
rect 16974 4257 17080 4279
rect 16974 4256 16976 4257
rect 12582 4189 12595 4223
rect 12629 4189 12663 4223
rect 12697 4189 12731 4223
rect 12765 4189 12799 4223
rect 12833 4189 12867 4223
rect 12901 4189 12935 4223
rect 12969 4189 13003 4223
rect 13037 4189 13071 4223
rect 13105 4189 13139 4223
rect 13173 4189 13207 4223
rect 13241 4189 13275 4223
rect 13309 4189 13343 4223
rect 13377 4189 13390 4223
rect 17010 4223 17044 4257
rect 17078 4256 17080 4257
rect 17007 4222 17045 4223
rect 17079 4222 17080 4256
rect 16974 4207 17080 4222
rect 19118 4257 19220 4273
rect 19158 4223 19186 4257
rect 23568 4254 23796 4289
rect 23568 4252 23597 4254
rect 19118 4207 19220 4223
rect 23568 4218 23593 4252
rect 23631 4220 23665 4254
rect 23699 4220 23733 4254
rect 23767 4252 23796 4254
rect 23627 4218 23665 4220
rect 23699 4218 23737 4220
rect 23771 4218 23796 4252
rect 12582 4153 13390 4189
rect 12582 4119 12595 4153
rect 12629 4119 12663 4153
rect 12697 4119 12731 4153
rect 12765 4119 12799 4153
rect 12833 4119 12867 4153
rect 12901 4119 12935 4153
rect 12969 4119 13003 4153
rect 13037 4119 13071 4153
rect 13105 4119 13139 4153
rect 13173 4119 13207 4153
rect 13241 4119 13275 4153
rect 13309 4119 13343 4153
rect 13377 4119 13390 4153
rect 12582 4083 13390 4119
rect 12582 4059 12595 4083
rect 12629 4059 12663 4083
rect 12697 4059 12731 4083
rect 12765 4059 12799 4083
rect 12833 4059 12867 4083
rect 12901 4059 12935 4083
rect 12969 4059 13003 4083
rect 13037 4059 13071 4083
rect 13105 4059 13139 4083
rect 13173 4059 13207 4083
rect 13241 4059 13275 4083
rect 13309 4059 13343 4083
rect 13377 4059 13390 4083
rect 23568 4185 23796 4218
rect 23568 4179 23597 4185
rect 23568 4145 23593 4179
rect 23631 4151 23665 4185
rect 23699 4151 23733 4185
rect 23767 4179 23796 4185
rect 23627 4145 23665 4151
rect 23699 4145 23737 4151
rect 23771 4145 23796 4179
rect 23568 4116 23796 4145
rect 23568 4106 23597 4116
rect 23767 4106 23796 4116
rect 23568 4072 23593 4106
rect 23771 4072 23796 4106
rect 12582 3881 12594 4059
rect 23568 4033 23597 4072
rect 23767 4033 23796 4072
rect 23568 3999 23593 4033
rect 23771 3999 23796 4033
rect 23568 3960 23597 3999
rect 23767 3960 23796 3999
rect 23568 3926 23593 3960
rect 23771 3926 23796 3960
rect 23568 3887 23597 3926
rect 23767 3887 23796 3926
rect 12582 3873 13390 3881
rect 12582 3839 12595 3873
rect 12629 3839 12663 3873
rect 12697 3839 12731 3873
rect 12765 3839 12799 3873
rect 12833 3839 12867 3873
rect 12901 3839 12935 3873
rect 12969 3839 13003 3873
rect 13037 3839 13071 3873
rect 13105 3839 13139 3873
rect 13173 3839 13207 3873
rect 13241 3839 13275 3873
rect 13309 3839 13343 3873
rect 13377 3839 13390 3873
rect 12582 3803 13390 3839
rect 12582 3769 12595 3803
rect 12629 3769 12663 3803
rect 12697 3769 12731 3803
rect 12765 3769 12799 3803
rect 12833 3769 12867 3803
rect 12901 3769 12935 3803
rect 12969 3769 13003 3803
rect 13037 3769 13071 3803
rect 13105 3769 13139 3803
rect 13173 3769 13207 3803
rect 13241 3769 13275 3803
rect 13309 3769 13343 3803
rect 13377 3769 13390 3803
rect 12582 3765 13390 3769
rect 23568 3853 23593 3887
rect 23771 3853 23796 3887
rect 23568 3814 23597 3853
rect 23767 3814 23796 3853
rect 23568 3780 23593 3814
rect 23771 3780 23796 3814
rect 12582 3731 12594 3765
rect 12628 3733 12667 3765
rect 12701 3733 12740 3765
rect 12774 3733 12813 3765
rect 12847 3733 12886 3765
rect 12920 3733 12959 3765
rect 12993 3733 13032 3765
rect 13066 3733 13105 3765
rect 12582 3699 12595 3731
rect 12629 3699 12663 3733
rect 12701 3731 12731 3733
rect 12774 3731 12799 3733
rect 12847 3731 12867 3733
rect 12920 3731 12935 3733
rect 12993 3731 13003 3733
rect 13066 3731 13071 3733
rect 12697 3699 12731 3731
rect 12765 3699 12799 3731
rect 12833 3699 12867 3731
rect 12901 3699 12935 3731
rect 12969 3699 13003 3731
rect 13037 3699 13071 3731
rect 13139 3733 13178 3765
rect 13212 3733 13251 3765
rect 13285 3733 13324 3765
rect 13358 3733 13397 3765
rect 13105 3699 13139 3731
rect 13173 3731 13178 3733
rect 13241 3731 13251 3733
rect 13309 3731 13324 3733
rect 13377 3731 13397 3733
rect 13431 3731 13470 3765
rect 13504 3731 13543 3765
rect 13577 3731 13616 3765
rect 13650 3731 13689 3765
rect 13723 3731 13762 3765
rect 13796 3731 13835 3765
rect 13869 3731 13908 3765
rect 13942 3731 13981 3765
rect 14015 3731 14054 3765
rect 14088 3731 14127 3765
rect 14161 3731 14200 3765
rect 14234 3731 14273 3765
rect 14307 3731 14346 3765
rect 14380 3731 14419 3765
rect 14453 3731 14492 3765
rect 14526 3731 14565 3765
rect 14599 3731 14638 3765
rect 14672 3731 14711 3765
rect 14745 3731 14784 3765
rect 14818 3731 14857 3765
rect 14891 3731 14930 3765
rect 14964 3731 15003 3765
rect 15037 3731 15076 3765
rect 15110 3731 15149 3765
rect 15183 3731 15222 3765
rect 15256 3731 15295 3765
rect 15329 3731 15368 3765
rect 15402 3731 15441 3765
rect 15475 3731 15514 3765
rect 15548 3731 15587 3765
rect 15621 3731 15660 3765
rect 15694 3731 15733 3765
rect 15767 3731 15806 3765
rect 15840 3731 15879 3765
rect 15913 3731 15952 3765
rect 15986 3731 16025 3765
rect 16059 3731 16098 3765
rect 16132 3731 16171 3765
rect 16205 3731 16244 3765
rect 16278 3731 16317 3765
rect 16351 3731 16390 3765
rect 13173 3699 13207 3731
rect 13241 3699 13275 3731
rect 13309 3699 13343 3731
rect 13377 3699 16424 3731
rect 12582 3693 16424 3699
rect 12582 3659 12594 3693
rect 12628 3663 12667 3693
rect 12701 3663 12740 3693
rect 12774 3663 12813 3693
rect 12847 3663 12886 3693
rect 12920 3663 12959 3693
rect 12993 3663 13032 3693
rect 13066 3663 13105 3693
rect 12582 3629 12595 3659
rect 12629 3629 12663 3663
rect 12701 3659 12731 3663
rect 12774 3659 12799 3663
rect 12847 3659 12867 3663
rect 12920 3659 12935 3663
rect 12993 3659 13003 3663
rect 13066 3659 13071 3663
rect 12697 3629 12731 3659
rect 12765 3629 12799 3659
rect 12833 3629 12867 3659
rect 12901 3629 12935 3659
rect 12969 3629 13003 3659
rect 13037 3629 13071 3659
rect 13139 3663 13178 3693
rect 13212 3663 13251 3693
rect 13285 3663 13324 3693
rect 13358 3663 13397 3693
rect 13105 3629 13139 3659
rect 13173 3659 13178 3663
rect 13241 3659 13251 3663
rect 13309 3659 13324 3663
rect 13377 3659 13397 3663
rect 13431 3659 13470 3693
rect 13504 3659 13543 3693
rect 13577 3659 13616 3693
rect 13650 3659 13689 3693
rect 13723 3659 13762 3693
rect 13796 3659 13835 3693
rect 13869 3659 13908 3693
rect 13942 3659 13981 3693
rect 14015 3659 14054 3693
rect 14088 3659 14127 3693
rect 14161 3659 14200 3693
rect 14234 3659 14273 3693
rect 14307 3659 14346 3693
rect 14380 3659 14419 3693
rect 14453 3659 14492 3693
rect 14526 3659 14565 3693
rect 14599 3659 14638 3693
rect 14672 3659 14711 3693
rect 14745 3659 14784 3693
rect 14818 3659 14857 3693
rect 14891 3659 14930 3693
rect 14964 3659 15003 3693
rect 15037 3659 15076 3693
rect 15110 3659 15149 3693
rect 15183 3659 15222 3693
rect 15256 3659 15295 3693
rect 15329 3659 15368 3693
rect 15402 3659 15441 3693
rect 15475 3659 15514 3693
rect 15548 3659 15587 3693
rect 15621 3659 15660 3693
rect 15694 3659 15733 3693
rect 15767 3659 15806 3693
rect 15840 3659 15879 3693
rect 15913 3659 15952 3693
rect 15986 3659 16025 3693
rect 16059 3659 16098 3693
rect 16132 3659 16171 3693
rect 16205 3659 16244 3693
rect 16278 3659 16317 3693
rect 16351 3659 16390 3693
rect 13173 3629 13207 3659
rect 13241 3629 13275 3659
rect 13309 3629 13343 3659
rect 13377 3629 16424 3659
rect 12582 3621 16424 3629
rect 12582 3587 12594 3621
rect 12628 3593 12667 3621
rect 12701 3593 12740 3621
rect 12774 3593 12813 3621
rect 12847 3593 12886 3621
rect 12920 3593 12959 3621
rect 12993 3593 13032 3621
rect 13066 3593 13105 3621
rect 12582 3559 12595 3587
rect 12629 3559 12663 3593
rect 12701 3587 12731 3593
rect 12774 3587 12799 3593
rect 12847 3587 12867 3593
rect 12920 3587 12935 3593
rect 12993 3587 13003 3593
rect 13066 3587 13071 3593
rect 12697 3559 12731 3587
rect 12765 3559 12799 3587
rect 12833 3559 12867 3587
rect 12901 3559 12935 3587
rect 12969 3559 13003 3587
rect 13037 3559 13071 3587
rect 13139 3593 13178 3621
rect 13212 3593 13251 3621
rect 13285 3593 13324 3621
rect 13358 3593 13397 3621
rect 13105 3559 13139 3587
rect 13173 3587 13178 3593
rect 13241 3587 13251 3593
rect 13309 3587 13324 3593
rect 13377 3587 13397 3593
rect 13431 3587 13470 3621
rect 13504 3587 13543 3621
rect 13577 3587 13616 3621
rect 13650 3587 13689 3621
rect 13723 3587 13762 3621
rect 13796 3587 13835 3621
rect 13869 3587 13908 3621
rect 13942 3587 13981 3621
rect 14015 3587 14054 3621
rect 14088 3587 14127 3621
rect 14161 3587 14200 3621
rect 14234 3587 14273 3621
rect 14307 3587 14346 3621
rect 14380 3587 14419 3621
rect 14453 3587 14492 3621
rect 14526 3587 14565 3621
rect 14599 3587 14638 3621
rect 14672 3587 14711 3621
rect 14745 3587 14784 3621
rect 14818 3587 14857 3621
rect 14891 3587 14930 3621
rect 14964 3587 15003 3621
rect 15037 3587 15076 3621
rect 15110 3587 15149 3621
rect 15183 3587 15222 3621
rect 15256 3587 15295 3621
rect 15329 3587 15368 3621
rect 15402 3587 15441 3621
rect 15475 3587 15514 3621
rect 15548 3587 15587 3621
rect 15621 3587 15660 3621
rect 15694 3587 15733 3621
rect 15767 3587 15806 3621
rect 15840 3587 15879 3621
rect 15913 3587 15952 3621
rect 15986 3587 16025 3621
rect 16059 3587 16098 3621
rect 16132 3587 16171 3621
rect 16205 3587 16244 3621
rect 16278 3587 16317 3621
rect 16351 3587 16390 3621
rect 23568 3741 23597 3780
rect 23767 3741 23796 3780
rect 23568 3707 23593 3741
rect 23771 3707 23796 3741
rect 23568 3668 23597 3707
rect 23767 3668 23796 3707
rect 23568 3634 23593 3668
rect 23771 3634 23796 3668
rect 23568 3595 23597 3634
rect 23767 3595 23796 3634
rect 13173 3559 13207 3587
rect 13241 3559 13275 3587
rect 13309 3559 13343 3587
rect 13377 3559 13390 3587
rect 12582 3523 13390 3559
rect 12582 3489 12595 3523
rect 12629 3489 12663 3523
rect 12697 3489 12731 3523
rect 12765 3489 12799 3523
rect 12833 3489 12867 3523
rect 12901 3489 12935 3523
rect 12969 3489 13003 3523
rect 13037 3489 13071 3523
rect 13105 3489 13139 3523
rect 13173 3489 13207 3523
rect 13241 3489 13275 3523
rect 13309 3489 13343 3523
rect 13377 3489 13390 3523
rect 12582 3475 13390 3489
rect 23568 3561 23593 3595
rect 23771 3561 23796 3595
rect 23568 3522 23597 3561
rect 23767 3522 23796 3561
rect 23568 3488 23593 3522
rect 23771 3488 23796 3522
rect 8643 3461 11590 3475
rect 8643 3460 10312 3461
rect 8677 3426 8711 3460
rect 8745 3426 8779 3460
rect 8813 3447 8847 3460
rect 8881 3447 8915 3460
rect 8949 3447 8983 3460
rect 9017 3447 9051 3460
rect 9085 3447 9119 3460
rect 8813 3426 8824 3447
rect 8881 3426 8897 3447
rect 8949 3426 8970 3447
rect 9017 3426 9043 3447
rect 9085 3426 9116 3447
rect 9153 3426 9187 3460
rect 9221 3447 9255 3460
rect 9289 3447 9323 3460
rect 9357 3447 9391 3460
rect 9425 3447 9459 3460
rect 9493 3447 9527 3460
rect 9561 3447 9595 3460
rect 9223 3426 9255 3447
rect 9296 3426 9323 3447
rect 9370 3426 9391 3447
rect 9444 3426 9459 3447
rect 9518 3426 9527 3447
rect 9592 3426 9595 3447
rect 9629 3447 9663 3460
rect 9697 3447 9731 3460
rect 9765 3447 9799 3460
rect 9833 3447 9867 3460
rect 9901 3447 9935 3460
rect 9969 3447 10003 3460
rect 9629 3426 9632 3447
rect 9697 3426 9706 3447
rect 9765 3426 9780 3447
rect 9833 3426 9854 3447
rect 9901 3426 9928 3447
rect 9969 3426 10002 3447
rect 10037 3426 10071 3460
rect 10105 3447 10139 3460
rect 10173 3447 10207 3460
rect 10241 3447 10312 3460
rect 10346 3447 10380 3461
rect 10414 3447 10448 3461
rect 10110 3426 10139 3447
rect 10184 3426 10207 3447
rect 8643 3413 8824 3426
rect 8858 3413 8897 3426
rect 8931 3413 8970 3426
rect 9004 3413 9043 3426
rect 9077 3413 9116 3426
rect 9150 3413 9189 3426
rect 9223 3413 9262 3426
rect 9296 3413 9336 3426
rect 9370 3413 9410 3426
rect 9444 3413 9484 3426
rect 9518 3413 9558 3426
rect 9592 3413 9632 3426
rect 9666 3413 9706 3426
rect 9740 3413 9780 3426
rect 9814 3413 9854 3426
rect 9888 3413 9928 3426
rect 9962 3413 10002 3426
rect 10036 3413 10076 3426
rect 10110 3413 10150 3426
rect 10184 3413 10224 3426
rect 10258 3413 10298 3447
rect 10346 3427 10372 3447
rect 10414 3427 10446 3447
rect 10482 3427 10516 3461
rect 10550 3447 10584 3461
rect 10618 3447 10652 3461
rect 10686 3447 10720 3461
rect 10754 3447 10788 3461
rect 10822 3447 10856 3461
rect 10554 3427 10584 3447
rect 10628 3427 10652 3447
rect 10702 3427 10720 3447
rect 10776 3427 10788 3447
rect 10850 3427 10856 3447
rect 10890 3447 10924 3461
rect 10332 3413 10372 3427
rect 10406 3413 10446 3427
rect 10480 3413 10520 3427
rect 10554 3413 10594 3427
rect 10628 3413 10668 3427
rect 10702 3413 10742 3427
rect 10776 3413 10816 3427
rect 10850 3413 10890 3427
rect 10958 3447 10992 3461
rect 11026 3447 11060 3461
rect 11094 3447 11128 3461
rect 11162 3447 11196 3461
rect 11230 3447 11264 3461
rect 10958 3427 10964 3447
rect 11026 3427 11038 3447
rect 11094 3427 11112 3447
rect 11162 3427 11186 3447
rect 11230 3427 11260 3447
rect 11298 3427 11332 3461
rect 11366 3447 11400 3461
rect 11434 3447 11468 3461
rect 11502 3447 11536 3461
rect 11570 3447 11590 3461
rect 11368 3427 11400 3447
rect 11442 3427 11468 3447
rect 11516 3427 11536 3447
rect 10924 3413 10964 3427
rect 10998 3413 11038 3427
rect 11072 3413 11112 3427
rect 11146 3413 11186 3427
rect 11220 3413 11260 3427
rect 11294 3413 11334 3427
rect 11368 3413 11408 3427
rect 11442 3413 11482 3427
rect 11516 3413 11556 3427
rect 8643 3391 11590 3413
rect 8643 3390 10312 3391
rect 8677 3356 8711 3390
rect 8745 3356 8779 3390
rect 8813 3375 8847 3390
rect 8881 3375 8915 3390
rect 8949 3375 8983 3390
rect 9017 3375 9051 3390
rect 9085 3375 9119 3390
rect 8813 3356 8824 3375
rect 8881 3356 8897 3375
rect 8949 3356 8970 3375
rect 9017 3356 9043 3375
rect 9085 3356 9116 3375
rect 9153 3356 9187 3390
rect 9221 3375 9255 3390
rect 9289 3375 9323 3390
rect 9357 3375 9391 3390
rect 9425 3375 9459 3390
rect 9493 3375 9527 3390
rect 9561 3375 9595 3390
rect 9223 3356 9255 3375
rect 9296 3356 9323 3375
rect 9370 3356 9391 3375
rect 9444 3356 9459 3375
rect 9518 3356 9527 3375
rect 9592 3356 9595 3375
rect 9629 3375 9663 3390
rect 9697 3375 9731 3390
rect 9765 3375 9799 3390
rect 9833 3375 9867 3390
rect 9901 3375 9935 3390
rect 9969 3375 10003 3390
rect 9629 3356 9632 3375
rect 9697 3356 9706 3375
rect 9765 3356 9780 3375
rect 9833 3356 9854 3375
rect 9901 3356 9928 3375
rect 9969 3356 10002 3375
rect 10037 3356 10071 3390
rect 10105 3375 10139 3390
rect 10173 3375 10207 3390
rect 10241 3375 10312 3390
rect 10346 3375 10380 3391
rect 10414 3375 10448 3391
rect 10110 3356 10139 3375
rect 10184 3356 10207 3375
rect 8643 3341 8824 3356
rect 8858 3341 8897 3356
rect 8931 3341 8970 3356
rect 9004 3341 9043 3356
rect 9077 3341 9116 3356
rect 9150 3341 9189 3356
rect 9223 3341 9262 3356
rect 9296 3341 9336 3356
rect 9370 3341 9410 3356
rect 9444 3341 9484 3356
rect 9518 3341 9558 3356
rect 9592 3341 9632 3356
rect 9666 3341 9706 3356
rect 9740 3341 9780 3356
rect 9814 3341 9854 3356
rect 9888 3341 9928 3356
rect 9962 3341 10002 3356
rect 10036 3341 10076 3356
rect 10110 3341 10150 3356
rect 10184 3341 10224 3356
rect 10258 3341 10298 3375
rect 10346 3357 10372 3375
rect 10414 3357 10446 3375
rect 10482 3357 10516 3391
rect 10550 3375 10584 3391
rect 10618 3375 10652 3391
rect 10686 3375 10720 3391
rect 10754 3375 10788 3391
rect 10822 3375 10856 3391
rect 10554 3357 10584 3375
rect 10628 3357 10652 3375
rect 10702 3357 10720 3375
rect 10776 3357 10788 3375
rect 10850 3357 10856 3375
rect 10890 3375 10924 3391
rect 10332 3341 10372 3357
rect 10406 3341 10446 3357
rect 10480 3341 10520 3357
rect 10554 3341 10594 3357
rect 10628 3341 10668 3357
rect 10702 3341 10742 3357
rect 10776 3341 10816 3357
rect 10850 3341 10890 3357
rect 10958 3375 10992 3391
rect 11026 3375 11060 3391
rect 11094 3375 11128 3391
rect 11162 3375 11196 3391
rect 11230 3375 11264 3391
rect 10958 3357 10964 3375
rect 11026 3357 11038 3375
rect 11094 3357 11112 3375
rect 11162 3357 11186 3375
rect 11230 3357 11260 3375
rect 11298 3357 11332 3391
rect 11366 3375 11400 3391
rect 11434 3375 11468 3391
rect 11502 3375 11536 3391
rect 11570 3375 11590 3391
rect 11368 3357 11400 3375
rect 11442 3357 11468 3375
rect 11516 3357 11536 3375
rect 10924 3341 10964 3357
rect 10998 3341 11038 3357
rect 11072 3341 11112 3357
rect 11146 3341 11186 3357
rect 11220 3341 11260 3357
rect 11294 3341 11334 3357
rect 11368 3341 11408 3357
rect 11442 3341 11482 3357
rect 11516 3341 11556 3357
rect 8643 3321 11590 3341
rect 8643 3320 10312 3321
rect 8677 3286 8711 3320
rect 8745 3286 8779 3320
rect 8813 3303 8847 3320
rect 8881 3303 8915 3320
rect 8949 3303 8983 3320
rect 9017 3303 9051 3320
rect 9085 3303 9119 3320
rect 8813 3286 8824 3303
rect 8881 3286 8897 3303
rect 8949 3286 8970 3303
rect 9017 3286 9043 3303
rect 9085 3286 9116 3303
rect 9153 3286 9187 3320
rect 9221 3303 9255 3320
rect 9289 3303 9323 3320
rect 9357 3303 9391 3320
rect 9425 3303 9459 3320
rect 9493 3303 9527 3320
rect 9561 3303 9595 3320
rect 9223 3286 9255 3303
rect 9296 3286 9323 3303
rect 9370 3286 9391 3303
rect 9444 3286 9459 3303
rect 9518 3286 9527 3303
rect 9592 3286 9595 3303
rect 9629 3303 9663 3320
rect 9697 3303 9731 3320
rect 9765 3303 9799 3320
rect 9833 3303 9867 3320
rect 9901 3303 9935 3320
rect 9969 3303 10003 3320
rect 9629 3286 9632 3303
rect 9697 3286 9706 3303
rect 9765 3286 9780 3303
rect 9833 3286 9854 3303
rect 9901 3286 9928 3303
rect 9969 3286 10002 3303
rect 10037 3286 10071 3320
rect 10105 3303 10139 3320
rect 10173 3303 10207 3320
rect 10241 3303 10312 3320
rect 10346 3303 10380 3321
rect 10414 3303 10448 3321
rect 10110 3286 10139 3303
rect 10184 3286 10207 3303
rect 8643 3269 8824 3286
rect 8858 3269 8897 3286
rect 8931 3269 8970 3286
rect 9004 3269 9043 3286
rect 9077 3269 9116 3286
rect 9150 3269 9189 3286
rect 9223 3269 9262 3286
rect 9296 3269 9336 3286
rect 9370 3269 9410 3286
rect 9444 3269 9484 3286
rect 9518 3269 9558 3286
rect 9592 3269 9632 3286
rect 9666 3269 9706 3286
rect 9740 3269 9780 3286
rect 9814 3269 9854 3286
rect 9888 3269 9928 3286
rect 9962 3269 10002 3286
rect 10036 3269 10076 3286
rect 10110 3269 10150 3286
rect 10184 3269 10224 3286
rect 10258 3269 10298 3303
rect 10346 3287 10372 3303
rect 10414 3287 10446 3303
rect 10482 3287 10516 3321
rect 10550 3303 10584 3321
rect 10618 3303 10652 3321
rect 10686 3303 10720 3321
rect 10754 3303 10788 3321
rect 10822 3303 10856 3321
rect 10554 3287 10584 3303
rect 10628 3287 10652 3303
rect 10702 3287 10720 3303
rect 10776 3287 10788 3303
rect 10850 3287 10856 3303
rect 10890 3303 10924 3321
rect 10332 3269 10372 3287
rect 10406 3269 10446 3287
rect 10480 3269 10520 3287
rect 10554 3269 10594 3287
rect 10628 3269 10668 3287
rect 10702 3269 10742 3287
rect 10776 3269 10816 3287
rect 10850 3269 10890 3287
rect 10958 3303 10992 3321
rect 11026 3303 11060 3321
rect 11094 3303 11128 3321
rect 11162 3303 11196 3321
rect 11230 3303 11264 3321
rect 10958 3287 10964 3303
rect 11026 3287 11038 3303
rect 11094 3287 11112 3303
rect 11162 3287 11186 3303
rect 11230 3287 11260 3303
rect 11298 3287 11332 3321
rect 11366 3303 11400 3321
rect 11434 3303 11468 3321
rect 11502 3303 11536 3321
rect 11570 3303 11590 3321
rect 11368 3287 11400 3303
rect 11442 3287 11468 3303
rect 11516 3287 11536 3303
rect 10924 3269 10964 3287
rect 10998 3269 11038 3287
rect 11072 3269 11112 3287
rect 11146 3269 11186 3287
rect 11220 3269 11260 3287
rect 11294 3269 11334 3287
rect 11368 3269 11408 3287
rect 11442 3269 11482 3287
rect 11516 3269 11556 3287
rect 8643 3251 11590 3269
rect 8643 3250 10312 3251
rect 8677 3216 8711 3250
rect 8745 3216 8779 3250
rect 8813 3216 8847 3250
rect 8881 3216 8915 3250
rect 8949 3216 8983 3250
rect 9017 3216 9051 3250
rect 9085 3216 9119 3250
rect 9153 3216 9187 3250
rect 9221 3216 9255 3250
rect 9289 3216 9323 3250
rect 9357 3216 9391 3250
rect 9425 3216 9459 3250
rect 9493 3216 9527 3250
rect 9561 3216 9595 3250
rect 9629 3216 9663 3250
rect 9697 3216 9731 3250
rect 9765 3216 9799 3250
rect 9833 3216 9867 3250
rect 9901 3216 9935 3250
rect 9969 3216 10003 3250
rect 10037 3216 10071 3250
rect 10105 3216 10139 3250
rect 10173 3216 10207 3250
rect 10241 3217 10312 3250
rect 10346 3217 10380 3251
rect 10414 3217 10448 3251
rect 10482 3217 10516 3251
rect 10550 3217 10584 3251
rect 10618 3217 10652 3251
rect 10686 3217 10720 3251
rect 10754 3217 10788 3251
rect 10822 3217 10856 3251
rect 10890 3217 10924 3251
rect 10958 3217 10992 3251
rect 11026 3217 11060 3251
rect 11094 3217 11128 3251
rect 11162 3217 11196 3251
rect 11230 3217 11264 3251
rect 11298 3217 11332 3251
rect 11366 3217 11400 3251
rect 11434 3217 11468 3251
rect 11502 3217 11536 3251
rect 11570 3241 11590 3251
rect 12582 3471 16424 3475
rect 12582 3437 12594 3471
rect 12628 3453 12667 3471
rect 12701 3453 12740 3471
rect 12774 3453 12813 3471
rect 12847 3453 12886 3471
rect 12920 3453 12959 3471
rect 12993 3453 13032 3471
rect 13066 3453 13105 3471
rect 12582 3419 12595 3437
rect 12629 3419 12663 3453
rect 12701 3437 12731 3453
rect 12774 3437 12799 3453
rect 12847 3437 12867 3453
rect 12920 3437 12935 3453
rect 12993 3437 13003 3453
rect 13066 3437 13071 3453
rect 12697 3419 12731 3437
rect 12765 3419 12799 3437
rect 12833 3419 12867 3437
rect 12901 3419 12935 3437
rect 12969 3419 13003 3437
rect 13037 3419 13071 3437
rect 13139 3453 13178 3471
rect 13212 3453 13251 3471
rect 13285 3453 13324 3471
rect 13358 3453 13397 3471
rect 13105 3419 13139 3437
rect 13173 3437 13178 3453
rect 13241 3437 13251 3453
rect 13309 3437 13324 3453
rect 13377 3437 13397 3453
rect 13431 3437 13470 3471
rect 13504 3437 13543 3471
rect 13577 3437 13616 3471
rect 13650 3437 13689 3471
rect 13723 3437 13762 3471
rect 13796 3437 13835 3471
rect 13869 3437 13908 3471
rect 13942 3437 13981 3471
rect 14015 3437 14054 3471
rect 14088 3437 14127 3471
rect 14161 3437 14200 3471
rect 14234 3437 14273 3471
rect 14307 3437 14346 3471
rect 14380 3437 14419 3471
rect 14453 3437 14492 3471
rect 14526 3437 14565 3471
rect 14599 3437 14638 3471
rect 14672 3437 14711 3471
rect 14745 3437 14784 3471
rect 14818 3437 14857 3471
rect 14891 3437 14930 3471
rect 14964 3437 15003 3471
rect 15037 3437 15076 3471
rect 15110 3437 15149 3471
rect 15183 3437 15222 3471
rect 15256 3437 15295 3471
rect 15329 3437 15368 3471
rect 15402 3437 15441 3471
rect 15475 3437 15514 3471
rect 15548 3437 15587 3471
rect 15621 3437 15660 3471
rect 15694 3437 15733 3471
rect 15767 3437 15806 3471
rect 15840 3437 15879 3471
rect 15913 3437 15952 3471
rect 15986 3437 16025 3471
rect 16059 3437 16098 3471
rect 16132 3437 16171 3471
rect 16205 3437 16244 3471
rect 16278 3437 16317 3471
rect 16351 3437 16390 3471
rect 13173 3419 13207 3437
rect 13241 3419 13275 3437
rect 13309 3419 13343 3437
rect 13377 3419 16424 3437
rect 12582 3399 16424 3419
rect 12582 3365 12594 3399
rect 12628 3383 12667 3399
rect 12701 3383 12740 3399
rect 12774 3383 12813 3399
rect 12847 3383 12886 3399
rect 12920 3383 12959 3399
rect 12993 3383 13032 3399
rect 13066 3383 13105 3399
rect 12582 3349 12595 3365
rect 12629 3349 12663 3383
rect 12701 3365 12731 3383
rect 12774 3365 12799 3383
rect 12847 3365 12867 3383
rect 12920 3365 12935 3383
rect 12993 3365 13003 3383
rect 13066 3365 13071 3383
rect 12697 3349 12731 3365
rect 12765 3349 12799 3365
rect 12833 3349 12867 3365
rect 12901 3349 12935 3365
rect 12969 3349 13003 3365
rect 13037 3349 13071 3365
rect 13139 3383 13178 3399
rect 13212 3383 13251 3399
rect 13285 3383 13324 3399
rect 13358 3383 13397 3399
rect 13105 3349 13139 3365
rect 13173 3365 13178 3383
rect 13241 3365 13251 3383
rect 13309 3365 13324 3383
rect 13377 3365 13397 3383
rect 13431 3365 13470 3399
rect 13504 3365 13543 3399
rect 13577 3365 13616 3399
rect 13650 3365 13689 3399
rect 13723 3365 13762 3399
rect 13796 3365 13835 3399
rect 13869 3365 13908 3399
rect 13942 3365 13981 3399
rect 14015 3365 14054 3399
rect 14088 3365 14127 3399
rect 14161 3365 14200 3399
rect 14234 3365 14273 3399
rect 14307 3365 14346 3399
rect 14380 3365 14419 3399
rect 14453 3365 14492 3399
rect 14526 3365 14565 3399
rect 14599 3365 14638 3399
rect 14672 3365 14711 3399
rect 14745 3365 14784 3399
rect 14818 3365 14857 3399
rect 14891 3365 14930 3399
rect 14964 3365 15003 3399
rect 15037 3365 15076 3399
rect 15110 3365 15149 3399
rect 15183 3365 15222 3399
rect 15256 3365 15295 3399
rect 15329 3365 15368 3399
rect 15402 3365 15441 3399
rect 15475 3365 15514 3399
rect 15548 3365 15587 3399
rect 15621 3365 15660 3399
rect 15694 3365 15733 3399
rect 15767 3365 15806 3399
rect 15840 3365 15879 3399
rect 15913 3365 15952 3399
rect 15986 3365 16025 3399
rect 16059 3365 16098 3399
rect 16132 3365 16171 3399
rect 16205 3365 16244 3399
rect 16278 3365 16317 3399
rect 16351 3365 16390 3399
rect 13173 3349 13207 3365
rect 13241 3349 13275 3365
rect 13309 3349 13343 3365
rect 13377 3349 16424 3365
rect 12582 3327 16424 3349
rect 12582 3293 12594 3327
rect 12628 3313 12667 3327
rect 12701 3313 12740 3327
rect 12774 3313 12813 3327
rect 12847 3313 12886 3327
rect 12920 3313 12959 3327
rect 12993 3313 13032 3327
rect 13066 3313 13105 3327
rect 12582 3279 12595 3293
rect 12629 3279 12663 3313
rect 12701 3293 12731 3313
rect 12774 3293 12799 3313
rect 12847 3293 12867 3313
rect 12920 3293 12935 3313
rect 12993 3293 13003 3313
rect 13066 3293 13071 3313
rect 12697 3279 12731 3293
rect 12765 3279 12799 3293
rect 12833 3279 12867 3293
rect 12901 3279 12935 3293
rect 12969 3279 13003 3293
rect 13037 3279 13071 3293
rect 13139 3313 13178 3327
rect 13212 3313 13251 3327
rect 13285 3313 13324 3327
rect 13358 3313 13397 3327
rect 13105 3279 13139 3293
rect 13173 3293 13178 3313
rect 13241 3293 13251 3313
rect 13309 3293 13324 3313
rect 13377 3293 13397 3313
rect 13431 3293 13470 3327
rect 13504 3293 13543 3327
rect 13577 3293 13616 3327
rect 13650 3293 13689 3327
rect 13723 3293 13762 3327
rect 13796 3293 13835 3327
rect 13869 3293 13908 3327
rect 13942 3293 13981 3327
rect 14015 3293 14054 3327
rect 14088 3293 14127 3327
rect 14161 3293 14200 3327
rect 14234 3293 14273 3327
rect 14307 3293 14346 3327
rect 14380 3293 14419 3327
rect 14453 3293 14492 3327
rect 14526 3293 14565 3327
rect 14599 3293 14638 3327
rect 14672 3293 14711 3327
rect 14745 3293 14784 3327
rect 14818 3293 14857 3327
rect 14891 3293 14930 3327
rect 14964 3293 15003 3327
rect 15037 3293 15076 3327
rect 15110 3293 15149 3327
rect 15183 3293 15222 3327
rect 15256 3293 15295 3327
rect 15329 3293 15368 3327
rect 15402 3293 15441 3327
rect 15475 3293 15514 3327
rect 15548 3293 15587 3327
rect 15621 3293 15660 3327
rect 15694 3293 15733 3327
rect 15767 3293 15806 3327
rect 15840 3293 15879 3327
rect 15913 3293 15952 3327
rect 15986 3293 16025 3327
rect 16059 3293 16098 3327
rect 16132 3293 16171 3327
rect 16205 3293 16244 3327
rect 16278 3293 16317 3327
rect 16351 3293 16390 3327
rect 13173 3279 13207 3293
rect 13241 3279 13275 3293
rect 13309 3279 13343 3293
rect 13377 3279 16424 3293
rect 12582 3255 16424 3279
rect 11570 3217 11589 3241
rect 10241 3216 11589 3217
rect 8643 3181 11589 3216
rect 8643 3180 10312 3181
rect 8677 3146 8711 3180
rect 8745 3146 8779 3180
rect 8813 3146 8847 3180
rect 8881 3146 8915 3180
rect 8949 3146 8983 3180
rect 9017 3146 9051 3180
rect 9085 3146 9119 3180
rect 9153 3146 9187 3180
rect 9221 3146 9255 3180
rect 9289 3146 9323 3180
rect 9357 3146 9391 3180
rect 9425 3146 9459 3180
rect 9493 3146 9527 3180
rect 9561 3146 9595 3180
rect 9629 3146 9663 3180
rect 9697 3146 9731 3180
rect 9765 3146 9799 3180
rect 9833 3146 9867 3180
rect 9901 3146 9935 3180
rect 9969 3146 10003 3180
rect 10037 3146 10071 3180
rect 10105 3146 10139 3180
rect 10173 3146 10207 3180
rect 10241 3147 10312 3180
rect 10346 3147 10380 3181
rect 10414 3147 10448 3181
rect 10482 3147 10516 3181
rect 10550 3147 10584 3181
rect 10618 3147 10652 3181
rect 10686 3147 10720 3181
rect 10754 3147 10788 3181
rect 10822 3147 10856 3181
rect 10890 3147 10924 3181
rect 10958 3147 10992 3181
rect 11026 3147 11060 3181
rect 11094 3147 11128 3181
rect 11162 3147 11196 3181
rect 11230 3147 11264 3181
rect 11298 3147 11332 3181
rect 11366 3147 11400 3181
rect 11434 3147 11468 3181
rect 11502 3147 11536 3181
rect 11570 3147 11589 3181
rect 10241 3146 11589 3147
rect 8643 3111 11589 3146
rect 8643 3110 10312 3111
rect 8677 3076 8711 3110
rect 8745 3076 8779 3110
rect 8813 3076 8847 3110
rect 8881 3076 8915 3110
rect 8949 3076 8983 3110
rect 9017 3076 9051 3110
rect 9085 3076 9119 3110
rect 9153 3076 9187 3110
rect 9221 3076 9255 3110
rect 9289 3076 9323 3110
rect 9357 3076 9391 3110
rect 9425 3076 9459 3110
rect 9493 3076 9527 3110
rect 9561 3076 9595 3110
rect 9629 3076 9663 3110
rect 9697 3076 9731 3110
rect 9765 3076 9799 3110
rect 9833 3076 9867 3110
rect 9901 3076 9935 3110
rect 9969 3076 10003 3110
rect 10037 3076 10071 3110
rect 10105 3076 10139 3110
rect 10173 3076 10207 3110
rect 10241 3077 10312 3110
rect 10346 3077 10380 3111
rect 10414 3077 10448 3111
rect 10482 3077 10516 3111
rect 10550 3077 10584 3111
rect 10618 3077 10652 3111
rect 10686 3077 10720 3111
rect 10754 3077 10788 3111
rect 10822 3077 10856 3111
rect 10890 3077 10924 3111
rect 10958 3077 10992 3111
rect 11026 3077 11060 3111
rect 11094 3077 11128 3111
rect 11162 3077 11196 3111
rect 11230 3077 11264 3111
rect 11298 3077 11332 3111
rect 11366 3077 11400 3111
rect 11434 3077 11468 3111
rect 11502 3077 11536 3111
rect 11570 3077 11589 3111
rect 10241 3076 11589 3077
rect 8643 3041 11589 3076
rect 8643 3040 10312 3041
rect 8677 3006 8711 3040
rect 8745 3006 8779 3040
rect 8813 3006 8847 3040
rect 8881 3006 8915 3040
rect 8949 3006 8983 3040
rect 9017 3006 9051 3040
rect 9085 3006 9119 3040
rect 9153 3006 9187 3040
rect 9221 3006 9255 3040
rect 9289 3006 9323 3040
rect 9357 3006 9391 3040
rect 9425 3006 9459 3040
rect 9493 3006 9527 3040
rect 9561 3006 9595 3040
rect 9629 3006 9663 3040
rect 9697 3006 9731 3040
rect 9765 3006 9799 3040
rect 9833 3006 9867 3040
rect 9901 3006 9935 3040
rect 9969 3006 10003 3040
rect 10037 3006 10071 3040
rect 10105 3006 10139 3040
rect 10173 3006 10207 3040
rect 10241 3007 10312 3040
rect 10346 3007 10380 3041
rect 10414 3007 10448 3041
rect 10482 3007 10516 3041
rect 10550 3007 10584 3041
rect 10618 3007 10652 3041
rect 10686 3007 10720 3041
rect 10754 3007 10788 3041
rect 10822 3007 10856 3041
rect 10890 3007 10924 3041
rect 10958 3007 10992 3041
rect 11026 3007 11060 3041
rect 11094 3007 11128 3041
rect 11162 3007 11196 3041
rect 11230 3007 11264 3041
rect 11298 3007 11332 3041
rect 11366 3007 11400 3041
rect 11434 3007 11468 3041
rect 11502 3007 11536 3041
rect 11570 3007 11589 3041
rect 10241 3006 11589 3007
rect 8643 2971 11589 3006
rect 8643 2970 10312 2971
rect 8677 2936 8711 2970
rect 8745 2936 8779 2970
rect 8813 2936 8847 2970
rect 8881 2936 8915 2970
rect 8949 2936 8983 2970
rect 9017 2936 9051 2970
rect 9085 2936 9119 2970
rect 9153 2936 9187 2970
rect 9221 2936 9255 2970
rect 9289 2936 9323 2970
rect 9357 2936 9391 2970
rect 9425 2936 9459 2970
rect 9493 2936 9527 2970
rect 9561 2936 9595 2970
rect 9629 2936 9663 2970
rect 9697 2936 9731 2970
rect 9765 2936 9799 2970
rect 9833 2936 9867 2970
rect 9901 2936 9935 2970
rect 9969 2936 10003 2970
rect 10037 2936 10071 2970
rect 10105 2936 10139 2970
rect 10173 2936 10207 2970
rect 10241 2937 10312 2970
rect 10346 2937 10380 2971
rect 10414 2937 10448 2971
rect 10482 2937 10516 2971
rect 10550 2937 10584 2971
rect 10618 2937 10652 2971
rect 10686 2937 10720 2971
rect 10754 2937 10788 2971
rect 10822 2937 10856 2971
rect 10890 2937 10924 2971
rect 10958 2937 10992 2971
rect 11026 2937 11060 2971
rect 11094 2937 11128 2971
rect 11162 2937 11196 2971
rect 11230 2937 11264 2971
rect 11298 2937 11332 2971
rect 11366 2937 11400 2971
rect 11434 2937 11468 2971
rect 11502 2937 11536 2971
rect 11570 2937 11589 2971
rect 12582 3221 12594 3255
rect 12628 3243 12667 3255
rect 12701 3243 12740 3255
rect 12774 3243 12813 3255
rect 12847 3243 12886 3255
rect 12920 3243 12959 3255
rect 12993 3243 13032 3255
rect 13066 3243 13105 3255
rect 12582 3209 12595 3221
rect 12629 3209 12663 3243
rect 12701 3221 12731 3243
rect 12774 3221 12799 3243
rect 12847 3221 12867 3243
rect 12920 3221 12935 3243
rect 12993 3221 13003 3243
rect 13066 3221 13071 3243
rect 12697 3209 12731 3221
rect 12765 3209 12799 3221
rect 12833 3209 12867 3221
rect 12901 3209 12935 3221
rect 12969 3209 13003 3221
rect 13037 3209 13071 3221
rect 13139 3243 13178 3255
rect 13212 3243 13251 3255
rect 13285 3243 13324 3255
rect 13358 3243 13397 3255
rect 13105 3209 13139 3221
rect 13173 3221 13178 3243
rect 13241 3221 13251 3243
rect 13309 3221 13324 3243
rect 13377 3221 13397 3243
rect 13431 3221 13470 3255
rect 13504 3221 13543 3255
rect 13577 3221 13616 3255
rect 13650 3221 13689 3255
rect 13723 3221 13762 3255
rect 13796 3221 13835 3255
rect 13869 3221 13908 3255
rect 13942 3221 13981 3255
rect 14015 3221 14054 3255
rect 14088 3221 14127 3255
rect 14161 3221 14200 3255
rect 14234 3221 14273 3255
rect 14307 3221 14346 3255
rect 14380 3221 14419 3255
rect 14453 3221 14492 3255
rect 14526 3221 14565 3255
rect 14599 3221 14638 3255
rect 14672 3221 14711 3255
rect 14745 3221 14784 3255
rect 14818 3221 14857 3255
rect 14891 3221 14930 3255
rect 14964 3221 15003 3255
rect 15037 3221 15076 3255
rect 15110 3221 15149 3255
rect 15183 3221 15222 3255
rect 15256 3221 15295 3255
rect 15329 3221 15368 3255
rect 15402 3221 15441 3255
rect 15475 3221 15514 3255
rect 15548 3221 15587 3255
rect 15621 3221 15660 3255
rect 15694 3221 15733 3255
rect 15767 3221 15806 3255
rect 15840 3221 15879 3255
rect 15913 3221 15952 3255
rect 15986 3221 16025 3255
rect 16059 3221 16098 3255
rect 16132 3221 16171 3255
rect 16205 3221 16244 3255
rect 16278 3221 16317 3255
rect 16351 3221 16390 3255
rect 13173 3209 13207 3221
rect 13241 3209 13275 3221
rect 13309 3209 13343 3221
rect 13377 3217 16424 3221
rect 23568 3449 23597 3488
rect 23767 3449 23796 3488
rect 23568 3415 23593 3449
rect 23771 3415 23796 3449
rect 23568 3376 23597 3415
rect 23767 3376 23796 3415
rect 23568 3342 23593 3376
rect 23771 3342 23796 3376
rect 23568 3303 23597 3342
rect 23767 3303 23796 3342
rect 23568 3269 23593 3303
rect 23771 3269 23796 3303
rect 23568 3230 23597 3269
rect 23767 3230 23796 3269
rect 13377 3209 13390 3217
rect 12582 3173 13390 3209
rect 12582 3139 12595 3173
rect 12629 3139 12663 3173
rect 12697 3139 12731 3173
rect 12765 3139 12799 3173
rect 12833 3139 12867 3173
rect 12901 3139 12935 3173
rect 12969 3139 13003 3173
rect 13037 3139 13071 3173
rect 13105 3139 13139 3173
rect 13173 3139 13207 3173
rect 13241 3139 13275 3173
rect 13309 3139 13343 3173
rect 13377 3139 13390 3173
rect 12582 3103 13390 3139
rect 12582 3069 12595 3103
rect 12629 3069 12663 3103
rect 12697 3069 12731 3103
rect 12765 3069 12799 3103
rect 12833 3069 12867 3103
rect 12901 3069 12935 3103
rect 12969 3069 13003 3103
rect 13037 3069 13071 3103
rect 13105 3069 13139 3103
rect 13173 3069 13207 3103
rect 13241 3069 13275 3103
rect 13309 3069 13343 3103
rect 13377 3069 13390 3103
rect 12582 3033 13390 3069
rect 12582 2999 12595 3033
rect 12629 2999 12663 3033
rect 12697 2999 12731 3033
rect 12765 2999 12799 3033
rect 12833 2999 12867 3033
rect 12901 2999 12935 3033
rect 12969 2999 13003 3033
rect 13037 2999 13071 3033
rect 13105 2999 13139 3033
rect 13173 2999 13207 3033
rect 13241 2999 13275 3033
rect 13309 2999 13343 3033
rect 13377 2999 13390 3033
rect 12582 2964 13390 2999
rect 10241 2936 11589 2937
rect 8643 2901 11589 2936
rect 11684 2914 12488 2959
rect 12582 2930 12595 2964
rect 12629 2930 12663 2964
rect 12697 2930 12731 2964
rect 12765 2930 12799 2964
rect 12833 2930 12867 2964
rect 12901 2930 12935 2964
rect 12969 2930 13003 2964
rect 13037 2930 13071 2964
rect 13105 2930 13139 2964
rect 13173 2930 13207 2964
rect 13241 2930 13275 2964
rect 13309 2930 13343 2964
rect 13377 2930 13390 2964
rect 8643 2900 10312 2901
rect 8677 2866 8711 2900
rect 8745 2866 8779 2900
rect 8813 2866 8847 2900
rect 8881 2866 8915 2900
rect 8949 2866 8983 2900
rect 9017 2866 9051 2900
rect 9085 2866 9119 2900
rect 9153 2866 9187 2900
rect 9221 2866 9255 2900
rect 9289 2866 9323 2900
rect 9357 2866 9391 2900
rect 9425 2866 9459 2900
rect 9493 2866 9527 2900
rect 9561 2866 9595 2900
rect 9629 2866 9663 2900
rect 9697 2866 9731 2900
rect 9765 2866 9799 2900
rect 9833 2866 9867 2900
rect 9901 2866 9935 2900
rect 9969 2866 10003 2900
rect 10037 2866 10071 2900
rect 10105 2866 10139 2900
rect 10173 2866 10207 2900
rect 10241 2867 10312 2900
rect 10346 2867 10380 2901
rect 10414 2867 10448 2901
rect 10482 2867 10516 2901
rect 10550 2867 10584 2901
rect 10618 2867 10652 2901
rect 10686 2867 10720 2901
rect 10754 2867 10788 2901
rect 10822 2867 10856 2901
rect 10890 2867 10924 2901
rect 10958 2867 10992 2901
rect 11026 2867 11060 2901
rect 11094 2867 11128 2901
rect 11162 2867 11196 2901
rect 11230 2867 11264 2901
rect 11298 2867 11332 2901
rect 11366 2867 11400 2901
rect 11434 2867 11468 2901
rect 11502 2867 11536 2901
rect 11570 2867 11589 2901
rect 10241 2866 11589 2867
rect 8643 2831 11589 2866
rect 8643 2830 10312 2831
rect 8677 2796 8711 2830
rect 8745 2796 8779 2830
rect 8813 2796 8847 2830
rect 8881 2796 8915 2830
rect 8949 2796 8983 2830
rect 9017 2796 9051 2830
rect 9085 2796 9119 2830
rect 9153 2796 9187 2830
rect 9221 2796 9255 2830
rect 9289 2796 9323 2830
rect 9357 2796 9391 2830
rect 9425 2796 9459 2830
rect 9493 2796 9527 2830
rect 9561 2796 9595 2830
rect 9629 2796 9663 2830
rect 9697 2796 9731 2830
rect 9765 2796 9799 2830
rect 9833 2796 9867 2830
rect 9901 2796 9935 2830
rect 9969 2796 10003 2830
rect 10037 2796 10071 2830
rect 10105 2796 10139 2830
rect 10173 2796 10207 2830
rect 10241 2797 10312 2830
rect 10346 2797 10380 2831
rect 10414 2797 10448 2831
rect 10482 2797 10516 2831
rect 10550 2797 10584 2831
rect 10618 2797 10652 2831
rect 10686 2797 10720 2831
rect 10754 2797 10788 2831
rect 10822 2797 10856 2831
rect 10890 2797 10924 2831
rect 10958 2797 10992 2831
rect 11026 2797 11060 2831
rect 11094 2797 11128 2831
rect 11162 2797 11196 2831
rect 11230 2797 11264 2831
rect 11298 2797 11332 2831
rect 11366 2797 11400 2831
rect 11434 2797 11468 2831
rect 11502 2797 11536 2831
rect 11570 2797 11589 2831
rect 10241 2796 11589 2797
rect 8643 2761 11589 2796
rect 8677 2727 8711 2761
rect 8745 2727 8779 2761
rect 8813 2727 8847 2761
rect 8881 2727 8915 2761
rect 8949 2727 8983 2761
rect 9017 2727 9051 2761
rect 9085 2727 9119 2761
rect 9153 2727 9187 2761
rect 9221 2727 9255 2761
rect 9289 2727 9323 2761
rect 9357 2727 9391 2761
rect 9425 2727 9459 2761
rect 9493 2727 9527 2761
rect 9561 2727 9595 2761
rect 9629 2727 9663 2761
rect 9697 2727 9731 2761
rect 9765 2727 9799 2761
rect 9833 2727 9867 2761
rect 9901 2727 9935 2761
rect 9969 2727 10003 2761
rect 10037 2727 10071 2761
rect 10105 2727 10139 2761
rect 10173 2727 10207 2761
rect 10241 2727 10312 2761
rect 10346 2727 10380 2761
rect 10414 2727 10448 2761
rect 10482 2727 10516 2761
rect 10550 2727 10584 2761
rect 10618 2727 10652 2761
rect 10686 2727 10720 2761
rect 10754 2727 10788 2761
rect 10822 2727 10856 2761
rect 10890 2727 10924 2761
rect 10958 2727 10992 2761
rect 11026 2727 11060 2761
rect 11094 2727 11128 2761
rect 11162 2727 11196 2761
rect 11230 2727 11264 2761
rect 11298 2727 11332 2761
rect 11366 2727 11400 2761
rect 11434 2727 11468 2761
rect 11502 2727 11536 2761
rect 11570 2730 11589 2761
rect 12582 2895 13390 2930
rect 12582 2861 12595 2895
rect 12629 2861 12663 2895
rect 12697 2861 12731 2895
rect 12765 2861 12799 2895
rect 12833 2861 12867 2895
rect 12901 2861 12935 2895
rect 12969 2861 13003 2895
rect 13037 2861 13071 2895
rect 13105 2861 13139 2895
rect 13173 2861 13207 2895
rect 13241 2861 13275 2895
rect 13309 2861 13343 2895
rect 13377 2861 13390 2895
rect 12582 2826 13390 2861
rect 12582 2792 12595 2826
rect 12629 2792 12663 2826
rect 12697 2792 12731 2826
rect 12765 2792 12799 2826
rect 12833 2792 12867 2826
rect 12901 2792 12935 2826
rect 12969 2792 13003 2826
rect 13037 2792 13071 2826
rect 13105 2792 13139 2826
rect 13173 2792 13207 2826
rect 13241 2792 13275 2826
rect 13309 2792 13343 2826
rect 13377 2792 13390 2826
rect 12582 2757 13390 2792
rect 12582 2730 12595 2757
rect 11570 2727 12595 2730
rect 8643 2702 12595 2727
rect 13377 2730 13390 2757
rect 23568 3196 23593 3230
rect 23771 3196 23796 3230
rect 23568 3156 23597 3196
rect 23767 3156 23796 3196
rect 23568 3122 23593 3156
rect 23771 3122 23796 3156
rect 23568 3082 23597 3122
rect 23767 3082 23796 3122
rect 23568 3048 23593 3082
rect 23771 3048 23796 3082
rect 23568 3008 23597 3048
rect 23767 3008 23796 3048
rect 23568 2974 23593 3008
rect 23771 2974 23796 3008
rect 23568 2934 23597 2974
rect 23767 2934 23796 2974
rect 23568 2900 23593 2934
rect 23771 2900 23796 2934
rect 23568 2860 23597 2900
rect 23767 2860 23796 2900
rect 23568 2826 23593 2860
rect 23771 2826 23796 2860
rect 23568 2786 23597 2826
rect 23767 2786 23796 2826
rect 23568 2752 23593 2786
rect 23771 2752 23796 2786
rect 13377 2723 13458 2730
rect 8643 2692 11198 2702
rect 11232 2692 11272 2702
rect 11306 2692 11346 2702
rect 11380 2692 11420 2702
rect 11454 2692 11494 2702
rect 11528 2692 11568 2702
rect 8677 2658 8711 2692
rect 8745 2658 8779 2692
rect 8813 2658 8847 2692
rect 8881 2658 8915 2692
rect 8949 2658 8983 2692
rect 9017 2658 9051 2692
rect 9085 2658 9119 2692
rect 9153 2658 9187 2692
rect 9221 2658 9255 2692
rect 9289 2658 9323 2692
rect 9357 2658 9391 2692
rect 9425 2658 9459 2692
rect 9493 2658 9527 2692
rect 9561 2658 9595 2692
rect 9629 2658 9663 2692
rect 9697 2658 9731 2692
rect 9765 2658 9799 2692
rect 9833 2658 9867 2692
rect 9901 2658 9935 2692
rect 9969 2658 10003 2692
rect 10037 2658 10071 2692
rect 10105 2658 10139 2692
rect 10173 2658 10207 2692
rect 10241 2658 10312 2692
rect 10346 2658 10380 2692
rect 10414 2658 10448 2692
rect 10482 2658 10516 2692
rect 10550 2658 10584 2692
rect 10618 2658 10652 2692
rect 10686 2658 10720 2692
rect 10754 2658 10788 2692
rect 10822 2658 10856 2692
rect 10890 2658 10924 2692
rect 10958 2658 10992 2692
rect 11026 2658 11060 2692
rect 11094 2658 11128 2692
rect 11162 2658 11196 2692
rect 11232 2668 11264 2692
rect 11306 2668 11332 2692
rect 11380 2668 11400 2692
rect 11454 2668 11468 2692
rect 11528 2668 11536 2692
rect 11602 2668 11642 2702
rect 11676 2699 11716 2702
rect 11750 2699 11790 2702
rect 11824 2699 11864 2702
rect 11898 2699 11938 2702
rect 11972 2699 12012 2702
rect 12046 2699 12087 2702
rect 12121 2699 12162 2702
rect 11686 2668 11716 2699
rect 11230 2658 11264 2668
rect 11298 2658 11332 2668
rect 11366 2658 11400 2668
rect 11434 2658 11468 2668
rect 11502 2658 11536 2668
rect 11570 2665 11652 2668
rect 11686 2665 11720 2668
rect 11754 2665 11788 2699
rect 11824 2668 11856 2699
rect 11898 2668 11924 2699
rect 11972 2668 11992 2699
rect 12046 2668 12060 2699
rect 12121 2668 12128 2699
rect 11822 2665 11856 2668
rect 11890 2665 11924 2668
rect 11958 2665 11992 2668
rect 12026 2665 12060 2668
rect 12094 2665 12128 2668
rect 12196 2699 12237 2702
rect 12271 2699 12312 2702
rect 12346 2699 12387 2702
rect 12421 2699 12462 2702
rect 12496 2699 12537 2702
rect 12162 2665 12196 2668
rect 12230 2668 12237 2699
rect 12298 2668 12312 2699
rect 12366 2668 12387 2699
rect 12434 2668 12462 2699
rect 12502 2668 12537 2699
rect 12571 2689 12595 2702
rect 12571 2668 12573 2689
rect 12230 2665 12264 2668
rect 12298 2665 12332 2668
rect 12366 2665 12400 2668
rect 12434 2665 12468 2668
rect 12502 2665 12573 2668
rect 11570 2658 12573 2665
rect 8643 2655 12573 2658
rect 13355 2655 13458 2723
rect 8643 2630 13458 2655
rect 8643 2623 11198 2630
rect 11232 2623 11272 2630
rect 11306 2623 11346 2630
rect 11380 2623 11420 2630
rect 11454 2623 11494 2630
rect 11528 2623 11568 2630
rect 8677 2589 8711 2623
rect 8745 2589 8779 2623
rect 8813 2589 8847 2623
rect 8881 2589 8915 2623
rect 8949 2589 8983 2623
rect 9017 2589 9051 2623
rect 9085 2589 9119 2623
rect 9153 2589 9187 2623
rect 9221 2589 9255 2623
rect 9289 2589 9323 2623
rect 9357 2589 9391 2623
rect 9425 2589 9459 2623
rect 9493 2589 9527 2623
rect 9561 2589 9595 2623
rect 9629 2589 9663 2623
rect 9697 2589 9731 2623
rect 9765 2589 9799 2623
rect 9833 2589 9867 2623
rect 9901 2589 9935 2623
rect 9969 2589 10003 2623
rect 10037 2589 10071 2623
rect 10105 2589 10139 2623
rect 10173 2589 10207 2623
rect 10241 2589 10312 2623
rect 10346 2589 10380 2623
rect 10414 2589 10448 2623
rect 10482 2589 10516 2623
rect 10550 2589 10584 2623
rect 10618 2589 10652 2623
rect 10686 2589 10720 2623
rect 10754 2589 10788 2623
rect 10822 2589 10856 2623
rect 10890 2589 10924 2623
rect 10958 2589 10992 2623
rect 11026 2589 11060 2623
rect 11094 2589 11128 2623
rect 11162 2589 11196 2623
rect 11232 2596 11264 2623
rect 11306 2596 11332 2623
rect 11380 2596 11400 2623
rect 11454 2596 11468 2623
rect 11528 2596 11536 2623
rect 11602 2596 11642 2630
rect 11676 2629 11716 2630
rect 11750 2629 11790 2630
rect 11824 2629 11864 2630
rect 11898 2629 11938 2630
rect 11972 2629 12012 2630
rect 12046 2629 12087 2630
rect 12121 2629 12162 2630
rect 11686 2596 11716 2629
rect 11230 2589 11264 2596
rect 11298 2589 11332 2596
rect 11366 2589 11400 2596
rect 11434 2589 11468 2596
rect 11502 2589 11536 2596
rect 11570 2595 11652 2596
rect 11686 2595 11720 2596
rect 11754 2595 11788 2629
rect 11824 2596 11856 2629
rect 11898 2596 11924 2629
rect 11972 2596 11992 2629
rect 12046 2596 12060 2629
rect 12121 2596 12128 2629
rect 11822 2595 11856 2596
rect 11890 2595 11924 2596
rect 11958 2595 11992 2596
rect 12026 2595 12060 2596
rect 12094 2595 12128 2596
rect 12196 2629 12237 2630
rect 12271 2629 12312 2630
rect 12346 2629 12387 2630
rect 12421 2629 12462 2630
rect 12496 2629 12537 2630
rect 12162 2595 12196 2596
rect 12230 2596 12237 2629
rect 12298 2596 12312 2629
rect 12366 2596 12387 2629
rect 12434 2596 12462 2629
rect 12502 2596 12537 2629
rect 12571 2620 12612 2630
rect 12646 2620 12687 2630
rect 12721 2620 12762 2630
rect 12796 2620 12837 2630
rect 12871 2620 12912 2630
rect 12946 2620 12987 2630
rect 13021 2620 13062 2630
rect 13096 2620 13137 2630
rect 13171 2620 13212 2630
rect 13246 2620 13458 2630
rect 12571 2596 12573 2620
rect 12230 2595 12264 2596
rect 12298 2595 12332 2596
rect 12366 2595 12400 2596
rect 12434 2595 12468 2596
rect 12502 2595 12573 2596
rect 11570 2589 12573 2595
rect 8643 2586 12573 2589
rect 12607 2596 12612 2620
rect 12675 2596 12687 2620
rect 12743 2596 12762 2620
rect 12811 2596 12837 2620
rect 12879 2596 12912 2620
rect 12607 2586 12641 2596
rect 12675 2586 12709 2596
rect 12743 2586 12777 2596
rect 12811 2586 12845 2596
rect 12879 2586 12913 2596
rect 12947 2586 12981 2620
rect 13021 2596 13049 2620
rect 13096 2596 13117 2620
rect 13171 2596 13185 2620
rect 13246 2596 13253 2620
rect 13015 2586 13049 2596
rect 13083 2586 13117 2596
rect 13151 2586 13185 2596
rect 13219 2586 13253 2596
rect 13287 2586 13321 2620
rect 13355 2586 13458 2620
rect 8643 2559 13458 2586
rect 8643 2558 11652 2559
rect 11686 2558 11720 2559
rect 8643 2554 11198 2558
rect 11232 2554 11272 2558
rect 11306 2554 11346 2558
rect 11380 2554 11420 2558
rect 11454 2554 11494 2558
rect 11528 2554 11568 2558
rect 8677 2520 8711 2554
rect 8745 2520 8779 2554
rect 8813 2520 8847 2554
rect 8881 2520 8915 2554
rect 8949 2520 8983 2554
rect 9017 2520 9051 2554
rect 9085 2520 9119 2554
rect 9153 2520 9187 2554
rect 9221 2520 9255 2554
rect 9289 2520 9323 2554
rect 9357 2520 9391 2554
rect 9425 2520 9459 2554
rect 9493 2520 9527 2554
rect 9561 2520 9595 2554
rect 9629 2520 9663 2554
rect 9697 2520 9731 2554
rect 9765 2520 9799 2554
rect 9833 2520 9867 2554
rect 9901 2520 9935 2554
rect 9969 2520 10003 2554
rect 10037 2520 10071 2554
rect 10105 2520 10139 2554
rect 10173 2520 10207 2554
rect 10241 2520 10312 2554
rect 10346 2520 10380 2554
rect 10414 2520 10448 2554
rect 10482 2520 10516 2554
rect 10550 2520 10584 2554
rect 10618 2520 10652 2554
rect 10686 2520 10720 2554
rect 10754 2520 10788 2554
rect 10822 2520 10856 2554
rect 10890 2520 10924 2554
rect 10958 2520 10992 2554
rect 11026 2520 11060 2554
rect 11094 2520 11128 2554
rect 11162 2520 11196 2554
rect 11232 2524 11264 2554
rect 11306 2524 11332 2554
rect 11380 2524 11400 2554
rect 11454 2524 11468 2554
rect 11528 2524 11536 2554
rect 11602 2524 11642 2558
rect 11686 2525 11716 2558
rect 11754 2525 11788 2559
rect 11822 2558 11856 2559
rect 11890 2558 11924 2559
rect 11958 2558 11992 2559
rect 12026 2558 12060 2559
rect 12094 2558 12128 2559
rect 11824 2525 11856 2558
rect 11898 2525 11924 2558
rect 11972 2525 11992 2558
rect 12046 2525 12060 2558
rect 12121 2525 12128 2558
rect 12162 2558 12196 2559
rect 11676 2524 11716 2525
rect 11750 2524 11790 2525
rect 11824 2524 11864 2525
rect 11898 2524 11938 2525
rect 11972 2524 12012 2525
rect 12046 2524 12087 2525
rect 12121 2524 12162 2525
rect 12230 2558 12264 2559
rect 12298 2558 12332 2559
rect 12366 2558 12400 2559
rect 12434 2558 12468 2559
rect 12502 2558 13458 2559
rect 12230 2525 12237 2558
rect 12298 2525 12312 2558
rect 12366 2525 12387 2558
rect 12434 2525 12462 2558
rect 12502 2525 12537 2558
rect 12196 2524 12237 2525
rect 12271 2524 12312 2525
rect 12346 2524 12387 2525
rect 12421 2524 12462 2525
rect 12496 2524 12537 2525
rect 12571 2551 12612 2558
rect 12646 2551 12687 2558
rect 12721 2551 12762 2558
rect 12796 2551 12837 2558
rect 12871 2551 12912 2558
rect 12946 2551 12987 2558
rect 13021 2551 13062 2558
rect 13096 2551 13137 2558
rect 13171 2551 13212 2558
rect 13246 2551 13458 2558
rect 12571 2524 12573 2551
rect 11230 2520 11264 2524
rect 11298 2520 11332 2524
rect 11366 2520 11400 2524
rect 11434 2520 11468 2524
rect 11502 2520 11536 2524
rect 11570 2520 12573 2524
rect 8643 2517 12573 2520
rect 12607 2524 12612 2551
rect 12675 2524 12687 2551
rect 12743 2524 12762 2551
rect 12811 2524 12837 2551
rect 12879 2524 12912 2551
rect 12607 2517 12641 2524
rect 12675 2517 12709 2524
rect 12743 2517 12777 2524
rect 12811 2517 12845 2524
rect 12879 2517 12913 2524
rect 12947 2517 12981 2551
rect 13021 2524 13049 2551
rect 13096 2524 13117 2551
rect 13171 2524 13185 2551
rect 13246 2524 13253 2551
rect 13015 2517 13049 2524
rect 13083 2517 13117 2524
rect 13151 2517 13185 2524
rect 13219 2517 13253 2524
rect 13287 2517 13321 2551
rect 13355 2517 13458 2551
rect 8643 2489 13458 2517
rect 8643 2485 11652 2489
rect 8677 2451 8711 2485
rect 8745 2451 8779 2485
rect 8813 2451 8847 2485
rect 8881 2451 8915 2485
rect 8949 2451 8983 2485
rect 9017 2451 9051 2485
rect 9085 2451 9119 2485
rect 9153 2451 9187 2485
rect 9221 2451 9255 2485
rect 9289 2451 9323 2485
rect 9357 2451 9391 2485
rect 9425 2451 9459 2485
rect 9493 2451 9527 2485
rect 9561 2451 9595 2485
rect 9629 2451 9663 2485
rect 9697 2451 9731 2485
rect 9765 2451 9799 2485
rect 9833 2451 9867 2485
rect 9901 2451 9935 2485
rect 9969 2451 10003 2485
rect 10037 2451 10071 2485
rect 10105 2451 10139 2485
rect 10173 2451 10207 2485
rect 10241 2451 10312 2485
rect 10346 2451 10380 2485
rect 10414 2451 10448 2485
rect 10482 2451 10516 2485
rect 10550 2451 10584 2485
rect 10618 2451 10652 2485
rect 10686 2451 10720 2485
rect 10754 2451 10788 2485
rect 10822 2451 10856 2485
rect 10890 2451 10924 2485
rect 10958 2451 10992 2485
rect 11026 2451 11060 2485
rect 11094 2451 11128 2485
rect 11162 2451 11196 2485
rect 11230 2451 11264 2485
rect 11298 2451 11332 2485
rect 11366 2451 11400 2485
rect 11434 2451 11468 2485
rect 11502 2451 11536 2485
rect 11570 2455 11652 2485
rect 11686 2455 11720 2489
rect 11754 2455 11788 2489
rect 11822 2455 11856 2489
rect 11890 2455 11924 2489
rect 11958 2455 11992 2489
rect 12026 2455 12060 2489
rect 12094 2455 12128 2489
rect 12162 2455 12196 2489
rect 12230 2455 12264 2489
rect 12298 2455 12332 2489
rect 12366 2455 12400 2489
rect 12434 2455 12468 2489
rect 12502 2482 13458 2489
rect 12502 2455 12573 2482
rect 11570 2451 12573 2455
rect 8643 2448 12573 2451
rect 12607 2448 12641 2482
rect 12675 2448 12709 2482
rect 12743 2448 12777 2482
rect 12811 2448 12845 2482
rect 12879 2448 12913 2482
rect 12947 2448 12981 2482
rect 13015 2448 13049 2482
rect 13083 2448 13117 2482
rect 13151 2448 13185 2482
rect 13219 2448 13253 2482
rect 13287 2448 13321 2482
rect 13355 2448 13458 2482
rect 8643 2419 13458 2448
rect 8643 2416 11652 2419
rect 8677 2382 8711 2416
rect 8745 2382 8779 2416
rect 8813 2382 8847 2416
rect 8881 2382 8915 2416
rect 8949 2382 8983 2416
rect 9017 2382 9051 2416
rect 9085 2382 9119 2416
rect 9153 2382 9187 2416
rect 9221 2382 9255 2416
rect 9289 2382 9323 2416
rect 9357 2382 9391 2416
rect 9425 2382 9459 2416
rect 9493 2382 9527 2416
rect 9561 2382 9595 2416
rect 9629 2382 9663 2416
rect 9697 2382 9731 2416
rect 9765 2382 9799 2416
rect 9833 2382 9867 2416
rect 9901 2382 9935 2416
rect 9969 2382 10003 2416
rect 10037 2382 10071 2416
rect 10105 2382 10139 2416
rect 10173 2382 10207 2416
rect 10241 2382 10312 2416
rect 10346 2382 10380 2416
rect 10414 2382 10448 2416
rect 10482 2382 10516 2416
rect 10550 2382 10584 2416
rect 10618 2382 10652 2416
rect 10686 2382 10720 2416
rect 10754 2382 10788 2416
rect 10822 2382 10856 2416
rect 10890 2382 10924 2416
rect 10958 2382 10992 2416
rect 11026 2382 11060 2416
rect 11094 2382 11128 2416
rect 11162 2382 11196 2416
rect 11230 2382 11264 2416
rect 11298 2382 11332 2416
rect 11366 2382 11400 2416
rect 11434 2382 11468 2416
rect 11502 2382 11536 2416
rect 11570 2385 11652 2416
rect 11686 2385 11720 2419
rect 11754 2385 11788 2419
rect 11822 2385 11856 2419
rect 11890 2385 11924 2419
rect 11958 2385 11992 2419
rect 12026 2385 12060 2419
rect 12094 2385 12128 2419
rect 12162 2385 12196 2419
rect 12230 2385 12264 2419
rect 12298 2385 12332 2419
rect 12366 2385 12400 2419
rect 12434 2385 12468 2419
rect 12502 2413 13458 2419
rect 12502 2385 12573 2413
rect 11570 2382 12573 2385
rect 8643 2379 12573 2382
rect 12607 2379 12641 2413
rect 12675 2379 12709 2413
rect 12743 2379 12777 2413
rect 12811 2379 12845 2413
rect 12879 2379 12913 2413
rect 12947 2379 12981 2413
rect 13015 2379 13049 2413
rect 13083 2379 13117 2413
rect 13151 2379 13185 2413
rect 13219 2379 13253 2413
rect 13287 2379 13321 2413
rect 13355 2379 13458 2413
rect 8643 2349 13458 2379
rect 8643 2347 11652 2349
rect 8677 2313 8711 2347
rect 8745 2313 8779 2347
rect 8813 2313 8847 2347
rect 8881 2313 8915 2347
rect 8949 2313 8983 2347
rect 9017 2313 9051 2347
rect 9085 2313 9119 2347
rect 9153 2313 9187 2347
rect 9221 2313 9255 2347
rect 9289 2313 9323 2347
rect 9357 2313 9391 2347
rect 9425 2313 9459 2347
rect 9493 2313 9527 2347
rect 9561 2313 9595 2347
rect 9629 2313 9663 2347
rect 9697 2313 9731 2347
rect 9765 2313 9799 2347
rect 9833 2313 9867 2347
rect 9901 2313 9935 2347
rect 9969 2313 10003 2347
rect 10037 2313 10071 2347
rect 10105 2313 10139 2347
rect 10173 2313 10207 2347
rect 10241 2313 10312 2347
rect 10346 2313 10380 2347
rect 10414 2313 10448 2347
rect 10482 2313 10516 2347
rect 10550 2313 10584 2347
rect 10618 2313 10652 2347
rect 10686 2313 10720 2347
rect 10754 2313 10788 2347
rect 10822 2313 10856 2347
rect 10890 2313 10924 2347
rect 10958 2313 10992 2347
rect 11026 2313 11060 2347
rect 11094 2313 11128 2347
rect 11162 2313 11196 2347
rect 11230 2313 11264 2347
rect 11298 2313 11332 2347
rect 11366 2313 11400 2347
rect 11434 2313 11468 2347
rect 11502 2313 11536 2347
rect 11570 2315 11652 2347
rect 11686 2315 11720 2349
rect 11754 2315 11788 2349
rect 11822 2315 11856 2349
rect 11890 2315 11924 2349
rect 11958 2315 11992 2349
rect 12026 2315 12060 2349
rect 12094 2315 12128 2349
rect 12162 2315 12196 2349
rect 12230 2315 12264 2349
rect 12298 2315 12332 2349
rect 12366 2315 12400 2349
rect 12434 2315 12468 2349
rect 12502 2344 13458 2349
rect 12502 2315 12573 2344
rect 11570 2313 12573 2315
rect 8643 2310 12573 2313
rect 12607 2310 12641 2344
rect 12675 2310 12709 2344
rect 12743 2310 12777 2344
rect 12811 2310 12845 2344
rect 12879 2310 12913 2344
rect 12947 2310 12981 2344
rect 13015 2310 13049 2344
rect 13083 2310 13117 2344
rect 13151 2310 13185 2344
rect 13219 2310 13253 2344
rect 13287 2310 13321 2344
rect 13355 2310 13458 2344
rect 8643 2279 13458 2310
rect 8643 2278 11652 2279
rect 8677 2244 8711 2278
rect 8745 2244 8779 2278
rect 8813 2244 8847 2278
rect 8881 2244 8915 2278
rect 8949 2244 8983 2278
rect 9017 2244 9051 2278
rect 9085 2244 9119 2278
rect 9153 2244 9187 2278
rect 9221 2244 9255 2278
rect 9289 2244 9323 2278
rect 9357 2244 9391 2278
rect 9425 2244 9459 2278
rect 9493 2244 9527 2278
rect 9561 2244 9595 2278
rect 9629 2244 9663 2278
rect 9697 2244 9731 2278
rect 9765 2244 9799 2278
rect 9833 2244 9867 2278
rect 9901 2244 9935 2278
rect 9969 2244 10003 2278
rect 10037 2244 10071 2278
rect 10105 2244 10139 2278
rect 10173 2244 10207 2278
rect 10241 2244 10312 2278
rect 10346 2244 10380 2278
rect 10414 2244 10448 2278
rect 10482 2244 10516 2278
rect 10550 2244 10584 2278
rect 10618 2244 10652 2278
rect 10686 2244 10720 2278
rect 10754 2244 10788 2278
rect 10822 2244 10856 2278
rect 10890 2244 10924 2278
rect 10958 2244 10992 2278
rect 11026 2244 11060 2278
rect 11094 2244 11128 2278
rect 11162 2244 11196 2278
rect 11230 2244 11264 2278
rect 11298 2244 11332 2278
rect 11366 2244 11400 2278
rect 11434 2244 11468 2278
rect 11502 2244 11536 2278
rect 11570 2245 11652 2278
rect 11686 2245 11720 2279
rect 11754 2245 11788 2279
rect 11822 2245 11856 2279
rect 11890 2245 11924 2279
rect 11958 2245 11992 2279
rect 12026 2245 12060 2279
rect 12094 2245 12128 2279
rect 12162 2245 12196 2279
rect 12230 2245 12264 2279
rect 12298 2245 12332 2279
rect 12366 2245 12400 2279
rect 12434 2245 12468 2279
rect 12502 2275 13458 2279
rect 12502 2245 12573 2275
rect 11570 2244 12573 2245
rect 8643 2241 12573 2244
rect 12607 2241 12641 2275
rect 12675 2241 12709 2275
rect 12743 2241 12777 2275
rect 12811 2241 12845 2275
rect 12879 2241 12913 2275
rect 12947 2241 12981 2275
rect 13015 2241 13049 2275
rect 13083 2241 13117 2275
rect 13151 2241 13185 2275
rect 13219 2241 13253 2275
rect 13287 2241 13321 2275
rect 13355 2241 13458 2275
rect 8643 2209 13458 2241
rect 8677 2175 8711 2209
rect 8745 2175 8779 2209
rect 8813 2175 8847 2209
rect 8881 2175 8915 2209
rect 8949 2175 8983 2209
rect 9017 2175 9051 2209
rect 9085 2175 9119 2209
rect 9153 2175 9187 2209
rect 9221 2175 9255 2209
rect 9289 2175 9323 2209
rect 9357 2175 9391 2209
rect 9425 2175 9459 2209
rect 9493 2175 9527 2209
rect 9561 2175 9595 2209
rect 9629 2175 9663 2209
rect 9697 2175 9731 2209
rect 9765 2175 9799 2209
rect 9833 2175 9867 2209
rect 9901 2175 9935 2209
rect 9969 2175 10003 2209
rect 10037 2175 10071 2209
rect 10105 2175 10139 2209
rect 10173 2175 10207 2209
rect 10241 2175 10312 2209
rect 10346 2175 10380 2209
rect 10414 2175 10448 2209
rect 10482 2175 10516 2209
rect 10550 2175 10584 2209
rect 10618 2175 10652 2209
rect 10686 2175 10720 2209
rect 10754 2175 10788 2209
rect 10822 2175 10856 2209
rect 10890 2175 10924 2209
rect 10958 2175 10992 2209
rect 11026 2175 11060 2209
rect 11094 2175 11128 2209
rect 11162 2175 11196 2209
rect 11230 2175 11264 2209
rect 11298 2175 11332 2209
rect 11366 2175 11400 2209
rect 11434 2175 11468 2209
rect 11502 2175 11536 2209
rect 11570 2175 11652 2209
rect 11686 2175 11720 2209
rect 11754 2175 11788 2209
rect 11822 2175 11856 2209
rect 11890 2175 11924 2209
rect 11958 2175 11992 2209
rect 12026 2175 12060 2209
rect 12094 2175 12128 2209
rect 12162 2175 12196 2209
rect 12230 2175 12264 2209
rect 12298 2175 12332 2209
rect 12366 2175 12400 2209
rect 12434 2175 12468 2209
rect 12502 2206 13458 2209
rect 12502 2175 12573 2206
rect 8643 2172 12573 2175
rect 12607 2172 12641 2206
rect 12675 2172 12709 2206
rect 12743 2172 12777 2206
rect 12811 2172 12845 2206
rect 12879 2172 12913 2206
rect 12947 2172 12981 2206
rect 13015 2172 13049 2206
rect 13083 2172 13117 2206
rect 13151 2172 13185 2206
rect 13219 2172 13253 2206
rect 13287 2172 13321 2206
rect 13355 2172 13458 2206
rect 8643 2154 13458 2172
rect 8643 2140 11319 2154
rect 11713 2140 11752 2154
rect 11786 2140 11825 2154
rect 11859 2140 11898 2154
rect 11932 2140 11971 2154
rect 12005 2140 12044 2154
rect 12078 2140 12117 2154
rect 12151 2140 12190 2154
rect 12224 2140 12263 2154
rect 12297 2140 12336 2154
rect 12370 2140 12409 2154
rect 12443 2140 12482 2154
rect 8677 2106 8711 2140
rect 8745 2106 8779 2140
rect 8813 2106 8847 2140
rect 8881 2106 8915 2140
rect 8949 2106 8983 2140
rect 9017 2106 9051 2140
rect 9085 2106 9119 2140
rect 9153 2106 9187 2140
rect 9221 2106 9255 2140
rect 9289 2106 9323 2140
rect 9357 2106 9391 2140
rect 9425 2106 9459 2140
rect 9493 2106 9527 2140
rect 9561 2106 9595 2140
rect 9629 2106 9663 2140
rect 9697 2106 9731 2140
rect 9765 2106 9799 2140
rect 9833 2106 9867 2140
rect 9901 2106 9935 2140
rect 9969 2106 10003 2140
rect 10037 2106 10071 2140
rect 10105 2106 10139 2140
rect 10173 2106 10207 2140
rect 10241 2106 10312 2140
rect 10346 2106 10380 2140
rect 10414 2106 10448 2140
rect 10482 2106 10516 2140
rect 10550 2106 10584 2140
rect 10618 2106 10652 2140
rect 10686 2106 10720 2140
rect 10754 2106 10788 2140
rect 10822 2106 10856 2140
rect 10890 2106 10924 2140
rect 10958 2106 10992 2140
rect 11026 2106 11060 2140
rect 11094 2106 11128 2140
rect 11162 2106 11196 2140
rect 11230 2106 11264 2140
rect 11298 2106 11319 2140
rect 11713 2106 11720 2140
rect 11786 2120 11788 2140
rect 11754 2106 11788 2120
rect 11822 2120 11825 2140
rect 11890 2120 11898 2140
rect 11958 2120 11971 2140
rect 12026 2120 12044 2140
rect 12094 2120 12117 2140
rect 12162 2120 12190 2140
rect 12230 2120 12263 2140
rect 11822 2106 11856 2120
rect 11890 2106 11924 2120
rect 11958 2106 11992 2120
rect 12026 2106 12060 2120
rect 12094 2106 12128 2120
rect 12162 2106 12196 2120
rect 12230 2106 12264 2120
rect 12298 2106 12332 2140
rect 12370 2120 12400 2140
rect 12443 2120 12468 2140
rect 12516 2120 12555 2154
rect 12589 2137 12628 2154
rect 12662 2137 12701 2154
rect 12735 2137 12774 2154
rect 12808 2137 12847 2154
rect 12881 2137 12920 2154
rect 12954 2137 12993 2154
rect 13027 2137 13066 2154
rect 13100 2137 13139 2154
rect 13173 2137 13212 2154
rect 13246 2137 13458 2154
rect 12607 2120 12628 2137
rect 12675 2120 12701 2137
rect 12743 2120 12774 2137
rect 12366 2106 12400 2120
rect 12434 2106 12468 2120
rect 12502 2106 12573 2120
rect 8643 2071 11319 2106
rect 11713 2103 12573 2106
rect 12607 2103 12641 2120
rect 12675 2103 12709 2120
rect 12743 2103 12777 2120
rect 12811 2103 12845 2137
rect 12881 2120 12913 2137
rect 12954 2120 12981 2137
rect 13027 2120 13049 2137
rect 13100 2120 13117 2137
rect 13173 2120 13185 2137
rect 13246 2120 13253 2137
rect 12879 2103 12913 2120
rect 12947 2103 12981 2120
rect 13015 2103 13049 2120
rect 13083 2103 13117 2120
rect 13151 2103 13185 2120
rect 13219 2103 13253 2120
rect 13287 2103 13321 2137
rect 13355 2103 13458 2137
rect 11713 2082 13458 2103
rect 11713 2071 11752 2082
rect 11786 2071 11825 2082
rect 11859 2071 11898 2082
rect 11932 2071 11971 2082
rect 12005 2071 12044 2082
rect 12078 2071 12117 2082
rect 12151 2071 12190 2082
rect 12224 2071 12263 2082
rect 12297 2071 12336 2082
rect 12370 2071 12409 2082
rect 12443 2071 12482 2082
rect 8677 2037 8711 2071
rect 8745 2037 8779 2071
rect 8813 2037 8847 2071
rect 8881 2037 8915 2071
rect 8949 2037 8983 2071
rect 9017 2037 9051 2071
rect 9085 2037 9119 2071
rect 9153 2037 9187 2071
rect 9221 2037 9255 2071
rect 9289 2037 9323 2071
rect 9357 2037 9391 2071
rect 9425 2037 9459 2071
rect 9493 2037 9527 2071
rect 9561 2037 9595 2071
rect 9629 2037 9663 2071
rect 9697 2037 9731 2071
rect 9765 2037 9799 2071
rect 9833 2037 9867 2071
rect 9901 2037 9935 2071
rect 9969 2037 10003 2071
rect 10037 2037 10071 2071
rect 10105 2037 10139 2071
rect 10173 2037 10207 2071
rect 10241 2037 10312 2071
rect 10346 2037 10380 2071
rect 10414 2037 10448 2071
rect 10482 2037 10516 2071
rect 10550 2037 10584 2071
rect 10618 2037 10652 2071
rect 10686 2037 10720 2071
rect 10754 2037 10788 2071
rect 10822 2037 10856 2071
rect 10890 2037 10924 2071
rect 10958 2037 10992 2071
rect 11026 2037 11060 2071
rect 11094 2037 11128 2071
rect 11162 2037 11196 2071
rect 11230 2037 11264 2071
rect 11298 2037 11319 2071
rect 11713 2037 11720 2071
rect 11786 2048 11788 2071
rect 11754 2037 11788 2048
rect 11822 2048 11825 2071
rect 11890 2048 11898 2071
rect 11958 2048 11971 2071
rect 12026 2048 12044 2071
rect 12094 2048 12117 2071
rect 12162 2048 12190 2071
rect 12230 2048 12263 2071
rect 11822 2037 11856 2048
rect 11890 2037 11924 2048
rect 11958 2037 11992 2048
rect 12026 2037 12060 2048
rect 12094 2037 12128 2048
rect 12162 2037 12196 2048
rect 12230 2037 12264 2048
rect 12298 2037 12332 2071
rect 12370 2048 12400 2071
rect 12443 2048 12468 2071
rect 12516 2048 12555 2082
rect 12589 2068 12628 2082
rect 12662 2068 12701 2082
rect 12735 2068 12774 2082
rect 12808 2068 12847 2082
rect 12881 2068 12920 2082
rect 12954 2068 12993 2082
rect 13027 2068 13066 2082
rect 13100 2068 13139 2082
rect 13173 2068 13212 2082
rect 13246 2068 13458 2082
rect 23568 2712 23597 2752
rect 23767 2712 23796 2752
rect 23568 2678 23593 2712
rect 23771 2678 23796 2712
rect 23568 2638 23597 2678
rect 23767 2638 23796 2678
rect 23568 2604 23593 2638
rect 23771 2604 23796 2638
rect 23568 2564 23597 2604
rect 23767 2564 23796 2604
rect 23568 2530 23593 2564
rect 23771 2530 23796 2564
rect 23568 2490 23597 2530
rect 23767 2490 23796 2530
rect 23568 2456 23593 2490
rect 23771 2456 23796 2490
rect 23568 2416 23597 2456
rect 23767 2416 23796 2456
rect 23568 2382 23593 2416
rect 23771 2382 23796 2416
rect 23568 2342 23597 2382
rect 23767 2342 23796 2382
rect 23568 2308 23593 2342
rect 23771 2308 23796 2342
rect 23568 2268 23597 2308
rect 23767 2268 23796 2308
rect 23568 2234 23593 2268
rect 23771 2234 23796 2268
rect 23568 2194 23597 2234
rect 23767 2194 23796 2234
rect 23568 2160 23593 2194
rect 23771 2160 23796 2194
rect 23568 2120 23597 2160
rect 23767 2120 23796 2160
rect 23568 2086 23593 2120
rect 23627 2086 23665 2110
rect 23699 2086 23737 2110
rect 23771 2086 23796 2120
rect 23568 2076 23796 2086
rect 12607 2048 12628 2068
rect 12675 2048 12701 2068
rect 12743 2048 12774 2068
rect 12366 2037 12400 2048
rect 12434 2037 12468 2048
rect 12502 2037 12573 2048
rect 4998 1798 5104 2032
rect 8643 2002 11319 2037
rect 11713 2034 12573 2037
rect 12607 2034 12641 2048
rect 12675 2034 12709 2048
rect 12743 2034 12777 2048
rect 12811 2034 12845 2068
rect 12881 2048 12913 2068
rect 12954 2048 12981 2068
rect 13027 2048 13049 2068
rect 13100 2048 13117 2068
rect 13173 2048 13185 2068
rect 13246 2048 13253 2068
rect 12879 2034 12913 2048
rect 12947 2034 12981 2048
rect 13015 2034 13049 2048
rect 13083 2034 13117 2048
rect 13151 2034 13185 2048
rect 13219 2034 13253 2048
rect 13287 2034 13321 2068
rect 13355 2034 13458 2068
rect 11713 2010 13458 2034
rect 11713 2002 11752 2010
rect 11786 2002 11825 2010
rect 11859 2002 11898 2010
rect 11932 2002 11971 2010
rect 12005 2002 12044 2010
rect 12078 2002 12117 2010
rect 12151 2002 12190 2010
rect 12224 2002 12263 2010
rect 12297 2002 12336 2010
rect 12370 2002 12409 2010
rect 12443 2002 12482 2010
rect 8677 1968 8711 2002
rect 8745 1975 8779 2002
rect 8745 1968 8774 1975
rect 8813 1968 8847 2002
rect 8881 1968 8915 2002
rect 8949 1975 8983 2002
rect 9017 1975 9051 2002
rect 9085 1975 9119 2002
rect 9153 1975 9187 2002
rect 9221 1975 9255 2002
rect 9289 1975 9323 2002
rect 8954 1968 8983 1975
rect 9027 1968 9051 1975
rect 9100 1968 9119 1975
rect 9173 1968 9187 1975
rect 9246 1968 9255 1975
rect 9319 1968 9323 1975
rect 9357 1975 9391 2002
rect 9425 1975 9459 2002
rect 9493 1975 9527 2002
rect 9561 1975 9595 2002
rect 9629 1975 9663 2002
rect 9697 1975 9731 2002
rect 9765 1975 9799 2002
rect 9357 1968 9358 1975
rect 9425 1968 9431 1975
rect 9493 1968 9504 1975
rect 9561 1968 9577 1975
rect 9629 1968 9650 1975
rect 9697 1968 9723 1975
rect 9765 1968 9796 1975
rect 9833 1968 9867 2002
rect 9901 1975 9935 2002
rect 9969 1975 10003 2002
rect 10037 1975 10071 2002
rect 10105 1975 10139 2002
rect 10173 1975 10207 2002
rect 10241 1975 10312 2002
rect 9903 1968 9935 1975
rect 9976 1968 10003 1975
rect 10049 1968 10071 1975
rect 10122 1968 10139 1975
rect 10195 1968 10207 1975
rect 8643 1941 8774 1968
rect 8808 1941 8847 1968
rect 8881 1941 8920 1968
rect 8954 1941 8993 1968
rect 9027 1941 9066 1968
rect 9100 1941 9139 1968
rect 9173 1941 9212 1968
rect 9246 1941 9285 1968
rect 9319 1941 9358 1968
rect 9392 1941 9431 1968
rect 9465 1941 9504 1968
rect 9538 1941 9577 1968
rect 9611 1941 9650 1968
rect 9684 1941 9723 1968
rect 9757 1941 9796 1968
rect 9830 1941 9869 1968
rect 9903 1941 9942 1968
rect 9976 1941 10015 1968
rect 10049 1941 10088 1968
rect 10122 1941 10161 1968
rect 10195 1941 10234 1968
rect 10268 1941 10307 1975
rect 10346 1968 10380 2002
rect 10414 1968 10448 2002
rect 10482 1975 10516 2002
rect 10550 1975 10584 2002
rect 10618 1975 10652 2002
rect 10686 1975 10720 2002
rect 10754 1975 10788 2002
rect 10822 1975 10856 2002
rect 10890 1975 10924 2002
rect 10958 1975 10992 2002
rect 11026 1975 11060 2002
rect 11094 1975 11128 2002
rect 11162 1975 11196 2002
rect 11230 1975 11264 2002
rect 11298 1975 11319 2002
rect 10487 1968 10516 1975
rect 10560 1968 10584 1975
rect 11713 1968 11720 2002
rect 11786 1976 11788 2002
rect 11754 1968 11788 1976
rect 11822 1976 11825 2002
rect 11890 1976 11898 2002
rect 11958 1976 11971 2002
rect 12026 1976 12044 2002
rect 12094 1976 12117 2002
rect 12162 1976 12190 2002
rect 12230 1976 12263 2002
rect 11822 1968 11856 1976
rect 11890 1968 11924 1976
rect 11958 1968 11992 1976
rect 12026 1968 12060 1976
rect 12094 1968 12128 1976
rect 12162 1968 12196 1976
rect 12230 1968 12264 1976
rect 12298 1968 12332 2002
rect 12370 1976 12400 2002
rect 12443 1976 12468 2002
rect 12516 1976 12555 2010
rect 12589 1999 12628 2010
rect 12662 1999 12701 2010
rect 12735 1999 12774 2010
rect 12808 1999 12847 2010
rect 12881 1999 12920 2010
rect 12954 1999 12993 2010
rect 13027 1999 13066 2010
rect 13100 1999 13139 2010
rect 13173 1999 13212 2010
rect 13246 1999 13458 2010
rect 12607 1976 12628 1999
rect 12675 1976 12701 1999
rect 12743 1976 12774 1999
rect 12366 1968 12400 1976
rect 12434 1968 12468 1976
rect 12502 1968 12573 1976
rect 10341 1941 10380 1968
rect 10414 1941 10453 1968
rect 10487 1941 10526 1968
rect 10560 1941 10599 1968
rect 8643 1933 10599 1941
rect 11713 1965 12573 1968
rect 12607 1965 12641 1976
rect 12675 1965 12709 1976
rect 12743 1965 12777 1976
rect 12811 1965 12845 1999
rect 12881 1976 12913 1999
rect 12954 1976 12981 1999
rect 13027 1976 13049 1999
rect 13100 1976 13117 1999
rect 13173 1976 13185 1999
rect 13246 1976 13253 1999
rect 12879 1965 12913 1976
rect 12947 1965 12981 1976
rect 13015 1965 13049 1976
rect 13083 1965 13117 1976
rect 13151 1965 13185 1976
rect 13219 1965 13253 1976
rect 13287 1965 13321 1999
rect 13355 1965 13458 1999
rect 11713 1938 13458 1965
rect 11713 1933 11752 1938
rect 11786 1933 11825 1938
rect 11859 1933 11898 1938
rect 11932 1933 11971 1938
rect 12005 1933 12044 1938
rect 12078 1933 12117 1938
rect 12151 1933 12190 1938
rect 12224 1933 12263 1938
rect 12297 1933 12336 1938
rect 12370 1933 12409 1938
rect 12443 1933 12482 1938
rect 8677 1899 8711 1933
rect 8745 1903 8779 1933
rect 8745 1899 8774 1903
rect 8813 1899 8847 1933
rect 8881 1899 8915 1933
rect 8949 1903 8983 1933
rect 9017 1903 9051 1933
rect 9085 1903 9119 1933
rect 9153 1903 9187 1933
rect 9221 1903 9255 1933
rect 9289 1903 9323 1933
rect 8954 1899 8983 1903
rect 9027 1899 9051 1903
rect 9100 1899 9119 1903
rect 9173 1899 9187 1903
rect 9246 1899 9255 1903
rect 9319 1899 9323 1903
rect 9357 1903 9391 1933
rect 9425 1903 9459 1933
rect 9493 1903 9527 1933
rect 9561 1903 9595 1933
rect 9629 1903 9663 1933
rect 9697 1903 9731 1933
rect 9765 1903 9799 1933
rect 9357 1899 9358 1903
rect 9425 1899 9431 1903
rect 9493 1899 9504 1903
rect 9561 1899 9577 1903
rect 9629 1899 9650 1903
rect 9697 1899 9723 1903
rect 9765 1899 9796 1903
rect 9833 1899 9867 1933
rect 9901 1903 9935 1933
rect 9969 1903 10003 1933
rect 10037 1903 10071 1933
rect 10105 1903 10139 1933
rect 10173 1903 10207 1933
rect 10241 1903 10312 1933
rect 9903 1899 9935 1903
rect 9976 1899 10003 1903
rect 10049 1899 10071 1903
rect 10122 1899 10139 1903
rect 10195 1899 10207 1903
rect 8643 1869 8774 1899
rect 8808 1869 8847 1899
rect 8881 1869 8920 1899
rect 8954 1869 8993 1899
rect 9027 1869 9066 1899
rect 9100 1869 9139 1899
rect 9173 1869 9212 1899
rect 9246 1869 9285 1899
rect 9319 1869 9358 1899
rect 9392 1869 9431 1899
rect 9465 1869 9504 1899
rect 9538 1869 9577 1899
rect 9611 1869 9650 1899
rect 9684 1869 9723 1899
rect 9757 1869 9796 1899
rect 9830 1869 9869 1899
rect 9903 1869 9942 1899
rect 9976 1869 10015 1899
rect 10049 1869 10088 1899
rect 10122 1869 10161 1899
rect 10195 1869 10234 1899
rect 10268 1869 10307 1903
rect 10346 1899 10380 1933
rect 10414 1899 10448 1933
rect 10482 1903 10516 1933
rect 10550 1903 10584 1933
rect 10487 1899 10516 1903
rect 10560 1899 10584 1903
rect 11713 1899 11720 1933
rect 11786 1904 11788 1933
rect 11754 1899 11788 1904
rect 11822 1904 11825 1933
rect 11890 1904 11898 1933
rect 11958 1904 11971 1933
rect 12026 1904 12044 1933
rect 12094 1904 12117 1933
rect 12162 1904 12190 1933
rect 12230 1904 12263 1933
rect 11822 1899 11856 1904
rect 11890 1899 11924 1904
rect 11958 1899 11992 1904
rect 12026 1899 12060 1904
rect 12094 1899 12128 1904
rect 12162 1899 12196 1904
rect 12230 1899 12264 1904
rect 12298 1899 12332 1933
rect 12370 1904 12400 1933
rect 12443 1904 12468 1933
rect 12516 1904 12555 1938
rect 12589 1930 12628 1938
rect 12662 1930 12701 1938
rect 12735 1930 12774 1938
rect 12808 1930 12847 1938
rect 12881 1930 12920 1938
rect 12954 1930 12993 1938
rect 13027 1930 13066 1938
rect 13100 1930 13139 1938
rect 13173 1930 13212 1938
rect 13246 1930 13458 1938
rect 12607 1904 12628 1930
rect 12675 1904 12701 1930
rect 12743 1904 12774 1930
rect 12366 1899 12400 1904
rect 12434 1899 12468 1904
rect 12502 1899 12573 1904
rect 10341 1869 10380 1899
rect 10414 1869 10453 1899
rect 10487 1869 10526 1899
rect 10560 1869 10599 1899
rect 11713 1896 12573 1899
rect 12607 1896 12641 1904
rect 12675 1896 12709 1904
rect 12743 1896 12777 1904
rect 12811 1896 12845 1930
rect 12881 1904 12913 1930
rect 12954 1904 12981 1930
rect 13027 1904 13049 1930
rect 13100 1904 13117 1930
rect 13173 1904 13185 1930
rect 13246 1904 13253 1930
rect 12879 1896 12913 1904
rect 12947 1896 12981 1904
rect 13015 1896 13049 1904
rect 13083 1896 13117 1904
rect 13151 1896 13185 1904
rect 13219 1896 13253 1904
rect 13287 1896 13321 1930
rect 13355 1896 13458 1930
rect 8643 1864 11319 1869
rect 11713 1866 13458 1896
rect 11713 1864 11752 1866
rect 11786 1864 11825 1866
rect 11859 1864 11898 1866
rect 11932 1864 11971 1866
rect 12005 1864 12044 1866
rect 12078 1864 12117 1866
rect 12151 1864 12190 1866
rect 12224 1864 12263 1866
rect 12297 1864 12336 1866
rect 12370 1864 12409 1866
rect 12443 1864 12482 1866
rect 8677 1830 8711 1864
rect 8745 1830 8779 1864
rect 8813 1830 8847 1864
rect 8881 1830 8915 1864
rect 8949 1830 8983 1864
rect 9017 1830 9051 1864
rect 9085 1830 9119 1864
rect 9153 1830 9187 1864
rect 9221 1830 9255 1864
rect 9289 1830 9323 1864
rect 9357 1830 9391 1864
rect 9425 1830 9459 1864
rect 9493 1830 9527 1864
rect 9561 1830 9595 1864
rect 9629 1830 9663 1864
rect 9697 1830 9731 1864
rect 9765 1830 9799 1864
rect 9833 1830 9867 1864
rect 9901 1830 9935 1864
rect 9969 1830 10003 1864
rect 10037 1830 10071 1864
rect 10105 1830 10139 1864
rect 10173 1830 10207 1864
rect 10241 1830 10312 1864
rect 10346 1830 10380 1864
rect 10414 1830 10448 1864
rect 10482 1830 10516 1864
rect 10550 1830 10584 1864
rect 10618 1830 10652 1864
rect 10686 1830 10720 1864
rect 10754 1830 10788 1864
rect 10822 1830 10856 1864
rect 10890 1830 10924 1864
rect 10958 1830 10992 1864
rect 11026 1830 11060 1864
rect 11094 1830 11128 1864
rect 11162 1830 11196 1864
rect 11230 1830 11264 1864
rect 11298 1830 11319 1864
rect 11713 1830 11720 1864
rect 11786 1832 11788 1864
rect 11754 1830 11788 1832
rect 11822 1832 11825 1864
rect 11890 1832 11898 1864
rect 11958 1832 11971 1864
rect 12026 1832 12044 1864
rect 12094 1832 12117 1864
rect 12162 1832 12190 1864
rect 12230 1832 12263 1864
rect 11822 1830 11856 1832
rect 11890 1830 11924 1832
rect 11958 1830 11992 1832
rect 12026 1830 12060 1832
rect 12094 1830 12128 1832
rect 12162 1830 12196 1832
rect 12230 1830 12264 1832
rect 12298 1830 12332 1864
rect 12370 1832 12400 1864
rect 12443 1832 12468 1864
rect 12516 1832 12555 1866
rect 12589 1861 12628 1866
rect 12662 1861 12701 1866
rect 12735 1861 12774 1866
rect 12808 1861 12847 1866
rect 12881 1861 12920 1866
rect 12954 1861 12993 1866
rect 13027 1861 13066 1866
rect 13100 1861 13139 1866
rect 13173 1861 13212 1866
rect 13246 1861 13458 1866
rect 12366 1830 12400 1832
rect 12434 1830 12468 1832
rect 12502 1830 12573 1832
rect 1460 1793 1575 1796
rect 1460 1772 1507 1793
rect 1541 1772 1575 1793
rect 1609 1772 1643 1796
rect 1491 1759 1507 1772
rect 1563 1762 1575 1772
rect 1635 1762 1643 1772
rect 1491 1738 1529 1759
rect 1563 1738 1601 1762
rect 1635 1738 1677 1762
rect 1460 1727 1677 1738
rect 1460 1725 1575 1727
rect 1460 1699 1507 1725
rect 1541 1699 1575 1725
rect 1609 1699 1643 1727
rect 1491 1691 1507 1699
rect 1563 1693 1575 1699
rect 1635 1693 1643 1699
rect 1491 1665 1529 1691
rect 1563 1665 1601 1693
rect 1635 1665 1677 1693
rect 1460 1658 1677 1665
rect 1460 1657 1575 1658
rect 1460 1626 1507 1657
rect 1541 1626 1575 1657
rect 1609 1626 1643 1658
rect 1491 1623 1507 1626
rect 1563 1624 1575 1626
rect 1635 1624 1643 1626
rect 1491 1592 1529 1623
rect 1563 1592 1601 1624
rect 1635 1592 1677 1624
rect 1460 1589 1677 1592
rect 8643 1795 11319 1830
rect 11713 1795 12573 1830
rect 8677 1761 8711 1795
rect 8745 1761 8779 1795
rect 8813 1761 8847 1795
rect 8881 1761 8915 1795
rect 8949 1761 8983 1795
rect 9017 1761 9051 1795
rect 9085 1761 9119 1795
rect 9153 1761 9187 1795
rect 9221 1761 9255 1795
rect 9289 1761 9323 1795
rect 9357 1761 9391 1795
rect 9425 1761 9459 1795
rect 9493 1761 9527 1795
rect 9561 1761 9595 1795
rect 9629 1761 9663 1795
rect 9697 1761 9731 1795
rect 9765 1761 9799 1795
rect 9833 1761 9867 1795
rect 9901 1761 9935 1795
rect 9969 1761 10003 1795
rect 10037 1761 10071 1795
rect 10105 1761 10139 1795
rect 10173 1761 10207 1795
rect 10241 1761 10312 1795
rect 10346 1761 10380 1795
rect 10414 1761 10448 1795
rect 10482 1761 10516 1795
rect 10550 1761 10584 1795
rect 10618 1761 10652 1795
rect 10686 1761 10720 1795
rect 10754 1761 10788 1795
rect 10822 1761 10856 1795
rect 10890 1761 10924 1795
rect 10958 1761 10992 1795
rect 11026 1761 11060 1795
rect 11094 1761 11128 1795
rect 11162 1761 11196 1795
rect 11230 1761 11264 1795
rect 11298 1761 11319 1795
rect 11713 1761 11720 1795
rect 11754 1794 11788 1795
rect 11786 1761 11788 1794
rect 11822 1794 11856 1795
rect 11890 1794 11924 1795
rect 11958 1794 11992 1795
rect 12026 1794 12060 1795
rect 12094 1794 12128 1795
rect 12162 1794 12196 1795
rect 12230 1794 12264 1795
rect 11822 1761 11825 1794
rect 11890 1761 11898 1794
rect 11958 1761 11971 1794
rect 12026 1761 12044 1794
rect 12094 1761 12117 1794
rect 12162 1761 12190 1794
rect 12230 1761 12263 1794
rect 12298 1761 12332 1795
rect 12366 1794 12400 1795
rect 12434 1794 12468 1795
rect 12502 1794 12573 1795
rect 12370 1761 12400 1794
rect 12443 1761 12468 1794
rect 8643 1760 11319 1761
rect 11713 1760 11752 1761
rect 11786 1760 11825 1761
rect 11859 1760 11898 1761
rect 11932 1760 11971 1761
rect 12005 1760 12044 1761
rect 12078 1760 12117 1761
rect 12151 1760 12190 1761
rect 12224 1760 12263 1761
rect 12297 1760 12336 1761
rect 12370 1760 12409 1761
rect 12443 1760 12482 1761
rect 12516 1760 12555 1794
rect 8643 1726 12573 1760
rect 8677 1692 8711 1726
rect 8745 1692 8779 1726
rect 8813 1692 8847 1726
rect 8881 1692 8915 1726
rect 8949 1692 8983 1726
rect 9017 1692 9051 1726
rect 9085 1692 9119 1726
rect 9153 1692 9187 1726
rect 9221 1692 9255 1726
rect 9289 1692 9323 1726
rect 9357 1692 9391 1726
rect 9425 1692 9459 1726
rect 9493 1692 9527 1726
rect 9561 1692 9595 1726
rect 9629 1692 9663 1726
rect 9697 1692 9731 1726
rect 9765 1692 9799 1726
rect 9833 1692 9867 1726
rect 9901 1692 9935 1726
rect 9969 1692 10003 1726
rect 10037 1692 10071 1726
rect 10105 1692 10139 1726
rect 10173 1692 10207 1726
rect 10241 1692 10312 1726
rect 10346 1692 10380 1726
rect 10414 1692 10448 1726
rect 10482 1692 10516 1726
rect 10550 1692 10584 1726
rect 10618 1692 10652 1726
rect 10686 1692 10720 1726
rect 10754 1692 10788 1726
rect 10822 1692 10856 1726
rect 10890 1692 10924 1726
rect 10958 1692 10992 1726
rect 11026 1692 11060 1726
rect 11094 1692 11128 1726
rect 11162 1692 11196 1726
rect 11230 1692 11264 1726
rect 11298 1692 11332 1726
rect 11366 1692 11400 1726
rect 11434 1692 11468 1726
rect 11502 1692 11536 1726
rect 11570 1692 11652 1726
rect 11686 1692 11720 1726
rect 11754 1692 11788 1726
rect 11822 1692 11856 1726
rect 11890 1692 11924 1726
rect 11958 1692 11992 1726
rect 12026 1692 12060 1726
rect 12094 1692 12128 1726
rect 12162 1692 12196 1726
rect 12230 1692 12264 1726
rect 12298 1692 12332 1726
rect 12366 1692 12400 1726
rect 12434 1692 12468 1726
rect 12502 1692 12573 1726
rect 8643 1657 12573 1692
rect 8677 1623 8711 1657
rect 8745 1623 8779 1657
rect 8813 1623 8847 1657
rect 8881 1623 8915 1657
rect 8949 1623 8983 1657
rect 9017 1623 9051 1657
rect 9085 1623 9119 1657
rect 9153 1623 9187 1657
rect 9221 1623 9255 1657
rect 9289 1623 9323 1657
rect 9357 1623 9391 1657
rect 9425 1623 9459 1657
rect 9493 1623 9527 1657
rect 9561 1623 9595 1657
rect 9629 1623 9663 1657
rect 9697 1623 9731 1657
rect 9765 1623 9799 1657
rect 9833 1623 9867 1657
rect 9901 1623 9935 1657
rect 9969 1623 10003 1657
rect 10037 1623 10071 1657
rect 10105 1623 10139 1657
rect 10173 1623 10207 1657
rect 10241 1623 10312 1657
rect 10346 1623 10380 1657
rect 10414 1623 10448 1657
rect 10482 1623 10516 1657
rect 10550 1623 10584 1657
rect 10618 1623 10652 1657
rect 10686 1623 10720 1657
rect 10754 1623 10788 1657
rect 10822 1623 10856 1657
rect 10890 1623 10924 1657
rect 10958 1623 10992 1657
rect 11026 1623 11060 1657
rect 11094 1623 11128 1657
rect 11162 1623 11196 1657
rect 11230 1623 11264 1657
rect 11298 1623 11332 1657
rect 11366 1623 11400 1657
rect 11434 1623 11468 1657
rect 11502 1623 11536 1657
rect 11570 1623 11652 1657
rect 11686 1623 11720 1657
rect 11754 1623 11788 1657
rect 11822 1623 11856 1657
rect 11890 1623 11924 1657
rect 11958 1623 11992 1657
rect 12026 1623 12060 1657
rect 12094 1623 12128 1657
rect 12162 1623 12196 1657
rect 12230 1623 12264 1657
rect 12298 1623 12332 1657
rect 12366 1623 12400 1657
rect 12434 1623 12468 1657
rect 12502 1623 12573 1657
rect 13355 1623 13458 1861
rect 8643 1589 13458 1623
rect 1460 1555 1507 1589
rect 1541 1555 1575 1589
rect 1609 1555 1643 1589
rect 1460 1553 1677 1555
rect 1491 1519 1529 1553
rect 1563 1521 1601 1553
rect 1635 1521 1677 1553
rect 8388 1555 8412 1589
rect 8446 1557 8482 1589
rect 8516 1557 8552 1589
rect 8586 1557 8622 1589
rect 8468 1555 8482 1557
rect 8543 1555 8552 1557
rect 8618 1555 8622 1557
rect 8656 1557 8692 1589
rect 8726 1557 8762 1589
rect 8796 1557 8832 1589
rect 8866 1557 8902 1589
rect 8936 1557 8972 1589
rect 9006 1557 9043 1589
rect 9077 1557 9114 1589
rect 9148 1557 9185 1589
rect 8656 1555 8659 1557
rect 8726 1555 8734 1557
rect 8796 1555 8809 1557
rect 8866 1555 8884 1557
rect 8936 1555 8959 1557
rect 9006 1555 9034 1557
rect 9077 1555 9109 1557
rect 9148 1555 9184 1557
rect 9219 1555 9256 1589
rect 9290 1557 9327 1589
rect 9361 1557 9398 1589
rect 9432 1557 9469 1589
rect 9503 1557 9540 1589
rect 9574 1557 9611 1589
rect 9645 1557 9682 1589
rect 9716 1557 9753 1589
rect 9787 1557 9824 1589
rect 9293 1555 9327 1557
rect 9368 1555 9398 1557
rect 9443 1555 9469 1557
rect 9518 1555 9540 1557
rect 9593 1555 9611 1557
rect 9668 1555 9682 1557
rect 9743 1555 9753 1557
rect 9818 1555 9824 1557
rect 9858 1557 9895 1589
rect 9858 1555 9860 1557
rect 8388 1523 8434 1555
rect 8468 1523 8509 1555
rect 8543 1523 8584 1555
rect 8618 1523 8659 1555
rect 8693 1523 8734 1555
rect 8768 1523 8809 1555
rect 8843 1523 8884 1555
rect 8918 1523 8959 1555
rect 8993 1523 9034 1555
rect 9068 1523 9109 1555
rect 9143 1523 9184 1555
rect 9218 1523 9259 1555
rect 9293 1523 9334 1555
rect 9368 1523 9409 1555
rect 9443 1523 9484 1555
rect 9518 1523 9559 1555
rect 9593 1523 9634 1555
rect 9668 1523 9709 1555
rect 9743 1523 9784 1555
rect 9818 1523 9860 1555
rect 9894 1555 9895 1557
rect 9929 1557 9966 1589
rect 10000 1583 13458 1589
rect 13728 2052 14489 2076
rect 13728 2018 13751 2052
rect 13785 2018 13819 2052
rect 13853 2018 13887 2052
rect 13921 2018 13955 2052
rect 13989 2018 14023 2052
rect 14057 2018 14091 2052
rect 14125 2018 14159 2052
rect 14193 2018 14227 2052
rect 14261 2018 14295 2052
rect 14329 2018 14363 2052
rect 14397 2042 14489 2052
rect 14523 2042 14567 2076
rect 14601 2061 23796 2076
rect 14601 2042 14701 2061
rect 14397 2018 14701 2042
rect 13728 2008 14701 2018
rect 13728 1980 14545 2008
rect 13728 1946 13751 1980
rect 13785 1946 13819 1980
rect 13853 1946 13887 1980
rect 13921 1946 13955 1980
rect 13989 1946 14023 1980
rect 14057 1946 14091 1980
rect 14125 1946 14159 1980
rect 14193 1946 14227 1980
rect 14261 1946 14295 1980
rect 14329 1946 14363 1980
rect 14397 1974 14545 1980
rect 14579 1974 14701 2008
rect 14397 1968 14701 1974
rect 14397 1946 14455 1968
rect 13728 1934 14455 1946
rect 14489 1939 14701 1968
rect 14489 1934 14523 1939
rect 13728 1908 14523 1934
rect 13728 1874 13751 1908
rect 13785 1874 13819 1908
rect 13853 1874 13887 1908
rect 13921 1874 13955 1908
rect 13989 1874 14023 1908
rect 14057 1874 14091 1908
rect 14125 1874 14159 1908
rect 14193 1874 14227 1908
rect 14261 1874 14295 1908
rect 14329 1874 14363 1908
rect 14397 1905 14523 1908
rect 14557 1916 14701 1939
rect 14557 1905 14591 1916
rect 14397 1897 14591 1905
rect 14397 1874 14455 1897
rect 13728 1863 14455 1874
rect 14489 1882 14591 1897
rect 14625 1882 14701 1916
rect 14489 1870 14701 1882
rect 14489 1863 14523 1870
rect 13728 1836 14523 1863
rect 14557 1846 14701 1870
rect 14557 1836 14591 1846
rect 13728 1802 13751 1836
rect 13785 1802 13819 1836
rect 13853 1802 13887 1836
rect 13921 1802 13955 1836
rect 13989 1802 14023 1836
rect 14057 1802 14091 1836
rect 14125 1802 14159 1836
rect 14193 1802 14227 1836
rect 14261 1802 14295 1836
rect 14329 1802 14363 1836
rect 14397 1826 14591 1836
rect 14397 1802 14455 1826
rect 13728 1792 14455 1802
rect 14489 1812 14591 1826
rect 14625 1812 14701 1846
rect 14489 1801 14701 1812
rect 14489 1792 14523 1801
rect 13728 1767 14523 1792
rect 14557 1776 14701 1801
rect 14557 1767 14591 1776
rect 13728 1764 14591 1767
rect 13728 1730 13751 1764
rect 13785 1730 13819 1764
rect 13853 1730 13887 1764
rect 13921 1730 13955 1764
rect 13989 1730 14023 1764
rect 14057 1730 14091 1764
rect 14125 1730 14159 1764
rect 14193 1730 14227 1764
rect 14261 1730 14295 1764
rect 14329 1730 14363 1764
rect 14397 1755 14591 1764
rect 14397 1730 14455 1755
rect 13728 1721 14455 1730
rect 14489 1742 14591 1755
rect 14625 1742 14701 1776
rect 14489 1732 14701 1742
rect 14489 1721 14523 1732
rect 13728 1698 14523 1721
rect 14557 1706 14701 1732
rect 14557 1698 14591 1706
rect 13728 1692 14591 1698
rect 13728 1658 13751 1692
rect 13785 1658 13819 1692
rect 13853 1658 13887 1692
rect 13921 1658 13955 1692
rect 13989 1658 14023 1692
rect 14057 1658 14091 1692
rect 14125 1658 14159 1692
rect 14193 1658 14227 1692
rect 14261 1658 14295 1692
rect 14329 1658 14363 1692
rect 14397 1684 14591 1692
rect 14397 1658 14455 1684
rect 13728 1650 14455 1658
rect 14489 1672 14591 1684
rect 14625 1672 14701 1706
rect 14489 1663 14701 1672
rect 14489 1650 14523 1663
rect 13728 1629 14523 1650
rect 14557 1636 14701 1663
rect 14557 1629 14591 1636
rect 13728 1620 14591 1629
rect 13728 1586 13751 1620
rect 13785 1586 13819 1620
rect 13853 1586 13887 1620
rect 13921 1586 13955 1620
rect 13989 1586 14023 1620
rect 14057 1586 14091 1620
rect 14125 1586 14159 1620
rect 14193 1586 14227 1620
rect 14261 1586 14295 1620
rect 14329 1586 14363 1620
rect 14397 1613 14591 1620
rect 14397 1586 14455 1613
rect 10000 1557 10024 1583
rect 13728 1579 14455 1586
rect 14489 1602 14591 1613
rect 14625 1602 14701 1636
rect 14489 1594 14701 1602
rect 14489 1579 14523 1594
rect 13728 1560 14523 1579
rect 14557 1566 14701 1594
rect 14557 1560 14591 1566
rect 9929 1555 9936 1557
rect 10000 1555 10012 1557
rect 9894 1523 9936 1555
rect 9970 1523 10012 1555
rect 8388 1521 10046 1523
rect 1460 1487 1531 1519
rect 1565 1487 1600 1521
rect 1635 1519 1669 1521
rect 1634 1487 1669 1519
rect 1703 1487 1738 1521
rect 1772 1487 1807 1521
rect 1841 1487 1876 1521
rect 1910 1487 1945 1521
rect 1979 1487 2014 1521
rect 2048 1487 2083 1521
rect 2117 1487 2152 1521
rect 2186 1487 2221 1521
rect 2255 1487 2290 1521
rect 2324 1487 2359 1521
rect 2393 1487 2428 1521
rect 2462 1487 2497 1521
rect 2531 1487 2566 1521
rect 2600 1487 2635 1521
rect 2669 1487 2704 1521
rect 2738 1487 2773 1521
rect 2807 1487 2842 1521
rect 2876 1487 2911 1521
rect 2945 1487 2980 1521
rect 3014 1487 3049 1521
rect 3083 1487 3118 1521
rect 3152 1487 3187 1521
rect 3221 1487 3256 1521
rect 3290 1487 3325 1521
rect 3359 1487 3394 1521
rect 3428 1487 3463 1521
rect 3497 1487 3532 1521
rect 3566 1487 3601 1521
rect 3635 1487 3670 1521
rect 3704 1487 3739 1521
rect 3773 1487 3808 1521
rect 3842 1487 3877 1521
rect 3911 1487 3946 1521
rect 3980 1487 4015 1521
rect 4049 1487 4084 1521
rect 4118 1487 4153 1521
rect 4187 1487 4222 1521
rect 4256 1487 4291 1521
rect 4325 1487 4360 1521
rect 4394 1487 4429 1521
rect 4463 1487 4498 1521
rect 4532 1487 4567 1521
rect 4601 1487 4636 1521
rect 4670 1487 4705 1521
rect 4739 1487 4774 1521
rect 4808 1487 4843 1521
rect 4877 1487 4912 1521
rect 4946 1487 4981 1521
rect 5015 1487 5050 1521
rect 5084 1487 5119 1521
rect 5153 1487 5188 1521
rect 5222 1487 5257 1521
rect 5291 1487 5326 1521
rect 5360 1487 5395 1521
rect 5429 1487 5464 1521
rect 5498 1487 5533 1521
rect 5567 1487 5602 1521
rect 5636 1487 5671 1521
rect 5705 1487 5740 1521
rect 5774 1487 5809 1521
rect 5843 1487 5878 1521
rect 5912 1487 5947 1521
rect 5981 1487 6016 1521
rect 6050 1487 6085 1521
rect 6119 1487 6154 1521
rect 1460 1480 6154 1487
rect 8364 1487 8412 1521
rect 8446 1487 8482 1521
rect 8516 1487 8552 1521
rect 8586 1487 8622 1521
rect 8656 1487 8692 1521
rect 8726 1487 8762 1521
rect 8796 1487 8832 1521
rect 8866 1487 8902 1521
rect 8936 1487 8972 1521
rect 9006 1487 9043 1521
rect 9077 1487 9114 1521
rect 9148 1487 9185 1521
rect 9219 1487 9256 1521
rect 9290 1487 9327 1521
rect 9361 1487 9398 1521
rect 9432 1487 9469 1521
rect 9503 1487 9540 1521
rect 9574 1487 9611 1521
rect 9645 1487 9682 1521
rect 9716 1487 9753 1521
rect 9787 1487 9824 1521
rect 9858 1487 9895 1521
rect 9929 1487 9966 1521
rect 10000 1487 10046 1521
rect 8364 1485 10046 1487
rect 8364 1480 8434 1485
rect 1491 1446 1529 1480
rect 1563 1453 1601 1480
rect 1635 1453 1683 1480
rect 1717 1453 1757 1480
rect 1791 1453 1831 1480
rect 1865 1453 1905 1480
rect 1939 1453 1979 1480
rect 1460 1443 1531 1446
rect 1086 1419 1531 1443
rect 1565 1419 1600 1453
rect 1635 1446 1669 1453
rect 1717 1446 1738 1453
rect 1791 1446 1807 1453
rect 1865 1446 1876 1453
rect 1939 1446 1945 1453
rect 1634 1419 1669 1446
rect 1703 1419 1738 1446
rect 1772 1419 1807 1446
rect 1841 1419 1876 1446
rect 1910 1419 1945 1446
rect 2013 1453 2053 1480
rect 2087 1453 2127 1480
rect 2161 1453 2201 1480
rect 2235 1453 2276 1480
rect 2310 1453 2351 1480
rect 2385 1453 2426 1480
rect 2460 1453 2501 1480
rect 2535 1453 2576 1480
rect 2610 1453 2651 1480
rect 2685 1453 2726 1480
rect 2760 1453 2801 1480
rect 2835 1453 2876 1480
rect 2013 1446 2014 1453
rect 1979 1419 2014 1446
rect 2048 1446 2053 1453
rect 2117 1446 2127 1453
rect 2186 1446 2201 1453
rect 2255 1446 2276 1453
rect 2324 1446 2351 1453
rect 2393 1446 2426 1453
rect 2048 1419 2083 1446
rect 2117 1419 2152 1446
rect 2186 1419 2221 1446
rect 2255 1419 2290 1446
rect 2324 1419 2359 1446
rect 2393 1419 2428 1446
rect 2462 1419 2497 1453
rect 2535 1446 2566 1453
rect 2610 1446 2635 1453
rect 2685 1446 2704 1453
rect 2760 1446 2773 1453
rect 2835 1446 2842 1453
rect 2531 1419 2566 1446
rect 2600 1419 2635 1446
rect 2669 1419 2704 1446
rect 2738 1419 2773 1446
rect 2807 1419 2842 1446
rect 2910 1453 2951 1480
rect 2985 1453 6154 1480
rect 2910 1446 2911 1453
rect 2876 1419 2911 1446
rect 2945 1446 2951 1453
rect 2945 1419 2980 1446
rect 3014 1419 3049 1453
rect 3083 1419 3118 1453
rect 3152 1419 3187 1453
rect 3221 1419 3256 1453
rect 3290 1419 3325 1453
rect 3359 1419 3394 1453
rect 3428 1419 3463 1453
rect 3497 1419 3532 1453
rect 3566 1419 3601 1453
rect 3635 1419 3670 1453
rect 3704 1419 3739 1453
rect 3773 1419 3808 1453
rect 3842 1419 3877 1453
rect 3911 1419 3946 1453
rect 3980 1419 4015 1453
rect 4049 1419 4084 1453
rect 4118 1419 4153 1453
rect 4187 1419 4222 1453
rect 4256 1419 4291 1453
rect 4325 1419 4360 1453
rect 4394 1419 4429 1453
rect 4463 1419 4498 1453
rect 4532 1419 4567 1453
rect 4601 1419 4636 1453
rect 4670 1419 4705 1453
rect 4739 1419 4774 1453
rect 4808 1419 4843 1453
rect 4877 1419 4912 1453
rect 4946 1419 4981 1453
rect 5015 1419 5050 1453
rect 5084 1419 5119 1453
rect 5153 1419 5188 1453
rect 5222 1419 5257 1453
rect 5291 1419 5326 1453
rect 5360 1419 5395 1453
rect 5429 1419 5464 1453
rect 5498 1419 5533 1453
rect 5567 1419 5602 1453
rect 5636 1419 5671 1453
rect 5705 1419 5740 1453
rect 5774 1419 5809 1453
rect 5843 1419 5878 1453
rect 5912 1419 5947 1453
rect 5981 1419 6016 1453
rect 6050 1419 6085 1453
rect 6119 1419 6154 1453
rect 8396 1453 8434 1480
rect 8468 1453 8509 1485
rect 8543 1453 8584 1485
rect 8618 1453 8659 1485
rect 8693 1453 8734 1485
rect 8768 1453 8809 1485
rect 8843 1453 8884 1485
rect 8918 1453 8959 1485
rect 8993 1453 9034 1485
rect 9068 1453 9109 1485
rect 9143 1453 9184 1485
rect 9218 1453 9259 1485
rect 9293 1453 9334 1485
rect 9368 1453 9409 1485
rect 9443 1453 9484 1485
rect 9518 1453 9559 1485
rect 9593 1453 9634 1485
rect 9668 1453 9709 1485
rect 9743 1453 9784 1485
rect 9818 1453 9860 1485
rect 8396 1446 8412 1453
rect 8468 1451 8482 1453
rect 8543 1451 8552 1453
rect 8618 1451 8622 1453
rect 8364 1419 8412 1446
rect 8446 1419 8482 1451
rect 8516 1419 8552 1451
rect 8586 1419 8622 1451
rect 8656 1451 8659 1453
rect 8726 1451 8734 1453
rect 8796 1451 8809 1453
rect 8866 1451 8884 1453
rect 8936 1451 8959 1453
rect 9006 1451 9034 1453
rect 9077 1451 9109 1453
rect 9148 1451 9184 1453
rect 8656 1419 8692 1451
rect 8726 1419 8762 1451
rect 8796 1419 8832 1451
rect 8866 1419 8902 1451
rect 8936 1419 8972 1451
rect 9006 1419 9043 1451
rect 9077 1419 9114 1451
rect 9148 1419 9185 1451
rect 9219 1419 9256 1453
rect 9293 1451 9327 1453
rect 9368 1451 9398 1453
rect 9443 1451 9469 1453
rect 9518 1451 9540 1453
rect 9593 1451 9611 1453
rect 9668 1451 9682 1453
rect 9743 1451 9753 1453
rect 9818 1451 9824 1453
rect 9290 1419 9327 1451
rect 9361 1419 9398 1451
rect 9432 1419 9469 1451
rect 9503 1419 9540 1451
rect 9574 1419 9611 1451
rect 9645 1419 9682 1451
rect 9716 1419 9753 1451
rect 9787 1419 9824 1451
rect 9858 1451 9860 1453
rect 9894 1453 9936 1485
rect 9970 1453 10012 1485
rect 9894 1451 9895 1453
rect 9858 1419 9895 1451
rect 9929 1451 9936 1453
rect 10000 1451 10012 1453
rect 13728 1548 14591 1560
rect 13728 1514 13751 1548
rect 13785 1514 13819 1548
rect 13853 1514 13887 1548
rect 13921 1514 13955 1548
rect 13989 1514 14023 1548
rect 14057 1514 14091 1548
rect 14125 1514 14159 1548
rect 14193 1514 14227 1548
rect 14261 1514 14295 1548
rect 14329 1514 14363 1548
rect 14397 1541 14591 1548
rect 14397 1514 14455 1541
rect 13728 1507 14455 1514
rect 14489 1532 14591 1541
rect 14625 1532 14701 1566
rect 14489 1525 14701 1532
rect 14489 1507 14523 1525
rect 13728 1494 14523 1507
rect 14557 1496 14701 1525
rect 14557 1494 14591 1496
rect 14625 1494 14701 1496
rect 19563 2027 19598 2061
rect 19632 2027 19667 2061
rect 19701 2027 19736 2061
rect 19770 2027 19805 2061
rect 19839 2027 19874 2061
rect 19908 2027 19943 2061
rect 19977 2027 20012 2061
rect 20046 2027 20081 2061
rect 20115 2027 20150 2061
rect 20184 2027 20219 2061
rect 20253 2027 20288 2061
rect 20322 2027 20357 2061
rect 20391 2027 20426 2061
rect 20460 2027 20495 2061
rect 20529 2027 20564 2061
rect 20598 2027 20633 2061
rect 20667 2027 20702 2061
rect 20736 2027 20771 2061
rect 20805 2027 20840 2061
rect 20874 2027 20909 2061
rect 20943 2027 20978 2061
rect 21012 2027 21047 2061
rect 21081 2027 21116 2061
rect 21150 2027 21185 2061
rect 21219 2027 21254 2061
rect 21288 2027 21323 2061
rect 21357 2027 21392 2061
rect 21426 2027 21461 2061
rect 21495 2027 21530 2061
rect 21564 2027 21599 2061
rect 21633 2027 21668 2061
rect 21702 2027 21737 2061
rect 21771 2027 21806 2061
rect 21840 2027 21875 2061
rect 21909 2027 21944 2061
rect 21978 2027 22013 2061
rect 22047 2027 22082 2061
rect 22116 2027 22151 2061
rect 22185 2027 22220 2061
rect 22254 2027 22289 2061
rect 22323 2027 22358 2061
rect 22392 2027 22427 2061
rect 22461 2027 22496 2061
rect 22530 2027 22565 2061
rect 22599 2027 22634 2061
rect 22668 2027 22703 2061
rect 22737 2027 22772 2061
rect 22806 2027 22841 2061
rect 22875 2027 22910 2061
rect 22944 2027 22979 2061
rect 23013 2027 23048 2061
rect 23082 2027 23117 2061
rect 23151 2027 23186 2061
rect 23220 2027 23255 2061
rect 23289 2027 23324 2061
rect 23358 2027 23393 2061
rect 23427 2027 23462 2061
rect 23496 2027 23531 2061
rect 23565 2046 23600 2061
rect 23634 2046 23669 2061
rect 23703 2046 23738 2061
rect 23565 2027 23593 2046
rect 23634 2027 23665 2046
rect 23703 2027 23737 2046
rect 23772 2027 23796 2061
rect 19563 2012 23593 2027
rect 23627 2012 23665 2027
rect 23699 2012 23737 2027
rect 23771 2012 23796 2027
rect 19563 1993 23796 2012
rect 19563 1959 19598 1993
rect 19632 1959 19667 1993
rect 19701 1959 19736 1993
rect 19770 1959 19805 1993
rect 19839 1959 19874 1993
rect 19908 1959 19943 1993
rect 19977 1959 20012 1993
rect 20046 1959 20081 1993
rect 20115 1959 20150 1993
rect 20184 1959 20219 1993
rect 20253 1959 20288 1993
rect 20322 1959 20357 1993
rect 20391 1959 20426 1993
rect 20460 1959 20495 1993
rect 20529 1959 20564 1993
rect 20598 1959 20633 1993
rect 20667 1959 20702 1993
rect 20736 1959 20771 1993
rect 20805 1959 20840 1993
rect 20874 1959 20909 1993
rect 20943 1959 20978 1993
rect 21012 1959 21047 1993
rect 21081 1959 21116 1993
rect 21150 1959 21185 1993
rect 21219 1959 21254 1993
rect 21288 1959 21323 1993
rect 21357 1959 21392 1993
rect 21426 1959 21461 1993
rect 21495 1959 21530 1993
rect 21564 1959 21599 1993
rect 21633 1959 21668 1993
rect 21702 1959 21737 1993
rect 21771 1959 21806 1993
rect 21840 1959 21875 1993
rect 21909 1959 21944 1993
rect 21978 1959 22013 1993
rect 22047 1959 22082 1993
rect 22116 1959 22151 1993
rect 22185 1959 22220 1993
rect 22254 1959 22289 1993
rect 22323 1959 22358 1993
rect 22392 1959 22427 1993
rect 22461 1959 22496 1993
rect 22530 1959 22565 1993
rect 22599 1959 22634 1993
rect 22668 1959 22703 1993
rect 22737 1959 22772 1993
rect 22806 1959 22841 1993
rect 22875 1959 22910 1993
rect 22944 1959 22979 1993
rect 23013 1959 23048 1993
rect 23082 1959 23117 1993
rect 23151 1959 23186 1993
rect 23220 1959 23255 1993
rect 23289 1959 23324 1993
rect 23358 1959 23393 1993
rect 23427 1959 23462 1993
rect 23496 1959 23531 1993
rect 23565 1972 23600 1993
rect 23634 1972 23669 1993
rect 23703 1972 23738 1993
rect 23565 1959 23593 1972
rect 23634 1959 23665 1972
rect 23703 1959 23737 1972
rect 23772 1959 23796 1993
rect 19563 1938 23593 1959
rect 23627 1938 23665 1959
rect 23699 1938 23737 1959
rect 23771 1938 23796 1959
rect 19563 1925 23796 1938
rect 19563 1891 19598 1925
rect 19632 1891 19667 1925
rect 19701 1891 19736 1925
rect 19770 1891 19805 1925
rect 19839 1891 19874 1925
rect 19908 1891 19943 1925
rect 19977 1891 20012 1925
rect 20046 1891 20081 1925
rect 20115 1891 20150 1925
rect 20184 1891 20219 1925
rect 20253 1891 20288 1925
rect 20322 1891 20357 1925
rect 20391 1891 20426 1925
rect 20460 1891 20495 1925
rect 20529 1891 20564 1925
rect 20598 1891 20633 1925
rect 20667 1891 20702 1925
rect 20736 1891 20771 1925
rect 20805 1891 20840 1925
rect 20874 1891 20909 1925
rect 20943 1891 20978 1925
rect 21012 1891 21047 1925
rect 21081 1891 21116 1925
rect 21150 1891 21185 1925
rect 21219 1891 21254 1925
rect 21288 1891 21323 1925
rect 21357 1891 21392 1925
rect 21426 1891 21461 1925
rect 21495 1891 21530 1925
rect 21564 1891 21599 1925
rect 21633 1891 21668 1925
rect 21702 1891 21737 1925
rect 21771 1891 21806 1925
rect 21840 1891 21875 1925
rect 21909 1891 21944 1925
rect 21978 1891 22013 1925
rect 22047 1891 22082 1925
rect 22116 1891 22151 1925
rect 22185 1891 22220 1925
rect 22254 1891 22289 1925
rect 22323 1891 22358 1925
rect 22392 1891 22427 1925
rect 22461 1891 22496 1925
rect 22530 1891 22565 1925
rect 22599 1891 22634 1925
rect 22668 1891 22703 1925
rect 22737 1891 22772 1925
rect 22806 1891 22841 1925
rect 22875 1891 22910 1925
rect 22944 1891 22979 1925
rect 23013 1891 23048 1925
rect 23082 1891 23117 1925
rect 23151 1891 23186 1925
rect 23220 1891 23255 1925
rect 23289 1891 23324 1925
rect 23358 1891 23393 1925
rect 23427 1891 23462 1925
rect 23496 1891 23531 1925
rect 23565 1891 23600 1925
rect 23634 1891 23669 1925
rect 23703 1891 23738 1925
rect 23772 1891 23796 1925
rect 19563 1857 23796 1891
rect 19563 1823 19598 1857
rect 19632 1823 19667 1857
rect 19701 1823 19736 1857
rect 19770 1823 19805 1857
rect 19839 1823 19874 1857
rect 19908 1823 19943 1857
rect 19977 1823 20012 1857
rect 20046 1823 20081 1857
rect 20115 1823 20150 1857
rect 20184 1823 20219 1857
rect 20253 1823 20288 1857
rect 20322 1823 20357 1857
rect 20391 1823 20426 1857
rect 20460 1823 20495 1857
rect 20529 1823 20564 1857
rect 20598 1823 20633 1857
rect 20667 1823 20702 1857
rect 20736 1823 20771 1857
rect 20805 1823 20840 1857
rect 20874 1823 20909 1857
rect 20943 1823 20978 1857
rect 21012 1823 21047 1857
rect 21081 1823 21116 1857
rect 21150 1823 21185 1857
rect 21219 1823 21254 1857
rect 21288 1823 21323 1857
rect 21357 1823 21392 1857
rect 21426 1823 21461 1857
rect 21495 1823 21530 1857
rect 21564 1823 21599 1857
rect 21633 1823 21668 1857
rect 21702 1823 21737 1857
rect 21771 1823 21806 1857
rect 21840 1823 21875 1857
rect 21909 1823 21944 1857
rect 21978 1823 22013 1857
rect 22047 1823 22082 1857
rect 22116 1823 22151 1857
rect 22185 1823 22220 1857
rect 22254 1823 22289 1857
rect 22323 1823 22358 1857
rect 22392 1823 22427 1857
rect 22461 1823 22496 1857
rect 22530 1823 22565 1857
rect 22599 1823 22634 1857
rect 22668 1823 22703 1857
rect 22737 1823 22772 1857
rect 22806 1823 22841 1857
rect 22875 1823 22910 1857
rect 22944 1823 22979 1857
rect 23013 1823 23048 1857
rect 23082 1823 23117 1857
rect 23151 1823 23186 1857
rect 23220 1823 23255 1857
rect 23289 1823 23324 1857
rect 23358 1823 23393 1857
rect 23427 1823 23462 1857
rect 23496 1823 23531 1857
rect 23565 1823 23600 1857
rect 23634 1823 23669 1857
rect 23703 1823 23738 1857
rect 23772 1823 23796 1857
rect 19563 1789 23796 1823
rect 19563 1755 19598 1789
rect 19632 1755 19667 1789
rect 19701 1755 19736 1789
rect 19770 1755 19805 1789
rect 19839 1755 19874 1789
rect 19908 1755 19943 1789
rect 19977 1755 20012 1789
rect 20046 1755 20081 1789
rect 20115 1755 20150 1789
rect 20184 1755 20219 1789
rect 20253 1755 20288 1789
rect 20322 1755 20357 1789
rect 20391 1755 20426 1789
rect 20460 1755 20495 1789
rect 20529 1755 20564 1789
rect 20598 1755 20633 1789
rect 20667 1755 20702 1789
rect 20736 1755 20771 1789
rect 20805 1755 20840 1789
rect 20874 1755 20909 1789
rect 20943 1755 20978 1789
rect 21012 1755 21047 1789
rect 21081 1755 21116 1789
rect 21150 1755 21185 1789
rect 21219 1755 21254 1789
rect 21288 1755 21323 1789
rect 21357 1755 21392 1789
rect 21426 1755 21461 1789
rect 21495 1755 21530 1789
rect 21564 1755 21599 1789
rect 21633 1755 21668 1789
rect 21702 1755 21737 1789
rect 21771 1755 21806 1789
rect 21840 1755 21875 1789
rect 21909 1755 21944 1789
rect 21978 1755 22013 1789
rect 22047 1755 22082 1789
rect 22116 1755 22151 1789
rect 22185 1755 22220 1789
rect 22254 1755 22289 1789
rect 22323 1755 22358 1789
rect 22392 1755 22427 1789
rect 22461 1755 22496 1789
rect 22530 1755 22565 1789
rect 22599 1755 22634 1789
rect 22668 1755 22703 1789
rect 22737 1755 22772 1789
rect 22806 1755 22841 1789
rect 22875 1755 22910 1789
rect 22944 1755 22979 1789
rect 23013 1755 23048 1789
rect 23082 1755 23117 1789
rect 23151 1755 23186 1789
rect 23220 1755 23255 1789
rect 23289 1755 23324 1789
rect 23358 1755 23393 1789
rect 23427 1755 23462 1789
rect 23496 1755 23531 1789
rect 23565 1755 23600 1789
rect 23634 1755 23669 1789
rect 23703 1755 23738 1789
rect 23772 1755 23796 1789
rect 19563 1721 23796 1755
rect 19563 1687 19598 1721
rect 19632 1687 19667 1721
rect 19701 1687 19736 1721
rect 19770 1687 19805 1721
rect 19839 1687 19874 1721
rect 19908 1687 19943 1721
rect 19977 1687 20012 1721
rect 20046 1687 20081 1721
rect 20115 1687 20150 1721
rect 20184 1687 20219 1721
rect 20253 1687 20288 1721
rect 20322 1687 20357 1721
rect 20391 1687 20426 1721
rect 20460 1687 20495 1721
rect 20529 1687 20564 1721
rect 20598 1687 20633 1721
rect 20667 1687 20702 1721
rect 20736 1687 20771 1721
rect 20805 1687 20840 1721
rect 20874 1687 20909 1721
rect 20943 1687 20978 1721
rect 21012 1687 21047 1721
rect 21081 1687 21116 1721
rect 21150 1687 21185 1721
rect 21219 1687 21254 1721
rect 21288 1687 21323 1721
rect 21357 1687 21392 1721
rect 21426 1687 21461 1721
rect 21495 1687 21530 1721
rect 21564 1687 21599 1721
rect 21633 1687 21668 1721
rect 21702 1687 21737 1721
rect 21771 1687 21806 1721
rect 21840 1687 21875 1721
rect 21909 1687 21944 1721
rect 21978 1687 22013 1721
rect 22047 1687 22082 1721
rect 22116 1687 22151 1721
rect 22185 1687 22220 1721
rect 22254 1687 22289 1721
rect 22323 1687 22358 1721
rect 22392 1687 22427 1721
rect 22461 1687 22496 1721
rect 22530 1687 22565 1721
rect 22599 1687 22634 1721
rect 22668 1687 22703 1721
rect 22737 1687 22772 1721
rect 22806 1687 22841 1721
rect 22875 1687 22910 1721
rect 22944 1687 22979 1721
rect 23013 1687 23048 1721
rect 23082 1687 23117 1721
rect 23151 1687 23186 1721
rect 23220 1687 23255 1721
rect 23289 1687 23324 1721
rect 23358 1687 23393 1721
rect 23427 1687 23462 1721
rect 23496 1687 23531 1721
rect 23565 1687 23600 1721
rect 23634 1687 23669 1721
rect 23703 1687 23738 1721
rect 23772 1687 23796 1721
rect 19563 1653 23796 1687
rect 19563 1619 19598 1653
rect 19632 1619 19667 1653
rect 19701 1619 19736 1653
rect 19770 1619 19805 1653
rect 19839 1619 19874 1653
rect 19908 1619 19943 1653
rect 19977 1619 20012 1653
rect 20046 1619 20081 1653
rect 20115 1619 20150 1653
rect 20184 1619 20219 1653
rect 20253 1619 20288 1653
rect 20322 1619 20357 1653
rect 20391 1619 20426 1653
rect 20460 1619 20495 1653
rect 20529 1619 20564 1653
rect 20598 1619 20633 1653
rect 20667 1619 20702 1653
rect 20736 1619 20771 1653
rect 20805 1619 20840 1653
rect 20874 1619 20909 1653
rect 20943 1619 20978 1653
rect 21012 1619 21047 1653
rect 21081 1619 21116 1653
rect 21150 1619 21185 1653
rect 21219 1619 21254 1653
rect 21288 1619 21323 1653
rect 21357 1619 21392 1653
rect 21426 1619 21461 1653
rect 21495 1619 21530 1653
rect 21564 1619 21599 1653
rect 21633 1619 21668 1653
rect 21702 1619 21737 1653
rect 21771 1619 21806 1653
rect 21840 1619 21875 1653
rect 21909 1619 21944 1653
rect 21978 1619 22013 1653
rect 22047 1619 22082 1653
rect 22116 1619 22151 1653
rect 22185 1619 22220 1653
rect 22254 1619 22289 1653
rect 22323 1619 22358 1653
rect 22392 1619 22427 1653
rect 22461 1619 22496 1653
rect 22530 1619 22565 1653
rect 22599 1619 22634 1653
rect 22668 1619 22703 1653
rect 22737 1619 22772 1653
rect 22806 1619 22841 1653
rect 22875 1619 22910 1653
rect 22944 1619 22979 1653
rect 23013 1619 23048 1653
rect 23082 1619 23117 1653
rect 23151 1619 23186 1653
rect 23220 1619 23255 1653
rect 23289 1619 23324 1653
rect 23358 1619 23393 1653
rect 23427 1619 23462 1653
rect 23496 1619 23531 1653
rect 23565 1619 23600 1653
rect 23634 1619 23669 1653
rect 23703 1619 23738 1653
rect 23772 1619 23796 1653
rect 19563 1585 23796 1619
rect 19563 1551 19598 1585
rect 19632 1551 19667 1585
rect 19701 1551 19736 1585
rect 19770 1551 19805 1585
rect 19839 1551 19874 1585
rect 19908 1551 19943 1585
rect 19977 1551 20012 1585
rect 20046 1551 20081 1585
rect 20115 1551 20150 1585
rect 20184 1551 20219 1585
rect 20253 1551 20288 1585
rect 20322 1551 20357 1585
rect 20391 1551 20426 1585
rect 20460 1551 20495 1585
rect 20529 1551 20564 1585
rect 20598 1551 20633 1585
rect 20667 1551 20702 1585
rect 20736 1551 20771 1585
rect 20805 1551 20840 1585
rect 20874 1551 20909 1585
rect 20943 1551 20978 1585
rect 21012 1551 21047 1585
rect 21081 1551 21116 1585
rect 21150 1551 21185 1585
rect 21219 1551 21254 1585
rect 21288 1551 21323 1585
rect 21357 1551 21392 1585
rect 21426 1551 21461 1585
rect 21495 1551 21530 1585
rect 21564 1551 21599 1585
rect 21633 1551 21668 1585
rect 21702 1551 21737 1585
rect 21771 1551 21806 1585
rect 21840 1551 21875 1585
rect 21909 1551 21944 1585
rect 21978 1551 22013 1585
rect 22047 1551 22082 1585
rect 22116 1551 22151 1585
rect 22185 1551 22220 1585
rect 22254 1551 22289 1585
rect 22323 1551 22358 1585
rect 22392 1551 22427 1585
rect 22461 1551 22496 1585
rect 22530 1551 22565 1585
rect 22599 1551 22634 1585
rect 22668 1551 22703 1585
rect 22737 1551 22772 1585
rect 22806 1551 22841 1585
rect 22875 1551 22910 1585
rect 22944 1551 22979 1585
rect 23013 1551 23048 1585
rect 23082 1551 23117 1585
rect 23151 1551 23186 1585
rect 23220 1551 23255 1585
rect 23289 1551 23324 1585
rect 23358 1551 23393 1585
rect 23427 1551 23462 1585
rect 23496 1551 23531 1585
rect 23565 1551 23600 1585
rect 23634 1551 23669 1585
rect 23703 1551 23738 1585
rect 23772 1551 23796 1585
rect 19563 1517 23796 1551
rect 19563 1494 19598 1517
rect 19632 1494 19667 1517
rect 19701 1494 19736 1517
rect 19770 1494 19805 1517
rect 19839 1494 19874 1517
rect 19908 1494 19943 1517
rect 19977 1494 20012 1517
rect 20046 1494 20081 1517
rect 20115 1494 20150 1517
rect 20184 1494 20219 1517
rect 20253 1494 20288 1517
rect 20322 1494 20357 1517
rect 20391 1494 20426 1517
rect 20460 1494 20495 1517
rect 20529 1494 20564 1517
rect 20598 1494 20633 1517
rect 20667 1494 20702 1517
rect 20736 1494 20771 1517
rect 20805 1494 20840 1517
rect 20874 1494 20909 1517
rect 20943 1494 20978 1517
rect 21012 1494 21047 1517
rect 21081 1494 21116 1517
rect 21150 1494 21185 1517
rect 21219 1494 21254 1517
rect 21288 1494 21323 1517
rect 21357 1494 21392 1517
rect 21426 1494 21461 1517
rect 21495 1494 21530 1517
rect 21564 1494 21599 1517
rect 21633 1494 21668 1517
rect 21702 1494 21737 1517
rect 21771 1494 21806 1517
rect 21840 1494 21875 1517
rect 21909 1494 21944 1517
rect 21978 1494 22013 1517
rect 22047 1494 22082 1517
rect 22116 1494 22151 1517
rect 22185 1494 22220 1517
rect 22254 1494 22289 1517
rect 22323 1494 22358 1517
rect 22392 1494 22427 1517
rect 22461 1494 22496 1517
rect 22530 1494 22565 1517
rect 22599 1494 22634 1517
rect 22668 1494 22703 1517
rect 22737 1494 22772 1517
rect 22806 1494 22841 1517
rect 22875 1494 22910 1517
rect 22944 1494 22979 1517
rect 23013 1494 23048 1517
rect 13728 1475 14493 1494
rect 14557 1491 14566 1494
rect 9929 1419 9966 1451
rect 10000 1425 10024 1451
rect 13728 1441 13751 1475
rect 13785 1441 13819 1475
rect 13853 1441 13887 1475
rect 13921 1441 13955 1475
rect 13989 1441 14023 1475
rect 14057 1441 14091 1475
rect 14125 1441 14159 1475
rect 14193 1441 14227 1475
rect 14261 1441 14295 1475
rect 14329 1441 14363 1475
rect 14397 1469 14493 1475
rect 14397 1441 14455 1469
rect 13728 1435 14455 1441
rect 14489 1460 14493 1469
rect 14527 1460 14566 1491
rect 14625 1462 14639 1494
rect 14600 1460 14639 1462
rect 14673 1460 14701 1494
rect 14489 1456 14701 1460
rect 14489 1435 14523 1456
rect 10000 1419 13559 1425
rect 1086 1408 13559 1419
rect 1086 1374 1683 1408
rect 1717 1374 1757 1408
rect 1791 1374 1831 1408
rect 1865 1374 1905 1408
rect 1939 1374 1979 1408
rect 2013 1374 2053 1408
rect 2087 1374 2127 1408
rect 2161 1374 2201 1408
rect 2235 1374 2276 1408
rect 2310 1374 2351 1408
rect 2385 1374 2426 1408
rect 2460 1374 2501 1408
rect 2535 1374 2576 1408
rect 2610 1374 2651 1408
rect 2685 1374 2726 1408
rect 2760 1374 2801 1408
rect 2835 1374 2876 1408
rect 2910 1374 2951 1408
rect 2985 1374 7117 1408
rect 7151 1374 7190 1408
rect 7224 1374 7263 1408
rect 7297 1374 7336 1408
rect 7370 1374 7409 1408
rect 7443 1374 7482 1408
rect 7516 1374 7555 1408
rect 7589 1374 7628 1408
rect 7662 1374 7701 1408
rect 7735 1374 7774 1408
rect 7808 1374 7847 1408
rect 7881 1374 7920 1408
rect 7954 1374 7993 1408
rect 8027 1374 8066 1408
rect 8100 1374 8140 1408
rect 8174 1374 8214 1408
rect 8248 1374 8288 1408
rect 8322 1374 8362 1408
rect 8396 1374 13559 1408
rect 1086 1317 13559 1374
rect 13728 1422 14523 1435
rect 14557 1426 14701 1456
rect 14557 1422 14591 1426
rect 14625 1422 14701 1426
rect 13728 1402 14493 1422
rect 13728 1368 13751 1402
rect 13785 1368 13819 1402
rect 13853 1368 13887 1402
rect 13921 1368 13955 1402
rect 13989 1368 14023 1402
rect 14057 1368 14091 1402
rect 14125 1368 14159 1402
rect 14193 1368 14227 1402
rect 14261 1368 14295 1402
rect 14329 1368 14363 1402
rect 14397 1397 14493 1402
rect 14397 1368 14455 1397
rect 13728 1363 14455 1368
rect 14489 1388 14493 1397
rect 14527 1388 14566 1422
rect 14625 1392 14639 1422
rect 14600 1388 14639 1392
rect 14673 1388 14701 1422
rect 14489 1387 14701 1388
rect 14489 1363 14523 1387
rect 13728 1353 14523 1363
rect 14557 1356 14701 1387
rect 14557 1353 14591 1356
rect 13728 1350 14591 1353
rect 14625 1350 14701 1356
rect 13728 1329 14493 1350
rect 696 1281 764 1297
rect 730 1259 764 1281
rect 13728 1267 13751 1329
rect 866 1261 13751 1267
rect 14397 1325 14493 1329
rect 14397 1291 14455 1325
rect 14489 1316 14493 1325
rect 14527 1318 14566 1350
rect 14625 1322 14639 1350
rect 14557 1316 14566 1318
rect 14600 1316 14639 1322
rect 14673 1316 14701 1350
rect 14489 1291 14523 1316
rect 14397 1284 14523 1291
rect 14557 1286 14701 1316
rect 14557 1284 14591 1286
rect 14397 1278 14591 1284
rect 14625 1278 14701 1286
rect 696 1225 728 1247
rect 762 1225 764 1259
rect 696 1212 764 1225
rect 934 1227 969 1261
rect 1003 1227 1038 1261
rect 1072 1227 1107 1261
rect 1141 1227 1176 1261
rect 1210 1227 1245 1261
rect 1279 1227 1314 1261
rect 1348 1227 1383 1261
rect 1417 1227 1452 1261
rect 1486 1227 1521 1261
rect 1555 1227 1590 1261
rect 1624 1227 1659 1261
rect 1693 1227 1728 1261
rect 1762 1227 1797 1261
rect 1831 1227 1866 1261
rect 1900 1227 1935 1261
rect 1969 1227 2004 1261
rect 2038 1227 2073 1261
rect 2107 1227 2142 1261
rect 2176 1227 2211 1261
rect 2245 1227 2280 1261
rect 2314 1227 2349 1261
rect 2383 1227 2418 1261
rect 2452 1227 2487 1261
rect 2521 1227 2556 1261
rect 2590 1227 2625 1261
rect 2659 1227 2694 1261
rect 2728 1227 2763 1261
rect 2797 1227 2832 1261
rect 2866 1227 2901 1261
rect 2935 1227 2970 1261
rect 3004 1227 3039 1261
rect 3073 1227 3108 1261
rect 3142 1227 3177 1261
rect 3211 1227 3246 1261
rect 3280 1227 3315 1261
rect 3349 1227 3384 1261
rect 3418 1227 3453 1261
rect 3487 1227 3522 1261
rect 3556 1227 3591 1261
rect 3625 1227 3660 1261
rect 3694 1227 3729 1261
rect 3763 1227 3798 1261
rect 3832 1227 3867 1261
rect 3901 1227 3936 1261
rect 3970 1227 4005 1261
rect 4039 1227 4074 1261
rect 4108 1227 4143 1261
rect 4177 1227 4212 1261
rect 4246 1227 4281 1261
rect 4315 1227 4350 1261
rect 4384 1227 4419 1261
rect 4453 1227 4488 1261
rect 4522 1227 4557 1261
rect 4591 1227 4626 1261
rect 4660 1227 4695 1261
rect 4729 1227 4764 1261
rect 4798 1227 4833 1261
rect 4867 1227 4902 1261
rect 4936 1227 4971 1261
rect 5005 1227 5040 1261
rect 5074 1227 5109 1261
rect 5143 1227 5178 1261
rect 5212 1227 5247 1261
rect 5281 1227 5316 1261
rect 5350 1227 5385 1261
rect 5419 1227 5454 1261
rect 5488 1227 5523 1261
rect 730 1187 764 1212
rect 934 1193 5523 1227
rect 696 1153 728 1178
rect 762 1153 764 1187
rect 696 1143 764 1153
rect 934 1159 969 1193
rect 1003 1159 1038 1193
rect 1072 1159 1107 1193
rect 1141 1159 1176 1193
rect 1210 1159 1245 1193
rect 1279 1159 1314 1193
rect 1348 1159 1383 1193
rect 1417 1159 1452 1193
rect 1486 1159 1521 1193
rect 1555 1159 1590 1193
rect 1624 1159 1659 1193
rect 1693 1159 1728 1193
rect 1762 1159 1797 1193
rect 1831 1159 1866 1193
rect 1900 1159 1935 1193
rect 1969 1159 2004 1193
rect 2038 1159 2073 1193
rect 2107 1159 2142 1193
rect 2176 1159 2211 1193
rect 2245 1159 2280 1193
rect 2314 1159 2349 1193
rect 2383 1159 2418 1193
rect 2452 1159 2487 1193
rect 2521 1159 2556 1193
rect 2590 1159 2625 1193
rect 2659 1159 2694 1193
rect 2728 1159 2763 1193
rect 2797 1159 2832 1193
rect 2866 1159 2901 1193
rect 2935 1159 2970 1193
rect 3004 1159 3039 1193
rect 3073 1159 3108 1193
rect 3142 1159 3177 1193
rect 3211 1159 3246 1193
rect 3280 1159 3315 1193
rect 3349 1159 3384 1193
rect 3418 1159 3453 1193
rect 3487 1159 3522 1193
rect 3556 1159 3591 1193
rect 3625 1159 3660 1193
rect 3694 1159 3729 1193
rect 3763 1159 3798 1193
rect 3832 1159 3867 1193
rect 3901 1159 3936 1193
rect 3970 1159 4005 1193
rect 4039 1159 4074 1193
rect 4108 1159 4143 1193
rect 4177 1159 4212 1193
rect 4246 1159 4281 1193
rect 4315 1159 4350 1193
rect 4384 1159 4419 1193
rect 4453 1159 4488 1193
rect 4522 1159 4557 1193
rect 4591 1159 4626 1193
rect 4660 1159 4695 1193
rect 4729 1159 4764 1193
rect 4798 1159 4833 1193
rect 4867 1159 4902 1193
rect 4936 1159 4971 1193
rect 5005 1159 5040 1193
rect 5074 1159 5109 1193
rect 5143 1159 5178 1193
rect 5212 1159 5247 1193
rect 5281 1159 5316 1193
rect 5350 1159 5385 1193
rect 5419 1159 5454 1193
rect 5488 1159 5523 1193
rect 730 1115 764 1143
rect 934 1125 5523 1159
rect 696 1081 728 1109
rect 762 1081 764 1115
rect 934 1091 969 1125
rect 1003 1091 1038 1125
rect 1072 1091 1107 1125
rect 1141 1091 1176 1125
rect 1210 1091 1245 1125
rect 1279 1091 1314 1125
rect 1348 1091 1383 1125
rect 1417 1091 1452 1125
rect 1486 1091 1521 1125
rect 1555 1091 1590 1125
rect 1624 1091 1659 1125
rect 1693 1091 1728 1125
rect 1762 1091 1797 1125
rect 1831 1091 1866 1125
rect 1900 1091 1935 1125
rect 1969 1091 2004 1125
rect 2038 1091 2073 1125
rect 2107 1091 2142 1125
rect 2176 1091 2211 1125
rect 2245 1091 2280 1125
rect 2314 1091 2349 1125
rect 2383 1091 2418 1125
rect 2452 1091 2487 1125
rect 2521 1091 2556 1125
rect 2590 1091 2625 1125
rect 2659 1091 2694 1125
rect 2728 1091 2763 1125
rect 2797 1091 2832 1125
rect 2866 1091 2901 1125
rect 2935 1091 2970 1125
rect 3004 1091 3039 1125
rect 3073 1091 3108 1125
rect 3142 1091 3177 1125
rect 3211 1091 3246 1125
rect 3280 1091 3315 1125
rect 3349 1091 3384 1125
rect 3418 1091 3453 1125
rect 3487 1091 3522 1125
rect 3556 1091 3591 1125
rect 3625 1091 3660 1125
rect 3694 1091 3729 1125
rect 3763 1091 3798 1125
rect 3832 1091 3867 1125
rect 3901 1091 3936 1125
rect 3970 1091 4005 1125
rect 4039 1091 4074 1125
rect 4108 1091 4143 1125
rect 4177 1091 4212 1125
rect 4246 1091 4281 1125
rect 4315 1091 4350 1125
rect 4384 1091 4419 1125
rect 4453 1091 4488 1125
rect 4522 1091 4557 1125
rect 4591 1091 4626 1125
rect 4660 1091 4695 1125
rect 4729 1091 4764 1125
rect 4798 1091 4833 1125
rect 4867 1091 4902 1125
rect 4936 1091 4971 1125
rect 5005 1091 5040 1125
rect 5074 1091 5109 1125
rect 5143 1091 5178 1125
rect 5212 1091 5247 1125
rect 5281 1091 5316 1125
rect 5350 1091 5385 1125
rect 5419 1091 5454 1125
rect 5488 1091 5523 1125
rect 14397 1253 14493 1278
rect 14397 1219 14455 1253
rect 14489 1244 14493 1253
rect 14527 1249 14566 1278
rect 14625 1252 14639 1278
rect 14557 1244 14566 1249
rect 14600 1244 14639 1252
rect 14673 1244 14701 1278
rect 14489 1219 14523 1244
rect 14397 1215 14523 1219
rect 14557 1216 14701 1244
rect 14557 1215 14591 1216
rect 14397 1206 14591 1215
rect 14625 1206 14701 1216
rect 14397 1181 14493 1206
rect 14397 1147 14455 1181
rect 14489 1172 14493 1181
rect 14527 1179 14566 1206
rect 14625 1182 14639 1206
rect 14557 1172 14566 1179
rect 14600 1172 14639 1182
rect 14673 1172 14701 1206
rect 23040 1483 23048 1494
rect 23082 1483 23117 1517
rect 23151 1483 23186 1517
rect 23220 1483 23255 1517
rect 23289 1483 23324 1517
rect 23358 1483 23393 1517
rect 23427 1483 23462 1517
rect 23496 1483 23531 1517
rect 23565 1483 23600 1517
rect 23634 1483 23669 1517
rect 23703 1483 23738 1517
rect 23772 1483 23796 1517
rect 23040 1449 23796 1483
rect 23040 1415 23048 1449
rect 23082 1415 23117 1449
rect 23151 1415 23186 1449
rect 23220 1415 23255 1449
rect 23289 1415 23324 1449
rect 23358 1415 23393 1449
rect 23427 1415 23462 1449
rect 23496 1415 23531 1449
rect 23565 1415 23600 1449
rect 23634 1415 23669 1449
rect 23703 1415 23738 1449
rect 23772 1415 23796 1449
rect 23040 1381 23796 1415
rect 23040 1347 23048 1381
rect 23082 1347 23117 1381
rect 23151 1347 23186 1381
rect 23220 1347 23255 1381
rect 23289 1347 23324 1381
rect 23358 1347 23393 1381
rect 23427 1347 23462 1381
rect 23496 1347 23531 1381
rect 23565 1347 23600 1381
rect 23634 1347 23669 1381
rect 23703 1347 23738 1381
rect 23772 1347 23796 1381
rect 23040 1313 23796 1347
rect 23040 1279 23048 1313
rect 23082 1279 23117 1313
rect 23151 1279 23186 1313
rect 23220 1279 23255 1313
rect 23289 1279 23324 1313
rect 23358 1279 23393 1313
rect 23427 1279 23462 1313
rect 23496 1279 23531 1313
rect 23565 1279 23600 1313
rect 23634 1279 23669 1313
rect 23703 1279 23738 1313
rect 23772 1279 23796 1313
rect 23040 1245 23796 1279
rect 23040 1211 23048 1245
rect 23082 1211 23117 1245
rect 23151 1211 23186 1245
rect 23220 1211 23255 1245
rect 23289 1211 23324 1245
rect 23358 1211 23393 1245
rect 23427 1211 23462 1245
rect 23496 1211 23531 1245
rect 23565 1211 23600 1245
rect 23634 1211 23669 1245
rect 23703 1211 23738 1245
rect 23772 1211 23796 1245
rect 23040 1177 23796 1211
rect 23040 1172 23048 1177
rect 14489 1147 14523 1172
rect 14397 1145 14523 1147
rect 14557 1146 14701 1172
rect 14557 1145 14591 1146
rect 14397 1134 14591 1145
rect 14625 1143 14701 1146
rect 19563 1143 19598 1172
rect 19632 1143 19667 1172
rect 19701 1143 19736 1172
rect 19770 1143 19805 1172
rect 19839 1143 19874 1172
rect 19908 1143 19943 1172
rect 19977 1143 20012 1172
rect 20046 1143 20081 1172
rect 20115 1143 20150 1172
rect 20184 1143 20219 1172
rect 20253 1143 20288 1172
rect 20322 1143 20357 1172
rect 20391 1143 20426 1172
rect 20460 1143 20495 1172
rect 20529 1143 20564 1172
rect 20598 1143 20633 1172
rect 20667 1143 20702 1172
rect 20736 1143 20771 1172
rect 20805 1143 20840 1172
rect 20874 1143 20909 1172
rect 20943 1143 20978 1172
rect 21012 1143 21047 1172
rect 21081 1143 21116 1172
rect 21150 1143 21185 1172
rect 21219 1143 21254 1172
rect 21288 1143 21323 1172
rect 21357 1143 21392 1172
rect 21426 1143 21461 1172
rect 21495 1143 21530 1172
rect 21564 1143 21599 1172
rect 21633 1143 21668 1172
rect 21702 1143 21737 1172
rect 21771 1143 21806 1172
rect 21840 1143 21875 1172
rect 21909 1143 21944 1172
rect 21978 1143 22013 1172
rect 22047 1143 22082 1172
rect 22116 1143 22151 1172
rect 22185 1143 22220 1172
rect 22254 1143 22289 1172
rect 22323 1143 22358 1172
rect 22392 1143 22427 1172
rect 22461 1143 22496 1172
rect 22530 1143 22565 1172
rect 22599 1143 22634 1172
rect 22668 1143 22703 1172
rect 22737 1143 22772 1172
rect 22806 1143 22841 1172
rect 22875 1143 22910 1172
rect 22944 1143 22979 1172
rect 23013 1143 23048 1172
rect 23082 1143 23117 1177
rect 23151 1143 23186 1177
rect 23220 1143 23255 1177
rect 23289 1143 23324 1177
rect 23358 1143 23393 1177
rect 23427 1143 23462 1177
rect 23496 1143 23531 1177
rect 23565 1143 23600 1177
rect 23634 1143 23669 1177
rect 23703 1143 23738 1177
rect 23772 1143 23796 1177
rect 14397 1109 14487 1134
rect 14521 1109 14559 1134
rect 14625 1128 23796 1143
rect 24119 5522 24540 5532
rect 24119 5488 24153 5522
rect 24187 5488 24221 5522
rect 24255 5488 24289 5522
rect 24323 5488 24357 5522
rect 24391 5488 24425 5522
rect 24459 5488 24493 5522
rect 24527 5488 24540 5522
rect 24119 5453 24540 5488
rect 24119 5419 24153 5453
rect 24187 5419 24221 5453
rect 24255 5419 24289 5453
rect 24323 5419 24357 5453
rect 24391 5419 24425 5453
rect 24459 5419 24493 5453
rect 24527 5419 24540 5453
rect 24119 5384 24540 5419
rect 24119 5350 24153 5384
rect 24187 5350 24221 5384
rect 24255 5350 24289 5384
rect 24323 5350 24357 5384
rect 24391 5350 24425 5384
rect 24459 5350 24493 5384
rect 24527 5350 24540 5384
rect 24119 5315 24540 5350
rect 24119 5281 24153 5315
rect 24187 5281 24221 5315
rect 24255 5281 24289 5315
rect 24323 5281 24357 5315
rect 24391 5281 24425 5315
rect 24459 5281 24493 5315
rect 24527 5281 24540 5315
rect 24119 5246 24540 5281
rect 24119 5212 24153 5246
rect 24187 5212 24221 5246
rect 24255 5212 24289 5246
rect 24323 5212 24357 5246
rect 24391 5212 24425 5246
rect 24459 5212 24493 5246
rect 24527 5212 24540 5246
rect 24119 5177 24540 5212
rect 24119 5143 24153 5177
rect 24187 5143 24221 5177
rect 24255 5143 24289 5177
rect 24323 5143 24357 5177
rect 24391 5143 24425 5177
rect 24459 5143 24493 5177
rect 24527 5143 24540 5177
rect 24119 5108 24540 5143
rect 24119 5074 24153 5108
rect 24187 5074 24221 5108
rect 24255 5074 24289 5108
rect 24323 5074 24357 5108
rect 24391 5074 24425 5108
rect 24459 5074 24493 5108
rect 24527 5074 24540 5108
rect 24119 5039 24540 5074
rect 24119 5005 24153 5039
rect 24187 5005 24221 5039
rect 24255 5005 24289 5039
rect 24323 5005 24357 5039
rect 24391 5005 24425 5039
rect 24459 5005 24493 5039
rect 24527 5005 24540 5039
rect 24119 4970 24540 5005
rect 24119 4936 24153 4970
rect 24187 4936 24221 4970
rect 24255 4936 24289 4970
rect 24323 4936 24357 4970
rect 24391 4936 24425 4970
rect 24459 4936 24493 4970
rect 24527 4936 24540 4970
rect 24119 4901 24540 4936
rect 24119 4867 24153 4901
rect 24187 4867 24221 4901
rect 24255 4867 24289 4901
rect 24323 4867 24357 4901
rect 24391 4867 24425 4901
rect 24459 4867 24493 4901
rect 24527 4867 24540 4901
rect 24119 4832 24540 4867
rect 24119 4798 24153 4832
rect 24187 4798 24221 4832
rect 24255 4798 24289 4832
rect 24323 4798 24357 4832
rect 24391 4798 24425 4832
rect 24459 4798 24493 4832
rect 24527 4798 24540 4832
rect 24119 4763 24540 4798
rect 24119 4729 24153 4763
rect 24187 4729 24221 4763
rect 24255 4729 24289 4763
rect 24323 4729 24357 4763
rect 24391 4729 24425 4763
rect 24459 4729 24493 4763
rect 24527 4729 24540 4763
rect 24119 4694 24540 4729
rect 24527 2348 24540 4694
rect 24119 2324 24540 2348
rect 14397 1091 14455 1109
rect 14521 1100 14523 1109
rect 696 1074 764 1081
rect 730 1043 764 1074
rect 866 1075 14455 1091
rect 14489 1075 14523 1100
rect 14557 1100 14559 1109
rect 14593 1100 14625 1112
rect 14557 1076 14625 1100
rect 14557 1075 14591 1076
rect 866 1053 14591 1075
rect 696 1009 728 1040
rect 762 1009 764 1043
rect 696 1005 764 1009
rect 866 1039 14559 1053
rect 866 1037 14523 1039
rect 866 1005 901 1037
rect 935 1005 970 1037
rect 1004 1005 1039 1037
rect 1073 1005 1108 1037
rect 1142 1005 1177 1037
rect 1211 1005 1246 1037
rect 1280 1005 1315 1037
rect 1349 1005 1384 1037
rect 1418 1005 1453 1037
rect 1487 1005 1522 1037
rect 1556 1005 1591 1037
rect 1625 1005 1660 1037
rect 1694 1005 1729 1037
rect 1763 1005 1798 1037
rect 1832 1005 1867 1037
rect 1901 1005 1936 1037
rect 1970 1005 2005 1037
rect 2039 1005 2074 1037
rect 2108 1005 2143 1037
rect 2177 1005 2212 1037
rect 2246 1005 2281 1037
rect 2315 1005 2350 1037
rect 2384 1005 2419 1037
rect 14489 1005 14523 1037
rect 14557 1019 14559 1039
rect 14593 1019 14625 1042
rect 14557 1006 14625 1019
rect 14557 1005 14591 1006
rect 730 1003 764 1005
rect 866 1003 873 1005
rect 935 1003 946 1005
rect 1004 1003 1019 1005
rect 1073 1003 1092 1005
rect 1142 1003 1165 1005
rect 1211 1003 1238 1005
rect 1280 1003 1311 1005
rect 730 971 800 1003
rect 834 971 873 1003
rect 907 971 946 1003
rect 980 971 1019 1003
rect 1053 971 1092 1003
rect 1126 971 1165 1003
rect 1199 971 1238 1003
rect 1272 971 1311 1003
rect 696 969 1311 971
rect 14521 972 14591 1005
rect 14521 971 14625 972
rect 14489 969 14559 971
rect 696 935 764 969
rect 798 935 833 969
rect 867 935 902 969
rect 936 935 971 969
rect 1005 935 1040 969
rect 1074 935 1109 969
rect 1143 935 1178 969
rect 1212 935 1247 969
rect 1281 935 1311 969
rect 696 933 1311 935
rect 696 901 766 933
rect 800 901 839 933
rect 873 901 912 933
rect 946 901 985 933
rect 1019 901 1057 933
rect 1091 901 1129 933
rect 1163 901 1201 933
rect 1235 901 1273 933
rect 1307 901 1311 933
rect 14557 937 14559 969
rect 14593 937 14625 971
rect 14557 935 14625 937
rect 696 867 730 901
rect 764 899 766 901
rect 833 899 839 901
rect 902 899 912 901
rect 971 899 985 901
rect 1040 899 1057 901
rect 1109 899 1129 901
rect 1178 899 1201 901
rect 1247 899 1273 901
rect 14523 901 14591 935
rect 764 867 799 899
rect 833 867 868 899
rect 902 867 937 899
rect 971 867 1006 899
rect 1040 867 1075 899
rect 1109 867 1144 899
rect 1178 867 1213 899
rect 1247 867 1282 899
rect 1316 867 1351 899
rect 1385 867 1420 899
rect 1454 867 1489 899
rect 1523 867 1558 899
rect 1592 867 1627 899
rect 1661 867 1696 899
rect 1730 867 1765 899
rect 1799 867 1834 899
rect 1868 867 1903 899
rect 1937 867 1972 899
rect 2006 867 2041 899
rect 2075 867 2110 899
rect 2144 867 2179 899
rect 2213 867 2248 899
rect 2282 867 2317 899
rect 14523 867 14625 901
rect 20507 944 20558 976
rect 20592 944 20627 976
rect 20507 910 20551 944
rect 20592 942 20625 944
rect 20661 942 20696 976
rect 20730 944 20765 976
rect 20799 944 20834 976
rect 20868 944 20903 976
rect 20937 944 20972 976
rect 21006 944 21041 976
rect 21075 944 21110 976
rect 21144 944 21179 976
rect 20733 942 20765 944
rect 20807 942 20834 944
rect 20881 942 20903 944
rect 20955 942 20972 944
rect 21029 942 21041 944
rect 21103 942 21110 944
rect 21177 942 21179 944
rect 21213 944 21248 976
rect 21282 944 21317 976
rect 21351 944 21386 976
rect 21420 944 21455 976
rect 21489 944 21524 976
rect 21558 944 21593 976
rect 21627 944 21662 976
rect 21213 942 21217 944
rect 21282 942 21291 944
rect 21351 942 21365 944
rect 21420 942 21439 944
rect 21489 942 21513 944
rect 21558 942 21587 944
rect 21627 942 21661 944
rect 21696 942 21731 976
rect 21765 944 21800 976
rect 21834 944 21869 976
rect 21903 944 21938 976
rect 21972 944 22007 976
rect 22041 944 22076 976
rect 22110 944 22145 976
rect 21769 942 21800 944
rect 21843 942 21869 944
rect 21917 942 21938 944
rect 21991 942 22007 944
rect 22065 942 22076 944
rect 22139 942 22145 944
rect 22179 944 22214 976
rect 20585 910 20625 942
rect 20659 910 20699 942
rect 20733 910 20773 942
rect 20807 910 20847 942
rect 20881 910 20921 942
rect 20955 910 20995 942
rect 21029 910 21069 942
rect 21103 910 21143 942
rect 21177 910 21217 942
rect 21251 910 21291 942
rect 21325 910 21365 942
rect 21399 910 21439 942
rect 21473 910 21513 942
rect 21547 910 21587 942
rect 21621 910 21661 942
rect 21695 910 21735 942
rect 21769 910 21809 942
rect 21843 910 21883 942
rect 21917 910 21957 942
rect 21991 910 22031 942
rect 22065 910 22105 942
rect 22139 910 22179 942
rect 22213 942 22214 944
rect 22248 944 22283 976
rect 22317 944 22352 976
rect 22386 944 22421 976
rect 22455 944 22490 976
rect 22524 944 22559 976
rect 22593 944 22628 976
rect 22662 944 22697 976
rect 22248 942 22253 944
rect 22317 942 22327 944
rect 22386 942 22401 944
rect 22455 942 22475 944
rect 22524 942 22549 944
rect 22593 942 22622 944
rect 22662 942 22695 944
rect 22731 942 22766 976
rect 22800 944 22835 976
rect 22869 944 22904 976
rect 22938 944 22973 976
rect 22802 942 22835 944
rect 22875 942 22904 944
rect 22213 910 22253 942
rect 22287 910 22327 942
rect 22361 910 22401 942
rect 22435 910 22475 942
rect 22509 910 22549 942
rect 22583 910 22622 942
rect 22656 910 22695 942
rect 22729 910 22768 942
rect 22802 910 22841 942
rect 22875 910 22914 942
rect 22948 910 22973 944
rect 20507 908 22973 910
rect 20507 874 20558 908
rect 20592 874 20627 908
rect 20661 874 20696 908
rect 20730 874 20765 908
rect 20799 874 20834 908
rect 20868 874 20903 908
rect 20937 874 20972 908
rect 21006 874 21041 908
rect 21075 874 21110 908
rect 21144 874 21179 908
rect 21213 874 21248 908
rect 21282 874 21317 908
rect 21351 874 21386 908
rect 21420 874 21455 908
rect 21489 874 21524 908
rect 21558 874 21593 908
rect 21627 874 21662 908
rect 21696 874 21731 908
rect 21765 874 21800 908
rect 21834 874 21869 908
rect 21903 874 21938 908
rect 21972 874 22007 908
rect 22041 874 22076 908
rect 22110 874 22145 908
rect 22179 874 22214 908
rect 22248 874 22283 908
rect 22317 874 22352 908
rect 22386 874 22421 908
rect 22455 874 22490 908
rect 22524 874 22559 908
rect 22593 874 22628 908
rect 22662 874 22697 908
rect 22731 874 22766 908
rect 22800 874 22835 908
rect 22869 874 22904 908
rect 22938 874 22973 908
rect 20507 872 22973 874
rect 278 855 448 857
rect 278 822 310 855
rect 344 822 382 855
rect 416 822 448 855
rect 344 821 346 822
rect 312 788 346 821
rect 380 821 382 822
rect 380 788 414 821
rect 20507 838 20551 872
rect 20585 840 20625 872
rect 20659 840 20699 872
rect 20733 840 20773 872
rect 20807 840 20847 872
rect 20881 840 20921 872
rect 20955 840 20995 872
rect 21029 840 21069 872
rect 21103 840 21143 872
rect 21177 840 21217 872
rect 21251 840 21291 872
rect 21325 840 21365 872
rect 21399 840 21439 872
rect 21473 840 21513 872
rect 21547 840 21587 872
rect 21621 840 21661 872
rect 21695 840 21735 872
rect 21769 840 21809 872
rect 21843 840 21883 872
rect 21917 840 21957 872
rect 21991 840 22031 872
rect 22065 840 22105 872
rect 22139 840 22179 872
rect 20592 838 20625 840
rect 20507 806 20558 838
rect 20592 806 20627 838
rect 20661 806 20696 840
rect 20733 838 20765 840
rect 20807 838 20834 840
rect 20881 838 20903 840
rect 20955 838 20972 840
rect 21029 838 21041 840
rect 21103 838 21110 840
rect 21177 838 21179 840
rect 20730 806 20765 838
rect 20799 806 20834 838
rect 20868 806 20903 838
rect 20937 806 20972 838
rect 21006 806 21041 838
rect 21075 806 21110 838
rect 21144 806 21179 838
rect 21213 838 21217 840
rect 21282 838 21291 840
rect 21351 838 21365 840
rect 21420 838 21439 840
rect 21489 838 21513 840
rect 21558 838 21587 840
rect 21627 838 21661 840
rect 21213 806 21248 838
rect 21282 806 21317 838
rect 21351 806 21386 838
rect 21420 806 21455 838
rect 21489 806 21524 838
rect 21558 806 21593 838
rect 21627 806 21662 838
rect 21696 806 21731 840
rect 21769 838 21800 840
rect 21843 838 21869 840
rect 21917 838 21938 840
rect 21991 838 22007 840
rect 22065 838 22076 840
rect 22139 838 22145 840
rect 21765 806 21800 838
rect 21834 806 21869 838
rect 21903 806 21938 838
rect 21972 806 22007 838
rect 22041 806 22076 838
rect 22110 806 22145 838
rect 22213 840 22253 872
rect 22287 840 22327 872
rect 22361 840 22401 872
rect 22435 840 22475 872
rect 22509 840 22549 872
rect 22583 840 22622 872
rect 22656 840 22695 872
rect 22729 840 22768 872
rect 22802 840 22841 872
rect 22875 840 22914 872
rect 22213 838 22214 840
rect 22179 806 22214 838
rect 22248 838 22253 840
rect 22317 838 22327 840
rect 22386 838 22401 840
rect 22455 838 22475 840
rect 22524 838 22549 840
rect 22593 838 22622 840
rect 22662 838 22695 840
rect 22248 806 22283 838
rect 22317 806 22352 838
rect 22386 806 22421 838
rect 22455 806 22490 838
rect 22524 806 22559 838
rect 22593 806 22628 838
rect 22662 806 22697 838
rect 22731 806 22766 840
rect 22802 838 22835 840
rect 22875 838 22904 840
rect 22948 838 22973 872
rect 22800 806 22835 838
rect 22869 806 22904 838
rect 22938 806 22973 838
rect 24095 806 24119 1010
rect 278 782 448 788
rect 278 753 310 782
rect 344 753 382 782
rect 416 753 448 782
rect 24272 772 24306 854
rect 25862 772 25896 854
rect 344 748 346 753
rect 312 719 346 748
rect 380 748 382 753
rect 380 719 414 748
rect 278 709 448 719
rect 278 684 310 709
rect 344 684 382 709
rect 416 684 448 709
rect 344 675 346 684
rect 312 650 346 675
rect 380 675 382 684
rect 380 650 414 675
rect 278 636 448 650
rect 278 615 310 636
rect 344 615 382 636
rect 416 615 448 636
rect 344 602 346 615
rect 312 581 346 602
rect 380 602 382 615
rect 380 581 414 602
rect 278 563 448 581
rect 278 546 310 563
rect 344 546 382 563
rect 416 546 448 563
rect 344 529 346 546
rect 312 512 346 529
rect 380 529 382 546
rect 380 512 414 529
rect 278 490 448 512
rect 278 477 310 490
rect 344 477 382 490
rect 416 477 448 490
rect 344 456 346 477
rect 312 443 346 456
rect 380 456 382 477
rect 380 443 414 456
rect 278 417 448 443
rect 278 408 310 417
rect 344 408 382 417
rect 416 408 448 417
rect 344 383 346 408
rect 312 374 346 383
rect 380 383 382 408
rect 380 374 414 383
rect 278 344 448 374
rect 278 339 310 344
rect 344 339 382 344
rect 416 339 448 344
rect 344 310 346 339
rect 312 305 346 310
rect 380 310 382 339
rect 380 305 414 310
rect 278 271 448 305
rect 278 270 310 271
rect 344 270 382 271
rect 416 270 448 271
rect 344 237 346 270
rect 312 236 346 237
rect 380 237 382 270
rect 380 236 414 237
rect 278 201 448 236
rect 312 198 346 201
rect 344 167 346 198
rect 380 198 414 201
rect 380 167 382 198
rect 278 164 310 167
rect 344 164 382 167
rect 416 164 448 167
rect 278 133 448 164
rect 21231 -1923 21269 -1889
rect 21303 -1923 21341 -1889
rect 21375 -1923 21413 -1889
rect 21447 -1923 21485 -1889
rect 21197 -1929 21519 -1923
<< viali >>
rect 22798 8985 22818 8997
rect 22818 8985 22852 8997
rect 22852 8985 22886 8997
rect 22886 8985 22920 8997
rect 22920 8985 22954 8997
rect 22954 8985 22988 8997
rect 22988 8985 23022 8997
rect 23022 8985 23056 8997
rect 23056 8985 23090 8997
rect 23090 8985 23124 8997
rect 23124 8985 23158 8997
rect 23158 8985 23192 8997
rect 23192 8985 23226 8997
rect 23226 8985 23260 8997
rect 23260 8985 23294 8997
rect 23294 8985 23328 8997
rect 23328 8985 23362 8997
rect 23362 8985 23396 8997
rect 23396 8985 23430 8997
rect 23430 8985 23464 8997
rect 23464 8985 23480 8997
rect 22798 8950 23480 8985
rect 22798 8916 22818 8950
rect 22818 8916 22852 8950
rect 22852 8916 22886 8950
rect 22886 8916 22920 8950
rect 22920 8916 22954 8950
rect 22954 8916 22988 8950
rect 22988 8916 23022 8950
rect 23022 8916 23056 8950
rect 23056 8916 23090 8950
rect 23090 8916 23124 8950
rect 23124 8916 23158 8950
rect 23158 8916 23192 8950
rect 23192 8916 23226 8950
rect 23226 8916 23260 8950
rect 23260 8916 23294 8950
rect 23294 8916 23328 8950
rect 23328 8916 23362 8950
rect 23362 8916 23396 8950
rect 23396 8916 23430 8950
rect 23430 8916 23464 8950
rect 23464 8916 23480 8950
rect 22798 8881 23480 8916
rect 22798 8847 22818 8881
rect 22818 8847 22852 8881
rect 22852 8847 22886 8881
rect 22886 8847 22920 8881
rect 22920 8847 22954 8881
rect 22954 8847 22988 8881
rect 22988 8847 23022 8881
rect 23022 8847 23056 8881
rect 23056 8847 23090 8881
rect 23090 8847 23124 8881
rect 23124 8847 23158 8881
rect 23158 8847 23192 8881
rect 23192 8847 23226 8881
rect 23226 8847 23260 8881
rect 23260 8847 23294 8881
rect 23294 8847 23328 8881
rect 23328 8847 23362 8881
rect 23362 8847 23396 8881
rect 23396 8847 23430 8881
rect 23430 8847 23464 8881
rect 23464 8847 23480 8881
rect 22798 8812 23480 8847
rect 22798 8778 22818 8812
rect 22818 8778 22852 8812
rect 22852 8778 22886 8812
rect 22886 8778 22920 8812
rect 22920 8778 22954 8812
rect 22954 8778 22988 8812
rect 22988 8778 23022 8812
rect 23022 8778 23056 8812
rect 23056 8778 23090 8812
rect 23090 8778 23124 8812
rect 23124 8778 23158 8812
rect 23158 8778 23192 8812
rect 23192 8778 23226 8812
rect 23226 8778 23260 8812
rect 23260 8778 23294 8812
rect 23294 8778 23328 8812
rect 23328 8778 23362 8812
rect 23362 8778 23396 8812
rect 23396 8778 23430 8812
rect 23430 8778 23464 8812
rect 23464 8778 23480 8812
rect 22798 8743 23480 8778
rect 22798 8709 22818 8743
rect 22818 8709 22852 8743
rect 22852 8709 22886 8743
rect 22886 8709 22920 8743
rect 22920 8709 22954 8743
rect 22954 8709 22988 8743
rect 22988 8709 23022 8743
rect 23022 8709 23056 8743
rect 23056 8709 23090 8743
rect 23090 8709 23124 8743
rect 23124 8709 23158 8743
rect 23158 8709 23192 8743
rect 23192 8709 23226 8743
rect 23226 8709 23260 8743
rect 23260 8709 23294 8743
rect 23294 8709 23328 8743
rect 23328 8709 23362 8743
rect 23362 8709 23396 8743
rect 23396 8709 23430 8743
rect 23430 8709 23464 8743
rect 23464 8709 23480 8743
rect 22798 8674 23480 8709
rect 22798 8640 22818 8674
rect 22818 8640 22852 8674
rect 22852 8640 22886 8674
rect 22886 8640 22920 8674
rect 22920 8640 22954 8674
rect 22954 8640 22988 8674
rect 22988 8640 23022 8674
rect 23022 8640 23056 8674
rect 23056 8640 23090 8674
rect 23090 8640 23124 8674
rect 23124 8640 23158 8674
rect 23158 8640 23192 8674
rect 23192 8640 23226 8674
rect 23226 8640 23260 8674
rect 23260 8640 23294 8674
rect 23294 8640 23328 8674
rect 23328 8640 23362 8674
rect 23362 8640 23396 8674
rect 23396 8640 23430 8674
rect 23430 8640 23464 8674
rect 23464 8640 23480 8674
rect 22798 8605 23480 8640
rect 22798 8603 22818 8605
rect 22818 8603 22852 8605
rect 22852 8603 22886 8605
rect 22886 8603 22920 8605
rect 22920 8603 22954 8605
rect 22954 8603 22988 8605
rect 22988 8603 23022 8605
rect 23022 8603 23056 8605
rect 23056 8603 23090 8605
rect 23090 8603 23124 8605
rect 23124 8603 23158 8605
rect 23158 8603 23192 8605
rect 23192 8603 23226 8605
rect 23226 8603 23260 8605
rect 23260 8603 23294 8605
rect 23294 8603 23328 8605
rect 23328 8603 23362 8605
rect 23362 8603 23396 8605
rect 23396 8603 23430 8605
rect 23430 8603 23464 8605
rect 23464 8603 23480 8605
rect 23781 8671 24370 8680
rect 24370 8671 24404 8680
rect 24404 8671 24438 8680
rect 24438 8671 24472 8680
rect 24472 8671 24506 8680
rect 24506 8671 24535 8680
rect 23781 8636 24535 8671
rect 22798 8536 22832 8564
rect 22870 8536 22904 8564
rect 22942 8536 22976 8564
rect 23014 8536 23048 8564
rect 23086 8536 23120 8564
rect 23158 8536 23192 8564
rect 23230 8536 23264 8564
rect 23302 8536 23336 8564
rect 23374 8536 23408 8564
rect 23446 8536 23480 8564
rect 22798 8530 22818 8536
rect 22818 8530 22832 8536
rect 22870 8530 22886 8536
rect 22886 8530 22904 8536
rect 22942 8530 22954 8536
rect 22954 8530 22976 8536
rect 23014 8530 23022 8536
rect 23022 8530 23048 8536
rect 23086 8530 23090 8536
rect 23090 8530 23120 8536
rect 23158 8530 23192 8536
rect 23230 8530 23260 8536
rect 23260 8530 23264 8536
rect 23302 8530 23328 8536
rect 23328 8530 23336 8536
rect 23374 8530 23396 8536
rect 23396 8530 23408 8536
rect 23446 8530 23464 8536
rect 23464 8530 23480 8536
rect 22798 8467 22832 8491
rect 22870 8467 22904 8491
rect 22942 8467 22976 8491
rect 23014 8467 23048 8491
rect 23086 8467 23120 8491
rect 23158 8467 23192 8491
rect 23230 8467 23264 8491
rect 23302 8467 23336 8491
rect 23374 8467 23408 8491
rect 23446 8467 23480 8491
rect 22798 8457 22818 8467
rect 22818 8457 22832 8467
rect 22870 8457 22886 8467
rect 22886 8457 22904 8467
rect 22942 8457 22954 8467
rect 22954 8457 22976 8467
rect 23014 8457 23022 8467
rect 23022 8457 23048 8467
rect 23086 8457 23090 8467
rect 23090 8457 23120 8467
rect 23158 8457 23192 8467
rect 23230 8457 23260 8467
rect 23260 8457 23264 8467
rect 23302 8457 23328 8467
rect 23328 8457 23336 8467
rect 23374 8457 23396 8467
rect 23396 8457 23408 8467
rect 23446 8457 23464 8467
rect 23464 8457 23480 8467
rect 22798 8398 22832 8418
rect 22870 8398 22904 8418
rect 22942 8398 22976 8418
rect 23014 8398 23048 8418
rect 23086 8398 23120 8418
rect 23158 8398 23192 8418
rect 23230 8398 23264 8418
rect 23302 8398 23336 8418
rect 23374 8398 23408 8418
rect 23446 8398 23480 8418
rect 22798 8384 22818 8398
rect 22818 8384 22832 8398
rect 22870 8384 22886 8398
rect 22886 8384 22904 8398
rect 22942 8384 22954 8398
rect 22954 8384 22976 8398
rect 23014 8384 23022 8398
rect 23022 8384 23048 8398
rect 23086 8384 23090 8398
rect 23090 8384 23120 8398
rect 23158 8384 23192 8398
rect 23230 8384 23260 8398
rect 23260 8384 23264 8398
rect 23302 8384 23328 8398
rect 23328 8384 23336 8398
rect 23374 8384 23396 8398
rect 23396 8384 23408 8398
rect 23446 8384 23464 8398
rect 23464 8384 23480 8398
rect 22798 8329 22832 8345
rect 22870 8329 22904 8345
rect 22942 8329 22976 8345
rect 23014 8329 23048 8345
rect 23086 8329 23120 8345
rect 23158 8329 23192 8345
rect 23230 8329 23264 8345
rect 23302 8329 23336 8345
rect 23374 8329 23408 8345
rect 23446 8329 23480 8345
rect 22798 8311 22818 8329
rect 22818 8311 22832 8329
rect 22870 8311 22886 8329
rect 22886 8311 22904 8329
rect 22942 8311 22954 8329
rect 22954 8311 22976 8329
rect 23014 8311 23022 8329
rect 23022 8311 23048 8329
rect 23086 8311 23090 8329
rect 23090 8311 23120 8329
rect 23158 8311 23192 8329
rect 23230 8311 23260 8329
rect 23260 8311 23264 8329
rect 23302 8311 23328 8329
rect 23328 8311 23336 8329
rect 23374 8311 23396 8329
rect 23396 8311 23408 8329
rect 23446 8311 23464 8329
rect 23464 8311 23480 8329
rect 22798 8260 22832 8272
rect 22870 8260 22904 8272
rect 22942 8260 22976 8272
rect 23014 8260 23048 8272
rect 23086 8260 23120 8272
rect 23158 8260 23192 8272
rect 23230 8260 23264 8272
rect 23302 8260 23336 8272
rect 23374 8260 23408 8272
rect 23446 8260 23480 8272
rect 22798 8238 22818 8260
rect 22818 8238 22832 8260
rect 22870 8238 22886 8260
rect 22886 8238 22904 8260
rect 22942 8238 22954 8260
rect 22954 8238 22976 8260
rect 23014 8238 23022 8260
rect 23022 8238 23048 8260
rect 23086 8238 23090 8260
rect 23090 8238 23120 8260
rect 23158 8238 23192 8260
rect 23230 8238 23260 8260
rect 23260 8238 23264 8260
rect 23302 8238 23328 8260
rect 23328 8238 23336 8260
rect 23374 8238 23396 8260
rect 23396 8238 23408 8260
rect 23446 8238 23464 8260
rect 23464 8238 23480 8260
rect 22798 8191 22832 8199
rect 22870 8191 22904 8199
rect 22942 8191 22976 8199
rect 23014 8191 23048 8199
rect 23086 8191 23120 8199
rect 23158 8191 23192 8199
rect 23230 8191 23264 8199
rect 23302 8191 23336 8199
rect 23374 8191 23408 8199
rect 23446 8191 23480 8199
rect 22798 8165 22818 8191
rect 22818 8165 22832 8191
rect 22870 8165 22886 8191
rect 22886 8165 22904 8191
rect 22942 8165 22954 8191
rect 22954 8165 22976 8191
rect 23014 8165 23022 8191
rect 23022 8165 23048 8191
rect 23086 8165 23090 8191
rect 23090 8165 23120 8191
rect 23158 8165 23192 8191
rect 23230 8165 23260 8191
rect 23260 8165 23264 8191
rect 23302 8165 23328 8191
rect 23328 8165 23336 8191
rect 23374 8165 23396 8191
rect 23396 8165 23408 8191
rect 23446 8165 23464 8191
rect 23464 8165 23480 8191
rect 22798 8122 22832 8126
rect 22870 8122 22904 8126
rect 22942 8122 22976 8126
rect 23014 8122 23048 8126
rect 23086 8122 23120 8126
rect 23158 8122 23192 8126
rect 23230 8122 23264 8126
rect 23302 8122 23336 8126
rect 23374 8122 23408 8126
rect 23446 8122 23480 8126
rect 22798 8092 22818 8122
rect 22818 8092 22832 8122
rect 22870 8092 22886 8122
rect 22886 8092 22904 8122
rect 22942 8092 22954 8122
rect 22954 8092 22976 8122
rect 23014 8092 23022 8122
rect 23022 8092 23048 8122
rect 23086 8092 23090 8122
rect 23090 8092 23120 8122
rect 23158 8092 23192 8122
rect 23230 8092 23260 8122
rect 23260 8092 23264 8122
rect 23302 8092 23328 8122
rect 23328 8092 23336 8122
rect 23374 8092 23396 8122
rect 23396 8092 23408 8122
rect 23446 8092 23464 8122
rect 23464 8092 23480 8122
rect 22798 8019 22818 8053
rect 22818 8019 22832 8053
rect 22870 8019 22886 8053
rect 22886 8019 22904 8053
rect 22942 8019 22954 8053
rect 22954 8019 22976 8053
rect 23014 8019 23022 8053
rect 23022 8019 23048 8053
rect 23086 8019 23090 8053
rect 23090 8019 23120 8053
rect 23158 8019 23192 8053
rect 23230 8019 23260 8053
rect 23260 8019 23264 8053
rect 23302 8019 23328 8053
rect 23328 8019 23336 8053
rect 23374 8019 23396 8053
rect 23396 8019 23408 8053
rect 23446 8019 23464 8053
rect 23464 8019 23480 8053
rect 22798 7950 22818 7980
rect 22818 7950 22832 7980
rect 22870 7950 22886 7980
rect 22886 7950 22904 7980
rect 22942 7950 22954 7980
rect 22954 7950 22976 7980
rect 23014 7950 23022 7980
rect 23022 7950 23048 7980
rect 23086 7950 23090 7980
rect 23090 7950 23120 7980
rect 23158 7950 23192 7980
rect 23230 7950 23260 7980
rect 23260 7950 23264 7980
rect 23302 7950 23328 7980
rect 23328 7950 23336 7980
rect 23374 7950 23396 7980
rect 23396 7950 23408 7980
rect 23446 7950 23464 7980
rect 23464 7950 23480 7980
rect 22798 7946 22832 7950
rect 22870 7946 22904 7950
rect 22942 7946 22976 7950
rect 23014 7946 23048 7950
rect 23086 7946 23120 7950
rect 23158 7946 23192 7950
rect 23230 7946 23264 7950
rect 23302 7946 23336 7950
rect 23374 7946 23408 7950
rect 23446 7946 23480 7950
rect 22798 7881 22818 7907
rect 22818 7881 22832 7907
rect 22870 7881 22886 7907
rect 22886 7881 22904 7907
rect 22942 7881 22954 7907
rect 22954 7881 22976 7907
rect 23014 7881 23022 7907
rect 23022 7881 23048 7907
rect 23086 7881 23090 7907
rect 23090 7881 23120 7907
rect 23158 7881 23192 7907
rect 23230 7881 23260 7907
rect 23260 7881 23264 7907
rect 23302 7881 23328 7907
rect 23328 7881 23336 7907
rect 23374 7881 23396 7907
rect 23396 7881 23408 7907
rect 23446 7881 23464 7907
rect 23464 7881 23480 7907
rect 22798 7873 22832 7881
rect 22870 7873 22904 7881
rect 22942 7873 22976 7881
rect 23014 7873 23048 7881
rect 23086 7873 23120 7881
rect 23158 7873 23192 7881
rect 23230 7873 23264 7881
rect 23302 7873 23336 7881
rect 23374 7873 23408 7881
rect 23446 7873 23480 7881
rect 22798 7812 22818 7834
rect 22818 7812 22832 7834
rect 22870 7812 22886 7834
rect 22886 7812 22904 7834
rect 22942 7812 22954 7834
rect 22954 7812 22976 7834
rect 23014 7812 23022 7834
rect 23022 7812 23048 7834
rect 23086 7812 23090 7834
rect 23090 7812 23120 7834
rect 23158 7812 23192 7834
rect 23230 7812 23260 7834
rect 23260 7812 23264 7834
rect 23302 7812 23328 7834
rect 23328 7812 23336 7834
rect 23374 7812 23396 7834
rect 23396 7812 23408 7834
rect 23446 7812 23464 7834
rect 23464 7812 23480 7834
rect 22798 7800 22832 7812
rect 22870 7800 22904 7812
rect 22942 7800 22976 7812
rect 23014 7800 23048 7812
rect 23086 7800 23120 7812
rect 23158 7800 23192 7812
rect 23230 7800 23264 7812
rect 23302 7800 23336 7812
rect 23374 7800 23408 7812
rect 23446 7800 23480 7812
rect 22798 7743 22818 7761
rect 22818 7743 22832 7761
rect 22870 7743 22886 7761
rect 22886 7743 22904 7761
rect 22942 7743 22954 7761
rect 22954 7743 22976 7761
rect 23014 7743 23022 7761
rect 23022 7743 23048 7761
rect 23086 7743 23090 7761
rect 23090 7743 23120 7761
rect 23158 7743 23192 7761
rect 23230 7743 23260 7761
rect 23260 7743 23264 7761
rect 23302 7743 23328 7761
rect 23328 7743 23336 7761
rect 23374 7743 23396 7761
rect 23396 7743 23408 7761
rect 23446 7743 23464 7761
rect 23464 7743 23480 7761
rect 22798 7727 22832 7743
rect 22870 7727 22904 7743
rect 22942 7727 22976 7743
rect 23014 7727 23048 7743
rect 23086 7727 23120 7743
rect 23158 7727 23192 7743
rect 23230 7727 23264 7743
rect 23302 7727 23336 7743
rect 23374 7727 23408 7743
rect 23446 7727 23480 7743
rect 22798 7674 22818 7688
rect 22818 7674 22832 7688
rect 22870 7674 22886 7688
rect 22886 7674 22904 7688
rect 22942 7674 22954 7688
rect 22954 7674 22976 7688
rect 23014 7674 23022 7688
rect 23022 7674 23048 7688
rect 23086 7674 23090 7688
rect 23090 7674 23120 7688
rect 23158 7674 23192 7688
rect 23230 7674 23260 7688
rect 23260 7674 23264 7688
rect 23302 7674 23328 7688
rect 23328 7674 23336 7688
rect 23374 7674 23396 7688
rect 23396 7674 23408 7688
rect 23446 7674 23464 7688
rect 23464 7674 23480 7688
rect 22798 7654 22832 7674
rect 22870 7654 22904 7674
rect 22942 7654 22976 7674
rect 23014 7654 23048 7674
rect 23086 7654 23120 7674
rect 23158 7654 23192 7674
rect 23230 7654 23264 7674
rect 23302 7654 23336 7674
rect 23374 7654 23408 7674
rect 23446 7654 23480 7674
rect 22798 7605 22818 7615
rect 22818 7605 22832 7615
rect 22870 7605 22886 7615
rect 22886 7605 22904 7615
rect 22942 7605 22954 7615
rect 22954 7605 22976 7615
rect 23014 7605 23022 7615
rect 23022 7605 23048 7615
rect 23086 7605 23090 7615
rect 23090 7605 23120 7615
rect 23158 7605 23192 7615
rect 23230 7605 23260 7615
rect 23260 7605 23264 7615
rect 23302 7605 23328 7615
rect 23328 7605 23336 7615
rect 23374 7605 23396 7615
rect 23396 7605 23408 7615
rect 23446 7605 23464 7615
rect 23464 7605 23480 7615
rect 22798 7581 22832 7605
rect 22870 7581 22904 7605
rect 22942 7581 22976 7605
rect 23014 7581 23048 7605
rect 23086 7581 23120 7605
rect 23158 7581 23192 7605
rect 23230 7581 23264 7605
rect 23302 7581 23336 7605
rect 23374 7581 23408 7605
rect 23446 7581 23480 7605
rect 22798 7536 22818 7542
rect 22818 7536 22832 7542
rect 22870 7536 22886 7542
rect 22886 7536 22904 7542
rect 22942 7536 22954 7542
rect 22954 7536 22976 7542
rect 23014 7536 23022 7542
rect 23022 7536 23048 7542
rect 23086 7536 23090 7542
rect 23090 7536 23120 7542
rect 23158 7536 23192 7542
rect 23230 7536 23260 7542
rect 23260 7536 23264 7542
rect 23302 7536 23328 7542
rect 23328 7536 23336 7542
rect 23374 7536 23396 7542
rect 23396 7536 23408 7542
rect 23446 7536 23464 7542
rect 23464 7536 23480 7542
rect 22798 7508 22832 7536
rect 22870 7508 22904 7536
rect 22942 7508 22976 7536
rect 23014 7508 23048 7536
rect 23086 7508 23120 7536
rect 23158 7508 23192 7536
rect 23230 7508 23264 7536
rect 23302 7508 23336 7536
rect 23374 7508 23408 7536
rect 23446 7508 23480 7536
rect 22798 7467 22818 7469
rect 22818 7467 22832 7469
rect 22870 7467 22886 7469
rect 22886 7467 22904 7469
rect 22942 7467 22954 7469
rect 22954 7467 22976 7469
rect 23014 7467 23022 7469
rect 23022 7467 23048 7469
rect 23086 7467 23090 7469
rect 23090 7467 23120 7469
rect 23158 7467 23192 7469
rect 23230 7467 23260 7469
rect 23260 7467 23264 7469
rect 23302 7467 23328 7469
rect 23328 7467 23336 7469
rect 23374 7467 23396 7469
rect 23396 7467 23408 7469
rect 23446 7467 23464 7469
rect 23464 7467 23480 7469
rect 22798 7435 22832 7467
rect 22870 7435 22904 7467
rect 22942 7435 22976 7467
rect 23014 7435 23048 7467
rect 23086 7435 23120 7467
rect 23158 7435 23192 7467
rect 23230 7435 23264 7467
rect 23302 7435 23336 7467
rect 23374 7435 23408 7467
rect 23446 7435 23480 7467
rect 22798 7363 22832 7396
rect 22870 7363 22904 7396
rect 22942 7363 22976 7396
rect 23014 7363 23048 7396
rect 23086 7363 23120 7396
rect 23158 7363 23192 7396
rect 23230 7363 23264 7396
rect 23302 7363 23336 7396
rect 23374 7363 23408 7396
rect 23446 7363 23480 7396
rect 22798 7362 22818 7363
rect 22818 7362 22832 7363
rect 22870 7362 22886 7363
rect 22886 7362 22904 7363
rect 22942 7362 22954 7363
rect 22954 7362 22976 7363
rect 23014 7362 23022 7363
rect 23022 7362 23048 7363
rect 23086 7362 23090 7363
rect 23090 7362 23120 7363
rect 23158 7362 23192 7363
rect 23230 7362 23260 7363
rect 23260 7362 23264 7363
rect 23302 7362 23328 7363
rect 23328 7362 23336 7363
rect 23374 7362 23396 7363
rect 23396 7362 23408 7363
rect 23446 7362 23464 7363
rect 23464 7362 23480 7363
rect 22798 7294 22832 7323
rect 22870 7294 22904 7323
rect 22942 7294 22976 7323
rect 23014 7294 23048 7323
rect 23086 7294 23120 7323
rect 23158 7294 23192 7323
rect 23230 7294 23264 7323
rect 23302 7294 23336 7323
rect 23374 7294 23408 7323
rect 23446 7294 23480 7323
rect 22798 7289 22818 7294
rect 22818 7289 22832 7294
rect 22870 7289 22886 7294
rect 22886 7289 22904 7294
rect 22942 7289 22954 7294
rect 22954 7289 22976 7294
rect 23014 7289 23022 7294
rect 23022 7289 23048 7294
rect 23086 7289 23090 7294
rect 23090 7289 23120 7294
rect 23158 7289 23192 7294
rect 23230 7289 23260 7294
rect 23260 7289 23264 7294
rect 23302 7289 23328 7294
rect 23328 7289 23336 7294
rect 23374 7289 23396 7294
rect 23396 7289 23408 7294
rect 23446 7289 23464 7294
rect 23464 7289 23480 7294
rect 22798 7225 22832 7250
rect 22870 7225 22904 7250
rect 22942 7225 22976 7250
rect 23014 7225 23048 7250
rect 23086 7225 23120 7250
rect 23158 7225 23192 7250
rect 23230 7225 23264 7250
rect 23302 7225 23336 7250
rect 23374 7225 23408 7250
rect 23446 7225 23480 7250
rect 22798 7216 22818 7225
rect 22818 7216 22832 7225
rect 22870 7216 22886 7225
rect 22886 7216 22904 7225
rect 22942 7216 22954 7225
rect 22954 7216 22976 7225
rect 23014 7216 23022 7225
rect 23022 7216 23048 7225
rect 23086 7216 23090 7225
rect 23090 7216 23120 7225
rect 23158 7216 23192 7225
rect 23230 7216 23260 7225
rect 23260 7216 23264 7225
rect 23302 7216 23328 7225
rect 23328 7216 23336 7225
rect 23374 7216 23396 7225
rect 23396 7216 23408 7225
rect 23446 7216 23464 7225
rect 23464 7216 23480 7225
rect 22798 7156 22832 7177
rect 22870 7156 22904 7177
rect 22942 7156 22976 7177
rect 23014 7156 23048 7177
rect 23086 7156 23120 7177
rect 23158 7156 23192 7177
rect 23230 7156 23264 7177
rect 23302 7156 23336 7177
rect 23374 7156 23408 7177
rect 23446 7156 23480 7177
rect 22798 7143 22818 7156
rect 22818 7143 22832 7156
rect 22870 7143 22886 7156
rect 22886 7143 22904 7156
rect 22942 7143 22954 7156
rect 22954 7143 22976 7156
rect 23014 7143 23022 7156
rect 23022 7143 23048 7156
rect 23086 7143 23090 7156
rect 23090 7143 23120 7156
rect 23158 7143 23192 7156
rect 23230 7143 23260 7156
rect 23260 7143 23264 7156
rect 23302 7143 23328 7156
rect 23328 7143 23336 7156
rect 23374 7143 23396 7156
rect 23396 7143 23408 7156
rect 23446 7143 23464 7156
rect 23464 7143 23480 7156
rect 22798 7087 22832 7104
rect 22870 7087 22904 7104
rect 22942 7087 22976 7104
rect 23014 7087 23048 7104
rect 23086 7087 23120 7104
rect 23158 7087 23192 7104
rect 23230 7087 23264 7104
rect 23302 7087 23336 7104
rect 23374 7087 23408 7104
rect 23446 7087 23480 7104
rect 22798 7070 22818 7087
rect 22818 7070 22832 7087
rect 22870 7070 22886 7087
rect 22886 7070 22904 7087
rect 22942 7070 22954 7087
rect 22954 7070 22976 7087
rect 23014 7070 23022 7087
rect 23022 7070 23048 7087
rect 23086 7070 23090 7087
rect 23090 7070 23120 7087
rect 23158 7070 23192 7087
rect 23230 7070 23260 7087
rect 23260 7070 23264 7087
rect 23302 7070 23328 7087
rect 23328 7070 23336 7087
rect 23374 7070 23396 7087
rect 23396 7070 23408 7087
rect 23446 7070 23464 7087
rect 23464 7070 23480 7087
rect 22798 7018 22832 7031
rect 22870 7018 22904 7031
rect 22942 7018 22976 7031
rect 23014 7018 23048 7031
rect 23086 7018 23120 7031
rect 23158 7018 23192 7031
rect 23230 7018 23264 7031
rect 23302 7018 23336 7031
rect 23374 7018 23408 7031
rect 23446 7018 23480 7031
rect 22798 6997 22818 7018
rect 22818 6997 22832 7018
rect 22870 6997 22886 7018
rect 22886 6997 22904 7018
rect 22942 6997 22954 7018
rect 22954 6997 22976 7018
rect 23014 6997 23022 7018
rect 23022 6997 23048 7018
rect 23086 6997 23090 7018
rect 23090 6997 23120 7018
rect 23158 6997 23192 7018
rect 23230 6997 23260 7018
rect 23260 6997 23264 7018
rect 23302 6997 23328 7018
rect 23328 6997 23336 7018
rect 23374 6997 23396 7018
rect 23396 6997 23408 7018
rect 23446 6997 23464 7018
rect 23464 6997 23480 7018
rect 22798 6949 22832 6958
rect 22870 6949 22904 6958
rect 22942 6949 22976 6958
rect 23014 6949 23048 6958
rect 23086 6949 23120 6958
rect 23158 6949 23192 6958
rect 23230 6949 23264 6958
rect 23302 6949 23336 6958
rect 23374 6949 23408 6958
rect 23446 6949 23480 6958
rect 22798 6924 22818 6949
rect 22818 6924 22832 6949
rect 22870 6924 22886 6949
rect 22886 6924 22904 6949
rect 22942 6924 22954 6949
rect 22954 6924 22976 6949
rect 23014 6924 23022 6949
rect 23022 6924 23048 6949
rect 23086 6924 23090 6949
rect 23090 6924 23120 6949
rect 23158 6924 23192 6949
rect 23230 6924 23260 6949
rect 23260 6924 23264 6949
rect 23302 6924 23328 6949
rect 23328 6924 23336 6949
rect 23374 6924 23396 6949
rect 23396 6924 23408 6949
rect 23446 6924 23464 6949
rect 23464 6924 23480 6949
rect 22798 6880 22832 6885
rect 22870 6880 22904 6885
rect 22942 6880 22976 6885
rect 23014 6880 23048 6885
rect 23086 6880 23120 6885
rect 23158 6880 23192 6885
rect 23230 6880 23264 6885
rect 23302 6880 23336 6885
rect 23374 6880 23408 6885
rect 23446 6880 23480 6885
rect 22798 6851 22818 6880
rect 22818 6851 22832 6880
rect 22870 6851 22886 6880
rect 22886 6851 22904 6880
rect 22942 6851 22954 6880
rect 22954 6851 22976 6880
rect 23014 6851 23022 6880
rect 23022 6851 23048 6880
rect 23086 6851 23090 6880
rect 23090 6851 23120 6880
rect 23158 6851 23192 6880
rect 23230 6851 23260 6880
rect 23260 6851 23264 6880
rect 23302 6851 23328 6880
rect 23328 6851 23336 6880
rect 23374 6851 23396 6880
rect 23396 6851 23408 6880
rect 23446 6851 23464 6880
rect 23464 6851 23480 6880
rect 22798 6811 22832 6812
rect 22870 6811 22904 6812
rect 22942 6811 22976 6812
rect 23014 6811 23048 6812
rect 23086 6811 23120 6812
rect 23158 6811 23192 6812
rect 23230 6811 23264 6812
rect 23302 6811 23336 6812
rect 23374 6811 23408 6812
rect 23446 6811 23480 6812
rect 22798 6778 22818 6811
rect 22818 6778 22832 6811
rect 22870 6778 22904 6811
rect 22942 6778 22976 6811
rect 23014 6778 23048 6811
rect 23086 6778 23120 6811
rect 23158 6778 23192 6811
rect 23230 6778 23264 6811
rect 23302 6778 23336 6811
rect 23374 6778 23408 6811
rect 23446 6778 23480 6811
rect 22798 6705 22818 6739
rect 22818 6705 22832 6739
rect 22870 6705 22904 6739
rect 22942 6705 22976 6739
rect 23014 6705 23048 6739
rect 23086 6705 23120 6739
rect 23158 6705 23192 6739
rect 23230 6705 23264 6739
rect 23302 6705 23336 6739
rect 23374 6705 23408 6739
rect 23446 6705 23480 6739
rect 22798 6632 22818 6666
rect 22818 6632 22832 6666
rect 22870 6632 22904 6666
rect 22942 6632 22976 6666
rect 23014 6632 23048 6666
rect 23086 6632 23120 6666
rect 23158 6632 23192 6666
rect 23230 6632 23264 6666
rect 23302 6632 23336 6666
rect 23374 6632 23408 6666
rect 23446 6632 23480 6666
rect 22798 6559 22818 6593
rect 22818 6559 22832 6593
rect 22870 6559 22904 6593
rect 22942 6559 22976 6593
rect 23014 6559 23048 6593
rect 23086 6559 23120 6593
rect 23158 6559 23192 6593
rect 23230 6559 23264 6593
rect 23302 6559 23336 6593
rect 23374 6559 23408 6593
rect 23446 6559 23480 6593
rect 22798 6486 22818 6520
rect 22818 6486 22832 6520
rect 22870 6486 22904 6520
rect 22942 6486 22976 6520
rect 23014 6486 23048 6520
rect 23086 6486 23120 6520
rect 23158 6486 23192 6520
rect 23230 6486 23264 6520
rect 23302 6486 23336 6520
rect 23374 6486 23408 6520
rect 23446 6486 23480 6520
rect 22798 6413 22818 6447
rect 22818 6413 22832 6447
rect 22870 6413 22904 6447
rect 22942 6413 22976 6447
rect 23014 6413 23048 6447
rect 23086 6413 23120 6447
rect 23158 6413 23192 6447
rect 23230 6413 23264 6447
rect 23302 6413 23336 6447
rect 23374 6413 23408 6447
rect 23446 6413 23480 6447
rect 22798 6340 22818 6374
rect 22818 6340 22832 6374
rect 22870 6340 22904 6374
rect 22942 6340 22976 6374
rect 23014 6340 23048 6374
rect 23086 6340 23120 6374
rect 23158 6340 23192 6374
rect 23230 6340 23264 6374
rect 23302 6340 23336 6374
rect 23374 6340 23408 6374
rect 23446 6340 23480 6374
rect 22798 6267 22818 6301
rect 22818 6267 22832 6301
rect 22870 6267 22904 6301
rect 22942 6267 22976 6301
rect 23014 6267 23048 6301
rect 23086 6267 23120 6301
rect 23158 6267 23192 6301
rect 23230 6267 23264 6301
rect 23302 6267 23336 6301
rect 23374 6267 23408 6301
rect 23446 6267 23480 6301
rect 22798 6194 22818 6228
rect 22818 6194 22832 6228
rect 22870 6194 22904 6228
rect 22942 6194 22976 6228
rect 23014 6194 23048 6228
rect 23086 6194 23120 6228
rect 23158 6194 23192 6228
rect 23230 6194 23264 6228
rect 23302 6194 23336 6228
rect 23374 6194 23408 6228
rect 23446 6194 23480 6228
rect 22798 6121 22818 6155
rect 22818 6121 22832 6155
rect 22870 6121 22904 6155
rect 22942 6121 22976 6155
rect 23014 6121 23048 6155
rect 23086 6121 23120 6155
rect 23158 6121 23192 6155
rect 23230 6121 23264 6155
rect 23302 6121 23336 6155
rect 23374 6121 23408 6155
rect 23446 6121 23480 6155
rect 22798 6048 22818 6082
rect 22818 6048 22832 6082
rect 22870 6048 22904 6082
rect 22942 6048 22976 6082
rect 23014 6048 23048 6082
rect 23086 6048 23120 6082
rect 23158 6048 23192 6082
rect 23230 6048 23264 6082
rect 23302 6048 23336 6082
rect 23374 6048 23408 6082
rect 23446 6048 23480 6082
rect 22798 5975 22818 6009
rect 22818 5975 22832 6009
rect 22870 5975 22904 6009
rect 22942 5975 22976 6009
rect 23014 5975 23048 6009
rect 23086 5975 23120 6009
rect 23158 5975 23192 6009
rect 23230 5975 23264 6009
rect 23302 5975 23336 6009
rect 23374 5975 23408 6009
rect 23446 5975 23480 6009
rect 22798 5902 22818 5936
rect 22818 5902 22832 5936
rect 22870 5902 22904 5936
rect 22942 5902 22976 5936
rect 23014 5902 23048 5936
rect 23086 5902 23120 5936
rect 23158 5902 23192 5936
rect 23230 5902 23264 5936
rect 23302 5902 23336 5936
rect 23374 5902 23408 5936
rect 23446 5902 23480 5936
rect 22798 5829 22818 5863
rect 22818 5829 22832 5863
rect 22870 5829 22904 5863
rect 22942 5829 22976 5863
rect 23014 5829 23048 5863
rect 23086 5829 23120 5863
rect 23158 5829 23192 5863
rect 23230 5829 23264 5863
rect 23302 5829 23336 5863
rect 23374 5829 23408 5863
rect 23446 5829 23480 5863
rect 22798 5756 22818 5790
rect 22818 5756 22832 5790
rect 22870 5756 22904 5790
rect 22942 5756 22976 5790
rect 23014 5756 23048 5790
rect 23086 5756 23120 5790
rect 23158 5756 23192 5790
rect 23230 5756 23264 5790
rect 23302 5756 23336 5790
rect 23374 5756 23408 5790
rect 23446 5756 23480 5790
rect 22798 5683 22818 5717
rect 22818 5683 22832 5717
rect 22870 5683 22904 5717
rect 22942 5683 22976 5717
rect 23014 5683 23048 5717
rect 23086 5683 23120 5717
rect 23158 5683 23192 5717
rect 23230 5683 23264 5717
rect 23302 5683 23336 5717
rect 23374 5683 23408 5717
rect 23446 5683 23480 5717
rect 22798 5610 22818 5644
rect 22818 5610 22832 5644
rect 22870 5610 22904 5644
rect 22942 5610 22976 5644
rect 23014 5610 23048 5644
rect 23086 5610 23120 5644
rect 23158 5610 23192 5644
rect 23230 5610 23264 5644
rect 23302 5610 23336 5644
rect 23374 5610 23408 5644
rect 23446 5610 23480 5644
rect 23781 8568 24370 8636
rect 24370 8568 24535 8636
rect 23781 8534 23789 8568
rect 23789 8534 23823 8568
rect 23823 8534 23857 8568
rect 23857 8534 23891 8568
rect 23891 8534 23925 8568
rect 23925 8534 23959 8568
rect 23959 8534 23993 8568
rect 23993 8534 24027 8568
rect 24027 8534 24061 8568
rect 24061 8534 24095 8568
rect 24095 8534 24129 8568
rect 24129 8534 24163 8568
rect 24163 8534 24197 8568
rect 24197 8534 24231 8568
rect 24231 8534 24265 8568
rect 24265 8534 24299 8568
rect 24299 8534 24333 8568
rect 24333 8534 24367 8568
rect 24367 8534 24535 8568
rect 23781 8499 24535 8534
rect 23781 8465 23789 8499
rect 23789 8465 23823 8499
rect 23823 8465 23857 8499
rect 23857 8465 23891 8499
rect 23891 8465 23925 8499
rect 23925 8465 23959 8499
rect 23959 8465 23993 8499
rect 23993 8465 24027 8499
rect 24027 8465 24061 8499
rect 24061 8465 24095 8499
rect 24095 8465 24129 8499
rect 24129 8465 24163 8499
rect 24163 8465 24197 8499
rect 24197 8465 24231 8499
rect 24231 8465 24265 8499
rect 24265 8465 24299 8499
rect 24299 8465 24333 8499
rect 24333 8465 24367 8499
rect 24367 8465 24401 8499
rect 24401 8465 24435 8499
rect 24435 8465 24469 8499
rect 24469 8465 24503 8499
rect 24503 8465 24535 8499
rect 23781 8430 24535 8465
rect 23781 8396 23789 8430
rect 23789 8396 23823 8430
rect 23823 8396 23857 8430
rect 23857 8396 23891 8430
rect 23891 8396 23925 8430
rect 23925 8396 23959 8430
rect 23959 8396 23993 8430
rect 23993 8396 24027 8430
rect 24027 8396 24061 8430
rect 24061 8396 24095 8430
rect 24095 8396 24129 8430
rect 24129 8396 24163 8430
rect 24163 8396 24197 8430
rect 24197 8396 24231 8430
rect 24231 8396 24265 8430
rect 24265 8396 24299 8430
rect 24299 8396 24333 8430
rect 24333 8396 24367 8430
rect 24367 8396 24401 8430
rect 24401 8396 24435 8430
rect 24435 8396 24469 8430
rect 24469 8396 24503 8430
rect 24503 8396 24535 8430
rect 23781 8361 24535 8396
rect 23781 8327 23789 8361
rect 23789 8327 23823 8361
rect 23823 8327 23857 8361
rect 23857 8327 23891 8361
rect 23891 8327 23925 8361
rect 23925 8327 23959 8361
rect 23959 8327 23993 8361
rect 23993 8327 24027 8361
rect 24027 8327 24061 8361
rect 24061 8327 24095 8361
rect 24095 8327 24129 8361
rect 24129 8327 24163 8361
rect 24163 8327 24197 8361
rect 24197 8327 24231 8361
rect 24231 8327 24265 8361
rect 24265 8327 24299 8361
rect 24299 8327 24333 8361
rect 24333 8327 24367 8361
rect 24367 8327 24401 8361
rect 24401 8327 24435 8361
rect 24435 8327 24469 8361
rect 24469 8327 24503 8361
rect 24503 8327 24535 8361
rect 23781 8292 24535 8327
rect 23781 8258 23789 8292
rect 23789 8258 23823 8292
rect 23823 8258 23857 8292
rect 23857 8258 23891 8292
rect 23891 8258 23925 8292
rect 23925 8258 23959 8292
rect 23959 8258 23993 8292
rect 23993 8258 24027 8292
rect 24027 8258 24061 8292
rect 24061 8258 24095 8292
rect 24095 8258 24129 8292
rect 24129 8258 24163 8292
rect 24163 8258 24197 8292
rect 24197 8258 24231 8292
rect 24231 8258 24265 8292
rect 24265 8258 24299 8292
rect 24299 8258 24333 8292
rect 24333 8258 24367 8292
rect 24367 8258 24401 8292
rect 24401 8258 24435 8292
rect 24435 8258 24469 8292
rect 24469 8258 24503 8292
rect 24503 8258 24535 8292
rect 23781 8223 24535 8258
rect 23781 8189 23789 8223
rect 23789 8189 23823 8223
rect 23823 8189 23857 8223
rect 23857 8189 23891 8223
rect 23891 8189 23925 8223
rect 23925 8189 23959 8223
rect 23959 8189 23993 8223
rect 23993 8189 24027 8223
rect 24027 8189 24061 8223
rect 24061 8189 24095 8223
rect 24095 8189 24129 8223
rect 24129 8189 24163 8223
rect 24163 8189 24197 8223
rect 24197 8189 24231 8223
rect 24231 8189 24265 8223
rect 24265 8189 24299 8223
rect 24299 8189 24333 8223
rect 24333 8189 24367 8223
rect 24367 8189 24401 8223
rect 24401 8189 24435 8223
rect 24435 8189 24469 8223
rect 24469 8189 24503 8223
rect 24503 8189 24535 8223
rect 23781 8154 24535 8189
rect 23781 8120 23789 8154
rect 23789 8120 23823 8154
rect 23823 8120 23857 8154
rect 23857 8120 23891 8154
rect 23891 8120 23925 8154
rect 23925 8120 23959 8154
rect 23959 8120 23993 8154
rect 23993 8120 24027 8154
rect 24027 8120 24061 8154
rect 24061 8120 24095 8154
rect 24095 8120 24129 8154
rect 24129 8120 24163 8154
rect 24163 8120 24197 8154
rect 24197 8120 24231 8154
rect 24231 8120 24265 8154
rect 24265 8120 24299 8154
rect 24299 8120 24333 8154
rect 24333 8120 24367 8154
rect 24367 8120 24401 8154
rect 24401 8120 24435 8154
rect 24435 8120 24469 8154
rect 24469 8120 24503 8154
rect 24503 8120 24535 8154
rect 23781 8085 24535 8120
rect 23781 8051 23789 8085
rect 23789 8051 23823 8085
rect 23823 8051 23857 8085
rect 23857 8051 23891 8085
rect 23891 8051 23925 8085
rect 23925 8051 23959 8085
rect 23959 8051 23993 8085
rect 23993 8051 24027 8085
rect 24027 8051 24061 8085
rect 24061 8051 24095 8085
rect 24095 8051 24129 8085
rect 24129 8051 24163 8085
rect 24163 8051 24197 8085
rect 24197 8051 24231 8085
rect 24231 8051 24265 8085
rect 24265 8051 24299 8085
rect 24299 8051 24333 8085
rect 24333 8051 24367 8085
rect 24367 8051 24401 8085
rect 24401 8051 24435 8085
rect 24435 8051 24469 8085
rect 24469 8051 24503 8085
rect 24503 8051 24535 8085
rect 23781 8016 24535 8051
rect 23781 7982 23789 8016
rect 23789 7982 23823 8016
rect 23823 7982 23857 8016
rect 23857 7982 23891 8016
rect 23891 7982 23925 8016
rect 23925 7982 23959 8016
rect 23959 7982 23993 8016
rect 23993 7982 24027 8016
rect 24027 7982 24061 8016
rect 24061 7982 24095 8016
rect 24095 7982 24129 8016
rect 24129 7982 24163 8016
rect 24163 7982 24197 8016
rect 24197 7982 24231 8016
rect 24231 7982 24265 8016
rect 24265 7982 24299 8016
rect 24299 7982 24333 8016
rect 24333 7982 24367 8016
rect 24367 7982 24401 8016
rect 24401 7982 24435 8016
rect 24435 7982 24469 8016
rect 24469 7982 24503 8016
rect 24503 7982 24535 8016
rect 23781 7947 24535 7982
rect 23781 7913 23789 7947
rect 23789 7913 23823 7947
rect 23823 7913 23857 7947
rect 23857 7913 23891 7947
rect 23891 7913 23925 7947
rect 23925 7913 23959 7947
rect 23959 7913 23993 7947
rect 23993 7913 24027 7947
rect 24027 7913 24061 7947
rect 24061 7913 24095 7947
rect 24095 7913 24129 7947
rect 24129 7913 24163 7947
rect 24163 7913 24197 7947
rect 24197 7913 24231 7947
rect 24231 7913 24265 7947
rect 24265 7913 24299 7947
rect 24299 7913 24333 7947
rect 24333 7913 24367 7947
rect 24367 7913 24401 7947
rect 24401 7913 24435 7947
rect 24435 7913 24469 7947
rect 24469 7913 24503 7947
rect 24503 7913 24535 7947
rect 23781 7878 24535 7913
rect 23781 7854 23789 7878
rect 23789 7854 23823 7878
rect 23823 7854 23857 7878
rect 23857 7854 23891 7878
rect 23891 7854 23925 7878
rect 23925 7854 23959 7878
rect 23959 7854 23993 7878
rect 23993 7854 24027 7878
rect 24027 7854 24061 7878
rect 24061 7854 24095 7878
rect 24095 7854 24129 7878
rect 24129 7854 24163 7878
rect 24163 7854 24197 7878
rect 24197 7854 24231 7878
rect 24231 7854 24265 7878
rect 24265 7854 24299 7878
rect 24299 7854 24333 7878
rect 24333 7854 24367 7878
rect 24367 7854 24401 7878
rect 24401 7854 24435 7878
rect 24435 7854 24469 7878
rect 24469 7854 24503 7878
rect 24503 7854 24535 7878
rect 23781 7809 23815 7815
rect 23853 7809 23887 7815
rect 23781 7781 23789 7809
rect 23789 7781 23815 7809
rect 23853 7781 23857 7809
rect 23857 7781 23887 7809
rect 23925 7781 23959 7815
rect 23997 7809 24031 7815
rect 24069 7809 24103 7815
rect 24141 7809 24175 7815
rect 24213 7809 24247 7815
rect 24285 7809 24319 7815
rect 24357 7809 24391 7815
rect 24429 7809 24463 7815
rect 24501 7809 24535 7815
rect 23997 7781 24027 7809
rect 24027 7781 24031 7809
rect 24069 7781 24095 7809
rect 24095 7781 24103 7809
rect 24141 7781 24163 7809
rect 24163 7781 24175 7809
rect 24213 7781 24231 7809
rect 24231 7781 24247 7809
rect 24285 7781 24299 7809
rect 24299 7781 24319 7809
rect 24357 7781 24367 7809
rect 24367 7781 24391 7809
rect 24429 7781 24435 7809
rect 24435 7781 24463 7809
rect 24501 7781 24503 7809
rect 24503 7781 24535 7809
rect 23781 7740 23815 7742
rect 23853 7740 23887 7742
rect 23781 7708 23789 7740
rect 23789 7708 23815 7740
rect 23853 7708 23857 7740
rect 23857 7708 23887 7740
rect 23925 7708 23959 7742
rect 23997 7740 24031 7742
rect 24069 7740 24103 7742
rect 24141 7740 24175 7742
rect 24213 7740 24247 7742
rect 24285 7740 24319 7742
rect 24357 7740 24391 7742
rect 24429 7740 24463 7742
rect 24501 7740 24535 7742
rect 23997 7708 24027 7740
rect 24027 7708 24031 7740
rect 24069 7708 24095 7740
rect 24095 7708 24103 7740
rect 24141 7708 24163 7740
rect 24163 7708 24175 7740
rect 24213 7708 24231 7740
rect 24231 7708 24247 7740
rect 24285 7708 24299 7740
rect 24299 7708 24319 7740
rect 24357 7708 24367 7740
rect 24367 7708 24391 7740
rect 24429 7708 24435 7740
rect 24435 7708 24463 7740
rect 24501 7708 24503 7740
rect 24503 7708 24535 7740
rect 23781 7637 23789 7669
rect 23789 7637 23815 7669
rect 23853 7637 23857 7669
rect 23857 7637 23887 7669
rect 23781 7635 23815 7637
rect 23853 7635 23887 7637
rect 23925 7635 23959 7669
rect 23997 7637 24027 7669
rect 24027 7637 24031 7669
rect 24069 7637 24095 7669
rect 24095 7637 24103 7669
rect 24141 7637 24163 7669
rect 24163 7637 24175 7669
rect 24213 7637 24231 7669
rect 24231 7637 24247 7669
rect 24285 7637 24299 7669
rect 24299 7637 24319 7669
rect 24357 7637 24367 7669
rect 24367 7637 24391 7669
rect 24429 7637 24435 7669
rect 24435 7637 24463 7669
rect 24501 7637 24503 7669
rect 24503 7637 24535 7669
rect 23997 7635 24031 7637
rect 24069 7635 24103 7637
rect 24141 7635 24175 7637
rect 24213 7635 24247 7637
rect 24285 7635 24319 7637
rect 24357 7635 24391 7637
rect 24429 7635 24463 7637
rect 24501 7635 24535 7637
rect 23781 7568 23789 7596
rect 23789 7568 23815 7596
rect 23853 7568 23857 7596
rect 23857 7568 23887 7596
rect 23781 7562 23815 7568
rect 23853 7562 23887 7568
rect 23925 7562 23959 7596
rect 23997 7568 24027 7596
rect 24027 7568 24031 7596
rect 24069 7568 24095 7596
rect 24095 7568 24103 7596
rect 24141 7568 24163 7596
rect 24163 7568 24175 7596
rect 24213 7568 24231 7596
rect 24231 7568 24247 7596
rect 24285 7568 24299 7596
rect 24299 7568 24319 7596
rect 24357 7568 24367 7596
rect 24367 7568 24391 7596
rect 24429 7568 24435 7596
rect 24435 7568 24463 7596
rect 24501 7568 24503 7596
rect 24503 7568 24535 7596
rect 23997 7562 24031 7568
rect 24069 7562 24103 7568
rect 24141 7562 24175 7568
rect 24213 7562 24247 7568
rect 24285 7562 24319 7568
rect 24357 7562 24391 7568
rect 24429 7562 24463 7568
rect 24501 7562 24535 7568
rect 23781 7499 23789 7523
rect 23789 7499 23815 7523
rect 23853 7499 23857 7523
rect 23857 7499 23887 7523
rect 23781 7489 23815 7499
rect 23853 7489 23887 7499
rect 23925 7489 23959 7523
rect 23997 7499 24027 7523
rect 24027 7499 24031 7523
rect 24069 7499 24095 7523
rect 24095 7499 24103 7523
rect 24141 7499 24163 7523
rect 24163 7499 24175 7523
rect 24213 7499 24231 7523
rect 24231 7499 24247 7523
rect 24285 7499 24299 7523
rect 24299 7499 24319 7523
rect 24357 7499 24367 7523
rect 24367 7499 24391 7523
rect 24429 7499 24435 7523
rect 24435 7499 24463 7523
rect 24501 7499 24503 7523
rect 24503 7499 24535 7523
rect 23997 7489 24031 7499
rect 24069 7489 24103 7499
rect 24141 7489 24175 7499
rect 24213 7489 24247 7499
rect 24285 7489 24319 7499
rect 24357 7489 24391 7499
rect 24429 7489 24463 7499
rect 24501 7489 24535 7499
rect 23781 7430 23789 7450
rect 23789 7430 23815 7450
rect 23853 7430 23857 7450
rect 23857 7430 23887 7450
rect 23781 7416 23815 7430
rect 23853 7416 23887 7430
rect 23925 7416 23959 7450
rect 23997 7430 24027 7450
rect 24027 7430 24031 7450
rect 24069 7430 24095 7450
rect 24095 7430 24103 7450
rect 24141 7430 24163 7450
rect 24163 7430 24175 7450
rect 24213 7430 24231 7450
rect 24231 7430 24247 7450
rect 24285 7430 24299 7450
rect 24299 7430 24319 7450
rect 24357 7430 24367 7450
rect 24367 7430 24391 7450
rect 24429 7430 24435 7450
rect 24435 7430 24463 7450
rect 24501 7430 24503 7450
rect 24503 7430 24535 7450
rect 23997 7416 24031 7430
rect 24069 7416 24103 7430
rect 24141 7416 24175 7430
rect 24213 7416 24247 7430
rect 24285 7416 24319 7430
rect 24357 7416 24391 7430
rect 24429 7416 24463 7430
rect 24501 7416 24535 7430
rect 23781 7361 23789 7377
rect 23789 7361 23815 7377
rect 23853 7361 23857 7377
rect 23857 7361 23887 7377
rect 23781 7343 23815 7361
rect 23853 7343 23887 7361
rect 23925 7343 23959 7377
rect 23997 7361 24027 7377
rect 24027 7361 24031 7377
rect 24069 7361 24095 7377
rect 24095 7361 24103 7377
rect 24141 7361 24163 7377
rect 24163 7361 24175 7377
rect 24213 7361 24231 7377
rect 24231 7361 24247 7377
rect 24285 7361 24299 7377
rect 24299 7361 24319 7377
rect 24357 7361 24367 7377
rect 24367 7361 24391 7377
rect 24429 7361 24435 7377
rect 24435 7361 24463 7377
rect 24501 7361 24503 7377
rect 24503 7361 24535 7377
rect 23997 7343 24031 7361
rect 24069 7343 24103 7361
rect 24141 7343 24175 7361
rect 24213 7343 24247 7361
rect 24285 7343 24319 7361
rect 24357 7343 24391 7361
rect 24429 7343 24463 7361
rect 24501 7343 24535 7361
rect 23781 7292 23789 7304
rect 23789 7292 23815 7304
rect 23853 7292 23857 7304
rect 23857 7292 23887 7304
rect 23781 7270 23815 7292
rect 23853 7270 23887 7292
rect 23925 7270 23959 7304
rect 23997 7292 24027 7304
rect 24027 7292 24031 7304
rect 24069 7292 24095 7304
rect 24095 7292 24103 7304
rect 24141 7292 24163 7304
rect 24163 7292 24175 7304
rect 24213 7292 24231 7304
rect 24231 7292 24247 7304
rect 24285 7292 24299 7304
rect 24299 7292 24319 7304
rect 24357 7292 24367 7304
rect 24367 7292 24391 7304
rect 24429 7292 24435 7304
rect 24435 7292 24463 7304
rect 24501 7292 24503 7304
rect 24503 7292 24535 7304
rect 23997 7270 24031 7292
rect 24069 7270 24103 7292
rect 24141 7270 24175 7292
rect 24213 7270 24247 7292
rect 24285 7270 24319 7292
rect 24357 7270 24391 7292
rect 24429 7270 24463 7292
rect 24501 7270 24535 7292
rect 23781 7223 23789 7231
rect 23789 7223 23815 7231
rect 23853 7223 23857 7231
rect 23857 7223 23887 7231
rect 23781 7197 23815 7223
rect 23853 7197 23887 7223
rect 23925 7197 23959 7231
rect 23997 7223 24027 7231
rect 24027 7223 24031 7231
rect 24069 7223 24095 7231
rect 24095 7223 24103 7231
rect 24141 7223 24163 7231
rect 24163 7223 24175 7231
rect 24213 7223 24231 7231
rect 24231 7223 24247 7231
rect 24285 7223 24299 7231
rect 24299 7223 24319 7231
rect 24357 7223 24367 7231
rect 24367 7223 24391 7231
rect 24429 7223 24435 7231
rect 24435 7223 24463 7231
rect 24501 7223 24503 7231
rect 24503 7223 24535 7231
rect 23997 7197 24031 7223
rect 24069 7197 24103 7223
rect 24141 7197 24175 7223
rect 24213 7197 24247 7223
rect 24285 7197 24319 7223
rect 24357 7197 24391 7223
rect 24429 7197 24463 7223
rect 24501 7197 24535 7223
rect 23781 7154 23789 7158
rect 23789 7154 23815 7158
rect 23853 7154 23857 7158
rect 23857 7154 23887 7158
rect 23781 7124 23815 7154
rect 23853 7124 23887 7154
rect 23925 7124 23959 7158
rect 23997 7154 24027 7158
rect 24027 7154 24031 7158
rect 24069 7154 24095 7158
rect 24095 7154 24103 7158
rect 24141 7154 24163 7158
rect 24163 7154 24175 7158
rect 24213 7154 24231 7158
rect 24231 7154 24247 7158
rect 24285 7154 24299 7158
rect 24299 7154 24319 7158
rect 24357 7154 24367 7158
rect 24367 7154 24391 7158
rect 24429 7154 24435 7158
rect 24435 7154 24463 7158
rect 24501 7154 24503 7158
rect 24503 7154 24535 7158
rect 23997 7124 24031 7154
rect 24069 7124 24103 7154
rect 24141 7124 24175 7154
rect 24213 7124 24247 7154
rect 24285 7124 24319 7154
rect 24357 7124 24391 7154
rect 24429 7124 24463 7154
rect 24501 7124 24535 7154
rect 23781 7051 23815 7085
rect 23853 7051 23887 7085
rect 23925 7051 23959 7085
rect 23997 7051 24031 7085
rect 24069 7051 24103 7085
rect 24141 7051 24175 7085
rect 24213 7051 24247 7085
rect 24285 7051 24319 7085
rect 24357 7051 24391 7085
rect 24429 7051 24463 7085
rect 24501 7051 24535 7085
rect 23781 6981 23815 7012
rect 23853 6981 23887 7012
rect 23781 6978 23789 6981
rect 23789 6978 23815 6981
rect 23853 6978 23857 6981
rect 23857 6978 23887 6981
rect 23925 6978 23959 7012
rect 23997 6981 24031 7012
rect 24069 6981 24103 7012
rect 24141 6981 24175 7012
rect 24213 6981 24247 7012
rect 24285 6981 24319 7012
rect 24357 6981 24391 7012
rect 24429 6981 24463 7012
rect 24501 6981 24535 7012
rect 23997 6978 24027 6981
rect 24027 6978 24031 6981
rect 24069 6978 24095 6981
rect 24095 6978 24103 6981
rect 24141 6978 24163 6981
rect 24163 6978 24175 6981
rect 24213 6978 24231 6981
rect 24231 6978 24247 6981
rect 24285 6978 24299 6981
rect 24299 6978 24319 6981
rect 24357 6978 24367 6981
rect 24367 6978 24391 6981
rect 24429 6978 24435 6981
rect 24435 6978 24463 6981
rect 24501 6978 24503 6981
rect 24503 6978 24535 6981
rect 23781 6912 23815 6939
rect 23853 6912 23887 6939
rect 23781 6905 23789 6912
rect 23789 6905 23815 6912
rect 23853 6905 23857 6912
rect 23857 6905 23887 6912
rect 23925 6905 23959 6939
rect 23997 6912 24031 6939
rect 24069 6912 24103 6939
rect 24141 6912 24175 6939
rect 24213 6912 24247 6939
rect 24285 6912 24319 6939
rect 24357 6912 24391 6939
rect 24429 6912 24463 6939
rect 24501 6912 24535 6939
rect 23997 6905 24027 6912
rect 24027 6905 24031 6912
rect 24069 6905 24095 6912
rect 24095 6905 24103 6912
rect 24141 6905 24163 6912
rect 24163 6905 24175 6912
rect 24213 6905 24231 6912
rect 24231 6905 24247 6912
rect 24285 6905 24299 6912
rect 24299 6905 24319 6912
rect 24357 6905 24367 6912
rect 24367 6905 24391 6912
rect 24429 6905 24435 6912
rect 24435 6905 24463 6912
rect 24501 6905 24503 6912
rect 24503 6905 24535 6912
rect 23781 6843 23815 6866
rect 23853 6843 23887 6866
rect 23781 6832 23789 6843
rect 23789 6832 23815 6843
rect 23853 6832 23857 6843
rect 23857 6832 23887 6843
rect 23925 6832 23959 6866
rect 23997 6843 24031 6866
rect 24069 6843 24103 6866
rect 24141 6843 24175 6866
rect 24213 6843 24247 6866
rect 24285 6843 24319 6866
rect 24357 6843 24391 6866
rect 24429 6843 24463 6866
rect 24501 6843 24535 6866
rect 23997 6832 24027 6843
rect 24027 6832 24031 6843
rect 24069 6832 24095 6843
rect 24095 6832 24103 6843
rect 24141 6832 24163 6843
rect 24163 6832 24175 6843
rect 24213 6832 24231 6843
rect 24231 6832 24247 6843
rect 24285 6832 24299 6843
rect 24299 6832 24319 6843
rect 24357 6832 24367 6843
rect 24367 6832 24391 6843
rect 24429 6832 24435 6843
rect 24435 6832 24463 6843
rect 24501 6832 24503 6843
rect 24503 6832 24535 6843
rect 23781 6774 23815 6793
rect 23853 6774 23887 6793
rect 23781 6759 23789 6774
rect 23789 6759 23815 6774
rect 23853 6759 23857 6774
rect 23857 6759 23887 6774
rect 23925 6759 23959 6793
rect 23997 6774 24031 6793
rect 24069 6774 24103 6793
rect 24141 6774 24175 6793
rect 24213 6774 24247 6793
rect 24285 6774 24319 6793
rect 24357 6774 24391 6793
rect 24429 6774 24463 6793
rect 24501 6774 24535 6793
rect 23997 6759 24027 6774
rect 24027 6759 24031 6774
rect 24069 6759 24095 6774
rect 24095 6759 24103 6774
rect 24141 6759 24163 6774
rect 24163 6759 24175 6774
rect 24213 6759 24231 6774
rect 24231 6759 24247 6774
rect 24285 6759 24299 6774
rect 24299 6759 24319 6774
rect 24357 6759 24367 6774
rect 24367 6759 24391 6774
rect 24429 6759 24435 6774
rect 24435 6759 24463 6774
rect 24501 6759 24503 6774
rect 24503 6759 24535 6774
rect 23781 6705 23815 6720
rect 23853 6705 23887 6720
rect 23781 6686 23789 6705
rect 23789 6686 23815 6705
rect 23853 6686 23857 6705
rect 23857 6686 23887 6705
rect 23925 6686 23959 6720
rect 23997 6705 24031 6720
rect 24069 6705 24103 6720
rect 24141 6705 24175 6720
rect 24213 6705 24247 6720
rect 24285 6705 24319 6720
rect 24357 6705 24391 6720
rect 24429 6705 24463 6720
rect 24501 6705 24535 6720
rect 23997 6686 24027 6705
rect 24027 6686 24031 6705
rect 24069 6686 24095 6705
rect 24095 6686 24103 6705
rect 24141 6686 24163 6705
rect 24163 6686 24175 6705
rect 24213 6686 24231 6705
rect 24231 6686 24247 6705
rect 24285 6686 24299 6705
rect 24299 6686 24319 6705
rect 24357 6686 24367 6705
rect 24367 6686 24391 6705
rect 24429 6686 24435 6705
rect 24435 6686 24463 6705
rect 24501 6686 24503 6705
rect 24503 6686 24535 6705
rect 23781 6636 23815 6647
rect 23853 6636 23887 6647
rect 23781 6613 23789 6636
rect 23789 6613 23815 6636
rect 23853 6613 23857 6636
rect 23857 6613 23887 6636
rect 23925 6613 23959 6647
rect 23997 6636 24031 6647
rect 24069 6636 24103 6647
rect 24141 6636 24175 6647
rect 24213 6636 24247 6647
rect 24285 6636 24319 6647
rect 24357 6636 24391 6647
rect 24429 6636 24463 6647
rect 24501 6636 24535 6647
rect 23997 6613 24027 6636
rect 24027 6613 24031 6636
rect 24069 6613 24095 6636
rect 24095 6613 24103 6636
rect 24141 6613 24163 6636
rect 24163 6613 24175 6636
rect 24213 6613 24231 6636
rect 24231 6613 24247 6636
rect 24285 6613 24299 6636
rect 24299 6613 24319 6636
rect 24357 6613 24367 6636
rect 24367 6613 24391 6636
rect 24429 6613 24435 6636
rect 24435 6613 24463 6636
rect 24501 6613 24503 6636
rect 24503 6613 24535 6636
rect 23781 6567 23815 6574
rect 23853 6567 23887 6574
rect 23781 6540 23789 6567
rect 23789 6540 23815 6567
rect 23853 6540 23857 6567
rect 23857 6540 23887 6567
rect 23925 6540 23959 6574
rect 23997 6567 24031 6574
rect 24069 6567 24103 6574
rect 24141 6567 24175 6574
rect 24213 6567 24247 6574
rect 24285 6567 24319 6574
rect 24357 6567 24391 6574
rect 24429 6567 24463 6574
rect 24501 6567 24535 6574
rect 23997 6540 24027 6567
rect 24027 6540 24031 6567
rect 24069 6540 24095 6567
rect 24095 6540 24103 6567
rect 24141 6540 24163 6567
rect 24163 6540 24175 6567
rect 24213 6540 24231 6567
rect 24231 6540 24247 6567
rect 24285 6540 24299 6567
rect 24299 6540 24319 6567
rect 24357 6540 24367 6567
rect 24367 6540 24391 6567
rect 24429 6540 24435 6567
rect 24435 6540 24463 6567
rect 24501 6540 24503 6567
rect 24503 6540 24535 6567
rect 23781 6498 23815 6501
rect 23853 6498 23887 6501
rect 23781 6467 23789 6498
rect 23789 6467 23815 6498
rect 23853 6467 23857 6498
rect 23857 6467 23887 6498
rect 23925 6467 23959 6501
rect 23997 6498 24031 6501
rect 24069 6498 24103 6501
rect 24141 6498 24175 6501
rect 24213 6498 24247 6501
rect 24285 6498 24319 6501
rect 24357 6498 24391 6501
rect 24429 6498 24463 6501
rect 24501 6498 24535 6501
rect 23997 6467 24027 6498
rect 24027 6467 24031 6498
rect 24069 6467 24095 6498
rect 24095 6467 24103 6498
rect 24141 6467 24163 6498
rect 24163 6467 24175 6498
rect 24213 6467 24231 6498
rect 24231 6467 24247 6498
rect 24285 6467 24299 6498
rect 24299 6467 24319 6498
rect 24357 6467 24367 6498
rect 24367 6467 24391 6498
rect 24429 6467 24435 6498
rect 24435 6467 24463 6498
rect 24501 6467 24503 6498
rect 24503 6467 24535 6498
rect 23781 6395 23789 6428
rect 23789 6395 23815 6428
rect 23853 6395 23857 6428
rect 23857 6395 23887 6428
rect 23781 6394 23815 6395
rect 23853 6394 23887 6395
rect 23925 6394 23959 6428
rect 23997 6395 24027 6428
rect 24027 6395 24031 6428
rect 24069 6395 24095 6428
rect 24095 6395 24103 6428
rect 24141 6395 24163 6428
rect 24163 6395 24175 6428
rect 24213 6395 24231 6428
rect 24231 6395 24247 6428
rect 24285 6395 24299 6428
rect 24299 6395 24319 6428
rect 24357 6395 24367 6428
rect 24367 6395 24391 6428
rect 24429 6395 24435 6428
rect 24435 6395 24463 6428
rect 24501 6395 24503 6428
rect 24503 6395 24535 6428
rect 23997 6394 24031 6395
rect 24069 6394 24103 6395
rect 24141 6394 24175 6395
rect 24213 6394 24247 6395
rect 24285 6394 24319 6395
rect 24357 6394 24391 6395
rect 24429 6394 24463 6395
rect 24501 6394 24535 6395
rect 23781 6326 23789 6355
rect 23789 6326 23815 6355
rect 23853 6326 23857 6355
rect 23857 6326 23887 6355
rect 23781 6321 23815 6326
rect 23853 6321 23887 6326
rect 23925 6321 23959 6355
rect 23997 6326 24027 6355
rect 24027 6326 24031 6355
rect 24069 6326 24095 6355
rect 24095 6326 24103 6355
rect 24141 6326 24163 6355
rect 24163 6326 24175 6355
rect 24213 6326 24231 6355
rect 24231 6326 24247 6355
rect 24285 6326 24299 6355
rect 24299 6326 24319 6355
rect 24357 6326 24367 6355
rect 24367 6326 24391 6355
rect 24429 6326 24435 6355
rect 24435 6326 24463 6355
rect 24501 6326 24503 6355
rect 24503 6326 24535 6355
rect 23997 6321 24031 6326
rect 24069 6321 24103 6326
rect 24141 6321 24175 6326
rect 24213 6321 24247 6326
rect 24285 6321 24319 6326
rect 24357 6321 24391 6326
rect 24429 6321 24463 6326
rect 24501 6321 24535 6326
rect 23781 6257 23789 6282
rect 23789 6257 23815 6282
rect 23853 6257 23857 6282
rect 23857 6257 23887 6282
rect 23781 6248 23815 6257
rect 23853 6248 23887 6257
rect 23925 6248 23959 6282
rect 23997 6257 24027 6282
rect 24027 6257 24031 6282
rect 24069 6257 24095 6282
rect 24095 6257 24103 6282
rect 24141 6257 24163 6282
rect 24163 6257 24175 6282
rect 24213 6257 24231 6282
rect 24231 6257 24247 6282
rect 24285 6257 24299 6282
rect 24299 6257 24319 6282
rect 24357 6257 24367 6282
rect 24367 6257 24391 6282
rect 24429 6257 24435 6282
rect 24435 6257 24463 6282
rect 24501 6257 24503 6282
rect 24503 6257 24535 6282
rect 23997 6248 24031 6257
rect 24069 6248 24103 6257
rect 24141 6248 24175 6257
rect 24213 6248 24247 6257
rect 24285 6248 24319 6257
rect 24357 6248 24391 6257
rect 24429 6248 24463 6257
rect 24501 6248 24535 6257
rect 23781 6188 23789 6209
rect 23789 6188 23815 6209
rect 23853 6188 23857 6209
rect 23857 6188 23887 6209
rect 23781 6175 23815 6188
rect 23853 6175 23887 6188
rect 23925 6175 23959 6209
rect 23997 6188 24027 6209
rect 24027 6188 24031 6209
rect 24069 6188 24095 6209
rect 24095 6188 24103 6209
rect 24141 6188 24163 6209
rect 24163 6188 24175 6209
rect 24213 6188 24231 6209
rect 24231 6188 24247 6209
rect 24285 6188 24299 6209
rect 24299 6188 24319 6209
rect 24357 6188 24367 6209
rect 24367 6188 24391 6209
rect 24429 6188 24435 6209
rect 24435 6188 24463 6209
rect 24501 6188 24503 6209
rect 24503 6188 24535 6209
rect 23997 6175 24031 6188
rect 24069 6175 24103 6188
rect 24141 6175 24175 6188
rect 24213 6175 24247 6188
rect 24285 6175 24319 6188
rect 24357 6175 24391 6188
rect 24429 6175 24463 6188
rect 24501 6175 24535 6188
rect 23781 6119 23789 6136
rect 23789 6119 23815 6136
rect 23853 6119 23857 6136
rect 23857 6119 23887 6136
rect 23781 6102 23815 6119
rect 23853 6102 23887 6119
rect 23925 6102 23959 6136
rect 23997 6119 24027 6136
rect 24027 6119 24031 6136
rect 24069 6119 24095 6136
rect 24095 6119 24103 6136
rect 24141 6119 24163 6136
rect 24163 6119 24175 6136
rect 24213 6119 24231 6136
rect 24231 6119 24247 6136
rect 24285 6119 24299 6136
rect 24299 6119 24319 6136
rect 24357 6119 24367 6136
rect 24367 6119 24391 6136
rect 24429 6119 24435 6136
rect 24435 6119 24463 6136
rect 24501 6119 24503 6136
rect 24503 6119 24535 6136
rect 23997 6102 24031 6119
rect 24069 6102 24103 6119
rect 24141 6102 24175 6119
rect 24213 6102 24247 6119
rect 24285 6102 24319 6119
rect 24357 6102 24391 6119
rect 24429 6102 24463 6119
rect 24501 6102 24535 6119
rect 23781 6050 23789 6063
rect 23789 6050 23815 6063
rect 23853 6050 23857 6063
rect 23857 6050 23887 6063
rect 23781 6029 23815 6050
rect 23853 6029 23887 6050
rect 23925 6029 23959 6063
rect 23997 6050 24027 6063
rect 24027 6050 24031 6063
rect 24069 6050 24095 6063
rect 24095 6050 24103 6063
rect 24141 6050 24163 6063
rect 24163 6050 24175 6063
rect 24213 6050 24231 6063
rect 24231 6050 24247 6063
rect 24285 6050 24299 6063
rect 24299 6050 24319 6063
rect 24357 6050 24367 6063
rect 24367 6050 24391 6063
rect 24429 6050 24435 6063
rect 24435 6050 24463 6063
rect 24501 6050 24503 6063
rect 24503 6050 24535 6063
rect 23997 6029 24031 6050
rect 24069 6029 24103 6050
rect 24141 6029 24175 6050
rect 24213 6029 24247 6050
rect 24285 6029 24319 6050
rect 24357 6029 24391 6050
rect 24429 6029 24463 6050
rect 24501 6029 24535 6050
rect 23781 5981 23789 5990
rect 23789 5981 23815 5990
rect 23853 5981 23857 5990
rect 23857 5981 23887 5990
rect 23781 5956 23815 5981
rect 23853 5956 23887 5981
rect 23925 5956 23959 5990
rect 23997 5981 24027 5990
rect 24027 5981 24031 5990
rect 24069 5981 24095 5990
rect 24095 5981 24103 5990
rect 24141 5981 24163 5990
rect 24163 5981 24175 5990
rect 24213 5981 24231 5990
rect 24231 5981 24247 5990
rect 24285 5981 24299 5990
rect 24299 5981 24319 5990
rect 24357 5981 24367 5990
rect 24367 5981 24391 5990
rect 24429 5981 24435 5990
rect 24435 5981 24463 5990
rect 24501 5981 24503 5990
rect 24503 5981 24535 5990
rect 23997 5956 24031 5981
rect 24069 5956 24103 5981
rect 24141 5956 24175 5981
rect 24213 5956 24247 5981
rect 24285 5956 24319 5981
rect 24357 5956 24391 5981
rect 24429 5956 24463 5981
rect 24501 5956 24535 5981
rect 23781 5912 23789 5917
rect 23789 5912 23815 5917
rect 23853 5912 23857 5917
rect 23857 5912 23887 5917
rect 23781 5883 23815 5912
rect 23853 5883 23887 5912
rect 23925 5883 23959 5917
rect 23997 5912 24027 5917
rect 24027 5912 24031 5917
rect 24069 5912 24095 5917
rect 24095 5912 24103 5917
rect 24141 5912 24163 5917
rect 24163 5912 24175 5917
rect 24213 5912 24231 5917
rect 24231 5912 24247 5917
rect 24285 5912 24299 5917
rect 24299 5912 24319 5917
rect 24357 5912 24367 5917
rect 24367 5912 24391 5917
rect 24429 5912 24435 5917
rect 24435 5912 24463 5917
rect 24501 5912 24503 5917
rect 24503 5912 24535 5917
rect 23997 5883 24031 5912
rect 24069 5883 24103 5912
rect 24141 5883 24175 5912
rect 24213 5883 24247 5912
rect 24285 5883 24319 5912
rect 24357 5883 24391 5912
rect 24429 5883 24463 5912
rect 24501 5883 24535 5912
rect 23781 5810 23815 5844
rect 23853 5810 23887 5844
rect 23925 5810 23959 5844
rect 23997 5810 24031 5844
rect 24069 5810 24103 5844
rect 24141 5810 24175 5844
rect 24213 5810 24247 5844
rect 24285 5810 24319 5844
rect 24357 5810 24391 5844
rect 24429 5810 24463 5844
rect 24501 5810 24535 5844
rect 23781 5737 23815 5771
rect 23853 5737 23887 5771
rect 23925 5737 23959 5771
rect 23997 5737 24031 5771
rect 24069 5737 24103 5771
rect 24141 5737 24175 5771
rect 24213 5737 24247 5771
rect 24285 5737 24319 5771
rect 24357 5737 24391 5771
rect 24429 5737 24463 5771
rect 24501 5737 24535 5771
rect 23781 5664 23815 5698
rect 23853 5664 23887 5698
rect 23925 5664 23959 5698
rect 23981 5664 24103 5698
rect 24141 5664 24175 5698
rect 24213 5664 24247 5698
rect 24285 5664 24319 5698
rect 24357 5664 24391 5698
rect 24429 5664 24463 5698
rect 24501 5664 24535 5698
rect 23981 5639 24087 5664
rect 22798 5537 22818 5571
rect 22818 5537 22832 5571
rect 22870 5537 22904 5571
rect 22942 5537 22976 5571
rect 23014 5537 23048 5571
rect 23086 5537 23120 5571
rect 23158 5537 23192 5571
rect 23230 5537 23264 5571
rect 23302 5537 23336 5571
rect 23374 5537 23408 5571
rect 23446 5537 23480 5571
rect 22798 5485 22818 5498
rect 22818 5485 22832 5498
rect 22870 5485 22904 5498
rect 22942 5485 22976 5498
rect 23014 5485 23048 5498
rect 23086 5485 23120 5498
rect 23158 5485 23192 5498
rect 23230 5485 23264 5498
rect 23302 5485 23336 5498
rect 23374 5485 23408 5498
rect 23446 5485 23480 5498
rect 22798 5464 22832 5485
rect 22870 5464 22904 5485
rect 22942 5464 22976 5485
rect 23014 5464 23048 5485
rect 23086 5464 23120 5485
rect 23158 5464 23192 5485
rect 23230 5464 23264 5485
rect 23302 5464 23336 5485
rect 23374 5464 23408 5485
rect 23446 5464 23480 5485
rect 23981 5532 24087 5639
rect 22798 5391 22832 5425
rect 22870 5391 22904 5425
rect 22942 5391 22944 5425
rect 22944 5391 22976 5425
rect 23014 5391 23048 5425
rect 23086 5406 23117 5425
rect 23117 5406 23120 5425
rect 23158 5406 23186 5425
rect 23186 5406 23192 5425
rect 23230 5406 23255 5425
rect 23255 5406 23264 5425
rect 23302 5406 23324 5425
rect 23324 5406 23336 5425
rect 23374 5406 23393 5425
rect 23393 5406 23408 5425
rect 23446 5406 23462 5425
rect 23462 5406 23480 5425
rect 23086 5391 23120 5406
rect 23158 5391 23192 5406
rect 23230 5391 23264 5406
rect 23302 5391 23336 5406
rect 23374 5391 23408 5406
rect 23446 5391 23480 5406
rect 22798 5318 22832 5352
rect 22870 5318 22904 5352
rect 22942 5318 22944 5352
rect 22944 5318 22976 5352
rect 23014 5318 23048 5352
rect 23086 5338 23117 5352
rect 23117 5338 23120 5352
rect 23158 5338 23186 5352
rect 23186 5338 23192 5352
rect 23230 5338 23255 5352
rect 23255 5338 23264 5352
rect 23302 5338 23324 5352
rect 23324 5338 23336 5352
rect 23374 5338 23393 5352
rect 23393 5338 23408 5352
rect 23446 5338 23462 5352
rect 23462 5338 23480 5352
rect 23086 5318 23120 5338
rect 23158 5318 23192 5338
rect 23230 5318 23264 5338
rect 23302 5318 23336 5338
rect 23374 5318 23408 5338
rect 23446 5318 23480 5338
rect 22782 5246 22816 5280
rect 22855 5246 22889 5280
rect 22928 5246 22944 5280
rect 22944 5246 22962 5280
rect 23001 5270 23013 5280
rect 23013 5270 23035 5280
rect 23074 5270 23082 5280
rect 23082 5270 23108 5280
rect 23147 5270 23151 5280
rect 23151 5270 23181 5280
rect 23001 5246 23035 5270
rect 23074 5246 23108 5270
rect 23147 5246 23181 5270
rect 23220 5246 23254 5280
rect 23294 5270 23324 5280
rect 23324 5270 23328 5280
rect 23368 5270 23393 5280
rect 23393 5270 23402 5280
rect 23442 5270 23462 5280
rect 23462 5270 23476 5280
rect 23516 5270 23531 5280
rect 23531 5270 23550 5280
rect 23593 5270 23600 5274
rect 23600 5270 23627 5274
rect 23665 5270 23669 5274
rect 23669 5270 23699 5274
rect 23737 5270 23738 5274
rect 23738 5270 23771 5274
rect 23294 5246 23328 5270
rect 23368 5246 23402 5270
rect 23442 5246 23476 5270
rect 23516 5246 23550 5270
rect 23593 5240 23627 5270
rect 23665 5240 23699 5270
rect 23737 5240 23771 5270
rect 22782 5174 22816 5208
rect 22855 5174 22889 5208
rect 22928 5174 22944 5208
rect 22944 5174 22962 5208
rect 23001 5202 23013 5208
rect 23013 5202 23035 5208
rect 23074 5202 23082 5208
rect 23082 5202 23108 5208
rect 23147 5202 23151 5208
rect 23151 5202 23181 5208
rect 23001 5174 23035 5202
rect 23074 5174 23108 5202
rect 23147 5174 23181 5202
rect 23220 5174 23254 5208
rect 23294 5202 23324 5208
rect 23324 5202 23328 5208
rect 23368 5202 23393 5208
rect 23393 5202 23402 5208
rect 23442 5202 23462 5208
rect 23462 5202 23476 5208
rect 23516 5202 23531 5208
rect 23531 5202 23550 5208
rect 23294 5174 23328 5202
rect 23368 5174 23402 5202
rect 23442 5174 23476 5202
rect 23516 5174 23550 5202
rect 23593 5168 23627 5201
rect 23665 5168 23699 5201
rect 23737 5168 23771 5201
rect 22782 5102 22816 5136
rect 22855 5102 22889 5136
rect 22928 5102 22944 5136
rect 22944 5102 22962 5136
rect 23001 5134 23013 5136
rect 23013 5134 23035 5136
rect 23074 5134 23082 5136
rect 23082 5134 23108 5136
rect 23147 5134 23151 5136
rect 23151 5134 23181 5136
rect 23001 5102 23035 5134
rect 23074 5102 23108 5134
rect 23147 5102 23181 5134
rect 23220 5102 23254 5136
rect 23593 5167 23600 5168
rect 23600 5167 23627 5168
rect 23665 5167 23669 5168
rect 23669 5167 23699 5168
rect 23737 5167 23738 5168
rect 23738 5167 23771 5168
rect 23294 5134 23324 5136
rect 23324 5134 23328 5136
rect 23368 5134 23393 5136
rect 23393 5134 23402 5136
rect 23442 5134 23462 5136
rect 23462 5134 23476 5136
rect 23516 5134 23531 5136
rect 23531 5134 23550 5136
rect 23294 5102 23328 5134
rect 23368 5102 23402 5134
rect 23442 5102 23476 5134
rect 23516 5102 23550 5134
rect 23593 5100 23627 5128
rect 23665 5100 23699 5128
rect 23737 5100 23771 5128
rect 23593 5094 23600 5100
rect 23600 5094 23627 5100
rect 23665 5094 23669 5100
rect 23669 5094 23699 5100
rect 23737 5094 23738 5100
rect 23738 5094 23771 5100
rect 22782 5030 22816 5064
rect 22855 5030 22889 5064
rect 22928 5030 22944 5064
rect 22944 5030 22962 5064
rect 23001 5032 23035 5064
rect 23074 5032 23108 5064
rect 23147 5032 23181 5064
rect 23001 5030 23013 5032
rect 23013 5030 23035 5032
rect 23074 5030 23082 5032
rect 23082 5030 23108 5032
rect 23147 5030 23151 5032
rect 23151 5030 23181 5032
rect 23220 5030 23254 5064
rect 23294 5032 23328 5064
rect 23368 5032 23402 5064
rect 23442 5032 23476 5064
rect 23516 5032 23550 5064
rect 23593 5032 23627 5055
rect 23665 5032 23699 5055
rect 23737 5032 23771 5055
rect 23294 5030 23324 5032
rect 23324 5030 23328 5032
rect 23368 5030 23393 5032
rect 23393 5030 23402 5032
rect 23442 5030 23462 5032
rect 23462 5030 23476 5032
rect 23516 5030 23531 5032
rect 23531 5030 23550 5032
rect 23593 5021 23600 5032
rect 23600 5021 23627 5032
rect 23665 5021 23669 5032
rect 23669 5021 23699 5032
rect 23737 5021 23738 5032
rect 23738 5021 23771 5032
rect 22782 4958 22816 4992
rect 22855 4958 22889 4992
rect 22928 4958 22944 4992
rect 22944 4958 22962 4992
rect 23001 4964 23035 4992
rect 23074 4964 23108 4992
rect 23147 4964 23181 4992
rect 23001 4958 23013 4964
rect 23013 4958 23035 4964
rect 23074 4958 23082 4964
rect 23082 4958 23108 4964
rect 23147 4958 23151 4964
rect 23151 4958 23181 4964
rect 23220 4958 23254 4992
rect 23294 4964 23328 4992
rect 23368 4964 23402 4992
rect 23442 4964 23476 4992
rect 23516 4964 23550 4992
rect 23593 4964 23627 4982
rect 23665 4964 23699 4982
rect 23737 4964 23771 4982
rect 23294 4958 23324 4964
rect 23324 4958 23328 4964
rect 23368 4958 23393 4964
rect 23393 4958 23402 4964
rect 23442 4958 23462 4964
rect 23462 4958 23476 4964
rect 23516 4958 23531 4964
rect 23531 4958 23550 4964
rect 23593 4948 23600 4964
rect 23600 4948 23627 4964
rect 23665 4948 23669 4964
rect 23669 4948 23699 4964
rect 23737 4948 23738 4964
rect 23738 4948 23771 4964
rect 23593 4896 23627 4909
rect 23665 4896 23699 4909
rect 23737 4896 23771 4909
rect 23593 4875 23600 4896
rect 23600 4875 23627 4896
rect 23665 4875 23669 4896
rect 23669 4875 23699 4896
rect 23737 4875 23738 4896
rect 23738 4875 23771 4896
rect 23593 4828 23627 4836
rect 23665 4828 23699 4836
rect 23737 4828 23771 4836
rect 23593 4802 23600 4828
rect 23600 4802 23627 4828
rect 23665 4802 23669 4828
rect 23669 4802 23699 4828
rect 23737 4802 23738 4828
rect 23738 4802 23771 4828
rect 728 4737 762 4746
rect 800 4737 834 4746
rect 728 4712 730 4737
rect 730 4712 762 4737
rect 800 4712 832 4737
rect 832 4712 834 4737
rect 728 4665 762 4673
rect 800 4665 834 4672
rect 728 4639 730 4665
rect 730 4639 762 4665
rect 800 4638 832 4665
rect 832 4638 834 4665
rect 728 4593 762 4600
rect 800 4593 834 4598
rect 728 4566 730 4593
rect 730 4566 762 4593
rect 800 4564 832 4593
rect 832 4564 834 4593
rect 23593 4737 23627 4763
rect 23665 4737 23699 4763
rect 23737 4737 23771 4763
rect 23593 4729 23597 4737
rect 23597 4729 23627 4737
rect 23665 4729 23699 4737
rect 23737 4729 23767 4737
rect 23767 4729 23771 4737
rect 23593 4668 23627 4690
rect 23665 4668 23699 4690
rect 23737 4668 23771 4690
rect 23593 4656 23597 4668
rect 23597 4656 23627 4668
rect 23665 4656 23699 4668
rect 23737 4656 23767 4668
rect 23767 4656 23771 4668
rect 23593 4599 23627 4617
rect 23665 4599 23699 4617
rect 23737 4599 23771 4617
rect 23593 4583 23597 4599
rect 23597 4583 23627 4599
rect 728 4521 762 4527
rect 800 4521 834 4524
rect 310 4449 312 4479
rect 312 4449 346 4479
rect 346 4449 380 4479
rect 380 4449 414 4479
rect 414 4449 416 4479
rect 310 4413 416 4449
rect 310 4379 312 4413
rect 312 4379 346 4413
rect 346 4379 380 4413
rect 380 4379 414 4413
rect 414 4379 416 4413
rect 310 4343 416 4379
rect 310 4309 312 4343
rect 312 4309 346 4343
rect 346 4309 380 4343
rect 380 4309 414 4343
rect 414 4309 416 4343
rect 310 4273 416 4309
rect 310 4239 312 4273
rect 312 4239 346 4273
rect 346 4239 380 4273
rect 380 4239 414 4273
rect 414 4239 416 4273
rect 310 4203 416 4239
rect 310 4169 312 4203
rect 312 4169 346 4203
rect 346 4169 380 4203
rect 380 4169 414 4203
rect 414 4169 416 4203
rect 310 4134 416 4169
rect 310 4100 312 4134
rect 312 4100 346 4134
rect 346 4100 380 4134
rect 380 4100 414 4134
rect 414 4100 416 4134
rect 310 4065 416 4100
rect 310 4031 312 4065
rect 312 4031 346 4065
rect 346 4031 380 4065
rect 380 4031 414 4065
rect 414 4031 416 4065
rect 310 3996 416 4031
rect 310 3962 312 3996
rect 312 3962 346 3996
rect 346 3962 380 3996
rect 380 3962 414 3996
rect 414 3962 416 3996
rect 310 3927 416 3962
rect 310 3893 312 3927
rect 312 3893 346 3927
rect 346 3893 380 3927
rect 380 3893 414 3927
rect 414 3893 416 3927
rect 310 3858 416 3893
rect 310 3824 312 3858
rect 312 3824 346 3858
rect 346 3824 380 3858
rect 380 3824 414 3858
rect 414 3824 416 3858
rect 310 3789 416 3824
rect 310 3755 312 3789
rect 312 3755 346 3789
rect 346 3755 380 3789
rect 380 3755 414 3789
rect 414 3755 416 3789
rect 310 3720 416 3755
rect 310 3686 312 3720
rect 312 3686 346 3720
rect 346 3686 380 3720
rect 380 3686 414 3720
rect 414 3686 416 3720
rect 310 3651 416 3686
rect 310 3617 312 3651
rect 312 3617 346 3651
rect 346 3617 380 3651
rect 380 3617 414 3651
rect 414 3617 416 3651
rect 310 3582 416 3617
rect 310 3548 312 3582
rect 312 3548 346 3582
rect 346 3548 380 3582
rect 380 3548 414 3582
rect 414 3548 416 3582
rect 310 3513 416 3548
rect 310 3479 312 3513
rect 312 3479 346 3513
rect 346 3479 380 3513
rect 380 3479 414 3513
rect 414 3479 416 3513
rect 310 3444 416 3479
rect 310 3410 312 3444
rect 312 3410 346 3444
rect 346 3410 380 3444
rect 380 3410 414 3444
rect 414 3410 416 3444
rect 310 3375 416 3410
rect 310 3341 312 3375
rect 312 3341 346 3375
rect 346 3341 380 3375
rect 380 3341 414 3375
rect 414 3341 416 3375
rect 310 3306 416 3341
rect 310 3272 312 3306
rect 312 3272 346 3306
rect 346 3272 380 3306
rect 380 3272 414 3306
rect 414 3272 416 3306
rect 310 3237 416 3272
rect 310 3203 312 3237
rect 312 3203 346 3237
rect 346 3203 380 3237
rect 380 3203 414 3237
rect 414 3203 416 3237
rect 310 3168 416 3203
rect 310 3134 312 3168
rect 312 3134 346 3168
rect 346 3134 380 3168
rect 380 3134 414 3168
rect 414 3134 416 3168
rect 310 3099 416 3134
rect 310 3065 312 3099
rect 312 3065 346 3099
rect 346 3065 380 3099
rect 380 3065 414 3099
rect 414 3065 416 3099
rect 310 3030 416 3065
rect 310 2996 312 3030
rect 312 2996 346 3030
rect 346 2996 380 3030
rect 380 2996 414 3030
rect 414 2996 416 3030
rect 310 2961 416 2996
rect 310 2927 312 2961
rect 312 2927 346 2961
rect 346 2927 380 2961
rect 380 2927 414 2961
rect 414 2927 416 2961
rect 310 2892 416 2927
rect 310 2858 312 2892
rect 312 2858 346 2892
rect 346 2858 380 2892
rect 380 2858 414 2892
rect 414 2858 416 2892
rect 310 2823 416 2858
rect 310 2789 312 2823
rect 312 2789 346 2823
rect 346 2789 380 2823
rect 380 2789 414 2823
rect 414 2789 416 2823
rect 310 2754 416 2789
rect 310 2720 312 2754
rect 312 2720 346 2754
rect 346 2720 380 2754
rect 380 2720 414 2754
rect 414 2720 416 2754
rect 310 2685 416 2720
rect 310 2651 312 2685
rect 312 2651 346 2685
rect 346 2651 380 2685
rect 380 2651 414 2685
rect 414 2651 416 2685
rect 310 2616 416 2651
rect 310 2582 312 2616
rect 312 2582 346 2616
rect 346 2582 380 2616
rect 380 2582 414 2616
rect 414 2582 416 2616
rect 310 2573 416 2582
rect 310 2513 312 2534
rect 312 2513 344 2534
rect 382 2513 414 2534
rect 414 2513 416 2534
rect 310 2500 344 2513
rect 382 2500 416 2513
rect 310 2444 312 2461
rect 312 2444 344 2461
rect 382 2444 414 2461
rect 414 2444 416 2461
rect 310 2427 344 2444
rect 382 2427 416 2444
rect 310 2375 312 2388
rect 312 2375 344 2388
rect 382 2375 414 2388
rect 414 2375 416 2388
rect 310 2354 344 2375
rect 382 2354 416 2375
rect 310 2306 312 2315
rect 312 2306 344 2315
rect 382 2306 414 2315
rect 414 2306 416 2315
rect 310 2281 344 2306
rect 382 2281 416 2306
rect 310 2237 312 2242
rect 312 2237 344 2242
rect 382 2237 414 2242
rect 414 2237 416 2242
rect 310 2208 344 2237
rect 382 2208 416 2237
rect 310 2168 312 2169
rect 312 2168 344 2169
rect 382 2168 414 2169
rect 414 2168 416 2169
rect 310 2135 344 2168
rect 382 2135 416 2168
rect 310 2064 344 2096
rect 382 2064 416 2096
rect 310 2062 312 2064
rect 312 2062 344 2064
rect 382 2062 414 2064
rect 414 2062 416 2064
rect 310 1995 344 2023
rect 382 1995 416 2023
rect 310 1989 312 1995
rect 312 1989 344 1995
rect 382 1989 414 1995
rect 414 1989 416 1995
rect 310 1926 344 1950
rect 382 1926 416 1950
rect 310 1916 312 1926
rect 312 1916 344 1926
rect 382 1916 414 1926
rect 414 1916 416 1926
rect 310 1857 344 1877
rect 382 1857 416 1877
rect 310 1843 312 1857
rect 312 1843 344 1857
rect 382 1843 414 1857
rect 414 1843 416 1857
rect 310 1788 344 1804
rect 382 1788 416 1804
rect 310 1770 312 1788
rect 312 1770 344 1788
rect 382 1770 414 1788
rect 414 1770 416 1788
rect 310 1719 344 1731
rect 382 1719 416 1731
rect 310 1697 312 1719
rect 312 1697 344 1719
rect 382 1697 414 1719
rect 414 1697 416 1719
rect 310 1650 344 1658
rect 382 1650 416 1658
rect 310 1624 312 1650
rect 312 1624 344 1650
rect 382 1624 414 1650
rect 414 1624 416 1650
rect 310 1581 344 1585
rect 382 1581 416 1585
rect 310 1551 312 1581
rect 312 1551 344 1581
rect 382 1551 414 1581
rect 414 1551 416 1581
rect 310 1478 312 1512
rect 312 1478 344 1512
rect 382 1478 414 1512
rect 414 1478 416 1512
rect 310 1409 312 1439
rect 312 1409 344 1439
rect 382 1409 414 1439
rect 414 1409 416 1439
rect 310 1405 344 1409
rect 382 1405 416 1409
rect 310 1340 312 1366
rect 312 1340 344 1366
rect 382 1340 414 1366
rect 414 1340 416 1366
rect 310 1332 344 1340
rect 382 1332 416 1340
rect 310 1271 312 1293
rect 312 1271 344 1293
rect 382 1271 414 1293
rect 414 1271 416 1293
rect 310 1259 344 1271
rect 382 1259 416 1271
rect 310 1202 312 1220
rect 312 1202 344 1220
rect 382 1202 414 1220
rect 414 1202 416 1220
rect 310 1186 344 1202
rect 382 1186 416 1202
rect 310 1133 312 1147
rect 312 1133 344 1147
rect 382 1133 414 1147
rect 414 1133 416 1147
rect 310 1113 344 1133
rect 382 1113 416 1133
rect 310 1064 312 1074
rect 312 1064 344 1074
rect 382 1064 414 1074
rect 414 1064 416 1074
rect 310 1040 344 1064
rect 382 1040 416 1064
rect 310 995 312 1001
rect 312 995 344 1001
rect 382 995 414 1001
rect 414 995 416 1001
rect 310 967 344 995
rect 382 967 416 995
rect 310 926 312 928
rect 312 926 344 928
rect 382 926 414 928
rect 414 926 416 928
rect 310 894 344 926
rect 382 894 416 926
rect 728 4493 730 4521
rect 730 4493 762 4521
rect 800 4490 832 4521
rect 832 4490 834 4521
rect 728 4449 762 4454
rect 800 4449 834 4450
rect 728 4420 730 4449
rect 730 4420 762 4449
rect 800 4416 832 4449
rect 832 4416 834 4449
rect 728 4377 762 4381
rect 728 4347 730 4377
rect 730 4347 762 4377
rect 800 4343 832 4376
rect 832 4343 834 4376
rect 800 4342 834 4343
rect 728 4305 762 4308
rect 728 4274 730 4305
rect 730 4274 762 4305
rect 800 4271 832 4302
rect 832 4271 834 4302
rect 800 4268 834 4271
rect 728 4233 762 4235
rect 728 4201 730 4233
rect 730 4201 762 4233
rect 800 4199 832 4228
rect 832 4199 834 4228
rect 800 4194 834 4199
rect 728 4161 762 4162
rect 728 4128 730 4161
rect 730 4128 762 4161
rect 800 4127 832 4154
rect 832 4127 834 4154
rect 800 4120 834 4127
rect 728 4055 730 4089
rect 730 4055 762 4089
rect 800 4055 832 4080
rect 832 4055 834 4080
rect 800 4046 834 4055
rect 728 3983 730 4016
rect 730 3983 762 4016
rect 800 3983 832 4006
rect 832 3983 834 4006
rect 728 3982 762 3983
rect 800 3972 834 3983
rect 728 3912 730 3943
rect 730 3912 762 3943
rect 800 3912 832 3932
rect 832 3912 834 3932
rect 728 3909 762 3912
rect 800 3898 834 3912
rect 728 3841 730 3870
rect 730 3841 762 3870
rect 800 3841 832 3858
rect 832 3841 834 3858
rect 728 3836 762 3841
rect 800 3824 834 3841
rect 728 3770 730 3797
rect 730 3770 762 3797
rect 800 3770 832 3784
rect 832 3770 834 3784
rect 728 3763 762 3770
rect 800 3750 834 3770
rect 728 3699 730 3724
rect 730 3699 762 3724
rect 800 3699 832 3710
rect 832 3699 834 3710
rect 728 3690 762 3699
rect 800 3676 834 3699
rect 728 3628 730 3651
rect 730 3628 762 3651
rect 800 3628 832 3636
rect 832 3628 834 3636
rect 728 3617 762 3628
rect 800 3602 834 3628
rect 728 3557 730 3578
rect 730 3557 762 3578
rect 800 3557 832 3562
rect 832 3557 834 3562
rect 728 3544 762 3557
rect 800 3528 834 3557
rect 728 3486 730 3505
rect 730 3486 762 3505
rect 800 3486 832 3488
rect 832 3486 834 3488
rect 728 3471 762 3486
rect 800 3454 834 3486
rect 728 3415 730 3432
rect 730 3415 762 3432
rect 728 3398 762 3415
rect 800 3380 834 3414
rect 728 3344 730 3359
rect 730 3344 762 3359
rect 728 3325 762 3344
rect 800 3307 834 3341
rect 728 3252 730 3286
rect 730 3252 762 3286
rect 800 3252 832 3268
rect 832 3252 834 3268
rect 800 3234 834 3252
rect 728 3182 730 3213
rect 730 3182 762 3213
rect 800 3183 832 3195
rect 832 3183 834 3195
rect 728 3179 762 3182
rect 800 3161 834 3183
rect 728 3112 730 3140
rect 730 3112 762 3140
rect 800 3114 832 3122
rect 832 3114 834 3122
rect 728 3106 762 3112
rect 800 3088 834 3114
rect 728 3042 730 3067
rect 730 3042 762 3067
rect 800 3045 832 3049
rect 832 3045 834 3049
rect 728 3033 762 3042
rect 800 3015 834 3045
rect 728 2972 730 2994
rect 730 2972 762 2994
rect 728 2960 762 2972
rect 800 2942 834 2976
rect 728 2903 730 2921
rect 730 2903 762 2921
rect 728 2887 762 2903
rect 800 2869 834 2903
rect 728 2834 730 2848
rect 730 2834 762 2848
rect 728 2814 762 2834
rect 800 2796 834 2830
rect 728 2765 730 2775
rect 730 2765 762 2775
rect 728 2741 762 2765
rect 800 2723 834 2757
rect 728 2696 730 2702
rect 730 2696 762 2702
rect 728 2668 762 2696
rect 800 2650 834 2684
rect 728 2627 730 2629
rect 730 2627 762 2629
rect 728 2595 762 2627
rect 800 2577 834 2611
rect 728 2523 762 2556
rect 728 2522 730 2523
rect 730 2522 762 2523
rect 800 2504 834 2538
rect 728 2454 762 2483
rect 728 2449 730 2454
rect 730 2449 762 2454
rect 800 2431 834 2465
rect 728 2385 762 2411
rect 728 2377 730 2385
rect 730 2377 762 2385
rect 800 2358 834 2392
rect 728 2316 762 2339
rect 728 2305 730 2316
rect 730 2305 762 2316
rect 800 2285 834 2319
rect 728 2247 762 2267
rect 728 2233 730 2247
rect 730 2233 762 2247
rect 800 2212 834 2246
rect 728 2178 762 2195
rect 728 2161 730 2178
rect 730 2161 762 2178
rect 800 2139 834 2173
rect 728 2109 762 2123
rect 728 2089 730 2109
rect 730 2089 762 2109
rect 800 2066 834 2100
rect 728 2040 762 2051
rect 728 2017 730 2040
rect 730 2017 762 2040
rect 800 1993 834 2027
rect 728 1971 762 1979
rect 728 1945 730 1971
rect 730 1945 762 1971
rect 800 1920 834 1954
rect 728 1902 762 1907
rect 728 1873 730 1902
rect 730 1873 762 1902
rect 800 1847 834 1881
rect 728 1833 762 1835
rect 728 1801 730 1833
rect 730 1801 762 1833
rect 800 1774 834 1808
rect 728 1730 730 1763
rect 730 1730 762 1763
rect 728 1729 762 1730
rect 800 1701 834 1735
rect 728 1661 730 1691
rect 730 1661 762 1691
rect 728 1657 762 1661
rect 800 1628 834 1662
rect 728 1592 730 1619
rect 730 1592 762 1619
rect 728 1585 762 1592
rect 800 1555 834 1589
rect 728 1523 730 1547
rect 730 1523 762 1547
rect 728 1513 762 1523
rect 800 1482 834 1516
rect 728 1454 730 1475
rect 730 1454 762 1475
rect 728 1441 762 1454
rect 800 1409 834 1443
rect 728 1385 730 1403
rect 730 1385 762 1403
rect 728 1369 762 1385
rect 800 1336 834 1370
rect 728 1316 730 1331
rect 730 1316 762 1331
rect 728 1297 762 1316
rect 1169 4447 1188 4479
rect 1188 4447 1203 4479
rect 1241 4447 1256 4479
rect 1256 4447 1275 4479
rect 1313 4447 1324 4479
rect 1324 4447 1347 4479
rect 1385 4447 1392 4479
rect 1392 4447 1419 4479
rect 1457 4447 1460 4479
rect 1460 4447 1491 4479
rect 1529 4471 1563 4479
rect 1601 4472 1635 4479
rect 1169 4445 1203 4447
rect 1241 4445 1275 4447
rect 1313 4445 1347 4447
rect 1385 4445 1419 4447
rect 1457 4445 1491 4447
rect 1529 4445 1541 4471
rect 1541 4445 1563 4471
rect 1601 4445 1635 4472
rect 1687 4451 1721 4485
rect 1760 4451 1794 4485
rect 1833 4451 1867 4485
rect 1906 4451 1940 4485
rect 1979 4451 2013 4485
rect 2052 4451 2086 4485
rect 2125 4451 2159 4485
rect 2198 4451 2232 4485
rect 2271 4451 2305 4485
rect 2344 4451 2378 4485
rect 2417 4451 2451 4485
rect 2490 4451 2524 4485
rect 2562 4451 2596 4485
rect 2634 4451 2668 4485
rect 2706 4451 2740 4485
rect 2778 4451 2812 4485
rect 2850 4451 2884 4485
rect 2922 4451 2956 4485
rect 2994 4451 3028 4485
rect 3066 4451 3100 4485
rect 3138 4451 3172 4485
rect 3210 4451 3244 4485
rect 3282 4451 3316 4485
rect 3354 4451 3388 4485
rect 3426 4451 3460 4485
rect 3498 4451 3532 4485
rect 3570 4451 3604 4485
rect 3642 4451 3676 4485
rect 3714 4451 3748 4485
rect 3786 4451 3820 4485
rect 3858 4451 3892 4485
rect 3930 4451 3964 4485
rect 4002 4451 4036 4485
rect 4074 4451 4108 4485
rect 4146 4451 4180 4485
rect 4218 4451 4252 4485
rect 4290 4451 4324 4485
rect 4362 4451 4396 4485
rect 4434 4451 4468 4485
rect 4506 4451 4540 4485
rect 4578 4451 4612 4485
rect 4650 4451 4684 4485
rect 4722 4451 4756 4485
rect 4794 4451 4828 4485
rect 4866 4451 4900 4485
rect 4938 4451 4972 4485
rect 5010 4451 5044 4485
rect 5082 4451 5116 4485
rect 5154 4451 5188 4485
rect 5226 4451 5260 4485
rect 5298 4451 5332 4485
rect 5370 4451 5404 4485
rect 5442 4451 5476 4485
rect 5514 4451 5548 4485
rect 5586 4451 5620 4485
rect 5658 4451 5692 4485
rect 5730 4451 5764 4485
rect 5802 4451 5836 4485
rect 5874 4451 5908 4485
rect 5946 4451 5980 4485
rect 6018 4451 6052 4485
rect 6090 4451 6124 4485
rect 6162 4451 6196 4485
rect 6234 4451 6268 4485
rect 6306 4451 6340 4485
rect 6378 4451 6412 4485
rect 6450 4451 6484 4485
rect 6522 4451 6556 4485
rect 6594 4451 6628 4485
rect 6666 4451 6700 4485
rect 6738 4451 6772 4485
rect 6810 4451 6844 4485
rect 6882 4451 6916 4485
rect 6954 4451 6988 4485
rect 7026 4451 7060 4485
rect 7098 4451 7132 4485
rect 7170 4451 7204 4485
rect 7242 4451 7276 4485
rect 7314 4451 7348 4485
rect 7386 4451 7420 4485
rect 7458 4451 7492 4485
rect 7530 4451 7564 4485
rect 7602 4451 7636 4485
rect 7674 4451 7708 4485
rect 7746 4451 7780 4485
rect 7818 4451 7852 4485
rect 7890 4451 7924 4485
rect 7962 4451 7996 4485
rect 8034 4451 8068 4485
rect 8106 4451 8140 4485
rect 8178 4451 8212 4485
rect 8250 4451 8284 4485
rect 8322 4451 8356 4485
rect 8394 4451 8428 4485
rect 8466 4451 8500 4485
rect 8538 4451 8572 4485
rect 8610 4451 8644 4485
rect 8682 4451 8716 4485
rect 8754 4472 8785 4485
rect 8785 4472 8788 4485
rect 8826 4472 8854 4485
rect 8854 4472 8860 4485
rect 8898 4472 8923 4485
rect 8923 4472 8932 4485
rect 8970 4472 8992 4485
rect 8992 4472 9004 4485
rect 9042 4472 9061 4485
rect 9061 4472 9076 4485
rect 9114 4472 9130 4485
rect 9130 4472 9148 4485
rect 9186 4472 9199 4485
rect 9199 4472 9220 4485
rect 9258 4472 9268 4485
rect 9268 4472 9292 4485
rect 9330 4472 9337 4485
rect 9337 4472 9364 4485
rect 9402 4472 9406 4485
rect 9406 4472 9436 4485
rect 9474 4472 9475 4485
rect 9475 4472 9508 4485
rect 23665 4583 23699 4599
rect 23737 4583 23767 4599
rect 23767 4583 23771 4599
rect 23593 4530 23627 4544
rect 23665 4530 23699 4544
rect 23737 4530 23771 4544
rect 23593 4510 23597 4530
rect 23597 4510 23627 4530
rect 23665 4510 23699 4530
rect 23737 4510 23767 4530
rect 23767 4510 23771 4530
rect 9546 4472 9578 4485
rect 9578 4472 9580 4485
rect 9618 4472 9647 4485
rect 9647 4472 9652 4485
rect 9690 4472 9716 4485
rect 9716 4472 9724 4485
rect 9762 4472 9785 4485
rect 9785 4472 9796 4485
rect 9834 4472 9854 4485
rect 9854 4472 9868 4485
rect 9906 4472 9923 4485
rect 9923 4472 9940 4485
rect 9978 4472 9992 4485
rect 9992 4472 10012 4485
rect 8754 4451 8788 4472
rect 8826 4451 8860 4472
rect 8898 4451 8932 4472
rect 8970 4451 9004 4472
rect 9042 4451 9076 4472
rect 9114 4451 9148 4472
rect 9186 4451 9220 4472
rect 9258 4451 9292 4472
rect 9330 4451 9364 4472
rect 9402 4451 9436 4472
rect 9474 4451 9508 4472
rect 9546 4451 9580 4472
rect 9618 4451 9652 4472
rect 9690 4451 9724 4472
rect 9762 4451 9796 4472
rect 9834 4451 9868 4472
rect 9906 4451 9940 4472
rect 9978 4451 10012 4472
rect 10050 4451 10084 4485
rect 10122 4451 10156 4485
rect 10194 4451 10228 4485
rect 10266 4451 10300 4485
rect 10338 4451 10372 4485
rect 10410 4451 10444 4485
rect 10482 4451 10516 4485
rect 10554 4451 10588 4485
rect 10626 4451 10660 4485
rect 10698 4451 10732 4485
rect 10770 4451 10804 4485
rect 10842 4451 10876 4485
rect 1169 4378 1188 4405
rect 1188 4378 1203 4405
rect 1241 4378 1256 4405
rect 1256 4378 1275 4405
rect 1313 4378 1324 4405
rect 1324 4378 1347 4405
rect 1385 4378 1392 4405
rect 1392 4378 1419 4405
rect 1457 4378 1460 4405
rect 1460 4378 1491 4405
rect 1529 4402 1563 4405
rect 1601 4402 1609 4405
rect 1609 4402 1635 4405
rect 23593 4461 23627 4471
rect 23665 4461 23699 4471
rect 23737 4461 23771 4471
rect 23593 4437 23597 4461
rect 23597 4437 23627 4461
rect 23665 4437 23699 4461
rect 23737 4437 23767 4461
rect 23767 4437 23771 4461
rect 1169 4371 1203 4378
rect 1241 4371 1275 4378
rect 1313 4371 1347 4378
rect 1385 4371 1419 4378
rect 1457 4371 1491 4378
rect 1529 4371 1541 4402
rect 1541 4371 1563 4402
rect 1601 4371 1635 4402
rect 1169 4309 1188 4331
rect 1188 4309 1203 4331
rect 1241 4309 1256 4331
rect 1256 4309 1275 4331
rect 1313 4309 1324 4331
rect 1324 4309 1347 4331
rect 1385 4309 1392 4331
rect 1392 4309 1419 4331
rect 1457 4309 1460 4331
rect 1460 4309 1491 4331
rect 1169 4297 1203 4309
rect 1241 4297 1275 4309
rect 1313 4297 1347 4309
rect 1385 4297 1419 4309
rect 1457 4297 1491 4309
rect 1529 4299 1541 4331
rect 1541 4299 1563 4331
rect 1529 4297 1563 4299
rect 1601 4297 1635 4331
rect 1169 4240 1188 4257
rect 1188 4240 1203 4257
rect 1241 4240 1256 4257
rect 1256 4240 1275 4257
rect 1313 4240 1324 4257
rect 1324 4240 1347 4257
rect 1385 4240 1392 4257
rect 1392 4240 1419 4257
rect 1457 4240 1460 4257
rect 1460 4240 1491 4257
rect 1169 4223 1203 4240
rect 1241 4223 1275 4240
rect 1313 4223 1347 4240
rect 1385 4223 1419 4240
rect 1457 4223 1491 4240
rect 1529 4230 1541 4257
rect 1541 4230 1563 4257
rect 1529 4223 1563 4230
rect 1601 4226 1635 4257
rect 1601 4223 1609 4226
rect 1609 4223 1635 4226
rect 1169 4171 1188 4183
rect 1188 4171 1203 4183
rect 1241 4171 1256 4183
rect 1256 4171 1275 4183
rect 1313 4171 1324 4183
rect 1324 4171 1347 4183
rect 1385 4171 1392 4183
rect 1392 4171 1419 4183
rect 1457 4171 1460 4183
rect 1460 4171 1491 4183
rect 1169 4149 1203 4171
rect 1241 4149 1275 4171
rect 1313 4149 1347 4171
rect 1385 4149 1419 4171
rect 1457 4149 1491 4171
rect 1529 4161 1541 4183
rect 1541 4161 1563 4183
rect 1529 4149 1563 4161
rect 1601 4156 1635 4183
rect 1601 4149 1609 4156
rect 1609 4149 1635 4156
rect 1169 4102 1188 4109
rect 1188 4102 1203 4109
rect 1241 4102 1256 4109
rect 1256 4102 1275 4109
rect 1313 4102 1324 4109
rect 1324 4102 1347 4109
rect 1385 4102 1392 4109
rect 1392 4102 1419 4109
rect 1457 4102 1460 4109
rect 1460 4102 1491 4109
rect 1169 4075 1203 4102
rect 1241 4075 1275 4102
rect 1313 4075 1347 4102
rect 1385 4075 1419 4102
rect 1457 4075 1491 4102
rect 1529 4092 1541 4109
rect 1541 4092 1563 4109
rect 1529 4075 1563 4092
rect 1601 4086 1635 4109
rect 1601 4075 1609 4086
rect 1609 4075 1635 4086
rect 1169 4033 1188 4035
rect 1188 4033 1203 4035
rect 1241 4033 1256 4035
rect 1256 4033 1275 4035
rect 1313 4033 1324 4035
rect 1324 4033 1347 4035
rect 1385 4033 1392 4035
rect 1392 4033 1419 4035
rect 1457 4033 1460 4035
rect 1460 4033 1491 4035
rect 1169 4001 1203 4033
rect 1241 4001 1275 4033
rect 1313 4001 1347 4033
rect 1385 4001 1419 4033
rect 1457 4001 1491 4033
rect 1529 4023 1541 4035
rect 1541 4023 1563 4035
rect 1529 4001 1563 4023
rect 1601 4016 1635 4035
rect 1601 4001 1609 4016
rect 1609 4001 1635 4016
rect 3946 4026 3978 4060
rect 3978 4026 3980 4060
rect 4018 4026 4046 4060
rect 4046 4026 4052 4060
rect 1169 3929 1203 3962
rect 1241 3929 1275 3962
rect 1313 3929 1347 3962
rect 1385 3929 1419 3962
rect 1457 3929 1491 3962
rect 1529 3954 1541 3962
rect 1541 3954 1563 3962
rect 1169 3928 1188 3929
rect 1188 3928 1203 3929
rect 1241 3928 1256 3929
rect 1256 3928 1275 3929
rect 1313 3928 1324 3929
rect 1324 3928 1347 3929
rect 1385 3928 1392 3929
rect 1392 3928 1419 3929
rect 1457 3928 1460 3929
rect 1460 3928 1491 3929
rect 1529 3928 1563 3954
rect 1601 3946 1635 3962
rect 1601 3928 1609 3946
rect 1609 3928 1635 3946
rect 1169 3860 1203 3889
rect 1241 3860 1275 3889
rect 1313 3860 1347 3889
rect 1385 3860 1419 3889
rect 1457 3860 1491 3889
rect 1529 3885 1541 3889
rect 1541 3885 1563 3889
rect 1169 3855 1188 3860
rect 1188 3855 1203 3860
rect 1241 3855 1256 3860
rect 1256 3855 1275 3860
rect 1313 3855 1324 3860
rect 1324 3855 1347 3860
rect 1385 3855 1392 3860
rect 1392 3855 1419 3860
rect 1457 3855 1460 3860
rect 1460 3855 1491 3860
rect 1529 3855 1563 3885
rect 1601 3876 1635 3889
rect 1601 3855 1609 3876
rect 1609 3855 1635 3876
rect 1169 3791 1203 3816
rect 1241 3791 1275 3816
rect 1313 3791 1347 3816
rect 1385 3791 1419 3816
rect 1457 3791 1491 3816
rect 1169 3782 1188 3791
rect 1188 3782 1203 3791
rect 1241 3782 1256 3791
rect 1256 3782 1275 3791
rect 1313 3782 1324 3791
rect 1324 3782 1347 3791
rect 1385 3782 1392 3791
rect 1392 3782 1419 3791
rect 1457 3782 1460 3791
rect 1460 3782 1491 3791
rect 1529 3782 1563 3816
rect 1601 3806 1635 3816
rect 1601 3782 1609 3806
rect 1609 3782 1635 3806
rect 1169 3722 1203 3743
rect 1241 3722 1275 3743
rect 1313 3722 1347 3743
rect 1385 3722 1419 3743
rect 1457 3722 1491 3743
rect 1169 3709 1188 3722
rect 1188 3709 1203 3722
rect 1241 3709 1256 3722
rect 1256 3709 1275 3722
rect 1313 3709 1324 3722
rect 1324 3709 1347 3722
rect 1385 3709 1392 3722
rect 1392 3709 1419 3722
rect 1457 3709 1460 3722
rect 1460 3709 1491 3722
rect 1529 3712 1563 3743
rect 1601 3736 1635 3743
rect 1529 3709 1541 3712
rect 1541 3709 1563 3712
rect 1601 3709 1609 3736
rect 1609 3709 1635 3736
rect 1169 3653 1203 3670
rect 1241 3653 1275 3670
rect 1313 3653 1347 3670
rect 1385 3653 1419 3670
rect 1457 3653 1491 3670
rect 1169 3636 1203 3653
rect 1241 3636 1275 3653
rect 1313 3636 1347 3653
rect 1385 3636 1419 3653
rect 1457 3636 1460 3653
rect 1460 3636 1491 3653
rect 1529 3643 1563 3670
rect 1601 3666 1635 3670
rect 1529 3636 1541 3643
rect 1541 3636 1563 3643
rect 1601 3636 1609 3666
rect 1609 3636 1635 3666
rect 1169 3563 1203 3597
rect 1241 3563 1275 3597
rect 1313 3563 1347 3597
rect 1385 3563 1419 3597
rect 1457 3563 1460 3597
rect 1460 3563 1491 3597
rect 1529 3574 1563 3597
rect 1601 3596 1635 3597
rect 1529 3563 1541 3574
rect 1541 3563 1563 3574
rect 1601 3563 1609 3596
rect 1609 3563 1635 3596
rect 1169 3490 1203 3524
rect 1241 3490 1275 3524
rect 1313 3490 1347 3524
rect 1385 3490 1419 3524
rect 1457 3490 1460 3524
rect 1460 3490 1491 3524
rect 1529 3505 1563 3524
rect 1529 3490 1541 3505
rect 1541 3490 1563 3505
rect 1601 3492 1609 3524
rect 1609 3492 1635 3524
rect 1601 3490 1635 3492
rect 1169 3417 1203 3451
rect 1241 3417 1275 3451
rect 1313 3417 1347 3451
rect 1385 3417 1419 3451
rect 1457 3417 1460 3451
rect 1460 3417 1491 3451
rect 1529 3436 1563 3451
rect 1529 3417 1541 3436
rect 1541 3417 1563 3436
rect 1601 3422 1609 3451
rect 1609 3422 1635 3451
rect 1601 3417 1635 3422
rect 1169 3344 1203 3378
rect 1241 3344 1275 3378
rect 1313 3344 1347 3378
rect 1385 3344 1419 3378
rect 1457 3344 1460 3378
rect 1460 3344 1491 3378
rect 1529 3367 1563 3378
rect 1529 3344 1541 3367
rect 1541 3344 1563 3367
rect 1601 3352 1609 3378
rect 1609 3352 1635 3378
rect 1601 3344 1635 3352
rect 1169 3271 1203 3305
rect 1241 3271 1275 3305
rect 1313 3271 1347 3305
rect 1385 3271 1419 3305
rect 1457 3271 1460 3305
rect 1460 3271 1491 3305
rect 1529 3298 1563 3305
rect 1529 3271 1541 3298
rect 1541 3271 1563 3298
rect 1601 3282 1609 3305
rect 1609 3282 1635 3305
rect 1601 3271 1635 3282
rect 1169 3198 1203 3232
rect 1241 3198 1275 3232
rect 1313 3198 1347 3232
rect 1385 3198 1419 3232
rect 1457 3198 1460 3232
rect 1460 3198 1491 3232
rect 1529 3229 1563 3232
rect 1529 3198 1541 3229
rect 1541 3198 1563 3229
rect 1601 3212 1609 3232
rect 1609 3212 1635 3232
rect 1712 3224 1740 3228
rect 1740 3224 1746 3228
rect 1785 3224 1809 3228
rect 1809 3224 1819 3228
rect 1858 3224 1878 3228
rect 1878 3224 1892 3228
rect 1931 3224 1947 3228
rect 1947 3224 1965 3228
rect 2004 3224 2016 3228
rect 2016 3224 2038 3228
rect 2077 3224 2085 3228
rect 2085 3224 2111 3228
rect 2150 3224 2154 3228
rect 2154 3224 2184 3228
rect 2223 3224 2257 3228
rect 2296 3224 2326 3228
rect 2326 3224 2330 3228
rect 2369 3224 2395 3228
rect 2395 3224 2403 3228
rect 2442 3224 2464 3228
rect 2464 3224 2476 3228
rect 2515 3224 2533 3228
rect 2533 3224 2549 3228
rect 2588 3224 2602 3228
rect 2602 3224 2622 3228
rect 2661 3224 2671 3228
rect 2671 3224 2695 3228
rect 2734 3224 2740 3228
rect 2740 3224 2768 3228
rect 2807 3224 2809 3228
rect 2809 3224 2844 3228
rect 1601 3198 1635 3212
rect 1712 3194 1746 3224
rect 1785 3194 1819 3224
rect 1858 3194 1892 3224
rect 1931 3194 1965 3224
rect 2004 3194 2038 3224
rect 2077 3194 2111 3224
rect 2150 3194 2184 3224
rect 2223 3194 2257 3224
rect 2296 3194 2330 3224
rect 2369 3194 2403 3224
rect 2442 3194 2476 3224
rect 2515 3194 2549 3224
rect 2588 3194 2622 3224
rect 2661 3194 2695 3224
rect 2734 3194 2768 3224
rect 2807 3190 2844 3224
rect 1169 3125 1203 3159
rect 1241 3125 1275 3159
rect 1313 3125 1347 3159
rect 1385 3125 1419 3159
rect 1457 3125 1460 3159
rect 1460 3125 1491 3159
rect 1529 3126 1541 3159
rect 1541 3126 1563 3159
rect 1601 3142 1609 3159
rect 1609 3142 1635 3159
rect 2807 3156 2809 3190
rect 2809 3156 2844 3190
rect 1529 3125 1563 3126
rect 1601 3125 1635 3142
rect 1712 3122 1746 3156
rect 1785 3122 1819 3156
rect 1858 3122 1892 3156
rect 1931 3122 1965 3156
rect 2004 3122 2038 3156
rect 2077 3122 2111 3156
rect 2150 3122 2184 3156
rect 2223 3122 2257 3156
rect 2296 3122 2330 3156
rect 2369 3122 2403 3156
rect 2442 3122 2476 3156
rect 2515 3122 2549 3156
rect 2588 3122 2622 3156
rect 2661 3122 2695 3156
rect 2734 3122 2768 3156
rect 2807 3122 2844 3156
rect 2844 3122 2985 3228
rect 1169 3052 1203 3086
rect 1241 3052 1275 3086
rect 1313 3052 1347 3086
rect 1385 3052 1419 3086
rect 1457 3052 1460 3086
rect 1460 3052 1491 3086
rect 1529 3057 1541 3086
rect 1541 3057 1563 3086
rect 1601 3073 1609 3086
rect 1609 3073 1635 3086
rect 1529 3052 1563 3057
rect 1601 3052 1635 3073
rect 1169 2979 1203 3013
rect 1241 2979 1275 3013
rect 1313 2979 1347 3013
rect 1385 2979 1419 3013
rect 1457 2979 1460 3013
rect 1460 2979 1491 3013
rect 1529 2988 1541 3013
rect 1541 2988 1563 3013
rect 1601 3004 1609 3013
rect 1609 3004 1635 3013
rect 1529 2979 1563 2988
rect 1601 2979 1635 3004
rect 1169 2906 1203 2940
rect 1241 2906 1275 2940
rect 1313 2906 1347 2940
rect 1385 2906 1419 2940
rect 1457 2906 1460 2940
rect 1460 2906 1491 2940
rect 1529 2919 1541 2940
rect 1541 2919 1563 2940
rect 1601 2935 1609 2940
rect 1609 2935 1635 2940
rect 1529 2906 1563 2919
rect 1601 2906 1635 2935
rect 1169 2833 1203 2867
rect 1241 2833 1275 2867
rect 1313 2833 1347 2867
rect 1385 2833 1419 2867
rect 1457 2833 1460 2867
rect 1460 2833 1491 2867
rect 1529 2850 1541 2867
rect 1541 2850 1563 2867
rect 1601 2866 1609 2867
rect 1609 2866 1635 2867
rect 1529 2833 1563 2850
rect 1601 2833 1635 2866
rect 1169 2760 1203 2794
rect 1241 2760 1275 2794
rect 1313 2760 1347 2794
rect 1385 2760 1419 2794
rect 1457 2760 1460 2794
rect 1460 2760 1491 2794
rect 1529 2781 1541 2794
rect 1541 2781 1563 2794
rect 1529 2760 1563 2781
rect 1601 2762 1635 2794
rect 1601 2760 1609 2762
rect 1609 2760 1635 2762
rect 1169 2687 1203 2721
rect 1241 2687 1275 2721
rect 1313 2687 1347 2721
rect 1385 2687 1419 2721
rect 1457 2687 1460 2721
rect 1460 2687 1491 2721
rect 1529 2712 1541 2721
rect 1541 2712 1563 2721
rect 1529 2687 1563 2712
rect 1601 2693 1635 2721
rect 1601 2687 1609 2693
rect 1609 2687 1635 2693
rect 1169 2614 1203 2648
rect 1241 2614 1275 2648
rect 1313 2614 1347 2648
rect 1385 2614 1419 2648
rect 1457 2614 1460 2648
rect 1460 2614 1491 2648
rect 1529 2643 1541 2648
rect 1541 2643 1563 2648
rect 1529 2614 1563 2643
rect 1601 2624 1635 2648
rect 1601 2614 1609 2624
rect 1609 2614 1635 2624
rect 1169 2541 1203 2575
rect 1241 2541 1275 2575
rect 1313 2541 1347 2575
rect 1385 2541 1419 2575
rect 1457 2541 1460 2575
rect 1460 2541 1491 2575
rect 1529 2541 1563 2575
rect 1601 2555 1635 2575
rect 1601 2541 1609 2555
rect 1609 2541 1635 2555
rect 1169 2468 1203 2502
rect 1241 2468 1275 2502
rect 1313 2468 1347 2502
rect 1385 2468 1419 2502
rect 1457 2468 1460 2502
rect 1460 2468 1491 2502
rect 1529 2473 1563 2502
rect 1601 2486 1635 2502
rect 1529 2468 1541 2473
rect 1541 2468 1563 2473
rect 1601 2468 1609 2486
rect 1609 2468 1635 2486
rect 1169 2395 1203 2429
rect 1241 2395 1275 2429
rect 1313 2395 1347 2429
rect 1385 2395 1419 2429
rect 1457 2395 1460 2429
rect 1460 2395 1491 2429
rect 1529 2405 1563 2429
rect 1601 2417 1635 2429
rect 1529 2395 1541 2405
rect 1541 2395 1563 2405
rect 1601 2395 1609 2417
rect 1609 2395 1635 2417
rect 7104 2375 7138 2409
rect 7179 2375 7213 2409
rect 7254 2375 7288 2409
rect 7329 2375 7363 2409
rect 7403 2375 7437 2409
rect 7477 2375 7511 2409
rect 7551 2375 7585 2409
rect 7625 2375 7659 2409
rect 7699 2375 7733 2409
rect 7773 2375 7807 2409
rect 7847 2375 7881 2409
rect 7921 2375 7955 2409
rect 7995 2375 8029 2409
rect 8069 2375 8103 2409
rect 8143 2375 8177 2409
rect 8217 2375 8251 2409
rect 8291 2375 8325 2409
rect 8365 2375 8399 2409
rect 8439 2375 8473 2409
rect 8513 2375 8547 2409
rect 1169 2322 1203 2356
rect 1241 2322 1275 2356
rect 1313 2322 1347 2356
rect 1385 2322 1419 2356
rect 1457 2322 1460 2356
rect 1460 2322 1491 2356
rect 1529 2337 1563 2356
rect 1601 2348 1635 2356
rect 1529 2322 1541 2337
rect 1541 2322 1563 2337
rect 1601 2322 1609 2348
rect 1609 2322 1635 2348
rect 1712 2327 1740 2330
rect 1740 2327 1746 2330
rect 1786 2327 1809 2330
rect 1809 2327 1820 2330
rect 1860 2327 1878 2330
rect 1878 2327 1894 2330
rect 1934 2327 1947 2330
rect 1947 2327 1968 2330
rect 2008 2327 2016 2330
rect 2016 2327 2042 2330
rect 2082 2327 2085 2330
rect 2085 2327 2116 2330
rect 2156 2327 2188 2330
rect 2188 2327 2190 2330
rect 2230 2327 2257 2330
rect 2257 2327 2264 2330
rect 2304 2327 2326 2330
rect 2326 2327 2338 2330
rect 2378 2327 2395 2330
rect 2395 2327 2412 2330
rect 2452 2327 2464 2330
rect 2464 2327 2486 2330
rect 2526 2327 2533 2330
rect 2533 2327 2560 2330
rect 2599 2327 2602 2330
rect 2602 2327 2633 2330
rect 1712 2296 1746 2327
rect 1786 2296 1820 2327
rect 1860 2296 1894 2327
rect 1934 2296 1968 2327
rect 2008 2296 2042 2327
rect 2082 2296 2116 2327
rect 2156 2296 2190 2327
rect 2230 2296 2264 2327
rect 2304 2296 2338 2327
rect 2378 2296 2412 2327
rect 2452 2296 2486 2327
rect 2526 2296 2560 2327
rect 2599 2296 2633 2327
rect 2672 2296 2706 2330
rect 2745 2327 2775 2330
rect 2775 2327 2779 2330
rect 2745 2296 2779 2327
rect 2818 2296 2844 2330
rect 2844 2296 2852 2330
rect 2891 2296 2925 2330
rect 2964 2296 2998 2330
rect 1169 2249 1203 2283
rect 1241 2249 1275 2283
rect 1313 2249 1347 2283
rect 1385 2249 1419 2283
rect 1457 2249 1460 2283
rect 1460 2249 1491 2283
rect 1529 2269 1563 2283
rect 1601 2279 1635 2283
rect 1529 2249 1541 2269
rect 1541 2249 1563 2269
rect 1601 2249 1609 2279
rect 1609 2249 1635 2279
rect 1712 2225 1746 2258
rect 1786 2225 1820 2258
rect 1860 2225 1894 2258
rect 1934 2225 1968 2258
rect 2008 2225 2042 2258
rect 2082 2225 2116 2258
rect 2156 2225 2190 2258
rect 2230 2225 2264 2258
rect 2304 2225 2338 2258
rect 2378 2225 2412 2258
rect 2452 2225 2486 2258
rect 2526 2225 2560 2258
rect 2599 2225 2633 2258
rect 1712 2224 1740 2225
rect 1740 2224 1746 2225
rect 1786 2224 1809 2225
rect 1809 2224 1820 2225
rect 1860 2224 1878 2225
rect 1878 2224 1894 2225
rect 1934 2224 1947 2225
rect 1947 2224 1968 2225
rect 2008 2224 2016 2225
rect 2016 2224 2042 2225
rect 2082 2224 2085 2225
rect 2085 2224 2116 2225
rect 1169 2176 1203 2210
rect 1241 2176 1275 2210
rect 1313 2176 1347 2210
rect 1385 2176 1419 2210
rect 1457 2176 1460 2210
rect 1460 2176 1491 2210
rect 1529 2201 1563 2210
rect 1529 2176 1541 2201
rect 1541 2176 1563 2201
rect 1601 2176 1609 2210
rect 1609 2176 1635 2210
rect 2156 2224 2188 2225
rect 2188 2224 2190 2225
rect 2230 2224 2257 2225
rect 2257 2224 2264 2225
rect 2304 2224 2326 2225
rect 2326 2224 2338 2225
rect 2378 2224 2395 2225
rect 2395 2224 2412 2225
rect 2452 2224 2464 2225
rect 2464 2224 2486 2225
rect 2526 2224 2533 2225
rect 2533 2224 2560 2225
rect 2599 2224 2602 2225
rect 2602 2224 2633 2225
rect 2672 2224 2706 2258
rect 2745 2225 2779 2258
rect 2745 2224 2775 2225
rect 2775 2224 2779 2225
rect 2818 2224 2844 2258
rect 2844 2224 2852 2258
rect 2891 2224 2925 2258
rect 2964 2224 2998 2258
rect 7104 2303 7138 2337
rect 7179 2303 7213 2337
rect 7254 2303 7288 2337
rect 7329 2303 7363 2337
rect 7403 2303 7437 2337
rect 7477 2303 7511 2337
rect 7551 2303 7585 2337
rect 7625 2303 7659 2337
rect 7699 2303 7733 2337
rect 7773 2303 7807 2337
rect 7847 2303 7881 2337
rect 7921 2303 7955 2337
rect 7995 2303 8029 2337
rect 8069 2303 8103 2337
rect 8143 2303 8177 2337
rect 8217 2303 8251 2337
rect 8291 2303 8325 2337
rect 8365 2303 8399 2337
rect 8439 2303 8473 2337
rect 8513 2303 8547 2337
rect 7104 2231 7138 2265
rect 7179 2231 7213 2265
rect 7254 2231 7288 2265
rect 7329 2231 7363 2265
rect 7403 2231 7437 2265
rect 7477 2231 7511 2265
rect 7551 2231 7585 2265
rect 7625 2231 7659 2265
rect 7699 2231 7733 2265
rect 7773 2231 7807 2265
rect 7847 2231 7881 2265
rect 7921 2231 7955 2265
rect 7995 2231 8029 2265
rect 8069 2231 8103 2265
rect 8143 2231 8177 2265
rect 8217 2231 8251 2265
rect 8291 2231 8325 2265
rect 8365 2231 8399 2265
rect 8439 2231 8473 2265
rect 8513 2231 8547 2265
rect 1169 2103 1203 2137
rect 1241 2103 1275 2137
rect 1313 2103 1347 2137
rect 1385 2103 1419 2137
rect 1457 2103 1460 2137
rect 1460 2103 1491 2137
rect 1529 2133 1563 2137
rect 1529 2103 1541 2133
rect 1541 2103 1563 2133
rect 1601 2107 1609 2137
rect 1609 2107 1635 2137
rect 1601 2103 1635 2107
rect 1169 2030 1203 2064
rect 1241 2030 1275 2064
rect 1313 2030 1347 2064
rect 1385 2030 1419 2064
rect 1457 2030 1460 2064
rect 1460 2030 1491 2064
rect 1529 2031 1541 2064
rect 1541 2031 1563 2064
rect 1601 2038 1609 2064
rect 1609 2038 1635 2064
rect 1529 2030 1563 2031
rect 1601 2030 1635 2038
rect 1169 1957 1203 1991
rect 1241 1957 1275 1991
rect 1313 1957 1347 1991
rect 1385 1957 1419 1991
rect 1457 1957 1460 1991
rect 1460 1957 1491 1991
rect 1529 1963 1541 1991
rect 1541 1963 1563 1991
rect 1601 1969 1609 1991
rect 1609 1969 1635 1991
rect 1529 1957 1563 1963
rect 1601 1957 1635 1969
rect 1169 1884 1203 1918
rect 1241 1884 1275 1918
rect 1313 1884 1347 1918
rect 1385 1884 1419 1918
rect 1457 1884 1460 1918
rect 1460 1884 1491 1918
rect 1529 1895 1541 1918
rect 1541 1895 1563 1918
rect 1601 1900 1609 1918
rect 1609 1900 1635 1918
rect 1529 1884 1563 1895
rect 1601 1884 1635 1900
rect 1169 1811 1203 1845
rect 1241 1811 1275 1845
rect 1313 1811 1347 1845
rect 1385 1811 1419 1845
rect 1457 1811 1460 1845
rect 1460 1811 1491 1845
rect 1529 1827 1541 1845
rect 1541 1827 1563 1845
rect 1601 1831 1609 1845
rect 1609 1831 1635 1845
rect 1529 1811 1563 1827
rect 1601 1811 1635 1831
rect 8824 3636 8847 3663
rect 8847 3636 8858 3663
rect 8898 3636 8915 3663
rect 8915 3636 8932 3663
rect 8972 3636 8983 3663
rect 8983 3636 9006 3663
rect 9046 3636 9051 3663
rect 9051 3636 9080 3663
rect 9120 3636 9153 3663
rect 9153 3636 9154 3663
rect 9194 3636 9221 3663
rect 9221 3636 9228 3663
rect 9268 3636 9289 3663
rect 9289 3636 9302 3663
rect 9342 3636 9357 3663
rect 9357 3636 9376 3663
rect 9416 3636 9425 3663
rect 9425 3636 9450 3663
rect 9490 3636 9493 3663
rect 9493 3636 9524 3663
rect 9564 3636 9595 3663
rect 9595 3636 9598 3663
rect 9638 3636 9663 3663
rect 9663 3636 9672 3663
rect 9712 3636 9731 3663
rect 9731 3636 9746 3663
rect 9786 3636 9799 3663
rect 9799 3636 9820 3663
rect 9860 3636 9867 3663
rect 9867 3636 9894 3663
rect 9934 3636 9935 3663
rect 9935 3636 9968 3663
rect 10008 3636 10037 3663
rect 10037 3636 10042 3663
rect 10082 3636 10105 3663
rect 10105 3636 10116 3663
rect 10156 3636 10173 3663
rect 10173 3636 10190 3663
rect 10230 3636 10241 3663
rect 10241 3636 10264 3663
rect 8824 3629 8858 3636
rect 8898 3629 8932 3636
rect 8972 3629 9006 3636
rect 9046 3629 9080 3636
rect 9120 3629 9154 3636
rect 9194 3629 9228 3636
rect 9268 3629 9302 3636
rect 9342 3629 9376 3636
rect 9416 3629 9450 3636
rect 9490 3629 9524 3636
rect 9564 3629 9598 3636
rect 9638 3629 9672 3636
rect 9712 3629 9746 3636
rect 9786 3629 9820 3636
rect 9860 3629 9894 3636
rect 9934 3629 9968 3636
rect 10008 3629 10042 3636
rect 10082 3629 10116 3636
rect 10156 3629 10190 3636
rect 10230 3629 10264 3636
rect 10304 3637 10312 3663
rect 10312 3637 10338 3663
rect 10378 3637 10380 3663
rect 10380 3637 10412 3663
rect 10452 3637 10482 3663
rect 10482 3637 10486 3663
rect 10526 3637 10550 3663
rect 10550 3637 10560 3663
rect 10600 3637 10618 3663
rect 10618 3637 10634 3663
rect 10674 3637 10686 3663
rect 10686 3637 10708 3663
rect 10748 3637 10754 3663
rect 10754 3637 10782 3663
rect 10304 3629 10338 3637
rect 10378 3629 10412 3637
rect 10452 3629 10486 3637
rect 10526 3629 10560 3637
rect 10600 3629 10634 3637
rect 10674 3629 10708 3637
rect 10748 3629 10782 3637
rect 10822 3629 10856 3663
rect 10896 3637 10924 3663
rect 10924 3637 10930 3663
rect 10970 3637 10992 3663
rect 10992 3637 11004 3663
rect 11043 3637 11060 3663
rect 11060 3637 11077 3663
rect 11116 3637 11128 3663
rect 11128 3637 11150 3663
rect 11189 3637 11196 3663
rect 11196 3637 11223 3663
rect 11262 3637 11264 3663
rect 11264 3637 11296 3663
rect 11335 3637 11366 3663
rect 11366 3637 11369 3663
rect 11408 3637 11434 3663
rect 11434 3637 11442 3663
rect 11481 3637 11502 3663
rect 11502 3637 11515 3663
rect 10896 3629 10930 3637
rect 10970 3629 11004 3637
rect 11043 3629 11077 3637
rect 11116 3629 11150 3637
rect 11189 3629 11223 3637
rect 11262 3629 11296 3637
rect 11335 3629 11369 3637
rect 11408 3629 11442 3637
rect 11481 3629 11515 3637
rect 8824 3566 8847 3591
rect 8847 3566 8858 3591
rect 8898 3566 8915 3591
rect 8915 3566 8932 3591
rect 8972 3566 8983 3591
rect 8983 3566 9006 3591
rect 9046 3566 9051 3591
rect 9051 3566 9080 3591
rect 9120 3566 9153 3591
rect 9153 3566 9154 3591
rect 9194 3566 9221 3591
rect 9221 3566 9228 3591
rect 9268 3566 9289 3591
rect 9289 3566 9302 3591
rect 9342 3566 9357 3591
rect 9357 3566 9376 3591
rect 9416 3566 9425 3591
rect 9425 3566 9450 3591
rect 9490 3566 9493 3591
rect 9493 3566 9524 3591
rect 9564 3566 9595 3591
rect 9595 3566 9598 3591
rect 9638 3566 9663 3591
rect 9663 3566 9672 3591
rect 9712 3566 9731 3591
rect 9731 3566 9746 3591
rect 9786 3566 9799 3591
rect 9799 3566 9820 3591
rect 9860 3566 9867 3591
rect 9867 3566 9894 3591
rect 9934 3566 9935 3591
rect 9935 3566 9968 3591
rect 10008 3566 10037 3591
rect 10037 3566 10042 3591
rect 10082 3566 10105 3591
rect 10105 3566 10116 3591
rect 10156 3566 10173 3591
rect 10173 3566 10190 3591
rect 10230 3566 10241 3591
rect 10241 3566 10264 3591
rect 8824 3557 8858 3566
rect 8898 3557 8932 3566
rect 8972 3557 9006 3566
rect 9046 3557 9080 3566
rect 9120 3557 9154 3566
rect 9194 3557 9228 3566
rect 9268 3557 9302 3566
rect 9342 3557 9376 3566
rect 9416 3557 9450 3566
rect 9490 3557 9524 3566
rect 9564 3557 9598 3566
rect 9638 3557 9672 3566
rect 9712 3557 9746 3566
rect 9786 3557 9820 3566
rect 9860 3557 9894 3566
rect 9934 3557 9968 3566
rect 10008 3557 10042 3566
rect 10082 3557 10116 3566
rect 10156 3557 10190 3566
rect 10230 3557 10264 3566
rect 10304 3567 10312 3591
rect 10312 3567 10338 3591
rect 10378 3567 10380 3591
rect 10380 3567 10412 3591
rect 10452 3567 10482 3591
rect 10482 3567 10486 3591
rect 10526 3567 10550 3591
rect 10550 3567 10560 3591
rect 10600 3567 10618 3591
rect 10618 3567 10634 3591
rect 10674 3567 10686 3591
rect 10686 3567 10708 3591
rect 10748 3567 10754 3591
rect 10754 3567 10782 3591
rect 10304 3557 10338 3567
rect 10378 3557 10412 3567
rect 10452 3557 10486 3567
rect 10526 3557 10560 3567
rect 10600 3557 10634 3567
rect 10674 3557 10708 3567
rect 10748 3557 10782 3567
rect 10822 3557 10856 3591
rect 10896 3567 10924 3591
rect 10924 3567 10930 3591
rect 10970 3567 10992 3591
rect 10992 3567 11004 3591
rect 11043 3567 11060 3591
rect 11060 3567 11077 3591
rect 11116 3567 11128 3591
rect 11128 3567 11150 3591
rect 11189 3567 11196 3591
rect 11196 3567 11223 3591
rect 11262 3567 11264 3591
rect 11264 3567 11296 3591
rect 11335 3567 11366 3591
rect 11366 3567 11369 3591
rect 11408 3567 11434 3591
rect 11434 3567 11442 3591
rect 11481 3567 11502 3591
rect 11502 3567 11515 3591
rect 10896 3557 10930 3567
rect 10970 3557 11004 3567
rect 11043 3557 11077 3567
rect 11116 3557 11150 3567
rect 11189 3557 11223 3567
rect 11262 3557 11296 3567
rect 11335 3557 11369 3567
rect 11408 3557 11442 3567
rect 11481 3557 11515 3567
rect 8824 3496 8847 3519
rect 8847 3496 8858 3519
rect 8898 3496 8915 3519
rect 8915 3496 8932 3519
rect 8972 3496 8983 3519
rect 8983 3496 9006 3519
rect 9046 3496 9051 3519
rect 9051 3496 9080 3519
rect 9120 3496 9153 3519
rect 9153 3496 9154 3519
rect 9194 3496 9221 3519
rect 9221 3496 9228 3519
rect 9268 3496 9289 3519
rect 9289 3496 9302 3519
rect 9342 3496 9357 3519
rect 9357 3496 9376 3519
rect 9416 3496 9425 3519
rect 9425 3496 9450 3519
rect 9490 3496 9493 3519
rect 9493 3496 9524 3519
rect 9564 3496 9595 3519
rect 9595 3496 9598 3519
rect 9638 3496 9663 3519
rect 9663 3496 9672 3519
rect 9712 3496 9731 3519
rect 9731 3496 9746 3519
rect 9786 3496 9799 3519
rect 9799 3496 9820 3519
rect 9860 3496 9867 3519
rect 9867 3496 9894 3519
rect 9934 3496 9935 3519
rect 9935 3496 9968 3519
rect 10008 3496 10037 3519
rect 10037 3496 10042 3519
rect 10082 3496 10105 3519
rect 10105 3496 10116 3519
rect 10156 3496 10173 3519
rect 10173 3496 10190 3519
rect 10230 3496 10241 3519
rect 10241 3496 10264 3519
rect 8824 3485 8858 3496
rect 8898 3485 8932 3496
rect 8972 3485 9006 3496
rect 9046 3485 9080 3496
rect 9120 3485 9154 3496
rect 9194 3485 9228 3496
rect 9268 3485 9302 3496
rect 9342 3485 9376 3496
rect 9416 3485 9450 3496
rect 9490 3485 9524 3496
rect 9564 3485 9598 3496
rect 9638 3485 9672 3496
rect 9712 3485 9746 3496
rect 9786 3485 9820 3496
rect 9860 3485 9894 3496
rect 9934 3485 9968 3496
rect 10008 3485 10042 3496
rect 10082 3485 10116 3496
rect 10156 3485 10190 3496
rect 10230 3485 10264 3496
rect 10304 3497 10312 3519
rect 10312 3497 10338 3519
rect 10378 3497 10380 3519
rect 10380 3497 10412 3519
rect 10452 3497 10482 3519
rect 10482 3497 10486 3519
rect 10526 3497 10550 3519
rect 10550 3497 10560 3519
rect 10600 3497 10618 3519
rect 10618 3497 10634 3519
rect 10674 3497 10686 3519
rect 10686 3497 10708 3519
rect 10748 3497 10754 3519
rect 10754 3497 10782 3519
rect 10304 3485 10338 3497
rect 10378 3485 10412 3497
rect 10452 3485 10486 3497
rect 10526 3485 10560 3497
rect 10600 3485 10634 3497
rect 10674 3485 10708 3497
rect 10748 3485 10782 3497
rect 10822 3485 10856 3519
rect 10896 3497 10924 3519
rect 10924 3497 10930 3519
rect 10970 3497 10992 3519
rect 10992 3497 11004 3519
rect 11043 3497 11060 3519
rect 11060 3497 11077 3519
rect 11116 3497 11128 3519
rect 11128 3497 11150 3519
rect 11189 3497 11196 3519
rect 11196 3497 11223 3519
rect 11262 3497 11264 3519
rect 11264 3497 11296 3519
rect 11335 3497 11366 3519
rect 11366 3497 11369 3519
rect 11408 3497 11434 3519
rect 11434 3497 11442 3519
rect 11481 3497 11502 3519
rect 11502 3497 11515 3519
rect 10896 3485 10930 3497
rect 10970 3485 11004 3497
rect 11043 3485 11077 3497
rect 11116 3485 11150 3497
rect 11189 3485 11223 3497
rect 11262 3485 11296 3497
rect 11335 3485 11369 3497
rect 11408 3485 11442 3497
rect 11481 3485 11515 3497
rect 23593 4392 23627 4398
rect 23665 4392 23699 4398
rect 23737 4392 23771 4398
rect 23593 4364 23597 4392
rect 23597 4364 23627 4392
rect 23665 4364 23699 4392
rect 23737 4364 23767 4392
rect 23767 4364 23771 4392
rect 23593 4323 23627 4325
rect 23665 4323 23699 4325
rect 23737 4323 23771 4325
rect 23593 4291 23597 4323
rect 23597 4291 23627 4323
rect 23665 4291 23699 4323
rect 23737 4291 23767 4323
rect 23767 4291 23771 4323
rect 16973 4223 16976 4256
rect 16976 4223 17007 4256
rect 17045 4223 17078 4256
rect 17078 4223 17079 4256
rect 16973 4222 17007 4223
rect 17045 4222 17079 4223
rect 19124 4223 19152 4257
rect 19152 4223 19158 4257
rect 19196 4223 19220 4257
rect 19220 4223 19230 4257
rect 23593 4220 23597 4252
rect 23597 4220 23627 4252
rect 23665 4220 23699 4252
rect 23737 4220 23767 4252
rect 23767 4220 23771 4252
rect 23593 4218 23627 4220
rect 23665 4218 23699 4220
rect 23737 4218 23771 4220
rect 23593 4151 23597 4179
rect 23597 4151 23627 4179
rect 23665 4151 23699 4179
rect 23737 4151 23767 4179
rect 23767 4151 23771 4179
rect 23593 4145 23627 4151
rect 23665 4145 23699 4151
rect 23737 4145 23771 4151
rect 23593 4072 23597 4106
rect 23597 4072 23627 4106
rect 23665 4072 23699 4106
rect 23737 4072 23767 4106
rect 23767 4072 23771 4106
rect 12594 4049 12595 4059
rect 12595 4049 12629 4059
rect 12629 4049 12663 4059
rect 12663 4049 12697 4059
rect 12697 4049 12731 4059
rect 12731 4049 12765 4059
rect 12765 4049 12799 4059
rect 12799 4049 12833 4059
rect 12833 4049 12867 4059
rect 12867 4049 12901 4059
rect 12901 4049 12935 4059
rect 12935 4049 12969 4059
rect 12969 4049 13003 4059
rect 13003 4049 13037 4059
rect 13037 4049 13071 4059
rect 13071 4049 13105 4059
rect 13105 4049 13139 4059
rect 13139 4049 13173 4059
rect 13173 4049 13207 4059
rect 13207 4049 13241 4059
rect 13241 4049 13275 4059
rect 13275 4049 13309 4059
rect 13309 4049 13343 4059
rect 13343 4049 13377 4059
rect 13377 4049 15580 4059
rect 12594 4013 15580 4049
rect 12594 3979 12595 4013
rect 12595 3979 12629 4013
rect 12629 3979 12663 4013
rect 12663 3979 12697 4013
rect 12697 3979 12731 4013
rect 12731 3979 12765 4013
rect 12765 3979 12799 4013
rect 12799 3979 12833 4013
rect 12833 3979 12867 4013
rect 12867 3979 12901 4013
rect 12901 3979 12935 4013
rect 12935 3979 12969 4013
rect 12969 3979 13003 4013
rect 13003 3979 13037 4013
rect 13037 3979 13071 4013
rect 13071 3979 13105 4013
rect 13105 3979 13139 4013
rect 13139 3979 13173 4013
rect 13173 3979 13207 4013
rect 13207 3979 13241 4013
rect 13241 3979 13275 4013
rect 13275 3979 13309 4013
rect 13309 3979 13343 4013
rect 13343 3979 13377 4013
rect 13377 3979 15580 4013
rect 12594 3943 15580 3979
rect 12594 3909 12595 3943
rect 12595 3909 12629 3943
rect 12629 3909 12663 3943
rect 12663 3909 12697 3943
rect 12697 3909 12731 3943
rect 12731 3909 12765 3943
rect 12765 3909 12799 3943
rect 12799 3909 12833 3943
rect 12833 3909 12867 3943
rect 12867 3909 12901 3943
rect 12901 3909 12935 3943
rect 12935 3909 12969 3943
rect 12969 3909 13003 3943
rect 13003 3909 13037 3943
rect 13037 3909 13071 3943
rect 13071 3909 13105 3943
rect 13105 3909 13139 3943
rect 13139 3909 13173 3943
rect 13173 3909 13207 3943
rect 13207 3909 13241 3943
rect 13241 3909 13275 3943
rect 13275 3909 13309 3943
rect 13309 3909 13343 3943
rect 13343 3909 13377 3943
rect 13377 3909 15580 3943
rect 12594 3881 15580 3909
rect 23593 3999 23597 4033
rect 23597 3999 23627 4033
rect 23665 3999 23699 4033
rect 23737 3999 23767 4033
rect 23767 3999 23771 4033
rect 23593 3926 23597 3960
rect 23597 3926 23627 3960
rect 23665 3926 23699 3960
rect 23737 3926 23767 3960
rect 23767 3926 23771 3960
rect 23593 3853 23597 3887
rect 23597 3853 23627 3887
rect 23665 3853 23699 3887
rect 23737 3853 23767 3887
rect 23767 3853 23771 3887
rect 23593 3780 23597 3814
rect 23597 3780 23627 3814
rect 23665 3780 23699 3814
rect 23737 3780 23767 3814
rect 23767 3780 23771 3814
rect 12594 3733 12628 3765
rect 12667 3733 12701 3765
rect 12740 3733 12774 3765
rect 12813 3733 12847 3765
rect 12886 3733 12920 3765
rect 12959 3733 12993 3765
rect 13032 3733 13066 3765
rect 12594 3731 12595 3733
rect 12595 3731 12628 3733
rect 12667 3731 12697 3733
rect 12697 3731 12701 3733
rect 12740 3731 12765 3733
rect 12765 3731 12774 3733
rect 12813 3731 12833 3733
rect 12833 3731 12847 3733
rect 12886 3731 12901 3733
rect 12901 3731 12920 3733
rect 12959 3731 12969 3733
rect 12969 3731 12993 3733
rect 13032 3731 13037 3733
rect 13037 3731 13066 3733
rect 13105 3731 13139 3765
rect 13178 3733 13212 3765
rect 13251 3733 13285 3765
rect 13324 3733 13358 3765
rect 13178 3731 13207 3733
rect 13207 3731 13212 3733
rect 13251 3731 13275 3733
rect 13275 3731 13285 3733
rect 13324 3731 13343 3733
rect 13343 3731 13358 3733
rect 13397 3731 13431 3765
rect 13470 3731 13504 3765
rect 13543 3731 13577 3765
rect 13616 3731 13650 3765
rect 13689 3731 13723 3765
rect 13762 3731 13796 3765
rect 13835 3731 13869 3765
rect 13908 3731 13942 3765
rect 13981 3731 14015 3765
rect 14054 3731 14088 3765
rect 14127 3731 14161 3765
rect 14200 3731 14234 3765
rect 14273 3731 14307 3765
rect 14346 3731 14380 3765
rect 14419 3731 14453 3765
rect 14492 3731 14526 3765
rect 14565 3731 14599 3765
rect 14638 3731 14672 3765
rect 14711 3731 14745 3765
rect 14784 3731 14818 3765
rect 14857 3731 14891 3765
rect 14930 3731 14964 3765
rect 15003 3731 15037 3765
rect 15076 3731 15110 3765
rect 15149 3731 15183 3765
rect 15222 3731 15256 3765
rect 15295 3731 15329 3765
rect 15368 3731 15402 3765
rect 15441 3731 15475 3765
rect 15514 3731 15548 3765
rect 15587 3731 15621 3765
rect 15660 3731 15694 3765
rect 15733 3731 15767 3765
rect 15806 3731 15840 3765
rect 15879 3731 15913 3765
rect 15952 3731 15986 3765
rect 16025 3731 16059 3765
rect 16098 3731 16132 3765
rect 16171 3731 16205 3765
rect 16244 3731 16278 3765
rect 16317 3731 16351 3765
rect 16390 3731 16424 3765
rect 12594 3663 12628 3693
rect 12667 3663 12701 3693
rect 12740 3663 12774 3693
rect 12813 3663 12847 3693
rect 12886 3663 12920 3693
rect 12959 3663 12993 3693
rect 13032 3663 13066 3693
rect 12594 3659 12595 3663
rect 12595 3659 12628 3663
rect 12667 3659 12697 3663
rect 12697 3659 12701 3663
rect 12740 3659 12765 3663
rect 12765 3659 12774 3663
rect 12813 3659 12833 3663
rect 12833 3659 12847 3663
rect 12886 3659 12901 3663
rect 12901 3659 12920 3663
rect 12959 3659 12969 3663
rect 12969 3659 12993 3663
rect 13032 3659 13037 3663
rect 13037 3659 13066 3663
rect 13105 3659 13139 3693
rect 13178 3663 13212 3693
rect 13251 3663 13285 3693
rect 13324 3663 13358 3693
rect 13178 3659 13207 3663
rect 13207 3659 13212 3663
rect 13251 3659 13275 3663
rect 13275 3659 13285 3663
rect 13324 3659 13343 3663
rect 13343 3659 13358 3663
rect 13397 3659 13431 3693
rect 13470 3659 13504 3693
rect 13543 3659 13577 3693
rect 13616 3659 13650 3693
rect 13689 3659 13723 3693
rect 13762 3659 13796 3693
rect 13835 3659 13869 3693
rect 13908 3659 13942 3693
rect 13981 3659 14015 3693
rect 14054 3659 14088 3693
rect 14127 3659 14161 3693
rect 14200 3659 14234 3693
rect 14273 3659 14307 3693
rect 14346 3659 14380 3693
rect 14419 3659 14453 3693
rect 14492 3659 14526 3693
rect 14565 3659 14599 3693
rect 14638 3659 14672 3693
rect 14711 3659 14745 3693
rect 14784 3659 14818 3693
rect 14857 3659 14891 3693
rect 14930 3659 14964 3693
rect 15003 3659 15037 3693
rect 15076 3659 15110 3693
rect 15149 3659 15183 3693
rect 15222 3659 15256 3693
rect 15295 3659 15329 3693
rect 15368 3659 15402 3693
rect 15441 3659 15475 3693
rect 15514 3659 15548 3693
rect 15587 3659 15621 3693
rect 15660 3659 15694 3693
rect 15733 3659 15767 3693
rect 15806 3659 15840 3693
rect 15879 3659 15913 3693
rect 15952 3659 15986 3693
rect 16025 3659 16059 3693
rect 16098 3659 16132 3693
rect 16171 3659 16205 3693
rect 16244 3659 16278 3693
rect 16317 3659 16351 3693
rect 16390 3659 16424 3693
rect 12594 3593 12628 3621
rect 12667 3593 12701 3621
rect 12740 3593 12774 3621
rect 12813 3593 12847 3621
rect 12886 3593 12920 3621
rect 12959 3593 12993 3621
rect 13032 3593 13066 3621
rect 12594 3587 12595 3593
rect 12595 3587 12628 3593
rect 12667 3587 12697 3593
rect 12697 3587 12701 3593
rect 12740 3587 12765 3593
rect 12765 3587 12774 3593
rect 12813 3587 12833 3593
rect 12833 3587 12847 3593
rect 12886 3587 12901 3593
rect 12901 3587 12920 3593
rect 12959 3587 12969 3593
rect 12969 3587 12993 3593
rect 13032 3587 13037 3593
rect 13037 3587 13066 3593
rect 13105 3587 13139 3621
rect 13178 3593 13212 3621
rect 13251 3593 13285 3621
rect 13324 3593 13358 3621
rect 13178 3587 13207 3593
rect 13207 3587 13212 3593
rect 13251 3587 13275 3593
rect 13275 3587 13285 3593
rect 13324 3587 13343 3593
rect 13343 3587 13358 3593
rect 13397 3587 13431 3621
rect 13470 3587 13504 3621
rect 13543 3587 13577 3621
rect 13616 3587 13650 3621
rect 13689 3587 13723 3621
rect 13762 3587 13796 3621
rect 13835 3587 13869 3621
rect 13908 3587 13942 3621
rect 13981 3587 14015 3621
rect 14054 3587 14088 3621
rect 14127 3587 14161 3621
rect 14200 3587 14234 3621
rect 14273 3587 14307 3621
rect 14346 3587 14380 3621
rect 14419 3587 14453 3621
rect 14492 3587 14526 3621
rect 14565 3587 14599 3621
rect 14638 3587 14672 3621
rect 14711 3587 14745 3621
rect 14784 3587 14818 3621
rect 14857 3587 14891 3621
rect 14930 3587 14964 3621
rect 15003 3587 15037 3621
rect 15076 3587 15110 3621
rect 15149 3587 15183 3621
rect 15222 3587 15256 3621
rect 15295 3587 15329 3621
rect 15368 3587 15402 3621
rect 15441 3587 15475 3621
rect 15514 3587 15548 3621
rect 15587 3587 15621 3621
rect 15660 3587 15694 3621
rect 15733 3587 15767 3621
rect 15806 3587 15840 3621
rect 15879 3587 15913 3621
rect 15952 3587 15986 3621
rect 16025 3587 16059 3621
rect 16098 3587 16132 3621
rect 16171 3587 16205 3621
rect 16244 3587 16278 3621
rect 16317 3587 16351 3621
rect 16390 3587 16424 3621
rect 23593 3707 23597 3741
rect 23597 3707 23627 3741
rect 23665 3707 23699 3741
rect 23737 3707 23767 3741
rect 23767 3707 23771 3741
rect 23593 3634 23597 3668
rect 23597 3634 23627 3668
rect 23665 3634 23699 3668
rect 23737 3634 23767 3668
rect 23767 3634 23771 3668
rect 23593 3561 23597 3595
rect 23597 3561 23627 3595
rect 23665 3561 23699 3595
rect 23737 3561 23767 3595
rect 23767 3561 23771 3595
rect 23593 3488 23597 3522
rect 23597 3488 23627 3522
rect 23665 3488 23699 3522
rect 23737 3488 23767 3522
rect 23767 3488 23771 3522
rect 8824 3426 8847 3447
rect 8847 3426 8858 3447
rect 8897 3426 8915 3447
rect 8915 3426 8931 3447
rect 8970 3426 8983 3447
rect 8983 3426 9004 3447
rect 9043 3426 9051 3447
rect 9051 3426 9077 3447
rect 9116 3426 9119 3447
rect 9119 3426 9150 3447
rect 9189 3426 9221 3447
rect 9221 3426 9223 3447
rect 9262 3426 9289 3447
rect 9289 3426 9296 3447
rect 9336 3426 9357 3447
rect 9357 3426 9370 3447
rect 9410 3426 9425 3447
rect 9425 3426 9444 3447
rect 9484 3426 9493 3447
rect 9493 3426 9518 3447
rect 9558 3426 9561 3447
rect 9561 3426 9592 3447
rect 9632 3426 9663 3447
rect 9663 3426 9666 3447
rect 9706 3426 9731 3447
rect 9731 3426 9740 3447
rect 9780 3426 9799 3447
rect 9799 3426 9814 3447
rect 9854 3426 9867 3447
rect 9867 3426 9888 3447
rect 9928 3426 9935 3447
rect 9935 3426 9962 3447
rect 10002 3426 10003 3447
rect 10003 3426 10036 3447
rect 10076 3426 10105 3447
rect 10105 3426 10110 3447
rect 10150 3426 10173 3447
rect 10173 3426 10184 3447
rect 10224 3426 10241 3447
rect 10241 3426 10258 3447
rect 8824 3413 8858 3426
rect 8897 3413 8931 3426
rect 8970 3413 9004 3426
rect 9043 3413 9077 3426
rect 9116 3413 9150 3426
rect 9189 3413 9223 3426
rect 9262 3413 9296 3426
rect 9336 3413 9370 3426
rect 9410 3413 9444 3426
rect 9484 3413 9518 3426
rect 9558 3413 9592 3426
rect 9632 3413 9666 3426
rect 9706 3413 9740 3426
rect 9780 3413 9814 3426
rect 9854 3413 9888 3426
rect 9928 3413 9962 3426
rect 10002 3413 10036 3426
rect 10076 3413 10110 3426
rect 10150 3413 10184 3426
rect 10224 3413 10258 3426
rect 10298 3427 10312 3447
rect 10312 3427 10332 3447
rect 10372 3427 10380 3447
rect 10380 3427 10406 3447
rect 10446 3427 10448 3447
rect 10448 3427 10480 3447
rect 10520 3427 10550 3447
rect 10550 3427 10554 3447
rect 10594 3427 10618 3447
rect 10618 3427 10628 3447
rect 10668 3427 10686 3447
rect 10686 3427 10702 3447
rect 10742 3427 10754 3447
rect 10754 3427 10776 3447
rect 10816 3427 10822 3447
rect 10822 3427 10850 3447
rect 10298 3413 10332 3427
rect 10372 3413 10406 3427
rect 10446 3413 10480 3427
rect 10520 3413 10554 3427
rect 10594 3413 10628 3427
rect 10668 3413 10702 3427
rect 10742 3413 10776 3427
rect 10816 3413 10850 3427
rect 10890 3413 10924 3447
rect 10964 3427 10992 3447
rect 10992 3427 10998 3447
rect 11038 3427 11060 3447
rect 11060 3427 11072 3447
rect 11112 3427 11128 3447
rect 11128 3427 11146 3447
rect 11186 3427 11196 3447
rect 11196 3427 11220 3447
rect 11260 3427 11264 3447
rect 11264 3427 11294 3447
rect 11334 3427 11366 3447
rect 11366 3427 11368 3447
rect 11408 3427 11434 3447
rect 11434 3427 11442 3447
rect 11482 3427 11502 3447
rect 11502 3427 11516 3447
rect 11556 3427 11570 3447
rect 11570 3427 11590 3447
rect 10964 3413 10998 3427
rect 11038 3413 11072 3427
rect 11112 3413 11146 3427
rect 11186 3413 11220 3427
rect 11260 3413 11294 3427
rect 11334 3413 11368 3427
rect 11408 3413 11442 3427
rect 11482 3413 11516 3427
rect 11556 3413 11590 3427
rect 8824 3356 8847 3375
rect 8847 3356 8858 3375
rect 8897 3356 8915 3375
rect 8915 3356 8931 3375
rect 8970 3356 8983 3375
rect 8983 3356 9004 3375
rect 9043 3356 9051 3375
rect 9051 3356 9077 3375
rect 9116 3356 9119 3375
rect 9119 3356 9150 3375
rect 9189 3356 9221 3375
rect 9221 3356 9223 3375
rect 9262 3356 9289 3375
rect 9289 3356 9296 3375
rect 9336 3356 9357 3375
rect 9357 3356 9370 3375
rect 9410 3356 9425 3375
rect 9425 3356 9444 3375
rect 9484 3356 9493 3375
rect 9493 3356 9518 3375
rect 9558 3356 9561 3375
rect 9561 3356 9592 3375
rect 9632 3356 9663 3375
rect 9663 3356 9666 3375
rect 9706 3356 9731 3375
rect 9731 3356 9740 3375
rect 9780 3356 9799 3375
rect 9799 3356 9814 3375
rect 9854 3356 9867 3375
rect 9867 3356 9888 3375
rect 9928 3356 9935 3375
rect 9935 3356 9962 3375
rect 10002 3356 10003 3375
rect 10003 3356 10036 3375
rect 10076 3356 10105 3375
rect 10105 3356 10110 3375
rect 10150 3356 10173 3375
rect 10173 3356 10184 3375
rect 10224 3356 10241 3375
rect 10241 3356 10258 3375
rect 8824 3341 8858 3356
rect 8897 3341 8931 3356
rect 8970 3341 9004 3356
rect 9043 3341 9077 3356
rect 9116 3341 9150 3356
rect 9189 3341 9223 3356
rect 9262 3341 9296 3356
rect 9336 3341 9370 3356
rect 9410 3341 9444 3356
rect 9484 3341 9518 3356
rect 9558 3341 9592 3356
rect 9632 3341 9666 3356
rect 9706 3341 9740 3356
rect 9780 3341 9814 3356
rect 9854 3341 9888 3356
rect 9928 3341 9962 3356
rect 10002 3341 10036 3356
rect 10076 3341 10110 3356
rect 10150 3341 10184 3356
rect 10224 3341 10258 3356
rect 10298 3357 10312 3375
rect 10312 3357 10332 3375
rect 10372 3357 10380 3375
rect 10380 3357 10406 3375
rect 10446 3357 10448 3375
rect 10448 3357 10480 3375
rect 10520 3357 10550 3375
rect 10550 3357 10554 3375
rect 10594 3357 10618 3375
rect 10618 3357 10628 3375
rect 10668 3357 10686 3375
rect 10686 3357 10702 3375
rect 10742 3357 10754 3375
rect 10754 3357 10776 3375
rect 10816 3357 10822 3375
rect 10822 3357 10850 3375
rect 10298 3341 10332 3357
rect 10372 3341 10406 3357
rect 10446 3341 10480 3357
rect 10520 3341 10554 3357
rect 10594 3341 10628 3357
rect 10668 3341 10702 3357
rect 10742 3341 10776 3357
rect 10816 3341 10850 3357
rect 10890 3341 10924 3375
rect 10964 3357 10992 3375
rect 10992 3357 10998 3375
rect 11038 3357 11060 3375
rect 11060 3357 11072 3375
rect 11112 3357 11128 3375
rect 11128 3357 11146 3375
rect 11186 3357 11196 3375
rect 11196 3357 11220 3375
rect 11260 3357 11264 3375
rect 11264 3357 11294 3375
rect 11334 3357 11366 3375
rect 11366 3357 11368 3375
rect 11408 3357 11434 3375
rect 11434 3357 11442 3375
rect 11482 3357 11502 3375
rect 11502 3357 11516 3375
rect 11556 3357 11570 3375
rect 11570 3357 11590 3375
rect 10964 3341 10998 3357
rect 11038 3341 11072 3357
rect 11112 3341 11146 3357
rect 11186 3341 11220 3357
rect 11260 3341 11294 3357
rect 11334 3341 11368 3357
rect 11408 3341 11442 3357
rect 11482 3341 11516 3357
rect 11556 3341 11590 3357
rect 8824 3286 8847 3303
rect 8847 3286 8858 3303
rect 8897 3286 8915 3303
rect 8915 3286 8931 3303
rect 8970 3286 8983 3303
rect 8983 3286 9004 3303
rect 9043 3286 9051 3303
rect 9051 3286 9077 3303
rect 9116 3286 9119 3303
rect 9119 3286 9150 3303
rect 9189 3286 9221 3303
rect 9221 3286 9223 3303
rect 9262 3286 9289 3303
rect 9289 3286 9296 3303
rect 9336 3286 9357 3303
rect 9357 3286 9370 3303
rect 9410 3286 9425 3303
rect 9425 3286 9444 3303
rect 9484 3286 9493 3303
rect 9493 3286 9518 3303
rect 9558 3286 9561 3303
rect 9561 3286 9592 3303
rect 9632 3286 9663 3303
rect 9663 3286 9666 3303
rect 9706 3286 9731 3303
rect 9731 3286 9740 3303
rect 9780 3286 9799 3303
rect 9799 3286 9814 3303
rect 9854 3286 9867 3303
rect 9867 3286 9888 3303
rect 9928 3286 9935 3303
rect 9935 3286 9962 3303
rect 10002 3286 10003 3303
rect 10003 3286 10036 3303
rect 10076 3286 10105 3303
rect 10105 3286 10110 3303
rect 10150 3286 10173 3303
rect 10173 3286 10184 3303
rect 10224 3286 10241 3303
rect 10241 3286 10258 3303
rect 8824 3269 8858 3286
rect 8897 3269 8931 3286
rect 8970 3269 9004 3286
rect 9043 3269 9077 3286
rect 9116 3269 9150 3286
rect 9189 3269 9223 3286
rect 9262 3269 9296 3286
rect 9336 3269 9370 3286
rect 9410 3269 9444 3286
rect 9484 3269 9518 3286
rect 9558 3269 9592 3286
rect 9632 3269 9666 3286
rect 9706 3269 9740 3286
rect 9780 3269 9814 3286
rect 9854 3269 9888 3286
rect 9928 3269 9962 3286
rect 10002 3269 10036 3286
rect 10076 3269 10110 3286
rect 10150 3269 10184 3286
rect 10224 3269 10258 3286
rect 10298 3287 10312 3303
rect 10312 3287 10332 3303
rect 10372 3287 10380 3303
rect 10380 3287 10406 3303
rect 10446 3287 10448 3303
rect 10448 3287 10480 3303
rect 10520 3287 10550 3303
rect 10550 3287 10554 3303
rect 10594 3287 10618 3303
rect 10618 3287 10628 3303
rect 10668 3287 10686 3303
rect 10686 3287 10702 3303
rect 10742 3287 10754 3303
rect 10754 3287 10776 3303
rect 10816 3287 10822 3303
rect 10822 3287 10850 3303
rect 10298 3269 10332 3287
rect 10372 3269 10406 3287
rect 10446 3269 10480 3287
rect 10520 3269 10554 3287
rect 10594 3269 10628 3287
rect 10668 3269 10702 3287
rect 10742 3269 10776 3287
rect 10816 3269 10850 3287
rect 10890 3269 10924 3303
rect 10964 3287 10992 3303
rect 10992 3287 10998 3303
rect 11038 3287 11060 3303
rect 11060 3287 11072 3303
rect 11112 3287 11128 3303
rect 11128 3287 11146 3303
rect 11186 3287 11196 3303
rect 11196 3287 11220 3303
rect 11260 3287 11264 3303
rect 11264 3287 11294 3303
rect 11334 3287 11366 3303
rect 11366 3287 11368 3303
rect 11408 3287 11434 3303
rect 11434 3287 11442 3303
rect 11482 3287 11502 3303
rect 11502 3287 11516 3303
rect 11556 3287 11570 3303
rect 11570 3287 11590 3303
rect 10964 3269 10998 3287
rect 11038 3269 11072 3287
rect 11112 3269 11146 3287
rect 11186 3269 11220 3287
rect 11260 3269 11294 3287
rect 11334 3269 11368 3287
rect 11408 3269 11442 3287
rect 11482 3269 11516 3287
rect 11556 3269 11590 3287
rect 12594 3453 12628 3471
rect 12667 3453 12701 3471
rect 12740 3453 12774 3471
rect 12813 3453 12847 3471
rect 12886 3453 12920 3471
rect 12959 3453 12993 3471
rect 13032 3453 13066 3471
rect 12594 3437 12595 3453
rect 12595 3437 12628 3453
rect 12667 3437 12697 3453
rect 12697 3437 12701 3453
rect 12740 3437 12765 3453
rect 12765 3437 12774 3453
rect 12813 3437 12833 3453
rect 12833 3437 12847 3453
rect 12886 3437 12901 3453
rect 12901 3437 12920 3453
rect 12959 3437 12969 3453
rect 12969 3437 12993 3453
rect 13032 3437 13037 3453
rect 13037 3437 13066 3453
rect 13105 3437 13139 3471
rect 13178 3453 13212 3471
rect 13251 3453 13285 3471
rect 13324 3453 13358 3471
rect 13178 3437 13207 3453
rect 13207 3437 13212 3453
rect 13251 3437 13275 3453
rect 13275 3437 13285 3453
rect 13324 3437 13343 3453
rect 13343 3437 13358 3453
rect 13397 3437 13431 3471
rect 13470 3437 13504 3471
rect 13543 3437 13577 3471
rect 13616 3437 13650 3471
rect 13689 3437 13723 3471
rect 13762 3437 13796 3471
rect 13835 3437 13869 3471
rect 13908 3437 13942 3471
rect 13981 3437 14015 3471
rect 14054 3437 14088 3471
rect 14127 3437 14161 3471
rect 14200 3437 14234 3471
rect 14273 3437 14307 3471
rect 14346 3437 14380 3471
rect 14419 3437 14453 3471
rect 14492 3437 14526 3471
rect 14565 3437 14599 3471
rect 14638 3437 14672 3471
rect 14711 3437 14745 3471
rect 14784 3437 14818 3471
rect 14857 3437 14891 3471
rect 14930 3437 14964 3471
rect 15003 3437 15037 3471
rect 15076 3437 15110 3471
rect 15149 3437 15183 3471
rect 15222 3437 15256 3471
rect 15295 3437 15329 3471
rect 15368 3437 15402 3471
rect 15441 3437 15475 3471
rect 15514 3437 15548 3471
rect 15587 3437 15621 3471
rect 15660 3437 15694 3471
rect 15733 3437 15767 3471
rect 15806 3437 15840 3471
rect 15879 3437 15913 3471
rect 15952 3437 15986 3471
rect 16025 3437 16059 3471
rect 16098 3437 16132 3471
rect 16171 3437 16205 3471
rect 16244 3437 16278 3471
rect 16317 3437 16351 3471
rect 16390 3437 16424 3471
rect 12594 3383 12628 3399
rect 12667 3383 12701 3399
rect 12740 3383 12774 3399
rect 12813 3383 12847 3399
rect 12886 3383 12920 3399
rect 12959 3383 12993 3399
rect 13032 3383 13066 3399
rect 12594 3365 12595 3383
rect 12595 3365 12628 3383
rect 12667 3365 12697 3383
rect 12697 3365 12701 3383
rect 12740 3365 12765 3383
rect 12765 3365 12774 3383
rect 12813 3365 12833 3383
rect 12833 3365 12847 3383
rect 12886 3365 12901 3383
rect 12901 3365 12920 3383
rect 12959 3365 12969 3383
rect 12969 3365 12993 3383
rect 13032 3365 13037 3383
rect 13037 3365 13066 3383
rect 13105 3365 13139 3399
rect 13178 3383 13212 3399
rect 13251 3383 13285 3399
rect 13324 3383 13358 3399
rect 13178 3365 13207 3383
rect 13207 3365 13212 3383
rect 13251 3365 13275 3383
rect 13275 3365 13285 3383
rect 13324 3365 13343 3383
rect 13343 3365 13358 3383
rect 13397 3365 13431 3399
rect 13470 3365 13504 3399
rect 13543 3365 13577 3399
rect 13616 3365 13650 3399
rect 13689 3365 13723 3399
rect 13762 3365 13796 3399
rect 13835 3365 13869 3399
rect 13908 3365 13942 3399
rect 13981 3365 14015 3399
rect 14054 3365 14088 3399
rect 14127 3365 14161 3399
rect 14200 3365 14234 3399
rect 14273 3365 14307 3399
rect 14346 3365 14380 3399
rect 14419 3365 14453 3399
rect 14492 3365 14526 3399
rect 14565 3365 14599 3399
rect 14638 3365 14672 3399
rect 14711 3365 14745 3399
rect 14784 3365 14818 3399
rect 14857 3365 14891 3399
rect 14930 3365 14964 3399
rect 15003 3365 15037 3399
rect 15076 3365 15110 3399
rect 15149 3365 15183 3399
rect 15222 3365 15256 3399
rect 15295 3365 15329 3399
rect 15368 3365 15402 3399
rect 15441 3365 15475 3399
rect 15514 3365 15548 3399
rect 15587 3365 15621 3399
rect 15660 3365 15694 3399
rect 15733 3365 15767 3399
rect 15806 3365 15840 3399
rect 15879 3365 15913 3399
rect 15952 3365 15986 3399
rect 16025 3365 16059 3399
rect 16098 3365 16132 3399
rect 16171 3365 16205 3399
rect 16244 3365 16278 3399
rect 16317 3365 16351 3399
rect 16390 3365 16424 3399
rect 12594 3313 12628 3327
rect 12667 3313 12701 3327
rect 12740 3313 12774 3327
rect 12813 3313 12847 3327
rect 12886 3313 12920 3327
rect 12959 3313 12993 3327
rect 13032 3313 13066 3327
rect 12594 3293 12595 3313
rect 12595 3293 12628 3313
rect 12667 3293 12697 3313
rect 12697 3293 12701 3313
rect 12740 3293 12765 3313
rect 12765 3293 12774 3313
rect 12813 3293 12833 3313
rect 12833 3293 12847 3313
rect 12886 3293 12901 3313
rect 12901 3293 12920 3313
rect 12959 3293 12969 3313
rect 12969 3293 12993 3313
rect 13032 3293 13037 3313
rect 13037 3293 13066 3313
rect 13105 3293 13139 3327
rect 13178 3313 13212 3327
rect 13251 3313 13285 3327
rect 13324 3313 13358 3327
rect 13178 3293 13207 3313
rect 13207 3293 13212 3313
rect 13251 3293 13275 3313
rect 13275 3293 13285 3313
rect 13324 3293 13343 3313
rect 13343 3293 13358 3313
rect 13397 3293 13431 3327
rect 13470 3293 13504 3327
rect 13543 3293 13577 3327
rect 13616 3293 13650 3327
rect 13689 3293 13723 3327
rect 13762 3293 13796 3327
rect 13835 3293 13869 3327
rect 13908 3293 13942 3327
rect 13981 3293 14015 3327
rect 14054 3293 14088 3327
rect 14127 3293 14161 3327
rect 14200 3293 14234 3327
rect 14273 3293 14307 3327
rect 14346 3293 14380 3327
rect 14419 3293 14453 3327
rect 14492 3293 14526 3327
rect 14565 3293 14599 3327
rect 14638 3293 14672 3327
rect 14711 3293 14745 3327
rect 14784 3293 14818 3327
rect 14857 3293 14891 3327
rect 14930 3293 14964 3327
rect 15003 3293 15037 3327
rect 15076 3293 15110 3327
rect 15149 3293 15183 3327
rect 15222 3293 15256 3327
rect 15295 3293 15329 3327
rect 15368 3293 15402 3327
rect 15441 3293 15475 3327
rect 15514 3293 15548 3327
rect 15587 3293 15621 3327
rect 15660 3293 15694 3327
rect 15733 3293 15767 3327
rect 15806 3293 15840 3327
rect 15879 3293 15913 3327
rect 15952 3293 15986 3327
rect 16025 3293 16059 3327
rect 16098 3293 16132 3327
rect 16171 3293 16205 3327
rect 16244 3293 16278 3327
rect 16317 3293 16351 3327
rect 16390 3293 16424 3327
rect 12594 3243 12628 3255
rect 12667 3243 12701 3255
rect 12740 3243 12774 3255
rect 12813 3243 12847 3255
rect 12886 3243 12920 3255
rect 12959 3243 12993 3255
rect 13032 3243 13066 3255
rect 12594 3221 12595 3243
rect 12595 3221 12628 3243
rect 12667 3221 12697 3243
rect 12697 3221 12701 3243
rect 12740 3221 12765 3243
rect 12765 3221 12774 3243
rect 12813 3221 12833 3243
rect 12833 3221 12847 3243
rect 12886 3221 12901 3243
rect 12901 3221 12920 3243
rect 12959 3221 12969 3243
rect 12969 3221 12993 3243
rect 13032 3221 13037 3243
rect 13037 3221 13066 3243
rect 13105 3221 13139 3255
rect 13178 3243 13212 3255
rect 13251 3243 13285 3255
rect 13324 3243 13358 3255
rect 13178 3221 13207 3243
rect 13207 3221 13212 3243
rect 13251 3221 13275 3243
rect 13275 3221 13285 3243
rect 13324 3221 13343 3243
rect 13343 3221 13358 3243
rect 13397 3221 13431 3255
rect 13470 3221 13504 3255
rect 13543 3221 13577 3255
rect 13616 3221 13650 3255
rect 13689 3221 13723 3255
rect 13762 3221 13796 3255
rect 13835 3221 13869 3255
rect 13908 3221 13942 3255
rect 13981 3221 14015 3255
rect 14054 3221 14088 3255
rect 14127 3221 14161 3255
rect 14200 3221 14234 3255
rect 14273 3221 14307 3255
rect 14346 3221 14380 3255
rect 14419 3221 14453 3255
rect 14492 3221 14526 3255
rect 14565 3221 14599 3255
rect 14638 3221 14672 3255
rect 14711 3221 14745 3255
rect 14784 3221 14818 3255
rect 14857 3221 14891 3255
rect 14930 3221 14964 3255
rect 15003 3221 15037 3255
rect 15076 3221 15110 3255
rect 15149 3221 15183 3255
rect 15222 3221 15256 3255
rect 15295 3221 15329 3255
rect 15368 3221 15402 3255
rect 15441 3221 15475 3255
rect 15514 3221 15548 3255
rect 15587 3221 15621 3255
rect 15660 3221 15694 3255
rect 15733 3221 15767 3255
rect 15806 3221 15840 3255
rect 15879 3221 15913 3255
rect 15952 3221 15986 3255
rect 16025 3221 16059 3255
rect 16098 3221 16132 3255
rect 16171 3221 16205 3255
rect 16244 3221 16278 3255
rect 16317 3221 16351 3255
rect 16390 3221 16424 3255
rect 23593 3415 23597 3449
rect 23597 3415 23627 3449
rect 23665 3415 23699 3449
rect 23737 3415 23767 3449
rect 23767 3415 23771 3449
rect 23593 3342 23597 3376
rect 23597 3342 23627 3376
rect 23665 3342 23699 3376
rect 23737 3342 23767 3376
rect 23767 3342 23771 3376
rect 23593 3269 23597 3303
rect 23597 3269 23627 3303
rect 23665 3269 23699 3303
rect 23737 3269 23767 3303
rect 23767 3269 23771 3303
rect 23593 3196 23597 3230
rect 23597 3196 23627 3230
rect 23665 3196 23699 3230
rect 23737 3196 23767 3230
rect 23767 3196 23771 3230
rect 23593 3122 23597 3156
rect 23597 3122 23627 3156
rect 23665 3122 23699 3156
rect 23737 3122 23767 3156
rect 23767 3122 23771 3156
rect 23593 3048 23597 3082
rect 23597 3048 23627 3082
rect 23665 3048 23699 3082
rect 23737 3048 23767 3082
rect 23767 3048 23771 3082
rect 23593 2974 23597 3008
rect 23597 2974 23627 3008
rect 23665 2974 23699 3008
rect 23737 2974 23767 3008
rect 23767 2974 23771 3008
rect 23593 2900 23597 2934
rect 23597 2900 23627 2934
rect 23665 2900 23699 2934
rect 23737 2900 23767 2934
rect 23767 2900 23771 2934
rect 23593 2826 23597 2860
rect 23597 2826 23627 2860
rect 23665 2826 23699 2860
rect 23737 2826 23767 2860
rect 23767 2826 23771 2860
rect 23593 2752 23597 2786
rect 23597 2752 23627 2786
rect 23665 2752 23699 2786
rect 23737 2752 23767 2786
rect 23767 2752 23771 2786
rect 11198 2692 11232 2702
rect 11272 2692 11306 2702
rect 11346 2692 11380 2702
rect 11420 2692 11454 2702
rect 11494 2692 11528 2702
rect 11568 2692 11602 2702
rect 11198 2668 11230 2692
rect 11230 2668 11232 2692
rect 11272 2668 11298 2692
rect 11298 2668 11306 2692
rect 11346 2668 11366 2692
rect 11366 2668 11380 2692
rect 11420 2668 11434 2692
rect 11434 2668 11454 2692
rect 11494 2668 11502 2692
rect 11502 2668 11528 2692
rect 11568 2668 11570 2692
rect 11570 2668 11602 2692
rect 11642 2699 11676 2702
rect 11716 2699 11750 2702
rect 11790 2699 11824 2702
rect 11864 2699 11898 2702
rect 11938 2699 11972 2702
rect 12012 2699 12046 2702
rect 12087 2699 12121 2702
rect 11642 2668 11652 2699
rect 11652 2668 11676 2699
rect 11716 2668 11720 2699
rect 11720 2668 11750 2699
rect 11790 2668 11822 2699
rect 11822 2668 11824 2699
rect 11864 2668 11890 2699
rect 11890 2668 11898 2699
rect 11938 2668 11958 2699
rect 11958 2668 11972 2699
rect 12012 2668 12026 2699
rect 12026 2668 12046 2699
rect 12087 2668 12094 2699
rect 12094 2668 12121 2699
rect 12162 2668 12196 2702
rect 12237 2699 12271 2702
rect 12312 2699 12346 2702
rect 12387 2699 12421 2702
rect 12462 2699 12496 2702
rect 12237 2668 12264 2699
rect 12264 2668 12271 2699
rect 12312 2668 12332 2699
rect 12332 2668 12346 2699
rect 12387 2668 12400 2699
rect 12400 2668 12421 2699
rect 12462 2668 12468 2699
rect 12468 2668 12496 2699
rect 12537 2668 12571 2702
rect 12612 2668 12646 2702
rect 12687 2668 12721 2702
rect 12762 2668 12796 2702
rect 12837 2668 12871 2702
rect 12912 2668 12946 2702
rect 12987 2668 13021 2702
rect 13062 2668 13096 2702
rect 13137 2668 13171 2702
rect 13212 2668 13246 2702
rect 11198 2623 11232 2630
rect 11272 2623 11306 2630
rect 11346 2623 11380 2630
rect 11420 2623 11454 2630
rect 11494 2623 11528 2630
rect 11568 2623 11602 2630
rect 11198 2596 11230 2623
rect 11230 2596 11232 2623
rect 11272 2596 11298 2623
rect 11298 2596 11306 2623
rect 11346 2596 11366 2623
rect 11366 2596 11380 2623
rect 11420 2596 11434 2623
rect 11434 2596 11454 2623
rect 11494 2596 11502 2623
rect 11502 2596 11528 2623
rect 11568 2596 11570 2623
rect 11570 2596 11602 2623
rect 11642 2629 11676 2630
rect 11716 2629 11750 2630
rect 11790 2629 11824 2630
rect 11864 2629 11898 2630
rect 11938 2629 11972 2630
rect 12012 2629 12046 2630
rect 12087 2629 12121 2630
rect 11642 2596 11652 2629
rect 11652 2596 11676 2629
rect 11716 2596 11720 2629
rect 11720 2596 11750 2629
rect 11790 2596 11822 2629
rect 11822 2596 11824 2629
rect 11864 2596 11890 2629
rect 11890 2596 11898 2629
rect 11938 2596 11958 2629
rect 11958 2596 11972 2629
rect 12012 2596 12026 2629
rect 12026 2596 12046 2629
rect 12087 2596 12094 2629
rect 12094 2596 12121 2629
rect 12162 2596 12196 2630
rect 12237 2629 12271 2630
rect 12312 2629 12346 2630
rect 12387 2629 12421 2630
rect 12462 2629 12496 2630
rect 12237 2596 12264 2629
rect 12264 2596 12271 2629
rect 12312 2596 12332 2629
rect 12332 2596 12346 2629
rect 12387 2596 12400 2629
rect 12400 2596 12421 2629
rect 12462 2596 12468 2629
rect 12468 2596 12496 2629
rect 12537 2596 12571 2630
rect 12612 2620 12646 2630
rect 12687 2620 12721 2630
rect 12762 2620 12796 2630
rect 12837 2620 12871 2630
rect 12912 2620 12946 2630
rect 12987 2620 13021 2630
rect 13062 2620 13096 2630
rect 13137 2620 13171 2630
rect 13212 2620 13246 2630
rect 12612 2596 12641 2620
rect 12641 2596 12646 2620
rect 12687 2596 12709 2620
rect 12709 2596 12721 2620
rect 12762 2596 12777 2620
rect 12777 2596 12796 2620
rect 12837 2596 12845 2620
rect 12845 2596 12871 2620
rect 12912 2596 12913 2620
rect 12913 2596 12946 2620
rect 12987 2596 13015 2620
rect 13015 2596 13021 2620
rect 13062 2596 13083 2620
rect 13083 2596 13096 2620
rect 13137 2596 13151 2620
rect 13151 2596 13171 2620
rect 13212 2596 13219 2620
rect 13219 2596 13246 2620
rect 11198 2554 11232 2558
rect 11272 2554 11306 2558
rect 11346 2554 11380 2558
rect 11420 2554 11454 2558
rect 11494 2554 11528 2558
rect 11568 2554 11602 2558
rect 11198 2524 11230 2554
rect 11230 2524 11232 2554
rect 11272 2524 11298 2554
rect 11298 2524 11306 2554
rect 11346 2524 11366 2554
rect 11366 2524 11380 2554
rect 11420 2524 11434 2554
rect 11434 2524 11454 2554
rect 11494 2524 11502 2554
rect 11502 2524 11528 2554
rect 11568 2524 11570 2554
rect 11570 2524 11602 2554
rect 11642 2525 11652 2558
rect 11652 2525 11676 2558
rect 11716 2525 11720 2558
rect 11720 2525 11750 2558
rect 11790 2525 11822 2558
rect 11822 2525 11824 2558
rect 11864 2525 11890 2558
rect 11890 2525 11898 2558
rect 11938 2525 11958 2558
rect 11958 2525 11972 2558
rect 12012 2525 12026 2558
rect 12026 2525 12046 2558
rect 12087 2525 12094 2558
rect 12094 2525 12121 2558
rect 11642 2524 11676 2525
rect 11716 2524 11750 2525
rect 11790 2524 11824 2525
rect 11864 2524 11898 2525
rect 11938 2524 11972 2525
rect 12012 2524 12046 2525
rect 12087 2524 12121 2525
rect 12162 2524 12196 2558
rect 12237 2525 12264 2558
rect 12264 2525 12271 2558
rect 12312 2525 12332 2558
rect 12332 2525 12346 2558
rect 12387 2525 12400 2558
rect 12400 2525 12421 2558
rect 12462 2525 12468 2558
rect 12468 2525 12496 2558
rect 12237 2524 12271 2525
rect 12312 2524 12346 2525
rect 12387 2524 12421 2525
rect 12462 2524 12496 2525
rect 12537 2524 12571 2558
rect 12612 2551 12646 2558
rect 12687 2551 12721 2558
rect 12762 2551 12796 2558
rect 12837 2551 12871 2558
rect 12912 2551 12946 2558
rect 12987 2551 13021 2558
rect 13062 2551 13096 2558
rect 13137 2551 13171 2558
rect 13212 2551 13246 2558
rect 12612 2524 12641 2551
rect 12641 2524 12646 2551
rect 12687 2524 12709 2551
rect 12709 2524 12721 2551
rect 12762 2524 12777 2551
rect 12777 2524 12796 2551
rect 12837 2524 12845 2551
rect 12845 2524 12871 2551
rect 12912 2524 12913 2551
rect 12913 2524 12946 2551
rect 12987 2524 13015 2551
rect 13015 2524 13021 2551
rect 13062 2524 13083 2551
rect 13083 2524 13096 2551
rect 13137 2524 13151 2551
rect 13151 2524 13171 2551
rect 13212 2524 13219 2551
rect 13219 2524 13246 2551
rect 11319 2140 11713 2154
rect 11752 2140 11786 2154
rect 11825 2140 11859 2154
rect 11898 2140 11932 2154
rect 11971 2140 12005 2154
rect 12044 2140 12078 2154
rect 12117 2140 12151 2154
rect 12190 2140 12224 2154
rect 12263 2140 12297 2154
rect 12336 2140 12370 2154
rect 12409 2140 12443 2154
rect 12482 2140 12516 2154
rect 11319 2106 11332 2140
rect 11332 2106 11366 2140
rect 11366 2106 11400 2140
rect 11400 2106 11434 2140
rect 11434 2106 11468 2140
rect 11468 2106 11502 2140
rect 11502 2106 11536 2140
rect 11536 2106 11570 2140
rect 11570 2106 11652 2140
rect 11652 2106 11686 2140
rect 11686 2106 11713 2140
rect 11752 2120 11754 2140
rect 11754 2120 11786 2140
rect 11825 2120 11856 2140
rect 11856 2120 11859 2140
rect 11898 2120 11924 2140
rect 11924 2120 11932 2140
rect 11971 2120 11992 2140
rect 11992 2120 12005 2140
rect 12044 2120 12060 2140
rect 12060 2120 12078 2140
rect 12117 2120 12128 2140
rect 12128 2120 12151 2140
rect 12190 2120 12196 2140
rect 12196 2120 12224 2140
rect 12263 2120 12264 2140
rect 12264 2120 12297 2140
rect 12336 2120 12366 2140
rect 12366 2120 12370 2140
rect 12409 2120 12434 2140
rect 12434 2120 12443 2140
rect 12482 2120 12502 2140
rect 12502 2120 12516 2140
rect 12555 2137 12589 2154
rect 12628 2137 12662 2154
rect 12701 2137 12735 2154
rect 12774 2137 12808 2154
rect 12847 2137 12881 2154
rect 12920 2137 12954 2154
rect 12993 2137 13027 2154
rect 13066 2137 13100 2154
rect 13139 2137 13173 2154
rect 13212 2137 13246 2154
rect 12555 2120 12573 2137
rect 12573 2120 12589 2137
rect 12628 2120 12641 2137
rect 12641 2120 12662 2137
rect 12701 2120 12709 2137
rect 12709 2120 12735 2137
rect 12774 2120 12777 2137
rect 12777 2120 12808 2137
rect 11319 2071 11713 2106
rect 12847 2120 12879 2137
rect 12879 2120 12881 2137
rect 12920 2120 12947 2137
rect 12947 2120 12954 2137
rect 12993 2120 13015 2137
rect 13015 2120 13027 2137
rect 13066 2120 13083 2137
rect 13083 2120 13100 2137
rect 13139 2120 13151 2137
rect 13151 2120 13173 2137
rect 13212 2120 13219 2137
rect 13219 2120 13246 2137
rect 11752 2071 11786 2082
rect 11825 2071 11859 2082
rect 11898 2071 11932 2082
rect 11971 2071 12005 2082
rect 12044 2071 12078 2082
rect 12117 2071 12151 2082
rect 12190 2071 12224 2082
rect 12263 2071 12297 2082
rect 12336 2071 12370 2082
rect 12409 2071 12443 2082
rect 12482 2071 12516 2082
rect 11319 2037 11332 2071
rect 11332 2037 11366 2071
rect 11366 2037 11400 2071
rect 11400 2037 11434 2071
rect 11434 2037 11468 2071
rect 11468 2037 11502 2071
rect 11502 2037 11536 2071
rect 11536 2037 11570 2071
rect 11570 2037 11652 2071
rect 11652 2037 11686 2071
rect 11686 2037 11713 2071
rect 11752 2048 11754 2071
rect 11754 2048 11786 2071
rect 11825 2048 11856 2071
rect 11856 2048 11859 2071
rect 11898 2048 11924 2071
rect 11924 2048 11932 2071
rect 11971 2048 11992 2071
rect 11992 2048 12005 2071
rect 12044 2048 12060 2071
rect 12060 2048 12078 2071
rect 12117 2048 12128 2071
rect 12128 2048 12151 2071
rect 12190 2048 12196 2071
rect 12196 2048 12224 2071
rect 12263 2048 12264 2071
rect 12264 2048 12297 2071
rect 12336 2048 12366 2071
rect 12366 2048 12370 2071
rect 12409 2048 12434 2071
rect 12434 2048 12443 2071
rect 12482 2048 12502 2071
rect 12502 2048 12516 2071
rect 12555 2068 12589 2082
rect 12628 2068 12662 2082
rect 12701 2068 12735 2082
rect 12774 2068 12808 2082
rect 12847 2068 12881 2082
rect 12920 2068 12954 2082
rect 12993 2068 13027 2082
rect 13066 2068 13100 2082
rect 13139 2068 13173 2082
rect 13212 2068 13246 2082
rect 23593 2678 23597 2712
rect 23597 2678 23627 2712
rect 23665 2678 23699 2712
rect 23737 2678 23767 2712
rect 23767 2678 23771 2712
rect 23593 2604 23597 2638
rect 23597 2604 23627 2638
rect 23665 2604 23699 2638
rect 23737 2604 23767 2638
rect 23767 2604 23771 2638
rect 23593 2530 23597 2564
rect 23597 2530 23627 2564
rect 23665 2530 23699 2564
rect 23737 2530 23767 2564
rect 23767 2530 23771 2564
rect 23593 2456 23597 2490
rect 23597 2456 23627 2490
rect 23665 2456 23699 2490
rect 23737 2456 23767 2490
rect 23767 2456 23771 2490
rect 23593 2382 23597 2416
rect 23597 2382 23627 2416
rect 23665 2382 23699 2416
rect 23737 2382 23767 2416
rect 23767 2382 23771 2416
rect 23593 2308 23597 2342
rect 23597 2308 23627 2342
rect 23665 2308 23699 2342
rect 23737 2308 23767 2342
rect 23767 2308 23771 2342
rect 23593 2234 23597 2268
rect 23597 2234 23627 2268
rect 23665 2234 23699 2268
rect 23737 2234 23767 2268
rect 23767 2234 23771 2268
rect 23593 2160 23597 2194
rect 23597 2160 23627 2194
rect 23665 2160 23699 2194
rect 23737 2160 23767 2194
rect 23767 2160 23771 2194
rect 23593 2110 23597 2120
rect 23597 2110 23627 2120
rect 23665 2110 23699 2120
rect 23737 2110 23767 2120
rect 23767 2110 23771 2120
rect 23593 2086 23627 2110
rect 23665 2086 23699 2110
rect 23737 2086 23771 2110
rect 12555 2048 12573 2068
rect 12573 2048 12589 2068
rect 12628 2048 12641 2068
rect 12641 2048 12662 2068
rect 12701 2048 12709 2068
rect 12709 2048 12735 2068
rect 12774 2048 12777 2068
rect 12777 2048 12808 2068
rect 11319 2002 11713 2037
rect 12847 2048 12879 2068
rect 12879 2048 12881 2068
rect 12920 2048 12947 2068
rect 12947 2048 12954 2068
rect 12993 2048 13015 2068
rect 13015 2048 13027 2068
rect 13066 2048 13083 2068
rect 13083 2048 13100 2068
rect 13139 2048 13151 2068
rect 13151 2048 13173 2068
rect 13212 2048 13219 2068
rect 13219 2048 13246 2068
rect 11752 2002 11786 2010
rect 11825 2002 11859 2010
rect 11898 2002 11932 2010
rect 11971 2002 12005 2010
rect 12044 2002 12078 2010
rect 12117 2002 12151 2010
rect 12190 2002 12224 2010
rect 12263 2002 12297 2010
rect 12336 2002 12370 2010
rect 12409 2002 12443 2010
rect 12482 2002 12516 2010
rect 8774 1968 8779 1975
rect 8779 1968 8808 1975
rect 8847 1968 8881 1975
rect 8920 1968 8949 1975
rect 8949 1968 8954 1975
rect 8993 1968 9017 1975
rect 9017 1968 9027 1975
rect 9066 1968 9085 1975
rect 9085 1968 9100 1975
rect 9139 1968 9153 1975
rect 9153 1968 9173 1975
rect 9212 1968 9221 1975
rect 9221 1968 9246 1975
rect 9285 1968 9289 1975
rect 9289 1968 9319 1975
rect 9358 1968 9391 1975
rect 9391 1968 9392 1975
rect 9431 1968 9459 1975
rect 9459 1968 9465 1975
rect 9504 1968 9527 1975
rect 9527 1968 9538 1975
rect 9577 1968 9595 1975
rect 9595 1968 9611 1975
rect 9650 1968 9663 1975
rect 9663 1968 9684 1975
rect 9723 1968 9731 1975
rect 9731 1968 9757 1975
rect 9796 1968 9799 1975
rect 9799 1968 9830 1975
rect 9869 1968 9901 1975
rect 9901 1968 9903 1975
rect 9942 1968 9969 1975
rect 9969 1968 9976 1975
rect 10015 1968 10037 1975
rect 10037 1968 10049 1975
rect 10088 1968 10105 1975
rect 10105 1968 10122 1975
rect 10161 1968 10173 1975
rect 10173 1968 10195 1975
rect 10234 1968 10241 1975
rect 10241 1968 10268 1975
rect 8774 1941 8808 1968
rect 8847 1941 8881 1968
rect 8920 1941 8954 1968
rect 8993 1941 9027 1968
rect 9066 1941 9100 1968
rect 9139 1941 9173 1968
rect 9212 1941 9246 1968
rect 9285 1941 9319 1968
rect 9358 1941 9392 1968
rect 9431 1941 9465 1968
rect 9504 1941 9538 1968
rect 9577 1941 9611 1968
rect 9650 1941 9684 1968
rect 9723 1941 9757 1968
rect 9796 1941 9830 1968
rect 9869 1941 9903 1968
rect 9942 1941 9976 1968
rect 10015 1941 10049 1968
rect 10088 1941 10122 1968
rect 10161 1941 10195 1968
rect 10234 1941 10268 1968
rect 10307 1968 10312 1975
rect 10312 1968 10341 1975
rect 10380 1968 10414 1975
rect 11319 1975 11332 2002
rect 10453 1968 10482 1975
rect 10482 1968 10487 1975
rect 10526 1968 10550 1975
rect 10550 1968 10560 1975
rect 10599 1968 10618 1975
rect 10618 1968 10652 1975
rect 10652 1968 10686 1975
rect 10686 1968 10720 1975
rect 10720 1968 10754 1975
rect 10754 1968 10788 1975
rect 10788 1968 10822 1975
rect 10822 1968 10856 1975
rect 10856 1968 10890 1975
rect 10890 1968 10924 1975
rect 10924 1968 10958 1975
rect 10958 1968 10992 1975
rect 10992 1968 11026 1975
rect 11026 1968 11060 1975
rect 11060 1968 11094 1975
rect 11094 1968 11128 1975
rect 11128 1968 11162 1975
rect 11162 1968 11196 1975
rect 11196 1968 11230 1975
rect 11230 1968 11264 1975
rect 11264 1968 11298 1975
rect 11298 1968 11332 1975
rect 11332 1968 11366 2002
rect 11366 1968 11400 2002
rect 11400 1968 11434 2002
rect 11434 1968 11468 2002
rect 11468 1968 11502 2002
rect 11502 1968 11536 2002
rect 11536 1968 11570 2002
rect 11570 1968 11652 2002
rect 11652 1968 11686 2002
rect 11686 1968 11713 2002
rect 11752 1976 11754 2002
rect 11754 1976 11786 2002
rect 11825 1976 11856 2002
rect 11856 1976 11859 2002
rect 11898 1976 11924 2002
rect 11924 1976 11932 2002
rect 11971 1976 11992 2002
rect 11992 1976 12005 2002
rect 12044 1976 12060 2002
rect 12060 1976 12078 2002
rect 12117 1976 12128 2002
rect 12128 1976 12151 2002
rect 12190 1976 12196 2002
rect 12196 1976 12224 2002
rect 12263 1976 12264 2002
rect 12264 1976 12297 2002
rect 12336 1976 12366 2002
rect 12366 1976 12370 2002
rect 12409 1976 12434 2002
rect 12434 1976 12443 2002
rect 12482 1976 12502 2002
rect 12502 1976 12516 2002
rect 12555 1999 12589 2010
rect 12628 1999 12662 2010
rect 12701 1999 12735 2010
rect 12774 1999 12808 2010
rect 12847 1999 12881 2010
rect 12920 1999 12954 2010
rect 12993 1999 13027 2010
rect 13066 1999 13100 2010
rect 13139 1999 13173 2010
rect 13212 1999 13246 2010
rect 12555 1976 12573 1999
rect 12573 1976 12589 1999
rect 12628 1976 12641 1999
rect 12641 1976 12662 1999
rect 12701 1976 12709 1999
rect 12709 1976 12735 1999
rect 12774 1976 12777 1999
rect 12777 1976 12808 1999
rect 10307 1941 10341 1968
rect 10380 1941 10414 1968
rect 10453 1941 10487 1968
rect 10526 1941 10560 1968
rect 10599 1933 11713 1968
rect 12847 1976 12879 1999
rect 12879 1976 12881 1999
rect 12920 1976 12947 1999
rect 12947 1976 12954 1999
rect 12993 1976 13015 1999
rect 13015 1976 13027 1999
rect 13066 1976 13083 1999
rect 13083 1976 13100 1999
rect 13139 1976 13151 1999
rect 13151 1976 13173 1999
rect 13212 1976 13219 1999
rect 13219 1976 13246 1999
rect 11752 1933 11786 1938
rect 11825 1933 11859 1938
rect 11898 1933 11932 1938
rect 11971 1933 12005 1938
rect 12044 1933 12078 1938
rect 12117 1933 12151 1938
rect 12190 1933 12224 1938
rect 12263 1933 12297 1938
rect 12336 1933 12370 1938
rect 12409 1933 12443 1938
rect 12482 1933 12516 1938
rect 8774 1899 8779 1903
rect 8779 1899 8808 1903
rect 8847 1899 8881 1903
rect 8920 1899 8949 1903
rect 8949 1899 8954 1903
rect 8993 1899 9017 1903
rect 9017 1899 9027 1903
rect 9066 1899 9085 1903
rect 9085 1899 9100 1903
rect 9139 1899 9153 1903
rect 9153 1899 9173 1903
rect 9212 1899 9221 1903
rect 9221 1899 9246 1903
rect 9285 1899 9289 1903
rect 9289 1899 9319 1903
rect 9358 1899 9391 1903
rect 9391 1899 9392 1903
rect 9431 1899 9459 1903
rect 9459 1899 9465 1903
rect 9504 1899 9527 1903
rect 9527 1899 9538 1903
rect 9577 1899 9595 1903
rect 9595 1899 9611 1903
rect 9650 1899 9663 1903
rect 9663 1899 9684 1903
rect 9723 1899 9731 1903
rect 9731 1899 9757 1903
rect 9796 1899 9799 1903
rect 9799 1899 9830 1903
rect 9869 1899 9901 1903
rect 9901 1899 9903 1903
rect 9942 1899 9969 1903
rect 9969 1899 9976 1903
rect 10015 1899 10037 1903
rect 10037 1899 10049 1903
rect 10088 1899 10105 1903
rect 10105 1899 10122 1903
rect 10161 1899 10173 1903
rect 10173 1899 10195 1903
rect 10234 1899 10241 1903
rect 10241 1899 10268 1903
rect 8774 1869 8808 1899
rect 8847 1869 8881 1899
rect 8920 1869 8954 1899
rect 8993 1869 9027 1899
rect 9066 1869 9100 1899
rect 9139 1869 9173 1899
rect 9212 1869 9246 1899
rect 9285 1869 9319 1899
rect 9358 1869 9392 1899
rect 9431 1869 9465 1899
rect 9504 1869 9538 1899
rect 9577 1869 9611 1899
rect 9650 1869 9684 1899
rect 9723 1869 9757 1899
rect 9796 1869 9830 1899
rect 9869 1869 9903 1899
rect 9942 1869 9976 1899
rect 10015 1869 10049 1899
rect 10088 1869 10122 1899
rect 10161 1869 10195 1899
rect 10234 1869 10268 1899
rect 10307 1899 10312 1903
rect 10312 1899 10341 1903
rect 10380 1899 10414 1903
rect 10453 1899 10482 1903
rect 10482 1899 10487 1903
rect 10526 1899 10550 1903
rect 10550 1899 10560 1903
rect 10599 1899 10618 1933
rect 10618 1899 10652 1933
rect 10652 1899 10686 1933
rect 10686 1899 10720 1933
rect 10720 1899 10754 1933
rect 10754 1899 10788 1933
rect 10788 1899 10822 1933
rect 10822 1899 10856 1933
rect 10856 1899 10890 1933
rect 10890 1899 10924 1933
rect 10924 1899 10958 1933
rect 10958 1899 10992 1933
rect 10992 1899 11026 1933
rect 11026 1899 11060 1933
rect 11060 1899 11094 1933
rect 11094 1899 11128 1933
rect 11128 1899 11162 1933
rect 11162 1899 11196 1933
rect 11196 1899 11230 1933
rect 11230 1899 11264 1933
rect 11264 1899 11298 1933
rect 11298 1899 11332 1933
rect 11332 1899 11366 1933
rect 11366 1899 11400 1933
rect 11400 1899 11434 1933
rect 11434 1899 11468 1933
rect 11468 1899 11502 1933
rect 11502 1899 11536 1933
rect 11536 1899 11570 1933
rect 11570 1899 11652 1933
rect 11652 1899 11686 1933
rect 11686 1899 11713 1933
rect 11752 1904 11754 1933
rect 11754 1904 11786 1933
rect 11825 1904 11856 1933
rect 11856 1904 11859 1933
rect 11898 1904 11924 1933
rect 11924 1904 11932 1933
rect 11971 1904 11992 1933
rect 11992 1904 12005 1933
rect 12044 1904 12060 1933
rect 12060 1904 12078 1933
rect 12117 1904 12128 1933
rect 12128 1904 12151 1933
rect 12190 1904 12196 1933
rect 12196 1904 12224 1933
rect 12263 1904 12264 1933
rect 12264 1904 12297 1933
rect 12336 1904 12366 1933
rect 12366 1904 12370 1933
rect 12409 1904 12434 1933
rect 12434 1904 12443 1933
rect 12482 1904 12502 1933
rect 12502 1904 12516 1933
rect 12555 1930 12589 1938
rect 12628 1930 12662 1938
rect 12701 1930 12735 1938
rect 12774 1930 12808 1938
rect 12847 1930 12881 1938
rect 12920 1930 12954 1938
rect 12993 1930 13027 1938
rect 13066 1930 13100 1938
rect 13139 1930 13173 1938
rect 13212 1930 13246 1938
rect 12555 1904 12573 1930
rect 12573 1904 12589 1930
rect 12628 1904 12641 1930
rect 12641 1904 12662 1930
rect 12701 1904 12709 1930
rect 12709 1904 12735 1930
rect 12774 1904 12777 1930
rect 12777 1904 12808 1930
rect 10307 1869 10341 1899
rect 10380 1869 10414 1899
rect 10453 1869 10487 1899
rect 10526 1869 10560 1899
rect 10599 1869 11713 1899
rect 12847 1904 12879 1930
rect 12879 1904 12881 1930
rect 12920 1904 12947 1930
rect 12947 1904 12954 1930
rect 12993 1904 13015 1930
rect 13015 1904 13027 1930
rect 13066 1904 13083 1930
rect 13083 1904 13100 1930
rect 13139 1904 13151 1930
rect 13151 1904 13173 1930
rect 13212 1904 13219 1930
rect 13219 1904 13246 1930
rect 11319 1864 11713 1869
rect 11752 1864 11786 1866
rect 11825 1864 11859 1866
rect 11898 1864 11932 1866
rect 11971 1864 12005 1866
rect 12044 1864 12078 1866
rect 12117 1864 12151 1866
rect 12190 1864 12224 1866
rect 12263 1864 12297 1866
rect 12336 1864 12370 1866
rect 12409 1864 12443 1866
rect 12482 1864 12516 1866
rect 11319 1830 11332 1864
rect 11332 1830 11366 1864
rect 11366 1830 11400 1864
rect 11400 1830 11434 1864
rect 11434 1830 11468 1864
rect 11468 1830 11502 1864
rect 11502 1830 11536 1864
rect 11536 1830 11570 1864
rect 11570 1830 11652 1864
rect 11652 1830 11686 1864
rect 11686 1830 11713 1864
rect 11752 1832 11754 1864
rect 11754 1832 11786 1864
rect 11825 1832 11856 1864
rect 11856 1832 11859 1864
rect 11898 1832 11924 1864
rect 11924 1832 11932 1864
rect 11971 1832 11992 1864
rect 11992 1832 12005 1864
rect 12044 1832 12060 1864
rect 12060 1832 12078 1864
rect 12117 1832 12128 1864
rect 12128 1832 12151 1864
rect 12190 1832 12196 1864
rect 12196 1832 12224 1864
rect 12263 1832 12264 1864
rect 12264 1832 12297 1864
rect 12336 1832 12366 1864
rect 12366 1832 12370 1864
rect 12409 1832 12434 1864
rect 12434 1832 12443 1864
rect 12482 1832 12502 1864
rect 12502 1832 12516 1864
rect 12555 1861 12589 1866
rect 12628 1861 12662 1866
rect 12701 1861 12735 1866
rect 12774 1861 12808 1866
rect 12847 1861 12881 1866
rect 12920 1861 12954 1866
rect 12993 1861 13027 1866
rect 13066 1861 13100 1866
rect 13139 1861 13173 1866
rect 13212 1861 13246 1866
rect 12555 1832 12573 1861
rect 12573 1832 12589 1861
rect 12628 1832 12662 1861
rect 12701 1832 12735 1861
rect 12774 1832 12808 1861
rect 12847 1832 12881 1861
rect 12920 1832 12954 1861
rect 12993 1832 13027 1861
rect 13066 1832 13100 1861
rect 13139 1832 13173 1861
rect 13212 1832 13246 1861
rect 1169 1738 1203 1772
rect 1241 1738 1275 1772
rect 1313 1738 1347 1772
rect 1385 1738 1419 1772
rect 1457 1738 1460 1772
rect 1460 1738 1491 1772
rect 1529 1759 1541 1772
rect 1541 1759 1563 1772
rect 1601 1762 1609 1772
rect 1609 1762 1635 1772
rect 1529 1738 1563 1759
rect 1601 1738 1635 1762
rect 1169 1665 1203 1699
rect 1241 1665 1275 1699
rect 1313 1665 1347 1699
rect 1385 1665 1419 1699
rect 1457 1665 1460 1699
rect 1460 1665 1491 1699
rect 1529 1691 1541 1699
rect 1541 1691 1563 1699
rect 1601 1693 1609 1699
rect 1609 1693 1635 1699
rect 1529 1665 1563 1691
rect 1601 1665 1635 1693
rect 1169 1592 1203 1626
rect 1241 1592 1275 1626
rect 1313 1592 1347 1626
rect 1385 1592 1419 1626
rect 1457 1592 1460 1626
rect 1460 1592 1491 1626
rect 1529 1623 1541 1626
rect 1541 1623 1563 1626
rect 1601 1624 1609 1626
rect 1609 1624 1635 1626
rect 1529 1592 1563 1623
rect 1601 1592 1635 1624
rect 11319 1795 11713 1830
rect 11319 1761 11332 1795
rect 11332 1761 11366 1795
rect 11366 1761 11400 1795
rect 11400 1761 11434 1795
rect 11434 1761 11468 1795
rect 11468 1761 11502 1795
rect 11502 1761 11536 1795
rect 11536 1761 11570 1795
rect 11570 1761 11652 1795
rect 11652 1761 11686 1795
rect 11686 1761 11713 1795
rect 11752 1761 11754 1794
rect 11754 1761 11786 1794
rect 11825 1761 11856 1794
rect 11856 1761 11859 1794
rect 11898 1761 11924 1794
rect 11924 1761 11932 1794
rect 11971 1761 11992 1794
rect 11992 1761 12005 1794
rect 12044 1761 12060 1794
rect 12060 1761 12078 1794
rect 12117 1761 12128 1794
rect 12128 1761 12151 1794
rect 12190 1761 12196 1794
rect 12196 1761 12224 1794
rect 12263 1761 12264 1794
rect 12264 1761 12297 1794
rect 12336 1761 12366 1794
rect 12366 1761 12370 1794
rect 12409 1761 12434 1794
rect 12434 1761 12443 1794
rect 12482 1761 12502 1794
rect 12502 1761 12516 1794
rect 11319 1760 11713 1761
rect 11752 1760 11786 1761
rect 11825 1760 11859 1761
rect 11898 1760 11932 1761
rect 11971 1760 12005 1761
rect 12044 1760 12078 1761
rect 12117 1760 12151 1761
rect 12190 1760 12224 1761
rect 12263 1760 12297 1761
rect 12336 1760 12370 1761
rect 12409 1760 12443 1761
rect 12482 1760 12516 1761
rect 12555 1760 12573 1794
rect 12573 1760 12589 1794
rect 12628 1760 12662 1794
rect 12701 1760 12735 1794
rect 12774 1760 12808 1794
rect 12847 1760 12881 1794
rect 12920 1760 12954 1794
rect 12993 1760 13027 1794
rect 13066 1760 13100 1794
rect 13139 1760 13173 1794
rect 13212 1760 13246 1794
rect 1169 1519 1203 1553
rect 1241 1519 1275 1553
rect 1313 1519 1347 1553
rect 1385 1519 1419 1553
rect 1457 1519 1460 1553
rect 1460 1519 1491 1553
rect 1529 1521 1563 1553
rect 1601 1521 1635 1553
rect 8434 1555 8446 1557
rect 8446 1555 8468 1557
rect 8509 1555 8516 1557
rect 8516 1555 8543 1557
rect 8584 1555 8586 1557
rect 8586 1555 8618 1557
rect 8659 1555 8692 1557
rect 8692 1555 8693 1557
rect 8734 1555 8762 1557
rect 8762 1555 8768 1557
rect 8809 1555 8832 1557
rect 8832 1555 8843 1557
rect 8884 1555 8902 1557
rect 8902 1555 8918 1557
rect 8959 1555 8972 1557
rect 8972 1555 8993 1557
rect 9034 1555 9043 1557
rect 9043 1555 9068 1557
rect 9109 1555 9114 1557
rect 9114 1555 9143 1557
rect 9184 1555 9185 1557
rect 9185 1555 9218 1557
rect 9259 1555 9290 1557
rect 9290 1555 9293 1557
rect 9334 1555 9361 1557
rect 9361 1555 9368 1557
rect 9409 1555 9432 1557
rect 9432 1555 9443 1557
rect 9484 1555 9503 1557
rect 9503 1555 9518 1557
rect 9559 1555 9574 1557
rect 9574 1555 9593 1557
rect 9634 1555 9645 1557
rect 9645 1555 9668 1557
rect 9709 1555 9716 1557
rect 9716 1555 9743 1557
rect 9784 1555 9787 1557
rect 9787 1555 9818 1557
rect 8434 1523 8468 1555
rect 8509 1523 8543 1555
rect 8584 1523 8618 1555
rect 8659 1523 8693 1555
rect 8734 1523 8768 1555
rect 8809 1523 8843 1555
rect 8884 1523 8918 1555
rect 8959 1523 8993 1555
rect 9034 1523 9068 1555
rect 9109 1523 9143 1555
rect 9184 1523 9218 1555
rect 9259 1523 9293 1555
rect 9334 1523 9368 1555
rect 9409 1523 9443 1555
rect 9484 1523 9518 1555
rect 9559 1523 9593 1555
rect 9634 1523 9668 1555
rect 9709 1523 9743 1555
rect 9784 1523 9818 1555
rect 9860 1523 9894 1557
rect 9936 1555 9966 1557
rect 9966 1555 9970 1557
rect 9936 1523 9970 1555
rect 10012 1523 10046 1557
rect 1529 1519 1531 1521
rect 1531 1519 1563 1521
rect 1601 1519 1634 1521
rect 1634 1519 1635 1521
rect 1169 1446 1203 1480
rect 1241 1446 1275 1480
rect 1313 1446 1347 1480
rect 1385 1446 1419 1480
rect 1457 1446 1460 1480
rect 1460 1446 1491 1480
rect 1529 1453 1563 1480
rect 1601 1453 1635 1480
rect 1683 1453 1717 1480
rect 1757 1453 1791 1480
rect 1831 1453 1865 1480
rect 1905 1453 1939 1480
rect 1529 1446 1531 1453
rect 1531 1446 1563 1453
rect 1601 1446 1634 1453
rect 1634 1446 1635 1453
rect 1683 1446 1703 1453
rect 1703 1446 1717 1453
rect 1757 1446 1772 1453
rect 1772 1446 1791 1453
rect 1831 1446 1841 1453
rect 1841 1446 1865 1453
rect 1905 1446 1910 1453
rect 1910 1446 1939 1453
rect 1979 1446 2013 1480
rect 2053 1453 2087 1480
rect 2127 1453 2161 1480
rect 2201 1453 2235 1480
rect 2276 1453 2310 1480
rect 2351 1453 2385 1480
rect 2426 1453 2460 1480
rect 2501 1453 2535 1480
rect 2576 1453 2610 1480
rect 2651 1453 2685 1480
rect 2726 1453 2760 1480
rect 2801 1453 2835 1480
rect 2053 1446 2083 1453
rect 2083 1446 2087 1453
rect 2127 1446 2152 1453
rect 2152 1446 2161 1453
rect 2201 1446 2221 1453
rect 2221 1446 2235 1453
rect 2276 1446 2290 1453
rect 2290 1446 2310 1453
rect 2351 1446 2359 1453
rect 2359 1446 2385 1453
rect 2426 1446 2428 1453
rect 2428 1446 2460 1453
rect 2501 1446 2531 1453
rect 2531 1446 2535 1453
rect 2576 1446 2600 1453
rect 2600 1446 2610 1453
rect 2651 1446 2669 1453
rect 2669 1446 2685 1453
rect 2726 1446 2738 1453
rect 2738 1446 2760 1453
rect 2801 1446 2807 1453
rect 2807 1446 2835 1453
rect 2876 1446 2910 1480
rect 2951 1453 2985 1480
rect 2951 1446 2980 1453
rect 2980 1446 2985 1453
rect 7117 1446 7151 1480
rect 7190 1446 7224 1480
rect 7263 1446 7297 1480
rect 7336 1446 7370 1480
rect 7409 1446 7443 1480
rect 7482 1446 7516 1480
rect 7555 1446 7589 1480
rect 7628 1446 7662 1480
rect 7701 1446 7735 1480
rect 7774 1446 7808 1480
rect 7847 1446 7881 1480
rect 7920 1446 7954 1480
rect 7993 1446 8027 1480
rect 8066 1446 8100 1480
rect 8140 1446 8174 1480
rect 8214 1446 8248 1480
rect 8288 1446 8322 1480
rect 8362 1446 8364 1480
rect 8364 1446 8396 1480
rect 8434 1453 8468 1485
rect 8509 1453 8543 1485
rect 8584 1453 8618 1485
rect 8659 1453 8693 1485
rect 8734 1453 8768 1485
rect 8809 1453 8843 1485
rect 8884 1453 8918 1485
rect 8959 1453 8993 1485
rect 9034 1453 9068 1485
rect 9109 1453 9143 1485
rect 9184 1453 9218 1485
rect 9259 1453 9293 1485
rect 9334 1453 9368 1485
rect 9409 1453 9443 1485
rect 9484 1453 9518 1485
rect 9559 1453 9593 1485
rect 9634 1453 9668 1485
rect 9709 1453 9743 1485
rect 9784 1453 9818 1485
rect 8434 1451 8446 1453
rect 8446 1451 8468 1453
rect 8509 1451 8516 1453
rect 8516 1451 8543 1453
rect 8584 1451 8586 1453
rect 8586 1451 8618 1453
rect 8659 1451 8692 1453
rect 8692 1451 8693 1453
rect 8734 1451 8762 1453
rect 8762 1451 8768 1453
rect 8809 1451 8832 1453
rect 8832 1451 8843 1453
rect 8884 1451 8902 1453
rect 8902 1451 8918 1453
rect 8959 1451 8972 1453
rect 8972 1451 8993 1453
rect 9034 1451 9043 1453
rect 9043 1451 9068 1453
rect 9109 1451 9114 1453
rect 9114 1451 9143 1453
rect 9184 1451 9185 1453
rect 9185 1451 9218 1453
rect 9259 1451 9290 1453
rect 9290 1451 9293 1453
rect 9334 1451 9361 1453
rect 9361 1451 9368 1453
rect 9409 1451 9432 1453
rect 9432 1451 9443 1453
rect 9484 1451 9503 1453
rect 9503 1451 9518 1453
rect 9559 1451 9574 1453
rect 9574 1451 9593 1453
rect 9634 1451 9645 1453
rect 9645 1451 9668 1453
rect 9709 1451 9716 1453
rect 9716 1451 9743 1453
rect 9784 1451 9787 1453
rect 9787 1451 9818 1453
rect 9860 1451 9894 1485
rect 9936 1453 9970 1485
rect 9936 1451 9966 1453
rect 9966 1451 9970 1453
rect 10012 1451 10046 1485
rect 23593 2027 23600 2046
rect 23600 2027 23627 2046
rect 23665 2027 23669 2046
rect 23669 2027 23699 2046
rect 23737 2027 23738 2046
rect 23738 2027 23771 2046
rect 23593 2012 23627 2027
rect 23665 2012 23699 2027
rect 23737 2012 23771 2027
rect 23593 1959 23600 1972
rect 23600 1959 23627 1972
rect 23665 1959 23669 1972
rect 23669 1959 23699 1972
rect 23737 1959 23738 1972
rect 23738 1959 23771 1972
rect 23593 1938 23627 1959
rect 23665 1938 23699 1959
rect 23737 1938 23771 1959
rect 14493 1491 14523 1494
rect 14523 1491 14527 1494
rect 14493 1460 14527 1491
rect 14566 1462 14591 1494
rect 14591 1462 14600 1494
rect 14566 1460 14600 1462
rect 14639 1460 14673 1494
rect 14712 1460 14746 1494
rect 14785 1460 14819 1494
rect 14858 1460 14892 1494
rect 14931 1460 14965 1494
rect 15004 1460 15038 1494
rect 15077 1460 15111 1494
rect 15150 1460 15184 1494
rect 15223 1460 15257 1494
rect 15296 1460 15330 1494
rect 15369 1460 15403 1494
rect 15442 1460 15476 1494
rect 15515 1460 15549 1494
rect 15588 1460 15622 1494
rect 15661 1460 15695 1494
rect 1683 1374 1717 1408
rect 1757 1374 1791 1408
rect 1831 1374 1865 1408
rect 1905 1374 1939 1408
rect 1979 1374 2013 1408
rect 2053 1374 2087 1408
rect 2127 1374 2161 1408
rect 2201 1374 2235 1408
rect 2276 1374 2310 1408
rect 2351 1374 2385 1408
rect 2426 1374 2460 1408
rect 2501 1374 2535 1408
rect 2576 1374 2610 1408
rect 2651 1374 2685 1408
rect 2726 1374 2760 1408
rect 2801 1374 2835 1408
rect 2876 1374 2910 1408
rect 2951 1374 2985 1408
rect 7117 1374 7151 1408
rect 7190 1374 7224 1408
rect 7263 1374 7297 1408
rect 7336 1374 7370 1408
rect 7409 1374 7443 1408
rect 7482 1374 7516 1408
rect 7555 1374 7589 1408
rect 7628 1374 7662 1408
rect 7701 1374 7735 1408
rect 7774 1374 7808 1408
rect 7847 1374 7881 1408
rect 7920 1374 7954 1408
rect 7993 1374 8027 1408
rect 8066 1374 8100 1408
rect 8140 1374 8174 1408
rect 8214 1374 8248 1408
rect 8288 1374 8322 1408
rect 8362 1374 8396 1408
rect 14493 1388 14527 1422
rect 14566 1392 14591 1422
rect 14591 1392 14600 1422
rect 14566 1388 14600 1392
rect 14639 1388 14673 1422
rect 14712 1388 14746 1422
rect 14785 1388 14819 1422
rect 14858 1388 14892 1422
rect 14931 1388 14965 1422
rect 15004 1388 15038 1422
rect 15077 1388 15111 1422
rect 15150 1388 15184 1422
rect 15223 1388 15257 1422
rect 15296 1388 15330 1422
rect 15369 1388 15403 1422
rect 15442 1388 15476 1422
rect 15515 1388 15549 1422
rect 15588 1388 15622 1422
rect 15661 1388 15695 1422
rect 800 1263 834 1297
rect 14493 1318 14527 1350
rect 14566 1322 14591 1350
rect 14591 1322 14600 1350
rect 14493 1316 14523 1318
rect 14523 1316 14527 1318
rect 14566 1316 14600 1322
rect 14639 1316 14673 1350
rect 14712 1316 14746 1350
rect 14785 1316 14819 1350
rect 14858 1316 14892 1350
rect 14931 1316 14965 1350
rect 15004 1316 15038 1350
rect 15077 1316 15111 1350
rect 15150 1316 15184 1350
rect 15223 1316 15257 1350
rect 15296 1316 15330 1350
rect 15369 1316 15403 1350
rect 15442 1316 15476 1350
rect 15515 1316 15549 1350
rect 15588 1316 15622 1350
rect 15661 1316 15695 1350
rect 728 1247 730 1259
rect 730 1247 762 1259
rect 728 1225 762 1247
rect 800 1190 834 1224
rect 728 1178 730 1187
rect 730 1178 762 1187
rect 728 1153 762 1178
rect 800 1117 834 1151
rect 728 1109 730 1115
rect 730 1109 762 1115
rect 728 1081 762 1109
rect 14493 1249 14527 1278
rect 14566 1252 14591 1278
rect 14591 1252 14600 1278
rect 14493 1244 14523 1249
rect 14523 1244 14527 1249
rect 14566 1244 14600 1252
rect 14639 1244 14673 1278
rect 14712 1244 14746 1278
rect 14785 1244 14819 1278
rect 14858 1244 14892 1278
rect 14931 1244 14965 1278
rect 15004 1244 15038 1278
rect 15077 1244 15111 1278
rect 15150 1244 15184 1278
rect 15223 1244 15257 1278
rect 15296 1244 15330 1278
rect 15369 1244 15403 1278
rect 15442 1244 15476 1278
rect 15515 1244 15549 1278
rect 15588 1244 15622 1278
rect 15661 1244 15695 1278
rect 14493 1179 14527 1206
rect 14566 1182 14591 1206
rect 14591 1182 14600 1206
rect 14493 1172 14523 1179
rect 14523 1172 14527 1179
rect 14566 1172 14600 1182
rect 14639 1172 14673 1206
rect 14712 1172 14746 1206
rect 14785 1172 14819 1206
rect 14858 1172 14892 1206
rect 14931 1172 14965 1206
rect 15004 1172 15038 1206
rect 15077 1172 15111 1206
rect 15150 1172 15184 1206
rect 15223 1172 15257 1206
rect 15296 1172 15330 1206
rect 15369 1172 15403 1206
rect 15442 1172 15476 1206
rect 15515 1172 15549 1206
rect 15588 1172 15622 1206
rect 15661 1172 15695 1206
rect 15734 1172 19563 1494
rect 19563 1483 19598 1494
rect 19598 1483 19632 1494
rect 19632 1483 19667 1494
rect 19667 1483 19701 1494
rect 19701 1483 19736 1494
rect 19736 1483 19770 1494
rect 19770 1483 19805 1494
rect 19805 1483 19839 1494
rect 19839 1483 19874 1494
rect 19874 1483 19908 1494
rect 19908 1483 19943 1494
rect 19943 1483 19977 1494
rect 19977 1483 20012 1494
rect 20012 1483 20046 1494
rect 20046 1483 20081 1494
rect 20081 1483 20115 1494
rect 20115 1483 20150 1494
rect 20150 1483 20184 1494
rect 20184 1483 20219 1494
rect 20219 1483 20253 1494
rect 20253 1483 20288 1494
rect 20288 1483 20322 1494
rect 20322 1483 20357 1494
rect 20357 1483 20391 1494
rect 20391 1483 20426 1494
rect 20426 1483 20460 1494
rect 20460 1483 20495 1494
rect 20495 1483 20529 1494
rect 20529 1483 20564 1494
rect 20564 1483 20598 1494
rect 20598 1483 20633 1494
rect 20633 1483 20667 1494
rect 20667 1483 20702 1494
rect 20702 1483 20736 1494
rect 20736 1483 20771 1494
rect 20771 1483 20805 1494
rect 20805 1483 20840 1494
rect 20840 1483 20874 1494
rect 20874 1483 20909 1494
rect 20909 1483 20943 1494
rect 20943 1483 20978 1494
rect 20978 1483 21012 1494
rect 21012 1483 21047 1494
rect 21047 1483 21081 1494
rect 21081 1483 21116 1494
rect 21116 1483 21150 1494
rect 21150 1483 21185 1494
rect 21185 1483 21219 1494
rect 21219 1483 21254 1494
rect 21254 1483 21288 1494
rect 21288 1483 21323 1494
rect 21323 1483 21357 1494
rect 21357 1483 21392 1494
rect 21392 1483 21426 1494
rect 21426 1483 21461 1494
rect 21461 1483 21495 1494
rect 21495 1483 21530 1494
rect 21530 1483 21564 1494
rect 21564 1483 21599 1494
rect 21599 1483 21633 1494
rect 21633 1483 21668 1494
rect 21668 1483 21702 1494
rect 21702 1483 21737 1494
rect 21737 1483 21771 1494
rect 21771 1483 21806 1494
rect 21806 1483 21840 1494
rect 21840 1483 21875 1494
rect 21875 1483 21909 1494
rect 21909 1483 21944 1494
rect 21944 1483 21978 1494
rect 21978 1483 22013 1494
rect 22013 1483 22047 1494
rect 22047 1483 22082 1494
rect 22082 1483 22116 1494
rect 22116 1483 22151 1494
rect 22151 1483 22185 1494
rect 22185 1483 22220 1494
rect 22220 1483 22254 1494
rect 22254 1483 22289 1494
rect 22289 1483 22323 1494
rect 22323 1483 22358 1494
rect 22358 1483 22392 1494
rect 22392 1483 22427 1494
rect 22427 1483 22461 1494
rect 22461 1483 22496 1494
rect 22496 1483 22530 1494
rect 22530 1483 22565 1494
rect 22565 1483 22599 1494
rect 22599 1483 22634 1494
rect 22634 1483 22668 1494
rect 22668 1483 22703 1494
rect 22703 1483 22737 1494
rect 22737 1483 22772 1494
rect 22772 1483 22806 1494
rect 22806 1483 22841 1494
rect 22841 1483 22875 1494
rect 22875 1483 22910 1494
rect 22910 1483 22944 1494
rect 22944 1483 22979 1494
rect 22979 1483 23013 1494
rect 23013 1483 23040 1494
rect 19563 1449 23040 1483
rect 19563 1415 19598 1449
rect 19598 1415 19632 1449
rect 19632 1415 19667 1449
rect 19667 1415 19701 1449
rect 19701 1415 19736 1449
rect 19736 1415 19770 1449
rect 19770 1415 19805 1449
rect 19805 1415 19839 1449
rect 19839 1415 19874 1449
rect 19874 1415 19908 1449
rect 19908 1415 19943 1449
rect 19943 1415 19977 1449
rect 19977 1415 20012 1449
rect 20012 1415 20046 1449
rect 20046 1415 20081 1449
rect 20081 1415 20115 1449
rect 20115 1415 20150 1449
rect 20150 1415 20184 1449
rect 20184 1415 20219 1449
rect 20219 1415 20253 1449
rect 20253 1415 20288 1449
rect 20288 1415 20322 1449
rect 20322 1415 20357 1449
rect 20357 1415 20391 1449
rect 20391 1415 20426 1449
rect 20426 1415 20460 1449
rect 20460 1415 20495 1449
rect 20495 1415 20529 1449
rect 20529 1415 20564 1449
rect 20564 1415 20598 1449
rect 20598 1415 20633 1449
rect 20633 1415 20667 1449
rect 20667 1415 20702 1449
rect 20702 1415 20736 1449
rect 20736 1415 20771 1449
rect 20771 1415 20805 1449
rect 20805 1415 20840 1449
rect 20840 1415 20874 1449
rect 20874 1415 20909 1449
rect 20909 1415 20943 1449
rect 20943 1415 20978 1449
rect 20978 1415 21012 1449
rect 21012 1415 21047 1449
rect 21047 1415 21081 1449
rect 21081 1415 21116 1449
rect 21116 1415 21150 1449
rect 21150 1415 21185 1449
rect 21185 1415 21219 1449
rect 21219 1415 21254 1449
rect 21254 1415 21288 1449
rect 21288 1415 21323 1449
rect 21323 1415 21357 1449
rect 21357 1415 21392 1449
rect 21392 1415 21426 1449
rect 21426 1415 21461 1449
rect 21461 1415 21495 1449
rect 21495 1415 21530 1449
rect 21530 1415 21564 1449
rect 21564 1415 21599 1449
rect 21599 1415 21633 1449
rect 21633 1415 21668 1449
rect 21668 1415 21702 1449
rect 21702 1415 21737 1449
rect 21737 1415 21771 1449
rect 21771 1415 21806 1449
rect 21806 1415 21840 1449
rect 21840 1415 21875 1449
rect 21875 1415 21909 1449
rect 21909 1415 21944 1449
rect 21944 1415 21978 1449
rect 21978 1415 22013 1449
rect 22013 1415 22047 1449
rect 22047 1415 22082 1449
rect 22082 1415 22116 1449
rect 22116 1415 22151 1449
rect 22151 1415 22185 1449
rect 22185 1415 22220 1449
rect 22220 1415 22254 1449
rect 22254 1415 22289 1449
rect 22289 1415 22323 1449
rect 22323 1415 22358 1449
rect 22358 1415 22392 1449
rect 22392 1415 22427 1449
rect 22427 1415 22461 1449
rect 22461 1415 22496 1449
rect 22496 1415 22530 1449
rect 22530 1415 22565 1449
rect 22565 1415 22599 1449
rect 22599 1415 22634 1449
rect 22634 1415 22668 1449
rect 22668 1415 22703 1449
rect 22703 1415 22737 1449
rect 22737 1415 22772 1449
rect 22772 1415 22806 1449
rect 22806 1415 22841 1449
rect 22841 1415 22875 1449
rect 22875 1415 22910 1449
rect 22910 1415 22944 1449
rect 22944 1415 22979 1449
rect 22979 1415 23013 1449
rect 23013 1415 23040 1449
rect 19563 1381 23040 1415
rect 19563 1347 19598 1381
rect 19598 1347 19632 1381
rect 19632 1347 19667 1381
rect 19667 1347 19701 1381
rect 19701 1347 19736 1381
rect 19736 1347 19770 1381
rect 19770 1347 19805 1381
rect 19805 1347 19839 1381
rect 19839 1347 19874 1381
rect 19874 1347 19908 1381
rect 19908 1347 19943 1381
rect 19943 1347 19977 1381
rect 19977 1347 20012 1381
rect 20012 1347 20046 1381
rect 20046 1347 20081 1381
rect 20081 1347 20115 1381
rect 20115 1347 20150 1381
rect 20150 1347 20184 1381
rect 20184 1347 20219 1381
rect 20219 1347 20253 1381
rect 20253 1347 20288 1381
rect 20288 1347 20322 1381
rect 20322 1347 20357 1381
rect 20357 1347 20391 1381
rect 20391 1347 20426 1381
rect 20426 1347 20460 1381
rect 20460 1347 20495 1381
rect 20495 1347 20529 1381
rect 20529 1347 20564 1381
rect 20564 1347 20598 1381
rect 20598 1347 20633 1381
rect 20633 1347 20667 1381
rect 20667 1347 20702 1381
rect 20702 1347 20736 1381
rect 20736 1347 20771 1381
rect 20771 1347 20805 1381
rect 20805 1347 20840 1381
rect 20840 1347 20874 1381
rect 20874 1347 20909 1381
rect 20909 1347 20943 1381
rect 20943 1347 20978 1381
rect 20978 1347 21012 1381
rect 21012 1347 21047 1381
rect 21047 1347 21081 1381
rect 21081 1347 21116 1381
rect 21116 1347 21150 1381
rect 21150 1347 21185 1381
rect 21185 1347 21219 1381
rect 21219 1347 21254 1381
rect 21254 1347 21288 1381
rect 21288 1347 21323 1381
rect 21323 1347 21357 1381
rect 21357 1347 21392 1381
rect 21392 1347 21426 1381
rect 21426 1347 21461 1381
rect 21461 1347 21495 1381
rect 21495 1347 21530 1381
rect 21530 1347 21564 1381
rect 21564 1347 21599 1381
rect 21599 1347 21633 1381
rect 21633 1347 21668 1381
rect 21668 1347 21702 1381
rect 21702 1347 21737 1381
rect 21737 1347 21771 1381
rect 21771 1347 21806 1381
rect 21806 1347 21840 1381
rect 21840 1347 21875 1381
rect 21875 1347 21909 1381
rect 21909 1347 21944 1381
rect 21944 1347 21978 1381
rect 21978 1347 22013 1381
rect 22013 1347 22047 1381
rect 22047 1347 22082 1381
rect 22082 1347 22116 1381
rect 22116 1347 22151 1381
rect 22151 1347 22185 1381
rect 22185 1347 22220 1381
rect 22220 1347 22254 1381
rect 22254 1347 22289 1381
rect 22289 1347 22323 1381
rect 22323 1347 22358 1381
rect 22358 1347 22392 1381
rect 22392 1347 22427 1381
rect 22427 1347 22461 1381
rect 22461 1347 22496 1381
rect 22496 1347 22530 1381
rect 22530 1347 22565 1381
rect 22565 1347 22599 1381
rect 22599 1347 22634 1381
rect 22634 1347 22668 1381
rect 22668 1347 22703 1381
rect 22703 1347 22737 1381
rect 22737 1347 22772 1381
rect 22772 1347 22806 1381
rect 22806 1347 22841 1381
rect 22841 1347 22875 1381
rect 22875 1347 22910 1381
rect 22910 1347 22944 1381
rect 22944 1347 22979 1381
rect 22979 1347 23013 1381
rect 23013 1347 23040 1381
rect 19563 1313 23040 1347
rect 19563 1279 19598 1313
rect 19598 1279 19632 1313
rect 19632 1279 19667 1313
rect 19667 1279 19701 1313
rect 19701 1279 19736 1313
rect 19736 1279 19770 1313
rect 19770 1279 19805 1313
rect 19805 1279 19839 1313
rect 19839 1279 19874 1313
rect 19874 1279 19908 1313
rect 19908 1279 19943 1313
rect 19943 1279 19977 1313
rect 19977 1279 20012 1313
rect 20012 1279 20046 1313
rect 20046 1279 20081 1313
rect 20081 1279 20115 1313
rect 20115 1279 20150 1313
rect 20150 1279 20184 1313
rect 20184 1279 20219 1313
rect 20219 1279 20253 1313
rect 20253 1279 20288 1313
rect 20288 1279 20322 1313
rect 20322 1279 20357 1313
rect 20357 1279 20391 1313
rect 20391 1279 20426 1313
rect 20426 1279 20460 1313
rect 20460 1279 20495 1313
rect 20495 1279 20529 1313
rect 20529 1279 20564 1313
rect 20564 1279 20598 1313
rect 20598 1279 20633 1313
rect 20633 1279 20667 1313
rect 20667 1279 20702 1313
rect 20702 1279 20736 1313
rect 20736 1279 20771 1313
rect 20771 1279 20805 1313
rect 20805 1279 20840 1313
rect 20840 1279 20874 1313
rect 20874 1279 20909 1313
rect 20909 1279 20943 1313
rect 20943 1279 20978 1313
rect 20978 1279 21012 1313
rect 21012 1279 21047 1313
rect 21047 1279 21081 1313
rect 21081 1279 21116 1313
rect 21116 1279 21150 1313
rect 21150 1279 21185 1313
rect 21185 1279 21219 1313
rect 21219 1279 21254 1313
rect 21254 1279 21288 1313
rect 21288 1279 21323 1313
rect 21323 1279 21357 1313
rect 21357 1279 21392 1313
rect 21392 1279 21426 1313
rect 21426 1279 21461 1313
rect 21461 1279 21495 1313
rect 21495 1279 21530 1313
rect 21530 1279 21564 1313
rect 21564 1279 21599 1313
rect 21599 1279 21633 1313
rect 21633 1279 21668 1313
rect 21668 1279 21702 1313
rect 21702 1279 21737 1313
rect 21737 1279 21771 1313
rect 21771 1279 21806 1313
rect 21806 1279 21840 1313
rect 21840 1279 21875 1313
rect 21875 1279 21909 1313
rect 21909 1279 21944 1313
rect 21944 1279 21978 1313
rect 21978 1279 22013 1313
rect 22013 1279 22047 1313
rect 22047 1279 22082 1313
rect 22082 1279 22116 1313
rect 22116 1279 22151 1313
rect 22151 1279 22185 1313
rect 22185 1279 22220 1313
rect 22220 1279 22254 1313
rect 22254 1279 22289 1313
rect 22289 1279 22323 1313
rect 22323 1279 22358 1313
rect 22358 1279 22392 1313
rect 22392 1279 22427 1313
rect 22427 1279 22461 1313
rect 22461 1279 22496 1313
rect 22496 1279 22530 1313
rect 22530 1279 22565 1313
rect 22565 1279 22599 1313
rect 22599 1279 22634 1313
rect 22634 1279 22668 1313
rect 22668 1279 22703 1313
rect 22703 1279 22737 1313
rect 22737 1279 22772 1313
rect 22772 1279 22806 1313
rect 22806 1279 22841 1313
rect 22841 1279 22875 1313
rect 22875 1279 22910 1313
rect 22910 1279 22944 1313
rect 22944 1279 22979 1313
rect 22979 1279 23013 1313
rect 23013 1279 23040 1313
rect 19563 1245 23040 1279
rect 19563 1211 19598 1245
rect 19598 1211 19632 1245
rect 19632 1211 19667 1245
rect 19667 1211 19701 1245
rect 19701 1211 19736 1245
rect 19736 1211 19770 1245
rect 19770 1211 19805 1245
rect 19805 1211 19839 1245
rect 19839 1211 19874 1245
rect 19874 1211 19908 1245
rect 19908 1211 19943 1245
rect 19943 1211 19977 1245
rect 19977 1211 20012 1245
rect 20012 1211 20046 1245
rect 20046 1211 20081 1245
rect 20081 1211 20115 1245
rect 20115 1211 20150 1245
rect 20150 1211 20184 1245
rect 20184 1211 20219 1245
rect 20219 1211 20253 1245
rect 20253 1211 20288 1245
rect 20288 1211 20322 1245
rect 20322 1211 20357 1245
rect 20357 1211 20391 1245
rect 20391 1211 20426 1245
rect 20426 1211 20460 1245
rect 20460 1211 20495 1245
rect 20495 1211 20529 1245
rect 20529 1211 20564 1245
rect 20564 1211 20598 1245
rect 20598 1211 20633 1245
rect 20633 1211 20667 1245
rect 20667 1211 20702 1245
rect 20702 1211 20736 1245
rect 20736 1211 20771 1245
rect 20771 1211 20805 1245
rect 20805 1211 20840 1245
rect 20840 1211 20874 1245
rect 20874 1211 20909 1245
rect 20909 1211 20943 1245
rect 20943 1211 20978 1245
rect 20978 1211 21012 1245
rect 21012 1211 21047 1245
rect 21047 1211 21081 1245
rect 21081 1211 21116 1245
rect 21116 1211 21150 1245
rect 21150 1211 21185 1245
rect 21185 1211 21219 1245
rect 21219 1211 21254 1245
rect 21254 1211 21288 1245
rect 21288 1211 21323 1245
rect 21323 1211 21357 1245
rect 21357 1211 21392 1245
rect 21392 1211 21426 1245
rect 21426 1211 21461 1245
rect 21461 1211 21495 1245
rect 21495 1211 21530 1245
rect 21530 1211 21564 1245
rect 21564 1211 21599 1245
rect 21599 1211 21633 1245
rect 21633 1211 21668 1245
rect 21668 1211 21702 1245
rect 21702 1211 21737 1245
rect 21737 1211 21771 1245
rect 21771 1211 21806 1245
rect 21806 1211 21840 1245
rect 21840 1211 21875 1245
rect 21875 1211 21909 1245
rect 21909 1211 21944 1245
rect 21944 1211 21978 1245
rect 21978 1211 22013 1245
rect 22013 1211 22047 1245
rect 22047 1211 22082 1245
rect 22082 1211 22116 1245
rect 22116 1211 22151 1245
rect 22151 1211 22185 1245
rect 22185 1211 22220 1245
rect 22220 1211 22254 1245
rect 22254 1211 22289 1245
rect 22289 1211 22323 1245
rect 22323 1211 22358 1245
rect 22358 1211 22392 1245
rect 22392 1211 22427 1245
rect 22427 1211 22461 1245
rect 22461 1211 22496 1245
rect 22496 1211 22530 1245
rect 22530 1211 22565 1245
rect 22565 1211 22599 1245
rect 22599 1211 22634 1245
rect 22634 1211 22668 1245
rect 22668 1211 22703 1245
rect 22703 1211 22737 1245
rect 22737 1211 22772 1245
rect 22772 1211 22806 1245
rect 22806 1211 22841 1245
rect 22841 1211 22875 1245
rect 22875 1211 22910 1245
rect 22910 1211 22944 1245
rect 22944 1211 22979 1245
rect 22979 1211 23013 1245
rect 23013 1211 23040 1245
rect 19563 1177 23040 1211
rect 19563 1172 19598 1177
rect 19598 1172 19632 1177
rect 19632 1172 19667 1177
rect 19667 1172 19701 1177
rect 19701 1172 19736 1177
rect 19736 1172 19770 1177
rect 19770 1172 19805 1177
rect 19805 1172 19839 1177
rect 19839 1172 19874 1177
rect 19874 1172 19908 1177
rect 19908 1172 19943 1177
rect 19943 1172 19977 1177
rect 19977 1172 20012 1177
rect 20012 1172 20046 1177
rect 20046 1172 20081 1177
rect 20081 1172 20115 1177
rect 20115 1172 20150 1177
rect 20150 1172 20184 1177
rect 20184 1172 20219 1177
rect 20219 1172 20253 1177
rect 20253 1172 20288 1177
rect 20288 1172 20322 1177
rect 20322 1172 20357 1177
rect 20357 1172 20391 1177
rect 20391 1172 20426 1177
rect 20426 1172 20460 1177
rect 20460 1172 20495 1177
rect 20495 1172 20529 1177
rect 20529 1172 20564 1177
rect 20564 1172 20598 1177
rect 20598 1172 20633 1177
rect 20633 1172 20667 1177
rect 20667 1172 20702 1177
rect 20702 1172 20736 1177
rect 20736 1172 20771 1177
rect 20771 1172 20805 1177
rect 20805 1172 20840 1177
rect 20840 1172 20874 1177
rect 20874 1172 20909 1177
rect 20909 1172 20943 1177
rect 20943 1172 20978 1177
rect 20978 1172 21012 1177
rect 21012 1172 21047 1177
rect 21047 1172 21081 1177
rect 21081 1172 21116 1177
rect 21116 1172 21150 1177
rect 21150 1172 21185 1177
rect 21185 1172 21219 1177
rect 21219 1172 21254 1177
rect 21254 1172 21288 1177
rect 21288 1172 21323 1177
rect 21323 1172 21357 1177
rect 21357 1172 21392 1177
rect 21392 1172 21426 1177
rect 21426 1172 21461 1177
rect 21461 1172 21495 1177
rect 21495 1172 21530 1177
rect 21530 1172 21564 1177
rect 21564 1172 21599 1177
rect 21599 1172 21633 1177
rect 21633 1172 21668 1177
rect 21668 1172 21702 1177
rect 21702 1172 21737 1177
rect 21737 1172 21771 1177
rect 21771 1172 21806 1177
rect 21806 1172 21840 1177
rect 21840 1172 21875 1177
rect 21875 1172 21909 1177
rect 21909 1172 21944 1177
rect 21944 1172 21978 1177
rect 21978 1172 22013 1177
rect 22013 1172 22047 1177
rect 22047 1172 22082 1177
rect 22082 1172 22116 1177
rect 22116 1172 22151 1177
rect 22151 1172 22185 1177
rect 22185 1172 22220 1177
rect 22220 1172 22254 1177
rect 22254 1172 22289 1177
rect 22289 1172 22323 1177
rect 22323 1172 22358 1177
rect 22358 1172 22392 1177
rect 22392 1172 22427 1177
rect 22427 1172 22461 1177
rect 22461 1172 22496 1177
rect 22496 1172 22530 1177
rect 22530 1172 22565 1177
rect 22565 1172 22599 1177
rect 22599 1172 22634 1177
rect 22634 1172 22668 1177
rect 22668 1172 22703 1177
rect 22703 1172 22737 1177
rect 22737 1172 22772 1177
rect 22772 1172 22806 1177
rect 22806 1172 22841 1177
rect 22841 1172 22875 1177
rect 22875 1172 22910 1177
rect 22910 1172 22944 1177
rect 22944 1172 22979 1177
rect 22979 1172 23013 1177
rect 23013 1172 23040 1177
rect 14487 1109 14521 1134
rect 14559 1112 14591 1134
rect 14591 1112 14593 1134
rect 23981 4800 24087 5532
rect 23981 4727 24015 4761
rect 24053 4727 24087 4761
rect 23981 4654 24015 4688
rect 24053 4654 24087 4688
rect 23981 4581 24015 4615
rect 24053 4581 24087 4615
rect 23981 4508 24015 4542
rect 24053 4508 24087 4542
rect 23981 4435 24015 4469
rect 24053 4435 24087 4469
rect 23981 4362 24015 4396
rect 24053 4362 24087 4396
rect 23981 4289 24015 4323
rect 24053 4289 24087 4323
rect 23981 4216 24015 4250
rect 24053 4216 24087 4250
rect 23981 4143 24015 4177
rect 24053 4143 24087 4177
rect 23981 4070 24015 4104
rect 24053 4070 24087 4104
rect 23981 3997 24015 4031
rect 24053 3997 24087 4031
rect 23981 3924 24015 3958
rect 24053 3924 24087 3958
rect 23981 3851 24015 3885
rect 24053 3851 24087 3885
rect 23981 3778 24015 3812
rect 24053 3778 24087 3812
rect 23981 3705 24015 3739
rect 24053 3705 24087 3739
rect 23981 3632 24015 3666
rect 24053 3632 24087 3666
rect 23981 3559 24015 3593
rect 24053 3559 24087 3593
rect 23981 3486 24015 3520
rect 24053 3486 24087 3520
rect 23981 3413 24015 3447
rect 24053 3413 24087 3447
rect 23981 3340 24015 3374
rect 24053 3340 24087 3374
rect 23981 3267 24015 3301
rect 24053 3267 24087 3301
rect 23981 3194 24015 3228
rect 24053 3194 24087 3228
rect 23981 3121 24015 3155
rect 24053 3121 24087 3155
rect 23981 3048 24015 3082
rect 24053 3048 24087 3082
rect 23981 2975 24015 3009
rect 24053 2975 24087 3009
rect 23981 2902 24015 2936
rect 24053 2902 24087 2936
rect 23981 2829 24015 2863
rect 24053 2829 24087 2863
rect 23981 2756 24015 2790
rect 24053 2756 24087 2790
rect 23981 2683 24015 2717
rect 24053 2683 24087 2717
rect 23981 2610 24015 2644
rect 24053 2610 24087 2644
rect 23981 2537 24015 2571
rect 24053 2537 24087 2571
rect 23981 2464 24015 2498
rect 24053 2464 24087 2498
rect 23981 2391 24015 2425
rect 24053 2391 24087 2425
rect 23981 2318 24015 2352
rect 24053 2318 24087 2352
rect 23981 2245 24015 2279
rect 24053 2245 24087 2279
rect 23981 2172 24015 2206
rect 24053 2172 24087 2206
rect 23981 2099 24015 2133
rect 24053 2099 24087 2133
rect 23981 2026 24015 2060
rect 24053 2026 24087 2060
rect 23981 1953 24015 1987
rect 24053 1953 24087 1987
rect 23981 1880 24015 1914
rect 24053 1880 24087 1914
rect 23981 1807 24015 1841
rect 24053 1807 24087 1841
rect 23981 1734 24015 1768
rect 24053 1734 24087 1768
rect 14487 1100 14489 1109
rect 14489 1100 14521 1109
rect 800 1044 834 1078
rect 14559 1100 14593 1112
rect 728 1040 730 1043
rect 730 1040 762 1043
rect 728 1009 762 1040
rect 14559 1042 14591 1053
rect 14591 1042 14593 1053
rect 14559 1019 14593 1042
rect 800 1003 834 1005
rect 873 1003 901 1005
rect 901 1003 907 1005
rect 946 1003 970 1005
rect 970 1003 980 1005
rect 1019 1003 1039 1005
rect 1039 1003 1053 1005
rect 1092 1003 1108 1005
rect 1108 1003 1126 1005
rect 1165 1003 1177 1005
rect 1177 1003 1199 1005
rect 1238 1003 1246 1005
rect 1246 1003 1272 1005
rect 1311 1003 1315 1005
rect 1315 1003 1349 1005
rect 1349 1003 1384 1005
rect 1384 1003 1418 1005
rect 1418 1003 1453 1005
rect 1453 1003 1487 1005
rect 1487 1003 1522 1005
rect 1522 1003 1556 1005
rect 1556 1003 1591 1005
rect 1591 1003 1625 1005
rect 1625 1003 1660 1005
rect 1660 1003 1694 1005
rect 1694 1003 1729 1005
rect 1729 1003 1763 1005
rect 1763 1003 1798 1005
rect 1798 1003 1832 1005
rect 1832 1003 1867 1005
rect 1867 1003 1901 1005
rect 1901 1003 1936 1005
rect 1936 1003 1970 1005
rect 1970 1003 2005 1005
rect 2005 1003 2039 1005
rect 2039 1003 2074 1005
rect 2074 1003 2108 1005
rect 2108 1003 2143 1005
rect 2143 1003 2177 1005
rect 2177 1003 2212 1005
rect 2212 1003 2246 1005
rect 2246 1003 2281 1005
rect 2281 1003 2315 1005
rect 2315 1003 2350 1005
rect 2350 1003 2384 1005
rect 2384 1003 2419 1005
rect 800 971 834 1003
rect 873 971 907 1003
rect 946 971 980 1003
rect 1019 971 1053 1003
rect 1092 971 1126 1003
rect 1165 971 1199 1003
rect 1238 971 1272 1003
rect 1311 969 2419 1003
rect 2419 969 14483 1005
rect 14487 971 14489 1005
rect 14489 971 14521 1005
rect 1311 935 1316 969
rect 1316 935 1350 969
rect 1350 935 1385 969
rect 1385 935 1419 969
rect 1419 935 1454 969
rect 1454 935 1488 969
rect 1488 935 1523 969
rect 1523 935 1557 969
rect 1557 935 1592 969
rect 1592 935 1626 969
rect 1626 935 1661 969
rect 1661 935 1695 969
rect 1695 935 1730 969
rect 1730 935 1764 969
rect 1764 935 1799 969
rect 1799 935 1833 969
rect 1833 935 1868 969
rect 1868 935 1902 969
rect 1902 935 1937 969
rect 1937 935 1971 969
rect 1971 935 2006 969
rect 2006 935 2040 969
rect 2040 935 2075 969
rect 2075 935 2109 969
rect 2109 935 2144 969
rect 2144 935 2178 969
rect 2178 935 2213 969
rect 2213 935 2247 969
rect 2247 935 2282 969
rect 2282 935 2316 969
rect 2316 935 2351 969
rect 766 901 800 933
rect 839 901 873 933
rect 912 901 946 933
rect 985 901 1019 933
rect 1057 901 1091 933
rect 1129 901 1163 933
rect 1201 901 1235 933
rect 1273 901 1307 933
rect 1311 901 2351 935
rect 2351 901 14483 969
rect 14559 937 14593 971
rect 766 899 799 901
rect 799 899 800 901
rect 839 899 868 901
rect 868 899 873 901
rect 912 899 937 901
rect 937 899 946 901
rect 985 899 1006 901
rect 1006 899 1019 901
rect 1057 899 1075 901
rect 1075 899 1091 901
rect 1129 899 1144 901
rect 1144 899 1163 901
rect 1201 899 1213 901
rect 1213 899 1235 901
rect 1273 899 1282 901
rect 1282 899 1307 901
rect 1311 899 1316 901
rect 1316 899 1351 901
rect 1351 899 1385 901
rect 1385 899 1420 901
rect 1420 899 1454 901
rect 1454 899 1489 901
rect 1489 899 1523 901
rect 1523 899 1558 901
rect 1558 899 1592 901
rect 1592 899 1627 901
rect 1627 899 1661 901
rect 1661 899 1696 901
rect 1696 899 1730 901
rect 1730 899 1765 901
rect 1765 899 1799 901
rect 1799 899 1834 901
rect 1834 899 1868 901
rect 1868 899 1903 901
rect 1903 899 1937 901
rect 1937 899 1972 901
rect 1972 899 2006 901
rect 2006 899 2041 901
rect 2041 899 2075 901
rect 2075 899 2110 901
rect 2110 899 2144 901
rect 2144 899 2179 901
rect 2179 899 2213 901
rect 2213 899 2248 901
rect 2248 899 2282 901
rect 2282 899 2317 901
rect 2317 899 14483 901
rect 20551 942 20558 944
rect 20558 942 20585 944
rect 20625 942 20627 944
rect 20627 942 20659 944
rect 20699 942 20730 944
rect 20730 942 20733 944
rect 20773 942 20799 944
rect 20799 942 20807 944
rect 20847 942 20868 944
rect 20868 942 20881 944
rect 20921 942 20937 944
rect 20937 942 20955 944
rect 20995 942 21006 944
rect 21006 942 21029 944
rect 21069 942 21075 944
rect 21075 942 21103 944
rect 21143 942 21144 944
rect 21144 942 21177 944
rect 21217 942 21248 944
rect 21248 942 21251 944
rect 21291 942 21317 944
rect 21317 942 21325 944
rect 21365 942 21386 944
rect 21386 942 21399 944
rect 21439 942 21455 944
rect 21455 942 21473 944
rect 21513 942 21524 944
rect 21524 942 21547 944
rect 21587 942 21593 944
rect 21593 942 21621 944
rect 21661 942 21662 944
rect 21662 942 21695 944
rect 21735 942 21765 944
rect 21765 942 21769 944
rect 21809 942 21834 944
rect 21834 942 21843 944
rect 21883 942 21903 944
rect 21903 942 21917 944
rect 21957 942 21972 944
rect 21972 942 21991 944
rect 22031 942 22041 944
rect 22041 942 22065 944
rect 22105 942 22110 944
rect 22110 942 22139 944
rect 20551 910 20585 942
rect 20625 910 20659 942
rect 20699 910 20733 942
rect 20773 910 20807 942
rect 20847 910 20881 942
rect 20921 910 20955 942
rect 20995 910 21029 942
rect 21069 910 21103 942
rect 21143 910 21177 942
rect 21217 910 21251 942
rect 21291 910 21325 942
rect 21365 910 21399 942
rect 21439 910 21473 942
rect 21513 910 21547 942
rect 21587 910 21621 942
rect 21661 910 21695 942
rect 21735 910 21769 942
rect 21809 910 21843 942
rect 21883 910 21917 942
rect 21957 910 21991 942
rect 22031 910 22065 942
rect 22105 910 22139 942
rect 22179 910 22213 944
rect 22253 942 22283 944
rect 22283 942 22287 944
rect 22327 942 22352 944
rect 22352 942 22361 944
rect 22401 942 22421 944
rect 22421 942 22435 944
rect 22475 942 22490 944
rect 22490 942 22509 944
rect 22549 942 22559 944
rect 22559 942 22583 944
rect 22622 942 22628 944
rect 22628 942 22656 944
rect 22695 942 22697 944
rect 22697 942 22729 944
rect 22768 942 22800 944
rect 22800 942 22802 944
rect 22841 942 22869 944
rect 22869 942 22875 944
rect 22914 942 22938 944
rect 22938 942 22948 944
rect 22253 910 22287 942
rect 22327 910 22361 942
rect 22401 910 22435 942
rect 22475 910 22509 942
rect 22549 910 22583 942
rect 22622 910 22656 942
rect 22695 910 22729 942
rect 22768 910 22802 942
rect 22841 910 22875 942
rect 22914 910 22948 942
rect 22987 910 23021 944
rect 23060 910 23094 944
rect 23133 910 23167 944
rect 23206 910 23240 944
rect 23279 910 23313 944
rect 23352 910 23386 944
rect 23425 910 23459 944
rect 23498 910 23532 944
rect 23571 910 23605 944
rect 23644 910 23678 944
rect 23717 910 23751 944
rect 310 822 344 855
rect 382 822 416 855
rect 310 821 312 822
rect 312 821 344 822
rect 382 821 414 822
rect 414 821 416 822
rect 20551 840 20585 872
rect 20625 840 20659 872
rect 20699 840 20733 872
rect 20773 840 20807 872
rect 20847 840 20881 872
rect 20921 840 20955 872
rect 20995 840 21029 872
rect 21069 840 21103 872
rect 21143 840 21177 872
rect 21217 840 21251 872
rect 21291 840 21325 872
rect 21365 840 21399 872
rect 21439 840 21473 872
rect 21513 840 21547 872
rect 21587 840 21621 872
rect 21661 840 21695 872
rect 21735 840 21769 872
rect 21809 840 21843 872
rect 21883 840 21917 872
rect 21957 840 21991 872
rect 22031 840 22065 872
rect 22105 840 22139 872
rect 20551 838 20558 840
rect 20558 838 20585 840
rect 20625 838 20627 840
rect 20627 838 20659 840
rect 20699 838 20730 840
rect 20730 838 20733 840
rect 20773 838 20799 840
rect 20799 838 20807 840
rect 20847 838 20868 840
rect 20868 838 20881 840
rect 20921 838 20937 840
rect 20937 838 20955 840
rect 20995 838 21006 840
rect 21006 838 21029 840
rect 21069 838 21075 840
rect 21075 838 21103 840
rect 21143 838 21144 840
rect 21144 838 21177 840
rect 21217 838 21248 840
rect 21248 838 21251 840
rect 21291 838 21317 840
rect 21317 838 21325 840
rect 21365 838 21386 840
rect 21386 838 21399 840
rect 21439 838 21455 840
rect 21455 838 21473 840
rect 21513 838 21524 840
rect 21524 838 21547 840
rect 21587 838 21593 840
rect 21593 838 21621 840
rect 21661 838 21662 840
rect 21662 838 21695 840
rect 21735 838 21765 840
rect 21765 838 21769 840
rect 21809 838 21834 840
rect 21834 838 21843 840
rect 21883 838 21903 840
rect 21903 838 21917 840
rect 21957 838 21972 840
rect 21972 838 21991 840
rect 22031 838 22041 840
rect 22041 838 22065 840
rect 22105 838 22110 840
rect 22110 838 22139 840
rect 22179 838 22213 872
rect 22253 840 22287 872
rect 22327 840 22361 872
rect 22401 840 22435 872
rect 22475 840 22509 872
rect 22549 840 22583 872
rect 22622 840 22656 872
rect 22695 840 22729 872
rect 22768 840 22802 872
rect 22841 840 22875 872
rect 22914 840 22948 872
rect 22253 838 22283 840
rect 22283 838 22287 840
rect 22327 838 22352 840
rect 22352 838 22361 840
rect 22401 838 22421 840
rect 22421 838 22435 840
rect 22475 838 22490 840
rect 22490 838 22509 840
rect 22549 838 22559 840
rect 22559 838 22583 840
rect 22622 838 22628 840
rect 22628 838 22656 840
rect 22695 838 22697 840
rect 22697 838 22729 840
rect 22768 838 22800 840
rect 22800 838 22802 840
rect 22841 838 22869 840
rect 22869 838 22875 840
rect 22914 838 22938 840
rect 22938 838 22948 840
rect 22987 838 23021 872
rect 23060 838 23094 872
rect 23133 838 23167 872
rect 23206 838 23240 872
rect 23279 838 23313 872
rect 23352 838 23386 872
rect 23425 838 23459 872
rect 23498 838 23532 872
rect 23571 838 23605 872
rect 23644 838 23678 872
rect 23717 838 23751 872
rect 310 753 344 782
rect 382 753 416 782
rect 310 748 312 753
rect 312 748 344 753
rect 382 748 414 753
rect 414 748 416 753
rect 310 684 344 709
rect 382 684 416 709
rect 310 675 312 684
rect 312 675 344 684
rect 382 675 414 684
rect 414 675 416 684
rect 310 615 344 636
rect 382 615 416 636
rect 310 602 312 615
rect 312 602 344 615
rect 382 602 414 615
rect 414 602 416 615
rect 310 546 344 563
rect 382 546 416 563
rect 310 529 312 546
rect 312 529 344 546
rect 382 529 414 546
rect 414 529 416 546
rect 310 477 344 490
rect 382 477 416 490
rect 310 456 312 477
rect 312 456 344 477
rect 382 456 414 477
rect 414 456 416 477
rect 310 408 344 417
rect 382 408 416 417
rect 310 383 312 408
rect 312 383 344 408
rect 382 383 414 408
rect 414 383 416 408
rect 310 339 344 344
rect 382 339 416 344
rect 310 310 312 339
rect 312 310 344 339
rect 382 310 414 339
rect 414 310 416 339
rect 310 270 344 271
rect 382 270 416 271
rect 310 237 312 270
rect 312 237 344 270
rect 382 237 414 270
rect 414 237 416 270
rect 310 167 312 198
rect 312 167 344 198
rect 382 167 414 198
rect 414 167 416 198
rect 310 164 344 167
rect 382 164 416 167
rect 21197 -1923 21231 -1889
rect 21269 -1923 21303 -1889
rect 21341 -1923 21375 -1889
rect 21413 -1923 21447 -1889
rect 21485 -1923 21519 -1889
<< metal1 >>
rect 23743 13310 23795 13316
rect 23743 13246 23795 13258
rect 23743 13188 23795 13194
rect 24229 10991 24281 10997
rect 24229 10927 24281 10939
rect 24735 10905 24741 10957
rect 24793 10905 24805 10957
rect 24857 10905 27440 10957
rect 27492 10905 27504 10957
rect 27556 10905 27562 10957
tri 24195 10123 24229 10157 se
rect 24229 10124 24281 10875
rect 25294 10812 25300 10864
rect 25352 10812 25364 10864
rect 25416 10812 25672 10864
rect 25724 10812 25736 10864
rect 25788 10812 25794 10864
rect 25993 10820 25999 10872
rect 26051 10820 26091 10872
rect 26143 10820 26183 10872
rect 26235 10820 26275 10872
rect 26327 10820 26367 10872
rect 26419 10820 26425 10872
rect 25256 10504 25262 10556
rect 25314 10504 25326 10556
rect 25378 10504 25384 10556
rect 25705 10504 25711 10556
rect 25763 10504 25775 10556
rect 25827 10504 27505 10556
rect 27557 10504 27569 10556
rect 27621 10504 27627 10556
rect 25762 10444 25814 10450
rect 25762 10379 25814 10392
rect 25762 10314 25814 10327
rect 25762 10248 25814 10262
rect 25762 10190 25814 10196
tri 24281 10124 24314 10157 sw
rect 24229 10123 24314 10124
tri 24314 10123 24315 10124 sw
tri 25264 10123 25265 10124 se
rect 25265 10123 25408 10124
rect 24189 10071 24195 10123
rect 24247 10071 24259 10123
rect 24311 10071 24317 10123
tri 25213 10072 25264 10123 se
rect 25264 10072 25408 10123
rect 25460 10072 25472 10124
rect 25524 10072 28069 10124
rect 28121 10072 28133 10124
rect 28185 10072 28191 10124
tri 25212 10071 25213 10072 se
rect 25213 10071 25265 10072
tri 25179 10038 25212 10071 se
rect 25212 10038 25265 10071
tri 25265 10038 25299 10072 nw
tri 25128 9987 25179 10038 se
rect 25179 9987 25214 10038
tri 25214 9987 25265 10038 nw
rect 25128 9974 25201 9987
tri 25201 9974 25214 9987 nw
rect 16993 9761 19340 9879
tri 16993 9759 16995 9761 ne
rect 16995 9759 19338 9761
tri 19338 9759 19340 9761 nw
rect 20696 9875 21415 9876
rect 20696 9823 20702 9875
rect 20754 9823 20768 9875
rect 20820 9823 20834 9875
rect 20886 9823 20900 9875
rect 20952 9823 20966 9875
rect 21018 9823 21032 9875
rect 21084 9823 21097 9875
rect 21149 9823 21162 9875
rect 21214 9823 21227 9875
rect 21279 9823 21292 9875
rect 21344 9823 21357 9875
rect 21409 9823 21415 9875
rect 20696 9811 21415 9823
rect 20696 9759 20702 9811
rect 20754 9759 20768 9811
rect 20820 9759 20834 9811
rect 20886 9759 20900 9811
rect 20952 9759 20966 9811
rect 21018 9759 21032 9811
rect 21084 9759 21097 9811
rect 21149 9759 21162 9811
rect 21214 9759 21227 9811
rect 21279 9759 21292 9811
rect 21344 9759 21357 9811
rect 21409 9759 21415 9811
tri 16995 9736 17018 9759 ne
rect 17018 9687 19315 9759
tri 19315 9736 19338 9759 nw
rect 20696 9758 21415 9759
rect 17018 9635 17024 9687
rect 17076 9635 17090 9687
rect 17142 9635 17156 9687
rect 17208 9635 17222 9687
rect 17274 9635 17288 9687
rect 17340 9635 17354 9687
rect 17406 9635 17420 9687
rect 17472 9635 17486 9687
rect 17538 9635 17552 9687
rect 17604 9635 17618 9687
rect 17670 9635 17684 9687
rect 17736 9635 17750 9687
rect 17802 9635 17816 9687
rect 17868 9635 17882 9687
rect 17934 9635 17948 9687
rect 18000 9635 18014 9687
rect 18066 9635 18080 9687
rect 18132 9635 18146 9687
rect 18198 9635 18212 9687
rect 18264 9635 18278 9687
rect 18330 9635 18344 9687
rect 18396 9635 18410 9687
rect 18462 9635 18476 9687
rect 18528 9635 18542 9687
rect 18594 9635 18607 9687
rect 18659 9635 18672 9687
rect 18724 9635 18737 9687
rect 18789 9635 18802 9687
rect 18854 9635 18867 9687
rect 18919 9635 18932 9687
rect 18984 9635 18997 9687
rect 19049 9635 19062 9687
rect 19114 9635 19127 9687
rect 19179 9635 19192 9687
rect 19244 9635 19257 9687
rect 19309 9635 19315 9687
rect 17018 9623 19315 9635
rect 17018 9571 17024 9623
rect 17076 9571 17090 9623
rect 17142 9571 17156 9623
rect 17208 9571 17222 9623
rect 17274 9571 17288 9623
rect 17340 9571 17354 9623
rect 17406 9571 17420 9623
rect 17472 9571 17486 9623
rect 17538 9571 17552 9623
rect 17604 9571 17618 9623
rect 17670 9571 17684 9623
rect 17736 9571 17750 9623
rect 17802 9571 17816 9623
rect 17868 9571 17882 9623
rect 17934 9571 17948 9623
rect 18000 9571 18014 9623
rect 18066 9571 18080 9623
rect 18132 9571 18146 9623
rect 18198 9571 18212 9623
rect 18264 9571 18278 9623
rect 18330 9571 18344 9623
rect 18396 9571 18410 9623
rect 18462 9571 18476 9623
rect 18528 9571 18542 9623
rect 18594 9571 18607 9623
rect 18659 9571 18672 9623
rect 18724 9571 18737 9623
rect 18789 9571 18802 9623
rect 18854 9571 18867 9623
rect 18919 9571 18932 9623
rect 18984 9571 18997 9623
rect 19049 9571 19062 9623
rect 19114 9571 19127 9623
rect 19179 9571 19192 9623
rect 19244 9571 19257 9623
rect 19309 9571 19315 9623
tri 24273 9159 24396 9282 se
rect 24396 9159 24514 9428
rect 25128 9353 25190 9974
tri 25190 9963 25201 9974 nw
rect 25505 9922 25511 9974
rect 25563 9922 25575 9974
rect 25627 9922 27664 9974
rect 27716 9922 27728 9974
rect 27780 9922 27786 9974
tri 25479 9779 25480 9780 se
rect 25480 9779 27312 9780
rect 25241 9727 25247 9779
rect 25299 9727 25311 9779
rect 25363 9728 27312 9779
rect 27364 9728 27376 9780
rect 27428 9728 27434 9780
rect 25363 9727 25501 9728
tri 25501 9727 25502 9728 nw
rect 27341 9546 27395 9552
rect 27341 9494 27342 9546
rect 27394 9494 27395 9546
rect 27341 9482 27395 9494
rect 27341 9430 27342 9482
rect 27394 9476 27395 9482
tri 27395 9476 27471 9552 sw
rect 27394 9430 27922 9476
rect 27341 9424 27922 9430
rect 27974 9424 27986 9476
rect 28038 9424 28044 9476
tri 24265 9151 24273 9159 se
rect 24273 9151 24514 9159
tri 24514 9151 24522 9159 sw
tri 22740 9132 22759 9151 sw
tri 24246 9132 24265 9151 se
rect 24265 9132 24522 9151
tri 24522 9132 24541 9151 sw
rect 22740 9069 22759 9132
tri 22759 9069 22822 9132 sw
rect 23775 9126 24541 9132
rect 17018 9039 17029 9069
rect 17023 9017 17029 9039
rect 17081 9017 17095 9069
rect 17147 9017 17161 9069
rect 17213 9017 17227 9069
rect 17279 9017 17293 9069
rect 17345 9017 17359 9069
rect 17411 9017 17425 9069
rect 17477 9017 17491 9069
rect 17543 9017 17557 9069
rect 17609 9017 17623 9069
rect 17675 9017 17689 9069
rect 17741 9017 17755 9069
rect 17807 9017 17821 9069
rect 17873 9017 17887 9069
rect 17939 9017 17953 9069
rect 18005 9017 18019 9069
rect 18071 9017 18085 9069
rect 18137 9017 18151 9069
rect 18203 9017 18217 9069
rect 18269 9017 18282 9069
rect 18334 9017 18347 9069
rect 18399 9017 18412 9069
rect 18464 9017 18477 9069
rect 18529 9017 18542 9069
rect 18594 9017 18607 9069
rect 18659 9017 18672 9069
rect 18724 9017 18737 9069
rect 18789 9017 18802 9069
rect 18854 9017 18867 9069
rect 18919 9017 18932 9069
rect 18984 9017 18997 9069
rect 19049 9017 19062 9069
rect 19114 9017 19127 9069
rect 19179 9017 19192 9069
rect 19244 9017 19257 9069
rect 19309 9017 19315 9069
rect 22740 9064 22822 9069
tri 22822 9064 22827 9069 sw
tri 19315 9039 19340 9064 sw
rect 22740 9039 22827 9064
tri 22827 9039 22852 9064 sw
rect 17023 9005 19315 9017
rect 22740 9009 22852 9039
tri 22852 9009 22882 9039 sw
rect 17023 8953 17029 9005
rect 17081 8953 17095 9005
rect 17147 8953 17161 9005
rect 17213 8953 17227 9005
rect 17279 8953 17293 9005
rect 17345 8953 17359 9005
rect 17411 8953 17425 9005
rect 17477 8953 17491 9005
rect 17543 8953 17557 9005
rect 17609 8953 17623 9005
rect 17675 8953 17689 9005
rect 17741 8953 17755 9005
rect 17807 8953 17821 9005
rect 17873 8953 17887 9005
rect 17939 8953 17953 9005
rect 18005 8953 18019 9005
rect 18071 8953 18085 9005
rect 18137 8953 18151 9005
rect 18203 8953 18217 9005
rect 18269 8953 18282 9005
rect 18334 8953 18347 9005
rect 18399 8953 18412 9005
rect 18464 8953 18477 9005
rect 18529 8953 18542 9005
rect 18594 8953 18607 9005
rect 18659 8953 18672 9005
rect 18724 8953 18737 9005
rect 18789 8953 18802 9005
rect 18854 8953 18867 9005
rect 18919 8953 18932 9005
rect 18984 8953 18997 9005
rect 19049 8953 19062 9005
rect 19114 8953 19127 9005
rect 19179 8953 19192 9005
rect 19244 8953 19257 9005
rect 19309 8953 19315 9005
rect 20696 8953 20702 9005
rect 20754 8953 20768 9005
rect 20820 8953 20834 9005
rect 20886 8953 20900 9005
rect 20952 8953 20966 9005
rect 21018 8953 21032 9005
rect 21084 8953 21097 9005
rect 21149 8953 21162 9005
rect 21214 8953 21227 9005
rect 21279 8953 21292 9005
rect 21344 8953 21357 9005
rect 21409 8953 21415 9005
rect 20696 8941 21415 8953
rect 20696 8889 20702 8941
rect 20754 8889 20768 8941
rect 20820 8889 20834 8941
rect 20886 8889 20900 8941
rect 20952 8889 20966 8941
rect 21018 8889 21032 8941
rect 21084 8889 21097 8941
rect 21149 8889 21162 8941
rect 21214 8889 21227 8941
rect 21279 8889 21292 8941
rect 21344 8889 21357 8941
rect 21409 8889 21415 8941
rect 20696 8877 21415 8889
rect 20696 8825 20702 8877
rect 20754 8825 20768 8877
rect 20820 8825 20834 8877
rect 20886 8825 20900 8877
rect 20952 8825 20966 8877
rect 21018 8825 21032 8877
rect 21084 8825 21097 8877
rect 21149 8825 21162 8877
rect 21214 8825 21227 8877
rect 21279 8825 21292 8877
rect 21344 8825 21357 8877
rect 21409 8825 21415 8877
rect 17023 8762 17029 8814
rect 17081 8762 17095 8814
rect 17147 8762 17161 8814
rect 17213 8762 17227 8814
rect 17279 8762 17293 8814
rect 17345 8762 17359 8814
rect 17411 8762 17425 8814
rect 17477 8762 17491 8814
rect 17543 8762 17557 8814
rect 17609 8762 17623 8814
rect 17675 8762 17689 8814
rect 17741 8762 17755 8814
rect 17807 8762 17821 8814
rect 17873 8762 17887 8814
rect 17939 8762 17953 8814
rect 18005 8762 18019 8814
rect 18071 8762 18085 8814
rect 18137 8762 18151 8814
rect 18203 8762 18217 8814
rect 18269 8762 18282 8814
rect 18334 8762 18347 8814
rect 18399 8762 18412 8814
rect 18464 8762 18477 8814
rect 18529 8762 18542 8814
rect 18594 8762 18607 8814
rect 18659 8762 18672 8814
rect 18724 8762 18737 8814
rect 18789 8762 18802 8814
rect 18854 8762 18867 8814
rect 18919 8762 18932 8814
rect 18984 8762 18997 8814
rect 19049 8762 19062 8814
rect 19114 8762 19127 8814
rect 19179 8762 19192 8814
rect 19244 8762 19257 8814
rect 19309 8762 19315 8814
rect 17023 8750 19315 8762
rect 17023 8698 17029 8750
rect 17081 8698 17095 8750
rect 17147 8698 17161 8750
rect 17213 8698 17227 8750
rect 17279 8698 17293 8750
rect 17345 8698 17359 8750
rect 17411 8698 17425 8750
rect 17477 8698 17491 8750
rect 17543 8698 17557 8750
rect 17609 8698 17623 8750
rect 17675 8698 17689 8750
rect 17741 8698 17755 8750
rect 17807 8698 17821 8750
rect 17873 8698 17887 8750
rect 17939 8698 17953 8750
rect 18005 8698 18019 8750
rect 18071 8698 18085 8750
rect 18137 8698 18151 8750
rect 18203 8698 18217 8750
rect 18269 8698 18282 8750
rect 18334 8698 18347 8750
rect 18399 8698 18412 8750
rect 18464 8698 18477 8750
rect 18529 8698 18542 8750
rect 18594 8698 18607 8750
rect 18659 8698 18672 8750
rect 18724 8698 18737 8750
rect 18789 8698 18802 8750
rect 18854 8698 18867 8750
rect 18919 8698 18932 8750
rect 18984 8698 18997 8750
rect 19049 8698 19062 8750
rect 19114 8698 19127 8750
rect 19179 8698 19192 8750
rect 19244 8698 19257 8750
rect 19309 8698 19315 8750
rect 17023 8686 19315 8698
rect 17023 8634 17029 8686
rect 17081 8634 17095 8686
rect 17147 8634 17161 8686
rect 17213 8634 17227 8686
rect 17279 8634 17293 8686
rect 17345 8634 17359 8686
rect 17411 8634 17425 8686
rect 17477 8634 17491 8686
rect 17543 8634 17557 8686
rect 17609 8634 17623 8686
rect 17675 8634 17689 8686
rect 17741 8634 17755 8686
rect 17807 8634 17821 8686
rect 17873 8634 17887 8686
rect 17939 8634 17953 8686
rect 18005 8634 18019 8686
rect 18071 8634 18085 8686
rect 18137 8634 18151 8686
rect 18203 8634 18217 8686
rect 18269 8634 18282 8686
rect 18334 8634 18347 8686
rect 18399 8634 18412 8686
rect 18464 8634 18477 8686
rect 18529 8634 18542 8686
rect 18594 8634 18607 8686
rect 18659 8634 18672 8686
rect 18724 8634 18737 8686
rect 18789 8634 18802 8686
rect 18854 8634 18867 8686
rect 18919 8634 18932 8686
rect 18984 8634 18997 8686
rect 19049 8634 19062 8686
rect 19114 8634 19127 8686
rect 19179 8634 19192 8686
rect 19244 8634 19257 8686
rect 19309 8634 19315 8686
rect 20696 8813 21415 8825
rect 20696 8761 20702 8813
rect 20754 8761 20768 8813
rect 20820 8761 20834 8813
rect 20886 8761 20900 8813
rect 20952 8761 20966 8813
rect 21018 8761 21032 8813
rect 21084 8761 21097 8813
rect 21149 8761 21162 8813
rect 21214 8761 21227 8813
rect 21279 8761 21292 8813
rect 21344 8761 21357 8813
rect 21409 8761 21415 8813
rect 20696 8749 21415 8761
rect 20696 8697 20702 8749
rect 20754 8697 20768 8749
rect 20820 8697 20834 8749
rect 20886 8697 20900 8749
rect 20952 8697 20966 8749
rect 21018 8697 21032 8749
rect 21084 8697 21097 8749
rect 21149 8697 21162 8749
rect 21214 8697 21227 8749
rect 21279 8697 21292 8749
rect 21344 8697 21357 8749
rect 21409 8697 21415 8749
rect 20696 8685 21415 8697
rect 20696 8633 20702 8685
rect 20754 8633 20768 8685
rect 20820 8633 20834 8685
rect 20886 8633 20900 8685
rect 20952 8633 20966 8685
rect 21018 8633 21032 8685
rect 21084 8633 21097 8685
rect 21149 8633 21162 8685
rect 21214 8633 21227 8685
rect 21279 8633 21292 8685
rect 21344 8633 21357 8685
rect 21409 8633 21415 8685
rect 22716 8997 23486 9009
rect 22716 8603 22798 8997
rect 23480 8603 23486 8997
rect 20503 8523 20509 8575
rect 20561 8523 20573 8575
rect 20625 8523 20631 8575
rect 22716 8564 23486 8603
rect 22716 8530 22798 8564
rect 22832 8530 22870 8564
rect 22904 8530 22942 8564
rect 22976 8530 23014 8564
rect 23048 8530 23086 8564
rect 23120 8530 23158 8564
rect 23192 8530 23230 8564
rect 23264 8530 23302 8564
rect 23336 8530 23374 8564
rect 23408 8530 23446 8564
rect 23480 8530 23486 8564
rect 17023 8443 17029 8495
rect 17081 8443 17095 8495
rect 17147 8443 17161 8495
rect 17213 8443 17227 8495
rect 17279 8443 17293 8495
rect 17345 8443 17359 8495
rect 17411 8443 17425 8495
rect 17477 8443 17491 8495
rect 17543 8443 17557 8495
rect 17609 8443 17623 8495
rect 17675 8443 17689 8495
rect 17741 8443 17755 8495
rect 17807 8443 17821 8495
rect 17873 8443 17887 8495
rect 17939 8443 17953 8495
rect 18005 8443 18019 8495
rect 18071 8443 18085 8495
rect 18137 8443 18151 8495
rect 18203 8443 18217 8495
rect 18269 8443 18282 8495
rect 18334 8443 18347 8495
rect 18399 8443 18412 8495
rect 18464 8443 18477 8495
rect 18529 8443 18542 8495
rect 18594 8443 18607 8495
rect 18659 8443 18672 8495
rect 18724 8443 18737 8495
rect 18789 8443 18802 8495
rect 18854 8443 18867 8495
rect 18919 8443 18932 8495
rect 18984 8443 18997 8495
rect 19049 8443 19062 8495
rect 19114 8443 19127 8495
rect 19179 8443 19192 8495
rect 19244 8443 19257 8495
rect 19309 8443 19315 8495
rect 17023 8431 19315 8443
rect 17023 8379 17029 8431
rect 17081 8379 17095 8431
rect 17147 8379 17161 8431
rect 17213 8379 17227 8431
rect 17279 8379 17293 8431
rect 17345 8379 17359 8431
rect 17411 8379 17425 8431
rect 17477 8379 17491 8431
rect 17543 8379 17557 8431
rect 17609 8379 17623 8431
rect 17675 8379 17689 8431
rect 17741 8379 17755 8431
rect 17807 8379 17821 8431
rect 17873 8379 17887 8431
rect 17939 8379 17953 8431
rect 18005 8379 18019 8431
rect 18071 8379 18085 8431
rect 18137 8379 18151 8431
rect 18203 8379 18217 8431
rect 18269 8379 18282 8431
rect 18334 8379 18347 8431
rect 18399 8379 18412 8431
rect 18464 8379 18477 8431
rect 18529 8379 18542 8431
rect 18594 8379 18607 8431
rect 18659 8379 18672 8431
rect 18724 8379 18737 8431
rect 18789 8379 18802 8431
rect 18854 8379 18867 8431
rect 18919 8379 18932 8431
rect 18984 8379 18997 8431
rect 19049 8379 19062 8431
rect 19114 8379 19127 8431
rect 19179 8379 19192 8431
rect 19244 8379 19257 8431
rect 19309 8379 19315 8431
rect 17023 8367 19315 8379
rect 17023 8315 17029 8367
rect 17081 8315 17095 8367
rect 17147 8315 17161 8367
rect 17213 8315 17227 8367
rect 17279 8315 17293 8367
rect 17345 8315 17359 8367
rect 17411 8315 17425 8367
rect 17477 8315 17491 8367
rect 17543 8315 17557 8367
rect 17609 8315 17623 8367
rect 17675 8315 17689 8367
rect 17741 8315 17755 8367
rect 17807 8315 17821 8367
rect 17873 8315 17887 8367
rect 17939 8315 17953 8367
rect 18005 8315 18019 8367
rect 18071 8315 18085 8367
rect 18137 8315 18151 8367
rect 18203 8315 18217 8367
rect 18269 8315 18282 8367
rect 18334 8315 18347 8367
rect 18399 8315 18412 8367
rect 18464 8315 18477 8367
rect 18529 8315 18542 8367
rect 18594 8315 18607 8367
rect 18659 8315 18672 8367
rect 18724 8315 18737 8367
rect 18789 8315 18802 8367
rect 18854 8315 18867 8367
rect 18919 8315 18932 8367
rect 18984 8315 18997 8367
rect 19049 8315 19062 8367
rect 19114 8315 19127 8367
rect 19179 8315 19192 8367
rect 19244 8315 19257 8367
rect 19309 8315 19315 8367
rect 20696 8443 20702 8495
rect 20754 8443 20768 8495
rect 20820 8443 20834 8495
rect 20886 8443 20900 8495
rect 20952 8443 20966 8495
rect 21018 8443 21032 8495
rect 21084 8443 21097 8495
rect 21149 8443 21162 8495
rect 21214 8443 21227 8495
rect 21279 8443 21292 8495
rect 21344 8443 21357 8495
rect 21409 8443 21415 8495
rect 20696 8431 21415 8443
rect 20696 8379 20702 8431
rect 20754 8379 20768 8431
rect 20820 8379 20834 8431
rect 20886 8379 20900 8431
rect 20952 8379 20966 8431
rect 21018 8379 21032 8431
rect 21084 8379 21097 8431
rect 21149 8379 21162 8431
rect 21214 8379 21227 8431
rect 21279 8379 21292 8431
rect 21344 8379 21357 8431
rect 21409 8379 21415 8431
rect 20696 8367 21415 8379
rect 20696 8315 20702 8367
rect 20754 8315 20768 8367
rect 20820 8315 20834 8367
rect 20886 8315 20900 8367
rect 20952 8315 20966 8367
rect 21018 8315 21032 8367
rect 21084 8315 21097 8367
rect 21149 8315 21162 8367
rect 21214 8315 21227 8367
rect 21279 8315 21292 8367
rect 21344 8315 21357 8367
rect 21409 8315 21415 8367
rect 22716 8491 23486 8530
rect 22716 8457 22798 8491
rect 22832 8457 22870 8491
rect 22904 8457 22942 8491
rect 22976 8457 23014 8491
rect 23048 8457 23086 8491
rect 23120 8457 23158 8491
rect 23192 8457 23230 8491
rect 23264 8457 23302 8491
rect 23336 8457 23374 8491
rect 23408 8457 23446 8491
rect 23480 8457 23486 8491
rect 22716 8418 23486 8457
rect 22716 8384 22798 8418
rect 22832 8384 22870 8418
rect 22904 8384 22942 8418
rect 22976 8384 23014 8418
rect 23048 8384 23086 8418
rect 23120 8384 23158 8418
rect 23192 8384 23230 8418
rect 23264 8384 23302 8418
rect 23336 8384 23374 8418
rect 23408 8384 23446 8418
rect 23480 8384 23486 8418
rect 22716 8345 23486 8384
rect 22716 8311 22798 8345
rect 22832 8311 22870 8345
rect 22904 8311 22942 8345
rect 22976 8311 23014 8345
rect 23048 8311 23086 8345
rect 23120 8311 23158 8345
rect 23192 8311 23230 8345
rect 23264 8311 23302 8345
rect 23336 8311 23374 8345
rect 23408 8311 23446 8345
rect 23480 8311 23486 8345
rect 22716 8272 23486 8311
rect 22716 8238 22798 8272
rect 22832 8238 22870 8272
rect 22904 8238 22942 8272
rect 22976 8238 23014 8272
rect 23048 8238 23086 8272
rect 23120 8238 23158 8272
rect 23192 8238 23230 8272
rect 23264 8238 23302 8272
rect 23336 8238 23374 8272
rect 23408 8238 23446 8272
rect 23480 8238 23486 8272
rect 17023 8179 17029 8231
rect 17081 8179 17095 8231
rect 17147 8179 17161 8231
rect 17213 8179 17227 8231
rect 17279 8179 17293 8231
rect 17345 8179 17359 8231
rect 17411 8179 17425 8231
rect 17477 8179 17491 8231
rect 17543 8179 17557 8231
rect 17609 8179 17623 8231
rect 17675 8179 17689 8231
rect 17741 8179 17755 8231
rect 17807 8179 17821 8231
rect 17873 8179 17887 8231
rect 17939 8179 17953 8231
rect 18005 8179 18019 8231
rect 18071 8179 18085 8231
rect 18137 8179 18151 8231
rect 18203 8179 18217 8231
rect 18269 8179 18282 8231
rect 18334 8179 18347 8231
rect 18399 8179 18412 8231
rect 18464 8179 18477 8231
rect 18529 8179 18542 8231
rect 18594 8179 18607 8231
rect 18659 8179 18672 8231
rect 18724 8179 18737 8231
rect 18789 8179 18802 8231
rect 18854 8179 18867 8231
rect 18919 8179 18932 8231
rect 18984 8179 18997 8231
rect 19049 8179 19062 8231
rect 19114 8179 19127 8231
rect 19179 8179 19192 8231
rect 19244 8179 19257 8231
rect 19309 8179 19315 8231
rect 17023 8167 19315 8179
rect 17023 8115 17029 8167
rect 17081 8115 17095 8167
rect 17147 8115 17161 8167
rect 17213 8115 17227 8167
rect 17279 8115 17293 8167
rect 17345 8115 17359 8167
rect 17411 8115 17425 8167
rect 17477 8115 17491 8167
rect 17543 8115 17557 8167
rect 17609 8115 17623 8167
rect 17675 8115 17689 8167
rect 17741 8115 17755 8167
rect 17807 8115 17821 8167
rect 17873 8115 17887 8167
rect 17939 8115 17953 8167
rect 18005 8115 18019 8167
rect 18071 8115 18085 8167
rect 18137 8115 18151 8167
rect 18203 8115 18217 8167
rect 18269 8115 18282 8167
rect 18334 8115 18347 8167
rect 18399 8115 18412 8167
rect 18464 8115 18477 8167
rect 18529 8115 18542 8167
rect 18594 8115 18607 8167
rect 18659 8115 18672 8167
rect 18724 8115 18737 8167
rect 18789 8115 18802 8167
rect 18854 8115 18867 8167
rect 18919 8115 18932 8167
rect 18984 8115 18997 8167
rect 19049 8115 19062 8167
rect 19114 8115 19127 8167
rect 19179 8115 19192 8167
rect 19244 8115 19257 8167
rect 19309 8115 19315 8167
rect 17023 8103 19315 8115
rect 17023 8051 17029 8103
rect 17081 8051 17095 8103
rect 17147 8051 17161 8103
rect 17213 8051 17227 8103
rect 17279 8051 17293 8103
rect 17345 8051 17359 8103
rect 17411 8051 17425 8103
rect 17477 8051 17491 8103
rect 17543 8051 17557 8103
rect 17609 8051 17623 8103
rect 17675 8051 17689 8103
rect 17741 8051 17755 8103
rect 17807 8051 17821 8103
rect 17873 8051 17887 8103
rect 17939 8051 17953 8103
rect 18005 8051 18019 8103
rect 18071 8051 18085 8103
rect 18137 8051 18151 8103
rect 18203 8051 18217 8103
rect 18269 8051 18282 8103
rect 18334 8051 18347 8103
rect 18399 8051 18412 8103
rect 18464 8051 18477 8103
rect 18529 8051 18542 8103
rect 18594 8051 18607 8103
rect 18659 8051 18672 8103
rect 18724 8051 18737 8103
rect 18789 8051 18802 8103
rect 18854 8051 18867 8103
rect 18919 8051 18932 8103
rect 18984 8051 18997 8103
rect 19049 8051 19062 8103
rect 19114 8051 19127 8103
rect 19179 8051 19192 8103
rect 19244 8051 19257 8103
rect 19309 8051 19315 8103
rect 20696 8179 20702 8231
rect 20754 8179 20768 8231
rect 20820 8179 20834 8231
rect 20886 8179 20900 8231
rect 20952 8179 20966 8231
rect 21018 8179 21032 8231
rect 21084 8179 21097 8231
rect 21149 8179 21162 8231
rect 21214 8179 21227 8231
rect 21279 8179 21292 8231
rect 21344 8179 21357 8231
rect 21409 8179 21415 8231
rect 20696 8167 21415 8179
rect 20696 8115 20702 8167
rect 20754 8115 20768 8167
rect 20820 8115 20834 8167
rect 20886 8115 20900 8167
rect 20952 8115 20966 8167
rect 21018 8115 21032 8167
rect 21084 8115 21097 8167
rect 21149 8115 21162 8167
rect 21214 8115 21227 8167
rect 21279 8115 21292 8167
rect 21344 8115 21357 8167
rect 21409 8115 21415 8167
rect 20696 8103 21415 8115
rect 20696 8051 20702 8103
rect 20754 8051 20768 8103
rect 20820 8051 20834 8103
rect 20886 8051 20900 8103
rect 20952 8051 20966 8103
rect 21018 8051 21032 8103
rect 21084 8051 21097 8103
rect 21149 8051 21162 8103
rect 21214 8051 21227 8103
rect 21279 8051 21292 8103
rect 21344 8051 21357 8103
rect 21409 8051 21415 8103
rect 22716 8199 23486 8238
rect 22716 8165 22798 8199
rect 22832 8165 22870 8199
rect 22904 8165 22942 8199
rect 22976 8165 23014 8199
rect 23048 8165 23086 8199
rect 23120 8165 23158 8199
rect 23192 8165 23230 8199
rect 23264 8165 23302 8199
rect 23336 8165 23374 8199
rect 23408 8165 23446 8199
rect 23480 8165 23486 8199
rect 22716 8126 23486 8165
rect 22716 8092 22798 8126
rect 22832 8092 22870 8126
rect 22904 8092 22942 8126
rect 22976 8092 23014 8126
rect 23048 8092 23086 8126
rect 23120 8092 23158 8126
rect 23192 8092 23230 8126
rect 23264 8092 23302 8126
rect 23336 8092 23374 8126
rect 23408 8092 23446 8126
rect 23480 8092 23486 8126
rect 22716 8053 23486 8092
rect 22716 8019 22798 8053
rect 22832 8019 22870 8053
rect 22904 8019 22942 8053
rect 22976 8019 23014 8053
rect 23048 8019 23086 8053
rect 23120 8019 23158 8053
rect 23192 8019 23230 8053
rect 23264 8019 23302 8053
rect 23336 8019 23374 8053
rect 23408 8019 23446 8053
rect 23480 8019 23486 8053
rect 22716 7980 23486 8019
rect 17023 7915 17029 7967
rect 17081 7915 17095 7967
rect 17147 7915 17161 7967
rect 17213 7915 17227 7967
rect 17279 7915 17293 7967
rect 17345 7915 17359 7967
rect 17411 7915 17425 7967
rect 17477 7915 17491 7967
rect 17543 7915 17557 7967
rect 17609 7915 17623 7967
rect 17675 7915 17689 7967
rect 17741 7915 17755 7967
rect 17807 7915 17821 7967
rect 17873 7915 17887 7967
rect 17939 7915 17953 7967
rect 18005 7915 18019 7967
rect 18071 7915 18085 7967
rect 18137 7915 18151 7967
rect 18203 7915 18217 7967
rect 18269 7915 18282 7967
rect 18334 7915 18347 7967
rect 18399 7915 18412 7967
rect 18464 7915 18477 7967
rect 18529 7915 18542 7967
rect 18594 7915 18607 7967
rect 18659 7915 18672 7967
rect 18724 7915 18737 7967
rect 18789 7915 18802 7967
rect 18854 7915 18867 7967
rect 18919 7915 18932 7967
rect 18984 7915 18997 7967
rect 19049 7915 19062 7967
rect 19114 7915 19127 7967
rect 19179 7915 19192 7967
rect 19244 7915 19257 7967
rect 19309 7915 19315 7967
rect 17023 7903 19315 7915
rect 17023 7851 17029 7903
rect 17081 7851 17095 7903
rect 17147 7851 17161 7903
rect 17213 7851 17227 7903
rect 17279 7851 17293 7903
rect 17345 7851 17359 7903
rect 17411 7851 17425 7903
rect 17477 7851 17491 7903
rect 17543 7851 17557 7903
rect 17609 7851 17623 7903
rect 17675 7851 17689 7903
rect 17741 7851 17755 7903
rect 17807 7851 17821 7903
rect 17873 7851 17887 7903
rect 17939 7851 17953 7903
rect 18005 7851 18019 7903
rect 18071 7851 18085 7903
rect 18137 7851 18151 7903
rect 18203 7851 18217 7903
rect 18269 7851 18282 7903
rect 18334 7851 18347 7903
rect 18399 7851 18412 7903
rect 18464 7851 18477 7903
rect 18529 7851 18542 7903
rect 18594 7851 18607 7903
rect 18659 7851 18672 7903
rect 18724 7851 18737 7903
rect 18789 7851 18802 7903
rect 18854 7851 18867 7903
rect 18919 7851 18932 7903
rect 18984 7851 18997 7903
rect 19049 7851 19062 7903
rect 19114 7851 19127 7903
rect 19179 7851 19192 7903
rect 19244 7851 19257 7903
rect 19309 7851 19315 7903
rect 17023 7839 19315 7851
rect 17023 7787 17029 7839
rect 17081 7787 17095 7839
rect 17147 7787 17161 7839
rect 17213 7787 17227 7839
rect 17279 7787 17293 7839
rect 17345 7787 17359 7839
rect 17411 7787 17425 7839
rect 17477 7787 17491 7839
rect 17543 7787 17557 7839
rect 17609 7787 17623 7839
rect 17675 7787 17689 7839
rect 17741 7787 17755 7839
rect 17807 7787 17821 7839
rect 17873 7787 17887 7839
rect 17939 7787 17953 7839
rect 18005 7787 18019 7839
rect 18071 7787 18085 7839
rect 18137 7787 18151 7839
rect 18203 7787 18217 7839
rect 18269 7787 18282 7839
rect 18334 7787 18347 7839
rect 18399 7787 18412 7839
rect 18464 7787 18477 7839
rect 18529 7787 18542 7839
rect 18594 7787 18607 7839
rect 18659 7787 18672 7839
rect 18724 7787 18737 7839
rect 18789 7787 18802 7839
rect 18854 7787 18867 7839
rect 18919 7787 18932 7839
rect 18984 7787 18997 7839
rect 19049 7787 19062 7839
rect 19114 7787 19127 7839
rect 19179 7787 19192 7839
rect 19244 7787 19257 7839
rect 19309 7787 19315 7839
rect 20696 7915 20702 7967
rect 20754 7915 20768 7967
rect 20820 7915 20834 7967
rect 20886 7915 20900 7967
rect 20952 7915 20966 7967
rect 21018 7915 21032 7967
rect 21084 7915 21097 7967
rect 21149 7915 21162 7967
rect 21214 7915 21227 7967
rect 21279 7915 21292 7967
rect 21344 7915 21357 7967
rect 21409 7915 21415 7967
rect 20696 7903 21415 7915
rect 20696 7851 20702 7903
rect 20754 7851 20768 7903
rect 20820 7851 20834 7903
rect 20886 7851 20900 7903
rect 20952 7851 20966 7903
rect 21018 7851 21032 7903
rect 21084 7851 21097 7903
rect 21149 7851 21162 7903
rect 21214 7851 21227 7903
rect 21279 7851 21292 7903
rect 21344 7851 21357 7903
rect 21409 7851 21415 7903
rect 20696 7839 21415 7851
rect 20696 7787 20702 7839
rect 20754 7787 20768 7839
rect 20820 7787 20834 7839
rect 20886 7787 20900 7839
rect 20952 7787 20966 7839
rect 21018 7787 21032 7839
rect 21084 7787 21097 7839
rect 21149 7787 21162 7839
rect 21214 7787 21227 7839
rect 21279 7787 21292 7839
rect 21344 7787 21357 7839
rect 21409 7787 21415 7839
rect 22716 7946 22798 7980
rect 22832 7946 22870 7980
rect 22904 7946 22942 7980
rect 22976 7946 23014 7980
rect 23048 7946 23086 7980
rect 23120 7946 23158 7980
rect 23192 7946 23230 7980
rect 23264 7946 23302 7980
rect 23336 7946 23374 7980
rect 23408 7946 23446 7980
rect 23480 7946 23486 7980
rect 22716 7907 23486 7946
rect 22716 7873 22798 7907
rect 22832 7873 22870 7907
rect 22904 7873 22942 7907
rect 22976 7873 23014 7907
rect 23048 7873 23086 7907
rect 23120 7873 23158 7907
rect 23192 7873 23230 7907
rect 23264 7873 23302 7907
rect 23336 7873 23374 7907
rect 23408 7873 23446 7907
rect 23480 7873 23486 7907
rect 22716 7834 23486 7873
rect 22716 7800 22798 7834
rect 22832 7800 22870 7834
rect 22904 7800 22942 7834
rect 22976 7800 23014 7834
rect 23048 7800 23086 7834
rect 23120 7800 23158 7834
rect 23192 7800 23230 7834
rect 23264 7800 23302 7834
rect 23336 7800 23374 7834
rect 23408 7800 23446 7834
rect 23480 7800 23486 7834
rect 22716 7761 23486 7800
rect 22716 7727 22798 7761
rect 22832 7727 22870 7761
rect 22904 7727 22942 7761
rect 22976 7727 23014 7761
rect 23048 7727 23086 7761
rect 23120 7727 23158 7761
rect 23192 7727 23230 7761
rect 23264 7727 23302 7761
rect 23336 7727 23374 7761
rect 23408 7727 23446 7761
rect 23480 7727 23486 7761
rect 17023 7651 17029 7703
rect 17081 7651 17095 7703
rect 17147 7651 17161 7703
rect 17213 7651 17227 7703
rect 17279 7651 17293 7703
rect 17345 7651 17359 7703
rect 17411 7651 17425 7703
rect 17477 7651 17491 7703
rect 17543 7651 17557 7703
rect 17609 7651 17623 7703
rect 17675 7651 17689 7703
rect 17741 7651 17755 7703
rect 17807 7651 17821 7703
rect 17873 7651 17887 7703
rect 17939 7651 17953 7703
rect 18005 7651 18019 7703
rect 18071 7651 18085 7703
rect 18137 7651 18151 7703
rect 18203 7651 18217 7703
rect 18269 7651 18282 7703
rect 18334 7651 18347 7703
rect 18399 7651 18412 7703
rect 18464 7651 18477 7703
rect 18529 7651 18542 7703
rect 18594 7651 18607 7703
rect 18659 7651 18672 7703
rect 18724 7651 18737 7703
rect 18789 7651 18802 7703
rect 18854 7651 18867 7703
rect 18919 7651 18932 7703
rect 18984 7651 18997 7703
rect 19049 7651 19062 7703
rect 19114 7651 19127 7703
rect 19179 7651 19192 7703
rect 19244 7651 19257 7703
rect 19309 7651 19315 7703
rect 17023 7639 19315 7651
rect 17023 7587 17029 7639
rect 17081 7587 17095 7639
rect 17147 7587 17161 7639
rect 17213 7587 17227 7639
rect 17279 7587 17293 7639
rect 17345 7587 17359 7639
rect 17411 7587 17425 7639
rect 17477 7587 17491 7639
rect 17543 7587 17557 7639
rect 17609 7587 17623 7639
rect 17675 7587 17689 7639
rect 17741 7587 17755 7639
rect 17807 7587 17821 7639
rect 17873 7587 17887 7639
rect 17939 7587 17953 7639
rect 18005 7587 18019 7639
rect 18071 7587 18085 7639
rect 18137 7587 18151 7639
rect 18203 7587 18217 7639
rect 18269 7587 18282 7639
rect 18334 7587 18347 7639
rect 18399 7587 18412 7639
rect 18464 7587 18477 7639
rect 18529 7587 18542 7639
rect 18594 7587 18607 7639
rect 18659 7587 18672 7639
rect 18724 7587 18737 7639
rect 18789 7587 18802 7639
rect 18854 7587 18867 7639
rect 18919 7587 18932 7639
rect 18984 7587 18997 7639
rect 19049 7587 19062 7639
rect 19114 7587 19127 7639
rect 19179 7587 19192 7639
rect 19244 7587 19257 7639
rect 19309 7587 19315 7639
rect 17023 7575 19315 7587
rect 17023 7523 17029 7575
rect 17081 7523 17095 7575
rect 17147 7523 17161 7575
rect 17213 7523 17227 7575
rect 17279 7523 17293 7575
rect 17345 7523 17359 7575
rect 17411 7523 17425 7575
rect 17477 7523 17491 7575
rect 17543 7523 17557 7575
rect 17609 7523 17623 7575
rect 17675 7523 17689 7575
rect 17741 7523 17755 7575
rect 17807 7523 17821 7575
rect 17873 7523 17887 7575
rect 17939 7523 17953 7575
rect 18005 7523 18019 7575
rect 18071 7523 18085 7575
rect 18137 7523 18151 7575
rect 18203 7523 18217 7575
rect 18269 7523 18282 7575
rect 18334 7523 18347 7575
rect 18399 7523 18412 7575
rect 18464 7523 18477 7575
rect 18529 7523 18542 7575
rect 18594 7523 18607 7575
rect 18659 7523 18672 7575
rect 18724 7523 18737 7575
rect 18789 7523 18802 7575
rect 18854 7523 18867 7575
rect 18919 7523 18932 7575
rect 18984 7523 18997 7575
rect 19049 7523 19062 7575
rect 19114 7523 19127 7575
rect 19179 7523 19192 7575
rect 19244 7523 19257 7575
rect 19309 7523 19315 7575
rect 20696 7651 20702 7703
rect 20754 7651 20768 7703
rect 20820 7651 20834 7703
rect 20886 7651 20900 7703
rect 20952 7651 20966 7703
rect 21018 7651 21032 7703
rect 21084 7651 21097 7703
rect 21149 7651 21162 7703
rect 21214 7651 21227 7703
rect 21279 7651 21292 7703
rect 21344 7651 21357 7703
rect 21409 7651 21415 7703
rect 20696 7639 21415 7651
rect 20696 7587 20702 7639
rect 20754 7587 20768 7639
rect 20820 7587 20834 7639
rect 20886 7587 20900 7639
rect 20952 7587 20966 7639
rect 21018 7587 21032 7639
rect 21084 7587 21097 7639
rect 21149 7587 21162 7639
rect 21214 7587 21227 7639
rect 21279 7587 21292 7639
rect 21344 7587 21357 7639
rect 21409 7587 21415 7639
rect 20696 7575 21415 7587
rect 20696 7523 20702 7575
rect 20754 7523 20768 7575
rect 20820 7523 20834 7575
rect 20886 7523 20900 7575
rect 20952 7523 20966 7575
rect 21018 7523 21032 7575
rect 21084 7523 21097 7575
rect 21149 7523 21162 7575
rect 21214 7523 21227 7575
rect 21279 7523 21292 7575
rect 21344 7523 21357 7575
rect 21409 7523 21415 7575
rect 22716 7688 23486 7727
rect 22716 7654 22798 7688
rect 22832 7654 22870 7688
rect 22904 7654 22942 7688
rect 22976 7654 23014 7688
rect 23048 7654 23086 7688
rect 23120 7654 23158 7688
rect 23192 7654 23230 7688
rect 23264 7654 23302 7688
rect 23336 7654 23374 7688
rect 23408 7654 23446 7688
rect 23480 7654 23486 7688
rect 22716 7615 23486 7654
rect 22716 7581 22798 7615
rect 22832 7581 22870 7615
rect 22904 7581 22942 7615
rect 22976 7581 23014 7615
rect 23048 7581 23086 7615
rect 23120 7581 23158 7615
rect 23192 7581 23230 7615
rect 23264 7581 23302 7615
rect 23336 7581 23374 7615
rect 23408 7581 23446 7615
rect 23480 7581 23486 7615
rect 22716 7542 23486 7581
rect 22716 7508 22798 7542
rect 22832 7508 22870 7542
rect 22904 7508 22942 7542
rect 22976 7508 23014 7542
rect 23048 7508 23086 7542
rect 23120 7508 23158 7542
rect 23192 7508 23230 7542
rect 23264 7508 23302 7542
rect 23336 7508 23374 7542
rect 23408 7508 23446 7542
rect 23480 7508 23486 7542
rect 22716 7469 23486 7508
rect 17023 7387 17029 7439
rect 17081 7387 17095 7439
rect 17147 7387 17161 7439
rect 17213 7387 17227 7439
rect 17279 7387 17293 7439
rect 17345 7387 17359 7439
rect 17411 7387 17425 7439
rect 17477 7387 17491 7439
rect 17543 7387 17557 7439
rect 17609 7387 17623 7439
rect 17675 7387 17689 7439
rect 17741 7387 17755 7439
rect 17807 7387 17821 7439
rect 17873 7387 17887 7439
rect 17939 7387 17953 7439
rect 18005 7387 18019 7439
rect 18071 7387 18085 7439
rect 18137 7387 18151 7439
rect 18203 7387 18217 7439
rect 18269 7387 18282 7439
rect 18334 7387 18347 7439
rect 18399 7387 18412 7439
rect 18464 7387 18477 7439
rect 18529 7387 18542 7439
rect 18594 7387 18607 7439
rect 18659 7387 18672 7439
rect 18724 7387 18737 7439
rect 18789 7387 18802 7439
rect 18854 7387 18867 7439
rect 18919 7387 18932 7439
rect 18984 7387 18997 7439
rect 19049 7387 19062 7439
rect 19114 7387 19127 7439
rect 19179 7387 19192 7439
rect 19244 7387 19257 7439
rect 19309 7387 19315 7439
rect 17023 7375 19315 7387
rect 17023 7323 17029 7375
rect 17081 7323 17095 7375
rect 17147 7323 17161 7375
rect 17213 7323 17227 7375
rect 17279 7323 17293 7375
rect 17345 7323 17359 7375
rect 17411 7323 17425 7375
rect 17477 7323 17491 7375
rect 17543 7323 17557 7375
rect 17609 7323 17623 7375
rect 17675 7323 17689 7375
rect 17741 7323 17755 7375
rect 17807 7323 17821 7375
rect 17873 7323 17887 7375
rect 17939 7323 17953 7375
rect 18005 7323 18019 7375
rect 18071 7323 18085 7375
rect 18137 7323 18151 7375
rect 18203 7323 18217 7375
rect 18269 7323 18282 7375
rect 18334 7323 18347 7375
rect 18399 7323 18412 7375
rect 18464 7323 18477 7375
rect 18529 7323 18542 7375
rect 18594 7323 18607 7375
rect 18659 7323 18672 7375
rect 18724 7323 18737 7375
rect 18789 7323 18802 7375
rect 18854 7323 18867 7375
rect 18919 7323 18932 7375
rect 18984 7323 18997 7375
rect 19049 7323 19062 7375
rect 19114 7323 19127 7375
rect 19179 7323 19192 7375
rect 19244 7323 19257 7375
rect 19309 7323 19315 7375
rect 17023 7311 19315 7323
rect 17023 7259 17029 7311
rect 17081 7259 17095 7311
rect 17147 7259 17161 7311
rect 17213 7259 17227 7311
rect 17279 7259 17293 7311
rect 17345 7259 17359 7311
rect 17411 7259 17425 7311
rect 17477 7259 17491 7311
rect 17543 7259 17557 7311
rect 17609 7259 17623 7311
rect 17675 7259 17689 7311
rect 17741 7259 17755 7311
rect 17807 7259 17821 7311
rect 17873 7259 17887 7311
rect 17939 7259 17953 7311
rect 18005 7259 18019 7311
rect 18071 7259 18085 7311
rect 18137 7259 18151 7311
rect 18203 7259 18217 7311
rect 18269 7259 18282 7311
rect 18334 7259 18347 7311
rect 18399 7259 18412 7311
rect 18464 7259 18477 7311
rect 18529 7259 18542 7311
rect 18594 7259 18607 7311
rect 18659 7259 18672 7311
rect 18724 7259 18737 7311
rect 18789 7259 18802 7311
rect 18854 7259 18867 7311
rect 18919 7259 18932 7311
rect 18984 7259 18997 7311
rect 19049 7259 19062 7311
rect 19114 7259 19127 7311
rect 19179 7259 19192 7311
rect 19244 7259 19257 7311
rect 19309 7259 19315 7311
rect 20696 7387 20702 7439
rect 20754 7387 20768 7439
rect 20820 7387 20834 7439
rect 20886 7387 20900 7439
rect 20952 7387 20966 7439
rect 21018 7387 21032 7439
rect 21084 7387 21097 7439
rect 21149 7387 21162 7439
rect 21214 7387 21227 7439
rect 21279 7387 21292 7439
rect 21344 7387 21357 7439
rect 21409 7387 21415 7439
rect 20696 7375 21415 7387
rect 20696 7323 20702 7375
rect 20754 7323 20768 7375
rect 20820 7323 20834 7375
rect 20886 7323 20900 7375
rect 20952 7323 20966 7375
rect 21018 7323 21032 7375
rect 21084 7323 21097 7375
rect 21149 7323 21162 7375
rect 21214 7323 21227 7375
rect 21279 7323 21292 7375
rect 21344 7323 21357 7375
rect 21409 7323 21415 7375
rect 20696 7311 21415 7323
rect 20696 7259 20702 7311
rect 20754 7259 20768 7311
rect 20820 7259 20834 7311
rect 20886 7259 20900 7311
rect 20952 7259 20966 7311
rect 21018 7259 21032 7311
rect 21084 7259 21097 7311
rect 21149 7259 21162 7311
rect 21214 7259 21227 7311
rect 21279 7259 21292 7311
rect 21344 7259 21357 7311
rect 21409 7259 21415 7311
rect 22716 7435 22798 7469
rect 22832 7435 22870 7469
rect 22904 7435 22942 7469
rect 22976 7435 23014 7469
rect 23048 7435 23086 7469
rect 23120 7435 23158 7469
rect 23192 7435 23230 7469
rect 23264 7435 23302 7469
rect 23336 7435 23374 7469
rect 23408 7435 23446 7469
rect 23480 7435 23486 7469
rect 22716 7396 23486 7435
rect 22716 7362 22798 7396
rect 22832 7362 22870 7396
rect 22904 7362 22942 7396
rect 22976 7362 23014 7396
rect 23048 7362 23086 7396
rect 23120 7362 23158 7396
rect 23192 7362 23230 7396
rect 23264 7362 23302 7396
rect 23336 7362 23374 7396
rect 23408 7362 23446 7396
rect 23480 7362 23486 7396
rect 22716 7323 23486 7362
rect 22716 7289 22798 7323
rect 22832 7289 22870 7323
rect 22904 7289 22942 7323
rect 22976 7289 23014 7323
rect 23048 7289 23086 7323
rect 23120 7289 23158 7323
rect 23192 7289 23230 7323
rect 23264 7289 23302 7323
rect 23336 7289 23374 7323
rect 23408 7289 23446 7323
rect 23480 7289 23486 7323
rect 22716 7250 23486 7289
rect 22716 7216 22798 7250
rect 22832 7216 22870 7250
rect 22904 7216 22942 7250
rect 22976 7216 23014 7250
rect 23048 7216 23086 7250
rect 23120 7216 23158 7250
rect 23192 7216 23230 7250
rect 23264 7216 23302 7250
rect 23336 7216 23374 7250
rect 23408 7216 23446 7250
rect 23480 7216 23486 7250
rect 22716 7177 23486 7216
rect 17023 7123 17029 7175
rect 17081 7123 17095 7175
rect 17147 7123 17161 7175
rect 17213 7123 17227 7175
rect 17279 7123 17293 7175
rect 17345 7123 17359 7175
rect 17411 7123 17425 7175
rect 17477 7123 17491 7175
rect 17543 7123 17557 7175
rect 17609 7123 17623 7175
rect 17675 7123 17689 7175
rect 17741 7123 17755 7175
rect 17807 7123 17821 7175
rect 17873 7123 17887 7175
rect 17939 7123 17953 7175
rect 18005 7123 18019 7175
rect 18071 7123 18085 7175
rect 18137 7123 18151 7175
rect 18203 7123 18217 7175
rect 18269 7123 18282 7175
rect 18334 7123 18347 7175
rect 18399 7123 18412 7175
rect 18464 7123 18477 7175
rect 18529 7123 18542 7175
rect 18594 7123 18607 7175
rect 18659 7123 18672 7175
rect 18724 7123 18737 7175
rect 18789 7123 18802 7175
rect 18854 7123 18867 7175
rect 18919 7123 18932 7175
rect 18984 7123 18997 7175
rect 19049 7123 19062 7175
rect 19114 7123 19127 7175
rect 19179 7123 19192 7175
rect 19244 7123 19257 7175
rect 19309 7123 19315 7175
rect 17023 7111 19315 7123
rect 17023 7059 17029 7111
rect 17081 7059 17095 7111
rect 17147 7059 17161 7111
rect 17213 7059 17227 7111
rect 17279 7059 17293 7111
rect 17345 7059 17359 7111
rect 17411 7059 17425 7111
rect 17477 7059 17491 7111
rect 17543 7059 17557 7111
rect 17609 7059 17623 7111
rect 17675 7059 17689 7111
rect 17741 7059 17755 7111
rect 17807 7059 17821 7111
rect 17873 7059 17887 7111
rect 17939 7059 17953 7111
rect 18005 7059 18019 7111
rect 18071 7059 18085 7111
rect 18137 7059 18151 7111
rect 18203 7059 18217 7111
rect 18269 7059 18282 7111
rect 18334 7059 18347 7111
rect 18399 7059 18412 7111
rect 18464 7059 18477 7111
rect 18529 7059 18542 7111
rect 18594 7059 18607 7111
rect 18659 7059 18672 7111
rect 18724 7059 18737 7111
rect 18789 7059 18802 7111
rect 18854 7059 18867 7111
rect 18919 7059 18932 7111
rect 18984 7059 18997 7111
rect 19049 7059 19062 7111
rect 19114 7059 19127 7111
rect 19179 7059 19192 7111
rect 19244 7059 19257 7111
rect 19309 7059 19315 7111
rect 17023 7047 19315 7059
rect 17023 6995 17029 7047
rect 17081 6995 17095 7047
rect 17147 6995 17161 7047
rect 17213 6995 17227 7047
rect 17279 6995 17293 7047
rect 17345 6995 17359 7047
rect 17411 6995 17425 7047
rect 17477 6995 17491 7047
rect 17543 6995 17557 7047
rect 17609 6995 17623 7047
rect 17675 6995 17689 7047
rect 17741 6995 17755 7047
rect 17807 6995 17821 7047
rect 17873 6995 17887 7047
rect 17939 6995 17953 7047
rect 18005 6995 18019 7047
rect 18071 6995 18085 7047
rect 18137 6995 18151 7047
rect 18203 6995 18217 7047
rect 18269 6995 18282 7047
rect 18334 6995 18347 7047
rect 18399 6995 18412 7047
rect 18464 6995 18477 7047
rect 18529 6995 18542 7047
rect 18594 6995 18607 7047
rect 18659 6995 18672 7047
rect 18724 6995 18737 7047
rect 18789 6995 18802 7047
rect 18854 6995 18867 7047
rect 18919 6995 18932 7047
rect 18984 6995 18997 7047
rect 19049 6995 19062 7047
rect 19114 6995 19127 7047
rect 19179 6995 19192 7047
rect 19244 6995 19257 7047
rect 19309 6995 19315 7047
rect 20696 7123 20702 7175
rect 20754 7123 20768 7175
rect 20820 7123 20834 7175
rect 20886 7123 20900 7175
rect 20952 7123 20966 7175
rect 21018 7123 21032 7175
rect 21084 7123 21097 7175
rect 21149 7123 21162 7175
rect 21214 7123 21227 7175
rect 21279 7123 21292 7175
rect 21344 7123 21357 7175
rect 21409 7123 21415 7175
rect 20696 7111 21415 7123
rect 20696 7059 20702 7111
rect 20754 7059 20768 7111
rect 20820 7059 20834 7111
rect 20886 7059 20900 7111
rect 20952 7059 20966 7111
rect 21018 7059 21032 7111
rect 21084 7059 21097 7111
rect 21149 7059 21162 7111
rect 21214 7059 21227 7111
rect 21279 7059 21292 7111
rect 21344 7059 21357 7111
rect 21409 7059 21415 7111
rect 20696 7047 21415 7059
rect 20696 6995 20702 7047
rect 20754 6995 20768 7047
rect 20820 6995 20834 7047
rect 20886 6995 20900 7047
rect 20952 6995 20966 7047
rect 21018 6995 21032 7047
rect 21084 6995 21097 7047
rect 21149 6995 21162 7047
rect 21214 6995 21227 7047
rect 21279 6995 21292 7047
rect 21344 6995 21357 7047
rect 21409 6995 21415 7047
rect 22716 7143 22798 7177
rect 22832 7143 22870 7177
rect 22904 7143 22942 7177
rect 22976 7143 23014 7177
rect 23048 7143 23086 7177
rect 23120 7143 23158 7177
rect 23192 7143 23230 7177
rect 23264 7143 23302 7177
rect 23336 7143 23374 7177
rect 23408 7143 23446 7177
rect 23480 7143 23486 7177
rect 22716 7104 23486 7143
rect 22716 7070 22798 7104
rect 22832 7070 22870 7104
rect 22904 7070 22942 7104
rect 22976 7070 23014 7104
rect 23048 7070 23086 7104
rect 23120 7070 23158 7104
rect 23192 7070 23230 7104
rect 23264 7070 23302 7104
rect 23336 7070 23374 7104
rect 23408 7070 23446 7104
rect 23480 7070 23486 7104
rect 22716 7031 23486 7070
rect 22716 6997 22798 7031
rect 22832 6997 22870 7031
rect 22904 6997 22942 7031
rect 22976 6997 23014 7031
rect 23048 6997 23086 7031
rect 23120 6997 23158 7031
rect 23192 6997 23230 7031
rect 23264 6997 23302 7031
rect 23336 6997 23374 7031
rect 23408 6997 23446 7031
rect 23480 6997 23486 7031
rect 20975 6790 21921 6963
rect 22716 6958 23486 6997
rect 22716 6924 22798 6958
rect 22832 6924 22870 6958
rect 22904 6924 22942 6958
rect 22976 6924 23014 6958
rect 23048 6924 23086 6958
rect 23120 6924 23158 6958
rect 23192 6924 23230 6958
rect 23264 6924 23302 6958
rect 23336 6924 23374 6958
rect 23408 6924 23446 6958
rect 23480 6924 23486 6958
rect 22716 6885 23486 6924
rect 22716 6851 22798 6885
rect 22832 6851 22870 6885
rect 22904 6851 22942 6885
rect 22976 6851 23014 6885
rect 23048 6851 23086 6885
rect 23120 6851 23158 6885
rect 23192 6851 23230 6885
rect 23264 6851 23302 6885
rect 23336 6851 23374 6885
rect 23408 6851 23446 6885
rect 23480 6851 23486 6885
rect 22716 6812 23486 6851
rect 22716 6778 22798 6812
rect 22832 6778 22870 6812
rect 22904 6778 22942 6812
rect 22976 6778 23014 6812
rect 23048 6778 23086 6812
rect 23120 6778 23158 6812
rect 23192 6778 23230 6812
rect 23264 6778 23302 6812
rect 23336 6778 23374 6812
rect 23408 6778 23446 6812
rect 23480 6778 23486 6812
rect 22716 6739 23486 6778
rect 22716 6705 22798 6739
rect 22832 6705 22870 6739
rect 22904 6705 22942 6739
rect 22976 6705 23014 6739
rect 23048 6705 23086 6739
rect 23120 6705 23158 6739
rect 23192 6705 23230 6739
rect 23264 6705 23302 6739
rect 23336 6705 23374 6739
rect 23408 6705 23446 6739
rect 23480 6705 23486 6739
rect 20975 6526 21921 6699
rect 22716 6666 23486 6705
rect 22716 6632 22798 6666
rect 22832 6632 22870 6666
rect 22904 6632 22942 6666
rect 22976 6632 23014 6666
rect 23048 6632 23086 6666
rect 23120 6632 23158 6666
rect 23192 6632 23230 6666
rect 23264 6632 23302 6666
rect 23336 6632 23374 6666
rect 23408 6632 23446 6666
rect 23480 6632 23486 6666
rect 22716 6593 23486 6632
rect 22716 6559 22798 6593
rect 22832 6559 22870 6593
rect 22904 6559 22942 6593
rect 22976 6559 23014 6593
rect 23048 6559 23086 6593
rect 23120 6559 23158 6593
rect 23192 6559 23230 6593
rect 23264 6559 23302 6593
rect 23336 6559 23374 6593
rect 23408 6559 23446 6593
rect 23480 6559 23486 6593
rect 22716 6520 23486 6559
rect 22716 6486 22798 6520
rect 22832 6486 22870 6520
rect 22904 6486 22942 6520
rect 22976 6486 23014 6520
rect 23048 6486 23086 6520
rect 23120 6486 23158 6520
rect 23192 6486 23230 6520
rect 23264 6486 23302 6520
rect 23336 6486 23374 6520
rect 23408 6486 23446 6520
rect 23480 6486 23486 6520
rect 22716 6447 23486 6486
rect 20975 6265 21921 6438
rect 22716 6413 22798 6447
rect 22832 6413 22870 6447
rect 22904 6413 22942 6447
rect 22976 6413 23014 6447
rect 23048 6413 23086 6447
rect 23120 6413 23158 6447
rect 23192 6413 23230 6447
rect 23264 6413 23302 6447
rect 23336 6413 23374 6447
rect 23408 6413 23446 6447
rect 23480 6413 23486 6447
rect 22716 6374 23486 6413
rect 22716 6340 22798 6374
rect 22832 6340 22870 6374
rect 22904 6340 22942 6374
rect 22976 6340 23014 6374
rect 23048 6340 23086 6374
rect 23120 6340 23158 6374
rect 23192 6340 23230 6374
rect 23264 6340 23302 6374
rect 23336 6340 23374 6374
rect 23408 6340 23446 6374
rect 23480 6340 23486 6374
rect 22716 6301 23486 6340
rect 22716 6267 22798 6301
rect 22832 6267 22870 6301
rect 22904 6267 22942 6301
rect 22976 6267 23014 6301
rect 23048 6267 23086 6301
rect 23120 6267 23158 6301
rect 23192 6267 23230 6301
rect 23264 6267 23302 6301
rect 23336 6267 23374 6301
rect 23408 6267 23446 6301
rect 23480 6267 23486 6301
rect 22716 6228 23486 6267
rect 22716 6194 22798 6228
rect 22832 6194 22870 6228
rect 22904 6194 22942 6228
rect 22976 6194 23014 6228
rect 23048 6194 23086 6228
rect 23120 6194 23158 6228
rect 23192 6194 23230 6228
rect 23264 6194 23302 6228
rect 23336 6194 23374 6228
rect 23408 6194 23446 6228
rect 23480 6194 23486 6228
rect 20975 5999 21921 6172
rect 22716 6155 23486 6194
rect 22716 6121 22798 6155
rect 22832 6121 22870 6155
rect 22904 6121 22942 6155
rect 22976 6121 23014 6155
rect 23048 6121 23086 6155
rect 23120 6121 23158 6155
rect 23192 6121 23230 6155
rect 23264 6121 23302 6155
rect 23336 6121 23374 6155
rect 23408 6121 23446 6155
rect 23480 6121 23486 6155
rect 22716 6082 23486 6121
rect 22716 6048 22798 6082
rect 22832 6048 22870 6082
rect 22904 6048 22942 6082
rect 22976 6048 23014 6082
rect 23048 6048 23086 6082
rect 23120 6048 23158 6082
rect 23192 6048 23230 6082
rect 23264 6048 23302 6082
rect 23336 6048 23374 6082
rect 23408 6048 23446 6082
rect 23480 6048 23486 6082
rect 22716 6009 23486 6048
rect 22716 5975 22798 6009
rect 22832 5975 22870 6009
rect 22904 5975 22942 6009
rect 22976 5975 23014 6009
rect 23048 5975 23086 6009
rect 23120 5975 23158 6009
rect 23192 5975 23230 6009
rect 23264 5975 23302 6009
rect 23336 5975 23374 6009
rect 23408 5975 23446 6009
rect 23480 5975 23486 6009
rect 22716 5936 23486 5975
rect 20975 5734 21921 5907
rect 22716 5902 22798 5936
rect 22832 5902 22870 5936
rect 22904 5902 22942 5936
rect 22976 5902 23014 5936
rect 23048 5902 23086 5936
rect 23120 5902 23158 5936
rect 23192 5902 23230 5936
rect 23264 5902 23302 5936
rect 23336 5902 23374 5936
rect 23408 5902 23446 5936
rect 23480 5902 23486 5936
rect 22716 5863 23486 5902
rect 22716 5829 22798 5863
rect 22832 5829 22870 5863
rect 22904 5829 22942 5863
rect 22976 5829 23014 5863
rect 23048 5829 23086 5863
rect 23120 5829 23158 5863
rect 23192 5829 23230 5863
rect 23264 5829 23302 5863
rect 23336 5829 23374 5863
rect 23408 5829 23446 5863
rect 23480 5829 23486 5863
rect 22716 5790 23486 5829
rect 22716 5756 22798 5790
rect 22832 5756 22870 5790
rect 22904 5756 22942 5790
rect 22976 5756 23014 5790
rect 23048 5756 23086 5790
rect 23120 5756 23158 5790
rect 23192 5756 23230 5790
rect 23264 5756 23302 5790
rect 23336 5756 23374 5790
rect 23408 5756 23446 5790
rect 23480 5756 23486 5790
rect 22716 5717 23486 5756
rect 22716 5683 22798 5717
rect 22832 5683 22870 5717
rect 22904 5683 22942 5717
rect 22976 5683 23014 5717
rect 23048 5683 23086 5717
rect 23120 5683 23158 5717
rect 23192 5683 23230 5717
rect 23264 5683 23302 5717
rect 23336 5683 23374 5717
rect 23408 5683 23446 5717
rect 23480 5683 23486 5717
rect 22716 5644 23486 5683
rect 23775 8680 23941 9126
rect 24505 8680 24541 9126
rect 23775 7854 23781 8680
rect 24535 7854 24541 8680
rect 23775 7815 23941 7854
rect 24505 7815 24541 7854
rect 23775 7781 23781 7815
rect 23815 7781 23853 7815
rect 23887 7781 23925 7815
rect 24535 7781 24541 7815
rect 23775 7742 23941 7781
rect 24505 7742 24541 7781
rect 23775 7708 23781 7742
rect 23815 7708 23853 7742
rect 23887 7708 23925 7742
rect 24535 7708 24541 7742
rect 23775 7669 23941 7708
rect 24505 7669 24541 7708
rect 23775 7635 23781 7669
rect 23815 7635 23853 7669
rect 23887 7635 23925 7669
rect 24535 7635 24541 7669
rect 23775 7596 23941 7635
rect 24505 7596 24541 7635
rect 23775 7562 23781 7596
rect 23815 7562 23853 7596
rect 23887 7562 23925 7596
rect 24535 7562 24541 7596
rect 23775 7523 23941 7562
rect 24505 7523 24541 7562
rect 23775 7489 23781 7523
rect 23815 7489 23853 7523
rect 23887 7489 23925 7523
rect 24535 7489 24541 7523
rect 23775 7450 23941 7489
rect 24505 7450 24541 7489
rect 23775 7416 23781 7450
rect 23815 7416 23853 7450
rect 23887 7416 23925 7450
rect 24535 7416 24541 7450
rect 23775 7377 23941 7416
rect 24505 7377 24541 7416
rect 23775 7343 23781 7377
rect 23815 7343 23853 7377
rect 23887 7343 23925 7377
rect 24535 7343 24541 7377
rect 23775 7304 23941 7343
rect 24505 7304 24541 7343
rect 23775 7270 23781 7304
rect 23815 7270 23853 7304
rect 23887 7270 23925 7304
rect 24535 7270 24541 7304
rect 23775 7231 23941 7270
rect 24505 7231 24541 7270
rect 23775 7197 23781 7231
rect 23815 7197 23853 7231
rect 23887 7197 23925 7231
rect 23959 7205 23997 7218
rect 24031 7205 24069 7218
rect 24103 7205 24141 7218
rect 24175 7205 24213 7218
rect 24247 7205 24285 7218
rect 24319 7205 24357 7218
rect 24391 7205 24429 7218
rect 24463 7205 24501 7218
rect 23993 7197 23997 7205
rect 23775 7158 23941 7197
rect 23993 7158 24005 7197
rect 23775 7124 23781 7158
rect 23815 7124 23853 7158
rect 23887 7124 23925 7158
rect 23993 7153 23997 7158
rect 24057 7153 24069 7205
rect 24121 7153 24133 7205
rect 24185 7153 24197 7205
rect 24249 7153 24261 7205
rect 24319 7197 24325 7205
rect 24535 7197 24541 7231
rect 24313 7158 24325 7197
rect 24377 7158 24389 7197
rect 24441 7158 24453 7197
rect 24505 7158 24541 7197
rect 24319 7153 24325 7158
rect 23959 7140 23997 7153
rect 24031 7140 24069 7153
rect 24103 7140 24141 7153
rect 24175 7140 24213 7153
rect 24247 7140 24285 7153
rect 24319 7140 24357 7153
rect 24391 7140 24429 7153
rect 24463 7140 24501 7153
rect 23993 7124 23997 7140
rect 23775 7088 23941 7124
rect 23993 7088 24005 7124
rect 24057 7088 24069 7140
rect 24121 7088 24133 7140
rect 24185 7088 24197 7140
rect 24249 7088 24261 7140
rect 24319 7124 24325 7140
rect 24535 7124 24541 7158
rect 24313 7088 24325 7124
rect 24377 7088 24389 7124
rect 24441 7088 24453 7124
rect 24505 7088 24541 7124
rect 23775 7085 24541 7088
rect 23775 7051 23781 7085
rect 23815 7051 23853 7085
rect 23887 7051 23925 7085
rect 23959 7075 23997 7085
rect 24031 7075 24069 7085
rect 24103 7075 24141 7085
rect 24175 7075 24213 7085
rect 24247 7075 24285 7085
rect 24319 7075 24357 7085
rect 24391 7075 24429 7085
rect 24463 7075 24501 7085
rect 23993 7051 23997 7075
rect 23775 7023 23941 7051
rect 23993 7023 24005 7051
rect 24057 7023 24069 7075
rect 24121 7023 24133 7075
rect 24185 7023 24197 7075
rect 24249 7023 24261 7075
rect 24319 7051 24325 7075
rect 24535 7051 24541 7085
rect 24313 7023 24325 7051
rect 24377 7023 24389 7051
rect 24441 7023 24453 7051
rect 24505 7023 24541 7051
rect 23775 7012 24541 7023
rect 23775 6978 23781 7012
rect 23815 6978 23853 7012
rect 23887 6978 23925 7012
rect 23959 7010 23997 7012
rect 24031 7010 24069 7012
rect 24103 7010 24141 7012
rect 24175 7010 24213 7012
rect 24247 7010 24285 7012
rect 24319 7010 24357 7012
rect 24391 7010 24429 7012
rect 24463 7010 24501 7012
rect 23993 6978 23997 7010
rect 23775 6958 23941 6978
rect 23993 6958 24005 6978
rect 24057 6958 24069 7010
rect 24121 6958 24133 7010
rect 24185 6958 24197 7010
rect 24249 6958 24261 7010
rect 24319 6978 24325 7010
rect 24535 6978 24541 7012
rect 24313 6958 24325 6978
rect 24377 6958 24389 6978
rect 24441 6958 24453 6978
rect 24505 6958 24541 6978
rect 23775 6945 24541 6958
rect 25522 6948 25528 7000
rect 25580 6948 25592 7000
rect 25644 6948 28183 7000
rect 28235 6948 28271 7000
rect 28323 6948 28329 7000
rect 23775 6939 23941 6945
rect 23993 6939 24005 6945
rect 23775 6905 23781 6939
rect 23815 6905 23853 6939
rect 23887 6905 23925 6939
rect 23993 6905 23997 6939
rect 23775 6893 23941 6905
rect 23993 6893 24005 6905
rect 24057 6893 24069 6945
rect 24121 6893 24133 6945
rect 24185 6893 24197 6945
rect 24249 6893 24261 6945
rect 24313 6939 24325 6945
rect 24377 6939 24389 6945
rect 24441 6939 24453 6945
rect 24505 6939 24541 6945
rect 24319 6905 24325 6939
rect 24535 6905 24541 6939
rect 24313 6893 24325 6905
rect 24377 6893 24389 6905
rect 24441 6893 24453 6905
rect 24505 6893 24541 6905
rect 23775 6880 24541 6893
rect 23775 6866 23941 6880
rect 23993 6866 24005 6880
rect 23775 6832 23781 6866
rect 23815 6832 23853 6866
rect 23887 6832 23925 6866
rect 23993 6832 23997 6866
rect 23775 6828 23941 6832
rect 23993 6828 24005 6832
rect 24057 6828 24069 6880
rect 24121 6828 24133 6880
rect 24185 6828 24197 6880
rect 24249 6828 24261 6880
rect 24313 6866 24325 6880
rect 24377 6866 24389 6880
rect 24441 6866 24453 6880
rect 24505 6866 24541 6880
rect 24319 6832 24325 6866
rect 24535 6832 24541 6866
rect 24313 6828 24325 6832
rect 24377 6828 24389 6832
rect 24441 6828 24453 6832
rect 24505 6828 24541 6832
rect 23775 6815 24541 6828
rect 23775 6793 23941 6815
rect 23993 6793 24005 6815
rect 23775 6759 23781 6793
rect 23815 6759 23853 6793
rect 23887 6759 23925 6793
rect 23993 6763 23997 6793
rect 24057 6763 24069 6815
rect 24121 6763 24133 6815
rect 24185 6763 24197 6815
rect 24249 6763 24261 6815
rect 24313 6793 24325 6815
rect 24377 6793 24389 6815
rect 24441 6793 24453 6815
rect 24505 6793 24541 6815
rect 24319 6763 24325 6793
rect 23959 6759 23997 6763
rect 24031 6759 24069 6763
rect 24103 6759 24141 6763
rect 24175 6759 24213 6763
rect 24247 6759 24285 6763
rect 24319 6759 24357 6763
rect 24391 6759 24429 6763
rect 24463 6759 24501 6763
rect 24535 6759 24541 6793
rect 23775 6750 24541 6759
rect 23775 6720 23941 6750
rect 23993 6720 24005 6750
rect 23775 6686 23781 6720
rect 23815 6686 23853 6720
rect 23887 6686 23925 6720
rect 23993 6698 23997 6720
rect 24057 6698 24069 6750
rect 24121 6698 24133 6750
rect 24185 6698 24197 6750
rect 24249 6698 24261 6750
rect 24313 6720 24325 6750
rect 24377 6720 24389 6750
rect 24441 6720 24453 6750
rect 24505 6720 24541 6750
rect 24319 6698 24325 6720
rect 23959 6686 23997 6698
rect 24031 6686 24069 6698
rect 24103 6686 24141 6698
rect 24175 6686 24213 6698
rect 24247 6686 24285 6698
rect 24319 6686 24357 6698
rect 24391 6686 24429 6698
rect 24463 6686 24501 6698
rect 24535 6686 24541 6720
rect 23775 6685 24541 6686
rect 23775 6647 23941 6685
rect 23993 6647 24005 6685
rect 23775 6613 23781 6647
rect 23815 6613 23853 6647
rect 23887 6613 23925 6647
rect 23993 6633 23997 6647
rect 24057 6633 24069 6685
rect 24121 6633 24133 6685
rect 24185 6633 24197 6685
rect 24249 6633 24261 6685
rect 24313 6647 24325 6685
rect 24377 6647 24389 6685
rect 24441 6647 24453 6685
rect 24505 6647 24541 6685
rect 24319 6633 24325 6647
rect 23959 6620 23997 6633
rect 24031 6620 24069 6633
rect 24103 6620 24141 6633
rect 24175 6620 24213 6633
rect 24247 6620 24285 6633
rect 24319 6620 24357 6633
rect 24391 6620 24429 6633
rect 24463 6620 24501 6633
rect 23993 6613 23997 6620
rect 23775 6574 23941 6613
rect 23993 6574 24005 6613
rect 23775 6540 23781 6574
rect 23815 6540 23853 6574
rect 23887 6540 23925 6574
rect 23993 6568 23997 6574
rect 24057 6568 24069 6620
rect 24121 6568 24133 6620
rect 24185 6568 24197 6620
rect 24249 6568 24261 6620
rect 24319 6613 24325 6620
rect 24535 6613 24541 6647
rect 24313 6574 24325 6613
rect 24377 6574 24389 6613
rect 24441 6574 24453 6613
rect 24505 6574 24541 6613
rect 24319 6568 24325 6574
rect 23959 6555 23997 6568
rect 24031 6555 24069 6568
rect 24103 6555 24141 6568
rect 24175 6555 24213 6568
rect 24247 6555 24285 6568
rect 24319 6555 24357 6568
rect 24391 6555 24429 6568
rect 24463 6555 24501 6568
rect 23993 6540 23997 6555
rect 23775 6503 23941 6540
rect 23993 6503 24005 6540
rect 24057 6503 24069 6555
rect 24121 6503 24133 6555
rect 24185 6503 24197 6555
rect 24249 6503 24261 6555
rect 24319 6540 24325 6555
rect 24535 6540 24541 6574
rect 24313 6503 24325 6540
rect 24377 6503 24389 6540
rect 24441 6503 24453 6540
rect 24505 6503 24541 6540
rect 23775 6501 24541 6503
rect 23775 6467 23781 6501
rect 23815 6467 23853 6501
rect 23887 6467 23925 6501
rect 23959 6490 23997 6501
rect 24031 6490 24069 6501
rect 24103 6490 24141 6501
rect 24175 6490 24213 6501
rect 24247 6490 24285 6501
rect 24319 6490 24357 6501
rect 24391 6490 24429 6501
rect 24463 6490 24501 6501
rect 23993 6467 23997 6490
rect 23775 6438 23941 6467
rect 23993 6438 24005 6467
rect 24057 6438 24069 6490
rect 24121 6438 24133 6490
rect 24185 6438 24197 6490
rect 24249 6438 24261 6490
rect 24319 6467 24325 6490
rect 24535 6467 24541 6501
rect 24313 6438 24325 6467
rect 24377 6438 24389 6467
rect 24441 6438 24453 6467
rect 24505 6438 24541 6467
rect 23775 6428 24541 6438
rect 23775 6394 23781 6428
rect 23815 6394 23853 6428
rect 23887 6394 23925 6428
rect 23959 6425 23997 6428
rect 24031 6425 24069 6428
rect 24103 6425 24141 6428
rect 24175 6425 24213 6428
rect 24247 6425 24285 6428
rect 24319 6425 24357 6428
rect 24391 6425 24429 6428
rect 24463 6425 24501 6428
rect 23993 6394 23997 6425
rect 23775 6373 23941 6394
rect 23993 6373 24005 6394
rect 24057 6373 24069 6425
rect 24121 6373 24133 6425
rect 24185 6373 24197 6425
rect 24249 6373 24261 6425
rect 24319 6394 24325 6425
rect 24535 6394 24541 6428
rect 24313 6373 24325 6394
rect 24377 6373 24389 6394
rect 24441 6373 24453 6394
rect 24505 6373 24541 6394
rect 23775 6360 24541 6373
rect 23775 6355 23941 6360
rect 23993 6355 24005 6360
rect 23775 6321 23781 6355
rect 23815 6321 23853 6355
rect 23887 6321 23925 6355
rect 23993 6321 23997 6355
rect 23775 6308 23941 6321
rect 23993 6308 24005 6321
rect 24057 6308 24069 6360
rect 24121 6308 24133 6360
rect 24185 6308 24197 6360
rect 24249 6308 24261 6360
rect 24313 6355 24325 6360
rect 24377 6355 24389 6360
rect 24441 6355 24453 6360
rect 24505 6355 24541 6360
rect 24319 6321 24325 6355
rect 24535 6321 24541 6355
rect 24313 6308 24325 6321
rect 24377 6308 24389 6321
rect 24441 6308 24453 6321
rect 24505 6308 24541 6321
rect 23775 6295 24541 6308
rect 23775 6282 23941 6295
rect 23993 6282 24005 6295
rect 23775 6248 23781 6282
rect 23815 6248 23853 6282
rect 23887 6248 23925 6282
rect 23993 6248 23997 6282
rect 23775 6243 23941 6248
rect 23993 6243 24005 6248
rect 24057 6243 24069 6295
rect 24121 6243 24133 6295
rect 24185 6243 24197 6295
rect 24249 6243 24261 6295
rect 24313 6282 24325 6295
rect 24377 6282 24389 6295
rect 24441 6282 24453 6295
rect 24505 6282 24541 6295
rect 24319 6248 24325 6282
rect 24535 6248 24541 6282
rect 24313 6243 24325 6248
rect 24377 6243 24389 6248
rect 24441 6243 24453 6248
rect 24505 6243 24541 6248
rect 23775 6230 24541 6243
rect 23775 6209 23941 6230
rect 23993 6209 24005 6230
rect 23775 6175 23781 6209
rect 23815 6175 23853 6209
rect 23887 6175 23925 6209
rect 23993 6178 23997 6209
rect 24057 6178 24069 6230
rect 24121 6178 24133 6230
rect 24185 6178 24197 6230
rect 24249 6178 24261 6230
rect 24313 6209 24325 6230
rect 24377 6209 24389 6230
rect 24441 6209 24453 6230
rect 24505 6209 24541 6230
rect 24319 6178 24325 6209
rect 23959 6175 23997 6178
rect 24031 6175 24069 6178
rect 24103 6175 24141 6178
rect 24175 6175 24213 6178
rect 24247 6175 24285 6178
rect 24319 6175 24357 6178
rect 24391 6175 24429 6178
rect 24463 6175 24501 6178
rect 24535 6175 24541 6209
rect 23775 6165 24541 6175
rect 23775 6136 23941 6165
rect 23993 6136 24005 6165
rect 23775 6102 23781 6136
rect 23815 6102 23853 6136
rect 23887 6102 23925 6136
rect 23993 6113 23997 6136
rect 24057 6113 24069 6165
rect 24121 6113 24133 6165
rect 24185 6113 24197 6165
rect 24249 6113 24261 6165
rect 24313 6136 24325 6165
rect 24377 6136 24389 6165
rect 24441 6136 24453 6165
rect 24505 6136 24541 6165
rect 24319 6113 24325 6136
rect 23959 6102 23997 6113
rect 24031 6102 24069 6113
rect 24103 6102 24141 6113
rect 24175 6102 24213 6113
rect 24247 6102 24285 6113
rect 24319 6102 24357 6113
rect 24391 6102 24429 6113
rect 24463 6102 24501 6113
rect 24535 6102 24541 6136
rect 23775 6100 24541 6102
rect 23775 6063 23941 6100
rect 23993 6063 24005 6100
rect 23775 6029 23781 6063
rect 23815 6029 23853 6063
rect 23887 6029 23925 6063
rect 23993 6048 23997 6063
rect 24057 6048 24069 6100
rect 24121 6048 24133 6100
rect 24185 6048 24197 6100
rect 24249 6048 24261 6100
rect 24313 6063 24325 6100
rect 24377 6063 24389 6100
rect 24441 6063 24453 6100
rect 24505 6063 24541 6100
rect 24319 6048 24325 6063
rect 23959 6035 23997 6048
rect 24031 6035 24069 6048
rect 24103 6035 24141 6048
rect 24175 6035 24213 6048
rect 24247 6035 24285 6048
rect 24319 6035 24357 6048
rect 24391 6035 24429 6048
rect 24463 6035 24501 6048
rect 23993 6029 23997 6035
rect 23775 5990 23941 6029
rect 23993 5990 24005 6029
rect 23775 5956 23781 5990
rect 23815 5956 23853 5990
rect 23887 5956 23925 5990
rect 23993 5983 23997 5990
rect 24057 5983 24069 6035
rect 24121 5983 24133 6035
rect 24185 5983 24197 6035
rect 24249 5983 24261 6035
rect 24319 6029 24325 6035
rect 24535 6029 24541 6063
rect 24313 5990 24325 6029
rect 24377 5990 24389 6029
rect 24441 5990 24453 6029
rect 24505 5990 24541 6029
rect 24319 5983 24325 5990
rect 23959 5970 23997 5983
rect 24031 5970 24069 5983
rect 24103 5970 24141 5983
rect 24175 5970 24213 5983
rect 24247 5970 24285 5983
rect 24319 5970 24357 5983
rect 24391 5970 24429 5983
rect 24463 5970 24501 5983
rect 23993 5956 23997 5970
rect 23775 5918 23941 5956
rect 23993 5918 24005 5956
rect 24057 5918 24069 5970
rect 24121 5918 24133 5970
rect 24185 5918 24197 5970
rect 24249 5918 24261 5970
rect 24319 5956 24325 5970
rect 24535 5956 24541 5990
rect 24313 5918 24325 5956
rect 24377 5918 24389 5956
rect 24441 5918 24453 5956
rect 24505 5918 24541 5956
rect 23775 5917 24541 5918
rect 23775 5883 23781 5917
rect 23815 5883 23853 5917
rect 23887 5883 23925 5917
rect 23959 5905 23997 5917
rect 24031 5905 24069 5917
rect 24103 5905 24141 5917
rect 24175 5905 24213 5917
rect 24247 5905 24285 5917
rect 24319 5905 24357 5917
rect 24391 5905 24429 5917
rect 24463 5905 24501 5917
rect 23993 5883 23997 5905
rect 23775 5853 23941 5883
rect 23993 5853 24005 5883
rect 24057 5853 24069 5905
rect 24121 5853 24133 5905
rect 24185 5853 24197 5905
rect 24249 5853 24261 5905
rect 24319 5883 24325 5905
rect 24535 5883 24541 5917
rect 24313 5853 24325 5883
rect 24377 5853 24389 5883
rect 24441 5853 24453 5883
rect 24505 5853 24541 5883
rect 23775 5844 24541 5853
rect 23775 5810 23781 5844
rect 23815 5810 23853 5844
rect 23887 5810 23925 5844
rect 23959 5840 23997 5844
rect 24031 5840 24069 5844
rect 24103 5840 24141 5844
rect 24175 5840 24213 5844
rect 24247 5840 24285 5844
rect 24319 5840 24357 5844
rect 24391 5840 24429 5844
rect 24463 5840 24501 5844
rect 23993 5810 23997 5840
rect 23775 5788 23941 5810
rect 23993 5788 24005 5810
rect 24057 5788 24069 5840
rect 24121 5788 24133 5840
rect 24185 5788 24197 5840
rect 24249 5788 24261 5840
rect 24319 5810 24325 5840
rect 24535 5810 24541 5844
rect 24313 5788 24325 5810
rect 24377 5788 24389 5810
rect 24441 5788 24453 5810
rect 24505 5788 24541 5810
rect 23775 5775 24541 5788
rect 23775 5771 23941 5775
rect 23993 5771 24005 5775
rect 23775 5737 23781 5771
rect 23815 5737 23853 5771
rect 23887 5737 23925 5771
rect 23993 5737 23997 5771
rect 23775 5723 23941 5737
rect 23993 5723 24005 5737
rect 24057 5723 24069 5775
rect 24121 5723 24133 5775
rect 24185 5723 24197 5775
rect 24249 5723 24261 5775
rect 24313 5771 24325 5775
rect 24377 5771 24389 5775
rect 24441 5771 24453 5775
rect 24505 5771 24541 5775
rect 24319 5737 24325 5771
rect 24535 5737 24541 5771
rect 24313 5723 24325 5737
rect 24377 5723 24389 5737
rect 24441 5723 24453 5737
rect 24505 5723 24541 5737
rect 23775 5710 24541 5723
rect 23775 5698 23941 5710
rect 23993 5698 24005 5710
rect 24057 5698 24069 5710
rect 23775 5664 23781 5698
rect 23815 5664 23853 5698
rect 23887 5664 23925 5698
rect 23775 5658 23941 5664
rect 24121 5658 24133 5710
rect 24185 5658 24197 5710
rect 24249 5658 24261 5710
rect 24313 5698 24325 5710
rect 24377 5698 24389 5710
rect 24441 5698 24453 5710
rect 24505 5698 24541 5710
rect 24319 5664 24325 5698
rect 24535 5664 24541 5698
rect 24313 5658 24325 5664
rect 24377 5658 24389 5664
rect 24441 5658 24453 5664
rect 24505 5658 24541 5664
rect 23775 5652 23981 5658
rect 20975 5470 21921 5643
rect 22716 5610 22798 5644
rect 22832 5610 22870 5644
rect 22904 5610 22942 5644
rect 22976 5610 23014 5644
rect 23048 5610 23086 5644
rect 23120 5610 23158 5644
rect 23192 5610 23230 5644
rect 23264 5610 23302 5644
rect 23336 5610 23374 5644
rect 23408 5610 23446 5644
rect 23480 5610 23486 5644
rect 22716 5571 23486 5610
rect 22716 5537 22798 5571
rect 22832 5537 22870 5571
rect 22904 5537 22942 5571
rect 22976 5537 23014 5571
rect 23048 5537 23086 5571
rect 23120 5537 23158 5571
rect 23192 5537 23230 5571
rect 23264 5537 23302 5571
rect 23336 5537 23374 5571
rect 23408 5537 23446 5571
rect 23480 5537 23486 5571
rect 22716 5498 23486 5537
tri 23801 5510 23943 5652 ne
rect 22716 5464 22798 5498
rect 22832 5464 22870 5498
rect 22904 5464 22942 5498
rect 22976 5464 23014 5498
rect 23048 5464 23086 5498
rect 23120 5464 23158 5498
rect 23192 5464 23230 5498
rect 23264 5464 23302 5498
rect 23336 5464 23374 5498
rect 23408 5464 23446 5498
rect 23480 5464 23486 5498
rect 22716 5427 23486 5464
tri 23486 5427 23487 5428 sw
rect 17481 5375 17487 5427
rect 17539 5375 17551 5427
rect 17603 5375 17609 5427
rect 20508 5375 20514 5427
rect 20566 5375 20578 5427
rect 20630 5375 20636 5427
rect 22716 5425 23487 5427
rect 22716 5391 22798 5425
rect 22832 5391 22870 5425
rect 22904 5391 22942 5425
rect 22976 5391 23014 5425
rect 23048 5391 23086 5425
rect 23120 5391 23158 5425
rect 23192 5391 23230 5425
rect 23264 5391 23302 5425
rect 23336 5391 23374 5425
rect 23408 5391 23446 5425
rect 23480 5391 23487 5425
rect 22716 5375 23487 5391
tri 23487 5375 23539 5427 sw
rect 22716 5352 23539 5375
rect 22716 5318 22798 5352
rect 22832 5318 22870 5352
rect 22904 5318 22942 5352
rect 22976 5318 23014 5352
rect 23048 5318 23086 5352
rect 23120 5318 23158 5352
rect 23192 5318 23230 5352
rect 23264 5318 23302 5352
rect 23336 5318 23374 5352
rect 23408 5318 23446 5352
rect 23480 5318 23539 5352
rect 22716 5286 23539 5318
tri 23539 5286 23628 5375 sw
rect 12413 5232 12419 5284
rect 12471 5232 12490 5284
rect 12542 5232 12561 5284
rect 12613 5232 12632 5284
rect 12684 5232 12703 5284
rect 12755 5232 12773 5284
rect 12825 5232 12831 5284
rect 22716 5280 23802 5286
rect 22716 5275 22782 5280
tri 16546 5246 16551 5251 se
rect 16551 5246 16603 5251
tri 16540 5240 16546 5246 se
rect 16546 5245 16603 5246
rect 16546 5240 16551 5245
rect 12413 5220 12831 5232
tri 16521 5221 16540 5240 se
rect 16540 5221 16551 5240
rect 12413 5168 12419 5220
rect 12471 5168 12490 5220
rect 12542 5168 12561 5220
rect 12613 5168 12632 5220
rect 12684 5168 12703 5220
rect 12755 5168 12773 5220
rect 12825 5168 12831 5220
tri 16454 5208 16467 5221 se
rect 16467 5208 16551 5221
tri 16420 5174 16454 5208 se
rect 16454 5193 16551 5208
rect 16454 5178 16603 5193
rect 16454 5174 16551 5178
tri 16414 5168 16420 5174 se
rect 16420 5168 16551 5174
tri 16413 5167 16414 5168 se
rect 16414 5167 16551 5168
tri 16382 5136 16413 5167 se
rect 16413 5136 16551 5167
tri 16366 5120 16382 5136 se
rect 16382 5126 16551 5136
rect 16382 5120 16603 5126
rect 16874 5246 16926 5248
tri 16926 5246 16928 5248 sw
rect 22740 5246 22782 5275
rect 22816 5246 22855 5280
rect 22889 5246 22928 5280
rect 22962 5246 23001 5280
rect 23035 5246 23074 5280
rect 23108 5246 23147 5280
rect 23181 5246 23220 5280
rect 23254 5246 23294 5280
rect 23328 5246 23368 5280
rect 23402 5246 23442 5280
rect 23476 5246 23516 5280
rect 23550 5274 23802 5280
rect 23550 5246 23593 5274
rect 16874 5242 16928 5246
rect 16926 5240 16928 5242
tri 16928 5240 16934 5246 sw
rect 22740 5240 23593 5246
rect 23627 5240 23665 5274
rect 23699 5240 23737 5274
rect 23771 5240 23802 5274
rect 16926 5211 16934 5240
tri 16934 5211 16963 5240 sw
rect 16926 5208 17095 5211
tri 17095 5208 17098 5211 sw
rect 22740 5208 23802 5240
rect 16926 5190 17098 5208
rect 16874 5178 17098 5190
rect 16926 5174 17098 5178
tri 17098 5174 17132 5208 sw
rect 22740 5174 22782 5208
rect 22816 5174 22855 5208
rect 22889 5174 22928 5208
rect 22962 5174 23001 5208
rect 23035 5174 23074 5208
rect 23108 5174 23147 5208
rect 23181 5174 23220 5208
rect 23254 5174 23294 5208
rect 23328 5174 23368 5208
rect 23402 5174 23442 5208
rect 23476 5174 23516 5208
rect 23550 5201 23802 5208
rect 23550 5174 23593 5201
rect 16926 5167 17132 5174
tri 17132 5167 17139 5174 sw
rect 22740 5167 23593 5174
rect 23627 5167 23665 5201
rect 23699 5167 23737 5201
rect 23771 5167 23802 5201
rect 16926 5144 17139 5167
tri 17139 5144 17162 5167 sw
rect 16926 5130 20336 5144
rect 16926 5126 20214 5130
rect 16874 5120 20214 5126
tri 16348 5102 16366 5120 se
rect 16366 5102 16472 5120
tri 16472 5102 16490 5120 nw
tri 17048 5102 17066 5120 ne
rect 17066 5102 20214 5120
tri 16343 5097 16348 5102 se
rect 16348 5097 16467 5102
tri 16467 5097 16472 5102 nw
tri 17066 5097 17071 5102 ne
rect 17071 5097 20214 5102
tri 16340 5094 16343 5097 se
rect 16343 5094 16464 5097
tri 16464 5094 16467 5097 nw
tri 17071 5094 17074 5097 ne
rect 17074 5094 20214 5097
tri 16324 5078 16340 5094 se
rect 16340 5078 16448 5094
tri 16448 5078 16464 5094 nw
tri 17074 5078 17090 5094 ne
rect 17090 5078 20214 5094
rect 20266 5078 20278 5130
rect 20330 5078 20336 5130
tri 16313 5067 16324 5078 se
rect 16324 5067 16434 5078
rect 14217 5064 16434 5067
tri 16434 5064 16448 5078 nw
tri 17090 5064 17104 5078 ne
rect 17104 5064 20336 5078
rect 22740 5136 23802 5167
rect 22740 5102 22782 5136
rect 22816 5102 22855 5136
rect 22889 5102 22928 5136
rect 22962 5102 23001 5136
rect 23035 5102 23074 5136
rect 23108 5102 23147 5136
rect 23181 5102 23220 5136
rect 23254 5102 23294 5136
rect 23328 5102 23368 5136
rect 23402 5102 23442 5136
rect 23476 5102 23516 5136
rect 23550 5128 23802 5136
rect 23550 5102 23593 5128
rect 22740 5094 23593 5102
rect 23627 5094 23665 5128
rect 23699 5094 23737 5128
rect 23771 5094 23802 5128
rect 22740 5064 23802 5094
rect 14217 5044 16407 5064
rect 14217 4992 14223 5044
rect 14275 4992 14290 5044
rect 14342 5037 16407 5044
tri 16407 5037 16434 5064 nw
rect 14342 5030 16400 5037
tri 16400 5030 16407 5037 nw
rect 14342 5029 16399 5030
tri 16399 5029 16400 5030 nw
rect 14342 5021 16391 5029
tri 16391 5021 16399 5029 nw
rect 14342 4992 16362 5021
tri 16362 4992 16391 5021 nw
rect 14217 4969 16339 4992
tri 16339 4969 16362 4992 nw
rect 16926 4985 16932 5037
rect 16984 4985 16996 5037
rect 17048 5030 17054 5037
tri 17054 5030 17061 5037 sw
rect 22740 5030 22782 5064
rect 22816 5030 22855 5064
rect 22889 5030 22928 5064
rect 22962 5030 23001 5064
rect 23035 5030 23074 5064
rect 23108 5030 23147 5064
rect 23181 5030 23220 5064
rect 23254 5030 23294 5064
rect 23328 5030 23368 5064
rect 23402 5030 23442 5064
rect 23476 5030 23516 5064
rect 23550 5055 23802 5064
rect 23550 5030 23593 5055
rect 17048 5029 17061 5030
tri 17061 5029 17062 5030 sw
rect 17048 5025 20336 5029
rect 17048 4985 20214 5025
tri 17038 4969 17054 4985 ne
rect 17054 4973 20214 4985
rect 20266 4973 20278 5025
rect 20330 4973 20336 5025
rect 17054 4969 20336 4973
rect 22740 5021 23593 5030
rect 23627 5021 23665 5055
rect 23699 5021 23737 5055
rect 23771 5021 23802 5055
rect 22740 4992 23802 5021
rect 14217 4967 16337 4969
tri 16337 4967 16339 4969 nw
tri 16682 4915 16707 4940 se
rect 16707 4915 16792 4968
rect 22740 4958 22782 4992
rect 22816 4958 22855 4992
rect 22889 4958 22928 4992
rect 22962 4958 23001 4992
rect 23035 4958 23074 4992
rect 23108 4958 23147 4992
rect 23181 4958 23220 4992
rect 23254 4958 23294 4992
rect 23328 4958 23368 4992
rect 23402 4958 23442 4992
rect 23476 4958 23516 4992
rect 23550 4982 23802 4992
rect 23550 4958 23593 4982
rect 22740 4952 23593 4958
rect 22740 4948 22878 4952
tri 22878 4948 22882 4952 nw
tri 23420 4948 23424 4952 ne
rect 23424 4948 23593 4952
rect 23627 4948 23665 4982
rect 23699 4948 23737 4982
rect 23771 4948 23802 4982
rect 22740 4915 22845 4948
tri 22845 4915 22878 4948 nw
tri 23424 4915 23457 4948 ne
rect 23457 4915 23802 4948
rect 697 4791 865 4858
rect 14430 4797 16900 4915
rect 22740 4909 22839 4915
tri 22839 4909 22845 4915 nw
tri 23457 4909 23463 4915 ne
rect 23463 4909 23802 4915
rect 22740 4905 22835 4909
tri 22835 4905 22839 4909 nw
tri 23463 4905 23467 4909 ne
rect 23467 4905 23593 4909
rect 22198 4819 22571 4905
rect 22740 4875 22805 4905
tri 22805 4875 22835 4905 nw
tri 23467 4875 23497 4905 ne
rect 23497 4875 23593 4905
rect 23627 4875 23665 4909
rect 23699 4875 23737 4909
rect 23771 4875 23802 4909
rect 22740 4836 22766 4875
tri 22766 4836 22805 4875 nw
tri 23497 4836 23536 4875 ne
rect 23536 4836 23802 4875
rect 22740 4819 22749 4836
tri 22749 4819 22766 4836 nw
tri 23536 4819 23553 4836 ne
rect 23553 4819 23593 4836
tri 22740 4810 22749 4819 nw
tri 23553 4810 23562 4819 ne
rect 23562 4802 23593 4819
rect 23627 4802 23665 4836
rect 23699 4802 23737 4836
rect 23771 4802 23802 4836
tri 697 4766 722 4791 ne
rect 722 4746 840 4791
tri 840 4766 865 4791 nw
rect 722 4712 728 4746
rect 762 4712 800 4746
rect 834 4712 840 4746
rect 722 4673 840 4712
rect 23562 4763 23802 4802
rect 23562 4729 23593 4763
rect 23627 4729 23665 4763
rect 23699 4729 23737 4763
rect 23771 4729 23802 4763
rect 722 4639 728 4673
rect 762 4672 840 4673
rect 762 4639 800 4672
rect 722 4638 800 4639
rect 834 4638 840 4672
rect 722 4600 840 4638
rect 13292 4676 14489 4700
rect 13292 4624 13322 4676
rect 13374 4624 13389 4676
rect 13441 4624 14200 4676
rect 14252 4624 14267 4676
rect 14319 4624 14489 4676
rect 13292 4600 14489 4624
rect 23562 4690 23802 4729
rect 23562 4656 23593 4690
rect 23627 4656 23665 4690
rect 23699 4656 23737 4690
rect 23771 4656 23802 4690
rect 23562 4617 23802 4656
rect 722 4566 728 4600
rect 762 4598 840 4600
rect 762 4566 800 4598
rect 722 4564 800 4566
rect 834 4564 840 4598
rect 722 4527 840 4564
rect 23562 4583 23593 4617
rect 23627 4583 23665 4617
rect 23699 4583 23737 4617
rect 23771 4583 23802 4617
rect 722 4493 728 4527
rect 762 4524 840 4527
rect 762 4493 800 4524
rect 258 4479 422 4491
rect 258 4373 310 4479
tri 279 4348 304 4373 ne
rect 304 2573 310 4373
rect 416 2573 422 4479
rect 304 2534 422 2573
rect 304 2500 310 2534
rect 344 2500 382 2534
rect 416 2500 422 2534
rect 304 2461 422 2500
rect 304 2427 310 2461
rect 344 2427 382 2461
rect 416 2427 422 2461
rect 304 2388 422 2427
rect 304 2354 310 2388
rect 344 2354 382 2388
rect 416 2354 422 2388
rect 304 2315 422 2354
rect 304 2281 310 2315
rect 344 2281 382 2315
rect 416 2281 422 2315
rect 304 2242 422 2281
rect 304 2208 310 2242
rect 344 2208 382 2242
rect 416 2208 422 2242
rect 304 2169 422 2208
rect 304 2135 310 2169
rect 344 2135 382 2169
rect 416 2135 422 2169
rect 304 2096 422 2135
rect 304 2062 310 2096
rect 344 2062 382 2096
rect 416 2062 422 2096
rect 304 2023 422 2062
rect 304 1989 310 2023
rect 344 1989 382 2023
rect 416 1989 422 2023
rect 304 1950 422 1989
rect 304 1916 310 1950
rect 344 1916 382 1950
rect 416 1916 422 1950
rect 304 1877 422 1916
rect 304 1843 310 1877
rect 344 1843 382 1877
rect 416 1843 422 1877
rect 304 1804 422 1843
rect 304 1770 310 1804
rect 344 1770 382 1804
rect 416 1770 422 1804
rect 304 1731 422 1770
rect 304 1697 310 1731
rect 344 1697 382 1731
rect 416 1697 422 1731
rect 304 1658 422 1697
rect 304 1624 310 1658
rect 344 1624 382 1658
rect 416 1624 422 1658
rect 304 1585 422 1624
rect 304 1551 310 1585
rect 344 1551 382 1585
rect 416 1551 422 1585
rect 304 1512 422 1551
rect 304 1478 310 1512
rect 344 1478 382 1512
rect 416 1478 422 1512
rect 304 1439 422 1478
rect 304 1405 310 1439
rect 344 1405 382 1439
rect 416 1405 422 1439
rect 304 1366 422 1405
rect 304 1332 310 1366
rect 344 1332 382 1366
rect 416 1332 422 1366
rect 304 1293 422 1332
rect 304 1259 310 1293
rect 344 1259 382 1293
rect 416 1259 422 1293
rect 304 1220 422 1259
rect 304 1186 310 1220
rect 344 1186 382 1220
rect 416 1186 422 1220
rect 304 1147 422 1186
rect 304 1113 310 1147
rect 344 1113 382 1147
rect 416 1113 422 1147
rect 304 1074 422 1113
rect 304 1040 310 1074
rect 344 1040 382 1074
rect 416 1040 422 1074
rect 304 1001 422 1040
rect 304 967 310 1001
rect 344 967 382 1001
rect 416 967 422 1001
rect 304 928 422 967
rect 304 894 310 928
rect 344 894 382 928
rect 416 894 422 928
rect 304 855 422 894
rect 722 4490 800 4493
rect 834 4490 840 4524
tri 10896 4510 10902 4516 se
tri 10894 4508 10896 4510 se
rect 10896 4508 10902 4510
tri 10877 4491 10894 4508 se
rect 10894 4491 10902 4508
rect 722 4454 840 4490
rect 722 4420 728 4454
rect 762 4450 840 4454
rect 762 4420 800 4450
rect 722 4416 800 4420
rect 834 4416 840 4450
rect 722 4381 840 4416
rect 722 4347 728 4381
rect 762 4376 840 4381
rect 762 4347 800 4376
rect 722 4342 800 4347
rect 834 4342 840 4376
rect 722 4308 840 4342
rect 722 4274 728 4308
rect 762 4302 840 4308
rect 762 4274 800 4302
rect 722 4268 800 4274
rect 834 4268 840 4302
rect 722 4235 840 4268
rect 722 4201 728 4235
rect 762 4228 840 4235
rect 762 4201 800 4228
rect 722 4194 800 4201
rect 834 4194 840 4228
rect 722 4162 840 4194
rect 722 4128 728 4162
rect 762 4154 840 4162
rect 762 4128 800 4154
rect 722 4120 800 4128
rect 834 4120 840 4154
rect 722 4089 840 4120
rect 722 4055 728 4089
rect 762 4080 840 4089
rect 762 4055 800 4080
rect 722 4046 800 4055
rect 834 4046 840 4080
rect 722 4016 840 4046
rect 722 3982 728 4016
rect 762 4006 840 4016
rect 762 3982 800 4006
rect 722 3972 800 3982
rect 834 3972 840 4006
rect 722 3943 840 3972
rect 722 3909 728 3943
rect 762 3932 840 3943
rect 762 3909 800 3932
rect 722 3898 800 3909
rect 834 3898 840 3932
rect 722 3870 840 3898
rect 722 3836 728 3870
rect 762 3858 840 3870
rect 762 3836 800 3858
rect 722 3824 800 3836
rect 834 3824 840 3858
rect 722 3797 840 3824
rect 722 3763 728 3797
rect 762 3784 840 3797
rect 762 3763 800 3784
rect 722 3750 800 3763
rect 834 3750 840 3784
rect 722 3724 840 3750
rect 722 3690 728 3724
rect 762 3710 840 3724
rect 762 3690 800 3710
rect 722 3676 800 3690
rect 834 3676 840 3710
rect 722 3651 840 3676
rect 722 3617 728 3651
rect 762 3636 840 3651
rect 762 3617 800 3636
rect 722 3602 800 3617
rect 834 3602 840 3636
rect 722 3578 840 3602
rect 722 3544 728 3578
rect 762 3562 840 3578
rect 762 3544 800 3562
rect 722 3528 800 3544
rect 834 3528 840 3562
rect 722 3505 840 3528
rect 722 3471 728 3505
rect 762 3488 840 3505
rect 762 3471 800 3488
rect 722 3454 800 3471
rect 834 3454 840 3488
rect 722 3432 840 3454
rect 722 3398 728 3432
rect 762 3414 840 3432
rect 762 3398 800 3414
rect 722 3380 800 3398
rect 834 3380 840 3414
rect 722 3359 840 3380
rect 722 3325 728 3359
rect 762 3341 840 3359
rect 762 3325 800 3341
rect 722 3307 800 3325
rect 834 3307 840 3341
rect 722 3286 840 3307
rect 722 3252 728 3286
rect 762 3268 840 3286
rect 762 3252 800 3268
rect 722 3234 800 3252
rect 834 3234 840 3268
rect 722 3213 840 3234
rect 722 3179 728 3213
rect 762 3195 840 3213
rect 762 3179 800 3195
rect 722 3161 800 3179
rect 834 3161 840 3195
rect 722 3140 840 3161
rect 722 3106 728 3140
rect 762 3122 840 3140
rect 762 3106 800 3122
rect 722 3088 800 3106
rect 834 3088 840 3122
rect 722 3067 840 3088
rect 722 3033 728 3067
rect 762 3049 840 3067
rect 762 3033 800 3049
rect 722 3015 800 3033
rect 834 3015 840 3049
rect 722 2994 840 3015
rect 722 2960 728 2994
rect 762 2976 840 2994
rect 762 2960 800 2976
rect 722 2942 800 2960
rect 834 2942 840 2976
rect 722 2921 840 2942
rect 722 2887 728 2921
rect 762 2903 840 2921
rect 762 2887 800 2903
rect 722 2869 800 2887
rect 834 2869 840 2903
rect 722 2848 840 2869
rect 722 2814 728 2848
rect 762 2830 840 2848
rect 762 2814 800 2830
rect 722 2796 800 2814
rect 834 2796 840 2830
rect 722 2775 840 2796
rect 722 2741 728 2775
rect 762 2757 840 2775
rect 762 2741 800 2757
rect 722 2723 800 2741
rect 834 2723 840 2757
rect 722 2702 840 2723
rect 722 2668 728 2702
rect 762 2684 840 2702
rect 762 2668 800 2684
rect 722 2650 800 2668
rect 834 2650 840 2684
rect 722 2629 840 2650
rect 722 2595 728 2629
rect 762 2611 840 2629
rect 762 2595 800 2611
rect 722 2577 800 2595
rect 834 2577 840 2611
rect 722 2556 840 2577
rect 722 2522 728 2556
rect 762 2538 840 2556
rect 762 2522 800 2538
rect 722 2504 800 2522
rect 834 2504 840 2538
rect 722 2483 840 2504
rect 722 2449 728 2483
rect 762 2465 840 2483
rect 762 2449 800 2465
rect 722 2431 800 2449
rect 834 2431 840 2465
rect 722 2411 840 2431
rect 722 2377 728 2411
rect 762 2392 840 2411
rect 762 2377 800 2392
rect 722 2358 800 2377
rect 834 2358 840 2392
rect 722 2339 840 2358
rect 722 2305 728 2339
rect 762 2319 840 2339
rect 762 2305 800 2319
rect 722 2285 800 2305
rect 834 2285 840 2319
rect 722 2267 840 2285
rect 722 2233 728 2267
rect 762 2246 840 2267
rect 762 2233 800 2246
rect 722 2212 800 2233
rect 834 2212 840 2246
rect 722 2195 840 2212
rect 722 2161 728 2195
rect 762 2173 840 2195
rect 762 2161 800 2173
rect 722 2139 800 2161
rect 834 2139 840 2173
rect 722 2123 840 2139
rect 722 2089 728 2123
rect 762 2100 840 2123
rect 762 2089 800 2100
rect 722 2066 800 2089
rect 834 2066 840 2100
rect 722 2051 840 2066
rect 722 2017 728 2051
rect 762 2027 840 2051
rect 762 2017 800 2027
rect 722 1993 800 2017
rect 834 1993 840 2027
rect 722 1979 840 1993
rect 722 1945 728 1979
rect 762 1954 840 1979
rect 762 1945 800 1954
rect 722 1920 800 1945
rect 834 1920 840 1954
rect 722 1907 840 1920
rect 722 1873 728 1907
rect 762 1881 840 1907
rect 762 1873 800 1881
rect 722 1847 800 1873
rect 834 1847 840 1881
rect 722 1835 840 1847
rect 722 1801 728 1835
rect 762 1808 840 1835
rect 762 1801 800 1808
rect 722 1774 800 1801
rect 834 1774 840 1808
rect 722 1763 840 1774
rect 722 1729 728 1763
rect 762 1735 840 1763
rect 762 1729 800 1735
rect 722 1701 800 1729
rect 834 1701 840 1735
rect 722 1691 840 1701
rect 722 1657 728 1691
rect 762 1662 840 1691
rect 762 1657 800 1662
rect 722 1628 800 1657
rect 834 1628 840 1662
rect 722 1619 840 1628
rect 722 1585 728 1619
rect 762 1589 840 1619
rect 762 1585 800 1589
rect 722 1555 800 1585
rect 834 1555 840 1589
rect 722 1547 840 1555
rect 722 1513 728 1547
rect 762 1516 840 1547
rect 762 1513 800 1516
rect 722 1482 800 1513
rect 834 1482 840 1516
rect 722 1475 840 1482
rect 722 1441 728 1475
rect 762 1443 840 1475
rect 762 1441 800 1443
rect 722 1409 800 1441
rect 834 1409 840 1443
rect 722 1403 840 1409
rect 722 1369 728 1403
rect 762 1370 840 1403
rect 762 1369 800 1370
rect 722 1336 800 1369
rect 834 1336 840 1370
rect 1153 4485 10902 4491
rect 1153 4479 1687 4485
rect 1153 4445 1169 4479
rect 1203 4445 1241 4479
rect 1275 4445 1313 4479
rect 1347 4445 1385 4479
rect 1419 4445 1457 4479
rect 1491 4445 1529 4479
rect 1563 4445 1601 4479
rect 1635 4451 1687 4479
rect 1721 4451 1760 4485
rect 1794 4451 1833 4485
rect 1867 4451 1906 4485
rect 1940 4451 1979 4485
rect 2013 4451 2052 4485
rect 2086 4451 2125 4485
rect 2159 4451 2198 4485
rect 2232 4451 2271 4485
rect 2305 4451 2344 4485
rect 2378 4451 2417 4485
rect 2451 4451 2490 4485
rect 2524 4451 2562 4485
rect 2596 4451 2634 4485
rect 2668 4451 2706 4485
rect 2740 4451 2778 4485
rect 2812 4451 2850 4485
rect 2884 4451 2922 4485
rect 2956 4451 2994 4485
rect 3028 4451 3066 4485
rect 3100 4451 3138 4485
rect 3172 4451 3210 4485
rect 3244 4451 3282 4485
rect 3316 4451 3354 4485
rect 3388 4451 3426 4485
rect 3460 4451 3498 4485
rect 3532 4451 3570 4485
rect 3604 4451 3642 4485
rect 3676 4451 3714 4485
rect 3748 4451 3786 4485
rect 3820 4451 3858 4485
rect 3892 4451 3930 4485
rect 3964 4451 4002 4485
rect 4036 4451 4074 4485
rect 4108 4451 4146 4485
rect 4180 4451 4218 4485
rect 4252 4451 4290 4485
rect 4324 4451 4362 4485
rect 4396 4451 4434 4485
rect 4468 4451 4506 4485
rect 4540 4451 4578 4485
rect 4612 4451 4650 4485
rect 4684 4451 4722 4485
rect 4756 4451 4794 4485
rect 4828 4451 4866 4485
rect 4900 4451 4938 4485
rect 4972 4451 5010 4485
rect 5044 4451 5082 4485
rect 5116 4451 5154 4485
rect 5188 4451 5226 4485
rect 5260 4451 5298 4485
rect 5332 4451 5370 4485
rect 5404 4451 5442 4485
rect 5476 4451 5514 4485
rect 5548 4451 5586 4485
rect 5620 4451 5658 4485
rect 5692 4451 5730 4485
rect 5764 4451 5802 4485
rect 5836 4451 5874 4485
rect 5908 4451 5946 4485
rect 5980 4451 6018 4485
rect 6052 4451 6090 4485
rect 6124 4451 6162 4485
rect 6196 4451 6234 4485
rect 6268 4451 6306 4485
rect 6340 4451 6378 4485
rect 6412 4451 6450 4485
rect 6484 4451 6522 4485
rect 6556 4451 6594 4485
rect 6628 4451 6666 4485
rect 6700 4451 6738 4485
rect 6772 4451 6810 4485
rect 6844 4451 6882 4485
rect 6916 4451 6954 4485
rect 6988 4451 7026 4485
rect 7060 4451 7098 4485
rect 7132 4451 7170 4485
rect 7204 4451 7242 4485
rect 7276 4451 7314 4485
rect 7348 4451 7386 4485
rect 7420 4451 7458 4485
rect 7492 4451 7530 4485
rect 7564 4451 7602 4485
rect 7636 4451 7674 4485
rect 7708 4451 7746 4485
rect 7780 4451 7818 4485
rect 7852 4451 7890 4485
rect 7924 4451 7962 4485
rect 7996 4451 8034 4485
rect 8068 4451 8106 4485
rect 8140 4451 8178 4485
rect 8212 4451 8250 4485
rect 8284 4451 8322 4485
rect 8356 4451 8394 4485
rect 8428 4451 8466 4485
rect 8500 4451 8538 4485
rect 8572 4451 8610 4485
rect 8644 4451 8682 4485
rect 8716 4451 8754 4485
rect 8788 4451 8826 4485
rect 8860 4451 8898 4485
rect 8932 4451 8970 4485
rect 9004 4451 9042 4485
rect 9076 4451 9114 4485
rect 9148 4451 9186 4485
rect 9220 4451 9258 4485
rect 9292 4451 9330 4485
rect 9364 4451 9402 4485
rect 9436 4451 9474 4485
rect 9508 4451 9546 4485
rect 9580 4451 9618 4485
rect 9652 4451 9690 4485
rect 9724 4451 9762 4485
rect 9796 4451 9834 4485
rect 9868 4451 9906 4485
rect 9940 4451 9978 4485
rect 10012 4451 10050 4485
rect 10084 4451 10122 4485
rect 10156 4451 10194 4485
rect 10228 4451 10266 4485
rect 10300 4451 10338 4485
rect 10372 4451 10410 4485
rect 10444 4451 10482 4485
rect 10516 4451 10554 4485
rect 10588 4451 10626 4485
rect 10660 4451 10698 4485
rect 10732 4451 10770 4485
rect 10804 4451 10842 4485
rect 10876 4451 10902 4485
rect 1635 4445 10902 4451
rect 1153 4437 1785 4445
tri 1785 4437 1793 4445 nw
tri 10888 4437 10896 4445 ne
rect 10896 4437 10902 4445
rect 1153 4435 1783 4437
tri 1783 4435 1785 4437 nw
tri 10896 4435 10898 4437 ne
rect 10898 4435 10902 4437
rect 1153 4431 1779 4435
tri 1779 4431 1783 4435 nw
tri 10898 4431 10902 4435 ne
rect 12413 4495 12419 4547
rect 12471 4495 12490 4547
rect 12542 4495 12561 4547
rect 12613 4495 12632 4547
rect 12684 4495 12703 4547
rect 12755 4495 12773 4547
rect 12825 4495 12831 4547
rect 12413 4483 12831 4495
rect 12413 4431 12419 4483
rect 12471 4431 12490 4483
rect 12542 4431 12561 4483
rect 12613 4431 12632 4483
rect 12684 4431 12703 4483
rect 12755 4431 12773 4483
rect 12825 4431 12831 4483
rect 23562 4544 23802 4583
rect 23562 4510 23593 4544
rect 23627 4510 23665 4544
rect 23699 4510 23737 4544
rect 23771 4510 23802 4544
rect 23562 4471 23802 4510
rect 23562 4437 23593 4471
rect 23627 4437 23665 4471
rect 23699 4437 23737 4471
rect 23771 4437 23802 4471
rect 1153 4405 1746 4431
rect 1153 4371 1169 4405
rect 1203 4371 1241 4405
rect 1275 4371 1313 4405
rect 1347 4371 1385 4405
rect 1419 4371 1457 4405
rect 1491 4371 1529 4405
rect 1563 4371 1601 4405
rect 1635 4398 1746 4405
tri 1746 4398 1779 4431 nw
tri 11524 4398 11529 4403 se
rect 11529 4398 14462 4403
rect 1635 4385 1733 4398
tri 1733 4385 1746 4398 nw
tri 11511 4385 11524 4398 se
rect 11524 4385 14462 4398
rect 1635 4371 1712 4385
rect 1153 4364 1712 4371
tri 1712 4364 1733 4385 nw
tri 11490 4364 11511 4385 se
rect 11511 4364 14340 4385
rect 1153 4362 1710 4364
tri 1710 4362 1712 4364 nw
tri 11488 4362 11490 4364 se
rect 11490 4362 14340 4364
rect 1153 4331 1673 4362
rect 1153 4297 1169 4331
rect 1203 4297 1241 4331
rect 1275 4297 1313 4331
rect 1347 4297 1385 4331
rect 1419 4297 1457 4331
rect 1491 4297 1529 4331
rect 1563 4297 1601 4331
rect 1635 4325 1673 4331
tri 1673 4325 1710 4362 nw
tri 11451 4325 11488 4362 se
rect 11488 4325 14340 4362
rect 1635 4297 1651 4325
tri 1651 4303 1673 4325 nw
tri 11429 4303 11451 4325 se
rect 11451 4303 14340 4325
rect 1153 4257 1651 4297
tri 11417 4291 11429 4303 se
rect 11429 4291 14340 4303
tri 11415 4289 11417 4291 se
rect 11417 4289 14340 4291
tri 11395 4269 11415 4289 se
rect 11415 4269 14340 4289
rect 14456 4269 14462 4385
rect 23562 4398 23802 4437
rect 23562 4364 23593 4398
rect 23627 4364 23665 4398
rect 23699 4364 23737 4398
rect 23771 4364 23802 4398
rect 23562 4325 23802 4364
rect 23562 4291 23593 4325
rect 23627 4291 23665 4325
rect 23699 4291 23737 4325
rect 23771 4291 23802 4325
tri 11388 4262 11395 4269 se
rect 11395 4262 11578 4269
tri 11578 4262 11585 4269 nw
rect 19118 4264 23191 4270
tri 11383 4257 11388 4262 se
rect 11388 4257 11573 4262
tri 11573 4257 11578 4262 nw
rect 1153 4223 1169 4257
rect 1203 4223 1241 4257
rect 1275 4223 1313 4257
rect 1347 4223 1385 4257
rect 1419 4223 1457 4257
rect 1491 4223 1529 4257
rect 1563 4223 1601 4257
rect 1635 4223 1651 4257
tri 11382 4256 11383 4257 se
rect 11383 4256 11572 4257
tri 11572 4256 11573 4257 nw
rect 1153 4183 1651 4223
tri 11348 4222 11382 4256 se
rect 11382 4222 11538 4256
tri 11538 4222 11572 4256 nw
tri 11344 4218 11348 4222 se
rect 11348 4218 11534 4222
tri 11534 4218 11538 4222 nw
tri 11342 4216 11344 4218 se
rect 11344 4216 11532 4218
tri 11532 4216 11534 4218 nw
tri 11340 4214 11342 4216 se
rect 11342 4214 11530 4216
tri 11530 4214 11532 4216 nw
tri 11339 4213 11340 4214 se
rect 11340 4213 11529 4214
tri 11529 4213 11530 4214 nw
rect 1153 4149 1169 4183
rect 1203 4149 1241 4183
rect 1275 4149 1313 4183
rect 1347 4149 1385 4183
rect 1419 4149 1457 4183
rect 1491 4149 1529 4183
rect 1563 4149 1601 4183
rect 1635 4149 1651 4183
tri 11305 4179 11339 4213 se
rect 11339 4179 11495 4213
tri 11495 4179 11529 4213 nw
rect 1153 4109 1651 4149
tri 11271 4145 11305 4179 se
rect 11305 4145 11461 4179
tri 11461 4145 11495 4179 nw
rect 1153 4075 1169 4109
rect 1203 4075 1241 4109
rect 1275 4075 1313 4109
rect 1347 4075 1385 4109
rect 1419 4075 1457 4109
rect 1491 4075 1529 4109
rect 1563 4075 1601 4109
rect 1635 4075 1651 4109
rect 1153 4035 1651 4075
rect 1153 4001 1169 4035
rect 1203 4001 1241 4035
rect 1275 4001 1313 4035
rect 1347 4001 1385 4035
rect 1419 4001 1457 4035
rect 1491 4001 1529 4035
rect 1563 4001 1601 4035
rect 1635 4001 1651 4035
rect 1153 3962 1651 4001
rect 3310 4143 11459 4145
tri 11459 4143 11461 4145 nw
rect 3310 4139 11455 4143
tri 11455 4139 11459 4143 nw
rect 3310 4133 11422 4139
rect 3310 4060 5862 4133
rect 3310 4026 3946 4060
rect 3980 4026 4018 4060
rect 4052 4026 5862 4060
rect 3310 4017 5862 4026
rect 5978 4106 11422 4133
tri 11422 4106 11455 4139 nw
rect 5978 4072 11388 4106
tri 11388 4072 11422 4106 nw
rect 11889 4084 12423 4214
rect 16892 4210 16898 4262
rect 16950 4210 16962 4262
rect 17014 4256 17091 4262
rect 17014 4222 17045 4256
rect 17079 4222 17091 4256
rect 17014 4210 17091 4222
rect 19118 4257 22947 4264
rect 19118 4223 19124 4257
rect 19158 4223 19196 4257
rect 19230 4223 22947 4257
rect 19118 4212 22947 4223
rect 22999 4212 23011 4264
rect 23063 4212 23075 4264
rect 23127 4212 23139 4264
rect 19118 4206 23191 4212
rect 23562 4252 23802 4291
rect 23562 4218 23593 4252
rect 23627 4218 23665 4252
rect 23699 4218 23737 4252
rect 23771 4218 23802 4252
rect 23562 4179 23802 4218
rect 16700 4145 17609 4149
rect 16700 4093 17487 4145
rect 17539 4093 17551 4145
rect 17603 4093 17609 4145
rect 16700 4089 17609 4093
rect 23562 4145 23593 4179
rect 23627 4145 23665 4179
rect 23699 4145 23737 4179
rect 23771 4145 23802 4179
rect 23562 4106 23802 4145
rect 11889 4072 12411 4084
tri 12411 4072 12423 4084 nw
rect 23562 4072 23593 4106
rect 23627 4072 23665 4106
rect 23699 4072 23737 4106
rect 23771 4072 23802 4106
rect 5978 4070 11386 4072
tri 11386 4070 11388 4072 nw
rect 11889 4070 12409 4072
tri 12409 4070 12411 4072 nw
rect 5978 4059 11375 4070
tri 11375 4059 11386 4070 nw
rect 11889 4069 12408 4070
tri 12408 4069 12409 4070 nw
rect 11889 4059 12398 4069
tri 12398 4059 12408 4069 nw
rect 12582 4063 15763 4069
rect 5978 4017 11327 4059
rect 3310 4011 11327 4017
tri 11327 4011 11375 4059 nw
rect 11889 4011 12350 4059
tri 12350 4011 12398 4059 nw
rect 12582 4011 12592 4063
rect 12644 4059 12684 4063
rect 12736 4059 12775 4063
rect 12827 4059 15763 4063
rect 15580 4057 15763 4059
rect 3310 3986 3660 4011
tri 3710 3986 3735 4011 nw
tri 3985 3986 4010 4011 ne
tri 4140 3986 4165 4011 nw
tri 6759 3986 6784 4011 ne
rect 6784 3986 7184 4011
tri 7184 3986 7209 4011 nw
tri 7459 3986 7484 4011 ne
tri 7614 3986 7639 4011 nw
rect 1153 3928 1169 3962
rect 1203 3928 1241 3962
rect 1275 3928 1313 3962
rect 1347 3928 1385 3962
rect 1419 3928 1457 3962
rect 1491 3928 1529 3962
rect 1563 3928 1601 3962
rect 1635 3928 1651 3962
rect 1153 3889 1651 3928
rect 1153 3855 1169 3889
rect 1203 3855 1241 3889
rect 1275 3855 1313 3889
rect 1347 3855 1385 3889
rect 1419 3855 1457 3889
rect 1491 3855 1529 3889
rect 1563 3855 1601 3889
rect 1635 3855 1651 3889
rect 1153 3816 1651 3855
rect 1153 3782 1169 3816
rect 1203 3782 1241 3816
rect 1275 3782 1313 3816
rect 1347 3782 1385 3816
rect 1419 3782 1457 3816
rect 1491 3782 1529 3816
rect 1563 3782 1601 3816
rect 1635 3782 1651 3816
rect 1153 3743 1651 3782
rect 11889 3881 12220 4011
tri 12220 3881 12350 4011 nw
rect 12582 3999 12594 4011
rect 15580 4005 15705 4057
rect 15757 4005 15763 4057
rect 12582 3947 12592 3999
rect 15580 3993 15763 4005
rect 12582 3935 12594 3947
rect 15580 3941 15705 3993
rect 15757 3941 15763 3993
rect 12582 3883 12592 3935
rect 15580 3929 15763 3941
rect 12582 3881 12594 3883
rect 15580 3881 15705 3929
rect 11889 3853 12192 3881
tri 12192 3853 12220 3881 nw
rect 12582 3877 15705 3881
rect 15757 3877 15763 3929
rect 12582 3875 15763 3877
rect 23562 4033 23802 4072
rect 23562 3999 23593 4033
rect 23627 3999 23665 4033
rect 23699 3999 23737 4033
rect 23771 3999 23802 4033
rect 23562 3960 23802 3999
rect 23562 3926 23593 3960
rect 23627 3926 23665 3960
rect 23699 3926 23737 3960
rect 23771 3926 23802 3960
rect 23562 3887 23802 3926
rect 12582 3853 12666 3875
tri 12666 3853 12688 3875 nw
tri 12930 3853 12952 3875 ne
rect 12952 3853 13101 3875
tri 13101 3853 13123 3875 nw
tri 13365 3853 13387 3875 ne
rect 13387 3853 13536 3875
tri 13536 3853 13558 3875 nw
tri 13800 3853 13822 3875 ne
rect 13822 3853 13971 3875
tri 13971 3853 13993 3875 nw
tri 14235 3853 14257 3875 ne
rect 14257 3853 14406 3875
tri 14406 3853 14428 3875 nw
tri 14670 3853 14692 3875 ne
rect 14692 3853 14841 3875
tri 14841 3853 14863 3875 nw
rect 23562 3853 23593 3887
rect 23627 3853 23665 3887
rect 23699 3853 23737 3887
rect 23771 3853 23802 3887
rect 11889 3851 12190 3853
tri 12190 3851 12192 3853 nw
rect 12582 3851 12664 3853
tri 12664 3851 12666 3853 nw
tri 12952 3851 12954 3853 ne
rect 12954 3851 13099 3853
tri 13099 3851 13101 3853 nw
tri 13387 3851 13389 3853 ne
rect 13389 3851 13534 3853
tri 13534 3851 13536 3853 nw
tri 13822 3851 13824 3853 ne
rect 13824 3851 13969 3853
tri 13969 3851 13971 3853 nw
tri 14257 3851 14259 3853 ne
rect 14259 3851 14404 3853
tri 14404 3851 14406 3853 nw
tri 14692 3851 14694 3853 ne
rect 14694 3851 14839 3853
tri 14839 3851 14841 3853 nw
rect 11889 3814 12153 3851
tri 12153 3814 12190 3851 nw
rect 11889 3780 12119 3814
tri 12119 3780 12153 3814 nw
rect 12582 3780 12663 3851
tri 12663 3850 12664 3851 nw
tri 12954 3850 12955 3851 ne
tri 12663 3780 12683 3800 sw
tri 12935 3780 12955 3800 se
rect 12955 3780 13098 3851
tri 13098 3850 13099 3851 nw
tri 13389 3850 13390 3851 ne
tri 13098 3780 13118 3800 sw
tri 13370 3780 13390 3800 se
rect 13390 3780 13533 3851
tri 13533 3850 13534 3851 nw
tri 13824 3850 13825 3851 ne
tri 13533 3780 13553 3800 sw
tri 13805 3780 13825 3800 se
rect 13825 3780 13968 3851
tri 13968 3850 13969 3851 nw
tri 14259 3850 14260 3851 ne
tri 13968 3780 13988 3800 sw
tri 14240 3780 14260 3800 se
rect 14260 3780 14403 3851
tri 14403 3850 14404 3851 nw
tri 14694 3850 14695 3851 ne
tri 14403 3780 14423 3800 sw
tri 14675 3780 14695 3800 se
rect 14695 3780 14838 3851
tri 14838 3850 14839 3851 nw
rect 23562 3814 23802 3853
rect 19972 3802 20038 3808
tri 14838 3780 14858 3800 sw
rect 11889 3778 12117 3780
tri 12117 3778 12119 3780 nw
rect 12582 3778 12683 3780
tri 12683 3778 12685 3780 sw
tri 12933 3778 12935 3780 se
rect 12935 3778 13118 3780
tri 13118 3778 13120 3780 sw
tri 13368 3778 13370 3780 se
rect 13370 3778 13553 3780
tri 13553 3778 13555 3780 sw
tri 13803 3778 13805 3780 se
rect 13805 3778 13988 3780
tri 13988 3778 13990 3780 sw
tri 14238 3778 14240 3780 se
rect 14240 3778 14423 3780
tri 14423 3778 14425 3780 sw
tri 14673 3778 14675 3780 se
rect 14675 3778 14858 3780
tri 14858 3778 14860 3780 sw
rect 11889 3766 12105 3778
tri 12105 3766 12117 3778 nw
rect 12582 3775 12685 3778
tri 12685 3775 12688 3778 sw
tri 12930 3775 12933 3778 se
rect 12933 3775 13120 3778
tri 13120 3775 13123 3778 sw
tri 13365 3775 13368 3778 se
rect 13368 3775 13555 3778
tri 13555 3775 13558 3778 sw
tri 13800 3775 13803 3778 se
rect 13803 3775 13990 3778
tri 13990 3775 13993 3778 sw
tri 14235 3775 14238 3778 se
rect 14238 3775 14425 3778
tri 14425 3775 14428 3778 sw
tri 14670 3775 14673 3778 se
rect 14673 3775 14860 3778
tri 14860 3775 14863 3778 sw
rect 12582 3769 16439 3775
rect 1153 3709 1169 3743
rect 1203 3709 1241 3743
rect 1275 3709 1313 3743
rect 1347 3709 1385 3743
rect 1419 3709 1457 3743
rect 1491 3709 1529 3743
rect 1563 3709 1601 3743
rect 1635 3709 1651 3743
rect 12582 3765 15723 3769
rect 12582 3764 12594 3765
rect 12628 3764 12667 3765
rect 12701 3764 12740 3765
rect 12582 3712 12592 3764
rect 12644 3731 12667 3764
rect 12736 3731 12740 3764
rect 12774 3764 12813 3765
rect 12774 3731 12775 3764
rect 12847 3731 12886 3765
rect 12920 3731 12959 3765
rect 12993 3731 13032 3765
rect 13066 3731 13105 3765
rect 13139 3731 13178 3765
rect 13212 3731 13251 3765
rect 13285 3731 13324 3765
rect 13358 3731 13397 3765
rect 13431 3731 13470 3765
rect 13504 3731 13543 3765
rect 13577 3731 13616 3765
rect 13650 3731 13689 3765
rect 13723 3731 13762 3765
rect 13796 3731 13835 3765
rect 13869 3731 13908 3765
rect 13942 3731 13981 3765
rect 14015 3731 14054 3765
rect 14088 3731 14127 3765
rect 14161 3731 14200 3765
rect 14234 3731 14273 3765
rect 14307 3731 14346 3765
rect 14380 3731 14419 3765
rect 14453 3731 14492 3765
rect 14526 3731 14565 3765
rect 14599 3731 14638 3765
rect 14672 3731 14711 3765
rect 14745 3731 14784 3765
rect 14818 3731 14857 3765
rect 14891 3731 14930 3765
rect 14964 3731 15003 3765
rect 15037 3731 15076 3765
rect 15110 3731 15149 3765
rect 15183 3731 15222 3765
rect 15256 3731 15295 3765
rect 15329 3731 15368 3765
rect 15402 3731 15441 3765
rect 15475 3731 15514 3765
rect 15548 3731 15587 3765
rect 15621 3731 15660 3765
rect 15694 3731 15723 3765
rect 12644 3712 12684 3731
rect 12736 3712 12775 3731
rect 12827 3717 15723 3731
rect 15775 3717 15787 3769
rect 15839 3765 15851 3769
rect 15903 3765 15915 3769
rect 15967 3765 15979 3769
rect 16031 3765 16043 3769
rect 16095 3765 16107 3769
rect 15840 3731 15851 3765
rect 15913 3731 15915 3765
rect 16095 3731 16098 3765
rect 15839 3717 15851 3731
rect 15903 3717 15915 3731
rect 15967 3717 15979 3731
rect 16031 3717 16043 3731
rect 16095 3717 16107 3731
rect 16159 3717 16171 3769
rect 16223 3717 16235 3769
rect 16287 3717 16299 3769
rect 16351 3717 16363 3769
rect 16415 3765 16439 3769
rect 16424 3731 16439 3765
rect 16415 3717 16439 3731
rect 12827 3712 16439 3717
rect 1153 3670 1651 3709
rect 1153 3636 1169 3670
rect 1203 3636 1241 3670
rect 1275 3636 1313 3670
rect 1347 3636 1385 3670
rect 1419 3636 1457 3670
rect 1491 3636 1529 3670
rect 1563 3636 1601 3670
rect 1635 3636 1651 3670
rect 8812 3707 11515 3711
tri 11515 3707 11519 3711 sw
rect 8812 3705 11519 3707
tri 11519 3705 11521 3707 sw
rect 8812 3697 11521 3705
tri 11521 3697 11529 3705 sw
rect 12582 3704 16439 3712
rect 12582 3700 15723 3704
rect 8812 3693 11529 3697
tri 11529 3693 11533 3697 sw
rect 8812 3663 11533 3693
rect 1153 3597 1651 3636
rect 1153 3563 1169 3597
rect 1203 3563 1241 3597
rect 1275 3563 1313 3597
rect 1347 3563 1385 3597
rect 1419 3563 1457 3597
rect 1491 3563 1529 3597
rect 1563 3563 1601 3597
rect 1635 3563 1651 3597
rect 2098 3594 2104 3646
rect 2156 3594 2168 3646
rect 2220 3594 2232 3646
rect 2284 3594 2296 3646
rect 2348 3594 2360 3646
rect 2412 3594 2424 3646
rect 2476 3594 3010 3646
rect 5338 3594 5344 3646
rect 5396 3594 5408 3646
rect 5460 3594 5472 3646
rect 5524 3594 6484 3646
rect 8812 3629 8824 3663
rect 8858 3629 8898 3663
rect 8932 3629 8972 3663
rect 9006 3629 9046 3663
rect 9080 3629 9120 3663
rect 9154 3629 9194 3663
rect 9228 3629 9268 3663
rect 9302 3629 9342 3663
rect 9376 3629 9416 3663
rect 9450 3629 9490 3663
rect 9524 3629 9564 3663
rect 9598 3629 9638 3663
rect 9672 3629 9712 3663
rect 9746 3629 9786 3663
rect 9820 3629 9860 3663
rect 9894 3629 9934 3663
rect 9968 3629 10008 3663
rect 10042 3629 10082 3663
rect 10116 3629 10156 3663
rect 10190 3629 10230 3663
rect 10264 3629 10304 3663
rect 10338 3629 10378 3663
rect 10412 3629 10452 3663
rect 10486 3629 10526 3663
rect 10560 3629 10600 3663
rect 10634 3629 10674 3663
rect 10708 3629 10748 3663
rect 10782 3629 10822 3663
rect 10856 3629 10896 3663
rect 10930 3629 10970 3663
rect 11004 3629 11043 3663
rect 11077 3629 11116 3663
rect 11150 3629 11189 3663
rect 11223 3629 11262 3663
rect 11296 3629 11335 3663
rect 11369 3629 11408 3663
rect 11442 3629 11481 3663
rect 11515 3659 11533 3663
tri 11533 3659 11567 3693 sw
rect 11515 3646 11567 3659
tri 11567 3646 11580 3659 sw
rect 12582 3648 12592 3700
rect 12644 3693 12684 3700
rect 12736 3693 12775 3700
rect 12827 3693 15723 3700
rect 12644 3659 12667 3693
rect 12736 3659 12740 3693
rect 12774 3659 12775 3693
rect 12847 3659 12886 3693
rect 12920 3659 12959 3693
rect 12993 3659 13032 3693
rect 13066 3659 13105 3693
rect 13139 3659 13178 3693
rect 13212 3659 13251 3693
rect 13285 3659 13324 3693
rect 13358 3659 13397 3693
rect 13431 3659 13470 3693
rect 13504 3659 13543 3693
rect 13577 3659 13616 3693
rect 13650 3659 13689 3693
rect 13723 3659 13762 3693
rect 13796 3659 13835 3693
rect 13869 3659 13908 3693
rect 13942 3659 13981 3693
rect 14015 3659 14054 3693
rect 14088 3659 14127 3693
rect 14161 3659 14200 3693
rect 14234 3659 14273 3693
rect 14307 3659 14346 3693
rect 14380 3659 14419 3693
rect 14453 3659 14492 3693
rect 14526 3659 14565 3693
rect 14599 3659 14638 3693
rect 14672 3659 14711 3693
rect 14745 3659 14784 3693
rect 14818 3659 14857 3693
rect 14891 3659 14930 3693
rect 14964 3659 15003 3693
rect 15037 3659 15076 3693
rect 15110 3659 15149 3693
rect 15183 3659 15222 3693
rect 15256 3659 15295 3693
rect 15329 3659 15368 3693
rect 15402 3659 15441 3693
rect 15475 3659 15514 3693
rect 15548 3659 15587 3693
rect 15621 3659 15660 3693
rect 15694 3659 15723 3693
rect 12644 3648 12684 3659
rect 12736 3648 12775 3659
rect 12827 3652 15723 3659
rect 15775 3652 15787 3704
rect 15839 3693 15851 3704
rect 15903 3693 15915 3704
rect 15967 3693 15979 3704
rect 16031 3693 16043 3704
rect 16095 3693 16107 3704
rect 15840 3659 15851 3693
rect 15913 3659 15915 3693
rect 16095 3659 16098 3693
rect 15839 3652 15851 3659
rect 15903 3652 15915 3659
rect 15967 3652 15979 3659
rect 16031 3652 16043 3659
rect 16095 3652 16107 3659
rect 16159 3652 16171 3704
rect 16223 3652 16235 3704
rect 16287 3652 16299 3704
rect 16351 3652 16363 3704
rect 16415 3693 16439 3704
rect 16424 3659 16439 3693
rect 16415 3652 16439 3659
rect 12827 3648 16439 3652
rect 11515 3634 11580 3646
tri 11580 3634 11592 3646 sw
rect 12582 3639 16439 3648
rect 12582 3636 15723 3639
rect 11515 3632 11592 3634
tri 11592 3632 11594 3634 sw
rect 11515 3629 11594 3632
rect 8812 3621 11594 3629
tri 11594 3621 11605 3632 sw
rect 8812 3594 11605 3621
tri 11605 3594 11632 3621 sw
rect 1153 3524 1651 3563
rect 1153 3490 1169 3524
rect 1203 3490 1241 3524
rect 1275 3490 1313 3524
rect 1347 3490 1385 3524
rect 1419 3490 1457 3524
rect 1491 3490 1529 3524
rect 1563 3490 1601 3524
rect 1635 3490 1651 3524
rect 1153 3451 1651 3490
rect 1153 3417 1169 3451
rect 1203 3417 1241 3451
rect 1275 3417 1313 3451
rect 1347 3417 1385 3451
rect 1419 3417 1457 3451
rect 1491 3417 1529 3451
rect 1563 3417 1601 3451
rect 1635 3417 1651 3451
rect 1153 3378 1651 3417
rect 1153 3344 1169 3378
rect 1203 3344 1241 3378
rect 1275 3344 1313 3378
rect 1347 3344 1385 3378
rect 1419 3344 1457 3378
rect 1491 3344 1529 3378
rect 1563 3344 1601 3378
rect 1635 3375 1651 3378
rect 8812 3591 11632 3594
rect 8812 3557 8824 3591
rect 8858 3557 8898 3591
rect 8932 3557 8972 3591
rect 9006 3557 9046 3591
rect 9080 3557 9120 3591
rect 9154 3557 9194 3591
rect 9228 3557 9268 3591
rect 9302 3557 9342 3591
rect 9376 3557 9416 3591
rect 9450 3557 9490 3591
rect 9524 3557 9564 3591
rect 9598 3557 9638 3591
rect 9672 3557 9712 3591
rect 9746 3557 9786 3591
rect 9820 3557 9860 3591
rect 9894 3557 9934 3591
rect 9968 3557 10008 3591
rect 10042 3557 10082 3591
rect 10116 3557 10156 3591
rect 10190 3557 10230 3591
rect 10264 3557 10304 3591
rect 10338 3557 10378 3591
rect 10412 3557 10452 3591
rect 10486 3557 10526 3591
rect 10560 3557 10600 3591
rect 10634 3557 10674 3591
rect 10708 3557 10748 3591
rect 10782 3557 10822 3591
rect 10856 3557 10896 3591
rect 10930 3557 10970 3591
rect 11004 3557 11043 3591
rect 11077 3557 11116 3591
rect 11150 3557 11189 3591
rect 11223 3557 11262 3591
rect 11296 3557 11335 3591
rect 11369 3557 11408 3591
rect 11442 3557 11481 3591
rect 11515 3587 11632 3591
tri 11632 3587 11639 3594 sw
rect 11515 3581 11639 3587
tri 11639 3581 11645 3587 sw
rect 12582 3584 12592 3636
rect 12644 3621 12684 3636
rect 12736 3621 12775 3636
rect 12827 3621 15723 3636
rect 12644 3587 12667 3621
rect 12736 3587 12740 3621
rect 12774 3587 12775 3621
rect 12847 3587 12886 3621
rect 12920 3587 12959 3621
rect 12993 3587 13032 3621
rect 13066 3587 13105 3621
rect 13139 3587 13178 3621
rect 13212 3587 13251 3621
rect 13285 3587 13324 3621
rect 13358 3587 13397 3621
rect 13431 3587 13470 3621
rect 13504 3587 13543 3621
rect 13577 3587 13616 3621
rect 13650 3587 13689 3621
rect 13723 3587 13762 3621
rect 13796 3587 13835 3621
rect 13869 3587 13908 3621
rect 13942 3587 13981 3621
rect 14015 3587 14054 3621
rect 14088 3587 14127 3621
rect 14161 3587 14200 3621
rect 14234 3587 14273 3621
rect 14307 3587 14346 3621
rect 14380 3587 14419 3621
rect 14453 3587 14492 3621
rect 14526 3587 14565 3621
rect 14599 3587 14638 3621
rect 14672 3587 14711 3621
rect 14745 3587 14784 3621
rect 14818 3587 14857 3621
rect 14891 3587 14930 3621
rect 14964 3587 15003 3621
rect 15037 3587 15076 3621
rect 15110 3587 15149 3621
rect 15183 3587 15222 3621
rect 15256 3587 15295 3621
rect 15329 3587 15368 3621
rect 15402 3587 15441 3621
rect 15475 3587 15514 3621
rect 15548 3587 15587 3621
rect 15621 3587 15660 3621
rect 15694 3587 15723 3621
rect 15775 3587 15787 3639
rect 15839 3621 15851 3639
rect 15903 3621 15915 3639
rect 15967 3621 15979 3639
rect 16031 3621 16043 3639
rect 16095 3621 16107 3639
rect 15840 3587 15851 3621
rect 15913 3587 15915 3621
rect 16095 3587 16098 3621
rect 16159 3587 16171 3639
rect 16223 3587 16235 3639
rect 16287 3587 16299 3639
rect 16351 3587 16363 3639
rect 16415 3621 16439 3639
rect 16424 3587 16439 3621
rect 12644 3584 12684 3587
rect 12736 3584 12775 3587
rect 12827 3584 16439 3587
rect 12582 3581 16439 3584
rect 19972 3750 19979 3802
rect 20031 3750 20038 3802
rect 19972 3737 20038 3750
rect 19972 3685 19979 3737
rect 20031 3685 20038 3737
rect 19972 3672 20038 3685
rect 19972 3620 19979 3672
rect 20031 3620 20038 3672
rect 19972 3607 20038 3620
rect 11515 3561 11645 3581
tri 11645 3561 11665 3581 sw
tri 12930 3561 12950 3581 ne
rect 12950 3561 13103 3581
tri 13103 3561 13123 3581 nw
tri 13365 3561 13385 3581 ne
rect 13385 3561 13538 3581
tri 13538 3561 13558 3581 nw
tri 13800 3561 13820 3581 ne
rect 13820 3561 13973 3581
tri 13973 3561 13993 3581 nw
tri 14235 3561 14255 3581 ne
rect 14255 3561 14408 3581
tri 14408 3561 14428 3581 nw
tri 14670 3561 14690 3581 ne
rect 14690 3561 14843 3581
tri 14843 3561 14863 3581 nw
rect 11515 3559 11665 3561
tri 11665 3559 11667 3561 sw
tri 12950 3559 12952 3561 ne
rect 12952 3559 13101 3561
tri 13101 3559 13103 3561 nw
tri 13385 3559 13387 3561 ne
rect 13387 3559 13536 3561
tri 13536 3559 13538 3561 nw
tri 13820 3559 13822 3561 ne
rect 13822 3559 13971 3561
tri 13971 3559 13973 3561 nw
tri 14255 3559 14257 3561 ne
rect 14257 3559 14406 3561
tri 14406 3559 14408 3561 nw
tri 14690 3559 14692 3561 ne
rect 14692 3559 14841 3561
tri 14841 3559 14843 3561 nw
rect 11515 3557 11667 3559
rect 8812 3556 11667 3557
tri 11667 3556 11670 3559 sw
tri 12952 3556 12955 3559 ne
rect 8812 3522 11670 3556
tri 11670 3522 11704 3556 sw
rect 8812 3519 11704 3522
rect 8812 3485 8824 3519
rect 8858 3485 8898 3519
rect 8932 3485 8972 3519
rect 9006 3485 9046 3519
rect 9080 3485 9120 3519
rect 9154 3485 9194 3519
rect 9228 3485 9268 3519
rect 9302 3485 9342 3519
rect 9376 3485 9416 3519
rect 9450 3485 9490 3519
rect 9524 3485 9564 3519
rect 9598 3485 9638 3519
rect 9672 3485 9712 3519
rect 9746 3485 9786 3519
rect 9820 3485 9860 3519
rect 9894 3485 9934 3519
rect 9968 3485 10008 3519
rect 10042 3485 10082 3519
rect 10116 3485 10156 3519
rect 10190 3485 10230 3519
rect 10264 3485 10304 3519
rect 10338 3485 10378 3519
rect 10412 3485 10452 3519
rect 10486 3485 10526 3519
rect 10560 3485 10600 3519
rect 10634 3485 10674 3519
rect 10708 3485 10748 3519
rect 10782 3485 10822 3519
rect 10856 3485 10896 3519
rect 10930 3485 10970 3519
rect 11004 3485 11043 3519
rect 11077 3485 11116 3519
rect 11150 3485 11189 3519
rect 11223 3485 11262 3519
rect 11296 3485 11335 3519
rect 11369 3485 11408 3519
rect 11442 3485 11481 3519
rect 11515 3506 11704 3519
tri 11704 3506 11720 3522 sw
rect 11515 3488 11720 3506
tri 11720 3488 11738 3506 sw
tri 12937 3488 12955 3506 se
rect 12955 3488 13098 3559
tri 13098 3556 13101 3559 nw
tri 13387 3556 13390 3559 ne
tri 13098 3488 13116 3506 sw
tri 13372 3488 13390 3506 se
rect 13390 3488 13533 3559
tri 13533 3556 13536 3559 nw
tri 13822 3556 13825 3559 ne
tri 13533 3488 13551 3506 sw
tri 13807 3488 13825 3506 se
rect 13825 3488 13968 3559
tri 13968 3556 13971 3559 nw
tri 14257 3556 14260 3559 ne
tri 13968 3488 13986 3506 sw
tri 14242 3488 14260 3506 se
rect 14260 3488 14403 3559
tri 14403 3556 14406 3559 nw
tri 14692 3556 14695 3559 ne
tri 14403 3488 14421 3506 sw
tri 14677 3488 14695 3506 se
rect 14695 3488 14838 3559
tri 14838 3556 14841 3559 nw
rect 19972 3555 19979 3607
rect 20031 3555 20038 3607
rect 19972 3542 20038 3555
tri 14838 3488 14856 3506 sw
rect 19972 3490 19979 3542
rect 20031 3490 20038 3542
rect 11515 3486 11738 3488
tri 11738 3486 11740 3488 sw
tri 12935 3486 12937 3488 se
rect 12937 3486 13116 3488
tri 13116 3486 13118 3488 sw
tri 13370 3486 13372 3488 se
rect 13372 3486 13551 3488
tri 13551 3486 13553 3488 sw
tri 13805 3486 13807 3488 se
rect 13807 3486 13986 3488
tri 13986 3486 13988 3488 sw
tri 14240 3486 14242 3488 se
rect 14242 3486 14421 3488
tri 14421 3486 14423 3488 sw
tri 14675 3486 14677 3488 se
rect 14677 3486 14856 3488
tri 14856 3486 14858 3488 sw
rect 11515 3485 11740 3486
rect 8812 3481 11740 3485
tri 11740 3481 11745 3486 sw
tri 12930 3481 12935 3486 se
rect 12935 3481 13118 3486
tri 13118 3481 13123 3486 sw
tri 13365 3481 13370 3486 se
rect 13370 3481 13553 3486
tri 13553 3481 13558 3486 sw
tri 13800 3481 13805 3486 se
rect 13805 3481 13988 3486
tri 13988 3481 13993 3486 sw
tri 14235 3481 14240 3486 se
rect 14240 3481 14423 3486
tri 14423 3481 14428 3486 sw
tri 14670 3481 14675 3486 se
rect 14675 3481 14858 3486
tri 14858 3481 14863 3486 sw
rect 8812 3475 16439 3481
rect 8812 3471 15723 3475
rect 8812 3468 12594 3471
rect 12628 3468 12667 3471
rect 12701 3468 12740 3471
rect 12774 3468 12813 3471
rect 8812 3447 12411 3468
rect 8812 3413 8824 3447
rect 8858 3413 8897 3447
rect 8931 3413 8970 3447
rect 9004 3413 9043 3447
rect 9077 3413 9116 3447
rect 9150 3413 9189 3447
rect 9223 3413 9262 3447
rect 9296 3413 9336 3447
rect 9370 3413 9410 3447
rect 9444 3413 9484 3447
rect 9518 3413 9558 3447
rect 9592 3413 9632 3447
rect 9666 3413 9706 3447
rect 9740 3413 9780 3447
rect 9814 3413 9854 3447
rect 9888 3413 9928 3447
rect 9962 3413 10002 3447
rect 10036 3413 10076 3447
rect 10110 3413 10150 3447
rect 10184 3413 10224 3447
rect 10258 3413 10298 3447
rect 10332 3413 10372 3447
rect 10406 3413 10446 3447
rect 10480 3413 10520 3447
rect 10554 3413 10594 3447
rect 10628 3413 10668 3447
rect 10702 3413 10742 3447
rect 10776 3413 10816 3447
rect 10850 3413 10890 3447
rect 10924 3413 10964 3447
rect 10998 3413 11038 3447
rect 11072 3413 11112 3447
rect 11146 3413 11186 3447
rect 11220 3413 11260 3447
rect 11294 3413 11334 3447
rect 11368 3413 11408 3447
rect 11442 3413 11482 3447
rect 11516 3413 11556 3447
rect 11590 3416 12411 3447
rect 12463 3416 12484 3468
rect 12536 3416 12556 3468
rect 12847 3437 12886 3471
rect 12920 3437 12959 3471
rect 12993 3437 13032 3471
rect 13066 3437 13105 3471
rect 13139 3437 13178 3471
rect 13212 3437 13251 3471
rect 13285 3437 13324 3471
rect 13358 3437 13397 3471
rect 13431 3437 13470 3471
rect 13504 3437 13543 3471
rect 13577 3437 13616 3471
rect 13650 3437 13689 3471
rect 13723 3437 13762 3471
rect 13796 3437 13835 3471
rect 13869 3437 13908 3471
rect 13942 3437 13981 3471
rect 14015 3437 14054 3471
rect 14088 3437 14127 3471
rect 14161 3437 14200 3471
rect 14234 3437 14273 3471
rect 14307 3437 14346 3471
rect 14380 3437 14419 3471
rect 14453 3437 14492 3471
rect 14526 3437 14565 3471
rect 14599 3437 14638 3471
rect 14672 3437 14711 3471
rect 14745 3437 14784 3471
rect 14818 3437 14857 3471
rect 14891 3437 14930 3471
rect 14964 3437 15003 3471
rect 15037 3437 15076 3471
rect 15110 3437 15149 3471
rect 15183 3437 15222 3471
rect 15256 3437 15295 3471
rect 15329 3437 15368 3471
rect 15402 3437 15441 3471
rect 15475 3437 15514 3471
rect 15548 3437 15587 3471
rect 15621 3437 15660 3471
rect 15694 3437 15723 3471
rect 12608 3416 12628 3437
rect 12680 3416 12700 3437
rect 12752 3416 12772 3437
rect 12824 3423 15723 3437
rect 15775 3423 15787 3475
rect 15839 3471 15851 3475
rect 15903 3471 15915 3475
rect 15967 3471 15979 3475
rect 16031 3471 16043 3475
rect 16095 3471 16107 3475
rect 15840 3437 15851 3471
rect 15913 3437 15915 3471
rect 16095 3437 16098 3471
rect 15839 3423 15851 3437
rect 15903 3423 15915 3437
rect 15967 3423 15979 3437
rect 16031 3423 16043 3437
rect 16095 3423 16107 3437
rect 16159 3423 16171 3475
rect 16223 3423 16235 3475
rect 16287 3423 16299 3475
rect 16351 3423 16363 3475
rect 16415 3471 16439 3475
rect 16424 3437 16439 3471
rect 16415 3423 16439 3437
rect 12824 3416 16439 3423
rect 11590 3413 16439 3416
rect 8812 3406 16439 3413
rect 8812 3404 15723 3406
tri 1651 3375 1652 3376 sw
rect 8812 3375 12411 3404
rect 1635 3344 1652 3375
rect 1153 3341 1652 3344
tri 1652 3341 1686 3375 sw
rect 8812 3341 8824 3375
rect 8858 3341 8897 3375
rect 8931 3341 8970 3375
rect 9004 3341 9043 3375
rect 9077 3341 9116 3375
rect 9150 3341 9189 3375
rect 9223 3341 9262 3375
rect 9296 3341 9336 3375
rect 9370 3341 9410 3375
rect 9444 3341 9484 3375
rect 9518 3341 9558 3375
rect 9592 3341 9632 3375
rect 9666 3341 9706 3375
rect 9740 3341 9780 3375
rect 9814 3341 9854 3375
rect 9888 3341 9928 3375
rect 9962 3341 10002 3375
rect 10036 3341 10076 3375
rect 10110 3341 10150 3375
rect 10184 3341 10224 3375
rect 10258 3341 10298 3375
rect 10332 3341 10372 3375
rect 10406 3341 10446 3375
rect 10480 3341 10520 3375
rect 10554 3341 10594 3375
rect 10628 3341 10668 3375
rect 10702 3341 10742 3375
rect 10776 3341 10816 3375
rect 10850 3341 10890 3375
rect 10924 3341 10964 3375
rect 10998 3341 11038 3375
rect 11072 3341 11112 3375
rect 11146 3341 11186 3375
rect 11220 3341 11260 3375
rect 11294 3341 11334 3375
rect 11368 3341 11408 3375
rect 11442 3341 11482 3375
rect 11516 3341 11556 3375
rect 11590 3352 12411 3375
rect 12463 3352 12484 3404
rect 12536 3352 12556 3404
rect 12608 3399 12628 3404
rect 12680 3399 12700 3404
rect 12752 3399 12772 3404
rect 12824 3399 15723 3404
rect 12847 3365 12886 3399
rect 12920 3365 12959 3399
rect 12993 3365 13032 3399
rect 13066 3365 13105 3399
rect 13139 3365 13178 3399
rect 13212 3365 13251 3399
rect 13285 3365 13324 3399
rect 13358 3365 13397 3399
rect 13431 3365 13470 3399
rect 13504 3365 13543 3399
rect 13577 3365 13616 3399
rect 13650 3365 13689 3399
rect 13723 3365 13762 3399
rect 13796 3365 13835 3399
rect 13869 3365 13908 3399
rect 13942 3365 13981 3399
rect 14015 3365 14054 3399
rect 14088 3365 14127 3399
rect 14161 3365 14200 3399
rect 14234 3365 14273 3399
rect 14307 3365 14346 3399
rect 14380 3365 14419 3399
rect 14453 3365 14492 3399
rect 14526 3365 14565 3399
rect 14599 3365 14638 3399
rect 14672 3365 14711 3399
rect 14745 3365 14784 3399
rect 14818 3365 14857 3399
rect 14891 3365 14930 3399
rect 14964 3365 15003 3399
rect 15037 3365 15076 3399
rect 15110 3365 15149 3399
rect 15183 3365 15222 3399
rect 15256 3365 15295 3399
rect 15329 3365 15368 3399
rect 15402 3365 15441 3399
rect 15475 3365 15514 3399
rect 15548 3365 15587 3399
rect 15621 3365 15660 3399
rect 15694 3365 15723 3399
rect 12608 3352 12628 3365
rect 12680 3352 12700 3365
rect 12752 3352 12772 3365
rect 12824 3354 15723 3365
rect 15775 3354 15787 3406
rect 15839 3399 15851 3406
rect 15903 3399 15915 3406
rect 15967 3399 15979 3406
rect 16031 3399 16043 3406
rect 16095 3399 16107 3406
rect 15840 3365 15851 3399
rect 15913 3365 15915 3399
rect 16095 3365 16098 3399
rect 15839 3354 15851 3365
rect 15903 3354 15915 3365
rect 15967 3354 15979 3365
rect 16031 3354 16043 3365
rect 16095 3354 16107 3365
rect 16159 3354 16171 3406
rect 16223 3354 16235 3406
rect 16287 3354 16299 3406
rect 16351 3354 16363 3406
rect 16415 3399 16439 3406
rect 16424 3365 16439 3399
rect 16415 3354 16439 3365
rect 12824 3352 16439 3354
rect 11590 3341 16439 3352
rect 1153 3340 1686 3341
tri 1686 3340 1687 3341 sw
rect 8812 3340 16439 3341
rect 1153 3327 1687 3340
tri 1687 3327 1700 3340 sw
rect 1153 3305 1700 3327
rect 1153 3271 1169 3305
rect 1203 3271 1241 3305
rect 1275 3271 1313 3305
rect 1347 3271 1385 3305
rect 1419 3271 1457 3305
rect 1491 3271 1529 3305
rect 1563 3271 1601 3305
rect 1635 3303 1700 3305
tri 1700 3303 1724 3327 sw
rect 8812 3303 12411 3340
rect 1635 3271 1724 3303
rect 1153 3269 1724 3271
tri 1724 3269 1758 3303 sw
rect 8812 3269 8824 3303
rect 8858 3269 8897 3303
rect 8931 3269 8970 3303
rect 9004 3269 9043 3303
rect 9077 3269 9116 3303
rect 9150 3269 9189 3303
rect 9223 3269 9262 3303
rect 9296 3269 9336 3303
rect 9370 3269 9410 3303
rect 9444 3269 9484 3303
rect 9518 3269 9558 3303
rect 9592 3269 9632 3303
rect 9666 3269 9706 3303
rect 9740 3269 9780 3303
rect 9814 3269 9854 3303
rect 9888 3269 9928 3303
rect 9962 3269 10002 3303
rect 10036 3269 10076 3303
rect 10110 3269 10150 3303
rect 10184 3269 10224 3303
rect 10258 3269 10298 3303
rect 10332 3269 10372 3303
rect 10406 3269 10446 3303
rect 10480 3269 10520 3303
rect 10554 3269 10594 3303
rect 10628 3269 10668 3303
rect 10702 3269 10742 3303
rect 10776 3269 10816 3303
rect 10850 3269 10890 3303
rect 10924 3269 10964 3303
rect 10998 3269 11038 3303
rect 11072 3269 11112 3303
rect 11146 3269 11186 3303
rect 11220 3269 11260 3303
rect 11294 3269 11334 3303
rect 11368 3269 11408 3303
rect 11442 3269 11482 3303
rect 11516 3269 11556 3303
rect 11590 3288 12411 3303
rect 12463 3288 12484 3340
rect 12536 3288 12556 3340
rect 12608 3327 12628 3340
rect 12680 3327 12700 3340
rect 12752 3327 12772 3340
rect 12824 3337 16439 3340
rect 12824 3327 15723 3337
rect 12847 3293 12886 3327
rect 12920 3293 12959 3327
rect 12993 3293 13032 3327
rect 13066 3293 13105 3327
rect 13139 3293 13178 3327
rect 13212 3293 13251 3327
rect 13285 3293 13324 3327
rect 13358 3293 13397 3327
rect 13431 3293 13470 3327
rect 13504 3293 13543 3327
rect 13577 3293 13616 3327
rect 13650 3293 13689 3327
rect 13723 3293 13762 3327
rect 13796 3293 13835 3327
rect 13869 3293 13908 3327
rect 13942 3293 13981 3327
rect 14015 3293 14054 3327
rect 14088 3293 14127 3327
rect 14161 3293 14200 3327
rect 14234 3293 14273 3327
rect 14307 3293 14346 3327
rect 14380 3293 14419 3327
rect 14453 3293 14492 3327
rect 14526 3293 14565 3327
rect 14599 3293 14638 3327
rect 14672 3293 14711 3327
rect 14745 3293 14784 3327
rect 14818 3293 14857 3327
rect 14891 3293 14930 3327
rect 14964 3293 15003 3327
rect 15037 3293 15076 3327
rect 15110 3293 15149 3327
rect 15183 3293 15222 3327
rect 15256 3293 15295 3327
rect 15329 3293 15368 3327
rect 15402 3293 15441 3327
rect 15475 3293 15514 3327
rect 15548 3293 15587 3327
rect 15621 3293 15660 3327
rect 15694 3293 15723 3327
rect 12608 3288 12628 3293
rect 12680 3288 12700 3293
rect 12752 3288 12772 3293
rect 12824 3288 15723 3293
rect 11590 3285 15723 3288
rect 15775 3285 15787 3337
rect 15839 3327 15851 3337
rect 15903 3327 15915 3337
rect 15967 3327 15979 3337
rect 16031 3327 16043 3337
rect 16095 3327 16107 3337
rect 15840 3293 15851 3327
rect 15913 3293 15915 3327
rect 16095 3293 16098 3327
rect 15839 3285 15851 3293
rect 15903 3285 15915 3293
rect 15967 3285 15979 3293
rect 16031 3285 16043 3293
rect 16095 3285 16107 3293
rect 16159 3285 16171 3337
rect 16223 3285 16235 3337
rect 16287 3285 16299 3337
rect 16351 3285 16363 3337
rect 16415 3327 16439 3337
rect 16424 3293 16439 3327
rect 16415 3285 16439 3293
rect 11590 3276 16439 3285
rect 11590 3269 12411 3276
rect 1153 3267 1758 3269
tri 1758 3267 1760 3269 sw
rect 1153 3255 1760 3267
tri 1760 3255 1772 3267 sw
rect 1153 3235 1772 3255
tri 1772 3235 1792 3255 sw
rect 8812 3235 12411 3269
rect 1153 3234 1792 3235
tri 1792 3234 1793 3235 sw
tri 11266 3234 11267 3235 ne
rect 11267 3234 12411 3235
rect 1153 3232 2997 3234
rect 1153 3198 1169 3232
rect 1203 3198 1241 3232
rect 1275 3198 1313 3232
rect 1347 3198 1385 3232
rect 1419 3198 1457 3232
rect 1491 3198 1529 3232
rect 1563 3198 1601 3232
rect 1635 3228 2997 3232
tri 11267 3229 11272 3234 ne
rect 11272 3229 12411 3234
rect 1635 3198 1712 3228
rect 1153 3194 1712 3198
rect 1746 3194 1785 3228
rect 1819 3194 1858 3228
rect 1892 3194 1931 3228
rect 1965 3194 2004 3228
rect 2038 3194 2077 3228
rect 2111 3194 2150 3228
rect 2184 3194 2223 3228
rect 2257 3194 2296 3228
rect 2330 3194 2369 3228
rect 2403 3194 2442 3228
rect 2476 3194 2515 3228
rect 2549 3194 2588 3228
rect 2622 3194 2661 3228
rect 2695 3194 2734 3228
rect 2768 3194 2807 3228
rect 1153 3159 2807 3194
rect 1153 3125 1169 3159
rect 1203 3125 1241 3159
rect 1275 3125 1313 3159
rect 1347 3125 1385 3159
rect 1419 3125 1457 3159
rect 1491 3125 1529 3159
rect 1563 3125 1601 3159
rect 1635 3156 2807 3159
rect 1635 3125 1712 3156
rect 1153 3122 1712 3125
rect 1746 3122 1785 3156
rect 1819 3122 1858 3156
rect 1892 3122 1931 3156
rect 1965 3122 2004 3156
rect 2038 3122 2077 3156
rect 2111 3122 2150 3156
rect 2184 3122 2223 3156
rect 2257 3122 2296 3156
rect 2330 3122 2369 3156
rect 2403 3122 2442 3156
rect 2476 3122 2515 3156
rect 2549 3122 2588 3156
rect 2622 3122 2661 3156
rect 2695 3122 2734 3156
rect 2768 3122 2807 3156
rect 2985 3122 2997 3228
rect 3718 3209 6778 3229
rect 7191 3221 8102 3229
tri 8102 3221 8110 3229 sw
tri 11272 3221 11280 3229 ne
rect 11280 3224 12411 3229
rect 12463 3224 12484 3276
rect 12536 3224 12556 3276
rect 12608 3255 12628 3276
rect 12680 3255 12700 3276
rect 12752 3255 12772 3276
rect 12824 3268 16439 3276
rect 12824 3255 15723 3268
rect 11280 3221 12594 3224
rect 12628 3221 12667 3224
rect 12701 3221 12740 3224
rect 12774 3221 12813 3224
rect 12847 3221 12886 3255
rect 12920 3221 12959 3255
rect 12993 3221 13032 3255
rect 13066 3221 13105 3255
rect 13139 3221 13178 3255
rect 13212 3221 13251 3255
rect 13285 3221 13324 3255
rect 13358 3221 13397 3255
rect 13431 3221 13470 3255
rect 13504 3221 13543 3255
rect 13577 3221 13616 3255
rect 13650 3221 13689 3255
rect 13723 3221 13762 3255
rect 13796 3221 13835 3255
rect 13869 3221 13908 3255
rect 13942 3221 13981 3255
rect 14015 3221 14054 3255
rect 14088 3221 14127 3255
rect 14161 3221 14200 3255
rect 14234 3221 14273 3255
rect 14307 3221 14346 3255
rect 14380 3221 14419 3255
rect 14453 3221 14492 3255
rect 14526 3221 14565 3255
rect 14599 3221 14638 3255
rect 14672 3221 14711 3255
rect 14745 3221 14784 3255
rect 14818 3221 14857 3255
rect 14891 3221 14930 3255
rect 14964 3221 15003 3255
rect 15037 3221 15076 3255
rect 15110 3221 15149 3255
rect 15183 3221 15222 3255
rect 15256 3221 15295 3255
rect 15329 3221 15368 3255
rect 15402 3221 15441 3255
rect 15475 3221 15514 3255
rect 15548 3221 15587 3255
rect 15621 3221 15660 3255
rect 15694 3221 15723 3255
rect 7191 3217 8110 3221
tri 8110 3217 8114 3221 sw
tri 11280 3217 11284 3221 ne
rect 11284 3217 15723 3221
rect 7191 3212 8114 3217
tri 8114 3212 8119 3217 sw
tri 11284 3212 11289 3217 ne
rect 11289 3216 15723 3217
rect 15775 3216 15787 3268
rect 15839 3255 15851 3268
rect 15903 3255 15915 3268
rect 15967 3255 15979 3268
rect 16031 3255 16043 3268
rect 16095 3255 16107 3268
rect 15840 3221 15851 3255
rect 15913 3221 15915 3255
rect 16095 3221 16098 3255
rect 15839 3216 15851 3221
rect 15903 3216 15915 3221
rect 15967 3216 15979 3221
rect 16031 3216 16043 3221
rect 16095 3216 16107 3221
rect 16159 3216 16171 3268
rect 16223 3216 16235 3268
rect 16287 3216 16299 3268
rect 16351 3216 16363 3268
rect 16415 3255 16439 3268
rect 16424 3221 16439 3255
rect 16415 3216 16439 3221
rect 11289 3212 16439 3216
rect 7191 3210 8119 3212
tri 8119 3210 8121 3212 sw
tri 11289 3210 11291 3212 ne
rect 11291 3210 16439 3212
rect 19972 3476 20038 3490
rect 19972 3424 19979 3476
rect 20031 3424 20038 3476
rect 19972 3410 20038 3424
rect 19972 3358 19979 3410
rect 20031 3358 20038 3410
rect 19972 3344 20038 3358
rect 19972 3292 19979 3344
rect 20031 3292 20038 3344
rect 19972 3278 20038 3292
rect 19972 3226 19979 3278
rect 20031 3226 20038 3278
rect 19972 3212 20038 3226
rect 7191 3209 8121 3210
rect 3718 3206 8121 3209
rect 3718 3192 4372 3206
rect 3297 3166 4372 3192
rect 3718 3154 4372 3166
rect 4424 3154 4436 3206
rect 4488 3196 8121 3206
tri 8121 3196 8135 3210 sw
rect 4488 3194 8135 3196
tri 8135 3194 8137 3196 sw
rect 4488 3156 8137 3194
tri 8137 3156 8175 3194 sw
rect 19972 3160 19979 3212
rect 20031 3160 20038 3212
rect 4488 3154 8175 3156
rect 3718 3150 8175 3154
rect 3718 3129 6388 3150
rect 6797 3148 8175 3150
tri 8175 3148 8183 3156 sw
rect 6797 3129 8183 3148
tri 8061 3122 8068 3129 ne
rect 8068 3122 8183 3129
tri 8183 3122 8209 3148 sw
rect 19972 3146 20038 3160
rect 1153 3116 2997 3122
tri 8068 3121 8069 3122 ne
rect 8069 3121 8209 3122
tri 8209 3121 8210 3122 sw
tri 8069 3116 8074 3121 ne
rect 8074 3116 8210 3121
tri 8210 3116 8215 3121 sw
rect 1153 3086 1759 3116
rect 1153 3052 1169 3086
rect 1203 3052 1241 3086
rect 1275 3052 1313 3086
rect 1347 3052 1385 3086
rect 1419 3052 1457 3086
rect 1491 3052 1529 3086
rect 1563 3052 1601 3086
rect 1635 3082 1759 3086
tri 1759 3082 1793 3116 nw
tri 8074 3082 8108 3116 ne
rect 8108 3082 8215 3116
tri 8215 3082 8249 3116 sw
rect 19972 3094 19979 3146
rect 20031 3094 20038 3146
rect 1635 3052 1725 3082
rect 1153 3048 1725 3052
tri 1725 3048 1759 3082 nw
tri 8108 3076 8114 3082 ne
rect 8114 3076 8249 3082
tri 8249 3076 8255 3082 sw
rect 19972 3080 20038 3094
tri 8114 3048 8142 3076 ne
rect 8142 3048 8255 3076
tri 8255 3048 8283 3076 sw
rect 1153 3013 1686 3048
rect 1153 2979 1169 3013
rect 1203 2979 1241 3013
rect 1275 2979 1313 3013
rect 1347 2979 1385 3013
rect 1419 2979 1457 3013
rect 1491 2979 1529 3013
rect 1563 2979 1601 3013
rect 1635 3009 1686 3013
tri 1686 3009 1725 3048 nw
tri 8142 3009 8181 3048 ne
rect 8181 3015 8283 3048
tri 8283 3015 8316 3048 sw
rect 19972 3028 19979 3080
rect 20031 3028 20038 3080
rect 8181 3009 8316 3015
tri 8316 3009 8322 3015 sw
tri 11270 3009 11276 3015 se
rect 11276 3009 13657 3015
rect 1635 3008 1685 3009
tri 1685 3008 1686 3009 nw
tri 8181 3008 8182 3009 ne
rect 8182 3008 8322 3009
tri 8322 3008 8323 3009 sw
tri 11269 3008 11270 3009 se
rect 11270 3008 13657 3009
rect 1635 2979 1651 3008
rect 1153 2940 1651 2979
tri 1651 2974 1685 3008 nw
tri 8182 2974 8216 3008 ne
rect 8216 2974 8323 3008
tri 8323 2974 8357 3008 sw
tri 11235 2974 11269 3008 se
rect 11269 2974 13657 3008
rect 1153 2906 1169 2940
rect 1203 2906 1241 2940
rect 1275 2906 1313 2940
rect 1347 2906 1385 2940
rect 1419 2906 1457 2940
rect 1491 2906 1529 2940
rect 1563 2906 1601 2940
rect 1635 2906 1651 2940
tri 8216 2936 8254 2974 ne
rect 8254 2936 8357 2974
tri 8357 2936 8395 2974 sw
tri 11197 2936 11235 2974 se
rect 11235 2936 13657 2974
tri 8254 2935 8255 2936 ne
rect 8255 2935 8395 2936
tri 8395 2935 8396 2936 sw
tri 11196 2935 11197 2936 se
rect 11197 2935 13657 2936
tri 8255 2934 8256 2935 ne
rect 8256 2934 13657 2935
rect 1153 2867 1651 2906
tri 8256 2900 8290 2934 ne
rect 8290 2900 13657 2934
tri 8290 2877 8313 2900 ne
rect 8313 2877 13657 2900
rect 19972 3014 20038 3028
rect 19972 2962 19979 3014
rect 20031 2962 20038 3014
rect 19972 2948 20038 2962
rect 19972 2896 19979 2948
rect 20031 2896 20038 2948
rect 19972 2882 20038 2896
rect 1153 2833 1169 2867
rect 1203 2833 1241 2867
rect 1275 2833 1313 2867
rect 1347 2833 1385 2867
rect 1419 2833 1457 2867
rect 1491 2833 1529 2867
rect 1563 2833 1601 2867
rect 1635 2833 1651 2867
tri 8313 2863 8327 2877 ne
rect 8327 2863 13657 2877
tri 8327 2860 8330 2863 ne
rect 8330 2860 13657 2863
tri 8330 2835 8355 2860 ne
rect 8355 2835 13657 2860
rect 1153 2794 1651 2833
rect 1153 2760 1169 2794
rect 1203 2760 1241 2794
rect 1275 2760 1313 2794
rect 1347 2760 1385 2794
rect 1419 2760 1457 2794
rect 1491 2760 1529 2794
rect 1563 2760 1601 2794
rect 1635 2760 1651 2794
rect 1153 2721 1651 2760
rect 1153 2687 1169 2721
rect 1203 2687 1241 2721
rect 1275 2687 1313 2721
rect 1347 2687 1385 2721
rect 1419 2687 1457 2721
rect 1491 2687 1529 2721
rect 1563 2687 1601 2721
rect 1635 2687 1651 2721
rect 2098 2712 2104 2764
rect 2156 2712 2168 2764
rect 2220 2712 2232 2764
rect 2284 2712 2296 2764
rect 2348 2712 2360 2764
rect 2412 2712 2424 2764
rect 2476 2712 3010 2764
rect 5038 2699 5064 2829
rect 13292 2786 13408 2792
rect 7092 2773 8004 2779
rect 7092 2721 7730 2773
rect 7782 2721 7794 2773
rect 7846 2721 8004 2773
rect 7092 2715 8004 2721
rect 11186 2702 13258 2736
rect 1153 2648 1651 2687
rect 1153 2614 1169 2648
rect 1203 2614 1241 2648
rect 1275 2614 1313 2648
rect 1347 2614 1385 2648
rect 1419 2614 1457 2648
rect 1491 2614 1529 2648
rect 1563 2614 1601 2648
rect 1635 2614 1651 2648
rect 1153 2575 1651 2614
rect 1153 2541 1169 2575
rect 1203 2541 1241 2575
rect 1275 2541 1313 2575
rect 1347 2541 1385 2575
rect 1419 2541 1457 2575
rect 1491 2541 1529 2575
rect 1563 2541 1601 2575
rect 1635 2541 1651 2575
rect 1153 2502 1651 2541
rect 1153 2468 1169 2502
rect 1203 2468 1241 2502
rect 1275 2468 1313 2502
rect 1347 2468 1385 2502
rect 1419 2468 1457 2502
rect 1491 2468 1529 2502
rect 1563 2468 1601 2502
rect 1635 2468 1651 2502
rect 11186 2668 11198 2702
rect 11232 2668 11272 2702
rect 11306 2668 11346 2702
rect 11380 2668 11420 2702
rect 11454 2668 11494 2702
rect 11528 2668 11568 2702
rect 11602 2668 11642 2702
rect 11676 2668 11716 2702
rect 11750 2668 11790 2702
rect 11824 2668 11864 2702
rect 11898 2668 11938 2702
rect 11972 2668 12012 2702
rect 12046 2668 12087 2702
rect 12121 2668 12162 2702
rect 12196 2668 12237 2702
rect 12271 2668 12312 2702
rect 12346 2668 12387 2702
rect 12421 2701 12462 2702
rect 12496 2701 12537 2702
rect 12571 2701 12612 2702
rect 12646 2701 12687 2702
rect 12721 2701 12762 2702
rect 12796 2701 12837 2702
rect 12610 2668 12612 2701
rect 12682 2668 12687 2701
rect 12754 2668 12762 2701
rect 12826 2668 12837 2701
rect 12871 2668 12912 2702
rect 12946 2668 12987 2702
rect 13021 2668 13062 2702
rect 13096 2668 13137 2702
rect 13171 2668 13212 2702
rect 13246 2668 13258 2702
rect 11186 2649 12414 2668
rect 12466 2649 12486 2668
rect 12538 2649 12558 2668
rect 12610 2649 12630 2668
rect 12682 2649 12702 2668
rect 12754 2649 12774 2668
rect 12826 2649 13258 2668
rect 13344 2734 13356 2786
rect 14334 2761 14340 2877
rect 14456 2863 16733 2877
tri 16733 2863 16747 2877 sw
rect 14456 2860 16747 2863
tri 16747 2860 16750 2863 sw
rect 14456 2846 16750 2860
tri 16750 2846 16764 2860 sw
rect 14456 2826 16764 2846
tri 16764 2826 16784 2846 sw
rect 14456 2807 16784 2826
tri 16784 2807 16803 2826 sw
rect 14456 2761 16803 2807
rect 17481 2794 17487 2846
rect 17539 2794 17551 2846
rect 17603 2794 17609 2846
rect 19972 2830 19979 2882
rect 20031 2830 20038 2882
rect 19972 2816 20038 2830
rect 19972 2764 19979 2816
rect 20031 2764 20038 2816
rect 13292 2719 13408 2734
rect 13344 2667 13356 2719
rect 13292 2661 13408 2667
rect 19972 2750 20038 2764
rect 19972 2698 19979 2750
rect 20031 2698 20038 2750
rect 19972 2684 20038 2698
rect 11186 2637 13258 2649
rect 11186 2630 12414 2637
rect 12466 2630 12486 2637
rect 12538 2630 12558 2637
rect 12610 2630 12630 2637
rect 12682 2630 12702 2637
rect 12754 2630 12774 2637
rect 12826 2630 13258 2637
rect 19972 2632 19979 2684
rect 20031 2632 20038 2684
rect 11186 2596 11198 2630
rect 11232 2596 11272 2630
rect 11306 2596 11346 2630
rect 11380 2596 11420 2630
rect 11454 2596 11494 2630
rect 11528 2596 11568 2630
rect 11602 2596 11642 2630
rect 11676 2596 11716 2630
rect 11750 2596 11790 2630
rect 11824 2596 11864 2630
rect 11898 2596 11938 2630
rect 11972 2596 12012 2630
rect 12046 2596 12087 2630
rect 12121 2596 12162 2630
rect 12196 2596 12237 2630
rect 12271 2596 12312 2630
rect 12346 2596 12387 2630
rect 12610 2596 12612 2630
rect 12682 2596 12687 2630
rect 12754 2596 12762 2630
rect 12826 2596 12837 2630
rect 12871 2596 12912 2630
rect 12946 2596 12987 2630
rect 13021 2596 13062 2630
rect 13096 2596 13137 2630
rect 13171 2596 13212 2630
rect 13246 2596 13258 2630
rect 11186 2585 12414 2596
rect 12466 2585 12486 2596
rect 12538 2585 12558 2596
rect 12610 2585 12630 2596
rect 12682 2585 12702 2596
rect 12754 2585 12774 2596
rect 12826 2585 13258 2596
rect 11186 2573 13258 2585
rect 11186 2558 12414 2573
rect 12466 2558 12486 2573
rect 12538 2558 12558 2573
rect 12610 2558 12630 2573
rect 12682 2558 12702 2573
rect 12754 2558 12774 2573
rect 12826 2558 13258 2573
rect 11186 2524 11198 2558
rect 11232 2524 11272 2558
rect 11306 2524 11346 2558
rect 11380 2524 11420 2558
rect 11454 2524 11494 2558
rect 11528 2524 11568 2558
rect 11602 2524 11642 2558
rect 11676 2524 11716 2558
rect 11750 2524 11790 2558
rect 11824 2524 11864 2558
rect 11898 2524 11938 2558
rect 11972 2524 12012 2558
rect 12046 2524 12087 2558
rect 12121 2524 12162 2558
rect 12196 2524 12237 2558
rect 12271 2524 12312 2558
rect 12346 2524 12387 2558
rect 12610 2524 12612 2558
rect 12682 2524 12687 2558
rect 12754 2524 12762 2558
rect 12826 2524 12837 2558
rect 12871 2524 12912 2558
rect 12946 2524 12987 2558
rect 13021 2524 13062 2558
rect 13096 2524 13137 2558
rect 13171 2524 13212 2558
rect 13246 2524 13258 2558
rect 11186 2521 12414 2524
rect 12466 2521 12486 2524
rect 12538 2521 12558 2524
rect 12610 2521 12630 2524
rect 12682 2521 12702 2524
rect 12754 2521 12774 2524
rect 12826 2521 13258 2524
rect 11186 2490 13258 2521
rect 13416 2558 13532 2564
rect 13468 2506 13480 2558
tri 13532 2530 13544 2542 sw
rect 13532 2517 13544 2530
tri 13544 2517 13557 2530 sw
rect 13532 2506 16501 2517
rect 13416 2491 16501 2506
rect 1153 2456 1651 2468
tri 1651 2456 1673 2478 sw
rect 1153 2433 1673 2456
tri 1673 2433 1696 2456 sw
rect 13468 2439 13480 2491
rect 13532 2465 16501 2491
rect 16553 2465 16565 2517
rect 16617 2465 16623 2517
rect 17263 2516 17269 2632
rect 17385 2516 17391 2632
rect 19972 2618 20038 2632
rect 19972 2566 19979 2618
rect 20031 2566 20038 2618
rect 19972 2552 20038 2566
rect 19972 2500 19979 2552
rect 20031 2500 20038 2552
rect 19972 2494 20038 2500
rect 20070 3802 20136 3808
rect 20070 3750 20077 3802
rect 20129 3750 20136 3802
rect 20070 3737 20136 3750
rect 20070 3685 20077 3737
rect 20129 3685 20136 3737
rect 20070 3672 20136 3685
rect 20070 3620 20077 3672
rect 20129 3620 20136 3672
rect 20070 3607 20136 3620
rect 20070 3555 20077 3607
rect 20129 3555 20136 3607
rect 20070 3542 20136 3555
rect 20070 3490 20077 3542
rect 20129 3490 20136 3542
rect 20070 3476 20136 3490
rect 20070 3424 20077 3476
rect 20129 3424 20136 3476
rect 20070 3410 20136 3424
rect 20070 3358 20077 3410
rect 20129 3358 20136 3410
rect 20070 3344 20136 3358
rect 20070 3292 20077 3344
rect 20129 3292 20136 3344
rect 20070 3278 20136 3292
rect 20070 3226 20077 3278
rect 20129 3226 20136 3278
rect 20070 3212 20136 3226
rect 20070 3160 20077 3212
rect 20129 3160 20136 3212
rect 20070 3146 20136 3160
rect 20070 3094 20077 3146
rect 20129 3094 20136 3146
rect 20070 3080 20136 3094
rect 20070 3028 20077 3080
rect 20129 3028 20136 3080
rect 20070 3014 20136 3028
rect 20070 2962 20077 3014
rect 20129 2962 20136 3014
rect 20070 2948 20136 2962
rect 20070 2896 20077 2948
rect 20129 2896 20136 2948
rect 20070 2882 20136 2896
rect 20070 2830 20077 2882
rect 20129 2830 20136 2882
rect 20070 2816 20136 2830
rect 20070 2764 20077 2816
rect 20129 2764 20136 2816
rect 20070 2750 20136 2764
rect 20070 2698 20077 2750
rect 20129 2698 20136 2750
rect 20070 2684 20136 2698
rect 20070 2632 20077 2684
rect 20129 2632 20136 2684
rect 20070 2618 20136 2632
rect 20070 2566 20077 2618
rect 20129 2566 20136 2618
rect 20070 2552 20136 2566
rect 20070 2500 20077 2552
rect 20129 2500 20136 2552
rect 20070 2494 20136 2500
rect 23562 3780 23593 3814
rect 23627 3780 23665 3814
rect 23699 3780 23737 3814
rect 23771 3780 23802 3814
rect 23562 3741 23802 3780
rect 23562 3707 23593 3741
rect 23627 3707 23665 3741
rect 23699 3707 23737 3741
rect 23771 3707 23802 3741
rect 23562 3668 23802 3707
rect 23562 3634 23593 3668
rect 23627 3634 23665 3668
rect 23699 3634 23737 3668
rect 23771 3634 23802 3668
rect 23562 3595 23802 3634
rect 23562 3561 23593 3595
rect 23627 3561 23665 3595
rect 23699 3561 23737 3595
rect 23771 3561 23802 3595
rect 23562 3522 23802 3561
rect 23562 3488 23593 3522
rect 23627 3488 23665 3522
rect 23699 3488 23737 3522
rect 23771 3488 23802 3522
rect 23562 3449 23802 3488
rect 23562 3415 23593 3449
rect 23627 3415 23665 3449
rect 23699 3415 23737 3449
rect 23771 3415 23802 3449
rect 23562 3376 23802 3415
rect 23562 3342 23593 3376
rect 23627 3342 23665 3376
rect 23699 3342 23737 3376
rect 23771 3342 23802 3376
rect 23562 3303 23802 3342
rect 23562 3269 23593 3303
rect 23627 3269 23665 3303
rect 23699 3269 23737 3303
rect 23771 3269 23802 3303
rect 23562 3230 23802 3269
rect 23562 3196 23593 3230
rect 23627 3196 23665 3230
rect 23699 3196 23737 3230
rect 23771 3196 23802 3230
rect 23562 3156 23802 3196
rect 23562 3122 23593 3156
rect 23627 3122 23665 3156
rect 23699 3122 23737 3156
rect 23771 3122 23802 3156
rect 23562 3082 23802 3122
rect 23562 3048 23593 3082
rect 23627 3048 23665 3082
rect 23699 3048 23737 3082
rect 23771 3048 23802 3082
rect 23562 3008 23802 3048
rect 23562 2974 23593 3008
rect 23627 2974 23665 3008
rect 23699 2974 23737 3008
rect 23771 2974 23802 3008
rect 23562 2934 23802 2974
rect 23562 2900 23593 2934
rect 23627 2900 23665 2934
rect 23699 2900 23737 2934
rect 23771 2900 23802 2934
rect 23562 2860 23802 2900
rect 23562 2826 23593 2860
rect 23627 2826 23665 2860
rect 23699 2826 23737 2860
rect 23771 2826 23802 2860
rect 23562 2786 23802 2826
rect 23562 2752 23593 2786
rect 23627 2752 23665 2786
rect 23699 2752 23737 2786
rect 23771 2752 23802 2786
rect 23562 2712 23802 2752
rect 23562 2678 23593 2712
rect 23627 2678 23665 2712
rect 23699 2678 23737 2712
rect 23771 2678 23802 2712
rect 23562 2638 23802 2678
rect 23562 2604 23593 2638
rect 23627 2604 23665 2638
rect 23699 2604 23737 2638
rect 23771 2604 23802 2638
rect 23562 2564 23802 2604
rect 23562 2530 23593 2564
rect 23627 2530 23665 2564
rect 23699 2530 23737 2564
rect 23771 2530 23802 2564
rect 23562 2490 23802 2530
rect 13532 2456 13548 2465
tri 13548 2456 13557 2465 nw
rect 23562 2456 23593 2490
rect 23627 2456 23665 2490
rect 23699 2456 23737 2490
rect 23771 2456 23802 2490
tri 13532 2440 13548 2456 nw
rect 13416 2433 13532 2439
rect 1153 2429 1696 2433
rect 1153 2395 1169 2429
rect 1203 2395 1241 2429
rect 1275 2395 1313 2429
rect 1347 2395 1385 2429
rect 1419 2395 1457 2429
rect 1491 2395 1529 2429
rect 1563 2395 1601 2429
rect 1635 2425 1696 2429
tri 1696 2425 1704 2433 sw
rect 1635 2416 1704 2425
tri 1704 2416 1713 2425 sw
rect 23562 2416 23802 2456
rect 1635 2415 1713 2416
tri 1713 2415 1714 2416 sw
rect 1635 2409 1714 2415
tri 1714 2409 1720 2415 sw
rect 7092 2409 8574 2415
rect 1635 2395 1720 2409
rect 1153 2375 1720 2395
tri 1720 2375 1754 2409 sw
rect 7092 2375 7104 2409
rect 7138 2375 7179 2409
rect 7213 2375 7254 2409
rect 7288 2375 7329 2409
rect 7363 2375 7403 2409
rect 7437 2375 7477 2409
rect 7511 2375 7551 2409
rect 7585 2375 7625 2409
rect 7659 2375 7699 2409
rect 7733 2375 7773 2409
rect 7807 2375 7847 2409
rect 7881 2375 7921 2409
rect 7955 2375 7995 2409
rect 8029 2375 8069 2409
rect 8103 2375 8143 2409
rect 8177 2375 8217 2409
rect 8251 2375 8291 2409
rect 8325 2375 8365 2409
rect 8399 2375 8439 2409
rect 8473 2375 8513 2409
rect 8547 2382 8574 2409
tri 13229 2399 13235 2405 se
rect 13235 2399 13351 2405
tri 8574 2382 8591 2399 sw
tri 13212 2382 13229 2399 se
rect 13229 2390 13351 2399
rect 13229 2382 13235 2390
rect 8547 2375 8591 2382
rect 1153 2356 1754 2375
rect 1153 2322 1169 2356
rect 1203 2322 1241 2356
rect 1275 2322 1313 2356
rect 1347 2322 1385 2356
rect 1419 2322 1457 2356
rect 1491 2322 1529 2356
rect 1563 2322 1601 2356
rect 1635 2352 1754 2356
tri 1754 2352 1777 2375 sw
rect 7092 2374 8591 2375
tri 8591 2374 8599 2382 sw
tri 13204 2374 13212 2382 se
rect 13212 2374 13235 2382
rect 3310 2352 3710 2372
tri 3710 2352 3730 2372 sw
tri 3990 2352 4010 2372 se
rect 1635 2342 1777 2352
tri 1777 2342 1787 2352 sw
rect 3310 2347 3730 2352
tri 3730 2347 3735 2352 sw
tri 3985 2347 3990 2352 se
rect 3990 2347 4010 2352
tri 4140 2352 4160 2372 sw
tri 5942 2352 5962 2372 se
rect 4140 2347 4160 2352
tri 4160 2347 4165 2352 sw
tri 5937 2347 5942 2352 se
rect 5942 2347 5962 2352
tri 6092 2352 6112 2372 sw
tri 6372 2352 6392 2372 se
rect 6392 2352 6792 2372
rect 6092 2347 6112 2352
tri 6112 2347 6117 2352 sw
tri 6367 2347 6372 2352 se
rect 6372 2347 6792 2352
rect 1635 2337 1787 2342
tri 1787 2337 1792 2342 sw
rect 1635 2336 1792 2337
tri 1792 2336 1793 2337 sw
rect 1635 2330 3010 2336
rect 1635 2322 1712 2330
rect 1153 2296 1712 2322
rect 1746 2296 1786 2330
rect 1820 2296 1860 2330
rect 1894 2296 1934 2330
rect 1968 2296 2008 2330
rect 2042 2296 2082 2330
rect 2116 2296 2156 2330
rect 2190 2296 2230 2330
rect 2264 2296 2304 2330
rect 2338 2296 2378 2330
rect 2412 2296 2452 2330
rect 2486 2296 2526 2330
rect 2560 2296 2599 2330
rect 2633 2296 2672 2330
rect 2706 2296 2745 2330
rect 2779 2296 2818 2330
rect 2852 2296 2891 2330
rect 2925 2296 2964 2330
rect 2998 2296 3010 2330
rect 1153 2283 3010 2296
rect 1153 2249 1169 2283
rect 1203 2249 1241 2283
rect 1275 2249 1313 2283
rect 1347 2249 1385 2283
rect 1419 2249 1457 2283
rect 1491 2249 1529 2283
rect 1563 2249 1601 2283
rect 1635 2258 3010 2283
rect 1635 2249 1712 2258
rect 1153 2224 1712 2249
rect 1746 2224 1786 2258
rect 1820 2224 1860 2258
rect 1894 2224 1934 2258
rect 1968 2224 2008 2258
rect 2042 2224 2082 2258
rect 2116 2224 2156 2258
rect 2190 2224 2230 2258
rect 2264 2224 2304 2258
rect 2338 2224 2378 2258
rect 2412 2224 2452 2258
rect 2486 2224 2526 2258
rect 2560 2224 2599 2258
rect 2633 2224 2672 2258
rect 2706 2224 2745 2258
rect 2779 2224 2818 2258
rect 2852 2224 2891 2258
rect 2925 2224 2964 2258
rect 2998 2224 3010 2258
rect 1153 2218 3010 2224
rect 3310 2331 6792 2347
rect 1153 2210 1784 2218
rect 1153 2176 1169 2210
rect 1203 2176 1241 2210
rect 1275 2176 1313 2210
rect 1347 2176 1385 2210
rect 1419 2176 1457 2210
rect 1491 2176 1529 2210
rect 1563 2176 1601 2210
rect 1635 2209 1784 2210
tri 1784 2209 1793 2218 nw
rect 3310 2215 5862 2331
rect 5978 2215 6792 2331
rect 7092 2338 13235 2374
rect 13287 2338 13299 2390
rect 7092 2337 13351 2338
rect 7092 2303 7104 2337
rect 7138 2303 7179 2337
rect 7213 2303 7254 2337
rect 7288 2303 7329 2337
rect 7363 2303 7403 2337
rect 7437 2303 7477 2337
rect 7511 2303 7551 2337
rect 7585 2303 7625 2337
rect 7659 2303 7699 2337
rect 7733 2303 7773 2337
rect 7807 2303 7847 2337
rect 7881 2303 7921 2337
rect 7955 2303 7995 2337
rect 8029 2303 8069 2337
rect 8103 2303 8143 2337
rect 8177 2303 8217 2337
rect 8251 2303 8291 2337
rect 8325 2303 8365 2337
rect 8399 2303 8439 2337
rect 8473 2303 8513 2337
rect 8547 2323 13351 2337
rect 8547 2303 13235 2323
rect 7092 2281 13235 2303
rect 7092 2279 8602 2281
tri 8602 2279 8604 2281 nw
tri 13219 2279 13221 2281 ne
rect 13221 2279 13235 2281
rect 7092 2268 8591 2279
tri 8591 2268 8602 2279 nw
tri 13221 2268 13232 2279 ne
rect 13232 2271 13235 2279
rect 13287 2271 13299 2323
rect 23562 2382 23593 2416
rect 23627 2382 23665 2416
rect 23699 2382 23737 2416
rect 23771 2382 23802 2416
rect 23562 2342 23802 2382
rect 23562 2308 23593 2342
rect 23627 2308 23665 2342
rect 23699 2308 23737 2342
rect 23771 2308 23802 2342
tri 23534 2279 23562 2307 se
rect 23562 2279 23802 2308
rect 13232 2268 13351 2271
tri 23523 2268 23534 2279 se
rect 23534 2268 23802 2279
rect 7092 2265 8574 2268
rect 7092 2231 7104 2265
rect 7138 2231 7179 2265
rect 7213 2231 7254 2265
rect 7288 2231 7329 2265
rect 7363 2231 7403 2265
rect 7437 2231 7477 2265
rect 7511 2231 7551 2265
rect 7585 2231 7625 2265
rect 7659 2231 7699 2265
rect 7733 2231 7773 2265
rect 7807 2231 7847 2265
rect 7881 2231 7921 2265
rect 7955 2231 7995 2265
rect 8029 2231 8069 2265
rect 8103 2231 8143 2265
rect 8177 2231 8217 2265
rect 8251 2231 8291 2265
rect 8325 2231 8365 2265
rect 8399 2231 8439 2265
rect 8473 2231 8513 2265
rect 8547 2231 8574 2265
tri 8574 2251 8591 2268 nw
tri 13232 2265 13235 2268 ne
rect 13235 2265 13351 2268
tri 23520 2265 23523 2268 se
rect 23523 2265 23593 2268
tri 23506 2251 23520 2265 se
rect 23520 2251 23593 2265
tri 23489 2234 23506 2251 se
rect 23506 2234 23593 2251
rect 23627 2234 23665 2268
rect 23699 2234 23737 2268
rect 23771 2234 23802 2268
rect 7092 2225 8574 2231
tri 23480 2225 23489 2234 se
rect 23489 2225 23802 2234
rect 1635 2206 1781 2209
tri 1781 2206 1784 2209 nw
rect 1635 2194 1769 2206
tri 1769 2194 1781 2206 nw
rect 3310 2203 6792 2215
tri 23461 2206 23480 2225 se
rect 23480 2206 23802 2225
tri 23458 2203 23461 2206 se
rect 23461 2203 23802 2206
rect 3710 2194 3726 2203
tri 3726 2194 3735 2203 nw
tri 3985 2194 3994 2203 ne
rect 3994 2194 4010 2203
rect 1635 2176 1735 2194
rect 1153 2160 1735 2176
tri 1735 2160 1769 2194 nw
tri 3710 2178 3726 2194 nw
tri 3994 2178 4010 2194 ne
rect 4140 2194 4156 2203
tri 4156 2194 4165 2203 nw
tri 5937 2194 5946 2203 ne
rect 5946 2194 5962 2203
tri 4140 2178 4156 2194 nw
tri 5946 2178 5962 2194 ne
rect 6092 2194 6108 2203
tri 6108 2194 6117 2203 nw
tri 6367 2194 6376 2203 ne
rect 6376 2194 6392 2203
tri 23449 2194 23458 2203 se
rect 23458 2194 23802 2203
tri 6092 2178 6108 2194 nw
tri 6376 2178 6392 2194 ne
tri 23433 2178 23449 2194 se
rect 23449 2178 23593 2194
tri 23415 2160 23433 2178 se
rect 23433 2160 23593 2178
rect 23627 2160 23665 2194
rect 23699 2160 23737 2194
rect 23771 2160 23802 2194
rect 1153 2154 1729 2160
tri 1729 2154 1735 2160 nw
rect 11307 2154 13258 2160
rect 1153 2137 1651 2154
rect 1153 2103 1169 2137
rect 1203 2103 1241 2137
rect 1275 2103 1313 2137
rect 1347 2103 1385 2137
rect 1419 2103 1457 2137
rect 1491 2103 1529 2137
rect 1563 2103 1601 2137
rect 1635 2103 1651 2137
rect 1153 2064 1651 2103
tri 1651 2076 1729 2154 nw
tri 11260 2076 11307 2123 se
rect 11307 2076 11319 2154
rect 1153 2030 1169 2064
rect 1203 2030 1241 2064
rect 1275 2030 1313 2064
rect 1347 2030 1385 2064
rect 1419 2030 1457 2064
rect 1491 2030 1529 2064
rect 1563 2030 1601 2064
rect 1635 2030 1651 2064
rect 1153 1991 1651 2030
rect 1153 1957 1169 1991
rect 1203 1957 1241 1991
rect 1275 1957 1313 1991
rect 1347 1957 1385 1991
rect 1419 1957 1457 1991
rect 1491 1957 1529 1991
rect 1563 1957 1601 1991
rect 1635 1957 1651 1991
tri 11165 1981 11260 2076 se
rect 11260 1981 11319 2076
rect 1153 1918 1651 1957
rect 1153 1884 1169 1918
rect 1203 1884 1241 1918
rect 1275 1884 1313 1918
rect 1347 1884 1385 1918
rect 1419 1884 1457 1918
rect 1491 1884 1529 1918
rect 1563 1884 1601 1918
rect 1635 1884 1651 1918
rect 1153 1845 1651 1884
rect 8762 1975 11319 1981
rect 11713 2120 11752 2154
rect 11786 2120 11825 2154
rect 11859 2120 11898 2154
rect 11932 2120 11971 2154
rect 12005 2120 12044 2154
rect 12078 2120 12117 2154
rect 12151 2120 12190 2154
rect 12224 2120 12263 2154
rect 12297 2120 12336 2154
rect 12370 2120 12409 2154
rect 12443 2143 12482 2154
rect 12516 2143 12555 2154
rect 12589 2143 12628 2154
rect 12662 2143 12701 2154
rect 12735 2143 12774 2154
rect 12808 2143 12847 2154
rect 12464 2120 12482 2143
rect 12538 2120 12555 2143
rect 12612 2120 12628 2143
rect 12686 2120 12701 2143
rect 12759 2120 12774 2143
rect 12832 2120 12847 2143
rect 12881 2120 12920 2154
rect 12954 2120 12993 2154
rect 13027 2120 13066 2154
rect 13100 2120 13139 2154
rect 13173 2120 13212 2154
rect 13246 2120 13258 2154
tri 23388 2133 23415 2160 se
rect 23415 2133 23802 2160
tri 23375 2120 23388 2133 se
rect 23388 2120 23802 2133
rect 11713 2091 12412 2120
rect 12464 2091 12486 2120
rect 12538 2091 12560 2120
rect 12612 2091 12634 2120
rect 12686 2091 12707 2120
rect 12759 2091 12780 2120
rect 12832 2091 13258 2120
tri 23353 2098 23375 2120 se
rect 23375 2098 23593 2120
rect 11713 2082 13258 2091
rect 11713 2048 11752 2082
rect 11786 2048 11825 2082
rect 11859 2048 11898 2082
rect 11932 2048 11971 2082
rect 12005 2048 12044 2082
rect 12078 2048 12117 2082
rect 12151 2048 12190 2082
rect 12224 2048 12263 2082
rect 12297 2048 12336 2082
rect 12370 2048 12409 2082
rect 12443 2079 12482 2082
rect 12516 2079 12555 2082
rect 12589 2079 12628 2082
rect 12662 2079 12701 2082
rect 12735 2079 12774 2082
rect 12808 2079 12847 2082
rect 12464 2048 12482 2079
rect 12538 2048 12555 2079
rect 12612 2048 12628 2079
rect 12686 2048 12701 2079
rect 12759 2048 12774 2079
rect 12832 2048 12847 2079
rect 12881 2048 12920 2082
rect 12954 2048 12993 2082
rect 13027 2048 13066 2082
rect 13100 2048 13139 2082
rect 13173 2048 13212 2082
rect 13246 2048 13258 2082
rect 11713 2027 12412 2048
rect 12464 2027 12486 2048
rect 12538 2027 12560 2048
rect 12612 2027 12634 2048
rect 12686 2027 12707 2048
rect 12759 2027 12780 2048
rect 12832 2027 13258 2048
rect 11713 2015 13258 2027
rect 11713 2010 12412 2015
rect 12464 2010 12486 2015
rect 12538 2010 12560 2015
rect 12612 2010 12634 2015
rect 12686 2010 12707 2015
rect 12759 2010 12780 2015
rect 12832 2010 13258 2015
rect 11713 1976 11752 2010
rect 11786 1976 11825 2010
rect 11859 1976 11898 2010
rect 11932 1976 11971 2010
rect 12005 1976 12044 2010
rect 12078 1976 12117 2010
rect 12151 1976 12190 2010
rect 12224 1976 12263 2010
rect 12297 1976 12336 2010
rect 12370 1976 12409 2010
rect 12464 1976 12482 2010
rect 12538 1976 12555 2010
rect 12612 1976 12628 2010
rect 12686 1976 12701 2010
rect 12759 1976 12774 2010
rect 12832 1976 12847 2010
rect 12881 1976 12920 2010
rect 12954 1976 12993 2010
rect 13027 1976 13066 2010
rect 13100 1976 13139 2010
rect 13173 1976 13212 2010
rect 13246 1976 13258 2010
rect 8762 1941 8774 1975
rect 8808 1941 8847 1975
rect 8881 1941 8920 1975
rect 8954 1941 8993 1975
rect 9027 1941 9066 1975
rect 9100 1941 9139 1975
rect 9173 1941 9212 1975
rect 9246 1941 9285 1975
rect 9319 1941 9358 1975
rect 9392 1941 9431 1975
rect 9465 1941 9504 1975
rect 9538 1941 9577 1975
rect 9611 1941 9650 1975
rect 9684 1941 9723 1975
rect 9757 1941 9796 1975
rect 9830 1941 9869 1975
rect 9903 1941 9942 1975
rect 9976 1941 10015 1975
rect 10049 1941 10088 1975
rect 10122 1941 10161 1975
rect 10195 1941 10234 1975
rect 10268 1941 10307 1975
rect 10341 1941 10380 1975
rect 10414 1941 10453 1975
rect 10487 1941 10526 1975
rect 10560 1941 10599 1975
rect 8762 1903 10599 1941
rect 8762 1869 8774 1903
rect 8808 1869 8847 1903
rect 8881 1869 8920 1903
rect 8954 1869 8993 1903
rect 9027 1869 9066 1903
rect 9100 1869 9139 1903
rect 9173 1869 9212 1903
rect 9246 1869 9285 1903
rect 9319 1869 9358 1903
rect 9392 1869 9431 1903
rect 9465 1869 9504 1903
rect 9538 1869 9577 1903
rect 9611 1869 9650 1903
rect 9684 1869 9723 1903
rect 9757 1869 9796 1903
rect 9830 1869 9869 1903
rect 9903 1869 9942 1903
rect 9976 1869 10015 1903
rect 10049 1869 10088 1903
rect 10122 1869 10161 1903
rect 10195 1869 10234 1903
rect 10268 1869 10307 1903
rect 10341 1869 10380 1903
rect 10414 1869 10453 1903
rect 10487 1869 10526 1903
rect 10560 1869 10599 1903
rect 11713 1963 12412 1976
rect 12464 1963 12486 1976
rect 12538 1963 12560 1976
rect 12612 1963 12634 1976
rect 12686 1963 12707 1976
rect 12759 1963 12780 1976
rect 12832 1963 13258 1976
rect 11713 1951 13258 1963
rect 11713 1938 12412 1951
rect 12464 1938 12486 1951
rect 12538 1938 12560 1951
rect 12612 1938 12634 1951
rect 12686 1938 12707 1951
rect 12759 1938 12780 1951
rect 12832 1938 13258 1951
rect 11713 1904 11752 1938
rect 11786 1904 11825 1938
rect 11859 1904 11898 1938
rect 11932 1904 11971 1938
rect 12005 1904 12044 1938
rect 12078 1904 12117 1938
rect 12151 1904 12190 1938
rect 12224 1904 12263 1938
rect 12297 1904 12336 1938
rect 12370 1904 12409 1938
rect 12464 1904 12482 1938
rect 12538 1904 12555 1938
rect 12612 1904 12628 1938
rect 12686 1904 12701 1938
rect 12759 1904 12774 1938
rect 12832 1904 12847 1938
rect 12881 1904 12920 1938
rect 12954 1904 12993 1938
rect 13027 1904 13066 1938
rect 13100 1904 13139 1938
rect 13173 1904 13212 1938
rect 13246 1904 13258 1938
rect 13604 1918 17052 2098
tri 23341 2086 23353 2098 se
rect 23353 2086 23593 2098
rect 23627 2086 23665 2120
rect 23699 2086 23737 2120
rect 23771 2086 23802 2120
tri 23315 2060 23341 2086 se
rect 23341 2060 23802 2086
tri 23301 2046 23315 2060 se
rect 23315 2046 23802 2060
tri 23267 2012 23301 2046 se
rect 23301 2012 23593 2046
rect 23627 2012 23665 2046
rect 23699 2012 23737 2046
rect 23771 2012 23802 2046
tri 23242 1987 23267 2012 se
rect 23267 1987 23802 2012
tri 23227 1972 23242 1987 se
rect 23242 1972 23802 1987
tri 23193 1938 23227 1972 se
rect 23227 1938 23593 1972
rect 23627 1938 23665 1972
rect 23699 1938 23737 1972
rect 23771 1938 23802 1972
tri 23173 1918 23193 1938 se
rect 23193 1918 23802 1938
tri 23169 1914 23173 1918 se
rect 23173 1916 23802 1918
rect 23173 1914 23800 1916
tri 23800 1914 23802 1916 nw
rect 23943 4800 23981 5652
rect 24087 5652 24541 5658
rect 24087 4800 24125 5652
tri 24125 5510 24267 5652 nw
rect 23943 4761 24125 4800
rect 23943 4727 23981 4761
rect 24015 4727 24053 4761
rect 24087 4727 24125 4761
rect 23943 4688 24125 4727
rect 23943 4654 23981 4688
rect 24015 4654 24053 4688
rect 24087 4654 24125 4688
rect 23943 4615 24125 4654
rect 23943 4581 23981 4615
rect 24015 4581 24053 4615
rect 24087 4581 24125 4615
rect 23943 4542 24125 4581
rect 23943 4508 23981 4542
rect 24015 4508 24053 4542
rect 24087 4508 24125 4542
rect 23943 4469 24125 4508
rect 23943 4435 23981 4469
rect 24015 4435 24053 4469
rect 24087 4435 24125 4469
rect 23943 4396 24125 4435
rect 23943 4362 23981 4396
rect 24015 4362 24053 4396
rect 24087 4362 24125 4396
rect 23943 4323 24125 4362
rect 23943 4289 23981 4323
rect 24015 4289 24053 4323
rect 24087 4289 24125 4323
rect 23943 4250 24125 4289
rect 23943 4216 23981 4250
rect 24015 4216 24053 4250
rect 24087 4216 24125 4250
rect 23943 4177 24125 4216
rect 23943 4143 23981 4177
rect 24015 4143 24053 4177
rect 24087 4143 24125 4177
rect 23943 4104 24125 4143
rect 23943 4070 23981 4104
rect 24015 4070 24053 4104
rect 24087 4070 24125 4104
rect 23943 4031 24125 4070
rect 23943 3997 23981 4031
rect 24015 3997 24053 4031
rect 24087 3997 24125 4031
rect 23943 3958 24125 3997
rect 23943 3924 23981 3958
rect 24015 3924 24053 3958
rect 24087 3924 24125 3958
rect 23943 3885 24125 3924
rect 23943 3851 23981 3885
rect 24015 3851 24053 3885
rect 24087 3851 24125 3885
rect 23943 3812 24125 3851
rect 23943 3778 23981 3812
rect 24015 3778 24053 3812
rect 24087 3778 24125 3812
rect 23943 3739 24125 3778
rect 23943 3705 23981 3739
rect 24015 3705 24053 3739
rect 24087 3705 24125 3739
rect 23943 3666 24125 3705
rect 23943 3632 23981 3666
rect 24015 3632 24053 3666
rect 24087 3632 24125 3666
rect 23943 3593 24125 3632
rect 23943 3559 23981 3593
rect 24015 3559 24053 3593
rect 24087 3559 24125 3593
rect 23943 3520 24125 3559
rect 23943 3486 23981 3520
rect 24015 3486 24053 3520
rect 24087 3486 24125 3520
rect 23943 3447 24125 3486
rect 23943 3413 23981 3447
rect 24015 3413 24053 3447
rect 24087 3413 24125 3447
rect 23943 3374 24125 3413
rect 23943 3340 23981 3374
rect 24015 3340 24053 3374
rect 24087 3340 24125 3374
rect 23943 3301 24125 3340
rect 23943 3267 23981 3301
rect 24015 3267 24053 3301
rect 24087 3267 24125 3301
rect 23943 3228 24125 3267
rect 23943 3194 23981 3228
rect 24015 3194 24053 3228
rect 24087 3194 24125 3228
rect 23943 3155 24125 3194
rect 23943 3121 23981 3155
rect 24015 3121 24053 3155
rect 24087 3121 24125 3155
rect 23943 3082 24125 3121
rect 23943 3048 23981 3082
rect 24015 3048 24053 3082
rect 24087 3048 24125 3082
rect 23943 3009 24125 3048
rect 23943 2975 23981 3009
rect 24015 2975 24053 3009
rect 24087 2975 24125 3009
rect 23943 2936 24125 2975
rect 23943 2902 23981 2936
rect 24015 2902 24053 2936
rect 24087 2902 24125 2936
rect 23943 2863 24125 2902
rect 23943 2829 23981 2863
rect 24015 2829 24053 2863
rect 24087 2829 24125 2863
rect 23943 2790 24125 2829
rect 23943 2756 23981 2790
rect 24015 2756 24053 2790
rect 24087 2756 24125 2790
rect 23943 2717 24125 2756
rect 23943 2683 23981 2717
rect 24015 2683 24053 2717
rect 24087 2683 24125 2717
rect 23943 2644 24125 2683
rect 23943 2610 23981 2644
rect 24015 2610 24053 2644
rect 24087 2610 24125 2644
rect 23943 2571 24125 2610
rect 23943 2537 23981 2571
rect 24015 2537 24053 2571
rect 24087 2537 24125 2571
rect 23943 2498 24125 2537
rect 23943 2464 23981 2498
rect 24015 2464 24053 2498
rect 24087 2464 24125 2498
rect 23943 2425 24125 2464
rect 23943 2391 23981 2425
rect 24015 2391 24053 2425
rect 24087 2391 24125 2425
rect 23943 2352 24125 2391
rect 23943 2318 23981 2352
rect 24015 2318 24053 2352
rect 24087 2318 24125 2352
rect 23943 2279 24125 2318
rect 23943 2245 23981 2279
rect 24015 2245 24053 2279
rect 24087 2245 24125 2279
rect 23943 2206 24125 2245
rect 23943 2172 23981 2206
rect 24015 2172 24053 2206
rect 24087 2172 24125 2206
rect 23943 2133 24125 2172
rect 23943 2099 23981 2133
rect 24015 2099 24053 2133
rect 24087 2099 24125 2133
rect 23943 2060 24125 2099
rect 23943 2026 23981 2060
rect 24015 2026 24053 2060
rect 24087 2026 24125 2060
rect 23943 1987 24125 2026
rect 23943 1953 23981 1987
rect 24015 1953 24053 1987
rect 24087 1953 24125 1987
rect 23943 1914 24125 1953
rect 11713 1899 12412 1904
rect 12464 1899 12486 1904
rect 12538 1899 12560 1904
rect 12612 1899 12634 1904
rect 12686 1899 12707 1904
rect 12759 1899 12780 1904
rect 12832 1899 13258 1904
rect 11713 1887 13258 1899
rect 8762 1863 11319 1869
tri 11198 1853 11208 1863 ne
rect 11208 1853 11319 1863
rect 1153 1811 1169 1845
rect 1203 1811 1241 1845
rect 1275 1811 1313 1845
rect 1347 1811 1385 1845
rect 1419 1811 1457 1845
rect 1491 1811 1529 1845
rect 1563 1811 1601 1845
rect 1635 1811 1651 1845
rect 1153 1772 1651 1811
rect 2098 1786 2104 1838
rect 2156 1786 2168 1838
rect 2220 1786 2232 1838
rect 2284 1786 2296 1838
rect 2348 1786 2360 1838
rect 2412 1786 2424 1838
rect 2476 1786 3010 1838
rect 1153 1738 1169 1772
rect 1203 1738 1241 1772
rect 1275 1738 1313 1772
rect 1347 1738 1385 1772
rect 1419 1738 1457 1772
rect 1491 1738 1529 1772
rect 1563 1738 1601 1772
rect 1635 1738 1651 1772
rect 1153 1699 1651 1738
rect 5031 1721 5071 1851
rect 7092 1847 8262 1853
rect 7092 1795 8146 1847
rect 8198 1795 8210 1847
rect 7092 1789 8262 1795
tri 11208 1789 11272 1853 ne
rect 11272 1789 11319 1853
tri 11272 1760 11301 1789 ne
rect 11301 1760 11319 1789
rect 11713 1866 12412 1887
rect 12464 1866 12486 1887
rect 12538 1866 12560 1887
rect 12612 1866 12634 1887
rect 12686 1866 12707 1887
rect 12759 1866 12780 1887
rect 12832 1866 13258 1887
tri 23135 1880 23169 1914 se
rect 23169 1880 23766 1914
tri 23766 1880 23800 1914 nw
rect 23943 1880 23981 1914
rect 24015 1880 24053 1914
rect 24087 1880 24125 1914
rect 11713 1832 11752 1866
rect 11786 1832 11825 1866
rect 11859 1832 11898 1866
rect 11932 1832 11971 1866
rect 12005 1832 12044 1866
rect 12078 1832 12117 1866
rect 12151 1832 12190 1866
rect 12224 1832 12263 1866
rect 12297 1832 12336 1866
rect 12370 1832 12409 1866
rect 12464 1835 12482 1866
rect 12538 1835 12555 1866
rect 12612 1835 12628 1866
rect 12686 1835 12701 1866
rect 12759 1835 12774 1866
rect 12832 1835 12847 1866
rect 12443 1832 12482 1835
rect 12516 1832 12555 1835
rect 12589 1832 12628 1835
rect 12662 1832 12701 1835
rect 12735 1832 12774 1835
rect 12808 1832 12847 1835
rect 12881 1832 12920 1866
rect 12954 1832 12993 1866
rect 13027 1832 13066 1866
rect 13100 1832 13139 1866
rect 13173 1832 13212 1866
rect 13246 1832 13258 1866
tri 23108 1853 23135 1880 se
rect 23135 1853 23727 1880
rect 11713 1823 13258 1832
rect 11713 1794 12412 1823
rect 12464 1794 12486 1823
rect 12538 1794 12560 1823
rect 12612 1794 12634 1823
rect 12686 1794 12707 1823
rect 12759 1794 12780 1823
rect 12832 1794 13258 1823
rect 11713 1760 11752 1794
rect 11786 1760 11825 1794
rect 11859 1760 11898 1794
rect 11932 1760 11971 1794
rect 12005 1760 12044 1794
rect 12078 1760 12117 1794
rect 12151 1760 12190 1794
rect 12224 1760 12263 1794
rect 12297 1760 12336 1794
rect 12370 1760 12409 1794
rect 12464 1771 12482 1794
rect 12538 1771 12555 1794
rect 12612 1771 12628 1794
rect 12686 1771 12701 1794
rect 12759 1771 12774 1794
rect 12832 1771 12847 1794
rect 12443 1760 12482 1771
rect 12516 1760 12555 1771
rect 12589 1760 12628 1771
rect 12662 1760 12701 1771
rect 12735 1760 12774 1771
rect 12808 1760 12847 1771
rect 12881 1760 12920 1794
rect 12954 1760 12993 1794
rect 13027 1760 13066 1794
rect 13100 1760 13139 1794
rect 13173 1760 13212 1794
rect 13246 1760 13258 1794
tri 11301 1754 11307 1760 ne
rect 11307 1754 13258 1760
rect 14251 1847 17609 1853
rect 14251 1795 17428 1847
rect 17480 1795 17492 1847
rect 17544 1795 17556 1847
rect 17608 1795 17609 1847
tri 23096 1841 23108 1853 se
rect 23108 1841 23727 1853
tri 23727 1841 23766 1880 nw
rect 23943 1841 24125 1880
tri 23062 1807 23096 1841 se
rect 23096 1807 23693 1841
tri 23693 1807 23727 1841 nw
rect 23943 1807 23981 1841
rect 24015 1807 24053 1841
rect 24087 1807 24125 1841
rect 14251 1735 17609 1795
tri 23023 1768 23062 1807 se
rect 23062 1768 23654 1807
tri 23654 1768 23693 1807 nw
rect 23943 1768 24125 1807
rect 1153 1665 1169 1699
rect 1203 1665 1241 1699
rect 1275 1665 1313 1699
rect 1347 1665 1385 1699
rect 1419 1665 1457 1699
rect 1491 1665 1529 1699
rect 1563 1665 1601 1699
rect 1635 1665 1651 1699
rect 14251 1683 17428 1735
rect 17480 1683 17492 1735
rect 17544 1683 17556 1735
rect 17608 1683 17609 1735
tri 22989 1734 23023 1768 se
rect 23023 1734 23620 1768
tri 23620 1734 23654 1768 nw
rect 23943 1734 23981 1768
rect 24015 1734 24053 1768
rect 24087 1734 24125 1768
tri 22977 1722 22989 1734 se
rect 22989 1722 23608 1734
tri 23608 1722 23620 1734 nw
rect 23943 1722 24125 1734
rect 14251 1673 17609 1683
tri 22932 1677 22977 1722 se
rect 22977 1677 23562 1722
tri 22931 1676 22932 1677 se
rect 22932 1676 23562 1677
tri 23562 1676 23608 1722 nw
tri 22928 1673 22931 1676 se
rect 22931 1673 23492 1676
rect 1153 1626 1651 1665
tri 22883 1628 22928 1673 se
rect 22928 1628 23492 1673
rect 1153 1592 1169 1626
rect 1203 1592 1241 1626
rect 1275 1592 1313 1626
rect 1347 1592 1385 1626
rect 1419 1592 1457 1626
rect 1491 1592 1529 1626
rect 1563 1592 1601 1626
rect 1635 1606 1651 1626
tri 1651 1606 1673 1628 sw
tri 22861 1606 22883 1628 se
rect 22883 1606 23492 1628
tri 23492 1606 23562 1676 nw
rect 1635 1592 1673 1606
rect 1153 1563 1673 1592
tri 1673 1563 1716 1606 sw
tri 22818 1563 22861 1606 se
rect 22861 1563 23386 1606
rect 1153 1557 1716 1563
tri 1716 1557 1722 1563 sw
tri 8416 1557 8422 1563 se
rect 8422 1557 10072 1563
rect 1153 1553 1722 1557
rect 1153 1519 1169 1553
rect 1203 1519 1241 1553
rect 1275 1519 1313 1553
rect 1347 1519 1385 1553
rect 1419 1519 1457 1553
rect 1491 1519 1529 1553
rect 1563 1519 1601 1553
rect 1635 1523 1722 1553
tri 1722 1523 1756 1557 sw
tri 8382 1523 8416 1557 se
rect 8416 1523 8434 1557
rect 8468 1523 8509 1557
rect 8543 1523 8584 1557
rect 8618 1523 8659 1557
rect 8693 1523 8734 1557
rect 8768 1523 8809 1557
rect 8843 1523 8884 1557
rect 8918 1523 8959 1557
rect 8993 1523 9034 1557
rect 9068 1523 9109 1557
rect 9143 1523 9184 1557
rect 9218 1523 9259 1557
rect 9293 1523 9334 1557
rect 9368 1523 9409 1557
rect 9443 1523 9484 1557
rect 9518 1523 9559 1557
rect 9593 1523 9634 1557
rect 9668 1523 9709 1557
rect 9743 1523 9784 1557
rect 9818 1523 9860 1557
rect 9894 1523 9936 1557
rect 9970 1523 10012 1557
rect 10046 1523 10072 1557
rect 1635 1519 1756 1523
rect 1153 1494 1756 1519
tri 1756 1494 1785 1523 sw
tri 8353 1494 8382 1523 se
rect 8382 1494 10072 1523
rect 1153 1486 1785 1494
tri 1785 1486 1793 1494 sw
tri 8345 1486 8353 1494 se
rect 8353 1486 10072 1494
rect 1153 1480 2997 1486
rect 1153 1446 1169 1480
rect 1203 1446 1241 1480
rect 1275 1446 1313 1480
rect 1347 1446 1385 1480
rect 1419 1446 1457 1480
rect 1491 1446 1529 1480
rect 1563 1446 1601 1480
rect 1635 1446 1683 1480
rect 1717 1446 1757 1480
rect 1791 1446 1831 1480
rect 1865 1446 1905 1480
rect 1939 1446 1979 1480
rect 2013 1446 2053 1480
rect 2087 1446 2127 1480
rect 2161 1446 2201 1480
rect 2235 1446 2276 1480
rect 2310 1446 2351 1480
rect 2385 1446 2426 1480
rect 2460 1446 2501 1480
rect 2535 1446 2576 1480
rect 2610 1446 2651 1480
rect 2685 1446 2726 1480
rect 2760 1446 2801 1480
rect 2835 1446 2876 1480
rect 2910 1446 2951 1480
rect 2985 1446 2997 1480
rect 1153 1408 2997 1446
rect 7105 1485 10072 1486
rect 7105 1480 8434 1485
rect 7105 1446 7117 1480
rect 7151 1446 7190 1480
rect 7224 1446 7263 1480
rect 7297 1446 7336 1480
rect 7370 1446 7409 1480
rect 7443 1446 7482 1480
rect 7516 1446 7555 1480
rect 7589 1446 7628 1480
rect 7662 1446 7701 1480
rect 7735 1446 7774 1480
rect 7808 1446 7847 1480
rect 7881 1446 7920 1480
rect 7954 1446 7993 1480
rect 8027 1446 8066 1480
rect 8100 1446 8140 1480
rect 8174 1446 8214 1480
rect 8248 1446 8288 1480
rect 8322 1446 8362 1480
rect 8396 1451 8434 1480
rect 8468 1451 8509 1485
rect 8543 1451 8584 1485
rect 8618 1451 8659 1485
rect 8693 1451 8734 1485
rect 8768 1451 8809 1485
rect 8843 1451 8884 1485
rect 8918 1451 8959 1485
rect 8993 1451 9034 1485
rect 9068 1451 9109 1485
rect 9143 1451 9184 1485
rect 9218 1451 9259 1485
rect 9293 1451 9334 1485
rect 9368 1451 9409 1485
rect 9443 1451 9484 1485
rect 9518 1451 9559 1485
rect 9593 1451 9634 1485
rect 9668 1451 9709 1485
rect 9743 1451 9784 1485
rect 9818 1451 9860 1485
rect 9894 1451 9936 1485
rect 9970 1451 10012 1485
rect 10046 1451 10072 1485
rect 8396 1446 10072 1451
rect 7105 1445 10072 1446
rect 12403 1562 12842 1563
rect 12403 1510 12409 1562
rect 12461 1510 12484 1562
rect 12536 1510 12559 1562
rect 12611 1510 12634 1562
rect 12686 1510 12709 1562
rect 12761 1510 12784 1562
rect 12836 1510 12842 1562
rect 12403 1498 12842 1510
tri 22755 1500 22818 1563 se
rect 22818 1500 23386 1563
tri 23386 1500 23492 1606 nw
rect 25689 1600 25765 1606
rect 25689 1548 25701 1600
rect 25753 1548 25765 1600
rect 25689 1525 25765 1548
rect 12403 1446 12409 1498
rect 12461 1446 12484 1498
rect 12536 1446 12559 1498
rect 12611 1446 12634 1498
rect 12686 1446 12709 1498
rect 12761 1446 12784 1498
rect 12836 1446 12842 1498
rect 12403 1445 12842 1446
rect 14481 1494 23277 1500
rect 14481 1460 14493 1494
rect 14527 1460 14566 1494
rect 14600 1460 14639 1494
rect 14673 1460 14712 1494
rect 14746 1460 14785 1494
rect 14819 1460 14858 1494
rect 14892 1460 14931 1494
rect 14965 1460 15004 1494
rect 15038 1460 15077 1494
rect 15111 1460 15150 1494
rect 15184 1460 15223 1494
rect 15257 1460 15296 1494
rect 15330 1460 15369 1494
rect 15403 1460 15442 1494
rect 15476 1460 15515 1494
rect 15549 1460 15588 1494
rect 15622 1460 15661 1494
rect 15695 1460 15734 1494
rect 7105 1422 8453 1445
tri 8453 1422 8476 1445 nw
rect 14481 1422 15734 1460
rect 3722 1414 6383 1421
rect 3722 1408 6805 1414
rect 1153 1374 1683 1408
rect 1717 1374 1757 1408
rect 1791 1374 1831 1408
rect 1865 1374 1905 1408
rect 1939 1374 1979 1408
rect 2013 1374 2053 1408
rect 2087 1374 2127 1408
rect 2161 1374 2201 1408
rect 2235 1374 2276 1408
rect 2310 1374 2351 1408
rect 2385 1374 2426 1408
rect 2460 1374 2501 1408
rect 2535 1374 2576 1408
rect 2610 1374 2651 1408
rect 2685 1374 2726 1408
rect 2760 1374 2801 1408
rect 2835 1374 2876 1408
rect 2910 1374 2951 1408
rect 2985 1374 2997 1408
rect 1153 1368 2997 1374
rect 3297 1390 6805 1408
rect 722 1331 840 1336
rect 722 1297 728 1331
rect 762 1297 840 1331
rect 3297 1338 4372 1390
rect 4424 1338 4436 1390
rect 4488 1338 6805 1390
rect 7105 1408 8419 1422
rect 7105 1374 7117 1408
rect 7151 1374 7190 1408
rect 7224 1374 7263 1408
rect 7297 1374 7336 1408
rect 7370 1374 7409 1408
rect 7443 1374 7482 1408
rect 7516 1374 7555 1408
rect 7589 1374 7628 1408
rect 7662 1374 7701 1408
rect 7735 1374 7774 1408
rect 7808 1374 7847 1408
rect 7881 1374 7920 1408
rect 7954 1374 7993 1408
rect 8027 1374 8066 1408
rect 8100 1374 8140 1408
rect 8174 1374 8214 1408
rect 8248 1374 8288 1408
rect 8322 1374 8362 1408
rect 8396 1388 8419 1408
tri 8419 1388 8453 1422 nw
rect 14481 1388 14493 1422
rect 14527 1388 14566 1422
rect 14600 1388 14639 1422
rect 14673 1388 14712 1422
rect 14746 1388 14785 1422
rect 14819 1388 14858 1422
rect 14892 1388 14931 1422
rect 14965 1388 15004 1422
rect 15038 1388 15077 1422
rect 15111 1388 15150 1422
rect 15184 1388 15223 1422
rect 15257 1388 15296 1422
rect 15330 1388 15369 1422
rect 15403 1388 15442 1422
rect 15476 1388 15515 1422
rect 15549 1388 15588 1422
rect 15622 1388 15661 1422
rect 15695 1388 15734 1422
rect 8396 1374 8408 1388
tri 8408 1377 8419 1388 nw
rect 7105 1368 8408 1374
rect 3297 1321 6805 1338
rect 14481 1350 15734 1388
rect 722 1263 800 1297
rect 834 1263 840 1297
rect 722 1259 840 1263
rect 722 1225 728 1259
rect 762 1225 840 1259
rect 722 1224 840 1225
rect 722 1190 800 1224
rect 834 1190 840 1224
rect 722 1187 840 1190
rect 722 1153 728 1187
rect 762 1153 840 1187
rect 722 1151 840 1153
rect 722 1117 800 1151
rect 834 1117 840 1151
rect 722 1115 840 1117
rect 722 1081 728 1115
rect 762 1081 840 1115
rect 722 1078 840 1081
rect 722 1044 800 1078
rect 834 1044 840 1078
rect 14481 1316 14493 1350
rect 14527 1316 14566 1350
rect 14600 1316 14639 1350
rect 14673 1316 14712 1350
rect 14746 1316 14785 1350
rect 14819 1316 14858 1350
rect 14892 1316 14931 1350
rect 14965 1316 15004 1350
rect 15038 1316 15077 1350
rect 15111 1316 15150 1350
rect 15184 1316 15223 1350
rect 15257 1316 15296 1350
rect 15330 1316 15369 1350
rect 15403 1316 15442 1350
rect 15476 1316 15515 1350
rect 15549 1316 15588 1350
rect 15622 1316 15661 1350
rect 15695 1316 15734 1350
rect 14481 1278 15734 1316
rect 14481 1244 14493 1278
rect 14527 1244 14566 1278
rect 14600 1244 14639 1278
rect 14673 1244 14712 1278
rect 14746 1244 14785 1278
rect 14819 1244 14858 1278
rect 14892 1244 14931 1278
rect 14965 1244 15004 1278
rect 15038 1244 15077 1278
rect 15111 1244 15150 1278
rect 15184 1244 15223 1278
rect 15257 1244 15296 1278
rect 15330 1244 15369 1278
rect 15403 1244 15442 1278
rect 15476 1244 15515 1278
rect 15549 1244 15588 1278
rect 15622 1244 15661 1278
rect 15695 1244 15734 1278
rect 14481 1206 15734 1244
rect 14481 1172 14493 1206
rect 14527 1172 14566 1206
rect 14600 1172 14639 1206
rect 14673 1172 14712 1206
rect 14746 1172 14785 1206
rect 14819 1172 14858 1206
rect 14892 1172 14931 1206
rect 14965 1172 15004 1206
rect 15038 1172 15077 1206
rect 15111 1172 15150 1206
rect 15184 1172 15223 1206
rect 15257 1172 15296 1206
rect 15330 1172 15369 1206
rect 15403 1172 15442 1206
rect 15476 1172 15515 1206
rect 15549 1172 15588 1206
rect 15622 1172 15661 1206
rect 15695 1172 15734 1206
rect 23040 1391 23277 1494
tri 23277 1391 23386 1500 nw
rect 25689 1473 25701 1525
rect 25753 1473 25765 1525
rect 25689 1449 25765 1473
rect 25689 1397 25701 1449
rect 25753 1397 25765 1449
rect 25689 1391 25765 1397
rect 23040 1213 23099 1391
tri 23099 1213 23277 1391 nw
rect 23040 1172 23052 1213
rect 14481 1166 23052 1172
tri 23052 1166 23099 1213 nw
rect 14481 1146 14721 1166
tri 14721 1146 14741 1166 nw
rect 14481 1134 14599 1146
rect 14481 1100 14487 1134
rect 14521 1100 14559 1134
rect 14593 1100 14599 1134
rect 14481 1053 14599 1100
rect 722 1043 840 1044
rect 722 1009 728 1043
rect 762 1021 840 1043
tri 840 1021 865 1046 sw
tri 14456 1021 14481 1046 se
rect 14481 1021 14559 1053
rect 762 1019 14559 1021
rect 14593 1019 14599 1053
tri 14599 1024 14721 1146 nw
rect 762 1009 14599 1019
rect 722 1005 14599 1009
rect 722 971 800 1005
rect 834 971 873 1005
rect 907 971 946 1005
rect 980 971 1019 1005
rect 1053 971 1092 1005
rect 1126 971 1165 1005
rect 1199 971 1238 1005
rect 1272 971 1311 1005
rect 722 933 1311 971
rect 722 899 766 933
rect 800 899 839 933
rect 873 899 912 933
rect 946 899 985 933
rect 1019 899 1057 933
rect 1091 899 1129 933
rect 1163 899 1201 933
rect 1235 899 1273 933
rect 1307 899 1311 933
rect 14483 971 14487 1005
rect 14521 971 14599 1005
rect 14483 937 14559 971
rect 14593 937 14599 971
tri 23528 950 23571 993 se
rect 23571 969 23577 1213
rect 23757 1033 23763 1213
rect 23693 969 23763 1033
rect 23571 957 23763 969
rect 23571 950 23577 957
rect 14483 899 14599 937
rect 722 893 14599 899
rect 20481 944 23577 950
rect 23629 944 23763 957
rect 20481 910 20551 944
rect 20585 910 20625 944
rect 20659 910 20699 944
rect 20733 910 20773 944
rect 20807 910 20847 944
rect 20881 910 20921 944
rect 20955 910 20995 944
rect 21029 910 21069 944
rect 21103 910 21143 944
rect 21177 910 21217 944
rect 21251 910 21291 944
rect 21325 910 21365 944
rect 21399 910 21439 944
rect 21473 910 21513 944
rect 21547 910 21587 944
rect 21621 910 21661 944
rect 21695 910 21735 944
rect 21769 910 21809 944
rect 21843 910 21883 944
rect 21917 910 21957 944
rect 21991 910 22031 944
rect 22065 910 22105 944
rect 22139 910 22179 944
rect 22213 910 22253 944
rect 22287 910 22327 944
rect 22361 910 22401 944
rect 22435 910 22475 944
rect 22509 910 22549 944
rect 22583 910 22622 944
rect 22656 910 22695 944
rect 22729 910 22768 944
rect 22802 910 22841 944
rect 22875 910 22914 944
rect 22948 910 22987 944
rect 23021 910 23060 944
rect 23094 910 23133 944
rect 23167 910 23206 944
rect 23240 910 23279 944
rect 23313 910 23352 944
rect 23386 910 23425 944
rect 23459 910 23498 944
rect 23532 910 23571 944
rect 23629 910 23644 944
rect 23678 910 23717 944
rect 23751 910 23763 944
rect 20481 905 23577 910
rect 23629 905 23763 910
rect 27009 1172 27372 1192
rect 27009 1120 27015 1172
rect 27067 1120 27090 1172
rect 27142 1120 27165 1172
rect 27217 1120 27240 1172
rect 27292 1120 27314 1172
rect 27366 1120 27372 1172
rect 27009 1108 27372 1120
rect 27009 1056 27015 1108
rect 27067 1056 27090 1108
rect 27142 1056 27165 1108
rect 27217 1056 27240 1108
rect 27292 1056 27314 1108
rect 27366 1056 27372 1108
rect 27009 1044 27372 1056
rect 27009 992 27015 1044
rect 27067 992 27090 1044
rect 27142 992 27165 1044
rect 27217 992 27240 1044
rect 27292 992 27314 1044
rect 27366 992 27372 1044
rect 27009 980 27372 992
rect 27009 928 27015 980
rect 27067 928 27090 980
rect 27142 928 27165 980
rect 27217 928 27240 980
rect 27292 928 27314 980
rect 27366 928 27372 980
rect 27009 908 27372 928
rect 304 821 310 855
rect 344 821 382 855
rect 416 821 422 855
rect 20481 872 23763 905
rect 20481 838 20551 872
rect 20585 838 20625 872
rect 20659 838 20699 872
rect 20733 838 20773 872
rect 20807 838 20847 872
rect 20881 838 20921 872
rect 20955 838 20995 872
rect 21029 838 21069 872
rect 21103 838 21143 872
rect 21177 838 21217 872
rect 21251 838 21291 872
rect 21325 838 21365 872
rect 21399 838 21439 872
rect 21473 838 21513 872
rect 21547 838 21587 872
rect 21621 838 21661 872
rect 21695 838 21735 872
rect 21769 838 21809 872
rect 21843 838 21883 872
rect 21917 838 21957 872
rect 21991 838 22031 872
rect 22065 838 22105 872
rect 22139 838 22179 872
rect 22213 838 22253 872
rect 22287 838 22327 872
rect 22361 838 22401 872
rect 22435 838 22475 872
rect 22509 838 22549 872
rect 22583 838 22622 872
rect 22656 838 22695 872
rect 22729 838 22768 872
rect 22802 838 22841 872
rect 22875 838 22914 872
rect 22948 838 22987 872
rect 23021 838 23060 872
rect 23094 838 23133 872
rect 23167 838 23206 872
rect 23240 838 23279 872
rect 23313 838 23352 872
rect 23386 838 23425 872
rect 23459 838 23498 872
rect 23532 838 23571 872
rect 23605 838 23644 872
rect 23678 838 23717 872
rect 23751 838 23763 872
rect 20481 832 23763 838
rect 304 782 422 821
rect 304 748 310 782
rect 344 748 382 782
rect 416 748 422 782
rect 304 709 422 748
rect 304 675 310 709
rect 344 675 382 709
rect 416 675 422 709
rect 304 636 422 675
rect 304 602 310 636
rect 344 602 382 636
rect 416 602 422 636
rect 304 563 422 602
rect 304 529 310 563
rect 344 529 382 563
rect 416 529 422 563
tri 14226 531 14251 556 se
rect 304 490 422 529
rect 304 456 310 490
rect 344 456 382 490
rect 416 456 422 490
rect 304 417 422 456
rect 304 383 310 417
rect 344 383 382 417
rect 416 383 422 417
rect 753 413 14371 531
rect 304 344 422 383
rect 304 310 310 344
rect 344 310 382 344
rect 416 310 422 344
rect 304 271 422 310
rect 304 237 310 271
rect 344 237 382 271
rect 416 237 422 271
rect 304 198 422 237
rect 304 164 310 198
rect 344 164 382 198
rect 416 164 422 198
tri 279 113 304 138 se
rect 304 113 422 164
tri 422 113 447 138 sw
rect 279 49 447 113
tri 21442 -1883 21467 -1858 se
rect 21467 -1883 21531 -1858
rect 21185 -1889 21531 -1883
rect 21185 -1923 21197 -1889
rect 21231 -1923 21269 -1889
rect 21303 -1923 21341 -1889
rect 21375 -1923 21413 -1889
rect 21447 -1923 21485 -1889
rect 21519 -1923 21531 -1889
rect 21185 -1929 21531 -1923
<< via1 >>
rect 23743 13258 23795 13310
rect 23743 13194 23795 13246
rect 24229 10939 24281 10991
rect 24229 10875 24281 10927
rect 24741 10905 24793 10957
rect 24805 10905 24857 10957
rect 27440 10905 27492 10957
rect 27504 10905 27556 10957
rect 25300 10812 25352 10864
rect 25364 10812 25416 10864
rect 25672 10812 25724 10864
rect 25736 10812 25788 10864
rect 25999 10820 26051 10872
rect 26091 10820 26143 10872
rect 26183 10820 26235 10872
rect 26275 10820 26327 10872
rect 26367 10820 26419 10872
rect 25262 10504 25314 10556
rect 25326 10504 25378 10556
rect 25711 10504 25763 10556
rect 25775 10504 25827 10556
rect 27505 10504 27557 10556
rect 27569 10504 27621 10556
rect 25762 10392 25814 10444
rect 25762 10327 25814 10379
rect 25762 10262 25814 10314
rect 25762 10196 25814 10248
rect 24195 10071 24247 10123
rect 24259 10071 24311 10123
rect 25408 10072 25460 10124
rect 25472 10072 25524 10124
rect 28069 10072 28121 10124
rect 28133 10072 28185 10124
rect 20702 9823 20754 9875
rect 20768 9823 20820 9875
rect 20834 9823 20886 9875
rect 20900 9823 20952 9875
rect 20966 9823 21018 9875
rect 21032 9823 21084 9875
rect 21097 9823 21149 9875
rect 21162 9823 21214 9875
rect 21227 9823 21279 9875
rect 21292 9823 21344 9875
rect 21357 9823 21409 9875
rect 20702 9759 20754 9811
rect 20768 9759 20820 9811
rect 20834 9759 20886 9811
rect 20900 9759 20952 9811
rect 20966 9759 21018 9811
rect 21032 9759 21084 9811
rect 21097 9759 21149 9811
rect 21162 9759 21214 9811
rect 21227 9759 21279 9811
rect 21292 9759 21344 9811
rect 21357 9759 21409 9811
rect 17024 9635 17076 9687
rect 17090 9635 17142 9687
rect 17156 9635 17208 9687
rect 17222 9635 17274 9687
rect 17288 9635 17340 9687
rect 17354 9635 17406 9687
rect 17420 9635 17472 9687
rect 17486 9635 17538 9687
rect 17552 9635 17604 9687
rect 17618 9635 17670 9687
rect 17684 9635 17736 9687
rect 17750 9635 17802 9687
rect 17816 9635 17868 9687
rect 17882 9635 17934 9687
rect 17948 9635 18000 9687
rect 18014 9635 18066 9687
rect 18080 9635 18132 9687
rect 18146 9635 18198 9687
rect 18212 9635 18264 9687
rect 18278 9635 18330 9687
rect 18344 9635 18396 9687
rect 18410 9635 18462 9687
rect 18476 9635 18528 9687
rect 18542 9635 18594 9687
rect 18607 9635 18659 9687
rect 18672 9635 18724 9687
rect 18737 9635 18789 9687
rect 18802 9635 18854 9687
rect 18867 9635 18919 9687
rect 18932 9635 18984 9687
rect 18997 9635 19049 9687
rect 19062 9635 19114 9687
rect 19127 9635 19179 9687
rect 19192 9635 19244 9687
rect 19257 9635 19309 9687
rect 17024 9571 17076 9623
rect 17090 9571 17142 9623
rect 17156 9571 17208 9623
rect 17222 9571 17274 9623
rect 17288 9571 17340 9623
rect 17354 9571 17406 9623
rect 17420 9571 17472 9623
rect 17486 9571 17538 9623
rect 17552 9571 17604 9623
rect 17618 9571 17670 9623
rect 17684 9571 17736 9623
rect 17750 9571 17802 9623
rect 17816 9571 17868 9623
rect 17882 9571 17934 9623
rect 17948 9571 18000 9623
rect 18014 9571 18066 9623
rect 18080 9571 18132 9623
rect 18146 9571 18198 9623
rect 18212 9571 18264 9623
rect 18278 9571 18330 9623
rect 18344 9571 18396 9623
rect 18410 9571 18462 9623
rect 18476 9571 18528 9623
rect 18542 9571 18594 9623
rect 18607 9571 18659 9623
rect 18672 9571 18724 9623
rect 18737 9571 18789 9623
rect 18802 9571 18854 9623
rect 18867 9571 18919 9623
rect 18932 9571 18984 9623
rect 18997 9571 19049 9623
rect 19062 9571 19114 9623
rect 19127 9571 19179 9623
rect 19192 9571 19244 9623
rect 19257 9571 19309 9623
rect 25511 9922 25563 9974
rect 25575 9922 25627 9974
rect 27664 9922 27716 9974
rect 27728 9922 27780 9974
rect 25247 9727 25299 9779
rect 25311 9727 25363 9779
rect 27312 9728 27364 9780
rect 27376 9728 27428 9780
rect 27342 9494 27394 9546
rect 27342 9430 27394 9482
rect 27922 9424 27974 9476
rect 27986 9424 28038 9476
rect 17029 9017 17081 9069
rect 17095 9017 17147 9069
rect 17161 9017 17213 9069
rect 17227 9017 17279 9069
rect 17293 9017 17345 9069
rect 17359 9017 17411 9069
rect 17425 9017 17477 9069
rect 17491 9017 17543 9069
rect 17557 9017 17609 9069
rect 17623 9017 17675 9069
rect 17689 9017 17741 9069
rect 17755 9017 17807 9069
rect 17821 9017 17873 9069
rect 17887 9017 17939 9069
rect 17953 9017 18005 9069
rect 18019 9017 18071 9069
rect 18085 9017 18137 9069
rect 18151 9017 18203 9069
rect 18217 9017 18269 9069
rect 18282 9017 18334 9069
rect 18347 9017 18399 9069
rect 18412 9017 18464 9069
rect 18477 9017 18529 9069
rect 18542 9017 18594 9069
rect 18607 9017 18659 9069
rect 18672 9017 18724 9069
rect 18737 9017 18789 9069
rect 18802 9017 18854 9069
rect 18867 9017 18919 9069
rect 18932 9017 18984 9069
rect 18997 9017 19049 9069
rect 19062 9017 19114 9069
rect 19127 9017 19179 9069
rect 19192 9017 19244 9069
rect 19257 9017 19309 9069
rect 17029 8953 17081 9005
rect 17095 8953 17147 9005
rect 17161 8953 17213 9005
rect 17227 8953 17279 9005
rect 17293 8953 17345 9005
rect 17359 8953 17411 9005
rect 17425 8953 17477 9005
rect 17491 8953 17543 9005
rect 17557 8953 17609 9005
rect 17623 8953 17675 9005
rect 17689 8953 17741 9005
rect 17755 8953 17807 9005
rect 17821 8953 17873 9005
rect 17887 8953 17939 9005
rect 17953 8953 18005 9005
rect 18019 8953 18071 9005
rect 18085 8953 18137 9005
rect 18151 8953 18203 9005
rect 18217 8953 18269 9005
rect 18282 8953 18334 9005
rect 18347 8953 18399 9005
rect 18412 8953 18464 9005
rect 18477 8953 18529 9005
rect 18542 8953 18594 9005
rect 18607 8953 18659 9005
rect 18672 8953 18724 9005
rect 18737 8953 18789 9005
rect 18802 8953 18854 9005
rect 18867 8953 18919 9005
rect 18932 8953 18984 9005
rect 18997 8953 19049 9005
rect 19062 8953 19114 9005
rect 19127 8953 19179 9005
rect 19192 8953 19244 9005
rect 19257 8953 19309 9005
rect 20702 8953 20754 9005
rect 20768 8953 20820 9005
rect 20834 8953 20886 9005
rect 20900 8953 20952 9005
rect 20966 8953 21018 9005
rect 21032 8953 21084 9005
rect 21097 8953 21149 9005
rect 21162 8953 21214 9005
rect 21227 8953 21279 9005
rect 21292 8953 21344 9005
rect 21357 8953 21409 9005
rect 20702 8889 20754 8941
rect 20768 8889 20820 8941
rect 20834 8889 20886 8941
rect 20900 8889 20952 8941
rect 20966 8889 21018 8941
rect 21032 8889 21084 8941
rect 21097 8889 21149 8941
rect 21162 8889 21214 8941
rect 21227 8889 21279 8941
rect 21292 8889 21344 8941
rect 21357 8889 21409 8941
rect 20702 8825 20754 8877
rect 20768 8825 20820 8877
rect 20834 8825 20886 8877
rect 20900 8825 20952 8877
rect 20966 8825 21018 8877
rect 21032 8825 21084 8877
rect 21097 8825 21149 8877
rect 21162 8825 21214 8877
rect 21227 8825 21279 8877
rect 21292 8825 21344 8877
rect 21357 8825 21409 8877
rect 17029 8762 17081 8814
rect 17095 8762 17147 8814
rect 17161 8762 17213 8814
rect 17227 8762 17279 8814
rect 17293 8762 17345 8814
rect 17359 8762 17411 8814
rect 17425 8762 17477 8814
rect 17491 8762 17543 8814
rect 17557 8762 17609 8814
rect 17623 8762 17675 8814
rect 17689 8762 17741 8814
rect 17755 8762 17807 8814
rect 17821 8762 17873 8814
rect 17887 8762 17939 8814
rect 17953 8762 18005 8814
rect 18019 8762 18071 8814
rect 18085 8762 18137 8814
rect 18151 8762 18203 8814
rect 18217 8762 18269 8814
rect 18282 8762 18334 8814
rect 18347 8762 18399 8814
rect 18412 8762 18464 8814
rect 18477 8762 18529 8814
rect 18542 8762 18594 8814
rect 18607 8762 18659 8814
rect 18672 8762 18724 8814
rect 18737 8762 18789 8814
rect 18802 8762 18854 8814
rect 18867 8762 18919 8814
rect 18932 8762 18984 8814
rect 18997 8762 19049 8814
rect 19062 8762 19114 8814
rect 19127 8762 19179 8814
rect 19192 8762 19244 8814
rect 19257 8762 19309 8814
rect 17029 8698 17081 8750
rect 17095 8698 17147 8750
rect 17161 8698 17213 8750
rect 17227 8698 17279 8750
rect 17293 8698 17345 8750
rect 17359 8698 17411 8750
rect 17425 8698 17477 8750
rect 17491 8698 17543 8750
rect 17557 8698 17609 8750
rect 17623 8698 17675 8750
rect 17689 8698 17741 8750
rect 17755 8698 17807 8750
rect 17821 8698 17873 8750
rect 17887 8698 17939 8750
rect 17953 8698 18005 8750
rect 18019 8698 18071 8750
rect 18085 8698 18137 8750
rect 18151 8698 18203 8750
rect 18217 8698 18269 8750
rect 18282 8698 18334 8750
rect 18347 8698 18399 8750
rect 18412 8698 18464 8750
rect 18477 8698 18529 8750
rect 18542 8698 18594 8750
rect 18607 8698 18659 8750
rect 18672 8698 18724 8750
rect 18737 8698 18789 8750
rect 18802 8698 18854 8750
rect 18867 8698 18919 8750
rect 18932 8698 18984 8750
rect 18997 8698 19049 8750
rect 19062 8698 19114 8750
rect 19127 8698 19179 8750
rect 19192 8698 19244 8750
rect 19257 8698 19309 8750
rect 17029 8634 17081 8686
rect 17095 8634 17147 8686
rect 17161 8634 17213 8686
rect 17227 8634 17279 8686
rect 17293 8634 17345 8686
rect 17359 8634 17411 8686
rect 17425 8634 17477 8686
rect 17491 8634 17543 8686
rect 17557 8634 17609 8686
rect 17623 8634 17675 8686
rect 17689 8634 17741 8686
rect 17755 8634 17807 8686
rect 17821 8634 17873 8686
rect 17887 8634 17939 8686
rect 17953 8634 18005 8686
rect 18019 8634 18071 8686
rect 18085 8634 18137 8686
rect 18151 8634 18203 8686
rect 18217 8634 18269 8686
rect 18282 8634 18334 8686
rect 18347 8634 18399 8686
rect 18412 8634 18464 8686
rect 18477 8634 18529 8686
rect 18542 8634 18594 8686
rect 18607 8634 18659 8686
rect 18672 8634 18724 8686
rect 18737 8634 18789 8686
rect 18802 8634 18854 8686
rect 18867 8634 18919 8686
rect 18932 8634 18984 8686
rect 18997 8634 19049 8686
rect 19062 8634 19114 8686
rect 19127 8634 19179 8686
rect 19192 8634 19244 8686
rect 19257 8634 19309 8686
rect 20702 8761 20754 8813
rect 20768 8761 20820 8813
rect 20834 8761 20886 8813
rect 20900 8761 20952 8813
rect 20966 8761 21018 8813
rect 21032 8761 21084 8813
rect 21097 8761 21149 8813
rect 21162 8761 21214 8813
rect 21227 8761 21279 8813
rect 21292 8761 21344 8813
rect 21357 8761 21409 8813
rect 20702 8697 20754 8749
rect 20768 8697 20820 8749
rect 20834 8697 20886 8749
rect 20900 8697 20952 8749
rect 20966 8697 21018 8749
rect 21032 8697 21084 8749
rect 21097 8697 21149 8749
rect 21162 8697 21214 8749
rect 21227 8697 21279 8749
rect 21292 8697 21344 8749
rect 21357 8697 21409 8749
rect 20702 8633 20754 8685
rect 20768 8633 20820 8685
rect 20834 8633 20886 8685
rect 20900 8633 20952 8685
rect 20966 8633 21018 8685
rect 21032 8633 21084 8685
rect 21097 8633 21149 8685
rect 21162 8633 21214 8685
rect 21227 8633 21279 8685
rect 21292 8633 21344 8685
rect 21357 8633 21409 8685
rect 20509 8523 20561 8575
rect 20573 8523 20625 8575
rect 17029 8443 17081 8495
rect 17095 8443 17147 8495
rect 17161 8443 17213 8495
rect 17227 8443 17279 8495
rect 17293 8443 17345 8495
rect 17359 8443 17411 8495
rect 17425 8443 17477 8495
rect 17491 8443 17543 8495
rect 17557 8443 17609 8495
rect 17623 8443 17675 8495
rect 17689 8443 17741 8495
rect 17755 8443 17807 8495
rect 17821 8443 17873 8495
rect 17887 8443 17939 8495
rect 17953 8443 18005 8495
rect 18019 8443 18071 8495
rect 18085 8443 18137 8495
rect 18151 8443 18203 8495
rect 18217 8443 18269 8495
rect 18282 8443 18334 8495
rect 18347 8443 18399 8495
rect 18412 8443 18464 8495
rect 18477 8443 18529 8495
rect 18542 8443 18594 8495
rect 18607 8443 18659 8495
rect 18672 8443 18724 8495
rect 18737 8443 18789 8495
rect 18802 8443 18854 8495
rect 18867 8443 18919 8495
rect 18932 8443 18984 8495
rect 18997 8443 19049 8495
rect 19062 8443 19114 8495
rect 19127 8443 19179 8495
rect 19192 8443 19244 8495
rect 19257 8443 19309 8495
rect 17029 8379 17081 8431
rect 17095 8379 17147 8431
rect 17161 8379 17213 8431
rect 17227 8379 17279 8431
rect 17293 8379 17345 8431
rect 17359 8379 17411 8431
rect 17425 8379 17477 8431
rect 17491 8379 17543 8431
rect 17557 8379 17609 8431
rect 17623 8379 17675 8431
rect 17689 8379 17741 8431
rect 17755 8379 17807 8431
rect 17821 8379 17873 8431
rect 17887 8379 17939 8431
rect 17953 8379 18005 8431
rect 18019 8379 18071 8431
rect 18085 8379 18137 8431
rect 18151 8379 18203 8431
rect 18217 8379 18269 8431
rect 18282 8379 18334 8431
rect 18347 8379 18399 8431
rect 18412 8379 18464 8431
rect 18477 8379 18529 8431
rect 18542 8379 18594 8431
rect 18607 8379 18659 8431
rect 18672 8379 18724 8431
rect 18737 8379 18789 8431
rect 18802 8379 18854 8431
rect 18867 8379 18919 8431
rect 18932 8379 18984 8431
rect 18997 8379 19049 8431
rect 19062 8379 19114 8431
rect 19127 8379 19179 8431
rect 19192 8379 19244 8431
rect 19257 8379 19309 8431
rect 17029 8315 17081 8367
rect 17095 8315 17147 8367
rect 17161 8315 17213 8367
rect 17227 8315 17279 8367
rect 17293 8315 17345 8367
rect 17359 8315 17411 8367
rect 17425 8315 17477 8367
rect 17491 8315 17543 8367
rect 17557 8315 17609 8367
rect 17623 8315 17675 8367
rect 17689 8315 17741 8367
rect 17755 8315 17807 8367
rect 17821 8315 17873 8367
rect 17887 8315 17939 8367
rect 17953 8315 18005 8367
rect 18019 8315 18071 8367
rect 18085 8315 18137 8367
rect 18151 8315 18203 8367
rect 18217 8315 18269 8367
rect 18282 8315 18334 8367
rect 18347 8315 18399 8367
rect 18412 8315 18464 8367
rect 18477 8315 18529 8367
rect 18542 8315 18594 8367
rect 18607 8315 18659 8367
rect 18672 8315 18724 8367
rect 18737 8315 18789 8367
rect 18802 8315 18854 8367
rect 18867 8315 18919 8367
rect 18932 8315 18984 8367
rect 18997 8315 19049 8367
rect 19062 8315 19114 8367
rect 19127 8315 19179 8367
rect 19192 8315 19244 8367
rect 19257 8315 19309 8367
rect 20702 8443 20754 8495
rect 20768 8443 20820 8495
rect 20834 8443 20886 8495
rect 20900 8443 20952 8495
rect 20966 8443 21018 8495
rect 21032 8443 21084 8495
rect 21097 8443 21149 8495
rect 21162 8443 21214 8495
rect 21227 8443 21279 8495
rect 21292 8443 21344 8495
rect 21357 8443 21409 8495
rect 20702 8379 20754 8431
rect 20768 8379 20820 8431
rect 20834 8379 20886 8431
rect 20900 8379 20952 8431
rect 20966 8379 21018 8431
rect 21032 8379 21084 8431
rect 21097 8379 21149 8431
rect 21162 8379 21214 8431
rect 21227 8379 21279 8431
rect 21292 8379 21344 8431
rect 21357 8379 21409 8431
rect 20702 8315 20754 8367
rect 20768 8315 20820 8367
rect 20834 8315 20886 8367
rect 20900 8315 20952 8367
rect 20966 8315 21018 8367
rect 21032 8315 21084 8367
rect 21097 8315 21149 8367
rect 21162 8315 21214 8367
rect 21227 8315 21279 8367
rect 21292 8315 21344 8367
rect 21357 8315 21409 8367
rect 17029 8179 17081 8231
rect 17095 8179 17147 8231
rect 17161 8179 17213 8231
rect 17227 8179 17279 8231
rect 17293 8179 17345 8231
rect 17359 8179 17411 8231
rect 17425 8179 17477 8231
rect 17491 8179 17543 8231
rect 17557 8179 17609 8231
rect 17623 8179 17675 8231
rect 17689 8179 17741 8231
rect 17755 8179 17807 8231
rect 17821 8179 17873 8231
rect 17887 8179 17939 8231
rect 17953 8179 18005 8231
rect 18019 8179 18071 8231
rect 18085 8179 18137 8231
rect 18151 8179 18203 8231
rect 18217 8179 18269 8231
rect 18282 8179 18334 8231
rect 18347 8179 18399 8231
rect 18412 8179 18464 8231
rect 18477 8179 18529 8231
rect 18542 8179 18594 8231
rect 18607 8179 18659 8231
rect 18672 8179 18724 8231
rect 18737 8179 18789 8231
rect 18802 8179 18854 8231
rect 18867 8179 18919 8231
rect 18932 8179 18984 8231
rect 18997 8179 19049 8231
rect 19062 8179 19114 8231
rect 19127 8179 19179 8231
rect 19192 8179 19244 8231
rect 19257 8179 19309 8231
rect 17029 8115 17081 8167
rect 17095 8115 17147 8167
rect 17161 8115 17213 8167
rect 17227 8115 17279 8167
rect 17293 8115 17345 8167
rect 17359 8115 17411 8167
rect 17425 8115 17477 8167
rect 17491 8115 17543 8167
rect 17557 8115 17609 8167
rect 17623 8115 17675 8167
rect 17689 8115 17741 8167
rect 17755 8115 17807 8167
rect 17821 8115 17873 8167
rect 17887 8115 17939 8167
rect 17953 8115 18005 8167
rect 18019 8115 18071 8167
rect 18085 8115 18137 8167
rect 18151 8115 18203 8167
rect 18217 8115 18269 8167
rect 18282 8115 18334 8167
rect 18347 8115 18399 8167
rect 18412 8115 18464 8167
rect 18477 8115 18529 8167
rect 18542 8115 18594 8167
rect 18607 8115 18659 8167
rect 18672 8115 18724 8167
rect 18737 8115 18789 8167
rect 18802 8115 18854 8167
rect 18867 8115 18919 8167
rect 18932 8115 18984 8167
rect 18997 8115 19049 8167
rect 19062 8115 19114 8167
rect 19127 8115 19179 8167
rect 19192 8115 19244 8167
rect 19257 8115 19309 8167
rect 17029 8051 17081 8103
rect 17095 8051 17147 8103
rect 17161 8051 17213 8103
rect 17227 8051 17279 8103
rect 17293 8051 17345 8103
rect 17359 8051 17411 8103
rect 17425 8051 17477 8103
rect 17491 8051 17543 8103
rect 17557 8051 17609 8103
rect 17623 8051 17675 8103
rect 17689 8051 17741 8103
rect 17755 8051 17807 8103
rect 17821 8051 17873 8103
rect 17887 8051 17939 8103
rect 17953 8051 18005 8103
rect 18019 8051 18071 8103
rect 18085 8051 18137 8103
rect 18151 8051 18203 8103
rect 18217 8051 18269 8103
rect 18282 8051 18334 8103
rect 18347 8051 18399 8103
rect 18412 8051 18464 8103
rect 18477 8051 18529 8103
rect 18542 8051 18594 8103
rect 18607 8051 18659 8103
rect 18672 8051 18724 8103
rect 18737 8051 18789 8103
rect 18802 8051 18854 8103
rect 18867 8051 18919 8103
rect 18932 8051 18984 8103
rect 18997 8051 19049 8103
rect 19062 8051 19114 8103
rect 19127 8051 19179 8103
rect 19192 8051 19244 8103
rect 19257 8051 19309 8103
rect 20702 8179 20754 8231
rect 20768 8179 20820 8231
rect 20834 8179 20886 8231
rect 20900 8179 20952 8231
rect 20966 8179 21018 8231
rect 21032 8179 21084 8231
rect 21097 8179 21149 8231
rect 21162 8179 21214 8231
rect 21227 8179 21279 8231
rect 21292 8179 21344 8231
rect 21357 8179 21409 8231
rect 20702 8115 20754 8167
rect 20768 8115 20820 8167
rect 20834 8115 20886 8167
rect 20900 8115 20952 8167
rect 20966 8115 21018 8167
rect 21032 8115 21084 8167
rect 21097 8115 21149 8167
rect 21162 8115 21214 8167
rect 21227 8115 21279 8167
rect 21292 8115 21344 8167
rect 21357 8115 21409 8167
rect 20702 8051 20754 8103
rect 20768 8051 20820 8103
rect 20834 8051 20886 8103
rect 20900 8051 20952 8103
rect 20966 8051 21018 8103
rect 21032 8051 21084 8103
rect 21097 8051 21149 8103
rect 21162 8051 21214 8103
rect 21227 8051 21279 8103
rect 21292 8051 21344 8103
rect 21357 8051 21409 8103
rect 17029 7915 17081 7967
rect 17095 7915 17147 7967
rect 17161 7915 17213 7967
rect 17227 7915 17279 7967
rect 17293 7915 17345 7967
rect 17359 7915 17411 7967
rect 17425 7915 17477 7967
rect 17491 7915 17543 7967
rect 17557 7915 17609 7967
rect 17623 7915 17675 7967
rect 17689 7915 17741 7967
rect 17755 7915 17807 7967
rect 17821 7915 17873 7967
rect 17887 7915 17939 7967
rect 17953 7915 18005 7967
rect 18019 7915 18071 7967
rect 18085 7915 18137 7967
rect 18151 7915 18203 7967
rect 18217 7915 18269 7967
rect 18282 7915 18334 7967
rect 18347 7915 18399 7967
rect 18412 7915 18464 7967
rect 18477 7915 18529 7967
rect 18542 7915 18594 7967
rect 18607 7915 18659 7967
rect 18672 7915 18724 7967
rect 18737 7915 18789 7967
rect 18802 7915 18854 7967
rect 18867 7915 18919 7967
rect 18932 7915 18984 7967
rect 18997 7915 19049 7967
rect 19062 7915 19114 7967
rect 19127 7915 19179 7967
rect 19192 7915 19244 7967
rect 19257 7915 19309 7967
rect 17029 7851 17081 7903
rect 17095 7851 17147 7903
rect 17161 7851 17213 7903
rect 17227 7851 17279 7903
rect 17293 7851 17345 7903
rect 17359 7851 17411 7903
rect 17425 7851 17477 7903
rect 17491 7851 17543 7903
rect 17557 7851 17609 7903
rect 17623 7851 17675 7903
rect 17689 7851 17741 7903
rect 17755 7851 17807 7903
rect 17821 7851 17873 7903
rect 17887 7851 17939 7903
rect 17953 7851 18005 7903
rect 18019 7851 18071 7903
rect 18085 7851 18137 7903
rect 18151 7851 18203 7903
rect 18217 7851 18269 7903
rect 18282 7851 18334 7903
rect 18347 7851 18399 7903
rect 18412 7851 18464 7903
rect 18477 7851 18529 7903
rect 18542 7851 18594 7903
rect 18607 7851 18659 7903
rect 18672 7851 18724 7903
rect 18737 7851 18789 7903
rect 18802 7851 18854 7903
rect 18867 7851 18919 7903
rect 18932 7851 18984 7903
rect 18997 7851 19049 7903
rect 19062 7851 19114 7903
rect 19127 7851 19179 7903
rect 19192 7851 19244 7903
rect 19257 7851 19309 7903
rect 17029 7787 17081 7839
rect 17095 7787 17147 7839
rect 17161 7787 17213 7839
rect 17227 7787 17279 7839
rect 17293 7787 17345 7839
rect 17359 7787 17411 7839
rect 17425 7787 17477 7839
rect 17491 7787 17543 7839
rect 17557 7787 17609 7839
rect 17623 7787 17675 7839
rect 17689 7787 17741 7839
rect 17755 7787 17807 7839
rect 17821 7787 17873 7839
rect 17887 7787 17939 7839
rect 17953 7787 18005 7839
rect 18019 7787 18071 7839
rect 18085 7787 18137 7839
rect 18151 7787 18203 7839
rect 18217 7787 18269 7839
rect 18282 7787 18334 7839
rect 18347 7787 18399 7839
rect 18412 7787 18464 7839
rect 18477 7787 18529 7839
rect 18542 7787 18594 7839
rect 18607 7787 18659 7839
rect 18672 7787 18724 7839
rect 18737 7787 18789 7839
rect 18802 7787 18854 7839
rect 18867 7787 18919 7839
rect 18932 7787 18984 7839
rect 18997 7787 19049 7839
rect 19062 7787 19114 7839
rect 19127 7787 19179 7839
rect 19192 7787 19244 7839
rect 19257 7787 19309 7839
rect 20702 7915 20754 7967
rect 20768 7915 20820 7967
rect 20834 7915 20886 7967
rect 20900 7915 20952 7967
rect 20966 7915 21018 7967
rect 21032 7915 21084 7967
rect 21097 7915 21149 7967
rect 21162 7915 21214 7967
rect 21227 7915 21279 7967
rect 21292 7915 21344 7967
rect 21357 7915 21409 7967
rect 20702 7851 20754 7903
rect 20768 7851 20820 7903
rect 20834 7851 20886 7903
rect 20900 7851 20952 7903
rect 20966 7851 21018 7903
rect 21032 7851 21084 7903
rect 21097 7851 21149 7903
rect 21162 7851 21214 7903
rect 21227 7851 21279 7903
rect 21292 7851 21344 7903
rect 21357 7851 21409 7903
rect 20702 7787 20754 7839
rect 20768 7787 20820 7839
rect 20834 7787 20886 7839
rect 20900 7787 20952 7839
rect 20966 7787 21018 7839
rect 21032 7787 21084 7839
rect 21097 7787 21149 7839
rect 21162 7787 21214 7839
rect 21227 7787 21279 7839
rect 21292 7787 21344 7839
rect 21357 7787 21409 7839
rect 17029 7651 17081 7703
rect 17095 7651 17147 7703
rect 17161 7651 17213 7703
rect 17227 7651 17279 7703
rect 17293 7651 17345 7703
rect 17359 7651 17411 7703
rect 17425 7651 17477 7703
rect 17491 7651 17543 7703
rect 17557 7651 17609 7703
rect 17623 7651 17675 7703
rect 17689 7651 17741 7703
rect 17755 7651 17807 7703
rect 17821 7651 17873 7703
rect 17887 7651 17939 7703
rect 17953 7651 18005 7703
rect 18019 7651 18071 7703
rect 18085 7651 18137 7703
rect 18151 7651 18203 7703
rect 18217 7651 18269 7703
rect 18282 7651 18334 7703
rect 18347 7651 18399 7703
rect 18412 7651 18464 7703
rect 18477 7651 18529 7703
rect 18542 7651 18594 7703
rect 18607 7651 18659 7703
rect 18672 7651 18724 7703
rect 18737 7651 18789 7703
rect 18802 7651 18854 7703
rect 18867 7651 18919 7703
rect 18932 7651 18984 7703
rect 18997 7651 19049 7703
rect 19062 7651 19114 7703
rect 19127 7651 19179 7703
rect 19192 7651 19244 7703
rect 19257 7651 19309 7703
rect 17029 7587 17081 7639
rect 17095 7587 17147 7639
rect 17161 7587 17213 7639
rect 17227 7587 17279 7639
rect 17293 7587 17345 7639
rect 17359 7587 17411 7639
rect 17425 7587 17477 7639
rect 17491 7587 17543 7639
rect 17557 7587 17609 7639
rect 17623 7587 17675 7639
rect 17689 7587 17741 7639
rect 17755 7587 17807 7639
rect 17821 7587 17873 7639
rect 17887 7587 17939 7639
rect 17953 7587 18005 7639
rect 18019 7587 18071 7639
rect 18085 7587 18137 7639
rect 18151 7587 18203 7639
rect 18217 7587 18269 7639
rect 18282 7587 18334 7639
rect 18347 7587 18399 7639
rect 18412 7587 18464 7639
rect 18477 7587 18529 7639
rect 18542 7587 18594 7639
rect 18607 7587 18659 7639
rect 18672 7587 18724 7639
rect 18737 7587 18789 7639
rect 18802 7587 18854 7639
rect 18867 7587 18919 7639
rect 18932 7587 18984 7639
rect 18997 7587 19049 7639
rect 19062 7587 19114 7639
rect 19127 7587 19179 7639
rect 19192 7587 19244 7639
rect 19257 7587 19309 7639
rect 17029 7523 17081 7575
rect 17095 7523 17147 7575
rect 17161 7523 17213 7575
rect 17227 7523 17279 7575
rect 17293 7523 17345 7575
rect 17359 7523 17411 7575
rect 17425 7523 17477 7575
rect 17491 7523 17543 7575
rect 17557 7523 17609 7575
rect 17623 7523 17675 7575
rect 17689 7523 17741 7575
rect 17755 7523 17807 7575
rect 17821 7523 17873 7575
rect 17887 7523 17939 7575
rect 17953 7523 18005 7575
rect 18019 7523 18071 7575
rect 18085 7523 18137 7575
rect 18151 7523 18203 7575
rect 18217 7523 18269 7575
rect 18282 7523 18334 7575
rect 18347 7523 18399 7575
rect 18412 7523 18464 7575
rect 18477 7523 18529 7575
rect 18542 7523 18594 7575
rect 18607 7523 18659 7575
rect 18672 7523 18724 7575
rect 18737 7523 18789 7575
rect 18802 7523 18854 7575
rect 18867 7523 18919 7575
rect 18932 7523 18984 7575
rect 18997 7523 19049 7575
rect 19062 7523 19114 7575
rect 19127 7523 19179 7575
rect 19192 7523 19244 7575
rect 19257 7523 19309 7575
rect 20702 7651 20754 7703
rect 20768 7651 20820 7703
rect 20834 7651 20886 7703
rect 20900 7651 20952 7703
rect 20966 7651 21018 7703
rect 21032 7651 21084 7703
rect 21097 7651 21149 7703
rect 21162 7651 21214 7703
rect 21227 7651 21279 7703
rect 21292 7651 21344 7703
rect 21357 7651 21409 7703
rect 20702 7587 20754 7639
rect 20768 7587 20820 7639
rect 20834 7587 20886 7639
rect 20900 7587 20952 7639
rect 20966 7587 21018 7639
rect 21032 7587 21084 7639
rect 21097 7587 21149 7639
rect 21162 7587 21214 7639
rect 21227 7587 21279 7639
rect 21292 7587 21344 7639
rect 21357 7587 21409 7639
rect 20702 7523 20754 7575
rect 20768 7523 20820 7575
rect 20834 7523 20886 7575
rect 20900 7523 20952 7575
rect 20966 7523 21018 7575
rect 21032 7523 21084 7575
rect 21097 7523 21149 7575
rect 21162 7523 21214 7575
rect 21227 7523 21279 7575
rect 21292 7523 21344 7575
rect 21357 7523 21409 7575
rect 17029 7387 17081 7439
rect 17095 7387 17147 7439
rect 17161 7387 17213 7439
rect 17227 7387 17279 7439
rect 17293 7387 17345 7439
rect 17359 7387 17411 7439
rect 17425 7387 17477 7439
rect 17491 7387 17543 7439
rect 17557 7387 17609 7439
rect 17623 7387 17675 7439
rect 17689 7387 17741 7439
rect 17755 7387 17807 7439
rect 17821 7387 17873 7439
rect 17887 7387 17939 7439
rect 17953 7387 18005 7439
rect 18019 7387 18071 7439
rect 18085 7387 18137 7439
rect 18151 7387 18203 7439
rect 18217 7387 18269 7439
rect 18282 7387 18334 7439
rect 18347 7387 18399 7439
rect 18412 7387 18464 7439
rect 18477 7387 18529 7439
rect 18542 7387 18594 7439
rect 18607 7387 18659 7439
rect 18672 7387 18724 7439
rect 18737 7387 18789 7439
rect 18802 7387 18854 7439
rect 18867 7387 18919 7439
rect 18932 7387 18984 7439
rect 18997 7387 19049 7439
rect 19062 7387 19114 7439
rect 19127 7387 19179 7439
rect 19192 7387 19244 7439
rect 19257 7387 19309 7439
rect 17029 7323 17081 7375
rect 17095 7323 17147 7375
rect 17161 7323 17213 7375
rect 17227 7323 17279 7375
rect 17293 7323 17345 7375
rect 17359 7323 17411 7375
rect 17425 7323 17477 7375
rect 17491 7323 17543 7375
rect 17557 7323 17609 7375
rect 17623 7323 17675 7375
rect 17689 7323 17741 7375
rect 17755 7323 17807 7375
rect 17821 7323 17873 7375
rect 17887 7323 17939 7375
rect 17953 7323 18005 7375
rect 18019 7323 18071 7375
rect 18085 7323 18137 7375
rect 18151 7323 18203 7375
rect 18217 7323 18269 7375
rect 18282 7323 18334 7375
rect 18347 7323 18399 7375
rect 18412 7323 18464 7375
rect 18477 7323 18529 7375
rect 18542 7323 18594 7375
rect 18607 7323 18659 7375
rect 18672 7323 18724 7375
rect 18737 7323 18789 7375
rect 18802 7323 18854 7375
rect 18867 7323 18919 7375
rect 18932 7323 18984 7375
rect 18997 7323 19049 7375
rect 19062 7323 19114 7375
rect 19127 7323 19179 7375
rect 19192 7323 19244 7375
rect 19257 7323 19309 7375
rect 17029 7259 17081 7311
rect 17095 7259 17147 7311
rect 17161 7259 17213 7311
rect 17227 7259 17279 7311
rect 17293 7259 17345 7311
rect 17359 7259 17411 7311
rect 17425 7259 17477 7311
rect 17491 7259 17543 7311
rect 17557 7259 17609 7311
rect 17623 7259 17675 7311
rect 17689 7259 17741 7311
rect 17755 7259 17807 7311
rect 17821 7259 17873 7311
rect 17887 7259 17939 7311
rect 17953 7259 18005 7311
rect 18019 7259 18071 7311
rect 18085 7259 18137 7311
rect 18151 7259 18203 7311
rect 18217 7259 18269 7311
rect 18282 7259 18334 7311
rect 18347 7259 18399 7311
rect 18412 7259 18464 7311
rect 18477 7259 18529 7311
rect 18542 7259 18594 7311
rect 18607 7259 18659 7311
rect 18672 7259 18724 7311
rect 18737 7259 18789 7311
rect 18802 7259 18854 7311
rect 18867 7259 18919 7311
rect 18932 7259 18984 7311
rect 18997 7259 19049 7311
rect 19062 7259 19114 7311
rect 19127 7259 19179 7311
rect 19192 7259 19244 7311
rect 19257 7259 19309 7311
rect 20702 7387 20754 7439
rect 20768 7387 20820 7439
rect 20834 7387 20886 7439
rect 20900 7387 20952 7439
rect 20966 7387 21018 7439
rect 21032 7387 21084 7439
rect 21097 7387 21149 7439
rect 21162 7387 21214 7439
rect 21227 7387 21279 7439
rect 21292 7387 21344 7439
rect 21357 7387 21409 7439
rect 20702 7323 20754 7375
rect 20768 7323 20820 7375
rect 20834 7323 20886 7375
rect 20900 7323 20952 7375
rect 20966 7323 21018 7375
rect 21032 7323 21084 7375
rect 21097 7323 21149 7375
rect 21162 7323 21214 7375
rect 21227 7323 21279 7375
rect 21292 7323 21344 7375
rect 21357 7323 21409 7375
rect 20702 7259 20754 7311
rect 20768 7259 20820 7311
rect 20834 7259 20886 7311
rect 20900 7259 20952 7311
rect 20966 7259 21018 7311
rect 21032 7259 21084 7311
rect 21097 7259 21149 7311
rect 21162 7259 21214 7311
rect 21227 7259 21279 7311
rect 21292 7259 21344 7311
rect 21357 7259 21409 7311
rect 17029 7123 17081 7175
rect 17095 7123 17147 7175
rect 17161 7123 17213 7175
rect 17227 7123 17279 7175
rect 17293 7123 17345 7175
rect 17359 7123 17411 7175
rect 17425 7123 17477 7175
rect 17491 7123 17543 7175
rect 17557 7123 17609 7175
rect 17623 7123 17675 7175
rect 17689 7123 17741 7175
rect 17755 7123 17807 7175
rect 17821 7123 17873 7175
rect 17887 7123 17939 7175
rect 17953 7123 18005 7175
rect 18019 7123 18071 7175
rect 18085 7123 18137 7175
rect 18151 7123 18203 7175
rect 18217 7123 18269 7175
rect 18282 7123 18334 7175
rect 18347 7123 18399 7175
rect 18412 7123 18464 7175
rect 18477 7123 18529 7175
rect 18542 7123 18594 7175
rect 18607 7123 18659 7175
rect 18672 7123 18724 7175
rect 18737 7123 18789 7175
rect 18802 7123 18854 7175
rect 18867 7123 18919 7175
rect 18932 7123 18984 7175
rect 18997 7123 19049 7175
rect 19062 7123 19114 7175
rect 19127 7123 19179 7175
rect 19192 7123 19244 7175
rect 19257 7123 19309 7175
rect 17029 7059 17081 7111
rect 17095 7059 17147 7111
rect 17161 7059 17213 7111
rect 17227 7059 17279 7111
rect 17293 7059 17345 7111
rect 17359 7059 17411 7111
rect 17425 7059 17477 7111
rect 17491 7059 17543 7111
rect 17557 7059 17609 7111
rect 17623 7059 17675 7111
rect 17689 7059 17741 7111
rect 17755 7059 17807 7111
rect 17821 7059 17873 7111
rect 17887 7059 17939 7111
rect 17953 7059 18005 7111
rect 18019 7059 18071 7111
rect 18085 7059 18137 7111
rect 18151 7059 18203 7111
rect 18217 7059 18269 7111
rect 18282 7059 18334 7111
rect 18347 7059 18399 7111
rect 18412 7059 18464 7111
rect 18477 7059 18529 7111
rect 18542 7059 18594 7111
rect 18607 7059 18659 7111
rect 18672 7059 18724 7111
rect 18737 7059 18789 7111
rect 18802 7059 18854 7111
rect 18867 7059 18919 7111
rect 18932 7059 18984 7111
rect 18997 7059 19049 7111
rect 19062 7059 19114 7111
rect 19127 7059 19179 7111
rect 19192 7059 19244 7111
rect 19257 7059 19309 7111
rect 17029 6995 17081 7047
rect 17095 6995 17147 7047
rect 17161 6995 17213 7047
rect 17227 6995 17279 7047
rect 17293 6995 17345 7047
rect 17359 6995 17411 7047
rect 17425 6995 17477 7047
rect 17491 6995 17543 7047
rect 17557 6995 17609 7047
rect 17623 6995 17675 7047
rect 17689 6995 17741 7047
rect 17755 6995 17807 7047
rect 17821 6995 17873 7047
rect 17887 6995 17939 7047
rect 17953 6995 18005 7047
rect 18019 6995 18071 7047
rect 18085 6995 18137 7047
rect 18151 6995 18203 7047
rect 18217 6995 18269 7047
rect 18282 6995 18334 7047
rect 18347 6995 18399 7047
rect 18412 6995 18464 7047
rect 18477 6995 18529 7047
rect 18542 6995 18594 7047
rect 18607 6995 18659 7047
rect 18672 6995 18724 7047
rect 18737 6995 18789 7047
rect 18802 6995 18854 7047
rect 18867 6995 18919 7047
rect 18932 6995 18984 7047
rect 18997 6995 19049 7047
rect 19062 6995 19114 7047
rect 19127 6995 19179 7047
rect 19192 6995 19244 7047
rect 19257 6995 19309 7047
rect 20702 7123 20754 7175
rect 20768 7123 20820 7175
rect 20834 7123 20886 7175
rect 20900 7123 20952 7175
rect 20966 7123 21018 7175
rect 21032 7123 21084 7175
rect 21097 7123 21149 7175
rect 21162 7123 21214 7175
rect 21227 7123 21279 7175
rect 21292 7123 21344 7175
rect 21357 7123 21409 7175
rect 20702 7059 20754 7111
rect 20768 7059 20820 7111
rect 20834 7059 20886 7111
rect 20900 7059 20952 7111
rect 20966 7059 21018 7111
rect 21032 7059 21084 7111
rect 21097 7059 21149 7111
rect 21162 7059 21214 7111
rect 21227 7059 21279 7111
rect 21292 7059 21344 7111
rect 21357 7059 21409 7111
rect 20702 6995 20754 7047
rect 20768 6995 20820 7047
rect 20834 6995 20886 7047
rect 20900 6995 20952 7047
rect 20966 6995 21018 7047
rect 21032 6995 21084 7047
rect 21097 6995 21149 7047
rect 21162 6995 21214 7047
rect 21227 6995 21279 7047
rect 21292 6995 21344 7047
rect 21357 6995 21409 7047
rect 23941 8680 24505 9126
rect 23941 7854 24505 8680
rect 23941 7815 24505 7854
rect 23941 7781 23959 7815
rect 23959 7781 23997 7815
rect 23997 7781 24031 7815
rect 24031 7781 24069 7815
rect 24069 7781 24103 7815
rect 24103 7781 24141 7815
rect 24141 7781 24175 7815
rect 24175 7781 24213 7815
rect 24213 7781 24247 7815
rect 24247 7781 24285 7815
rect 24285 7781 24319 7815
rect 24319 7781 24357 7815
rect 24357 7781 24391 7815
rect 24391 7781 24429 7815
rect 24429 7781 24463 7815
rect 24463 7781 24501 7815
rect 24501 7781 24505 7815
rect 23941 7742 24505 7781
rect 23941 7708 23959 7742
rect 23959 7708 23997 7742
rect 23997 7708 24031 7742
rect 24031 7708 24069 7742
rect 24069 7708 24103 7742
rect 24103 7708 24141 7742
rect 24141 7708 24175 7742
rect 24175 7708 24213 7742
rect 24213 7708 24247 7742
rect 24247 7708 24285 7742
rect 24285 7708 24319 7742
rect 24319 7708 24357 7742
rect 24357 7708 24391 7742
rect 24391 7708 24429 7742
rect 24429 7708 24463 7742
rect 24463 7708 24501 7742
rect 24501 7708 24505 7742
rect 23941 7669 24505 7708
rect 23941 7635 23959 7669
rect 23959 7635 23997 7669
rect 23997 7635 24031 7669
rect 24031 7635 24069 7669
rect 24069 7635 24103 7669
rect 24103 7635 24141 7669
rect 24141 7635 24175 7669
rect 24175 7635 24213 7669
rect 24213 7635 24247 7669
rect 24247 7635 24285 7669
rect 24285 7635 24319 7669
rect 24319 7635 24357 7669
rect 24357 7635 24391 7669
rect 24391 7635 24429 7669
rect 24429 7635 24463 7669
rect 24463 7635 24501 7669
rect 24501 7635 24505 7669
rect 23941 7596 24505 7635
rect 23941 7562 23959 7596
rect 23959 7562 23997 7596
rect 23997 7562 24031 7596
rect 24031 7562 24069 7596
rect 24069 7562 24103 7596
rect 24103 7562 24141 7596
rect 24141 7562 24175 7596
rect 24175 7562 24213 7596
rect 24213 7562 24247 7596
rect 24247 7562 24285 7596
rect 24285 7562 24319 7596
rect 24319 7562 24357 7596
rect 24357 7562 24391 7596
rect 24391 7562 24429 7596
rect 24429 7562 24463 7596
rect 24463 7562 24501 7596
rect 24501 7562 24505 7596
rect 23941 7523 24505 7562
rect 23941 7489 23959 7523
rect 23959 7489 23997 7523
rect 23997 7489 24031 7523
rect 24031 7489 24069 7523
rect 24069 7489 24103 7523
rect 24103 7489 24141 7523
rect 24141 7489 24175 7523
rect 24175 7489 24213 7523
rect 24213 7489 24247 7523
rect 24247 7489 24285 7523
rect 24285 7489 24319 7523
rect 24319 7489 24357 7523
rect 24357 7489 24391 7523
rect 24391 7489 24429 7523
rect 24429 7489 24463 7523
rect 24463 7489 24501 7523
rect 24501 7489 24505 7523
rect 23941 7450 24505 7489
rect 23941 7416 23959 7450
rect 23959 7416 23997 7450
rect 23997 7416 24031 7450
rect 24031 7416 24069 7450
rect 24069 7416 24103 7450
rect 24103 7416 24141 7450
rect 24141 7416 24175 7450
rect 24175 7416 24213 7450
rect 24213 7416 24247 7450
rect 24247 7416 24285 7450
rect 24285 7416 24319 7450
rect 24319 7416 24357 7450
rect 24357 7416 24391 7450
rect 24391 7416 24429 7450
rect 24429 7416 24463 7450
rect 24463 7416 24501 7450
rect 24501 7416 24505 7450
rect 23941 7377 24505 7416
rect 23941 7343 23959 7377
rect 23959 7343 23997 7377
rect 23997 7343 24031 7377
rect 24031 7343 24069 7377
rect 24069 7343 24103 7377
rect 24103 7343 24141 7377
rect 24141 7343 24175 7377
rect 24175 7343 24213 7377
rect 24213 7343 24247 7377
rect 24247 7343 24285 7377
rect 24285 7343 24319 7377
rect 24319 7343 24357 7377
rect 24357 7343 24391 7377
rect 24391 7343 24429 7377
rect 24429 7343 24463 7377
rect 24463 7343 24501 7377
rect 24501 7343 24505 7377
rect 23941 7304 24505 7343
rect 23941 7270 23959 7304
rect 23959 7270 23997 7304
rect 23997 7270 24031 7304
rect 24031 7270 24069 7304
rect 24069 7270 24103 7304
rect 24103 7270 24141 7304
rect 24141 7270 24175 7304
rect 24175 7270 24213 7304
rect 24213 7270 24247 7304
rect 24247 7270 24285 7304
rect 24285 7270 24319 7304
rect 24319 7270 24357 7304
rect 24357 7270 24391 7304
rect 24391 7270 24429 7304
rect 24429 7270 24463 7304
rect 24463 7270 24501 7304
rect 24501 7270 24505 7304
rect 23941 7231 24505 7270
rect 23941 7218 23959 7231
rect 23959 7218 23997 7231
rect 23997 7218 24031 7231
rect 24031 7218 24069 7231
rect 24069 7218 24103 7231
rect 24103 7218 24141 7231
rect 24141 7218 24175 7231
rect 24175 7218 24213 7231
rect 24213 7218 24247 7231
rect 24247 7218 24285 7231
rect 24285 7218 24319 7231
rect 24319 7218 24357 7231
rect 24357 7218 24391 7231
rect 24391 7218 24429 7231
rect 24429 7218 24463 7231
rect 24463 7218 24501 7231
rect 24501 7218 24505 7231
rect 23941 7197 23959 7205
rect 23959 7197 23993 7205
rect 24005 7197 24031 7205
rect 24031 7197 24057 7205
rect 23941 7158 23993 7197
rect 24005 7158 24057 7197
rect 23941 7153 23959 7158
rect 23959 7153 23993 7158
rect 24005 7153 24031 7158
rect 24031 7153 24057 7158
rect 24069 7197 24103 7205
rect 24103 7197 24121 7205
rect 24069 7158 24121 7197
rect 24069 7153 24103 7158
rect 24103 7153 24121 7158
rect 24133 7197 24141 7205
rect 24141 7197 24175 7205
rect 24175 7197 24185 7205
rect 24133 7158 24185 7197
rect 24133 7153 24141 7158
rect 24141 7153 24175 7158
rect 24175 7153 24185 7158
rect 24197 7197 24213 7205
rect 24213 7197 24247 7205
rect 24247 7197 24249 7205
rect 24197 7158 24249 7197
rect 24197 7153 24213 7158
rect 24213 7153 24247 7158
rect 24247 7153 24249 7158
rect 24261 7197 24285 7205
rect 24285 7197 24313 7205
rect 24325 7197 24357 7205
rect 24357 7197 24377 7205
rect 24389 7197 24391 7205
rect 24391 7197 24429 7205
rect 24429 7197 24441 7205
rect 24453 7197 24463 7205
rect 24463 7197 24501 7205
rect 24501 7197 24505 7205
rect 24261 7158 24313 7197
rect 24325 7158 24377 7197
rect 24389 7158 24441 7197
rect 24453 7158 24505 7197
rect 24261 7153 24285 7158
rect 24285 7153 24313 7158
rect 24325 7153 24357 7158
rect 24357 7153 24377 7158
rect 24389 7153 24391 7158
rect 24391 7153 24429 7158
rect 24429 7153 24441 7158
rect 24453 7153 24463 7158
rect 24463 7153 24501 7158
rect 24501 7153 24505 7158
rect 23941 7124 23959 7140
rect 23959 7124 23993 7140
rect 24005 7124 24031 7140
rect 24031 7124 24057 7140
rect 23941 7088 23993 7124
rect 24005 7088 24057 7124
rect 24069 7124 24103 7140
rect 24103 7124 24121 7140
rect 24069 7088 24121 7124
rect 24133 7124 24141 7140
rect 24141 7124 24175 7140
rect 24175 7124 24185 7140
rect 24133 7088 24185 7124
rect 24197 7124 24213 7140
rect 24213 7124 24247 7140
rect 24247 7124 24249 7140
rect 24197 7088 24249 7124
rect 24261 7124 24285 7140
rect 24285 7124 24313 7140
rect 24325 7124 24357 7140
rect 24357 7124 24377 7140
rect 24389 7124 24391 7140
rect 24391 7124 24429 7140
rect 24429 7124 24441 7140
rect 24453 7124 24463 7140
rect 24463 7124 24501 7140
rect 24501 7124 24505 7140
rect 24261 7088 24313 7124
rect 24325 7088 24377 7124
rect 24389 7088 24441 7124
rect 24453 7088 24505 7124
rect 23941 7051 23959 7075
rect 23959 7051 23993 7075
rect 24005 7051 24031 7075
rect 24031 7051 24057 7075
rect 23941 7023 23993 7051
rect 24005 7023 24057 7051
rect 24069 7051 24103 7075
rect 24103 7051 24121 7075
rect 24069 7023 24121 7051
rect 24133 7051 24141 7075
rect 24141 7051 24175 7075
rect 24175 7051 24185 7075
rect 24133 7023 24185 7051
rect 24197 7051 24213 7075
rect 24213 7051 24247 7075
rect 24247 7051 24249 7075
rect 24197 7023 24249 7051
rect 24261 7051 24285 7075
rect 24285 7051 24313 7075
rect 24325 7051 24357 7075
rect 24357 7051 24377 7075
rect 24389 7051 24391 7075
rect 24391 7051 24429 7075
rect 24429 7051 24441 7075
rect 24453 7051 24463 7075
rect 24463 7051 24501 7075
rect 24501 7051 24505 7075
rect 24261 7023 24313 7051
rect 24325 7023 24377 7051
rect 24389 7023 24441 7051
rect 24453 7023 24505 7051
rect 23941 6978 23959 7010
rect 23959 6978 23993 7010
rect 24005 6978 24031 7010
rect 24031 6978 24057 7010
rect 23941 6958 23993 6978
rect 24005 6958 24057 6978
rect 24069 6978 24103 7010
rect 24103 6978 24121 7010
rect 24069 6958 24121 6978
rect 24133 6978 24141 7010
rect 24141 6978 24175 7010
rect 24175 6978 24185 7010
rect 24133 6958 24185 6978
rect 24197 6978 24213 7010
rect 24213 6978 24247 7010
rect 24247 6978 24249 7010
rect 24197 6958 24249 6978
rect 24261 6978 24285 7010
rect 24285 6978 24313 7010
rect 24325 6978 24357 7010
rect 24357 6978 24377 7010
rect 24389 6978 24391 7010
rect 24391 6978 24429 7010
rect 24429 6978 24441 7010
rect 24453 6978 24463 7010
rect 24463 6978 24501 7010
rect 24501 6978 24505 7010
rect 24261 6958 24313 6978
rect 24325 6958 24377 6978
rect 24389 6958 24441 6978
rect 24453 6958 24505 6978
rect 25528 6948 25580 7000
rect 25592 6948 25644 7000
rect 28183 6948 28235 7000
rect 28271 6948 28323 7000
rect 23941 6939 23993 6945
rect 24005 6939 24057 6945
rect 23941 6905 23959 6939
rect 23959 6905 23993 6939
rect 24005 6905 24031 6939
rect 24031 6905 24057 6939
rect 23941 6893 23993 6905
rect 24005 6893 24057 6905
rect 24069 6939 24121 6945
rect 24069 6905 24103 6939
rect 24103 6905 24121 6939
rect 24069 6893 24121 6905
rect 24133 6939 24185 6945
rect 24133 6905 24141 6939
rect 24141 6905 24175 6939
rect 24175 6905 24185 6939
rect 24133 6893 24185 6905
rect 24197 6939 24249 6945
rect 24197 6905 24213 6939
rect 24213 6905 24247 6939
rect 24247 6905 24249 6939
rect 24197 6893 24249 6905
rect 24261 6939 24313 6945
rect 24325 6939 24377 6945
rect 24389 6939 24441 6945
rect 24453 6939 24505 6945
rect 24261 6905 24285 6939
rect 24285 6905 24313 6939
rect 24325 6905 24357 6939
rect 24357 6905 24377 6939
rect 24389 6905 24391 6939
rect 24391 6905 24429 6939
rect 24429 6905 24441 6939
rect 24453 6905 24463 6939
rect 24463 6905 24501 6939
rect 24501 6905 24505 6939
rect 24261 6893 24313 6905
rect 24325 6893 24377 6905
rect 24389 6893 24441 6905
rect 24453 6893 24505 6905
rect 23941 6866 23993 6880
rect 24005 6866 24057 6880
rect 23941 6832 23959 6866
rect 23959 6832 23993 6866
rect 24005 6832 24031 6866
rect 24031 6832 24057 6866
rect 23941 6828 23993 6832
rect 24005 6828 24057 6832
rect 24069 6866 24121 6880
rect 24069 6832 24103 6866
rect 24103 6832 24121 6866
rect 24069 6828 24121 6832
rect 24133 6866 24185 6880
rect 24133 6832 24141 6866
rect 24141 6832 24175 6866
rect 24175 6832 24185 6866
rect 24133 6828 24185 6832
rect 24197 6866 24249 6880
rect 24197 6832 24213 6866
rect 24213 6832 24247 6866
rect 24247 6832 24249 6866
rect 24197 6828 24249 6832
rect 24261 6866 24313 6880
rect 24325 6866 24377 6880
rect 24389 6866 24441 6880
rect 24453 6866 24505 6880
rect 24261 6832 24285 6866
rect 24285 6832 24313 6866
rect 24325 6832 24357 6866
rect 24357 6832 24377 6866
rect 24389 6832 24391 6866
rect 24391 6832 24429 6866
rect 24429 6832 24441 6866
rect 24453 6832 24463 6866
rect 24463 6832 24501 6866
rect 24501 6832 24505 6866
rect 24261 6828 24313 6832
rect 24325 6828 24377 6832
rect 24389 6828 24441 6832
rect 24453 6828 24505 6832
rect 23941 6793 23993 6815
rect 24005 6793 24057 6815
rect 23941 6763 23959 6793
rect 23959 6763 23993 6793
rect 24005 6763 24031 6793
rect 24031 6763 24057 6793
rect 24069 6793 24121 6815
rect 24069 6763 24103 6793
rect 24103 6763 24121 6793
rect 24133 6793 24185 6815
rect 24133 6763 24141 6793
rect 24141 6763 24175 6793
rect 24175 6763 24185 6793
rect 24197 6793 24249 6815
rect 24197 6763 24213 6793
rect 24213 6763 24247 6793
rect 24247 6763 24249 6793
rect 24261 6793 24313 6815
rect 24325 6793 24377 6815
rect 24389 6793 24441 6815
rect 24453 6793 24505 6815
rect 24261 6763 24285 6793
rect 24285 6763 24313 6793
rect 24325 6763 24357 6793
rect 24357 6763 24377 6793
rect 24389 6763 24391 6793
rect 24391 6763 24429 6793
rect 24429 6763 24441 6793
rect 24453 6763 24463 6793
rect 24463 6763 24501 6793
rect 24501 6763 24505 6793
rect 23941 6720 23993 6750
rect 24005 6720 24057 6750
rect 23941 6698 23959 6720
rect 23959 6698 23993 6720
rect 24005 6698 24031 6720
rect 24031 6698 24057 6720
rect 24069 6720 24121 6750
rect 24069 6698 24103 6720
rect 24103 6698 24121 6720
rect 24133 6720 24185 6750
rect 24133 6698 24141 6720
rect 24141 6698 24175 6720
rect 24175 6698 24185 6720
rect 24197 6720 24249 6750
rect 24197 6698 24213 6720
rect 24213 6698 24247 6720
rect 24247 6698 24249 6720
rect 24261 6720 24313 6750
rect 24325 6720 24377 6750
rect 24389 6720 24441 6750
rect 24453 6720 24505 6750
rect 24261 6698 24285 6720
rect 24285 6698 24313 6720
rect 24325 6698 24357 6720
rect 24357 6698 24377 6720
rect 24389 6698 24391 6720
rect 24391 6698 24429 6720
rect 24429 6698 24441 6720
rect 24453 6698 24463 6720
rect 24463 6698 24501 6720
rect 24501 6698 24505 6720
rect 23941 6647 23993 6685
rect 24005 6647 24057 6685
rect 23941 6633 23959 6647
rect 23959 6633 23993 6647
rect 24005 6633 24031 6647
rect 24031 6633 24057 6647
rect 24069 6647 24121 6685
rect 24069 6633 24103 6647
rect 24103 6633 24121 6647
rect 24133 6647 24185 6685
rect 24133 6633 24141 6647
rect 24141 6633 24175 6647
rect 24175 6633 24185 6647
rect 24197 6647 24249 6685
rect 24197 6633 24213 6647
rect 24213 6633 24247 6647
rect 24247 6633 24249 6647
rect 24261 6647 24313 6685
rect 24325 6647 24377 6685
rect 24389 6647 24441 6685
rect 24453 6647 24505 6685
rect 24261 6633 24285 6647
rect 24285 6633 24313 6647
rect 24325 6633 24357 6647
rect 24357 6633 24377 6647
rect 24389 6633 24391 6647
rect 24391 6633 24429 6647
rect 24429 6633 24441 6647
rect 24453 6633 24463 6647
rect 24463 6633 24501 6647
rect 24501 6633 24505 6647
rect 23941 6613 23959 6620
rect 23959 6613 23993 6620
rect 24005 6613 24031 6620
rect 24031 6613 24057 6620
rect 23941 6574 23993 6613
rect 24005 6574 24057 6613
rect 23941 6568 23959 6574
rect 23959 6568 23993 6574
rect 24005 6568 24031 6574
rect 24031 6568 24057 6574
rect 24069 6613 24103 6620
rect 24103 6613 24121 6620
rect 24069 6574 24121 6613
rect 24069 6568 24103 6574
rect 24103 6568 24121 6574
rect 24133 6613 24141 6620
rect 24141 6613 24175 6620
rect 24175 6613 24185 6620
rect 24133 6574 24185 6613
rect 24133 6568 24141 6574
rect 24141 6568 24175 6574
rect 24175 6568 24185 6574
rect 24197 6613 24213 6620
rect 24213 6613 24247 6620
rect 24247 6613 24249 6620
rect 24197 6574 24249 6613
rect 24197 6568 24213 6574
rect 24213 6568 24247 6574
rect 24247 6568 24249 6574
rect 24261 6613 24285 6620
rect 24285 6613 24313 6620
rect 24325 6613 24357 6620
rect 24357 6613 24377 6620
rect 24389 6613 24391 6620
rect 24391 6613 24429 6620
rect 24429 6613 24441 6620
rect 24453 6613 24463 6620
rect 24463 6613 24501 6620
rect 24501 6613 24505 6620
rect 24261 6574 24313 6613
rect 24325 6574 24377 6613
rect 24389 6574 24441 6613
rect 24453 6574 24505 6613
rect 24261 6568 24285 6574
rect 24285 6568 24313 6574
rect 24325 6568 24357 6574
rect 24357 6568 24377 6574
rect 24389 6568 24391 6574
rect 24391 6568 24429 6574
rect 24429 6568 24441 6574
rect 24453 6568 24463 6574
rect 24463 6568 24501 6574
rect 24501 6568 24505 6574
rect 23941 6540 23959 6555
rect 23959 6540 23993 6555
rect 24005 6540 24031 6555
rect 24031 6540 24057 6555
rect 23941 6503 23993 6540
rect 24005 6503 24057 6540
rect 24069 6540 24103 6555
rect 24103 6540 24121 6555
rect 24069 6503 24121 6540
rect 24133 6540 24141 6555
rect 24141 6540 24175 6555
rect 24175 6540 24185 6555
rect 24133 6503 24185 6540
rect 24197 6540 24213 6555
rect 24213 6540 24247 6555
rect 24247 6540 24249 6555
rect 24197 6503 24249 6540
rect 24261 6540 24285 6555
rect 24285 6540 24313 6555
rect 24325 6540 24357 6555
rect 24357 6540 24377 6555
rect 24389 6540 24391 6555
rect 24391 6540 24429 6555
rect 24429 6540 24441 6555
rect 24453 6540 24463 6555
rect 24463 6540 24501 6555
rect 24501 6540 24505 6555
rect 24261 6503 24313 6540
rect 24325 6503 24377 6540
rect 24389 6503 24441 6540
rect 24453 6503 24505 6540
rect 23941 6467 23959 6490
rect 23959 6467 23993 6490
rect 24005 6467 24031 6490
rect 24031 6467 24057 6490
rect 23941 6438 23993 6467
rect 24005 6438 24057 6467
rect 24069 6467 24103 6490
rect 24103 6467 24121 6490
rect 24069 6438 24121 6467
rect 24133 6467 24141 6490
rect 24141 6467 24175 6490
rect 24175 6467 24185 6490
rect 24133 6438 24185 6467
rect 24197 6467 24213 6490
rect 24213 6467 24247 6490
rect 24247 6467 24249 6490
rect 24197 6438 24249 6467
rect 24261 6467 24285 6490
rect 24285 6467 24313 6490
rect 24325 6467 24357 6490
rect 24357 6467 24377 6490
rect 24389 6467 24391 6490
rect 24391 6467 24429 6490
rect 24429 6467 24441 6490
rect 24453 6467 24463 6490
rect 24463 6467 24501 6490
rect 24501 6467 24505 6490
rect 24261 6438 24313 6467
rect 24325 6438 24377 6467
rect 24389 6438 24441 6467
rect 24453 6438 24505 6467
rect 23941 6394 23959 6425
rect 23959 6394 23993 6425
rect 24005 6394 24031 6425
rect 24031 6394 24057 6425
rect 23941 6373 23993 6394
rect 24005 6373 24057 6394
rect 24069 6394 24103 6425
rect 24103 6394 24121 6425
rect 24069 6373 24121 6394
rect 24133 6394 24141 6425
rect 24141 6394 24175 6425
rect 24175 6394 24185 6425
rect 24133 6373 24185 6394
rect 24197 6394 24213 6425
rect 24213 6394 24247 6425
rect 24247 6394 24249 6425
rect 24197 6373 24249 6394
rect 24261 6394 24285 6425
rect 24285 6394 24313 6425
rect 24325 6394 24357 6425
rect 24357 6394 24377 6425
rect 24389 6394 24391 6425
rect 24391 6394 24429 6425
rect 24429 6394 24441 6425
rect 24453 6394 24463 6425
rect 24463 6394 24501 6425
rect 24501 6394 24505 6425
rect 24261 6373 24313 6394
rect 24325 6373 24377 6394
rect 24389 6373 24441 6394
rect 24453 6373 24505 6394
rect 23941 6355 23993 6360
rect 24005 6355 24057 6360
rect 23941 6321 23959 6355
rect 23959 6321 23993 6355
rect 24005 6321 24031 6355
rect 24031 6321 24057 6355
rect 23941 6308 23993 6321
rect 24005 6308 24057 6321
rect 24069 6355 24121 6360
rect 24069 6321 24103 6355
rect 24103 6321 24121 6355
rect 24069 6308 24121 6321
rect 24133 6355 24185 6360
rect 24133 6321 24141 6355
rect 24141 6321 24175 6355
rect 24175 6321 24185 6355
rect 24133 6308 24185 6321
rect 24197 6355 24249 6360
rect 24197 6321 24213 6355
rect 24213 6321 24247 6355
rect 24247 6321 24249 6355
rect 24197 6308 24249 6321
rect 24261 6355 24313 6360
rect 24325 6355 24377 6360
rect 24389 6355 24441 6360
rect 24453 6355 24505 6360
rect 24261 6321 24285 6355
rect 24285 6321 24313 6355
rect 24325 6321 24357 6355
rect 24357 6321 24377 6355
rect 24389 6321 24391 6355
rect 24391 6321 24429 6355
rect 24429 6321 24441 6355
rect 24453 6321 24463 6355
rect 24463 6321 24501 6355
rect 24501 6321 24505 6355
rect 24261 6308 24313 6321
rect 24325 6308 24377 6321
rect 24389 6308 24441 6321
rect 24453 6308 24505 6321
rect 23941 6282 23993 6295
rect 24005 6282 24057 6295
rect 23941 6248 23959 6282
rect 23959 6248 23993 6282
rect 24005 6248 24031 6282
rect 24031 6248 24057 6282
rect 23941 6243 23993 6248
rect 24005 6243 24057 6248
rect 24069 6282 24121 6295
rect 24069 6248 24103 6282
rect 24103 6248 24121 6282
rect 24069 6243 24121 6248
rect 24133 6282 24185 6295
rect 24133 6248 24141 6282
rect 24141 6248 24175 6282
rect 24175 6248 24185 6282
rect 24133 6243 24185 6248
rect 24197 6282 24249 6295
rect 24197 6248 24213 6282
rect 24213 6248 24247 6282
rect 24247 6248 24249 6282
rect 24197 6243 24249 6248
rect 24261 6282 24313 6295
rect 24325 6282 24377 6295
rect 24389 6282 24441 6295
rect 24453 6282 24505 6295
rect 24261 6248 24285 6282
rect 24285 6248 24313 6282
rect 24325 6248 24357 6282
rect 24357 6248 24377 6282
rect 24389 6248 24391 6282
rect 24391 6248 24429 6282
rect 24429 6248 24441 6282
rect 24453 6248 24463 6282
rect 24463 6248 24501 6282
rect 24501 6248 24505 6282
rect 24261 6243 24313 6248
rect 24325 6243 24377 6248
rect 24389 6243 24441 6248
rect 24453 6243 24505 6248
rect 23941 6209 23993 6230
rect 24005 6209 24057 6230
rect 23941 6178 23959 6209
rect 23959 6178 23993 6209
rect 24005 6178 24031 6209
rect 24031 6178 24057 6209
rect 24069 6209 24121 6230
rect 24069 6178 24103 6209
rect 24103 6178 24121 6209
rect 24133 6209 24185 6230
rect 24133 6178 24141 6209
rect 24141 6178 24175 6209
rect 24175 6178 24185 6209
rect 24197 6209 24249 6230
rect 24197 6178 24213 6209
rect 24213 6178 24247 6209
rect 24247 6178 24249 6209
rect 24261 6209 24313 6230
rect 24325 6209 24377 6230
rect 24389 6209 24441 6230
rect 24453 6209 24505 6230
rect 24261 6178 24285 6209
rect 24285 6178 24313 6209
rect 24325 6178 24357 6209
rect 24357 6178 24377 6209
rect 24389 6178 24391 6209
rect 24391 6178 24429 6209
rect 24429 6178 24441 6209
rect 24453 6178 24463 6209
rect 24463 6178 24501 6209
rect 24501 6178 24505 6209
rect 23941 6136 23993 6165
rect 24005 6136 24057 6165
rect 23941 6113 23959 6136
rect 23959 6113 23993 6136
rect 24005 6113 24031 6136
rect 24031 6113 24057 6136
rect 24069 6136 24121 6165
rect 24069 6113 24103 6136
rect 24103 6113 24121 6136
rect 24133 6136 24185 6165
rect 24133 6113 24141 6136
rect 24141 6113 24175 6136
rect 24175 6113 24185 6136
rect 24197 6136 24249 6165
rect 24197 6113 24213 6136
rect 24213 6113 24247 6136
rect 24247 6113 24249 6136
rect 24261 6136 24313 6165
rect 24325 6136 24377 6165
rect 24389 6136 24441 6165
rect 24453 6136 24505 6165
rect 24261 6113 24285 6136
rect 24285 6113 24313 6136
rect 24325 6113 24357 6136
rect 24357 6113 24377 6136
rect 24389 6113 24391 6136
rect 24391 6113 24429 6136
rect 24429 6113 24441 6136
rect 24453 6113 24463 6136
rect 24463 6113 24501 6136
rect 24501 6113 24505 6136
rect 23941 6063 23993 6100
rect 24005 6063 24057 6100
rect 23941 6048 23959 6063
rect 23959 6048 23993 6063
rect 24005 6048 24031 6063
rect 24031 6048 24057 6063
rect 24069 6063 24121 6100
rect 24069 6048 24103 6063
rect 24103 6048 24121 6063
rect 24133 6063 24185 6100
rect 24133 6048 24141 6063
rect 24141 6048 24175 6063
rect 24175 6048 24185 6063
rect 24197 6063 24249 6100
rect 24197 6048 24213 6063
rect 24213 6048 24247 6063
rect 24247 6048 24249 6063
rect 24261 6063 24313 6100
rect 24325 6063 24377 6100
rect 24389 6063 24441 6100
rect 24453 6063 24505 6100
rect 24261 6048 24285 6063
rect 24285 6048 24313 6063
rect 24325 6048 24357 6063
rect 24357 6048 24377 6063
rect 24389 6048 24391 6063
rect 24391 6048 24429 6063
rect 24429 6048 24441 6063
rect 24453 6048 24463 6063
rect 24463 6048 24501 6063
rect 24501 6048 24505 6063
rect 23941 6029 23959 6035
rect 23959 6029 23993 6035
rect 24005 6029 24031 6035
rect 24031 6029 24057 6035
rect 23941 5990 23993 6029
rect 24005 5990 24057 6029
rect 23941 5983 23959 5990
rect 23959 5983 23993 5990
rect 24005 5983 24031 5990
rect 24031 5983 24057 5990
rect 24069 6029 24103 6035
rect 24103 6029 24121 6035
rect 24069 5990 24121 6029
rect 24069 5983 24103 5990
rect 24103 5983 24121 5990
rect 24133 6029 24141 6035
rect 24141 6029 24175 6035
rect 24175 6029 24185 6035
rect 24133 5990 24185 6029
rect 24133 5983 24141 5990
rect 24141 5983 24175 5990
rect 24175 5983 24185 5990
rect 24197 6029 24213 6035
rect 24213 6029 24247 6035
rect 24247 6029 24249 6035
rect 24197 5990 24249 6029
rect 24197 5983 24213 5990
rect 24213 5983 24247 5990
rect 24247 5983 24249 5990
rect 24261 6029 24285 6035
rect 24285 6029 24313 6035
rect 24325 6029 24357 6035
rect 24357 6029 24377 6035
rect 24389 6029 24391 6035
rect 24391 6029 24429 6035
rect 24429 6029 24441 6035
rect 24453 6029 24463 6035
rect 24463 6029 24501 6035
rect 24501 6029 24505 6035
rect 24261 5990 24313 6029
rect 24325 5990 24377 6029
rect 24389 5990 24441 6029
rect 24453 5990 24505 6029
rect 24261 5983 24285 5990
rect 24285 5983 24313 5990
rect 24325 5983 24357 5990
rect 24357 5983 24377 5990
rect 24389 5983 24391 5990
rect 24391 5983 24429 5990
rect 24429 5983 24441 5990
rect 24453 5983 24463 5990
rect 24463 5983 24501 5990
rect 24501 5983 24505 5990
rect 23941 5956 23959 5970
rect 23959 5956 23993 5970
rect 24005 5956 24031 5970
rect 24031 5956 24057 5970
rect 23941 5918 23993 5956
rect 24005 5918 24057 5956
rect 24069 5956 24103 5970
rect 24103 5956 24121 5970
rect 24069 5918 24121 5956
rect 24133 5956 24141 5970
rect 24141 5956 24175 5970
rect 24175 5956 24185 5970
rect 24133 5918 24185 5956
rect 24197 5956 24213 5970
rect 24213 5956 24247 5970
rect 24247 5956 24249 5970
rect 24197 5918 24249 5956
rect 24261 5956 24285 5970
rect 24285 5956 24313 5970
rect 24325 5956 24357 5970
rect 24357 5956 24377 5970
rect 24389 5956 24391 5970
rect 24391 5956 24429 5970
rect 24429 5956 24441 5970
rect 24453 5956 24463 5970
rect 24463 5956 24501 5970
rect 24501 5956 24505 5970
rect 24261 5918 24313 5956
rect 24325 5918 24377 5956
rect 24389 5918 24441 5956
rect 24453 5918 24505 5956
rect 23941 5883 23959 5905
rect 23959 5883 23993 5905
rect 24005 5883 24031 5905
rect 24031 5883 24057 5905
rect 23941 5853 23993 5883
rect 24005 5853 24057 5883
rect 24069 5883 24103 5905
rect 24103 5883 24121 5905
rect 24069 5853 24121 5883
rect 24133 5883 24141 5905
rect 24141 5883 24175 5905
rect 24175 5883 24185 5905
rect 24133 5853 24185 5883
rect 24197 5883 24213 5905
rect 24213 5883 24247 5905
rect 24247 5883 24249 5905
rect 24197 5853 24249 5883
rect 24261 5883 24285 5905
rect 24285 5883 24313 5905
rect 24325 5883 24357 5905
rect 24357 5883 24377 5905
rect 24389 5883 24391 5905
rect 24391 5883 24429 5905
rect 24429 5883 24441 5905
rect 24453 5883 24463 5905
rect 24463 5883 24501 5905
rect 24501 5883 24505 5905
rect 24261 5853 24313 5883
rect 24325 5853 24377 5883
rect 24389 5853 24441 5883
rect 24453 5853 24505 5883
rect 23941 5810 23959 5840
rect 23959 5810 23993 5840
rect 24005 5810 24031 5840
rect 24031 5810 24057 5840
rect 23941 5788 23993 5810
rect 24005 5788 24057 5810
rect 24069 5810 24103 5840
rect 24103 5810 24121 5840
rect 24069 5788 24121 5810
rect 24133 5810 24141 5840
rect 24141 5810 24175 5840
rect 24175 5810 24185 5840
rect 24133 5788 24185 5810
rect 24197 5810 24213 5840
rect 24213 5810 24247 5840
rect 24247 5810 24249 5840
rect 24197 5788 24249 5810
rect 24261 5810 24285 5840
rect 24285 5810 24313 5840
rect 24325 5810 24357 5840
rect 24357 5810 24377 5840
rect 24389 5810 24391 5840
rect 24391 5810 24429 5840
rect 24429 5810 24441 5840
rect 24453 5810 24463 5840
rect 24463 5810 24501 5840
rect 24501 5810 24505 5840
rect 24261 5788 24313 5810
rect 24325 5788 24377 5810
rect 24389 5788 24441 5810
rect 24453 5788 24505 5810
rect 23941 5771 23993 5775
rect 24005 5771 24057 5775
rect 23941 5737 23959 5771
rect 23959 5737 23993 5771
rect 24005 5737 24031 5771
rect 24031 5737 24057 5771
rect 23941 5723 23993 5737
rect 24005 5723 24057 5737
rect 24069 5771 24121 5775
rect 24069 5737 24103 5771
rect 24103 5737 24121 5771
rect 24069 5723 24121 5737
rect 24133 5771 24185 5775
rect 24133 5737 24141 5771
rect 24141 5737 24175 5771
rect 24175 5737 24185 5771
rect 24133 5723 24185 5737
rect 24197 5771 24249 5775
rect 24197 5737 24213 5771
rect 24213 5737 24247 5771
rect 24247 5737 24249 5771
rect 24197 5723 24249 5737
rect 24261 5771 24313 5775
rect 24325 5771 24377 5775
rect 24389 5771 24441 5775
rect 24453 5771 24505 5775
rect 24261 5737 24285 5771
rect 24285 5737 24313 5771
rect 24325 5737 24357 5771
rect 24357 5737 24377 5771
rect 24389 5737 24391 5771
rect 24391 5737 24429 5771
rect 24429 5737 24441 5771
rect 24453 5737 24463 5771
rect 24463 5737 24501 5771
rect 24501 5737 24505 5771
rect 24261 5723 24313 5737
rect 24325 5723 24377 5737
rect 24389 5723 24441 5737
rect 24453 5723 24505 5737
rect 23941 5698 23993 5710
rect 24005 5698 24057 5710
rect 24069 5698 24121 5710
rect 23941 5664 23959 5698
rect 23959 5664 23981 5698
rect 23941 5658 23981 5664
rect 23981 5658 23993 5698
rect 24005 5658 24057 5698
rect 24069 5664 24103 5698
rect 24103 5664 24121 5698
rect 24069 5658 24087 5664
rect 24087 5658 24121 5664
rect 24133 5698 24185 5710
rect 24133 5664 24141 5698
rect 24141 5664 24175 5698
rect 24175 5664 24185 5698
rect 24133 5658 24185 5664
rect 24197 5698 24249 5710
rect 24197 5664 24213 5698
rect 24213 5664 24247 5698
rect 24247 5664 24249 5698
rect 24197 5658 24249 5664
rect 24261 5698 24313 5710
rect 24325 5698 24377 5710
rect 24389 5698 24441 5710
rect 24453 5698 24505 5710
rect 24261 5664 24285 5698
rect 24285 5664 24313 5698
rect 24325 5664 24357 5698
rect 24357 5664 24377 5698
rect 24389 5664 24391 5698
rect 24391 5664 24429 5698
rect 24429 5664 24441 5698
rect 24453 5664 24463 5698
rect 24463 5664 24501 5698
rect 24501 5664 24505 5698
rect 24261 5658 24313 5664
rect 24325 5658 24377 5664
rect 24389 5658 24441 5664
rect 24453 5658 24505 5664
rect 17487 5375 17539 5427
rect 17551 5375 17603 5427
rect 20514 5375 20566 5427
rect 20578 5375 20630 5427
rect 12419 5232 12471 5284
rect 12490 5232 12542 5284
rect 12561 5232 12613 5284
rect 12632 5232 12684 5284
rect 12703 5232 12755 5284
rect 12773 5232 12825 5284
rect 12419 5168 12471 5220
rect 12490 5168 12542 5220
rect 12561 5168 12613 5220
rect 12632 5168 12684 5220
rect 12703 5168 12755 5220
rect 12773 5168 12825 5220
rect 16551 5193 16603 5245
rect 16551 5126 16603 5178
rect 16874 5190 16926 5242
rect 16874 5126 16926 5178
rect 20214 5078 20266 5130
rect 20278 5078 20330 5130
rect 14223 4992 14275 5044
rect 14290 4992 14342 5044
rect 16932 4985 16984 5037
rect 16996 4985 17048 5037
rect 20214 4973 20266 5025
rect 20278 4973 20330 5025
rect 13322 4624 13374 4676
rect 13389 4624 13441 4676
rect 14200 4624 14252 4676
rect 14267 4624 14319 4676
rect 12419 4495 12471 4547
rect 12490 4495 12542 4547
rect 12561 4495 12613 4547
rect 12632 4495 12684 4547
rect 12703 4495 12755 4547
rect 12773 4495 12825 4547
rect 12419 4431 12471 4483
rect 12490 4431 12542 4483
rect 12561 4431 12613 4483
rect 12632 4431 12684 4483
rect 12703 4431 12755 4483
rect 12773 4431 12825 4483
rect 14340 4269 14456 4385
rect 5862 4017 5978 4133
rect 16898 4210 16950 4262
rect 16962 4256 17014 4262
rect 16962 4222 16973 4256
rect 16973 4222 17007 4256
rect 17007 4222 17014 4256
rect 16962 4210 17014 4222
rect 22947 4212 22999 4264
rect 23011 4212 23063 4264
rect 23075 4212 23127 4264
rect 23139 4212 23191 4264
rect 17487 4093 17539 4145
rect 17551 4093 17603 4145
rect 12592 4059 12644 4063
rect 12684 4059 12736 4063
rect 12775 4059 12827 4063
rect 12592 4011 12594 4059
rect 12594 4011 12644 4059
rect 12684 4011 12736 4059
rect 12775 4011 12827 4059
rect 15705 4005 15757 4057
rect 12592 3947 12594 3999
rect 12594 3947 12644 3999
rect 12684 3947 12736 3999
rect 12775 3947 12827 3999
rect 15705 3941 15757 3993
rect 12592 3883 12594 3935
rect 12594 3883 12644 3935
rect 12684 3883 12736 3935
rect 12775 3883 12827 3935
rect 15705 3877 15757 3929
rect 15723 3765 15775 3769
rect 12592 3731 12594 3764
rect 12594 3731 12628 3764
rect 12628 3731 12644 3764
rect 12684 3731 12701 3764
rect 12701 3731 12736 3764
rect 12775 3731 12813 3764
rect 12813 3731 12827 3764
rect 15723 3731 15733 3765
rect 15733 3731 15767 3765
rect 15767 3731 15775 3765
rect 12592 3712 12644 3731
rect 12684 3712 12736 3731
rect 12775 3712 12827 3731
rect 15723 3717 15775 3731
rect 15787 3765 15839 3769
rect 15851 3765 15903 3769
rect 15915 3765 15967 3769
rect 15979 3765 16031 3769
rect 16043 3765 16095 3769
rect 16107 3765 16159 3769
rect 15787 3731 15806 3765
rect 15806 3731 15839 3765
rect 15851 3731 15879 3765
rect 15879 3731 15903 3765
rect 15915 3731 15952 3765
rect 15952 3731 15967 3765
rect 15979 3731 15986 3765
rect 15986 3731 16025 3765
rect 16025 3731 16031 3765
rect 16043 3731 16059 3765
rect 16059 3731 16095 3765
rect 16107 3731 16132 3765
rect 16132 3731 16159 3765
rect 15787 3717 15839 3731
rect 15851 3717 15903 3731
rect 15915 3717 15967 3731
rect 15979 3717 16031 3731
rect 16043 3717 16095 3731
rect 16107 3717 16159 3731
rect 16171 3765 16223 3769
rect 16171 3731 16205 3765
rect 16205 3731 16223 3765
rect 16171 3717 16223 3731
rect 16235 3765 16287 3769
rect 16235 3731 16244 3765
rect 16244 3731 16278 3765
rect 16278 3731 16287 3765
rect 16235 3717 16287 3731
rect 16299 3765 16351 3769
rect 16299 3731 16317 3765
rect 16317 3731 16351 3765
rect 16299 3717 16351 3731
rect 16363 3765 16415 3769
rect 16363 3731 16390 3765
rect 16390 3731 16415 3765
rect 16363 3717 16415 3731
rect 2104 3594 2156 3646
rect 2168 3594 2220 3646
rect 2232 3594 2284 3646
rect 2296 3594 2348 3646
rect 2360 3594 2412 3646
rect 2424 3594 2476 3646
rect 5344 3594 5396 3646
rect 5408 3594 5460 3646
rect 5472 3594 5524 3646
rect 12592 3693 12644 3700
rect 12684 3693 12736 3700
rect 12775 3693 12827 3700
rect 15723 3693 15775 3704
rect 12592 3659 12594 3693
rect 12594 3659 12628 3693
rect 12628 3659 12644 3693
rect 12684 3659 12701 3693
rect 12701 3659 12736 3693
rect 12775 3659 12813 3693
rect 12813 3659 12827 3693
rect 15723 3659 15733 3693
rect 15733 3659 15767 3693
rect 15767 3659 15775 3693
rect 12592 3648 12644 3659
rect 12684 3648 12736 3659
rect 12775 3648 12827 3659
rect 15723 3652 15775 3659
rect 15787 3693 15839 3704
rect 15851 3693 15903 3704
rect 15915 3693 15967 3704
rect 15979 3693 16031 3704
rect 16043 3693 16095 3704
rect 16107 3693 16159 3704
rect 15787 3659 15806 3693
rect 15806 3659 15839 3693
rect 15851 3659 15879 3693
rect 15879 3659 15903 3693
rect 15915 3659 15952 3693
rect 15952 3659 15967 3693
rect 15979 3659 15986 3693
rect 15986 3659 16025 3693
rect 16025 3659 16031 3693
rect 16043 3659 16059 3693
rect 16059 3659 16095 3693
rect 16107 3659 16132 3693
rect 16132 3659 16159 3693
rect 15787 3652 15839 3659
rect 15851 3652 15903 3659
rect 15915 3652 15967 3659
rect 15979 3652 16031 3659
rect 16043 3652 16095 3659
rect 16107 3652 16159 3659
rect 16171 3693 16223 3704
rect 16171 3659 16205 3693
rect 16205 3659 16223 3693
rect 16171 3652 16223 3659
rect 16235 3693 16287 3704
rect 16235 3659 16244 3693
rect 16244 3659 16278 3693
rect 16278 3659 16287 3693
rect 16235 3652 16287 3659
rect 16299 3693 16351 3704
rect 16299 3659 16317 3693
rect 16317 3659 16351 3693
rect 16299 3652 16351 3659
rect 16363 3693 16415 3704
rect 16363 3659 16390 3693
rect 16390 3659 16415 3693
rect 16363 3652 16415 3659
rect 12592 3621 12644 3636
rect 12684 3621 12736 3636
rect 12775 3621 12827 3636
rect 15723 3621 15775 3639
rect 12592 3587 12594 3621
rect 12594 3587 12628 3621
rect 12628 3587 12644 3621
rect 12684 3587 12701 3621
rect 12701 3587 12736 3621
rect 12775 3587 12813 3621
rect 12813 3587 12827 3621
rect 15723 3587 15733 3621
rect 15733 3587 15767 3621
rect 15767 3587 15775 3621
rect 15787 3621 15839 3639
rect 15851 3621 15903 3639
rect 15915 3621 15967 3639
rect 15979 3621 16031 3639
rect 16043 3621 16095 3639
rect 16107 3621 16159 3639
rect 15787 3587 15806 3621
rect 15806 3587 15839 3621
rect 15851 3587 15879 3621
rect 15879 3587 15903 3621
rect 15915 3587 15952 3621
rect 15952 3587 15967 3621
rect 15979 3587 15986 3621
rect 15986 3587 16025 3621
rect 16025 3587 16031 3621
rect 16043 3587 16059 3621
rect 16059 3587 16095 3621
rect 16107 3587 16132 3621
rect 16132 3587 16159 3621
rect 16171 3621 16223 3639
rect 16171 3587 16205 3621
rect 16205 3587 16223 3621
rect 16235 3621 16287 3639
rect 16235 3587 16244 3621
rect 16244 3587 16278 3621
rect 16278 3587 16287 3621
rect 16299 3621 16351 3639
rect 16299 3587 16317 3621
rect 16317 3587 16351 3621
rect 16363 3621 16415 3639
rect 16363 3587 16390 3621
rect 16390 3587 16415 3621
rect 12592 3584 12644 3587
rect 12684 3584 12736 3587
rect 12775 3584 12827 3587
rect 19979 3750 20031 3802
rect 19979 3685 20031 3737
rect 19979 3620 20031 3672
rect 19979 3555 20031 3607
rect 19979 3490 20031 3542
rect 15723 3471 15775 3475
rect 12411 3416 12463 3468
rect 12484 3416 12536 3468
rect 12556 3437 12594 3468
rect 12594 3437 12608 3468
rect 12628 3437 12667 3468
rect 12667 3437 12680 3468
rect 12700 3437 12701 3468
rect 12701 3437 12740 3468
rect 12740 3437 12752 3468
rect 12772 3437 12774 3468
rect 12774 3437 12813 3468
rect 12813 3437 12824 3468
rect 15723 3437 15733 3471
rect 15733 3437 15767 3471
rect 15767 3437 15775 3471
rect 12556 3416 12608 3437
rect 12628 3416 12680 3437
rect 12700 3416 12752 3437
rect 12772 3416 12824 3437
rect 15723 3423 15775 3437
rect 15787 3471 15839 3475
rect 15851 3471 15903 3475
rect 15915 3471 15967 3475
rect 15979 3471 16031 3475
rect 16043 3471 16095 3475
rect 16107 3471 16159 3475
rect 15787 3437 15806 3471
rect 15806 3437 15839 3471
rect 15851 3437 15879 3471
rect 15879 3437 15903 3471
rect 15915 3437 15952 3471
rect 15952 3437 15967 3471
rect 15979 3437 15986 3471
rect 15986 3437 16025 3471
rect 16025 3437 16031 3471
rect 16043 3437 16059 3471
rect 16059 3437 16095 3471
rect 16107 3437 16132 3471
rect 16132 3437 16159 3471
rect 15787 3423 15839 3437
rect 15851 3423 15903 3437
rect 15915 3423 15967 3437
rect 15979 3423 16031 3437
rect 16043 3423 16095 3437
rect 16107 3423 16159 3437
rect 16171 3471 16223 3475
rect 16171 3437 16205 3471
rect 16205 3437 16223 3471
rect 16171 3423 16223 3437
rect 16235 3471 16287 3475
rect 16235 3437 16244 3471
rect 16244 3437 16278 3471
rect 16278 3437 16287 3471
rect 16235 3423 16287 3437
rect 16299 3471 16351 3475
rect 16299 3437 16317 3471
rect 16317 3437 16351 3471
rect 16299 3423 16351 3437
rect 16363 3471 16415 3475
rect 16363 3437 16390 3471
rect 16390 3437 16415 3471
rect 16363 3423 16415 3437
rect 12411 3352 12463 3404
rect 12484 3352 12536 3404
rect 12556 3399 12608 3404
rect 12628 3399 12680 3404
rect 12700 3399 12752 3404
rect 12772 3399 12824 3404
rect 15723 3399 15775 3406
rect 12556 3365 12594 3399
rect 12594 3365 12608 3399
rect 12628 3365 12667 3399
rect 12667 3365 12680 3399
rect 12700 3365 12701 3399
rect 12701 3365 12740 3399
rect 12740 3365 12752 3399
rect 12772 3365 12774 3399
rect 12774 3365 12813 3399
rect 12813 3365 12824 3399
rect 15723 3365 15733 3399
rect 15733 3365 15767 3399
rect 15767 3365 15775 3399
rect 12556 3352 12608 3365
rect 12628 3352 12680 3365
rect 12700 3352 12752 3365
rect 12772 3352 12824 3365
rect 15723 3354 15775 3365
rect 15787 3399 15839 3406
rect 15851 3399 15903 3406
rect 15915 3399 15967 3406
rect 15979 3399 16031 3406
rect 16043 3399 16095 3406
rect 16107 3399 16159 3406
rect 15787 3365 15806 3399
rect 15806 3365 15839 3399
rect 15851 3365 15879 3399
rect 15879 3365 15903 3399
rect 15915 3365 15952 3399
rect 15952 3365 15967 3399
rect 15979 3365 15986 3399
rect 15986 3365 16025 3399
rect 16025 3365 16031 3399
rect 16043 3365 16059 3399
rect 16059 3365 16095 3399
rect 16107 3365 16132 3399
rect 16132 3365 16159 3399
rect 15787 3354 15839 3365
rect 15851 3354 15903 3365
rect 15915 3354 15967 3365
rect 15979 3354 16031 3365
rect 16043 3354 16095 3365
rect 16107 3354 16159 3365
rect 16171 3399 16223 3406
rect 16171 3365 16205 3399
rect 16205 3365 16223 3399
rect 16171 3354 16223 3365
rect 16235 3399 16287 3406
rect 16235 3365 16244 3399
rect 16244 3365 16278 3399
rect 16278 3365 16287 3399
rect 16235 3354 16287 3365
rect 16299 3399 16351 3406
rect 16299 3365 16317 3399
rect 16317 3365 16351 3399
rect 16299 3354 16351 3365
rect 16363 3399 16415 3406
rect 16363 3365 16390 3399
rect 16390 3365 16415 3399
rect 16363 3354 16415 3365
rect 12411 3288 12463 3340
rect 12484 3288 12536 3340
rect 12556 3327 12608 3340
rect 12628 3327 12680 3340
rect 12700 3327 12752 3340
rect 12772 3327 12824 3340
rect 15723 3327 15775 3337
rect 12556 3293 12594 3327
rect 12594 3293 12608 3327
rect 12628 3293 12667 3327
rect 12667 3293 12680 3327
rect 12700 3293 12701 3327
rect 12701 3293 12740 3327
rect 12740 3293 12752 3327
rect 12772 3293 12774 3327
rect 12774 3293 12813 3327
rect 12813 3293 12824 3327
rect 15723 3293 15733 3327
rect 15733 3293 15767 3327
rect 15767 3293 15775 3327
rect 12556 3288 12608 3293
rect 12628 3288 12680 3293
rect 12700 3288 12752 3293
rect 12772 3288 12824 3293
rect 15723 3285 15775 3293
rect 15787 3327 15839 3337
rect 15851 3327 15903 3337
rect 15915 3327 15967 3337
rect 15979 3327 16031 3337
rect 16043 3327 16095 3337
rect 16107 3327 16159 3337
rect 15787 3293 15806 3327
rect 15806 3293 15839 3327
rect 15851 3293 15879 3327
rect 15879 3293 15903 3327
rect 15915 3293 15952 3327
rect 15952 3293 15967 3327
rect 15979 3293 15986 3327
rect 15986 3293 16025 3327
rect 16025 3293 16031 3327
rect 16043 3293 16059 3327
rect 16059 3293 16095 3327
rect 16107 3293 16132 3327
rect 16132 3293 16159 3327
rect 15787 3285 15839 3293
rect 15851 3285 15903 3293
rect 15915 3285 15967 3293
rect 15979 3285 16031 3293
rect 16043 3285 16095 3293
rect 16107 3285 16159 3293
rect 16171 3327 16223 3337
rect 16171 3293 16205 3327
rect 16205 3293 16223 3327
rect 16171 3285 16223 3293
rect 16235 3327 16287 3337
rect 16235 3293 16244 3327
rect 16244 3293 16278 3327
rect 16278 3293 16287 3327
rect 16235 3285 16287 3293
rect 16299 3327 16351 3337
rect 16299 3293 16317 3327
rect 16317 3293 16351 3327
rect 16299 3285 16351 3293
rect 16363 3327 16415 3337
rect 16363 3293 16390 3327
rect 16390 3293 16415 3327
rect 16363 3285 16415 3293
rect 12411 3224 12463 3276
rect 12484 3224 12536 3276
rect 12556 3255 12608 3276
rect 12628 3255 12680 3276
rect 12700 3255 12752 3276
rect 12772 3255 12824 3276
rect 15723 3255 15775 3268
rect 12556 3224 12594 3255
rect 12594 3224 12608 3255
rect 12628 3224 12667 3255
rect 12667 3224 12680 3255
rect 12700 3224 12701 3255
rect 12701 3224 12740 3255
rect 12740 3224 12752 3255
rect 12772 3224 12774 3255
rect 12774 3224 12813 3255
rect 12813 3224 12824 3255
rect 15723 3221 15733 3255
rect 15733 3221 15767 3255
rect 15767 3221 15775 3255
rect 15723 3216 15775 3221
rect 15787 3255 15839 3268
rect 15851 3255 15903 3268
rect 15915 3255 15967 3268
rect 15979 3255 16031 3268
rect 16043 3255 16095 3268
rect 16107 3255 16159 3268
rect 15787 3221 15806 3255
rect 15806 3221 15839 3255
rect 15851 3221 15879 3255
rect 15879 3221 15903 3255
rect 15915 3221 15952 3255
rect 15952 3221 15967 3255
rect 15979 3221 15986 3255
rect 15986 3221 16025 3255
rect 16025 3221 16031 3255
rect 16043 3221 16059 3255
rect 16059 3221 16095 3255
rect 16107 3221 16132 3255
rect 16132 3221 16159 3255
rect 15787 3216 15839 3221
rect 15851 3216 15903 3221
rect 15915 3216 15967 3221
rect 15979 3216 16031 3221
rect 16043 3216 16095 3221
rect 16107 3216 16159 3221
rect 16171 3255 16223 3268
rect 16171 3221 16205 3255
rect 16205 3221 16223 3255
rect 16171 3216 16223 3221
rect 16235 3255 16287 3268
rect 16235 3221 16244 3255
rect 16244 3221 16278 3255
rect 16278 3221 16287 3255
rect 16235 3216 16287 3221
rect 16299 3255 16351 3268
rect 16299 3221 16317 3255
rect 16317 3221 16351 3255
rect 16299 3216 16351 3221
rect 16363 3255 16415 3268
rect 16363 3221 16390 3255
rect 16390 3221 16415 3255
rect 16363 3216 16415 3221
rect 19979 3424 20031 3476
rect 19979 3358 20031 3410
rect 19979 3292 20031 3344
rect 19979 3226 20031 3278
rect 4372 3154 4424 3206
rect 4436 3154 4488 3206
rect 19979 3160 20031 3212
rect 19979 3094 20031 3146
rect 19979 3028 20031 3080
rect 19979 2962 20031 3014
rect 19979 2896 20031 2948
rect 2104 2712 2156 2764
rect 2168 2712 2220 2764
rect 2232 2712 2284 2764
rect 2296 2712 2348 2764
rect 2360 2712 2412 2764
rect 2424 2712 2476 2764
rect 7730 2721 7782 2773
rect 7794 2721 7846 2773
rect 12414 2668 12421 2701
rect 12421 2668 12462 2701
rect 12462 2668 12466 2701
rect 12486 2668 12496 2701
rect 12496 2668 12537 2701
rect 12537 2668 12538 2701
rect 12558 2668 12571 2701
rect 12571 2668 12610 2701
rect 12630 2668 12646 2701
rect 12646 2668 12682 2701
rect 12702 2668 12721 2701
rect 12721 2668 12754 2701
rect 12774 2668 12796 2701
rect 12796 2668 12826 2701
rect 12414 2649 12466 2668
rect 12486 2649 12538 2668
rect 12558 2649 12610 2668
rect 12630 2649 12682 2668
rect 12702 2649 12754 2668
rect 12774 2649 12826 2668
rect 13292 2734 13344 2786
rect 13356 2734 13408 2786
rect 14340 2761 14456 2877
rect 17487 2794 17539 2846
rect 17551 2794 17603 2846
rect 19979 2830 20031 2882
rect 19979 2764 20031 2816
rect 13292 2667 13344 2719
rect 13356 2667 13408 2719
rect 19979 2698 20031 2750
rect 12414 2630 12466 2637
rect 12486 2630 12538 2637
rect 12558 2630 12610 2637
rect 12630 2630 12682 2637
rect 12702 2630 12754 2637
rect 12774 2630 12826 2637
rect 19979 2632 20031 2684
rect 12414 2596 12421 2630
rect 12421 2596 12462 2630
rect 12462 2596 12466 2630
rect 12486 2596 12496 2630
rect 12496 2596 12537 2630
rect 12537 2596 12538 2630
rect 12558 2596 12571 2630
rect 12571 2596 12610 2630
rect 12630 2596 12646 2630
rect 12646 2596 12682 2630
rect 12702 2596 12721 2630
rect 12721 2596 12754 2630
rect 12774 2596 12796 2630
rect 12796 2596 12826 2630
rect 12414 2585 12466 2596
rect 12486 2585 12538 2596
rect 12558 2585 12610 2596
rect 12630 2585 12682 2596
rect 12702 2585 12754 2596
rect 12774 2585 12826 2596
rect 12414 2558 12466 2573
rect 12486 2558 12538 2573
rect 12558 2558 12610 2573
rect 12630 2558 12682 2573
rect 12702 2558 12754 2573
rect 12774 2558 12826 2573
rect 12414 2524 12421 2558
rect 12421 2524 12462 2558
rect 12462 2524 12466 2558
rect 12486 2524 12496 2558
rect 12496 2524 12537 2558
rect 12537 2524 12538 2558
rect 12558 2524 12571 2558
rect 12571 2524 12610 2558
rect 12630 2524 12646 2558
rect 12646 2524 12682 2558
rect 12702 2524 12721 2558
rect 12721 2524 12754 2558
rect 12774 2524 12796 2558
rect 12796 2524 12826 2558
rect 12414 2521 12466 2524
rect 12486 2521 12538 2524
rect 12558 2521 12610 2524
rect 12630 2521 12682 2524
rect 12702 2521 12754 2524
rect 12774 2521 12826 2524
rect 13416 2506 13468 2558
rect 13480 2506 13532 2558
rect 13416 2439 13468 2491
rect 13480 2439 13532 2491
rect 16501 2465 16553 2517
rect 16565 2465 16617 2517
rect 17269 2516 17385 2632
rect 19979 2566 20031 2618
rect 19979 2500 20031 2552
rect 20077 3750 20129 3802
rect 20077 3685 20129 3737
rect 20077 3620 20129 3672
rect 20077 3555 20129 3607
rect 20077 3490 20129 3542
rect 20077 3424 20129 3476
rect 20077 3358 20129 3410
rect 20077 3292 20129 3344
rect 20077 3226 20129 3278
rect 20077 3160 20129 3212
rect 20077 3094 20129 3146
rect 20077 3028 20129 3080
rect 20077 2962 20129 3014
rect 20077 2896 20129 2948
rect 20077 2830 20129 2882
rect 20077 2764 20129 2816
rect 20077 2698 20129 2750
rect 20077 2632 20129 2684
rect 20077 2566 20129 2618
rect 20077 2500 20129 2552
rect 5862 2215 5978 2331
rect 13235 2338 13287 2390
rect 13299 2338 13351 2390
rect 13235 2271 13287 2323
rect 13299 2271 13351 2323
rect 12412 2120 12443 2143
rect 12443 2120 12464 2143
rect 12486 2120 12516 2143
rect 12516 2120 12538 2143
rect 12560 2120 12589 2143
rect 12589 2120 12612 2143
rect 12634 2120 12662 2143
rect 12662 2120 12686 2143
rect 12707 2120 12735 2143
rect 12735 2120 12759 2143
rect 12780 2120 12808 2143
rect 12808 2120 12832 2143
rect 12412 2091 12464 2120
rect 12486 2091 12538 2120
rect 12560 2091 12612 2120
rect 12634 2091 12686 2120
rect 12707 2091 12759 2120
rect 12780 2091 12832 2120
rect 12412 2048 12443 2079
rect 12443 2048 12464 2079
rect 12486 2048 12516 2079
rect 12516 2048 12538 2079
rect 12560 2048 12589 2079
rect 12589 2048 12612 2079
rect 12634 2048 12662 2079
rect 12662 2048 12686 2079
rect 12707 2048 12735 2079
rect 12735 2048 12759 2079
rect 12780 2048 12808 2079
rect 12808 2048 12832 2079
rect 12412 2027 12464 2048
rect 12486 2027 12538 2048
rect 12560 2027 12612 2048
rect 12634 2027 12686 2048
rect 12707 2027 12759 2048
rect 12780 2027 12832 2048
rect 12412 2010 12464 2015
rect 12486 2010 12538 2015
rect 12560 2010 12612 2015
rect 12634 2010 12686 2015
rect 12707 2010 12759 2015
rect 12780 2010 12832 2015
rect 12412 1976 12443 2010
rect 12443 1976 12464 2010
rect 12486 1976 12516 2010
rect 12516 1976 12538 2010
rect 12560 1976 12589 2010
rect 12589 1976 12612 2010
rect 12634 1976 12662 2010
rect 12662 1976 12686 2010
rect 12707 1976 12735 2010
rect 12735 1976 12759 2010
rect 12780 1976 12808 2010
rect 12808 1976 12832 2010
rect 12412 1963 12464 1976
rect 12486 1963 12538 1976
rect 12560 1963 12612 1976
rect 12634 1963 12686 1976
rect 12707 1963 12759 1976
rect 12780 1963 12832 1976
rect 12412 1938 12464 1951
rect 12486 1938 12538 1951
rect 12560 1938 12612 1951
rect 12634 1938 12686 1951
rect 12707 1938 12759 1951
rect 12780 1938 12832 1951
rect 12412 1904 12443 1938
rect 12443 1904 12464 1938
rect 12486 1904 12516 1938
rect 12516 1904 12538 1938
rect 12560 1904 12589 1938
rect 12589 1904 12612 1938
rect 12634 1904 12662 1938
rect 12662 1904 12686 1938
rect 12707 1904 12735 1938
rect 12735 1904 12759 1938
rect 12780 1904 12808 1938
rect 12808 1904 12832 1938
rect 12412 1899 12464 1904
rect 12486 1899 12538 1904
rect 12560 1899 12612 1904
rect 12634 1899 12686 1904
rect 12707 1899 12759 1904
rect 12780 1899 12832 1904
rect 2104 1786 2156 1838
rect 2168 1786 2220 1838
rect 2232 1786 2284 1838
rect 2296 1786 2348 1838
rect 2360 1786 2412 1838
rect 2424 1786 2476 1838
rect 8146 1795 8198 1847
rect 8210 1795 8262 1847
rect 12412 1866 12464 1887
rect 12486 1866 12538 1887
rect 12560 1866 12612 1887
rect 12634 1866 12686 1887
rect 12707 1866 12759 1887
rect 12780 1866 12832 1887
rect 12412 1835 12443 1866
rect 12443 1835 12464 1866
rect 12486 1835 12516 1866
rect 12516 1835 12538 1866
rect 12560 1835 12589 1866
rect 12589 1835 12612 1866
rect 12634 1835 12662 1866
rect 12662 1835 12686 1866
rect 12707 1835 12735 1866
rect 12735 1835 12759 1866
rect 12780 1835 12808 1866
rect 12808 1835 12832 1866
rect 12412 1794 12464 1823
rect 12486 1794 12538 1823
rect 12560 1794 12612 1823
rect 12634 1794 12686 1823
rect 12707 1794 12759 1823
rect 12780 1794 12832 1823
rect 12412 1771 12443 1794
rect 12443 1771 12464 1794
rect 12486 1771 12516 1794
rect 12516 1771 12538 1794
rect 12560 1771 12589 1794
rect 12589 1771 12612 1794
rect 12634 1771 12662 1794
rect 12662 1771 12686 1794
rect 12707 1771 12735 1794
rect 12735 1771 12759 1794
rect 12780 1771 12808 1794
rect 12808 1771 12832 1794
rect 17428 1795 17480 1847
rect 17492 1795 17544 1847
rect 17556 1795 17608 1847
rect 17428 1683 17480 1735
rect 17492 1683 17544 1735
rect 17556 1683 17608 1735
rect 12409 1510 12461 1562
rect 12484 1510 12536 1562
rect 12559 1510 12611 1562
rect 12634 1510 12686 1562
rect 12709 1510 12761 1562
rect 12784 1510 12836 1562
rect 25701 1548 25753 1600
rect 12409 1446 12461 1498
rect 12484 1446 12536 1498
rect 12559 1446 12611 1498
rect 12634 1446 12686 1498
rect 12709 1446 12761 1498
rect 12784 1446 12836 1498
rect 4372 1338 4424 1390
rect 4436 1338 4488 1390
rect 25701 1473 25753 1525
rect 25701 1397 25753 1449
rect 23577 1033 23757 1213
rect 23577 969 23693 1033
rect 23577 944 23629 957
rect 23577 910 23605 944
rect 23605 910 23629 944
rect 23577 905 23629 910
rect 27015 1120 27067 1172
rect 27090 1120 27142 1172
rect 27165 1120 27217 1172
rect 27240 1120 27292 1172
rect 27314 1120 27366 1172
rect 27015 1056 27067 1108
rect 27090 1056 27142 1108
rect 27165 1056 27217 1108
rect 27240 1056 27292 1108
rect 27314 1056 27366 1108
rect 27015 992 27067 1044
rect 27090 992 27142 1044
rect 27165 992 27217 1044
rect 27240 992 27292 1044
rect 27314 992 27366 1044
rect 27015 928 27067 980
rect 27090 928 27142 980
rect 27165 928 27217 980
rect 27240 928 27292 980
rect 27314 928 27366 980
<< metal2 >>
rect 23743 13310 23795 13316
tri 23795 13275 23829 13309 sw
rect 23795 13258 29168 13275
rect 23743 13256 29168 13258
tri 29168 13256 29187 13275 sw
rect 23743 13246 29187 13256
rect 23795 13223 29187 13246
rect 23743 13188 23795 13194
tri 23795 13189 23829 13223 nw
tri 29146 13189 29180 13223 ne
rect 29180 13189 29187 13223
tri 29180 13188 29181 13189 ne
rect 29181 13188 29187 13189
tri 29187 13188 29255 13256 sw
tri 29181 13182 29187 13188 ne
rect 29187 13182 29255 13188
tri 29255 13182 29261 13188 sw
tri 29187 13108 29261 13182 ne
tri 29261 13108 29335 13182 sw
tri 29261 13086 29283 13108 ne
rect 24392 12365 24721 12603
tri 27147 11955 27203 12011 sw
rect 27147 11917 29057 11955
tri 29057 11917 29095 11955 sw
rect 27147 11903 29095 11917
tri 29035 11843 29095 11903 ne
tri 29095 11843 29169 11917 sw
tri 29095 11769 29169 11843 ne
tri 29169 11769 29243 11843 sw
tri 29169 11747 29191 11769 ne
rect 24229 10991 24281 10997
tri 24281 10957 24315 10991 sw
rect 24281 10939 24741 10957
rect 24229 10927 24741 10939
rect 24281 10905 24741 10927
rect 24793 10905 24805 10957
rect 24857 10905 24881 10957
rect 27434 10905 27440 10957
rect 27492 10905 27504 10957
rect 27556 10922 28968 10957
tri 28968 10922 29003 10957 sw
rect 27556 10905 29003 10922
tri 29003 10905 29020 10922 sw
rect 24281 10875 24282 10905
rect 24229 10872 24282 10875
tri 24282 10872 24315 10905 nw
tri 28946 10872 28979 10905 ne
rect 28979 10872 29020 10905
rect 24229 10869 24281 10872
tri 24281 10871 24282 10872 nw
rect 25294 10812 25300 10864
rect 25352 10812 25364 10864
rect 25416 10812 25422 10864
rect 25666 10812 25672 10864
rect 25724 10812 25736 10864
rect 25788 10812 25794 10864
rect 25993 10820 25999 10872
rect 26051 10820 26091 10872
rect 26143 10820 26183 10872
rect 26235 10820 26275 10872
rect 26327 10820 26367 10872
rect 26419 10820 26425 10872
tri 28979 10869 28982 10872 ne
rect 28982 10869 29020 10872
tri 29020 10869 29056 10905 sw
tri 28982 10864 28987 10869 ne
rect 28987 10864 29056 10869
tri 29056 10864 29061 10869 sw
tri 28987 10848 29003 10864 ne
rect 29003 10848 29061 10864
tri 29061 10848 29077 10864 sw
tri 29003 10820 29031 10848 ne
rect 29031 10820 29077 10848
tri 29031 10812 29039 10820 ne
rect 29039 10812 29077 10820
tri 29077 10812 29113 10848 sw
tri 25299 10779 25332 10812 ne
rect 25332 10779 25385 10812
tri 25385 10779 25418 10812 nw
tri 25671 10779 25704 10812 ne
rect 25704 10779 25756 10812
rect 25332 10684 25384 10779
tri 25384 10778 25385 10779 nw
tri 25704 10778 25705 10779 ne
tri 25299 10556 25332 10589 se
rect 25332 10556 25384 10682
tri 25189 10504 25241 10556 se
rect 25241 10504 25262 10556
rect 25314 10504 25326 10556
rect 25378 10504 25384 10556
tri 25543 10556 25577 10590 sw
tri 25671 10556 25705 10590 se
rect 25705 10556 25756 10779
tri 25756 10778 25790 10812 nw
tri 29039 10778 29073 10812 ne
rect 29073 10778 29113 10812
tri 29073 10774 29077 10778 ne
rect 29077 10774 29113 10778
tri 29113 10774 29151 10812 sw
tri 29077 10752 29099 10774 ne
tri 25756 10556 25790 10590 sw
rect 25543 10504 25711 10556
rect 25763 10504 25775 10556
rect 25827 10504 25833 10556
rect 27499 10504 27505 10556
rect 27557 10504 27569 10556
rect 27621 10504 28904 10556
tri 28904 10504 28956 10556 sw
tri 25155 10470 25189 10504 se
rect 25189 10470 25254 10504
tri 25254 10470 25288 10504 nw
rect 25543 10493 25566 10504
tri 25566 10493 25577 10504 nw
tri 28864 10493 28875 10504 ne
rect 28875 10493 28956 10504
tri 28956 10493 28967 10504 sw
tri 25543 10470 25566 10493 nw
tri 28875 10470 28898 10493 ne
rect 28898 10470 28967 10493
tri 25149 10464 25155 10470 se
rect 25155 10464 25248 10470
tri 25248 10464 25254 10470 nw
tri 28898 10464 28904 10470 ne
rect 28904 10464 28967 10470
tri 25142 10457 25149 10464 se
rect 25149 10457 25241 10464
tri 25241 10457 25248 10464 nw
tri 28904 10457 28911 10464 ne
rect 28911 10457 28967 10464
tri 25135 10450 25142 10457 se
rect 25142 10450 25234 10457
tri 25234 10450 25241 10457 nw
tri 28911 10450 28918 10457 ne
rect 28918 10450 28967 10457
tri 25129 10444 25135 10450 se
rect 25135 10444 25228 10450
tri 25228 10444 25234 10450 nw
rect 25757 10444 25818 10450
tri 25077 10392 25129 10444 se
rect 25129 10392 25176 10444
tri 25176 10392 25228 10444 nw
rect 25757 10392 25762 10444
rect 25814 10392 25818 10444
tri 28918 10401 28967 10450 ne
tri 28967 10401 29059 10493 sw
tri 25064 10379 25077 10392 se
rect 25077 10379 25163 10392
tri 25163 10379 25176 10392 nw
rect 25757 10379 25818 10392
tri 25060 10375 25064 10379 se
rect 25064 10375 25159 10379
tri 25159 10375 25163 10379 nw
tri 25026 10263 25060 10297 se
rect 25060 10263 25124 10375
tri 25124 10340 25159 10375 nw
rect 25757 10327 25762 10379
rect 25814 10327 25818 10379
tri 28967 10373 28995 10401 ne
rect 25757 10314 25818 10327
rect 20256 10262 25124 10263
tri 25124 10262 25125 10263 sw
rect 25757 10262 25762 10314
rect 25814 10262 25818 10314
rect 20256 10248 25125 10262
tri 25125 10248 25139 10262 sw
rect 25757 10248 25818 10262
rect 20256 10196 25139 10248
tri 25139 10196 25191 10248 sw
rect 25757 10196 25762 10248
rect 25814 10196 25818 10248
rect 25993 10225 26429 10300
rect 20256 10183 25191 10196
tri 25191 10183 25204 10196 sw
rect 17018 9635 17024 9687
rect 17076 9635 17090 9687
rect 17142 9635 17156 9687
rect 17208 9635 17222 9687
rect 17274 9635 17288 9687
rect 17340 9635 17354 9687
rect 17406 9635 17420 9687
rect 17472 9635 17486 9687
rect 17538 9635 17552 9687
rect 17604 9635 17618 9687
rect 17670 9635 17684 9687
rect 17736 9635 17750 9687
rect 17802 9635 17816 9687
rect 17868 9635 17882 9687
rect 17934 9635 17948 9687
rect 18000 9635 18014 9687
rect 18066 9635 18080 9687
rect 18132 9635 18146 9687
rect 18198 9635 18212 9687
rect 18264 9635 18278 9687
rect 18330 9635 18344 9687
rect 18396 9635 18410 9687
rect 18462 9635 18476 9687
rect 18528 9635 18542 9687
rect 18594 9635 18607 9687
rect 18659 9635 18672 9687
rect 18724 9635 18737 9687
rect 18789 9635 18802 9687
rect 18854 9635 18867 9687
rect 18919 9635 18932 9687
rect 18984 9635 18997 9687
rect 19049 9635 19062 9687
rect 19114 9635 19127 9687
rect 19179 9635 19192 9687
rect 19244 9635 19257 9687
rect 19309 9635 19315 9687
rect 17018 9623 19315 9635
rect 17018 9571 17024 9623
rect 17076 9571 17090 9623
rect 17142 9571 17156 9623
rect 17208 9571 17222 9623
rect 17274 9571 17288 9623
rect 17340 9571 17354 9623
rect 17406 9571 17420 9623
rect 17472 9571 17486 9623
rect 17538 9571 17552 9623
rect 17604 9571 17618 9623
rect 17670 9571 17684 9623
rect 17736 9571 17750 9623
rect 17802 9571 17816 9623
rect 17868 9571 17882 9623
rect 17934 9571 17948 9623
rect 18000 9571 18014 9623
rect 18066 9571 18080 9623
rect 18132 9571 18146 9623
rect 18198 9571 18212 9623
rect 18264 9571 18278 9623
rect 18330 9571 18344 9623
rect 18396 9571 18410 9623
rect 18462 9571 18476 9623
rect 18528 9571 18542 9623
rect 18594 9571 18607 9623
rect 18659 9571 18672 9623
rect 18724 9571 18737 9623
rect 18789 9571 18802 9623
rect 18854 9571 18867 9623
rect 18919 9571 18932 9623
rect 18984 9571 18997 9623
rect 19049 9571 19062 9623
rect 19114 9571 19127 9623
rect 19179 9571 19192 9623
rect 19244 9571 19257 9623
rect 19309 9571 19315 9623
rect 15699 8825 16439 9470
rect 17018 9069 17198 9571
tri 17198 9546 17223 9571 nw
tri 17523 9546 17548 9571 ne
tri 17198 9069 17223 9094 sw
tri 17523 9069 17548 9094 se
rect 17548 9069 17728 9571
tri 17728 9546 17753 9571 nw
tri 18041 9546 18066 9571 ne
tri 17728 9069 17753 9094 sw
tri 18041 9069 18066 9094 se
rect 18066 9069 18246 9571
tri 18246 9546 18271 9571 nw
tri 18584 9546 18609 9571 ne
tri 18246 9069 18271 9094 sw
tri 18584 9069 18609 9094 se
rect 18609 9069 18789 9571
tri 18789 9546 18814 9571 nw
tri 19110 9546 19135 9571 ne
tri 18789 9069 18814 9094 sw
tri 19110 9069 19135 9094 se
rect 19135 9069 19315 9571
rect 17018 9017 17029 9069
rect 17081 9017 17095 9069
rect 17147 9017 17161 9069
rect 17213 9017 17227 9069
rect 17279 9017 17293 9069
rect 17345 9017 17359 9069
rect 17411 9017 17425 9069
rect 17477 9017 17491 9069
rect 17543 9017 17557 9069
rect 17609 9017 17623 9069
rect 17675 9017 17689 9069
rect 17741 9017 17755 9069
rect 17807 9017 17821 9069
rect 17873 9017 17887 9069
rect 17939 9017 17953 9069
rect 18005 9017 18019 9069
rect 18071 9017 18085 9069
rect 18137 9017 18151 9069
rect 18203 9017 18217 9069
rect 18269 9017 18282 9069
rect 18334 9017 18347 9069
rect 18399 9017 18412 9069
rect 18464 9017 18477 9069
rect 18529 9017 18542 9069
rect 18594 9017 18607 9069
rect 18659 9017 18672 9069
rect 18724 9017 18737 9069
rect 18789 9017 18802 9069
rect 18854 9017 18867 9069
rect 18919 9017 18932 9069
rect 18984 9017 18997 9069
rect 19049 9017 19062 9069
rect 19114 9017 19127 9069
rect 19179 9017 19192 9069
rect 19244 9017 19257 9069
rect 19309 9017 19315 9069
rect 17018 9005 19315 9017
rect 17018 8953 17029 9005
rect 17081 8953 17095 9005
rect 17147 8953 17161 9005
rect 17213 8953 17227 9005
rect 17279 8953 17293 9005
rect 17345 8953 17359 9005
rect 17411 8953 17425 9005
rect 17477 8953 17491 9005
rect 17543 8953 17557 9005
rect 17609 8953 17623 9005
rect 17675 8953 17689 9005
rect 17741 8953 17755 9005
rect 17807 8953 17821 9005
rect 17873 8953 17887 9005
rect 17939 8953 17953 9005
rect 18005 8953 18019 9005
rect 18071 8953 18085 9005
rect 18137 8953 18151 9005
rect 18203 8953 18217 9005
rect 18269 8953 18282 9005
rect 18334 8953 18347 9005
rect 18399 8953 18412 9005
rect 18464 8953 18477 9005
rect 18529 8953 18542 9005
rect 18594 8953 18607 9005
rect 18659 8953 18672 9005
rect 18724 8953 18737 9005
rect 18789 8953 18802 9005
rect 18854 8953 18867 9005
rect 18919 8953 18932 9005
rect 18984 8953 18997 9005
rect 19049 8953 19062 9005
rect 19114 8953 19127 9005
rect 19179 8953 19192 9005
rect 19244 8953 19257 9005
rect 19309 8953 19315 9005
rect 17018 8941 17211 8953
tri 17211 8941 17223 8953 nw
tri 17523 8941 17535 8953 ne
rect 17535 8941 17741 8953
tri 17741 8941 17753 8953 nw
tri 18041 8941 18053 8953 ne
rect 18053 8941 18259 8953
tri 18259 8941 18271 8953 nw
tri 18584 8941 18596 8953 ne
rect 18596 8941 18802 8953
tri 18802 8941 18814 8953 nw
tri 19110 8941 19122 8953 ne
rect 19122 8941 19315 8953
tri 16439 8825 16453 8839 sw
tri 17004 8825 17018 8839 se
rect 17018 8825 17198 8941
tri 17198 8928 17211 8941 nw
tri 17535 8928 17548 8941 ne
tri 17198 8825 17212 8839 sw
tri 17534 8825 17548 8839 se
rect 17548 8825 17728 8941
tri 17728 8928 17741 8941 nw
tri 18053 8928 18066 8941 ne
tri 17728 8825 17742 8839 sw
tri 18052 8825 18066 8839 se
rect 18066 8825 18246 8941
tri 18246 8928 18259 8941 nw
tri 18596 8928 18609 8941 ne
tri 18246 8825 18260 8839 sw
tri 18595 8825 18609 8839 se
rect 18609 8825 18789 8941
tri 18789 8928 18802 8941 nw
tri 19122 8928 19135 8941 ne
tri 18789 8825 18803 8839 sw
tri 19121 8825 19135 8839 se
rect 19135 8825 19315 8941
rect 15699 8814 16453 8825
tri 16453 8814 16464 8825 sw
tri 16993 8814 17004 8825 se
rect 17004 8814 17212 8825
tri 17212 8814 17223 8825 sw
tri 17523 8814 17534 8825 se
rect 17534 8814 17742 8825
tri 17742 8814 17753 8825 sw
tri 18041 8814 18052 8825 se
rect 18052 8814 18260 8825
tri 18260 8814 18271 8825 sw
tri 18584 8814 18595 8825 se
rect 18595 8814 18803 8825
tri 18803 8814 18814 8825 sw
tri 19110 8814 19121 8825 se
rect 19121 8814 19315 8825
rect 15699 8762 17029 8814
rect 17081 8762 17095 8814
rect 17147 8762 17161 8814
rect 17213 8762 17227 8814
rect 17279 8762 17293 8814
rect 17345 8762 17359 8814
rect 17411 8762 17425 8814
rect 17477 8762 17491 8814
rect 17543 8762 17557 8814
rect 17609 8762 17623 8814
rect 17675 8762 17689 8814
rect 17741 8762 17755 8814
rect 17807 8762 17821 8814
rect 17873 8762 17887 8814
rect 17939 8762 17953 8814
rect 18005 8762 18019 8814
rect 18071 8762 18085 8814
rect 18137 8762 18151 8814
rect 18203 8762 18217 8814
rect 18269 8762 18282 8814
rect 18334 8762 18347 8814
rect 18399 8762 18412 8814
rect 18464 8762 18477 8814
rect 18529 8762 18542 8814
rect 18594 8762 18607 8814
rect 18659 8762 18672 8814
rect 18724 8762 18737 8814
rect 18789 8762 18802 8814
rect 18854 8762 18867 8814
rect 18919 8762 18932 8814
rect 18984 8762 18997 8814
rect 19049 8762 19062 8814
rect 19114 8762 19127 8814
rect 19179 8762 19192 8814
rect 19244 8762 19257 8814
rect 19309 8762 19315 8814
rect 15699 8750 19315 8762
rect 15699 8698 17029 8750
rect 17081 8698 17095 8750
rect 17147 8698 17161 8750
rect 17213 8698 17227 8750
rect 17279 8698 17293 8750
rect 17345 8698 17359 8750
rect 17411 8698 17425 8750
rect 17477 8698 17491 8750
rect 17543 8698 17557 8750
rect 17609 8698 17623 8750
rect 17675 8698 17689 8750
rect 17741 8698 17755 8750
rect 17807 8698 17821 8750
rect 17873 8698 17887 8750
rect 17939 8698 17953 8750
rect 18005 8698 18019 8750
rect 18071 8698 18085 8750
rect 18137 8698 18151 8750
rect 18203 8698 18217 8750
rect 18269 8698 18282 8750
rect 18334 8698 18347 8750
rect 18399 8698 18412 8750
rect 18464 8698 18477 8750
rect 18529 8698 18542 8750
rect 18594 8698 18607 8750
rect 18659 8698 18672 8750
rect 18724 8698 18737 8750
rect 18789 8698 18802 8750
rect 18854 8698 18867 8750
rect 18919 8698 18932 8750
rect 18984 8698 18997 8750
rect 19049 8698 19062 8750
rect 19114 8698 19127 8750
rect 19179 8698 19192 8750
rect 19244 8698 19257 8750
rect 19309 8698 19315 8750
rect 15699 8686 19315 8698
rect 15699 8634 17029 8686
rect 17081 8634 17095 8686
rect 17147 8634 17161 8686
rect 17213 8634 17227 8686
rect 17279 8634 17293 8686
rect 17345 8634 17359 8686
rect 17411 8634 17425 8686
rect 17477 8634 17491 8686
rect 17543 8634 17557 8686
rect 17609 8634 17623 8686
rect 17675 8634 17689 8686
rect 17741 8634 17755 8686
rect 17807 8634 17821 8686
rect 17873 8634 17887 8686
rect 17939 8634 17953 8686
rect 18005 8634 18019 8686
rect 18071 8634 18085 8686
rect 18137 8634 18151 8686
rect 18203 8634 18217 8686
rect 18269 8634 18282 8686
rect 18334 8634 18347 8686
rect 18399 8634 18412 8686
rect 18464 8634 18477 8686
rect 18529 8634 18542 8686
rect 18594 8634 18607 8686
rect 18659 8634 18672 8686
rect 18724 8634 18737 8686
rect 18789 8634 18802 8686
rect 18854 8634 18867 8686
rect 18919 8634 18932 8686
rect 18984 8634 18997 8686
rect 19049 8634 19062 8686
rect 19114 8634 19127 8686
rect 19179 8634 19192 8686
rect 19244 8634 19257 8686
rect 19309 8634 19315 8686
rect 15699 8633 16463 8634
tri 16463 8633 16464 8634 nw
tri 16993 8633 16994 8634 ne
rect 16994 8633 17222 8634
tri 17222 8633 17223 8634 nw
tri 17523 8633 17524 8634 ne
rect 17524 8633 17752 8634
tri 17752 8633 17753 8634 nw
tri 18041 8633 18042 8634 ne
rect 18042 8633 18270 8634
tri 18270 8633 18271 8634 nw
tri 18584 8633 18585 8634 ne
rect 18585 8633 18813 8634
tri 18813 8633 18814 8634 nw
tri 19110 8633 19111 8634 ne
rect 19111 8633 19315 8634
rect 15699 8495 16439 8633
tri 16439 8609 16463 8633 nw
tri 16994 8609 17018 8633 ne
tri 16439 8495 16464 8520 sw
tri 16993 8495 17018 8520 se
rect 17018 8495 17198 8633
tri 17198 8609 17222 8633 nw
tri 17524 8609 17548 8633 ne
tri 17198 8495 17223 8520 sw
tri 17523 8495 17548 8520 se
rect 17548 8495 17728 8633
tri 17728 8609 17752 8633 nw
tri 18042 8609 18066 8633 ne
tri 17728 8495 17753 8520 sw
tri 18041 8495 18066 8520 se
rect 18066 8495 18246 8633
tri 18246 8609 18270 8633 nw
tri 18585 8609 18609 8633 ne
tri 18246 8495 18271 8520 sw
tri 18584 8495 18609 8520 se
rect 18609 8495 18789 8633
tri 18789 8609 18813 8633 nw
tri 19111 8609 19135 8633 ne
tri 18789 8495 18814 8520 sw
tri 19110 8495 19135 8520 se
rect 19135 8495 19315 8633
rect 15699 8443 17029 8495
rect 17081 8443 17095 8495
rect 17147 8443 17161 8495
rect 17213 8443 17227 8495
rect 17279 8443 17293 8495
rect 17345 8443 17359 8495
rect 17411 8443 17425 8495
rect 17477 8443 17491 8495
rect 17543 8443 17557 8495
rect 17609 8443 17623 8495
rect 17675 8443 17689 8495
rect 17741 8443 17755 8495
rect 17807 8443 17821 8495
rect 17873 8443 17887 8495
rect 17939 8443 17953 8495
rect 18005 8443 18019 8495
rect 18071 8443 18085 8495
rect 18137 8443 18151 8495
rect 18203 8443 18217 8495
rect 18269 8443 18282 8495
rect 18334 8443 18347 8495
rect 18399 8443 18412 8495
rect 18464 8443 18477 8495
rect 18529 8443 18542 8495
rect 18594 8443 18607 8495
rect 18659 8443 18672 8495
rect 18724 8443 18737 8495
rect 18789 8443 18802 8495
rect 18854 8443 18867 8495
rect 18919 8443 18932 8495
rect 18984 8443 18997 8495
rect 19049 8443 19062 8495
rect 19114 8443 19127 8495
rect 19179 8443 19192 8495
rect 19244 8443 19257 8495
rect 19309 8443 19315 8495
rect 15699 8431 19315 8443
rect 15699 8379 17029 8431
rect 17081 8379 17095 8431
rect 17147 8379 17161 8431
rect 17213 8379 17227 8431
rect 17279 8379 17293 8431
rect 17345 8379 17359 8431
rect 17411 8379 17425 8431
rect 17477 8379 17491 8431
rect 17543 8379 17557 8431
rect 17609 8379 17623 8431
rect 17675 8379 17689 8431
rect 17741 8379 17755 8431
rect 17807 8379 17821 8431
rect 17873 8379 17887 8431
rect 17939 8379 17953 8431
rect 18005 8379 18019 8431
rect 18071 8379 18085 8431
rect 18137 8379 18151 8431
rect 18203 8379 18217 8431
rect 18269 8379 18282 8431
rect 18334 8379 18347 8431
rect 18399 8379 18412 8431
rect 18464 8379 18477 8431
rect 18529 8379 18542 8431
rect 18594 8379 18607 8431
rect 18659 8379 18672 8431
rect 18724 8379 18737 8431
rect 18789 8379 18802 8431
rect 18854 8379 18867 8431
rect 18919 8379 18932 8431
rect 18984 8379 18997 8431
rect 19049 8379 19062 8431
rect 19114 8379 19127 8431
rect 19179 8379 19192 8431
rect 19244 8379 19257 8431
rect 19309 8379 19315 8431
rect 15699 8367 19315 8379
rect 15699 8315 17029 8367
rect 17081 8315 17095 8367
rect 17147 8315 17161 8367
rect 17213 8315 17227 8367
rect 17279 8315 17293 8367
rect 17345 8315 17359 8367
rect 17411 8315 17425 8367
rect 17477 8315 17491 8367
rect 17543 8315 17557 8367
rect 17609 8315 17623 8367
rect 17675 8315 17689 8367
rect 17741 8315 17755 8367
rect 17807 8315 17821 8367
rect 17873 8315 17887 8367
rect 17939 8315 17953 8367
rect 18005 8315 18019 8367
rect 18071 8315 18085 8367
rect 18137 8315 18151 8367
rect 18203 8315 18217 8367
rect 18269 8315 18282 8367
rect 18334 8315 18347 8367
rect 18399 8315 18412 8367
rect 18464 8315 18477 8367
rect 18529 8315 18542 8367
rect 18594 8315 18607 8367
rect 18659 8315 18672 8367
rect 18724 8315 18737 8367
rect 18789 8315 18802 8367
rect 18854 8315 18867 8367
rect 18919 8315 18932 8367
rect 18984 8315 18997 8367
rect 19049 8315 19062 8367
rect 19114 8315 19127 8367
rect 19179 8315 19192 8367
rect 19244 8315 19257 8367
rect 19309 8315 19315 8367
rect 15699 8231 16439 8315
tri 16439 8290 16464 8315 nw
tri 16993 8290 17018 8315 ne
tri 16439 8231 16464 8256 sw
tri 16993 8231 17018 8256 se
rect 17018 8231 17198 8315
tri 17198 8290 17223 8315 nw
tri 17523 8290 17548 8315 ne
tri 17198 8231 17223 8256 sw
tri 17523 8231 17548 8256 se
rect 17548 8231 17728 8315
tri 17728 8290 17753 8315 nw
tri 18041 8290 18066 8315 ne
tri 17728 8231 17753 8256 sw
tri 18041 8231 18066 8256 se
rect 18066 8231 18246 8315
tri 18246 8290 18271 8315 nw
tri 18584 8290 18609 8315 ne
tri 18246 8231 18271 8256 sw
tri 18584 8231 18609 8256 se
rect 18609 8231 18789 8315
tri 18789 8290 18814 8315 nw
tri 19110 8290 19135 8315 ne
tri 18789 8231 18814 8256 sw
tri 19110 8231 19135 8256 se
rect 19135 8231 19315 8315
rect 15699 8179 17029 8231
rect 17081 8179 17095 8231
rect 17147 8179 17161 8231
rect 17213 8179 17227 8231
rect 17279 8179 17293 8231
rect 17345 8179 17359 8231
rect 17411 8179 17425 8231
rect 17477 8179 17491 8231
rect 17543 8179 17557 8231
rect 17609 8179 17623 8231
rect 17675 8179 17689 8231
rect 17741 8179 17755 8231
rect 17807 8179 17821 8231
rect 17873 8179 17887 8231
rect 17939 8179 17953 8231
rect 18005 8179 18019 8231
rect 18071 8179 18085 8231
rect 18137 8179 18151 8231
rect 18203 8179 18217 8231
rect 18269 8179 18282 8231
rect 18334 8179 18347 8231
rect 18399 8179 18412 8231
rect 18464 8179 18477 8231
rect 18529 8179 18542 8231
rect 18594 8179 18607 8231
rect 18659 8179 18672 8231
rect 18724 8179 18737 8231
rect 18789 8179 18802 8231
rect 18854 8179 18867 8231
rect 18919 8179 18932 8231
rect 18984 8179 18997 8231
rect 19049 8179 19062 8231
rect 19114 8179 19127 8231
rect 19179 8179 19192 8231
rect 19244 8179 19257 8231
rect 19309 8179 19315 8231
rect 15699 8167 19315 8179
rect 15699 8115 17029 8167
rect 17081 8115 17095 8167
rect 17147 8115 17161 8167
rect 17213 8115 17227 8167
rect 17279 8115 17293 8167
rect 17345 8115 17359 8167
rect 17411 8115 17425 8167
rect 17477 8115 17491 8167
rect 17543 8115 17557 8167
rect 17609 8115 17623 8167
rect 17675 8115 17689 8167
rect 17741 8115 17755 8167
rect 17807 8115 17821 8167
rect 17873 8115 17887 8167
rect 17939 8115 17953 8167
rect 18005 8115 18019 8167
rect 18071 8115 18085 8167
rect 18137 8115 18151 8167
rect 18203 8115 18217 8167
rect 18269 8115 18282 8167
rect 18334 8115 18347 8167
rect 18399 8115 18412 8167
rect 18464 8115 18477 8167
rect 18529 8115 18542 8167
rect 18594 8115 18607 8167
rect 18659 8115 18672 8167
rect 18724 8115 18737 8167
rect 18789 8115 18802 8167
rect 18854 8115 18867 8167
rect 18919 8115 18932 8167
rect 18984 8115 18997 8167
rect 19049 8115 19062 8167
rect 19114 8115 19127 8167
rect 19179 8115 19192 8167
rect 19244 8115 19257 8167
rect 19309 8115 19315 8167
rect 15699 8103 19315 8115
rect 15699 8051 17029 8103
rect 17081 8051 17095 8103
rect 17147 8051 17161 8103
rect 17213 8051 17227 8103
rect 17279 8051 17293 8103
rect 17345 8051 17359 8103
rect 17411 8051 17425 8103
rect 17477 8051 17491 8103
rect 17543 8051 17557 8103
rect 17609 8051 17623 8103
rect 17675 8051 17689 8103
rect 17741 8051 17755 8103
rect 17807 8051 17821 8103
rect 17873 8051 17887 8103
rect 17939 8051 17953 8103
rect 18005 8051 18019 8103
rect 18071 8051 18085 8103
rect 18137 8051 18151 8103
rect 18203 8051 18217 8103
rect 18269 8051 18282 8103
rect 18334 8051 18347 8103
rect 18399 8051 18412 8103
rect 18464 8051 18477 8103
rect 18529 8051 18542 8103
rect 18594 8051 18607 8103
rect 18659 8051 18672 8103
rect 18724 8051 18737 8103
rect 18789 8051 18802 8103
rect 18854 8051 18867 8103
rect 18919 8051 18932 8103
rect 18984 8051 18997 8103
rect 19049 8051 19062 8103
rect 19114 8051 19127 8103
rect 19179 8051 19192 8103
rect 19244 8051 19257 8103
rect 19309 8051 19315 8103
rect 15699 7967 16439 8051
tri 16439 8026 16464 8051 nw
tri 16993 8026 17018 8051 ne
tri 16439 7967 16464 7992 sw
tri 16993 7967 17018 7992 se
rect 17018 7967 17198 8051
tri 17198 8026 17223 8051 nw
tri 17523 8026 17548 8051 ne
tri 17198 7967 17223 7992 sw
tri 17523 7967 17548 7992 se
rect 17548 7967 17728 8051
tri 17728 8026 17753 8051 nw
tri 18041 8026 18066 8051 ne
tri 17728 7967 17753 7992 sw
tri 18041 7967 18066 7992 se
rect 18066 7967 18246 8051
tri 18246 8026 18271 8051 nw
tri 18584 8026 18609 8051 ne
tri 18246 7967 18271 7992 sw
tri 18584 7967 18609 7992 se
rect 18609 7967 18789 8051
tri 18789 8026 18814 8051 nw
tri 19110 8026 19135 8051 ne
tri 18789 7967 18814 7992 sw
tri 19110 7967 19135 7992 se
rect 19135 7967 19315 8051
rect 15699 7915 17029 7967
rect 17081 7915 17095 7967
rect 17147 7915 17161 7967
rect 17213 7915 17227 7967
rect 17279 7915 17293 7967
rect 17345 7915 17359 7967
rect 17411 7915 17425 7967
rect 17477 7915 17491 7967
rect 17543 7915 17557 7967
rect 17609 7915 17623 7967
rect 17675 7915 17689 7967
rect 17741 7915 17755 7967
rect 17807 7915 17821 7967
rect 17873 7915 17887 7967
rect 17939 7915 17953 7967
rect 18005 7915 18019 7967
rect 18071 7915 18085 7967
rect 18137 7915 18151 7967
rect 18203 7915 18217 7967
rect 18269 7915 18282 7967
rect 18334 7915 18347 7967
rect 18399 7915 18412 7967
rect 18464 7915 18477 7967
rect 18529 7915 18542 7967
rect 18594 7915 18607 7967
rect 18659 7915 18672 7967
rect 18724 7915 18737 7967
rect 18789 7915 18802 7967
rect 18854 7915 18867 7967
rect 18919 7915 18932 7967
rect 18984 7915 18997 7967
rect 19049 7915 19062 7967
rect 19114 7915 19127 7967
rect 19179 7915 19192 7967
rect 19244 7915 19257 7967
rect 19309 7915 19315 7967
rect 15699 7903 19315 7915
rect 15699 7851 17029 7903
rect 17081 7851 17095 7903
rect 17147 7851 17161 7903
rect 17213 7851 17227 7903
rect 17279 7851 17293 7903
rect 17345 7851 17359 7903
rect 17411 7851 17425 7903
rect 17477 7851 17491 7903
rect 17543 7851 17557 7903
rect 17609 7851 17623 7903
rect 17675 7851 17689 7903
rect 17741 7851 17755 7903
rect 17807 7851 17821 7903
rect 17873 7851 17887 7903
rect 17939 7851 17953 7903
rect 18005 7851 18019 7903
rect 18071 7851 18085 7903
rect 18137 7851 18151 7903
rect 18203 7851 18217 7903
rect 18269 7851 18282 7903
rect 18334 7851 18347 7903
rect 18399 7851 18412 7903
rect 18464 7851 18477 7903
rect 18529 7851 18542 7903
rect 18594 7851 18607 7903
rect 18659 7851 18672 7903
rect 18724 7851 18737 7903
rect 18789 7851 18802 7903
rect 18854 7851 18867 7903
rect 18919 7851 18932 7903
rect 18984 7851 18997 7903
rect 19049 7851 19062 7903
rect 19114 7851 19127 7903
rect 19179 7851 19192 7903
rect 19244 7851 19257 7903
rect 19309 7851 19315 7903
rect 15699 7839 19315 7851
rect 15699 7787 17029 7839
rect 17081 7787 17095 7839
rect 17147 7787 17161 7839
rect 17213 7787 17227 7839
rect 17279 7787 17293 7839
rect 17345 7787 17359 7839
rect 17411 7787 17425 7839
rect 17477 7787 17491 7839
rect 17543 7787 17557 7839
rect 17609 7787 17623 7839
rect 17675 7787 17689 7839
rect 17741 7787 17755 7839
rect 17807 7787 17821 7839
rect 17873 7787 17887 7839
rect 17939 7787 17953 7839
rect 18005 7787 18019 7839
rect 18071 7787 18085 7839
rect 18137 7787 18151 7839
rect 18203 7787 18217 7839
rect 18269 7787 18282 7839
rect 18334 7787 18347 7839
rect 18399 7787 18412 7839
rect 18464 7787 18477 7839
rect 18529 7787 18542 7839
rect 18594 7787 18607 7839
rect 18659 7787 18672 7839
rect 18724 7787 18737 7839
rect 18789 7787 18802 7839
rect 18854 7787 18867 7839
rect 18919 7787 18932 7839
rect 18984 7787 18997 7839
rect 19049 7787 19062 7839
rect 19114 7787 19127 7839
rect 19179 7787 19192 7839
rect 19244 7787 19257 7839
rect 19309 7787 19315 7839
rect 15699 7703 16439 7787
tri 16439 7762 16464 7787 nw
tri 16993 7762 17018 7787 ne
tri 16439 7703 16464 7728 sw
tri 16993 7703 17018 7728 se
rect 17018 7703 17198 7787
tri 17198 7762 17223 7787 nw
tri 17523 7762 17548 7787 ne
tri 17198 7703 17223 7728 sw
tri 17523 7703 17548 7728 se
rect 17548 7703 17728 7787
tri 17728 7762 17753 7787 nw
tri 18041 7762 18066 7787 ne
tri 17728 7703 17753 7728 sw
tri 18041 7703 18066 7728 se
rect 18066 7703 18246 7787
tri 18246 7762 18271 7787 nw
tri 18584 7762 18609 7787 ne
tri 18246 7703 18271 7728 sw
tri 18584 7703 18609 7728 se
rect 18609 7703 18789 7787
tri 18789 7762 18814 7787 nw
tri 19110 7762 19135 7787 ne
tri 18789 7703 18814 7728 sw
tri 19110 7703 19135 7728 se
rect 19135 7703 19315 7787
rect 15699 7651 17029 7703
rect 17081 7651 17095 7703
rect 17147 7651 17161 7703
rect 17213 7651 17227 7703
rect 17279 7651 17293 7703
rect 17345 7651 17359 7703
rect 17411 7651 17425 7703
rect 17477 7651 17491 7703
rect 17543 7651 17557 7703
rect 17609 7651 17623 7703
rect 17675 7651 17689 7703
rect 17741 7651 17755 7703
rect 17807 7651 17821 7703
rect 17873 7651 17887 7703
rect 17939 7651 17953 7703
rect 18005 7651 18019 7703
rect 18071 7651 18085 7703
rect 18137 7651 18151 7703
rect 18203 7651 18217 7703
rect 18269 7651 18282 7703
rect 18334 7651 18347 7703
rect 18399 7651 18412 7703
rect 18464 7651 18477 7703
rect 18529 7651 18542 7703
rect 18594 7651 18607 7703
rect 18659 7651 18672 7703
rect 18724 7651 18737 7703
rect 18789 7651 18802 7703
rect 18854 7651 18867 7703
rect 18919 7651 18932 7703
rect 18984 7651 18997 7703
rect 19049 7651 19062 7703
rect 19114 7651 19127 7703
rect 19179 7651 19192 7703
rect 19244 7651 19257 7703
rect 19309 7651 19315 7703
rect 15699 7639 19315 7651
rect 15699 7587 17029 7639
rect 17081 7587 17095 7639
rect 17147 7587 17161 7639
rect 17213 7587 17227 7639
rect 17279 7587 17293 7639
rect 17345 7587 17359 7639
rect 17411 7587 17425 7639
rect 17477 7587 17491 7639
rect 17543 7587 17557 7639
rect 17609 7587 17623 7639
rect 17675 7587 17689 7639
rect 17741 7587 17755 7639
rect 17807 7587 17821 7639
rect 17873 7587 17887 7639
rect 17939 7587 17953 7639
rect 18005 7587 18019 7639
rect 18071 7587 18085 7639
rect 18137 7587 18151 7639
rect 18203 7587 18217 7639
rect 18269 7587 18282 7639
rect 18334 7587 18347 7639
rect 18399 7587 18412 7639
rect 18464 7587 18477 7639
rect 18529 7587 18542 7639
rect 18594 7587 18607 7639
rect 18659 7587 18672 7639
rect 18724 7587 18737 7639
rect 18789 7587 18802 7639
rect 18854 7587 18867 7639
rect 18919 7587 18932 7639
rect 18984 7587 18997 7639
rect 19049 7587 19062 7639
rect 19114 7587 19127 7639
rect 19179 7587 19192 7639
rect 19244 7587 19257 7639
rect 19309 7587 19315 7639
rect 15699 7575 19315 7587
rect 15699 7523 17029 7575
rect 17081 7523 17095 7575
rect 17147 7523 17161 7575
rect 17213 7523 17227 7575
rect 17279 7523 17293 7575
rect 17345 7523 17359 7575
rect 17411 7523 17425 7575
rect 17477 7523 17491 7575
rect 17543 7523 17557 7575
rect 17609 7523 17623 7575
rect 17675 7523 17689 7575
rect 17741 7523 17755 7575
rect 17807 7523 17821 7575
rect 17873 7523 17887 7575
rect 17939 7523 17953 7575
rect 18005 7523 18019 7575
rect 18071 7523 18085 7575
rect 18137 7523 18151 7575
rect 18203 7523 18217 7575
rect 18269 7523 18282 7575
rect 18334 7523 18347 7575
rect 18399 7523 18412 7575
rect 18464 7523 18477 7575
rect 18529 7523 18542 7575
rect 18594 7523 18607 7575
rect 18659 7523 18672 7575
rect 18724 7523 18737 7575
rect 18789 7523 18802 7575
rect 18854 7523 18867 7575
rect 18919 7523 18932 7575
rect 18984 7523 18997 7575
rect 19049 7523 19062 7575
rect 19114 7523 19127 7575
rect 19179 7523 19192 7575
rect 19244 7523 19257 7575
rect 19309 7523 19315 7575
rect 15699 7439 16439 7523
tri 16439 7498 16464 7523 nw
tri 16993 7498 17018 7523 ne
tri 16439 7439 16464 7464 sw
tri 16993 7439 17018 7464 se
rect 17018 7439 17198 7523
tri 17198 7498 17223 7523 nw
tri 17523 7498 17548 7523 ne
tri 17198 7439 17223 7464 sw
tri 17523 7439 17548 7464 se
rect 17548 7439 17728 7523
tri 17728 7498 17753 7523 nw
tri 18041 7498 18066 7523 ne
tri 17728 7439 17753 7464 sw
tri 18041 7439 18066 7464 se
rect 18066 7439 18246 7523
tri 18246 7498 18271 7523 nw
tri 18584 7498 18609 7523 ne
tri 18246 7439 18271 7464 sw
tri 18584 7439 18609 7464 se
rect 18609 7439 18789 7523
tri 18789 7498 18814 7523 nw
tri 19110 7498 19135 7523 ne
tri 18789 7439 18814 7464 sw
tri 19110 7439 19135 7464 se
rect 19135 7439 19315 7523
rect 15699 7387 17029 7439
rect 17081 7387 17095 7439
rect 17147 7387 17161 7439
rect 17213 7387 17227 7439
rect 17279 7387 17293 7439
rect 17345 7387 17359 7439
rect 17411 7387 17425 7439
rect 17477 7387 17491 7439
rect 17543 7387 17557 7439
rect 17609 7387 17623 7439
rect 17675 7387 17689 7439
rect 17741 7387 17755 7439
rect 17807 7387 17821 7439
rect 17873 7387 17887 7439
rect 17939 7387 17953 7439
rect 18005 7387 18019 7439
rect 18071 7387 18085 7439
rect 18137 7387 18151 7439
rect 18203 7387 18217 7439
rect 18269 7387 18282 7439
rect 18334 7387 18347 7439
rect 18399 7387 18412 7439
rect 18464 7387 18477 7439
rect 18529 7387 18542 7439
rect 18594 7387 18607 7439
rect 18659 7387 18672 7439
rect 18724 7387 18737 7439
rect 18789 7387 18802 7439
rect 18854 7387 18867 7439
rect 18919 7387 18932 7439
rect 18984 7387 18997 7439
rect 19049 7387 19062 7439
rect 19114 7387 19127 7439
rect 19179 7387 19192 7439
rect 19244 7387 19257 7439
rect 19309 7387 19315 7439
rect 15699 7375 19315 7387
rect 15699 7323 17029 7375
rect 17081 7323 17095 7375
rect 17147 7323 17161 7375
rect 17213 7323 17227 7375
rect 17279 7323 17293 7375
rect 17345 7323 17359 7375
rect 17411 7323 17425 7375
rect 17477 7323 17491 7375
rect 17543 7323 17557 7375
rect 17609 7323 17623 7375
rect 17675 7323 17689 7375
rect 17741 7323 17755 7375
rect 17807 7323 17821 7375
rect 17873 7323 17887 7375
rect 17939 7323 17953 7375
rect 18005 7323 18019 7375
rect 18071 7323 18085 7375
rect 18137 7323 18151 7375
rect 18203 7323 18217 7375
rect 18269 7323 18282 7375
rect 18334 7323 18347 7375
rect 18399 7323 18412 7375
rect 18464 7323 18477 7375
rect 18529 7323 18542 7375
rect 18594 7323 18607 7375
rect 18659 7323 18672 7375
rect 18724 7323 18737 7375
rect 18789 7323 18802 7375
rect 18854 7323 18867 7375
rect 18919 7323 18932 7375
rect 18984 7323 18997 7375
rect 19049 7323 19062 7375
rect 19114 7323 19127 7375
rect 19179 7323 19192 7375
rect 19244 7323 19257 7375
rect 19309 7323 19315 7375
rect 15699 7311 19315 7323
rect 15699 7259 17029 7311
rect 17081 7259 17095 7311
rect 17147 7259 17161 7311
rect 17213 7259 17227 7311
rect 17279 7259 17293 7311
rect 17345 7259 17359 7311
rect 17411 7259 17425 7311
rect 17477 7259 17491 7311
rect 17543 7259 17557 7311
rect 17609 7259 17623 7311
rect 17675 7259 17689 7311
rect 17741 7259 17755 7311
rect 17807 7259 17821 7311
rect 17873 7259 17887 7311
rect 17939 7259 17953 7311
rect 18005 7259 18019 7311
rect 18071 7259 18085 7311
rect 18137 7259 18151 7311
rect 18203 7259 18217 7311
rect 18269 7259 18282 7311
rect 18334 7259 18347 7311
rect 18399 7259 18412 7311
rect 18464 7259 18477 7311
rect 18529 7259 18542 7311
rect 18594 7259 18607 7311
rect 18659 7259 18672 7311
rect 18724 7259 18737 7311
rect 18789 7259 18802 7311
rect 18854 7259 18867 7311
rect 18919 7259 18932 7311
rect 18984 7259 18997 7311
rect 19049 7259 19062 7311
rect 19114 7259 19127 7311
rect 19179 7259 19192 7311
rect 19244 7259 19257 7311
rect 19309 7259 19315 7311
rect 15699 7175 16439 7259
tri 16439 7234 16464 7259 nw
tri 16993 7234 17018 7259 ne
tri 16439 7175 16464 7200 sw
tri 16993 7175 17018 7200 se
rect 17018 7175 17198 7259
tri 17198 7234 17223 7259 nw
tri 17523 7234 17548 7259 ne
tri 17198 7175 17223 7200 sw
tri 17523 7175 17548 7200 se
rect 17548 7175 17728 7259
tri 17728 7234 17753 7259 nw
tri 18041 7234 18066 7259 ne
tri 17728 7175 17753 7200 sw
tri 18041 7175 18066 7200 se
rect 18066 7175 18246 7259
tri 18246 7234 18271 7259 nw
tri 18584 7234 18609 7259 ne
tri 18246 7175 18271 7200 sw
tri 18584 7175 18609 7200 se
rect 18609 7175 18789 7259
tri 18789 7234 18814 7259 nw
tri 19110 7234 19135 7259 ne
tri 18789 7175 18814 7200 sw
tri 19110 7175 19135 7200 se
rect 19135 7175 19315 7259
rect 15699 7123 17029 7175
rect 17081 7123 17095 7175
rect 17147 7123 17161 7175
rect 17213 7123 17227 7175
rect 17279 7123 17293 7175
rect 17345 7123 17359 7175
rect 17411 7123 17425 7175
rect 17477 7123 17491 7175
rect 17543 7123 17557 7175
rect 17609 7123 17623 7175
rect 17675 7123 17689 7175
rect 17741 7123 17755 7175
rect 17807 7123 17821 7175
rect 17873 7123 17887 7175
rect 17939 7123 17953 7175
rect 18005 7123 18019 7175
rect 18071 7123 18085 7175
rect 18137 7123 18151 7175
rect 18203 7123 18217 7175
rect 18269 7123 18282 7175
rect 18334 7123 18347 7175
rect 18399 7123 18412 7175
rect 18464 7123 18477 7175
rect 18529 7123 18542 7175
rect 18594 7123 18607 7175
rect 18659 7123 18672 7175
rect 18724 7123 18737 7175
rect 18789 7123 18802 7175
rect 18854 7123 18867 7175
rect 18919 7123 18932 7175
rect 18984 7123 18997 7175
rect 19049 7123 19062 7175
rect 19114 7123 19127 7175
rect 19179 7123 19192 7175
rect 19244 7123 19257 7175
rect 19309 7123 19315 7175
rect 15699 7111 19315 7123
rect 15699 7059 17029 7111
rect 17081 7059 17095 7111
rect 17147 7059 17161 7111
rect 17213 7059 17227 7111
rect 17279 7059 17293 7111
rect 17345 7059 17359 7111
rect 17411 7059 17425 7111
rect 17477 7059 17491 7111
rect 17543 7059 17557 7111
rect 17609 7059 17623 7111
rect 17675 7059 17689 7111
rect 17741 7059 17755 7111
rect 17807 7059 17821 7111
rect 17873 7059 17887 7111
rect 17939 7059 17953 7111
rect 18005 7059 18019 7111
rect 18071 7059 18085 7111
rect 18137 7059 18151 7111
rect 18203 7059 18217 7111
rect 18269 7059 18282 7111
rect 18334 7059 18347 7111
rect 18399 7059 18412 7111
rect 18464 7059 18477 7111
rect 18529 7059 18542 7111
rect 18594 7059 18607 7111
rect 18659 7059 18672 7111
rect 18724 7059 18737 7111
rect 18789 7059 18802 7111
rect 18854 7059 18867 7111
rect 18919 7059 18932 7111
rect 18984 7059 18997 7111
rect 19049 7059 19062 7111
rect 19114 7059 19127 7111
rect 19179 7059 19192 7111
rect 19244 7059 19257 7111
rect 19309 7059 19315 7111
rect 15699 7047 19315 7059
rect 15699 6995 17029 7047
rect 17081 6995 17095 7047
rect 17147 6995 17161 7047
rect 17213 6995 17227 7047
rect 17279 6995 17293 7047
rect 17345 6995 17359 7047
rect 17411 6995 17425 7047
rect 17477 6995 17491 7047
rect 17543 6995 17557 7047
rect 17609 6995 17623 7047
rect 17675 6995 17689 7047
rect 17741 6995 17755 7047
rect 17807 6995 17821 7047
rect 17873 6995 17887 7047
rect 17939 6995 17953 7047
rect 18005 6995 18019 7047
rect 18071 6995 18085 7047
rect 18137 6995 18151 7047
rect 18203 6995 18217 7047
rect 18269 6995 18282 7047
rect 18334 6995 18347 7047
rect 18399 6995 18412 7047
rect 18464 6995 18477 7047
rect 18529 6995 18542 7047
rect 18594 6995 18607 7047
rect 18659 6995 18672 7047
rect 18724 6995 18737 7047
rect 18789 6995 18802 7047
rect 18854 6995 18867 7047
rect 18919 6995 18932 7047
rect 18984 6995 18997 7047
rect 19049 6995 19062 7047
rect 19114 6995 19127 7047
rect 19179 6995 19192 7047
rect 19244 6995 19257 7047
rect 19309 6995 19315 7047
rect 12403 5284 12842 5292
rect 12403 5232 12419 5284
rect 12471 5232 12490 5284
rect 12542 5232 12561 5284
rect 12613 5232 12632 5284
rect 12684 5232 12703 5284
rect 12755 5232 12773 5284
rect 12825 5232 12842 5284
rect 12403 5220 12842 5232
rect 12403 5168 12419 5220
rect 12471 5168 12490 5220
rect 12542 5168 12561 5220
rect 12613 5168 12632 5220
rect 12684 5168 12703 5220
rect 12755 5168 12773 5220
rect 12825 5168 12842 5220
rect 5862 4133 5978 4139
rect -232 4011 4975 4014
tri 4975 4011 4978 4014 sw
rect -232 4005 4978 4011
tri 4978 4005 4984 4011 sw
rect -232 3999 4984 4005
tri 4984 3999 4990 4005 sw
rect -232 3962 4990 3999
tri 4953 3947 4968 3962 ne
rect 4968 3947 4990 3962
tri 4990 3947 5042 3999 sw
tri 4968 3942 4973 3947 ne
rect 4973 3942 5042 3947
tri 5042 3942 5047 3947 sw
tri 4973 3941 4974 3942 ne
rect 4974 3941 5047 3942
tri 5047 3941 5048 3942 sw
tri 4974 3940 4975 3941 ne
rect 4975 3940 5048 3941
tri 4975 3935 4980 3940 ne
rect 4980 3935 5048 3940
tri 5048 3935 5054 3941 sw
tri 4980 3883 5032 3935 ne
rect 5032 3883 5054 3935
tri 5054 3883 5106 3935 sw
tri 5032 3877 5038 3883 ne
rect 5038 3877 5106 3883
tri 5106 3877 5112 3883 sw
tri 5038 3868 5047 3877 ne
rect 5047 3868 5112 3877
tri 5112 3868 5121 3877 sw
tri 5047 3802 5113 3868 ne
rect 5113 3802 5121 3868
tri 5121 3802 5187 3868 sw
tri 5113 3794 5121 3802 ne
rect 5121 3794 5187 3802
tri 5187 3794 5195 3802 sw
tri 5121 3769 5146 3794 ne
rect 5146 3769 5195 3794
tri 5195 3769 5220 3794 sw
tri 5146 3764 5151 3769 ne
rect 5151 3764 5220 3769
tri 5220 3764 5225 3769 sw
tri 5151 3720 5195 3764 ne
rect 5195 3720 5225 3764
tri 5225 3720 5269 3764 sw
tri 5195 3712 5203 3720 ne
rect 5203 3712 5269 3720
tri 5269 3712 5277 3720 sw
tri 5203 3704 5211 3712 ne
rect 5211 3704 5277 3712
tri 5277 3704 5285 3712 sw
tri 5211 3700 5215 3704 ne
rect 5215 3700 5285 3704
tri 5285 3700 5289 3704 sw
tri 5215 3648 5267 3700 ne
rect 5267 3648 5289 3700
tri 5289 3648 5341 3700 sw
tri 5267 3646 5269 3648 ne
rect 5269 3646 5341 3648
tri 5341 3646 5343 3648 sw
rect -232 3594 2104 3646
rect 2156 3594 2168 3646
rect 2220 3594 2232 3646
rect 2284 3594 2296 3646
rect 2348 3594 2360 3646
rect 2412 3594 2424 3646
rect 2476 3594 2482 3646
tri 5269 3594 5321 3646 ne
rect 5321 3594 5344 3646
rect 5396 3594 5408 3646
rect 5460 3594 5472 3646
rect 5524 3594 5530 3646
rect 4372 3206 4488 3212
rect 4424 3154 4436 3206
rect -232 2712 2104 2764
rect 2156 2712 2168 2764
rect 2220 2712 2232 2764
rect 2284 2712 2296 2764
rect 2348 2712 2360 2764
rect 2412 2712 2424 2764
rect 2476 2712 2482 2764
rect -232 1786 2104 1838
rect 2156 1786 2168 1838
rect 2220 1786 2232 1838
rect 2284 1786 2296 1838
rect 2348 1786 2360 1838
rect 2412 1786 2424 1838
rect 2476 1786 2482 1838
rect 4372 1390 4488 3154
rect 5862 2331 5978 4017
rect 7730 2773 7846 4660
rect 7782 2721 7794 2773
rect 7730 2715 7846 2721
rect 5862 2209 5978 2215
rect 8146 1847 8262 4660
rect 8198 1795 8210 1847
rect 8146 1789 8262 1795
rect 12403 4547 12842 5168
rect 14217 4992 14223 5044
rect 14275 4992 14290 5044
rect 14342 4992 14348 5044
tri 14217 4985 14224 4992 ne
rect 14224 4985 14341 4992
tri 14341 4985 14348 4992 nw
tri 14224 4984 14225 4985 ne
rect 14225 4973 14329 4985
tri 14329 4973 14341 4985 nw
tri 14194 4676 14225 4707 se
rect 14225 4676 14325 4973
tri 14325 4969 14329 4973 nw
rect 12403 4495 12419 4547
rect 12471 4495 12490 4547
rect 12542 4495 12561 4547
rect 12613 4495 12632 4547
rect 12684 4495 12703 4547
rect 12755 4495 12773 4547
rect 12825 4495 12842 4547
rect 12403 4483 12842 4495
rect 12403 4431 12419 4483
rect 12471 4431 12490 4483
rect 12542 4431 12561 4483
rect 12613 4431 12632 4483
rect 12684 4431 12703 4483
rect 12755 4431 12773 4483
rect 12825 4431 12842 4483
rect 12403 4063 12842 4431
rect 12403 4011 12592 4063
rect 12644 4011 12684 4063
rect 12736 4011 12775 4063
rect 12827 4011 12842 4063
rect 12403 3999 12842 4011
rect 12403 3947 12592 3999
rect 12644 3947 12684 3999
rect 12736 3947 12775 3999
rect 12827 3947 12842 3999
rect 12403 3935 12842 3947
rect 12403 3883 12592 3935
rect 12644 3883 12684 3935
rect 12736 3883 12775 3935
rect 12827 3883 12842 3935
rect 12403 3764 12842 3883
rect 12403 3712 12592 3764
rect 12644 3712 12684 3764
rect 12736 3712 12775 3764
rect 12827 3712 12842 3764
rect 12403 3700 12842 3712
rect 12403 3648 12592 3700
rect 12644 3648 12684 3700
rect 12736 3648 12775 3700
rect 12827 3648 12842 3700
rect 12403 3636 12842 3648
rect 12403 3584 12592 3636
rect 12644 3584 12684 3636
rect 12736 3584 12775 3636
rect 12827 3584 12842 3636
rect 12403 3468 12842 3584
rect 12403 3416 12411 3468
rect 12463 3416 12484 3468
rect 12536 3416 12556 3468
rect 12608 3416 12628 3468
rect 12680 3416 12700 3468
rect 12752 3416 12772 3468
rect 12824 3416 12842 3468
rect 12403 3404 12842 3416
rect 12403 3352 12411 3404
rect 12463 3352 12484 3404
rect 12536 3352 12556 3404
rect 12608 3352 12628 3404
rect 12680 3352 12700 3404
rect 12752 3352 12772 3404
rect 12824 3352 12842 3404
rect 12403 3340 12842 3352
rect 12403 3288 12411 3340
rect 12463 3288 12484 3340
rect 12536 3288 12556 3340
rect 12608 3288 12628 3340
rect 12680 3288 12700 3340
rect 12752 3288 12772 3340
rect 12824 3288 12842 3340
rect 12403 3276 12842 3288
rect 12403 3224 12411 3276
rect 12463 3224 12484 3276
rect 12536 3224 12556 3276
rect 12608 3224 12628 3276
rect 12680 3224 12700 3276
rect 12752 3224 12772 3276
rect 12824 3224 12842 3276
rect 12403 2701 12842 3224
rect 12403 2649 12414 2701
rect 12466 2649 12486 2701
rect 12538 2649 12558 2701
rect 12610 2649 12630 2701
rect 12682 2649 12702 2701
rect 12754 2649 12774 2701
rect 12826 2649 12842 2701
rect 12403 2637 12842 2649
rect 12403 2585 12414 2637
rect 12466 2585 12486 2637
rect 12538 2585 12558 2637
rect 12610 2585 12630 2637
rect 12682 2585 12702 2637
rect 12754 2585 12774 2637
rect 12826 2585 12842 2637
rect 13292 4624 13322 4676
rect 13374 4624 13389 4676
rect 13441 4624 13447 4676
rect 14194 4624 14200 4676
rect 14252 4624 14267 4676
rect 14319 4624 14325 4676
rect 13292 2792 13392 4624
tri 13392 4589 13427 4624 nw
rect 14334 4269 14340 4385
rect 14456 4269 14462 4385
tri 13392 2792 13408 2808 sw
rect 13292 2786 13408 2792
rect 13344 2734 13356 2786
rect 13292 2719 13408 2734
rect 13344 2667 13356 2719
rect 13292 2648 13408 2667
rect 13292 2605 13408 2646
rect 12403 2573 12842 2585
rect 12403 2521 12414 2573
rect 12466 2521 12486 2573
rect 12538 2521 12558 2573
rect 12610 2521 12630 2573
rect 12682 2521 12702 2573
rect 12754 2521 12774 2573
rect 12826 2521 12842 2573
tri 13294 2558 13300 2564 se
rect 13300 2558 13399 2564
rect 12403 2143 12842 2521
tri 13242 2506 13294 2558 se
rect 13294 2506 13399 2558
tri 13235 2499 13242 2506 se
rect 13242 2499 13399 2506
rect 13235 2433 13399 2499
rect 13401 2558 13532 2564
rect 13401 2506 13416 2558
rect 13468 2506 13480 2558
rect 13401 2491 13532 2506
rect 13401 2439 13416 2491
rect 13468 2439 13480 2491
rect 13401 2433 13532 2439
rect 13235 2390 13351 2433
tri 13351 2396 13388 2433 nw
rect 13287 2338 13299 2390
rect 13235 2323 13351 2338
rect 13287 2271 13299 2323
rect 13235 2265 13351 2271
rect 12403 2091 12412 2143
rect 12464 2091 12486 2143
rect 12538 2091 12560 2143
rect 12612 2091 12634 2143
rect 12686 2091 12707 2143
rect 12759 2091 12780 2143
rect 12832 2091 12842 2143
rect 13561 2098 13753 2956
rect 14334 2877 14462 4269
rect 14334 2761 14340 2877
rect 14456 2761 14462 2877
rect 15699 4057 16439 6995
tri 16439 6970 16464 6995 nw
rect 17481 5375 17487 5427
rect 17539 5375 17551 5427
rect 17603 5375 17609 5427
rect 16551 5248 16603 5251
tri 16603 5248 16606 5251 sw
rect 16551 5245 16606 5248
rect 16603 5242 16606 5245
tri 16606 5242 16612 5248 sw
tri 16868 5242 16874 5248 se
rect 16874 5242 16926 5248
rect 16603 5220 16612 5242
tri 16612 5220 16634 5242 sw
tri 16846 5220 16868 5242 se
rect 16868 5220 16874 5242
rect 16603 5193 16874 5220
rect 16551 5190 16874 5193
rect 16551 5178 16926 5190
rect 16603 5126 16874 5178
rect 16551 5120 16926 5126
rect 16520 5037 17054 5045
rect 16520 4985 16932 5037
rect 16984 4985 16996 5037
rect 17048 4985 17054 5037
rect 16520 4973 16604 4985
tri 16604 4973 16616 4985 nw
tri 16495 4210 16520 4235 se
rect 16520 4210 16576 4973
tri 16576 4945 16604 4973 nw
rect 16892 4719 17020 4746
tri 16576 4210 16623 4257 sw
rect 16892 4210 16898 4262
rect 16950 4210 16962 4262
rect 17014 4210 17020 4262
rect 16947 4206 16968 4210
tri 16968 4206 16972 4210 nw
tri 16947 4185 16968 4206 nw
rect 15699 4005 15705 4057
rect 15757 4005 16439 4057
rect 15699 3993 16439 4005
rect 15699 3941 15705 3993
rect 15757 3941 16439 3993
rect 15699 3929 16439 3941
rect 15699 3877 15705 3929
rect 15757 3877 16439 3929
rect 15699 3769 16439 3877
rect 15699 3717 15723 3769
rect 15775 3717 15787 3769
rect 15839 3717 15851 3769
rect 15903 3717 15915 3769
rect 15967 3717 15979 3769
rect 16031 3717 16043 3769
rect 16095 3717 16107 3769
rect 16159 3717 16171 3769
rect 16223 3717 16235 3769
rect 16287 3717 16299 3769
rect 16351 3717 16363 3769
rect 16415 3717 16439 3769
rect 15699 3704 16439 3717
rect 15699 3652 15723 3704
rect 15775 3652 15787 3704
rect 15839 3652 15851 3704
rect 15903 3652 15915 3704
rect 15967 3652 15979 3704
rect 16031 3652 16043 3704
rect 16095 3652 16107 3704
rect 16159 3652 16171 3704
rect 16223 3652 16235 3704
rect 16287 3652 16299 3704
rect 16351 3652 16363 3704
rect 16415 3652 16439 3704
rect 15699 3639 16439 3652
rect 15699 3587 15723 3639
rect 15775 3587 15787 3639
rect 15839 3587 15851 3639
rect 15903 3587 15915 3639
rect 15967 3587 15979 3639
rect 16031 3587 16043 3639
rect 16095 3587 16107 3639
rect 16159 3587 16171 3639
rect 16223 3587 16235 3639
rect 16287 3587 16299 3639
rect 16351 3587 16363 3639
rect 16415 3587 16439 3639
rect 15699 3475 16439 3587
rect 15699 3423 15723 3475
rect 15775 3423 15787 3475
rect 15839 3423 15851 3475
rect 15903 3423 15915 3475
rect 15967 3423 15979 3475
rect 16031 3423 16043 3475
rect 16095 3423 16107 3475
rect 16159 3423 16171 3475
rect 16223 3423 16235 3475
rect 16287 3423 16299 3475
rect 16351 3423 16363 3475
rect 16415 3423 16439 3475
rect 15699 3406 16439 3423
rect 15699 3354 15723 3406
rect 15775 3354 15787 3406
rect 15839 3354 15851 3406
rect 15903 3354 15915 3406
rect 15967 3354 15979 3406
rect 16031 3354 16043 3406
rect 16095 3354 16107 3406
rect 16159 3354 16171 3406
rect 16223 3354 16235 3406
rect 16287 3354 16299 3406
rect 16351 3354 16363 3406
rect 16415 3354 16439 3406
rect 15699 3337 16439 3354
rect 15699 3285 15723 3337
rect 15775 3285 15787 3337
rect 15839 3285 15851 3337
rect 15903 3285 15915 3337
rect 15967 3285 15979 3337
rect 16031 3285 16043 3337
rect 16095 3285 16107 3337
rect 16159 3285 16171 3337
rect 16223 3285 16235 3337
rect 16287 3285 16299 3337
rect 16351 3285 16363 3337
rect 16415 3285 16439 3337
rect 15699 3268 16439 3285
rect 15699 3216 15723 3268
rect 15775 3216 15787 3268
rect 15839 3216 15851 3268
rect 15903 3216 15915 3268
rect 15967 3216 15979 3268
rect 16031 3216 16043 3268
rect 16095 3216 16107 3268
rect 16159 3216 16171 3268
rect 16223 3216 16235 3268
rect 16287 3216 16299 3268
rect 16351 3216 16363 3268
rect 16415 3216 16439 3268
rect 15699 2255 16439 3216
rect 17481 4145 17609 5375
tri 20208 5130 20256 5178 se
rect 20256 5130 20336 10183
tri 20336 10149 20370 10183 nw
tri 25107 10168 25122 10183 ne
rect 25122 10168 25204 10183
tri 25204 10168 25219 10183 sw
tri 25122 10166 25124 10168 ne
rect 25124 10166 25219 10168
tri 25124 10149 25141 10166 ne
rect 25141 10149 25219 10166
tri 25219 10149 25238 10168 sw
tri 25141 10127 25163 10149 ne
rect 25163 10127 25238 10149
tri 25238 10127 25260 10149 sw
rect 20392 10124 25090 10127
tri 25090 10124 25093 10127 sw
tri 25163 10124 25166 10127 ne
rect 25166 10124 25260 10127
tri 25260 10124 25263 10127 sw
rect 20392 10123 25093 10124
rect 20392 10071 24195 10123
rect 24247 10071 24259 10123
rect 24311 10093 25093 10123
tri 25093 10093 25124 10124 sw
tri 25166 10093 25197 10124 ne
rect 25197 10093 25263 10124
rect 24311 10072 25124 10093
tri 25124 10072 25145 10093 sw
tri 25197 10072 25218 10093 ne
rect 25218 10072 25263 10093
tri 25263 10072 25315 10124 sw
rect 25402 10072 25408 10124
rect 25460 10072 25472 10124
rect 25524 10072 25530 10124
rect 24311 10071 25145 10072
tri 25145 10071 25146 10072 sw
tri 25218 10071 25219 10072 ne
rect 25219 10071 25315 10072
tri 25315 10071 25316 10072 sw
rect 20392 10067 25146 10071
tri 25146 10067 25150 10071 sw
tri 25219 10067 25223 10071 ne
rect 25223 10067 25316 10071
tri 25316 10067 25320 10071 sw
tri 20377 5292 20392 5307 se
rect 20392 5292 20452 10067
tri 20452 10033 20486 10067 nw
tri 25063 10051 25079 10067 ne
rect 25079 10059 25150 10067
tri 25150 10059 25158 10067 sw
tri 25223 10059 25231 10067 ne
rect 25231 10059 25320 10067
tri 25320 10059 25328 10067 sw
rect 25079 10051 25158 10059
tri 25158 10051 25166 10059 sw
tri 25231 10051 25239 10059 ne
rect 25239 10051 25328 10059
tri 25328 10051 25336 10059 sw
tri 25079 10040 25090 10051 ne
rect 25090 10050 25166 10051
tri 25166 10050 25167 10051 sw
tri 25239 10050 25240 10051 ne
rect 25240 10050 25336 10051
tri 25336 10050 25337 10051 sw
rect 25090 10040 25167 10050
tri 25090 10033 25097 10040 ne
rect 25097 10033 25167 10040
tri 25167 10033 25184 10050 sw
tri 25240 10033 25257 10050 ne
rect 25257 10033 25337 10050
tri 25337 10033 25354 10050 sw
tri 25097 10011 25119 10033 ne
rect 25119 10011 25184 10033
tri 25184 10011 25206 10033 sw
tri 25257 10011 25279 10033 ne
rect 25279 10011 25354 10033
tri 25354 10011 25376 10033 sw
rect 20508 9992 25071 10011
tri 25071 9992 25090 10011 sw
tri 25119 9992 25138 10011 ne
rect 25138 9998 25206 10011
tri 25206 9998 25219 10011 sw
tri 25279 9998 25292 10011 ne
rect 25292 9998 25376 10011
rect 25138 9992 25219 9998
rect 20508 9974 25090 9992
tri 25090 9974 25108 9992 sw
tri 25138 9974 25156 9992 ne
rect 25156 9985 25219 9992
tri 25219 9985 25232 9998 sw
tri 25292 9985 25305 9998 ne
rect 25305 9985 25376 9998
tri 25376 9985 25402 10011 sw
rect 25156 9974 25232 9985
tri 25232 9974 25243 9985 sw
tri 25305 9974 25316 9985 ne
rect 25316 9974 25402 9985
tri 25402 9974 25413 9985 sw
rect 20508 9964 25108 9974
tri 25108 9964 25118 9974 sw
tri 25156 9964 25166 9974 ne
rect 25166 9964 25243 9974
tri 25243 9964 25253 9974 sw
tri 25316 9964 25326 9974 ne
rect 25326 9964 25511 9974
rect 20508 9953 25118 9964
tri 25118 9953 25129 9964 sw
tri 25166 9953 25177 9964 ne
rect 25177 9953 25253 9964
tri 25253 9953 25264 9964 sw
tri 25326 9953 25337 9964 ne
rect 25337 9953 25511 9964
rect 20508 9931 25129 9953
tri 25129 9931 25151 9953 sw
tri 25177 9931 25199 9953 ne
rect 25199 9931 25264 9953
tri 25264 9931 25286 9953 sw
tri 25337 9931 25359 9953 ne
rect 25359 9931 25511 9953
rect 20508 9922 20613 9931
tri 20613 9922 20622 9931 nw
tri 25038 9922 25047 9931 ne
rect 25047 9922 25151 9931
tri 25151 9922 25160 9931 sw
tri 25199 9922 25208 9931 ne
rect 25208 9922 25286 9931
tri 25286 9922 25295 9931 sw
tri 25359 9922 25368 9931 ne
rect 25368 9922 25511 9931
rect 25563 9922 25575 9974
rect 25627 9922 25633 9974
tri 20503 8575 20508 8580 se
rect 20508 8575 20588 9922
tri 20588 9897 20613 9922 nw
tri 25047 9897 25072 9922 ne
rect 25072 9916 25160 9922
tri 25160 9916 25166 9922 sw
tri 25208 9916 25214 9922 ne
rect 25214 9916 25295 9922
rect 25072 9897 25166 9916
tri 25166 9897 25185 9916 sw
tri 25214 9897 25233 9916 ne
rect 25233 9897 25295 9916
tri 25295 9897 25320 9922 sw
tri 25072 9875 25094 9897 ne
rect 25094 9887 25185 9897
tri 25185 9887 25195 9897 sw
tri 25233 9887 25243 9897 ne
rect 25243 9887 25320 9897
tri 25320 9887 25330 9897 sw
rect 25094 9877 25195 9887
tri 25195 9877 25205 9887 sw
tri 25243 9877 25253 9887 ne
rect 25253 9877 25330 9887
tri 25330 9877 25340 9887 sw
rect 25094 9875 25205 9877
tri 25205 9875 25207 9877 sw
tri 25253 9875 25255 9877 ne
rect 25255 9875 25611 9877
tri 25611 9875 25613 9877 sw
rect 20696 9823 20702 9875
rect 20754 9823 20768 9875
rect 20820 9823 20834 9875
rect 20886 9823 20900 9875
rect 20952 9823 20966 9875
rect 21018 9823 21032 9875
rect 21084 9823 21097 9875
rect 21149 9823 21162 9875
rect 21214 9823 21227 9875
rect 21279 9823 21292 9875
rect 21344 9823 21357 9875
rect 21409 9823 21415 9875
tri 25094 9840 25129 9875 ne
rect 25129 9840 25207 9875
tri 25207 9840 25242 9875 sw
tri 25255 9840 25290 9875 ne
rect 25290 9840 25613 9875
tri 25613 9840 25648 9875 sw
rect 25757 9840 25818 10196
rect 28063 10072 28069 10124
rect 28121 10072 28133 10124
rect 28185 10072 28816 10124
tri 28816 10072 28868 10124 sw
tri 28794 10067 28799 10072 ne
rect 28799 10067 28868 10072
tri 28868 10067 28873 10072 sw
tri 28799 10059 28807 10067 ne
rect 28807 10059 28873 10067
tri 28873 10059 28881 10067 sw
tri 28807 10050 28816 10059 ne
rect 28816 10050 28881 10059
tri 28816 10033 28833 10050 ne
rect 28833 10033 28881 10050
tri 28881 10033 28907 10059 sw
tri 28833 10011 28855 10033 ne
rect 28855 10011 28907 10033
tri 28907 10011 28929 10033 sw
tri 28855 9985 28881 10011 ne
rect 28881 9985 28929 10011
tri 28929 9985 28955 10011 sw
tri 28881 9974 28892 9985 ne
rect 28892 9974 28955 9985
rect 27658 9922 27664 9974
rect 27716 9922 27728 9974
rect 27780 9922 27786 9974
tri 28892 9963 28903 9974 ne
tri 27658 9887 27693 9922 ne
rect 27693 9887 27751 9922
tri 27751 9887 27786 9922 nw
tri 25818 9840 25827 9849 sw
rect 20696 9811 21415 9823
rect 20696 9759 20702 9811
rect 20754 9759 20768 9811
rect 20820 9759 20834 9811
rect 20886 9759 20900 9811
rect 20952 9759 20966 9811
rect 21018 9759 21032 9811
rect 21084 9759 21097 9811
rect 21149 9759 21162 9811
rect 21214 9759 21227 9811
rect 21279 9759 21292 9811
rect 21344 9759 21357 9811
rect 21409 9759 21415 9811
tri 25129 9780 25189 9840 ne
rect 25189 9832 25242 9840
tri 25242 9832 25250 9840 sw
tri 25290 9832 25298 9840 ne
rect 25298 9832 25648 9840
rect 25189 9780 25250 9832
tri 25250 9780 25302 9832 sw
tri 25581 9822 25591 9832 ne
rect 25591 9822 25648 9832
tri 25648 9822 25666 9840 sw
tri 25591 9802 25611 9822 ne
rect 25611 9802 25666 9822
tri 25611 9799 25614 9802 ne
tri 25189 9779 25190 9780 ne
rect 25190 9779 25302 9780
tri 25302 9779 25303 9780 sw
rect 20696 9005 21415 9759
tri 25190 9728 25241 9779 ne
rect 25241 9727 25247 9779
rect 25299 9727 25311 9779
rect 25363 9727 25369 9779
rect 25614 9526 25666 9802
rect 25757 9826 25827 9840
tri 25757 9796 25787 9826 ne
rect 25787 9796 25827 9826
tri 25827 9796 25871 9840 sw
tri 25787 9780 25803 9796 ne
rect 25803 9780 25871 9796
tri 25871 9780 25887 9796 sw
tri 25803 9765 25818 9780 ne
rect 25818 9765 25887 9780
tri 25818 9728 25855 9765 ne
rect 25855 9728 25887 9765
tri 25887 9728 25939 9780 sw
rect 27306 9728 27312 9780
rect 27364 9728 27376 9780
rect 27428 9728 27434 9780
tri 25855 9712 25871 9728 ne
rect 25871 9727 25939 9728
tri 25939 9727 25940 9728 sw
tri 27306 9727 27307 9728 ne
rect 27307 9727 27399 9728
rect 25871 9712 25940 9727
tri 25940 9712 25955 9727 sw
tri 27307 9712 27322 9727 ne
rect 27322 9712 27399 9727
tri 25871 9628 25955 9712 ne
tri 25955 9693 25974 9712 sw
tri 27322 9693 27341 9712 ne
rect 27341 9693 27399 9712
tri 27399 9693 27434 9728 nw
rect 25955 9628 25974 9693
tri 25974 9628 26039 9693 sw
tri 25955 9546 26037 9628 ne
rect 26037 9546 26039 9628
tri 26039 9546 26121 9628 sw
rect 27341 9546 27396 9693
tri 27396 9690 27399 9693 nw
tri 26037 9544 26039 9546 ne
rect 26039 9544 26121 9546
tri 26121 9544 26123 9546 sw
tri 26039 9526 26057 9544 ne
rect 26057 9526 26123 9544
tri 26057 9520 26063 9526 ne
rect 26063 9385 26123 9526
rect 27341 9494 27342 9546
rect 27394 9494 27396 9546
rect 27341 9491 27396 9494
rect 27341 9482 27395 9491
rect 27693 9490 27745 9887
tri 27745 9881 27751 9887 nw
tri 26123 9437 26157 9471 sw
rect 27341 9430 27342 9482
rect 27394 9430 27395 9482
rect 27341 9424 27395 9430
rect 27916 9424 27922 9476
rect 27974 9424 27986 9476
rect 28038 9450 28689 9476
tri 28689 9450 28715 9476 sw
rect 28038 9424 28715 9450
tri 28715 9424 28741 9450 sw
tri 28667 9385 28706 9424 ne
rect 28706 9385 28741 9424
tri 28706 9376 28715 9385 ne
rect 28715 9376 28741 9385
tri 28741 9376 28789 9424 sw
tri 28715 9302 28789 9376 ne
tri 28789 9302 28863 9376 sw
tri 28789 9280 28811 9302 ne
rect 20696 8953 20702 9005
rect 20754 8953 20768 9005
rect 20820 8953 20834 9005
rect 20886 8953 20900 9005
rect 20952 8953 20966 9005
rect 21018 8953 21032 9005
rect 21084 8953 21097 9005
rect 21149 8953 21162 9005
rect 21214 8953 21227 9005
rect 21279 8953 21292 9005
rect 21344 8953 21357 9005
rect 21409 8953 21415 9005
rect 20696 8941 21415 8953
rect 20696 8889 20702 8941
rect 20754 8889 20768 8941
rect 20820 8889 20834 8941
rect 20886 8889 20900 8941
rect 20952 8889 20966 8941
rect 21018 8889 21032 8941
rect 21084 8889 21097 8941
rect 21149 8889 21162 8941
rect 21214 8889 21227 8941
rect 21279 8889 21292 8941
rect 21344 8889 21357 8941
rect 21409 8889 21415 8941
rect 20696 8877 21415 8889
rect 20696 8825 20702 8877
rect 20754 8825 20768 8877
rect 20820 8825 20834 8877
rect 20886 8825 20900 8877
rect 20952 8825 20966 8877
rect 21018 8825 21032 8877
rect 21084 8825 21097 8877
rect 21149 8825 21162 8877
rect 21214 8825 21227 8877
rect 21279 8825 21292 8877
rect 21344 8825 21357 8877
rect 21409 8825 21415 8877
rect 20696 8813 21415 8825
rect 20696 8761 20702 8813
rect 20754 8761 20768 8813
rect 20820 8761 20834 8813
rect 20886 8761 20900 8813
rect 20952 8761 20966 8813
rect 21018 8761 21032 8813
rect 21084 8761 21097 8813
rect 21149 8761 21162 8813
rect 21214 8761 21227 8813
rect 21279 8761 21292 8813
rect 21344 8761 21357 8813
rect 21409 8761 21415 8813
rect 20696 8749 21415 8761
rect 20696 8697 20702 8749
rect 20754 8697 20768 8749
rect 20820 8697 20834 8749
rect 20886 8697 20900 8749
rect 20952 8697 20966 8749
rect 21018 8697 21032 8749
rect 21084 8697 21097 8749
rect 21149 8697 21162 8749
rect 21214 8697 21227 8749
rect 21279 8697 21292 8749
rect 21344 8697 21357 8749
rect 21409 8697 21415 8749
rect 20696 8685 21415 8697
rect 20696 8633 20702 8685
rect 20754 8633 20768 8685
rect 20820 8633 20834 8685
rect 20886 8633 20900 8685
rect 20952 8633 20966 8685
rect 21018 8633 21032 8685
rect 21084 8633 21097 8685
rect 21149 8633 21162 8685
rect 21214 8633 21227 8685
rect 21279 8633 21292 8685
rect 21344 8633 21357 8685
rect 21409 8633 21415 8685
tri 20588 8575 20631 8618 sw
rect 20503 8523 20509 8575
rect 20561 8523 20573 8575
rect 20625 8523 20631 8575
tri 20503 8518 20508 8523 ne
rect 20508 8495 20603 8523
tri 20603 8495 20631 8523 nw
rect 20696 8495 21415 8633
rect 20508 5427 20588 8495
tri 20588 8480 20603 8495 nw
rect 20696 8443 20702 8495
rect 20754 8443 20768 8495
rect 20820 8443 20834 8495
rect 20886 8443 20900 8495
rect 20952 8443 20966 8495
rect 21018 8443 21032 8495
rect 21084 8443 21097 8495
rect 21149 8443 21162 8495
rect 21214 8443 21227 8495
rect 21279 8443 21292 8495
rect 21344 8443 21357 8495
rect 21409 8443 21415 8495
rect 20696 8431 21415 8443
rect 20696 8379 20702 8431
rect 20754 8379 20768 8431
rect 20820 8379 20834 8431
rect 20886 8379 20900 8431
rect 20952 8379 20966 8431
rect 21018 8379 21032 8431
rect 21084 8379 21097 8431
rect 21149 8379 21162 8431
rect 21214 8379 21227 8431
rect 21279 8379 21292 8431
rect 21344 8379 21357 8431
rect 21409 8379 21415 8431
rect 20696 8367 21415 8379
rect 20696 8315 20702 8367
rect 20754 8315 20768 8367
rect 20820 8315 20834 8367
rect 20886 8315 20900 8367
rect 20952 8315 20966 8367
rect 21018 8315 21032 8367
rect 21084 8315 21097 8367
rect 21149 8315 21162 8367
rect 21214 8315 21227 8367
rect 21279 8315 21292 8367
rect 21344 8315 21357 8367
rect 21409 8315 21415 8367
rect 20696 8231 21415 8315
rect 20696 8179 20702 8231
rect 20754 8179 20768 8231
rect 20820 8179 20834 8231
rect 20886 8179 20900 8231
rect 20952 8179 20966 8231
rect 21018 8179 21032 8231
rect 21084 8179 21097 8231
rect 21149 8179 21162 8231
rect 21214 8179 21227 8231
rect 21279 8179 21292 8231
rect 21344 8179 21357 8231
rect 21409 8179 21415 8231
rect 20696 8167 21415 8179
rect 20696 8115 20702 8167
rect 20754 8115 20768 8167
rect 20820 8115 20834 8167
rect 20886 8115 20900 8167
rect 20952 8115 20966 8167
rect 21018 8115 21032 8167
rect 21084 8115 21097 8167
rect 21149 8115 21162 8167
rect 21214 8115 21227 8167
rect 21279 8115 21292 8167
rect 21344 8115 21357 8167
rect 21409 8115 21415 8167
rect 20696 8103 21415 8115
rect 20696 8051 20702 8103
rect 20754 8051 20768 8103
rect 20820 8051 20834 8103
rect 20886 8051 20900 8103
rect 20952 8051 20966 8103
rect 21018 8051 21032 8103
rect 21084 8051 21097 8103
rect 21149 8051 21162 8103
rect 21214 8051 21227 8103
rect 21279 8051 21292 8103
rect 21344 8051 21357 8103
rect 21409 8051 21415 8103
rect 20696 7967 21415 8051
rect 20696 7915 20702 7967
rect 20754 7915 20768 7967
rect 20820 7915 20834 7967
rect 20886 7915 20900 7967
rect 20952 7915 20966 7967
rect 21018 7915 21032 7967
rect 21084 7915 21097 7967
rect 21149 7915 21162 7967
rect 21214 7915 21227 7967
rect 21279 7915 21292 7967
rect 21344 7915 21357 7967
rect 21409 7915 21415 7967
rect 20696 7903 21415 7915
rect 20696 7851 20702 7903
rect 20754 7851 20768 7903
rect 20820 7851 20834 7903
rect 20886 7851 20900 7903
rect 20952 7851 20966 7903
rect 21018 7851 21032 7903
rect 21084 7851 21097 7903
rect 21149 7851 21162 7903
rect 21214 7851 21227 7903
rect 21279 7851 21292 7903
rect 21344 7851 21357 7903
rect 21409 7851 21415 7903
rect 20696 7839 21415 7851
rect 20696 7787 20702 7839
rect 20754 7787 20768 7839
rect 20820 7787 20834 7839
rect 20886 7787 20900 7839
rect 20952 7787 20966 7839
rect 21018 7787 21032 7839
rect 21084 7787 21097 7839
rect 21149 7787 21162 7839
rect 21214 7787 21227 7839
rect 21279 7787 21292 7839
rect 21344 7787 21357 7839
rect 21409 7787 21415 7839
rect 20696 7703 21415 7787
rect 20696 7651 20702 7703
rect 20754 7651 20768 7703
rect 20820 7651 20834 7703
rect 20886 7651 20900 7703
rect 20952 7651 20966 7703
rect 21018 7651 21032 7703
rect 21084 7651 21097 7703
rect 21149 7651 21162 7703
rect 21214 7651 21227 7703
rect 21279 7651 21292 7703
rect 21344 7651 21357 7703
rect 21409 7651 21415 7703
rect 20696 7639 21415 7651
rect 20696 7587 20702 7639
rect 20754 7587 20768 7639
rect 20820 7587 20834 7639
rect 20886 7587 20900 7639
rect 20952 7587 20966 7639
rect 21018 7587 21032 7639
rect 21084 7587 21097 7639
rect 21149 7587 21162 7639
rect 21214 7587 21227 7639
rect 21279 7587 21292 7639
rect 21344 7587 21357 7639
rect 21409 7587 21415 7639
rect 20696 7575 21415 7587
rect 20696 7523 20702 7575
rect 20754 7523 20768 7575
rect 20820 7523 20834 7575
rect 20886 7523 20900 7575
rect 20952 7523 20966 7575
rect 21018 7523 21032 7575
rect 21084 7523 21097 7575
rect 21149 7523 21162 7575
rect 21214 7523 21227 7575
rect 21279 7523 21292 7575
rect 21344 7523 21357 7575
rect 21409 7523 21415 7575
rect 20696 7439 21415 7523
rect 20696 7387 20702 7439
rect 20754 7387 20768 7439
rect 20820 7387 20834 7439
rect 20886 7387 20900 7439
rect 20952 7387 20966 7439
rect 21018 7387 21032 7439
rect 21084 7387 21097 7439
rect 21149 7387 21162 7439
rect 21214 7387 21227 7439
rect 21279 7387 21292 7439
rect 21344 7387 21357 7439
rect 21409 7387 21415 7439
rect 20696 7375 21415 7387
rect 20696 7323 20702 7375
rect 20754 7323 20768 7375
rect 20820 7323 20834 7375
rect 20886 7323 20900 7375
rect 20952 7323 20966 7375
rect 21018 7323 21032 7375
rect 21084 7323 21097 7375
rect 21149 7323 21162 7375
rect 21214 7323 21227 7375
rect 21279 7323 21292 7375
rect 21344 7323 21357 7375
rect 21409 7323 21415 7375
rect 20696 7311 21415 7323
rect 20696 7259 20702 7311
rect 20754 7259 20768 7311
rect 20820 7259 20834 7311
rect 20886 7259 20900 7311
rect 20952 7259 20966 7311
rect 21018 7259 21032 7311
rect 21084 7259 21097 7311
rect 21149 7259 21162 7311
rect 21214 7259 21227 7311
rect 21279 7259 21292 7311
rect 21344 7259 21357 7311
rect 21409 7259 21415 7311
rect 20696 7175 21415 7259
rect 20696 7123 20702 7175
rect 20754 7123 20768 7175
rect 20820 7123 20834 7175
rect 20886 7123 20900 7175
rect 20952 7123 20966 7175
rect 21018 7123 21032 7175
rect 21084 7123 21097 7175
rect 21149 7123 21162 7175
rect 21214 7123 21227 7175
rect 21279 7123 21292 7175
rect 21344 7123 21357 7175
rect 21409 7123 21415 7175
rect 20696 7111 21415 7123
rect 20696 7059 20702 7111
rect 20754 7059 20768 7111
rect 20820 7059 20834 7111
rect 20886 7059 20900 7111
rect 20952 7059 20966 7111
rect 21018 7059 21032 7111
rect 21084 7059 21097 7111
rect 21149 7059 21162 7111
rect 21214 7059 21227 7111
rect 21279 7059 21292 7111
rect 21344 7059 21357 7111
rect 21409 7059 21415 7111
rect 20696 7047 21415 7059
rect 20696 6995 20702 7047
rect 20754 6995 20768 7047
rect 20820 6995 20834 7047
rect 20886 6995 20900 7047
rect 20952 6995 20966 7047
rect 21018 6995 21032 7047
rect 21084 6995 21097 7047
rect 21149 6995 21162 7047
rect 21214 6995 21227 7047
rect 21279 6995 21292 7047
rect 21344 6995 21357 7047
rect 21409 6995 21415 7047
rect 23932 9126 24514 9132
rect 23932 7218 23941 9126
rect 24505 7218 24514 9126
rect 23932 7205 24514 7218
rect 23932 7153 23941 7205
rect 23993 7153 24005 7205
rect 24057 7153 24069 7205
rect 24121 7153 24133 7205
rect 24185 7153 24197 7205
rect 24249 7153 24261 7205
rect 24313 7153 24325 7205
rect 24377 7153 24389 7205
rect 24441 7153 24453 7205
rect 24505 7153 24514 7205
rect 23932 7140 24514 7153
rect 23932 7088 23941 7140
rect 23993 7088 24005 7140
rect 24057 7088 24069 7140
rect 24121 7088 24133 7140
rect 24185 7088 24197 7140
rect 24249 7088 24261 7140
rect 24313 7088 24325 7140
rect 24377 7088 24389 7140
rect 24441 7088 24453 7140
rect 24505 7088 24514 7140
rect 23932 7075 24514 7088
rect 23932 7023 23941 7075
rect 23993 7023 24005 7075
rect 24057 7023 24069 7075
rect 24121 7023 24133 7075
rect 24185 7023 24197 7075
rect 24249 7023 24261 7075
rect 24313 7023 24325 7075
rect 24377 7023 24389 7075
rect 24441 7023 24453 7075
rect 24505 7023 24514 7075
rect 23932 7010 24514 7023
rect 23932 6958 23941 7010
rect 23993 6958 24005 7010
rect 24057 6958 24069 7010
rect 24121 6958 24133 7010
rect 24185 6958 24197 7010
rect 24249 6958 24261 7010
rect 24313 6958 24325 7010
rect 24377 6958 24389 7010
rect 24441 6958 24453 7010
rect 24505 6958 24514 7010
rect 23932 6945 24514 6958
tri 25293 6948 25345 7000 se
rect 25345 6948 25528 7000
rect 25580 6948 25592 7000
rect 25644 6948 25650 7000
rect 28177 6948 28183 7000
rect 28235 6948 28271 7000
rect 28323 6997 28692 7000
tri 28692 6997 28695 7000 sw
rect 28323 6948 28695 6997
tri 28695 6948 28744 6997 sw
rect 23932 6893 23941 6945
rect 23993 6893 24005 6945
rect 24057 6893 24069 6945
rect 24121 6893 24133 6945
rect 24185 6893 24197 6945
rect 24249 6893 24261 6945
rect 24313 6893 24325 6945
rect 24377 6893 24389 6945
rect 24441 6893 24453 6945
rect 24505 6893 24514 6945
rect 23932 6880 24514 6893
rect 23932 6828 23941 6880
rect 23993 6828 24005 6880
rect 24057 6828 24069 6880
rect 24121 6828 24133 6880
rect 24185 6828 24197 6880
rect 24249 6828 24261 6880
rect 24313 6828 24325 6880
rect 24377 6828 24389 6880
rect 24441 6828 24453 6880
rect 24505 6828 24514 6880
rect 23932 6815 24514 6828
rect 23932 6763 23941 6815
rect 23993 6763 24005 6815
rect 24057 6763 24069 6815
rect 24121 6763 24133 6815
rect 24185 6763 24197 6815
rect 24249 6763 24261 6815
rect 24313 6763 24325 6815
rect 24377 6763 24389 6815
rect 24441 6763 24453 6815
rect 24505 6763 24514 6815
rect 23932 6750 24514 6763
rect 23932 6698 23941 6750
rect 23993 6698 24005 6750
rect 24057 6698 24069 6750
rect 24121 6698 24133 6750
rect 24185 6698 24197 6750
rect 24249 6698 24261 6750
rect 24313 6698 24325 6750
rect 24377 6698 24389 6750
rect 24441 6698 24453 6750
rect 24505 6698 24514 6750
rect 23932 6685 24514 6698
rect 23932 6633 23941 6685
rect 23993 6633 24005 6685
rect 24057 6633 24069 6685
rect 24121 6633 24133 6685
rect 24185 6633 24197 6685
rect 24249 6633 24261 6685
rect 24313 6633 24325 6685
rect 24377 6633 24389 6685
rect 24441 6633 24453 6685
rect 24505 6633 24514 6685
rect 23932 6620 24514 6633
rect 23932 6568 23941 6620
rect 23993 6568 24005 6620
rect 24057 6568 24069 6620
rect 24121 6568 24133 6620
rect 24185 6568 24197 6620
rect 24249 6568 24261 6620
rect 24313 6568 24325 6620
rect 24377 6568 24389 6620
rect 24441 6568 24453 6620
rect 24505 6568 24514 6620
rect 23932 6555 24514 6568
rect 23932 6503 23941 6555
rect 23993 6503 24005 6555
rect 24057 6503 24069 6555
rect 24121 6503 24133 6555
rect 24185 6503 24197 6555
rect 24249 6503 24261 6555
rect 24313 6503 24325 6555
rect 24377 6503 24389 6555
rect 24441 6503 24453 6555
rect 24505 6503 24514 6555
rect 23932 6490 24514 6503
rect 23932 6438 23941 6490
rect 23993 6438 24005 6490
rect 24057 6438 24069 6490
rect 24121 6438 24133 6490
rect 24185 6438 24197 6490
rect 24249 6438 24261 6490
rect 24313 6438 24325 6490
rect 24377 6438 24389 6490
rect 24441 6438 24453 6490
rect 24505 6438 24514 6490
rect 23932 6425 24514 6438
rect 23932 6373 23941 6425
rect 23993 6373 24005 6425
rect 24057 6373 24069 6425
rect 24121 6373 24133 6425
rect 24185 6373 24197 6425
rect 24249 6373 24261 6425
rect 24313 6373 24325 6425
rect 24377 6373 24389 6425
rect 24441 6373 24453 6425
rect 24505 6373 24514 6425
rect 23932 6360 24514 6373
rect 23932 6308 23941 6360
rect 23993 6308 24005 6360
rect 24057 6308 24069 6360
rect 24121 6308 24133 6360
rect 24185 6308 24197 6360
rect 24249 6308 24261 6360
rect 24313 6308 24325 6360
rect 24377 6308 24389 6360
rect 24441 6308 24453 6360
rect 24505 6308 24514 6360
rect 23932 6295 24514 6308
rect 23932 6243 23941 6295
rect 23993 6243 24005 6295
rect 24057 6243 24069 6295
rect 24121 6243 24133 6295
rect 24185 6243 24197 6295
rect 24249 6243 24261 6295
rect 24313 6243 24325 6295
rect 24377 6243 24389 6295
rect 24441 6243 24453 6295
rect 24505 6243 24514 6295
rect 23932 6230 24514 6243
rect 23932 6178 23941 6230
rect 23993 6178 24005 6230
rect 24057 6178 24069 6230
rect 24121 6178 24133 6230
rect 24185 6178 24197 6230
rect 24249 6178 24261 6230
rect 24313 6178 24325 6230
rect 24377 6178 24389 6230
rect 24441 6178 24453 6230
rect 24505 6178 24514 6230
rect 23932 6165 24514 6178
rect 23932 6113 23941 6165
rect 23993 6113 24005 6165
rect 24057 6113 24069 6165
rect 24121 6113 24133 6165
rect 24185 6113 24197 6165
rect 24249 6113 24261 6165
rect 24313 6113 24325 6165
rect 24377 6113 24389 6165
rect 24441 6113 24453 6165
rect 24505 6113 24514 6165
rect 23932 6100 24514 6113
rect 23932 6048 23941 6100
rect 23993 6048 24005 6100
rect 24057 6048 24069 6100
rect 24121 6048 24133 6100
rect 24185 6048 24197 6100
rect 24249 6048 24261 6100
rect 24313 6048 24325 6100
rect 24377 6048 24389 6100
rect 24441 6048 24453 6100
rect 24505 6048 24514 6100
rect 23932 6035 24514 6048
rect 23932 5983 23941 6035
rect 23993 5983 24005 6035
rect 24057 5983 24069 6035
rect 24121 5983 24133 6035
rect 24185 5983 24197 6035
rect 24249 5983 24261 6035
rect 24313 5983 24325 6035
rect 24377 5983 24389 6035
rect 24441 5983 24453 6035
rect 24505 5983 24514 6035
rect 23932 5970 24514 5983
rect 23932 5918 23941 5970
rect 23993 5918 24005 5970
rect 24057 5918 24069 5970
rect 24121 5918 24133 5970
rect 24185 5918 24197 5970
rect 24249 5918 24261 5970
rect 24313 5918 24325 5970
rect 24377 5918 24389 5970
rect 24441 5918 24453 5970
rect 24505 5918 24514 5970
rect 23932 5905 24514 5918
rect 23932 5853 23941 5905
rect 23993 5853 24005 5905
rect 24057 5853 24069 5905
rect 24121 5853 24133 5905
rect 24185 5853 24197 5905
rect 24249 5853 24261 5905
rect 24313 5853 24325 5905
rect 24377 5853 24389 5905
rect 24441 5853 24453 5905
rect 24505 5853 24514 5905
rect 23932 5840 24514 5853
rect 23932 5788 23941 5840
rect 23993 5788 24005 5840
rect 24057 5788 24069 5840
rect 24121 5788 24133 5840
rect 24185 5788 24197 5840
rect 24249 5788 24261 5840
rect 24313 5788 24325 5840
rect 24377 5788 24389 5840
rect 24441 5788 24453 5840
rect 24505 5788 24514 5840
rect 23932 5775 24514 5788
rect 23932 5723 23941 5775
rect 23993 5723 24005 5775
rect 24057 5723 24069 5775
rect 24121 5723 24133 5775
rect 24185 5723 24197 5775
rect 24249 5723 24261 5775
rect 24313 5723 24325 5775
rect 24377 5723 24389 5775
rect 24441 5723 24453 5775
rect 24505 5723 24514 5775
rect 23932 5710 24514 5723
rect 23932 5658 23941 5710
rect 23993 5658 24005 5710
rect 24057 5658 24069 5710
rect 24121 5658 24133 5710
rect 24185 5658 24197 5710
rect 24249 5658 24261 5710
rect 24313 5658 24325 5710
rect 24377 5658 24389 5710
rect 24441 5658 24453 5710
rect 24505 5658 24514 5710
tri 20588 5427 20636 5475 sw
rect 20508 5375 20514 5427
rect 20566 5375 20578 5427
rect 20630 5375 20636 5427
rect 20208 5078 20214 5130
rect 20266 5078 20278 5130
rect 20330 5078 20336 5130
tri 20371 5286 20377 5292 se
rect 20377 5286 20452 5292
rect 20371 5232 20452 5286
tri 20343 5025 20371 5053 se
rect 20371 5025 20423 5232
tri 20423 5203 20452 5232 nw
rect 20208 4973 20214 5025
rect 20266 4973 20278 5025
rect 20330 4973 20423 5025
tri 23907 4270 23932 4295 se
rect 23932 4270 24514 5658
rect 22941 4264 24514 4270
rect 22941 4212 22947 4264
rect 22999 4212 23011 4264
rect 23063 4212 23075 4264
rect 23127 4212 23139 4264
rect 23191 4212 24514 4264
rect 22941 4206 24514 4212
tri 23907 4181 23932 4206 ne
rect 17481 4093 17487 4145
rect 17539 4093 17551 4145
rect 17603 4093 17609 4145
rect 17481 2846 17609 4093
rect 17481 2794 17487 2846
rect 17539 2794 17551 2846
rect 17603 2794 17609 2846
tri 17443 2632 17481 2670 se
rect 17481 2632 17609 2794
rect 16495 2465 16501 2517
rect 16553 2465 16565 2517
rect 16617 2465 16623 2517
rect 17263 2516 17269 2632
rect 17385 2516 17411 2632
rect 17413 2516 17609 2632
tri 17443 2500 17459 2516 ne
rect 17459 2500 17609 2516
tri 17459 2494 17465 2500 ne
rect 17465 2494 17609 2500
rect 19972 3802 20038 3808
rect 19972 3750 19979 3802
rect 20031 3750 20038 3802
rect 19972 3737 20038 3750
rect 19972 3685 19979 3737
rect 20031 3685 20038 3737
rect 19972 3672 20038 3685
rect 19972 3620 19979 3672
rect 20031 3620 20038 3672
rect 19972 3607 20038 3620
rect 19972 3555 19979 3607
rect 20031 3555 20038 3607
rect 19972 3542 20038 3555
rect 19972 3490 19979 3542
rect 20031 3490 20038 3542
rect 19972 3476 20038 3490
rect 19972 3424 19979 3476
rect 20031 3424 20038 3476
rect 19972 3410 20038 3424
rect 19972 3358 19979 3410
rect 20031 3358 20038 3410
rect 19972 3344 20038 3358
rect 19972 3292 19979 3344
rect 20031 3292 20038 3344
rect 19972 3278 20038 3292
rect 19972 3226 19979 3278
rect 20031 3226 20038 3278
rect 19972 3212 20038 3226
rect 19972 3160 19979 3212
rect 20031 3160 20038 3212
rect 19972 3146 20038 3160
rect 19972 3094 19979 3146
rect 20031 3094 20038 3146
rect 19972 3080 20038 3094
rect 19972 3028 19979 3080
rect 20031 3028 20038 3080
rect 19972 3014 20038 3028
rect 19972 2962 19979 3014
rect 20031 2962 20038 3014
rect 19972 2948 20038 2962
rect 19972 2896 19979 2948
rect 20031 2896 20038 2948
rect 19972 2882 20038 2896
rect 19972 2830 19979 2882
rect 20031 2830 20038 2882
rect 19972 2816 20038 2830
rect 19972 2764 19979 2816
rect 20031 2764 20038 2816
rect 19972 2750 20038 2764
rect 19972 2698 19979 2750
rect 20031 2698 20038 2750
rect 19972 2684 20038 2698
rect 19972 2632 19979 2684
rect 20031 2632 20038 2684
rect 19972 2618 20038 2632
rect 19972 2566 19979 2618
rect 20031 2566 20038 2618
rect 19972 2552 20038 2566
rect 19972 2500 19979 2552
rect 20031 2500 20038 2552
rect 19972 2494 20038 2500
rect 20070 3802 20136 3808
rect 20070 3750 20077 3802
rect 20129 3750 20136 3802
rect 20070 3737 20136 3750
rect 20070 3685 20077 3737
rect 20129 3685 20136 3737
rect 20070 3672 20136 3685
rect 20070 3620 20077 3672
rect 20129 3620 20136 3672
rect 20070 3607 20136 3620
rect 20070 3555 20077 3607
rect 20129 3555 20136 3607
rect 20070 3542 20136 3555
rect 20070 3490 20077 3542
rect 20129 3490 20136 3542
rect 20070 3476 20136 3490
rect 20070 3424 20077 3476
rect 20129 3424 20136 3476
rect 20070 3410 20136 3424
rect 20070 3358 20077 3410
rect 20129 3358 20136 3410
rect 20070 3344 20136 3358
rect 20070 3292 20077 3344
rect 20129 3292 20136 3344
rect 20070 3278 20136 3292
rect 20070 3226 20077 3278
rect 20129 3226 20136 3278
rect 20070 3212 20136 3226
rect 20070 3160 20077 3212
rect 20129 3160 20136 3212
rect 20070 3146 20136 3160
rect 20070 3094 20077 3146
rect 20129 3094 20136 3146
rect 20070 3080 20136 3094
rect 20070 3028 20077 3080
rect 20129 3028 20136 3080
rect 20070 3014 20136 3028
rect 20070 2962 20077 3014
rect 20129 2962 20136 3014
rect 20070 2948 20136 2962
rect 20070 2896 20077 2948
rect 20129 2896 20136 2948
rect 20070 2882 20136 2896
rect 20070 2830 20077 2882
rect 20129 2830 20136 2882
rect 20070 2816 20136 2830
rect 20070 2764 20077 2816
rect 20129 2764 20136 2816
rect 20070 2750 20136 2764
rect 20070 2698 20077 2750
rect 20129 2698 20136 2750
rect 20070 2684 20136 2698
rect 20070 2632 20077 2684
rect 20129 2632 20136 2684
rect 20070 2618 20136 2632
rect 20070 2566 20077 2618
rect 20129 2566 20136 2618
rect 20070 2552 20136 2566
rect 20070 2500 20077 2552
rect 20129 2500 20136 2552
rect 20070 2494 20136 2500
rect 16651 2363 16791 2494
tri 16791 2469 16816 2494 nw
tri 17465 2478 17481 2494 ne
tri 16791 2363 16816 2388 sw
rect 12403 2079 12842 2091
rect 12403 2027 12412 2079
rect 12464 2027 12486 2079
rect 12538 2027 12560 2079
rect 12612 2027 12634 2079
rect 12686 2027 12707 2079
rect 12759 2027 12780 2079
rect 12832 2027 12842 2079
rect 12403 2015 12842 2027
rect 12403 1963 12412 2015
rect 12464 1963 12486 2015
rect 12538 1963 12560 2015
rect 12612 1963 12634 2015
rect 12686 1963 12707 2015
rect 12759 1963 12780 2015
rect 12832 1963 12842 2015
rect 12403 1951 12842 1963
rect 12403 1899 12412 1951
rect 12464 1899 12486 1951
rect 12538 1899 12560 1951
rect 12612 1899 12634 1951
rect 12686 1899 12707 1951
rect 12759 1899 12780 1951
rect 12832 1899 12842 1951
rect 16651 1925 16860 2363
rect 12403 1887 12842 1899
rect 12403 1835 12412 1887
rect 12464 1835 12486 1887
rect 12538 1835 12560 1887
rect 12612 1835 12634 1887
rect 12686 1835 12707 1887
rect 12759 1835 12780 1887
rect 12832 1835 12842 1887
tri 17428 1853 17481 1906 se
rect 17481 1853 17609 2494
rect 12403 1823 12842 1835
rect 12403 1771 12412 1823
rect 12464 1771 12486 1823
rect 12538 1771 12560 1823
rect 12612 1771 12634 1823
rect 12686 1771 12707 1823
rect 12759 1771 12780 1823
rect 12832 1771 12842 1823
rect 12403 1562 12842 1771
rect 12403 1510 12409 1562
rect 12461 1510 12484 1562
rect 12536 1510 12559 1562
rect 12611 1510 12634 1562
rect 12686 1510 12709 1562
rect 12761 1510 12784 1562
rect 12836 1510 12842 1562
rect 12403 1498 12842 1510
rect 12403 1446 12409 1498
rect 12461 1446 12484 1498
rect 12536 1446 12559 1498
rect 12611 1446 12634 1498
rect 12686 1446 12709 1498
rect 12761 1446 12784 1498
rect 12836 1446 12842 1498
rect 12403 1445 12842 1446
rect 4424 1338 4436 1390
rect 4372 1332 4488 1338
rect -232 833 75 949
rect 77 905 280 949
tri 280 905 324 949 sw
rect 77 833 324 905
tri 324 833 396 905 sw
tri 232 669 396 833 ne
tri 396 669 560 833 sw
tri 396 505 560 669 ne
tri 560 531 698 669 sw
rect 14251 593 14443 1853
rect 17428 1847 17609 1853
rect 23932 1853 24514 4206
tri 25289 6944 25293 6948 se
rect 25293 6944 25369 6948
tri 25369 6944 25373 6948 nw
tri 28678 6944 28682 6948 ne
rect 28682 6944 28744 6948
tri 28744 6944 28748 6948 sw
rect 25289 3287 25341 6944
tri 25341 6916 25369 6944 nw
tri 28682 6931 28695 6944 ne
rect 28695 6931 28748 6944
tri 28748 6931 28761 6944 sw
tri 28695 6916 28710 6931 ne
rect 28710 6916 28761 6931
tri 28710 6912 28714 6916 ne
rect 28714 6101 28761 6916
rect 28811 6190 28863 9302
rect 28903 6258 28955 9974
rect 28995 6351 29059 10401
rect 29099 6457 29151 10774
rect 29191 6522 29243 11769
rect 29283 6610 29335 13108
tri 29335 6610 29369 6644 sw
rect 29283 6592 29695 6610
tri 29283 6563 29312 6592 ne
rect 29312 6563 29695 6592
tri 29695 6563 29742 6610 sw
tri 29312 6562 29313 6563 ne
rect 29313 6562 29742 6563
tri 29675 6556 29681 6562 ne
rect 29681 6556 29742 6562
tri 29742 6556 29749 6563 sw
tri 29243 6522 29277 6556 sw
tri 29681 6522 29715 6556 ne
rect 29715 6522 29749 6556
tri 29749 6522 29783 6556 sw
rect 29191 6504 29657 6522
tri 29657 6504 29675 6522 sw
tri 29715 6504 29733 6522 ne
rect 29733 6504 29783 6522
tri 29191 6474 29221 6504 ne
rect 29221 6495 29675 6504
tri 29675 6495 29684 6504 sw
tri 29733 6495 29742 6504 ne
rect 29742 6495 29783 6504
tri 29783 6495 29810 6522 sw
rect 29221 6474 29684 6495
tri 29637 6468 29643 6474 ne
rect 29643 6468 29684 6474
tri 29151 6457 29162 6468 sw
tri 29643 6457 29654 6468 ne
rect 29654 6457 29684 6468
tri 29684 6457 29722 6495 sw
tri 29742 6457 29780 6495 ne
rect 29780 6457 29810 6495
tri 29810 6457 29848 6495 sw
rect 29099 6454 29162 6457
tri 29162 6454 29165 6457 sw
tri 29654 6454 29657 6457 ne
rect 29657 6454 29722 6457
rect 29099 6434 29165 6454
tri 29165 6434 29185 6454 sw
tri 29657 6434 29677 6454 ne
rect 29677 6437 29722 6454
tri 29722 6437 29742 6457 sw
tri 29780 6437 29800 6457 ne
rect 29800 6437 29848 6457
rect 29677 6434 29742 6437
rect 29099 6419 29619 6434
tri 29619 6419 29634 6434 sw
tri 29677 6419 29692 6434 ne
rect 29692 6427 29742 6434
tri 29742 6427 29752 6437 sw
tri 29800 6427 29810 6437 ne
rect 29810 6427 29848 6437
tri 29848 6427 29878 6457 sw
rect 29692 6419 29752 6427
rect 29099 6416 29634 6419
tri 29099 6386 29129 6416 ne
rect 29129 6409 29634 6416
tri 29634 6409 29644 6419 sw
tri 29692 6409 29702 6419 ne
rect 29702 6409 29752 6419
rect 29129 6389 29644 6409
tri 29644 6389 29664 6409 sw
tri 29702 6389 29722 6409 ne
rect 29722 6389 29752 6409
tri 29752 6389 29790 6427 sw
tri 29810 6389 29848 6427 ne
rect 29848 6389 29878 6427
tri 29878 6389 29916 6427 sw
rect 29129 6386 29664 6389
tri 29599 6380 29605 6386 ne
rect 29605 6380 29664 6386
tri 29059 6351 29088 6380 sw
tri 29605 6351 29634 6380 ne
rect 29634 6351 29664 6380
tri 29664 6351 29702 6389 sw
tri 29722 6351 29760 6389 ne
rect 29760 6369 29790 6389
tri 29790 6369 29810 6389 sw
tri 29848 6369 29868 6389 ne
rect 29868 6369 29916 6389
rect 29760 6359 29810 6369
tri 29810 6359 29820 6369 sw
tri 29868 6359 29878 6369 ne
rect 29878 6359 29916 6369
tri 29916 6359 29946 6389 sw
rect 29760 6351 29820 6359
rect 28995 6346 29088 6351
tri 29088 6346 29093 6351 sw
tri 29634 6346 29639 6351 ne
rect 29639 6346 29702 6351
rect 28995 6328 29581 6346
tri 28995 6313 29010 6328 ne
rect 29010 6313 29581 6328
tri 29581 6313 29614 6346 sw
tri 29639 6313 29672 6346 ne
rect 29672 6341 29702 6346
tri 29702 6341 29712 6351 sw
tri 29760 6341 29770 6351 ne
rect 29770 6341 29820 6351
rect 29672 6321 29712 6341
tri 29712 6321 29732 6341 sw
tri 29770 6321 29790 6341 ne
rect 29790 6321 29820 6341
tri 29820 6321 29858 6359 sw
tri 29878 6321 29916 6359 ne
rect 29916 6321 29946 6359
tri 29946 6321 29984 6359 sw
rect 29672 6313 29732 6321
tri 29010 6298 29025 6313 ne
rect 29025 6303 29614 6313
tri 29614 6303 29624 6313 sw
tri 29672 6303 29682 6313 ne
rect 29682 6303 29732 6313
rect 29025 6298 29624 6303
tri 29561 6292 29567 6298 ne
rect 29567 6292 29624 6298
tri 28955 6258 28989 6292 sw
tri 29567 6258 29601 6292 ne
rect 29601 6283 29624 6292
tri 29624 6283 29644 6303 sw
tri 29682 6283 29702 6303 ne
rect 29702 6283 29732 6303
tri 29732 6283 29770 6321 sw
tri 29790 6283 29828 6321 ne
rect 29828 6301 29858 6321
tri 29858 6301 29878 6321 sw
tri 29916 6301 29936 6321 ne
rect 29936 6301 29984 6321
rect 29828 6291 29878 6301
tri 29878 6291 29888 6301 sw
tri 29936 6291 29946 6301 ne
rect 29946 6291 29984 6301
tri 29984 6291 30014 6321 sw
rect 29828 6283 29888 6291
rect 29601 6258 29644 6283
rect 28903 6245 29543 6258
tri 29543 6245 29556 6258 sw
tri 29601 6245 29614 6258 ne
rect 29614 6245 29644 6258
tri 29644 6245 29682 6283 sw
tri 29702 6245 29740 6283 ne
rect 29740 6273 29770 6283
tri 29770 6273 29780 6283 sw
tri 29828 6273 29838 6283 ne
rect 29838 6273 29888 6283
rect 29740 6253 29780 6273
tri 29780 6253 29800 6273 sw
tri 29838 6253 29858 6273 ne
rect 29858 6253 29888 6273
tri 29888 6253 29926 6291 sw
tri 29946 6253 29984 6291 ne
rect 29984 6253 30014 6291
tri 30014 6253 30052 6291 sw
rect 29740 6245 29800 6253
rect 28903 6240 29556 6245
tri 28903 6210 28933 6240 ne
rect 28933 6210 29556 6240
tri 29523 6207 29526 6210 ne
rect 29526 6207 29556 6210
tri 29556 6207 29594 6245 sw
tri 29614 6207 29652 6245 ne
rect 29652 6235 29682 6245
tri 29682 6235 29692 6245 sw
tri 29740 6235 29750 6245 ne
rect 29750 6235 29800 6245
rect 29652 6215 29692 6235
tri 29692 6215 29712 6235 sw
tri 29750 6215 29770 6235 ne
rect 29770 6215 29800 6235
tri 29800 6215 29838 6253 sw
tri 29858 6215 29896 6253 ne
rect 29896 6233 29926 6253
tri 29926 6233 29946 6253 sw
tri 29984 6233 30004 6253 ne
rect 30004 6233 30052 6253
rect 29896 6223 29946 6233
tri 29946 6223 29956 6233 sw
tri 30004 6223 30014 6233 ne
rect 30014 6223 30052 6233
tri 30052 6223 30082 6253 sw
rect 29896 6215 29956 6223
rect 29652 6207 29712 6215
tri 29526 6203 29530 6207 ne
rect 29530 6203 29594 6207
tri 28863 6190 28876 6203 sw
tri 29530 6190 29543 6203 ne
rect 29543 6197 29594 6203
tri 29594 6197 29604 6207 sw
tri 29652 6197 29662 6207 ne
rect 29662 6197 29712 6207
rect 29543 6190 29604 6197
rect 28811 6170 28876 6190
tri 28876 6170 28896 6190 sw
tri 29543 6170 29563 6190 ne
rect 29563 6177 29604 6190
tri 29604 6177 29624 6197 sw
tri 29662 6177 29682 6197 ne
rect 29682 6177 29712 6197
tri 29712 6177 29750 6215 sw
tri 29770 6177 29808 6215 ne
rect 29808 6205 29838 6215
tri 29838 6205 29848 6215 sw
tri 29896 6205 29906 6215 ne
rect 29906 6205 29956 6215
rect 29808 6185 29848 6205
tri 29848 6185 29868 6205 sw
tri 29906 6185 29926 6205 ne
rect 29926 6185 29956 6205
tri 29956 6185 29994 6223 sw
tri 30014 6203 30034 6223 ne
rect 29808 6177 29868 6185
rect 29563 6170 29624 6177
rect 28811 6169 29505 6170
tri 29505 6169 29506 6170 sw
tri 29563 6169 29564 6170 ne
rect 29564 6169 29624 6170
rect 28811 6159 29506 6169
tri 29506 6159 29516 6169 sw
tri 29564 6159 29574 6169 ne
rect 29574 6159 29624 6169
rect 28811 6151 29516 6159
tri 28811 6122 28840 6151 ne
rect 28840 6139 29516 6151
tri 29516 6139 29536 6159 sw
tri 29574 6139 29594 6159 ne
rect 29594 6139 29624 6159
tri 29624 6139 29662 6177 sw
tri 29682 6139 29720 6177 ne
rect 29720 6167 29750 6177
tri 29750 6167 29760 6177 sw
tri 29808 6167 29818 6177 ne
rect 29818 6167 29868 6177
rect 29720 6147 29760 6167
tri 29760 6147 29780 6167 sw
tri 29818 6147 29838 6167 ne
rect 29838 6165 29868 6167
tri 29868 6165 29888 6185 sw
tri 29926 6165 29946 6185 ne
rect 29838 6147 29888 6165
tri 29888 6147 29906 6165 sw
rect 29720 6139 29780 6147
rect 28840 6122 29536 6139
tri 29485 6120 29487 6122 ne
rect 29487 6120 29536 6122
tri 28761 6101 28780 6120 sw
tri 29487 6101 29506 6120 ne
rect 29506 6101 29536 6120
tri 29536 6101 29574 6139 sw
tri 29594 6101 29632 6139 ne
rect 29632 6129 29662 6139
tri 29662 6129 29672 6139 sw
tri 29720 6129 29730 6139 ne
rect 29730 6129 29780 6139
rect 29632 6109 29672 6129
tri 29672 6109 29692 6129 sw
tri 29730 6109 29750 6129 ne
rect 29750 6127 29780 6129
tri 29780 6127 29800 6147 sw
tri 29838 6127 29858 6147 ne
rect 29750 6109 29800 6127
tri 29800 6109 29818 6127 sw
rect 29632 6101 29692 6109
rect 28714 6082 28780 6101
tri 28780 6082 28799 6101 sw
tri 29506 6082 29525 6101 ne
rect 29525 6091 29574 6101
tri 29574 6091 29584 6101 sw
tri 29632 6091 29642 6101 ne
rect 29642 6091 29692 6101
rect 29525 6082 29584 6091
rect 28714 6063 29467 6082
tri 29467 6063 29486 6082 sw
tri 29525 6063 29544 6082 ne
rect 29544 6071 29584 6082
tri 29584 6071 29604 6091 sw
tri 29642 6071 29662 6091 ne
rect 29662 6089 29692 6091
tri 29692 6089 29712 6109 sw
tri 29750 6089 29770 6109 ne
rect 29662 6071 29712 6089
tri 29712 6071 29730 6089 sw
rect 29544 6063 29604 6071
tri 28714 6034 28743 6063 ne
rect 28743 6053 29486 6063
tri 29486 6053 29496 6063 sw
tri 29544 6053 29554 6063 ne
rect 29554 6053 29604 6063
rect 28743 6034 29496 6053
tri 29447 5995 29486 6034 ne
rect 29486 6033 29496 6034
tri 29496 6033 29516 6053 sw
tri 29554 6033 29574 6053 ne
rect 29574 6051 29604 6053
tri 29604 6051 29624 6071 sw
tri 29662 6051 29682 6071 ne
rect 29574 6033 29624 6051
tri 29624 6033 29642 6051 sw
rect 29486 6013 29516 6033
tri 29516 6013 29536 6033 sw
tri 29574 6013 29594 6033 ne
rect 29486 5995 29536 6013
tri 29536 5995 29554 6013 sw
tri 29486 5975 29506 5995 ne
tri 25341 3287 25363 3309 sw
tri 25289 3213 25363 3287 ne
tri 25363 3213 25437 3287 sw
tri 25363 3212 25364 3213 ne
rect 25364 3212 25437 3213
tri 25364 3148 25428 3212 ne
rect 25428 3148 25437 3212
tri 25428 3139 25437 3148 ne
tri 25437 3139 25511 3213 sw
tri 25437 3065 25511 3139 ne
tri 25511 3065 25585 3139 sw
tri 25511 2991 25585 3065 ne
tri 25585 2991 25659 3065 sw
tri 25585 2956 25620 2991 ne
rect 25620 2956 25659 2991
tri 25620 2917 25659 2956 ne
tri 25659 2951 25699 2991 sw
rect 25659 2917 25699 2951
tri 25699 2917 25733 2951 sw
tri 25659 2877 25699 2917 ne
rect 25699 2899 25733 2917
tri 25733 2899 25751 2917 sw
tri 24514 1853 24571 1910 sw
rect 17480 1795 17492 1847
rect 17544 1795 17556 1847
rect 17608 1795 17609 1847
rect 17428 1735 17609 1795
rect 17480 1683 17492 1735
rect 17544 1683 17556 1735
rect 17608 1683 17609 1735
rect 17428 1677 17609 1683
rect 23161 788 23213 1852
rect 23932 1845 24571 1853
tri 24571 1845 24579 1853 sw
rect 23932 1616 24579 1845
tri 24579 1616 24808 1845 sw
rect 23932 1606 24808 1616
tri 24808 1606 24818 1616 sw
tri 25689 1606 25699 1616 se
rect 25699 1606 25751 2899
tri 25751 1606 25765 1620 sw
rect 23932 1600 24818 1606
tri 24818 1600 24824 1606 sw
rect 25689 1600 25765 1606
tri 23890 1548 23932 1590 se
rect 23932 1548 24824 1600
tri 24824 1548 24876 1600 sw
rect 25689 1548 25701 1600
rect 25753 1548 25765 1600
tri 23867 1525 23890 1548 se
rect 23890 1525 24876 1548
tri 24876 1525 24899 1548 sw
rect 25689 1525 25765 1548
tri 23815 1473 23867 1525 se
rect 23867 1516 24899 1525
tri 24899 1516 24908 1525 sw
rect 23867 1473 24908 1516
tri 24908 1473 24951 1516 sw
rect 25689 1473 25701 1525
rect 25753 1473 25765 1525
tri 23791 1449 23815 1473 se
rect 23815 1449 24951 1473
tri 24951 1449 24975 1473 sw
rect 25689 1449 25765 1473
tri 23739 1397 23791 1449 se
rect 23791 1397 24975 1449
tri 24975 1397 25027 1449 sw
rect 25689 1397 25701 1449
rect 25753 1397 25765 1449
tri 23665 1323 23739 1397 se
rect 23739 1391 25027 1397
rect 23739 1323 24071 1391
tri 24071 1323 24139 1391 nw
tri 24511 1323 24579 1391 ne
rect 24579 1323 25027 1391
tri 25027 1323 25101 1397 sw
rect 25689 1391 25765 1397
tri 23571 1229 23665 1323 se
rect 23665 1229 23977 1323
tri 23977 1229 24071 1323 nw
tri 24579 1229 24673 1323 ne
rect 24673 1229 25101 1323
rect 23571 1213 23961 1229
tri 23961 1213 23977 1229 nw
tri 24673 1213 24689 1229 ne
rect 24689 1213 25101 1229
rect 23571 969 23577 1213
rect 23757 1172 23920 1213
tri 23920 1172 23961 1213 nw
tri 24689 1172 24730 1213 ne
rect 24730 1172 25101 1213
rect 23757 1120 23868 1172
tri 23868 1120 23920 1172 nw
tri 24730 1120 24782 1172 ne
rect 24782 1120 25101 1172
rect 23757 1108 23856 1120
tri 23856 1108 23868 1120 nw
tri 24782 1108 24794 1120 ne
rect 24794 1108 25101 1120
rect 23757 1056 23804 1108
tri 23804 1056 23856 1108 nw
tri 24794 1056 24846 1108 ne
rect 24846 1056 25101 1108
rect 23757 1044 23792 1056
tri 23792 1044 23804 1056 nw
tri 24846 1044 24858 1056 ne
rect 24858 1044 25101 1056
rect 23757 1033 23781 1044
tri 23781 1033 23792 1044 nw
tri 24858 1033 24869 1044 ne
rect 24869 1033 25101 1044
rect 23693 992 23740 1033
tri 23740 992 23781 1033 nw
tri 24869 994 24908 1033 ne
rect 23693 980 23728 992
tri 23728 980 23740 992 nw
rect 23693 969 23717 980
tri 23717 969 23728 980 nw
rect 23571 957 23676 969
rect 23571 905 23577 957
rect 23629 928 23676 957
tri 23676 928 23717 969 nw
rect 23629 905 23653 928
tri 23653 905 23676 928 nw
rect 560 505 753 531
rect 24908 510 25101 1033
rect 27001 1172 27385 1516
rect 27001 1120 27015 1172
rect 27067 1120 27090 1172
rect 27142 1120 27165 1172
rect 27217 1120 27240 1172
rect 27292 1120 27314 1172
rect 27366 1120 27385 1172
rect 27001 1108 27385 1120
rect 27001 1056 27015 1108
rect 27067 1056 27090 1108
rect 27142 1056 27165 1108
rect 27217 1056 27240 1108
rect 27292 1056 27314 1108
rect 27366 1056 27385 1108
rect 27001 1044 27385 1056
rect 27001 992 27015 1044
rect 27067 992 27090 1044
rect 27142 992 27165 1044
rect 27217 992 27240 1044
rect 27292 992 27314 1044
rect 27366 992 27385 1044
rect 27001 980 27385 992
rect 27001 928 27015 980
rect 27067 928 27090 980
rect 27142 928 27165 980
rect 27217 928 27240 980
rect 27292 928 27314 980
rect 27366 928 27385 980
tri 560 415 650 505 ne
rect 650 415 753 505
rect 27001 -747 27385 928
tri 29502 339 29506 343 se
rect 29506 339 29554 5995
tri 29590 1263 29594 1267 se
rect 29594 1263 29642 6033
tri 29678 2187 29682 2191 se
rect 29682 2187 29730 6071
tri 29766 3111 29770 3115 se
rect 29770 3111 29818 6109
tri 29854 4035 29858 4039 se
rect 29858 4035 29906 6147
tri 29942 4959 29946 4963 se
rect 29946 4959 29994 6185
tri 30030 5883 30034 5887 se
rect 30034 5883 30082 6223
tri 30082 5883 30086 5887 sw
rect 30030 5874 30086 5883
rect 30030 5794 30086 5818
rect 30030 5729 30086 5738
tri 29994 4959 29998 4963 sw
rect 29942 4950 29998 4959
rect 29942 4870 29998 4894
rect 29942 4805 29998 4814
tri 29906 4035 29910 4039 sw
rect 29854 4026 29910 4035
rect 29854 3946 29910 3970
rect 29854 3881 29910 3890
tri 29854 3877 29858 3881 ne
rect 29858 3877 29906 3881
tri 29906 3877 29910 3881 nw
tri 29818 3111 29822 3115 sw
rect 29766 3102 29822 3111
rect 29766 3022 29822 3046
rect 29766 2957 29822 2966
tri 29730 2187 29734 2191 sw
rect 29678 2178 29734 2187
rect 29678 2098 29734 2122
rect 29678 2033 29734 2042
tri 29642 1263 29646 1267 sw
rect 29590 1254 29646 1263
rect 29590 1174 29646 1198
rect 29590 1109 29646 1118
tri 29554 339 29558 343 sw
rect 29502 330 29558 339
rect 29502 250 29558 274
rect 29502 185 29558 194
tri 27001 -833 27087 -747 ne
tri 27001 -1361 27087 -1275 se
rect 27087 -1361 27385 -747
rect 23583 -1899 23839 -1783
rect 24908 -1953 25101 -1909
rect 23037 -2275 23089 -2253
rect 23867 -2273 24123 -2103
rect 27001 -2273 27385 -1361
rect 28226 -2129 28278 -2077
rect 20884 -2464 20936 -2425
<< rmetal2 >>
rect 25332 10682 25384 10684
rect 13292 2646 13408 2648
rect 13399 2433 13401 2564
rect 17411 2516 17413 2632
rect 75 833 77 949
<< via2 >>
rect 30030 5818 30086 5874
rect 30030 5738 30086 5794
rect 29942 4894 29998 4950
rect 29942 4814 29998 4870
rect 29854 3970 29910 4026
rect 29854 3890 29910 3946
rect 29766 3046 29822 3102
rect 29766 2966 29822 3022
rect 29678 2122 29734 2178
rect 29678 2042 29734 2098
rect 29590 1198 29646 1254
rect 29590 1118 29646 1174
rect 29502 274 29558 330
rect 29502 194 29558 250
<< metal3 >>
rect 30025 5874 30091 5879
rect 30025 5873 30030 5874
rect 30086 5873 30091 5874
rect 30025 5809 30027 5873
rect 30025 5794 30091 5809
rect 30025 5793 30030 5794
rect 30086 5793 30091 5794
rect 30025 5733 30027 5793
tri 30025 5731 30027 5733 ne
rect 30027 5723 30091 5729
rect 29937 4950 30003 4955
rect 29937 4949 29942 4950
rect 29998 4949 30003 4950
rect 29937 4885 29939 4949
rect 29937 4870 30003 4885
rect 29937 4869 29942 4870
rect 29998 4869 30003 4870
rect 29937 4809 29939 4869
tri 29937 4807 29939 4809 ne
rect 29939 4799 30003 4805
rect 11695 3983 11921 4069
rect 29849 4026 29915 4031
rect 29849 4025 29854 4026
rect 29910 4025 29915 4026
rect 29849 3961 29851 4025
rect 29849 3946 29915 3961
rect 29849 3945 29854 3946
rect 29910 3945 29915 3946
rect 29849 3885 29851 3945
tri 29849 3883 29851 3885 ne
rect 29851 3875 29915 3881
rect 29761 3102 29827 3107
rect 29761 3101 29766 3102
rect 29822 3101 29827 3102
rect 29761 3037 29763 3101
rect 29761 3022 29827 3037
rect 29761 3021 29766 3022
rect 29822 3021 29827 3022
rect 29761 2961 29763 3021
tri 29761 2959 29763 2961 ne
rect 29763 2951 29827 2957
rect 29673 2178 29739 2183
rect 29673 2177 29678 2178
rect 29734 2177 29739 2178
rect 29673 2113 29675 2177
rect 29673 2098 29739 2113
rect 29673 2097 29678 2098
rect 29734 2097 29739 2098
rect 29673 2037 29675 2097
tri 29673 2035 29675 2037 ne
rect 29675 2027 29739 2033
rect 29585 1254 29651 1259
rect 29585 1253 29590 1254
rect 29646 1253 29651 1254
rect 29585 1189 29587 1253
rect 29585 1174 29651 1189
rect 29585 1173 29590 1174
rect 29646 1173 29651 1174
rect 29585 1113 29587 1173
tri 29585 1111 29587 1113 ne
rect 29587 1103 29651 1109
rect 29497 330 29563 335
rect 29497 329 29502 330
rect 29558 329 29563 330
rect 29497 265 29499 329
rect 29497 250 29563 265
rect 29497 249 29502 250
rect 29558 249 29563 250
rect 29497 189 29499 249
tri 29497 187 29499 189 ne
rect 29499 179 29563 185
<< via3 >>
rect 30027 5818 30030 5873
rect 30030 5818 30086 5873
rect 30086 5818 30091 5873
rect 30027 5809 30091 5818
rect 30027 5738 30030 5793
rect 30030 5738 30086 5793
rect 30086 5738 30091 5793
rect 30027 5729 30091 5738
rect 29939 4894 29942 4949
rect 29942 4894 29998 4949
rect 29998 4894 30003 4949
rect 29939 4885 30003 4894
rect 29939 4814 29942 4869
rect 29942 4814 29998 4869
rect 29998 4814 30003 4869
rect 29939 4805 30003 4814
rect 29851 3970 29854 4025
rect 29854 3970 29910 4025
rect 29910 3970 29915 4025
rect 29851 3961 29915 3970
rect 29851 3890 29854 3945
rect 29854 3890 29910 3945
rect 29910 3890 29915 3945
rect 29851 3881 29915 3890
rect 29763 3046 29766 3101
rect 29766 3046 29822 3101
rect 29822 3046 29827 3101
rect 29763 3037 29827 3046
rect 29763 2966 29766 3021
rect 29766 2966 29822 3021
rect 29822 2966 29827 3021
rect 29763 2957 29827 2966
rect 29675 2122 29678 2177
rect 29678 2122 29734 2177
rect 29734 2122 29739 2177
rect 29675 2113 29739 2122
rect 29675 2042 29678 2097
rect 29678 2042 29734 2097
rect 29734 2042 29739 2097
rect 29675 2033 29739 2042
rect 29587 1198 29590 1253
rect 29590 1198 29646 1253
rect 29646 1198 29651 1253
rect 29587 1189 29651 1198
rect 29587 1118 29590 1173
rect 29590 1118 29646 1173
rect 29646 1118 29651 1173
rect 29587 1109 29651 1118
rect 29499 274 29502 329
rect 29502 274 29558 329
rect 29558 274 29563 329
rect 29499 265 29563 274
rect 29499 194 29502 249
rect 29502 194 29558 249
rect 29558 194 29563 249
rect 29499 185 29563 194
<< metal4 >>
rect 29498 329 29536 330
rect 29498 265 29499 329
rect 29498 249 29536 265
rect 29498 185 29499 249
rect 29498 184 29536 185
tri 29498 146 29536 184 ne
<< via4 >>
rect 29536 5873 30092 5874
rect 29536 5809 30027 5873
rect 30027 5809 30091 5873
rect 30091 5809 30092 5873
rect 29536 5793 30092 5809
rect 29536 5729 30027 5793
rect 30027 5729 30091 5793
rect 30091 5729 30092 5793
rect 29536 5318 30092 5729
rect 29536 4949 30092 4950
rect 29536 4885 29939 4949
rect 29939 4885 30003 4949
rect 30003 4885 30092 4949
rect 29536 4869 30092 4885
rect 29536 4805 29939 4869
rect 29939 4805 30003 4869
rect 30003 4805 30092 4869
rect 29536 4394 30092 4805
rect 29536 4025 30092 4026
rect 29536 3961 29851 4025
rect 29851 3961 29915 4025
rect 29915 3961 30092 4025
rect 29536 3945 30092 3961
rect 29536 3881 29851 3945
rect 29851 3881 29915 3945
rect 29915 3881 30092 3945
rect 29536 3470 30092 3881
rect 29536 3101 30092 3102
rect 29536 3037 29763 3101
rect 29763 3037 29827 3101
rect 29827 3037 30092 3101
rect 29536 3021 30092 3037
rect 29536 2957 29763 3021
rect 29763 2957 29827 3021
rect 29827 2957 30092 3021
rect 29536 2546 30092 2957
rect 29536 2177 30092 2178
rect 29536 2113 29675 2177
rect 29675 2113 29739 2177
rect 29739 2113 30092 2177
rect 29536 2097 30092 2113
rect 29536 2033 29675 2097
rect 29675 2033 29739 2097
rect 29739 2033 30092 2097
rect 29536 1622 30092 2033
rect 29536 1253 30092 1254
rect 29536 1189 29587 1253
rect 29587 1189 29651 1253
rect 29651 1189 30092 1253
rect 29536 1173 30092 1189
rect 29536 1109 29587 1173
rect 29587 1109 29651 1173
rect 29651 1109 30092 1173
rect 29536 698 30092 1109
rect 29536 329 30092 330
rect 29536 265 29563 329
rect 29563 265 30092 329
rect 29536 249 30092 265
rect 29536 185 29563 249
rect 29563 185 30092 249
rect 29536 -226 30092 185
<< metal5 >>
rect 29512 5874 30116 5898
rect 29512 5318 29536 5874
rect 30092 5318 30116 5874
rect 29512 5294 30116 5318
rect 29512 4950 30116 4974
rect 29512 4394 29536 4950
rect 30092 4394 30116 4950
rect 29512 4370 30116 4394
rect 29512 4026 30116 4050
rect 29512 3470 29536 4026
rect 30092 3470 30116 4026
rect 29512 3446 30116 3470
rect 29512 3102 30116 3126
rect 29512 2546 29536 3102
rect 30092 2546 30116 3102
rect 29512 2522 30116 2546
rect 29512 2178 30116 2202
rect 29512 1622 29536 2178
rect 30092 1622 30116 2178
rect 29512 1598 30116 1622
rect 29512 1254 30116 1278
rect 29512 698 29536 1254
rect 30092 698 30116 1254
rect 29512 674 30116 698
rect 29512 330 30116 354
rect 29512 -226 29536 330
rect 30092 -226 30116 330
rect 29512 -250 30116 -226
<< comment >>
tri 26894 12551 26917 12552 se
rect 26917 12551 26964 12552
tri 26964 12551 26987 12552 sw
tri 26872 12549 26894 12551 se
rect 26894 12549 26987 12551
tri 26987 12549 27009 12551 sw
tri 26850 12546 26872 12549 se
rect 26872 12546 27009 12549
tri 27009 12546 27031 12549 sw
tri 26829 12543 26850 12546 se
rect 26850 12543 27031 12546
tri 27031 12543 27052 12546 sw
tri 26809 12539 26829 12543 se
rect 26829 12539 27052 12543
tri 27052 12539 27072 12543 sw
tri 26791 12535 26809 12539 se
rect 26809 12535 27072 12539
tri 27072 12535 27091 12539 sw
tri 26773 12530 26791 12535 se
rect 26791 12530 27091 12535
tri 27091 12530 27108 12535 sw
tri 26758 12525 26773 12530 se
rect 26773 12525 27108 12530
tri 27108 12525 27123 12530 sw
tri 26744 12519 26758 12525 se
rect 26758 12519 27123 12525
tri 27123 12519 27137 12525 sw
tri 26732 12512 26744 12519 se
rect 26744 12512 27137 12519
tri 27137 12512 27149 12519 sw
tri 26722 12506 26732 12512 se
rect 26732 12506 27149 12512
tri 27149 12506 27159 12512 sw
tri 26714 12499 26722 12506 se
rect 26722 12499 27159 12506
tri 27159 12499 27167 12506 sw
tri 26709 12492 26714 12499 se
rect 26714 12492 27167 12499
tri 27167 12492 27173 12499 sw
tri 26705 12484 26709 12492 se
rect 26709 12484 27173 12492
tri 27173 12484 27176 12492 sw
tri 26704 12477 26705 12484 se
tri 26704 12470 26705 12477 ne
rect 26705 12470 27176 12484
tri 27176 12477 27177 12484 sw
tri 27176 12470 27177 12477 nw
tri 26705 12462 26709 12470 ne
rect 26709 12462 27173 12470
tri 27173 12462 27176 12470 nw
tri 26709 12455 26714 12462 ne
rect 26714 12455 27167 12462
tri 27167 12455 27173 12462 nw
tri 26714 12448 26722 12455 ne
rect 26722 12448 27159 12455
tri 27159 12448 27167 12455 nw
tri 26722 12442 26732 12448 ne
rect 26732 12442 27149 12448
tri 27149 12442 27159 12448 nw
tri 26732 12435 26744 12442 ne
rect 26744 12435 27137 12442
tri 27137 12435 27149 12442 nw
tri 26744 12429 26758 12435 ne
rect 26758 12429 27123 12435
tri 27123 12429 27137 12435 nw
tri 26758 12424 26773 12429 ne
rect 26773 12424 27108 12429
tri 27108 12424 27123 12429 nw
tri 26773 12419 26791 12424 ne
rect 26791 12419 27091 12424
tri 27091 12419 27108 12424 nw
tri 26791 12415 26809 12419 ne
rect 26809 12415 27072 12419
tri 27072 12415 27091 12419 nw
tri 26809 12411 26829 12415 ne
rect 26829 12411 27052 12415
tri 27052 12411 27072 12415 nw
tri 26829 12408 26850 12411 ne
rect 26850 12408 27031 12411
tri 27031 12408 27052 12411 nw
tri 26850 12405 26872 12408 ne
rect 26872 12405 27009 12408
tri 27009 12405 27031 12408 nw
tri 26872 12403 26894 12405 ne
rect 26894 12403 26987 12405
tri 26987 12403 27009 12405 nw
tri 26894 12402 26917 12403 ne
rect 26917 12402 26964 12403
tri 26964 12402 26987 12403 nw
tri 25598 11882 25605 11883 se
tri 25605 11882 25612 11883 sw
tri 25590 11878 25598 11882 se
rect 25598 11878 25612 11882
tri 25612 11878 25620 11882 sw
tri 25583 11871 25590 11878 se
rect 25590 11871 25620 11878
tri 25620 11871 25627 11878 sw
tri 25576 11863 25583 11871 se
rect 25583 11863 25627 11871
tri 25627 11863 25634 11871 sw
tri 25570 11851 25576 11863 se
rect 25576 11851 25634 11863
tri 25634 11851 25640 11863 sw
tri 25563 11838 25570 11851 se
rect 25570 11838 25640 11851
tri 25640 11838 25647 11851 sw
tri 25557 11822 25563 11838 se
rect 25563 11822 25647 11838
tri 25647 11822 25653 11838 sw
tri 25552 11805 25557 11822 se
rect 25557 11805 25653 11822
tri 25653 11805 25658 11822 sw
tri 25547 11785 25552 11805 se
rect 25552 11785 25658 11805
tri 25658 11785 25663 11805 sw
tri 25543 11764 25547 11785 se
rect 25547 11764 25663 11785
tri 25663 11764 25667 11785 sw
tri 25539 11742 25543 11764 se
rect 25543 11742 25667 11764
tri 25667 11742 25671 11764 sw
tri 25536 11718 25539 11742 se
rect 25539 11718 25671 11742
tri 25671 11718 25674 11742 sw
tri 25533 11693 25536 11718 se
rect 25536 11693 25674 11718
tri 25674 11693 25677 11718 sw
tri 25531 11668 25533 11693 se
rect 25533 11668 25677 11693
tri 25677 11668 25679 11693 sw
tri 25530 11642 25531 11668 se
rect 25531 11642 25679 11668
tri 25679 11642 25680 11668 sw
rect 25530 11589 25680 11642
tri 25530 11563 25531 11589 ne
rect 25531 11563 25679 11589
tri 25679 11563 25680 11589 nw
tri 25531 11538 25533 11563 ne
rect 25533 11538 25677 11563
tri 25677 11538 25679 11563 nw
tri 25533 11513 25536 11538 ne
rect 25536 11513 25674 11538
tri 25674 11513 25677 11538 nw
tri 25536 11489 25539 11513 ne
rect 25539 11489 25671 11513
tri 25671 11489 25674 11513 nw
tri 25539 11467 25543 11489 ne
rect 25543 11467 25667 11489
tri 25667 11467 25671 11489 nw
tri 25543 11446 25547 11467 ne
rect 25547 11446 25663 11467
tri 25663 11446 25667 11467 nw
tri 25547 11426 25552 11446 ne
rect 25552 11426 25658 11446
tri 25658 11426 25663 11446 nw
tri 25552 11409 25557 11426 ne
rect 25557 11409 25653 11426
tri 25653 11409 25658 11426 nw
tri 25557 11393 25563 11409 ne
rect 25563 11393 25647 11409
tri 25647 11393 25653 11409 nw
tri 25563 11379 25570 11393 ne
rect 25570 11379 25640 11393
tri 25640 11379 25647 11393 nw
tri 25570 11368 25576 11379 ne
rect 25576 11368 25634 11379
tri 25634 11368 25640 11379 nw
tri 25576 11359 25583 11368 ne
rect 25583 11359 25627 11368
tri 25627 11359 25634 11368 nw
tri 25583 11353 25590 11359 ne
rect 25590 11353 25620 11359
tri 25620 11353 25627 11359 nw
tri 25590 11349 25598 11353 ne
rect 25598 11349 25612 11353
tri 25612 11349 25620 11353 nw
tri 25598 11348 25605 11349 ne
tri 25605 11348 25612 11349 nw
tri 26168 10971 26189 10972 se
rect 26189 10971 26232 10972
tri 26232 10971 26253 10972 sw
tri 26147 10970 26168 10971 se
rect 26168 10970 26253 10971
tri 26253 10970 26274 10971 sw
tri 26127 10968 26147 10970 se
rect 26147 10968 26274 10970
tri 26274 10968 26294 10970 sw
tri 26107 10966 26127 10968 se
rect 26127 10966 26294 10968
tri 26294 10966 26313 10968 sw
tri 26089 10964 26107 10966 se
rect 26107 10964 26313 10966
tri 26313 10964 26332 10966 sw
tri 26072 10961 26089 10964 se
rect 26089 10961 26332 10964
tri 26332 10961 26349 10964 sw
tri 26056 10957 26072 10961 se
rect 26072 10957 26349 10961
tri 26349 10957 26365 10961 sw
tri 26041 10954 26056 10957 se
rect 26056 10954 26365 10957
tri 26365 10954 26379 10957 sw
tri 26029 10950 26041 10954 se
rect 26041 10950 26379 10954
tri 26379 10950 26392 10954 sw
tri 26018 10946 26029 10950 se
rect 26029 10946 26392 10950
tri 26392 10946 26403 10950 sw
tri 26008 10942 26018 10946 se
rect 26018 10942 26403 10946
tri 26403 10942 26412 10946 sw
tri 26001 10937 26008 10942 se
rect 26008 10937 26412 10942
tri 26412 10937 26420 10942 sw
tri 25996 10932 26001 10937 se
rect 26001 10932 26420 10937
tri 26420 10932 26425 10937 sw
tri 25993 10928 25996 10932 se
rect 25996 10928 26425 10932
tri 26425 10928 26428 10932 sw
tri 25992 10923 25993 10928 se
tri 25992 10918 25993 10923 ne
rect 25993 10918 26428 10928
tri 26428 10923 26429 10928 sw
tri 26428 10918 26429 10923 nw
tri 25993 10913 25996 10918 ne
rect 25996 10913 26425 10918
tri 26425 10913 26428 10918 nw
tri 25996 10909 26001 10913 ne
rect 26001 10909 26420 10913
tri 26420 10909 26425 10913 nw
tri 26001 10904 26008 10909 ne
rect 26008 10904 26412 10909
tri 26412 10904 26420 10909 nw
tri 26008 10900 26018 10904 ne
rect 26018 10900 26403 10904
tri 26403 10900 26412 10904 nw
tri 26018 10896 26029 10900 ne
rect 26029 10896 26392 10900
tri 26392 10896 26403 10900 nw
tri 26029 10892 26041 10896 ne
rect 26041 10892 26379 10896
tri 26379 10892 26392 10896 nw
tri 26041 10888 26056 10892 ne
rect 26056 10888 26365 10892
tri 26365 10888 26379 10892 nw
tri 26056 10885 26072 10888 ne
rect 26072 10885 26349 10888
tri 26349 10885 26365 10888 nw
tri 26072 10882 26089 10885 ne
rect 26089 10882 26332 10885
tri 26332 10882 26349 10885 nw
tri 26089 10880 26107 10882 ne
rect 26107 10880 26313 10882
tri 26313 10880 26332 10882 nw
tri 26107 10878 26127 10880 ne
rect 26127 10878 26294 10880
tri 26294 10878 26313 10880 nw
tri 26127 10876 26147 10878 ne
rect 26147 10876 26274 10878
tri 26274 10876 26294 10878 nw
tri 26450 10876 26455 10877 se
tri 26455 10876 26460 10877 sw
tri 26147 10875 26168 10876 ne
rect 26168 10875 26253 10876
tri 26253 10875 26274 10876 nw
tri 26448 10875 26450 10876 se
rect 26450 10875 26460 10876
tri 26460 10875 26462 10876 sw
tri 26168 10874 26189 10875 ne
rect 26189 10874 26232 10875
tri 26232 10874 26253 10875 nw
tri 26447 10874 26448 10875 se
rect 26448 10874 26462 10875
tri 26462 10874 26463 10875 sw
tri 26445 10873 26447 10874 se
rect 26447 10873 26463 10874
tri 26463 10873 26465 10874 sw
tri 26441 10868 26445 10873 se
rect 26445 10868 26465 10873
tri 26465 10868 26469 10873 sw
tri 26436 10860 26441 10868 se
rect 26441 10860 26469 10868
tri 26469 10860 26474 10868 sw
tri 26432 10851 26436 10860 se
rect 26436 10851 26474 10860
tri 26474 10851 26478 10860 sw
tri 26428 10840 26432 10851 se
rect 26432 10840 26478 10851
tri 26478 10840 26482 10851 sw
tri 26424 10827 26428 10840 se
rect 26428 10827 26482 10840
tri 26482 10827 26486 10840 sw
tri 26420 10813 26424 10827 se
rect 26424 10813 26486 10827
tri 26486 10813 26490 10827 sw
tri 26417 10797 26420 10813 se
rect 26420 10797 26490 10813
tri 26490 10797 26493 10813 sw
tri 26414 10780 26417 10797 se
rect 26417 10780 26493 10797
tri 26493 10780 26496 10797 sw
tri 26412 10761 26414 10780 se
rect 26414 10761 26496 10780
tri 26496 10761 26498 10780 sw
tri 26410 10742 26412 10761 se
rect 26412 10742 26498 10761
tri 26498 10742 26500 10761 sw
tri 26408 10722 26410 10742 se
rect 26410 10722 26500 10742
tri 26500 10722 26502 10742 sw
tri 26407 10701 26408 10722 se
rect 26408 10701 26502 10722
tri 26502 10701 26503 10722 sw
tri 26406 10680 26407 10701 se
rect 26407 10680 26503 10701
tri 26503 10680 26504 10701 sw
rect 26406 10637 26504 10680
tri 26406 10616 26407 10637 ne
rect 26407 10616 26503 10637
tri 26503 10616 26504 10637 nw
tri 25623 10615 25646 10616 se
tri 25646 10615 25669 10616 sw
tri 25600 10614 25623 10615 se
rect 25623 10614 25669 10615
tri 25669 10614 25692 10615 sw
tri 25578 10613 25600 10614 se
rect 25600 10613 25692 10614
tri 25692 10613 25714 10614 sw
tri 25556 10610 25578 10613 se
rect 25578 10610 25714 10613
tri 25714 10610 25736 10613 sw
tri 25535 10607 25556 10610 se
rect 25556 10607 25736 10610
tri 25736 10607 25757 10610 sw
rect 26407 10607 26502 10616
tri 25515 10603 25535 10607 se
rect 25535 10603 25757 10607
tri 25757 10603 25776 10607 sw
tri 26407 10605 26408 10607 ne
tri 25497 10599 25515 10603 se
rect 25515 10599 25776 10603
tri 25776 10599 25795 10603 sw
tri 25480 10594 25497 10599 se
rect 25497 10594 25795 10599
tri 25795 10594 25812 10599 sw
rect 26408 10595 26502 10607
tri 26502 10595 26503 10616 nw
rect 26408 10594 26500 10595
tri 25464 10588 25480 10594 se
rect 25480 10588 25812 10594
tri 25812 10588 25827 10594 sw
tri 26408 10590 26409 10594 ne
tri 25450 10582 25464 10588 se
rect 25464 10582 25827 10588
tri 25827 10582 25841 10588 sw
rect 26409 10582 26500 10594
tri 25439 10576 25450 10582 se
rect 25450 10576 25841 10582
tri 25841 10576 25853 10582 sw
tri 26409 10577 26410 10582 ne
tri 25429 10570 25439 10576 se
rect 25439 10570 25853 10576
tri 25853 10570 25863 10576 sw
rect 26410 10575 26500 10582
tri 26500 10575 26502 10595 nw
rect 26410 10570 26498 10575
tri 25421 10563 25429 10570 se
rect 25429 10563 25863 10570
tri 25863 10563 25871 10570 sw
tri 26410 10563 26411 10570 ne
rect 26411 10563 26498 10570
tri 25415 10555 25421 10563 se
rect 25421 10555 25871 10563
tri 25871 10555 25876 10563 sw
tri 26411 10555 26412 10563 ne
rect 26412 10555 26498 10563
tri 26498 10555 26500 10575 nw
tri 25412 10548 25415 10555 se
rect 25415 10548 25876 10555
tri 25876 10548 25880 10555 sw
tri 26412 10549 26413 10555 ne
rect 26413 10548 26496 10555
tri 25411 10541 25412 10548 se
tri 25411 10533 25412 10541 ne
rect 25412 10533 25880 10548
tri 25880 10541 25881 10548 sw
tri 25880 10533 25881 10541 nw
tri 26413 10537 26414 10548 ne
rect 26414 10537 26496 10548
tri 26496 10537 26498 10555 nw
tri 26414 10533 26415 10537 ne
rect 26415 10533 26493 10537
tri 25412 10526 25415 10533 ne
rect 25415 10526 25876 10533
tri 25876 10526 25880 10533 nw
tri 26415 10527 26416 10533 ne
rect 26416 10526 26493 10533
tri 25415 10519 25421 10526 ne
rect 25421 10519 25871 10526
tri 25871 10519 25876 10526 nw
tri 26416 10520 26417 10526 ne
rect 26417 10520 26493 10526
tri 26493 10520 26496 10537 nw
rect 26417 10519 26490 10520
tri 25421 10512 25429 10519 ne
rect 25429 10512 25863 10519
tri 25863 10512 25871 10519 nw
tri 26417 10513 26419 10519 ne
rect 26419 10512 26490 10519
tri 25429 10505 25439 10512 ne
rect 25439 10505 25853 10512
tri 25853 10505 25863 10512 nw
tri 26419 10506 26420 10512 ne
tri 25439 10499 25450 10505 ne
rect 25450 10499 25841 10505
tri 25841 10499 25853 10505 nw
rect 26420 10504 26490 10512
tri 26490 10504 26493 10520 nw
tri 26420 10500 26421 10504 ne
rect 26421 10499 26486 10504
tri 25450 10493 25464 10499 ne
rect 25464 10493 25827 10499
tri 25827 10493 25841 10499 nw
tri 26421 10493 26423 10499 ne
rect 26423 10493 26486 10499
tri 25464 10488 25480 10493 ne
rect 25480 10488 25812 10493
tri 25812 10488 25827 10493 nw
tri 26423 10489 26424 10493 ne
rect 26424 10489 26486 10493
tri 26486 10489 26490 10504 nw
rect 26424 10488 26482 10489
tri 25480 10483 25497 10488 ne
rect 25497 10483 25795 10488
tri 25795 10483 25812 10488 nw
tri 26424 10483 26426 10488 ne
rect 26426 10483 26482 10488
tri 25497 10478 25515 10483 ne
rect 25515 10478 25776 10483
tri 25776 10478 25795 10483 nw
tri 26426 10479 26427 10483 ne
rect 26427 10478 26482 10483
tri 25515 10475 25535 10478 ne
rect 25535 10475 25757 10478
tri 25757 10475 25776 10478 nw
tri 26427 10477 26428 10478 ne
rect 26428 10477 26482 10478
tri 26482 10477 26486 10489 nw
rect 26428 10475 26478 10477
tri 25535 10472 25556 10475 ne
rect 25556 10472 25736 10475
tri 25736 10472 25757 10475 nw
tri 26428 10472 26430 10475 ne
rect 26430 10472 26478 10475
tri 25556 10469 25578 10472 ne
rect 25578 10469 25714 10472
tri 25714 10469 25736 10472 nw
tri 26430 10469 26431 10472 ne
tri 25578 10467 25600 10469 ne
rect 25600 10467 25692 10469
tri 25692 10467 25714 10469 nw
rect 26431 10467 26478 10472
tri 25600 10466 25623 10467 ne
rect 25623 10466 25669 10467
tri 25669 10466 25692 10467 nw
rect 26432 10466 26478 10467
tri 26478 10466 26482 10477 nw
tri 26432 10456 26436 10466 ne
rect 26436 10456 26474 10466
tri 26474 10456 26478 10466 nw
tri 26436 10449 26441 10456 ne
rect 26441 10449 26469 10456
tri 26469 10449 26474 10456 nw
tri 26441 10444 26445 10449 ne
rect 26445 10444 26465 10449
tri 26465 10444 26469 10449 nw
tri 26445 10441 26450 10444 ne
rect 26450 10441 26460 10444
tri 26460 10441 26465 10444 nw
tri 26450 10440 26455 10441 ne
tri 26455 10440 26460 10441 nw
tri 25503 10209 25522 10210 se
rect 25522 10209 25561 10210
tri 25561 10209 25580 10210 sw
tri 25484 10208 25503 10209 se
rect 25503 10208 25580 10209
tri 25580 10208 25599 10209 sw
tri 25466 10207 25484 10208 se
rect 25484 10207 25599 10208
tri 25599 10207 25617 10208 sw
tri 25448 10205 25466 10207 se
rect 25466 10205 25617 10207
tri 25617 10205 25635 10207 sw
tri 25432 10203 25448 10205 se
rect 25448 10203 25635 10205
tri 25635 10203 25651 10205 sw
tri 25416 10201 25432 10203 se
rect 25432 10201 25651 10203
tri 25651 10201 25667 10203 sw
tri 25402 10198 25416 10201 se
rect 25416 10198 25667 10201
tri 25667 10198 25681 10201 sw
tri 25389 10195 25402 10198 se
rect 25402 10195 25681 10198
tri 25681 10195 25694 10198 sw
tri 25377 10192 25389 10195 se
rect 25389 10192 25694 10195
tri 25694 10192 25706 10195 sw
tri 25367 10188 25377 10192 se
rect 25377 10188 25706 10192
tri 25706 10188 25716 10192 sw
tri 25359 10184 25367 10188 se
rect 25367 10184 25716 10188
tri 25716 10184 25724 10188 sw
tri 25353 10180 25359 10184 se
rect 25359 10180 25724 10184
tri 25724 10180 25731 10184 sw
tri 25348 10177 25353 10180 se
rect 25353 10177 25731 10180
tri 25731 10177 25735 10180 sw
tri 25345 10172 25348 10177 se
rect 25348 10172 25735 10177
tri 25735 10172 25738 10177 sw
tri 25344 10168 25345 10172 se
tri 25344 10164 25345 10168 ne
rect 25345 10164 25738 10172
tri 25738 10168 25739 10172 sw
tri 25738 10164 25739 10168 nw
tri 25345 10160 25348 10164 ne
rect 25348 10160 25735 10164
tri 25735 10160 25738 10164 nw
tri 25348 10156 25353 10160 ne
rect 25353 10156 25731 10160
tri 25731 10156 25735 10160 nw
tri 25353 10152 25359 10156 ne
rect 25359 10152 25724 10156
tri 25724 10152 25731 10156 nw
tri 25359 10149 25367 10152 ne
rect 25367 10149 25716 10152
tri 25716 10149 25724 10152 nw
tri 25367 10145 25377 10149 ne
rect 25377 10145 25706 10149
tri 25706 10145 25716 10149 nw
tri 25377 10142 25389 10145 ne
rect 25389 10142 25694 10145
tri 25694 10142 25706 10145 nw
tri 25389 10139 25402 10142 ne
rect 25402 10139 25681 10142
tri 25681 10139 25694 10142 nw
tri 25402 10136 25416 10139 ne
rect 25416 10136 25667 10139
tri 25667 10136 25681 10139 nw
tri 25416 10134 25432 10136 ne
rect 25432 10134 25651 10136
tri 25651 10134 25667 10136 nw
tri 25432 10132 25448 10134 ne
rect 25448 10132 25635 10134
tri 25635 10132 25651 10134 nw
tri 25448 10130 25466 10132 ne
rect 25466 10130 25617 10132
tri 25617 10130 25635 10132 nw
tri 25466 10129 25484 10130 ne
rect 25484 10129 25599 10130
tri 25599 10129 25617 10130 nw
tri 25484 10128 25503 10129 ne
rect 25503 10128 25580 10129
tri 25580 10128 25599 10129 nw
tri 25503 10127 25522 10128 ne
rect 25522 10127 25561 10128
tri 25561 10127 25580 10128 nw
tri 20509 8651 20533 8652 se
rect 20533 8651 20582 8652
tri 20582 8651 20607 8652 sw
tri 20485 8649 20509 8651 se
rect 20509 8649 20607 8651
tri 20607 8649 20630 8651 sw
tri 20462 8647 20485 8649 se
rect 20485 8647 20630 8649
tri 20630 8647 20654 8649 sw
tri 20440 8644 20462 8647 se
rect 20462 8644 20654 8647
tri 20654 8644 20676 8647 sw
tri 20419 8640 20440 8644 se
rect 20440 8640 20676 8644
tri 20676 8640 20697 8644 sw
tri 20399 8636 20419 8640 se
rect 20419 8636 20697 8640
tri 20697 8636 20717 8640 sw
tri 20381 8631 20399 8636 se
rect 20399 8631 20717 8636
tri 20717 8631 20735 8636 sw
tri 20364 8626 20381 8631 se
rect 20381 8626 20735 8631
tri 20735 8626 20751 8631 sw
tri 20350 8620 20364 8626 se
rect 20364 8620 20751 8626
tri 20751 8620 20766 8626 sw
tri 20337 8614 20350 8620 se
rect 20350 8614 20766 8620
tri 20766 8614 20778 8620 sw
tri 20327 8608 20337 8614 se
rect 20337 8608 20778 8614
tri 20778 8608 20789 8614 sw
tri 20318 8601 20327 8608 se
rect 20327 8601 20789 8608
tri 20789 8601 20797 8608 sw
tri 20312 8594 20318 8601 se
rect 20318 8594 20797 8601
tri 20797 8594 20803 8601 sw
tri 20309 8587 20312 8594 se
rect 20312 8587 20803 8594
tri 20803 8587 20807 8594 sw
tri 20308 8580 20309 8587 se
tri 20308 8573 20309 8580 ne
rect 20309 8573 20807 8587
tri 20807 8580 20808 8587 sw
tri 20807 8573 20808 8580 nw
tri 20309 8566 20312 8573 ne
rect 20312 8566 20803 8573
tri 20803 8566 20807 8573 nw
tri 20312 8560 20318 8566 ne
rect 20318 8560 20797 8566
tri 20797 8560 20803 8566 nw
tri 20318 8553 20327 8560 ne
rect 20327 8553 20789 8560
tri 20789 8553 20797 8560 nw
tri 20327 8547 20337 8553 ne
rect 20337 8547 20778 8553
tri 20778 8547 20789 8553 nw
tri 20337 8541 20350 8547 ne
rect 20350 8541 20766 8547
tri 20766 8541 20778 8547 nw
tri 20350 8535 20364 8541 ne
rect 20364 8535 20751 8541
tri 20751 8535 20766 8541 nw
tri 20364 8530 20381 8535 ne
rect 20381 8530 20735 8535
tri 20735 8530 20751 8535 nw
tri 20381 8525 20399 8530 ne
rect 20399 8525 20717 8530
tri 20717 8525 20735 8530 nw
tri 20399 8521 20419 8525 ne
rect 20419 8521 20697 8525
tri 20697 8521 20717 8525 nw
tri 20419 8517 20440 8521 ne
rect 20440 8517 20676 8521
tri 20676 8517 20697 8521 nw
tri 20440 8514 20462 8517 ne
rect 20462 8514 20654 8517
tri 20654 8514 20676 8517 nw
tri 20462 8512 20485 8514 ne
rect 20485 8512 20630 8514
tri 20630 8512 20654 8514 nw
tri 20485 8510 20509 8512 ne
rect 20509 8510 20607 8512
tri 20607 8510 20630 8512 nw
tri 20509 8509 20533 8510 ne
rect 20533 8509 20582 8510
tri 20582 8509 20607 8510 nw
tri 13371 5536 13386 5537 se
rect 13386 5536 13418 5537
tri 13418 5536 13433 5537 sw
tri 13340 5535 13355 5536 se
rect 13355 5535 13449 5536
tri 13449 5535 13464 5536 sw
tri 13326 5534 13340 5535 se
rect 13340 5534 13464 5535
tri 13464 5534 13478 5535 sw
tri 13313 5533 13326 5534 se
rect 13326 5533 13478 5534
tri 13478 5533 13491 5534 sw
tri 13300 5531 13313 5533 se
rect 13313 5531 13491 5533
tri 13491 5531 13504 5533 sw
tri 13288 5529 13300 5531 se
rect 13300 5529 13504 5531
tri 13504 5529 13516 5531 sw
tri 13278 5528 13288 5529 se
rect 13288 5528 13516 5529
tri 13516 5528 13526 5529 sw
tri 13268 5526 13278 5528 se
rect 13278 5526 13526 5528
tri 13526 5526 13536 5528 sw
tri 13260 5523 13268 5526 se
rect 13268 5523 13536 5526
tri 13536 5523 13544 5526 sw
tri 13253 5521 13260 5523 se
rect 13260 5521 13544 5523
tri 13544 5521 13551 5523 sw
tri 13248 5519 13253 5521 se
rect 13253 5519 13551 5521
tri 13551 5519 13556 5521 sw
tri 13244 5516 13248 5519 se
rect 13248 5516 13556 5519
tri 13556 5516 13560 5519 sw
tri 13242 5514 13244 5516 se
rect 13244 5514 13560 5516
tri 13560 5514 13562 5516 sw
tri 13241 5511 13242 5514 se
tri 13241 5509 13242 5511 ne
rect 13242 5509 13562 5514
tri 13562 5511 13563 5514 sw
tri 13562 5509 13563 5511 nw
tri 13242 5506 13244 5509 ne
rect 13244 5506 13560 5509
tri 13560 5506 13562 5509 nw
tri 13244 5504 13248 5506 ne
rect 13248 5504 13556 5506
tri 13556 5504 13560 5506 nw
tri 13248 5502 13253 5504 ne
rect 13253 5502 13551 5504
tri 13551 5502 13556 5504 nw
tri 13253 5499 13260 5502 ne
rect 13260 5499 13544 5502
tri 13544 5499 13551 5502 nw
tri 13260 5497 13268 5499 ne
rect 13268 5497 13536 5499
tri 13536 5497 13544 5499 nw
tri 13268 5495 13278 5497 ne
rect 13278 5495 13526 5497
tri 13526 5495 13536 5497 nw
tri 13278 5493 13288 5495 ne
rect 13288 5493 13516 5495
tri 13516 5493 13526 5495 nw
tri 13288 5492 13300 5493 ne
rect 13300 5492 13504 5493
tri 13504 5492 13516 5493 nw
tri 13300 5490 13313 5492 ne
rect 13313 5490 13491 5492
tri 13491 5490 13504 5492 nw
tri 13313 5489 13326 5490 ne
rect 13326 5489 13478 5490
tri 13478 5489 13491 5490 nw
tri 13326 5488 13340 5489 ne
rect 13340 5488 13464 5489
tri 13464 5488 13478 5489 nw
tri 13340 5487 13355 5488 ne
rect 13355 5487 13449 5488
tri 13449 5487 13464 5488 nw
tri 13355 5486 13371 5487 ne
rect 13371 5486 13433 5487
tri 13433 5486 13449 5487 nw
tri 13283 5469 13298 5470 se
rect 13298 5469 13330 5470
tri 13330 5469 13345 5470 sw
tri 13252 5468 13267 5469 se
rect 13267 5468 13361 5469
tri 13361 5468 13376 5469 sw
tri 13238 5467 13252 5468 se
rect 13252 5467 13376 5468
tri 13376 5467 13390 5468 sw
tri 13225 5466 13238 5467 se
rect 13238 5466 13390 5467
tri 13390 5466 13403 5467 sw
tri 13212 5464 13225 5466 se
rect 13225 5464 13403 5466
tri 13403 5464 13416 5466 sw
tri 13200 5462 13212 5464 se
rect 13212 5462 13416 5464
tri 13416 5462 13428 5464 sw
tri 13190 5461 13200 5462 se
rect 13200 5461 13428 5462
tri 13428 5461 13438 5462 sw
tri 13180 5459 13190 5461 se
rect 13190 5459 13438 5461
tri 13438 5459 13448 5461 sw
tri 13172 5456 13180 5459 se
rect 13180 5456 13448 5459
tri 13448 5456 13456 5459 sw
tri 13165 5454 13172 5456 se
rect 13172 5454 13456 5456
tri 13456 5454 13463 5456 sw
tri 13160 5452 13165 5454 se
rect 13165 5452 13463 5454
tri 13463 5452 13468 5454 sw
tri 13156 5449 13160 5452 se
rect 13160 5449 13468 5452
tri 13468 5449 13472 5452 sw
tri 13154 5447 13156 5449 se
rect 13156 5447 13472 5449
tri 13472 5447 13474 5449 sw
tri 13153 5444 13154 5447 se
tri 13153 5442 13154 5444 ne
rect 13154 5442 13474 5447
tri 13474 5444 13475 5447 sw
tri 13474 5442 13475 5444 nw
tri 13154 5439 13156 5442 ne
rect 13156 5439 13472 5442
tri 13472 5439 13474 5442 nw
tri 13156 5437 13160 5439 ne
rect 13160 5437 13468 5439
tri 13468 5437 13472 5439 nw
tri 13160 5435 13165 5437 ne
rect 13165 5435 13463 5437
tri 13463 5435 13468 5437 nw
tri 13165 5432 13172 5435 ne
rect 13172 5432 13456 5435
tri 13456 5432 13463 5435 nw
tri 13172 5430 13180 5432 ne
rect 13180 5430 13448 5432
tri 13448 5430 13456 5432 nw
tri 13180 5428 13190 5430 ne
rect 13190 5428 13438 5430
tri 13438 5428 13448 5430 nw
tri 13190 5426 13200 5428 ne
rect 13200 5426 13428 5428
tri 13428 5426 13438 5428 nw
tri 13200 5425 13212 5426 ne
rect 13212 5425 13416 5426
tri 13416 5425 13428 5426 nw
tri 13212 5423 13225 5425 ne
rect 13225 5423 13403 5425
tri 13403 5423 13416 5425 nw
tri 13225 5422 13238 5423 ne
rect 13238 5422 13390 5423
tri 13390 5422 13403 5423 nw
tri 13238 5421 13252 5422 ne
rect 13252 5421 13376 5422
tri 13376 5421 13390 5422 nw
tri 13252 5420 13267 5421 ne
rect 13267 5420 13361 5421
tri 13361 5420 13376 5421 nw
tri 13267 5419 13283 5420 ne
rect 13283 5419 13345 5420
tri 13345 5419 13361 5420 nw
tri 14981 4925 14989 4926 se
tri 14989 4925 14997 4926 sw
tri 15190 4925 15198 4926 se
tri 15198 4925 15206 4926 sw
tri 14972 4922 14981 4925 se
rect 14981 4922 14997 4925
tri 14997 4922 15006 4925 sw
tri 15181 4922 15190 4925 se
rect 15190 4922 15206 4925
tri 15206 4922 15215 4925 sw
tri 14964 4916 14972 4922 se
rect 14972 4916 15006 4922
tri 15006 4916 15014 4922 sw
tri 15173 4916 15181 4922 se
rect 15181 4916 15215 4922
tri 15215 4916 15223 4922 sw
tri 14956 4908 14964 4916 se
rect 14964 4908 15014 4916
tri 15014 4908 15022 4916 sw
tri 15165 4908 15173 4916 se
rect 15173 4908 15223 4916
tri 15223 4908 15231 4916 sw
tri 14949 4899 14956 4908 se
rect 14956 4899 15022 4908
tri 15022 4899 15029 4908 sw
tri 15158 4899 15165 4908 se
rect 15165 4899 15231 4908
tri 15231 4899 15238 4908 sw
tri 14942 4887 14949 4899 se
rect 14949 4887 15029 4899
tri 15029 4887 15036 4899 sw
tri 15151 4887 15158 4899 se
rect 15158 4887 15238 4899
tri 15238 4887 15245 4899 sw
tri 14935 4873 14942 4887 se
rect 14942 4873 15036 4887
tri 15036 4873 15043 4887 sw
tri 15144 4873 15151 4887 se
rect 15151 4873 15245 4887
tri 15245 4873 15252 4887 sw
tri 14929 4858 14935 4873 se
rect 14935 4858 15043 4873
tri 15043 4858 15049 4873 sw
tri 15138 4858 15144 4873 se
rect 15144 4858 15252 4873
tri 15252 4858 15258 4873 sw
tri 14923 4841 14929 4858 se
rect 14929 4841 15049 4858
tri 15049 4841 15055 4858 sw
tri 15132 4841 15138 4858 se
rect 15138 4841 15258 4858
tri 15258 4841 15264 4858 sw
tri 14918 4823 14923 4841 se
rect 14923 4823 15055 4841
tri 15055 4823 15060 4841 sw
tri 15127 4823 15132 4841 se
rect 15132 4823 15264 4841
tri 15264 4823 15269 4841 sw
tri 14914 4803 14918 4823 se
rect 14918 4803 15060 4823
tri 15060 4803 15064 4823 sw
tri 15123 4803 15127 4823 se
rect 15127 4803 15269 4823
tri 15269 4803 15273 4823 sw
tri 14910 4782 14914 4803 se
rect 14914 4782 15064 4803
tri 15064 4782 15068 4803 sw
tri 15119 4782 15123 4803 se
rect 15123 4782 15273 4803
tri 15273 4782 15277 4803 sw
tri 14907 4761 14910 4782 se
rect 14910 4761 15068 4782
tri 15068 4761 15071 4782 sw
tri 15116 4761 15119 4782 se
rect 15119 4761 15277 4782
tri 15277 4761 15280 4782 sw
tri 14905 4739 14907 4761 se
rect 14907 4739 15071 4761
tri 15071 4739 15073 4761 sw
tri 15114 4739 15116 4761 se
rect 15116 4739 15280 4761
tri 15280 4739 15282 4761 sw
tri 14904 4716 14905 4739 se
rect 14905 4716 15073 4739
tri 15073 4716 15074 4739 sw
rect 14904 4671 15074 4716
tri 14904 4648 14905 4671 ne
rect 14905 4648 15073 4671
tri 15073 4648 15074 4671 nw
tri 15113 4716 15114 4739 se
rect 15114 4716 15282 4739
tri 15282 4716 15283 4739 sw
rect 15113 4671 15283 4716
tri 15113 4648 15114 4671 ne
rect 15114 4648 15282 4671
tri 15282 4648 15283 4671 nw
tri 14905 4626 14907 4648 ne
rect 14907 4626 15071 4648
tri 15071 4626 15073 4648 nw
tri 15114 4626 15116 4648 ne
rect 15116 4626 15280 4648
tri 15280 4626 15282 4648 nw
tri 14907 4604 14910 4626 ne
rect 14910 4604 15068 4626
tri 15068 4604 15071 4626 nw
tri 15116 4604 15119 4626 ne
rect 15119 4604 15277 4626
tri 15277 4604 15280 4626 nw
tri 14910 4584 14914 4604 ne
rect 14914 4584 15064 4604
tri 15064 4584 15068 4604 nw
tri 15119 4584 15123 4604 ne
rect 15123 4584 15273 4604
tri 15273 4584 15277 4604 nw
tri 14914 4564 14918 4584 ne
rect 14918 4564 15060 4584
tri 15060 4564 15064 4584 nw
tri 15123 4564 15127 4584 ne
rect 15127 4564 15269 4584
tri 15269 4564 15273 4584 nw
tri 14918 4546 14923 4564 ne
rect 14923 4546 15055 4564
tri 15055 4546 15060 4564 nw
tri 15127 4546 15132 4564 ne
rect 15132 4546 15264 4564
tri 15264 4546 15269 4564 nw
tri 14923 4529 14929 4546 ne
rect 14929 4529 15049 4546
tri 15049 4529 15055 4546 nw
tri 15132 4529 15138 4546 ne
rect 15138 4529 15258 4546
tri 15258 4529 15264 4546 nw
tri 14929 4513 14935 4529 ne
rect 14935 4513 15043 4529
tri 15043 4513 15049 4529 nw
tri 15138 4513 15144 4529 ne
rect 15144 4513 15252 4529
tri 15252 4513 15258 4529 nw
tri 14935 4500 14942 4513 ne
rect 14942 4500 15036 4513
tri 15036 4500 15043 4513 nw
tri 15144 4500 15151 4513 ne
rect 15151 4500 15245 4513
tri 15245 4500 15252 4513 nw
tri 14942 4488 14949 4500 ne
rect 14949 4488 15029 4500
tri 15029 4488 15036 4500 nw
tri 15151 4488 15158 4500 ne
rect 15158 4488 15238 4500
tri 15238 4488 15245 4500 nw
tri 14949 4478 14956 4488 ne
rect 14956 4478 15022 4488
tri 15022 4478 15029 4488 nw
tri 15158 4478 15165 4488 ne
rect 15165 4478 15231 4488
tri 15231 4478 15238 4488 nw
tri 14956 4471 14964 4478 ne
rect 14964 4471 15014 4478
tri 15014 4471 15022 4478 nw
tri 15165 4471 15173 4478 ne
rect 15173 4471 15223 4478
tri 15223 4471 15231 4478 nw
tri 14964 4465 14972 4471 ne
rect 14972 4465 15006 4471
tri 15006 4465 15014 4471 nw
tri 15173 4465 15181 4471 ne
rect 15181 4465 15215 4471
tri 15215 4465 15223 4471 nw
tri 14972 4462 14981 4465 ne
rect 14981 4462 14997 4465
tri 14997 4462 15006 4465 nw
tri 15181 4462 15190 4465 ne
rect 15190 4462 15206 4465
tri 15206 4462 15215 4465 nw
tri 14981 4461 14989 4462 ne
tri 14989 4461 14997 4462 nw
tri 15190 4461 15198 4462 ne
tri 15198 4461 15206 4462 nw
tri 20046 3538 20051 3540 se
tri 20051 3538 20056 3540 sw
tri 20041 3532 20046 3538 se
rect 20046 3532 20056 3538
tri 20056 3532 20061 3538 sw
tri 20036 3523 20041 3532 se
rect 20041 3523 20061 3532
tri 20061 3523 20066 3532 sw
tri 20032 3510 20036 3523 se
rect 20036 3510 20066 3523
tri 20066 3510 20070 3523 sw
tri 20027 3494 20032 3510 se
rect 20032 3494 20070 3510
tri 20070 3494 20075 3510 sw
tri 20023 3475 20027 3494 se
rect 20027 3475 20075 3494
tri 20075 3475 20079 3494 sw
tri 20019 3452 20023 3475 se
rect 20023 3452 20079 3475
tri 20079 3452 20083 3475 sw
tri 20016 3427 20019 3452 se
rect 20019 3427 20083 3452
tri 20083 3427 20086 3452 sw
tri 20012 3399 20016 3427 se
rect 20016 3399 20086 3427
tri 20086 3399 20090 3427 sw
tri 20009 3369 20012 3399 se
rect 20012 3369 20090 3399
tri 20090 3369 20093 3399 sw
tri 20007 3336 20009 3369 se
rect 20009 3336 20093 3369
tri 20093 3336 20095 3369 sw
tri 20005 3302 20007 3336 se
rect 20007 3302 20095 3336
tri 20095 3302 20097 3336 sw
tri 20003 3266 20005 3302 se
rect 20005 3266 20097 3302
tri 20097 3266 20099 3302 sw
tri 20002 3230 20003 3266 se
rect 20003 3230 20099 3266
tri 20099 3230 20100 3266 sw
tri 20001 3192 20002 3230 se
rect 20002 3192 20100 3230
tri 20100 3192 20101 3230 sw
tri 13336 3160 13343 3162 se
tri 13343 3160 13349 3162 sw
tri 13330 3153 13336 3160 se
rect 13336 3153 13349 3160
tri 13349 3153 13356 3160 sw
tri 13324 3142 13330 3153 se
rect 13330 3142 13356 3153
tri 13356 3142 13362 3153 sw
tri 13318 3126 13324 3142 se
rect 13324 3126 13362 3142
tri 13362 3126 13368 3142 sw
tri 13312 3107 13318 3126 se
rect 13318 3107 13368 3126
tri 13368 3107 13374 3126 sw
rect 20001 3117 20101 3192
rect 20001 3107 20100 3117
tri 13307 3083 13312 3107 se
rect 13312 3083 13374 3107
tri 13374 3083 13379 3107 sw
tri 20001 3088 20002 3107 ne
tri 13301 3056 13307 3083 se
rect 13307 3056 13379 3083
tri 13379 3056 13384 3083 sw
rect 20002 3079 20100 3107
tri 20100 3079 20101 3117 nw
tri 20002 3061 20003 3079 ne
tri 13297 3025 13301 3056 se
rect 13301 3025 13384 3056
tri 13384 3025 13389 3056 sw
rect 20003 3043 20099 3079
tri 20099 3043 20100 3079 nw
tri 20003 3025 20004 3043 ne
rect 20004 3025 20097 3043
tri 13292 2990 13297 3025 se
rect 13297 2990 13389 3025
tri 13389 2990 13393 3025 sw
tri 20004 3007 20005 3025 ne
rect 20005 3007 20097 3025
tri 20097 3007 20099 3043 nw
tri 20005 2991 20006 3007 ne
rect 20006 2990 20095 3007
tri 13289 2953 13292 2990 se
rect 13292 2957 13393 2990
tri 13393 2957 13397 2990 sw
tri 20006 2973 20007 2990 ne
rect 20007 2973 20095 2990
tri 20095 2973 20097 3007 nw
tri 20007 2959 20008 2973 ne
rect 13292 2953 13397 2957
tri 13483 2955 13490 2957 se
tri 13490 2955 13496 2957 sw
rect 20008 2955 20093 2973
tri 13482 2953 13483 2955 se
rect 13483 2953 13496 2955
tri 13285 2914 13289 2953 se
rect 13289 2939 13397 2953
tri 13477 2948 13482 2953 se
rect 13482 2948 13496 2953
tri 13496 2948 13503 2955 sw
tri 20008 2951 20009 2955 ne
tri 13397 2939 13398 2948 sw
rect 13289 2923 13398 2939
tri 13471 2937 13477 2948 se
rect 13477 2937 13503 2948
tri 13503 2937 13509 2948 sw
rect 20009 2940 20093 2955
tri 20093 2940 20095 2973 nw
tri 20009 2938 20010 2940 ne
rect 20010 2937 20090 2940
tri 13398 2923 13400 2937 sw
rect 13289 2914 13400 2923
tri 13465 2922 13471 2937 se
rect 13471 2922 13509 2937
tri 13509 2922 13515 2937 sw
tri 20010 2922 20011 2937 ne
rect 20011 2922 20090 2937
tri 13462 2914 13465 2922 se
rect 13465 2914 13515 2922
tri 13283 2872 13285 2914 se
rect 13285 2904 13400 2914
tri 13400 2904 13401 2914 sw
rect 13285 2882 13401 2904
tri 13459 2903 13462 2914 se
rect 13462 2903 13515 2914
tri 13515 2903 13521 2922 sw
tri 20011 2910 20012 2922 ne
rect 20012 2910 20090 2922
tri 20090 2910 20093 2940 nw
tri 20012 2903 20013 2910 ne
rect 20013 2903 20086 2910
tri 13401 2882 13402 2903 sw
rect 13285 2872 13402 2882
tri 13454 2879 13459 2903 se
rect 13459 2879 13521 2903
tri 13521 2879 13526 2903 sw
tri 20013 2882 20016 2903 ne
rect 20016 2882 20086 2903
tri 20086 2882 20090 2910 nw
rect 20016 2879 20083 2882
tri 13402 2872 13403 2879 sw
tri 13452 2872 13454 2879 se
rect 13454 2872 13526 2879
tri 13280 2829 13283 2872 se
rect 13283 2852 13403 2872
tri 13403 2852 13404 2872 sw
tri 13448 2852 13452 2872 se
rect 13452 2852 13526 2872
tri 13526 2852 13531 2879 sw
tri 20016 2856 20019 2879 ne
rect 20019 2856 20083 2879
tri 20083 2856 20086 2882 nw
tri 20019 2853 20020 2856 ne
rect 20020 2852 20079 2856
rect 13283 2829 13404 2852
tri 13404 2829 13405 2852 sw
tri 13279 2784 13280 2829 se
rect 13280 2790 13405 2829
tri 13445 2829 13448 2852 se
rect 13448 2829 13531 2852
tri 13444 2822 13445 2828 se
rect 13445 2822 13531 2829
tri 13531 2822 13536 2852 sw
tri 20020 2834 20023 2852 ne
rect 20023 2834 20079 2852
tri 20079 2834 20083 2856 nw
tri 20023 2823 20026 2834 ne
rect 20026 2822 20075 2834
tri 13405 2790 13407 2822 sw
rect 13280 2784 13407 2790
tri 13439 2788 13444 2822 se
rect 13444 2788 13536 2822
tri 13536 2788 13540 2822 sw
tri 20026 2815 20027 2822 ne
rect 20027 2815 20075 2822
tri 20075 2815 20079 2834 nw
tri 20027 2798 20032 2815 ne
rect 20032 2798 20070 2815
tri 20070 2798 20075 2815 nw
tri 20032 2789 20035 2798 ne
rect 20035 2788 20066 2798
tri 13278 2738 13279 2784 se
rect 13279 2738 13407 2784
tri 13436 2752 13439 2784 se
rect 13439 2752 13540 2788
tri 13540 2752 13544 2788 sw
tri 20035 2786 20036 2788 ne
rect 20036 2786 20066 2788
tri 20066 2786 20070 2798 nw
tri 20036 2776 20041 2786 ne
rect 20041 2776 20061 2786
tri 20061 2776 20066 2786 nw
tri 20041 2771 20046 2776 ne
rect 20046 2771 20056 2776
tri 20056 2771 20061 2776 nw
tri 20046 2769 20051 2771 ne
tri 20051 2769 20056 2771 nw
tri 13407 2738 13408 2752 sw
tri 13434 2738 13436 2752 se
rect 13436 2738 13544 2752
rect 13278 2646 13408 2738
tri 13432 2713 13434 2738 se
rect 13434 2713 13544 2738
tri 13544 2713 13547 2752 sw
tri 13430 2672 13432 2713 se
rect 13432 2672 13547 2713
tri 13547 2672 13550 2713 sw
tri 17373 2680 17401 2682 se
rect 17401 2680 17458 2682
tri 17458 2680 17486 2682 sw
tri 17346 2678 17373 2680 se
rect 17373 2678 17486 2680
tri 17486 2678 17514 2680 sw
tri 17319 2675 17346 2678 se
rect 17346 2675 17514 2678
tri 17514 2675 17540 2678 sw
tri 17304 2672 17319 2675 se
rect 17319 2672 17540 2675
tri 17540 2672 17556 2675 sw
rect 13278 2629 13407 2646
tri 13407 2635 13408 2646 nw
tri 13428 2646 13430 2672 se
rect 13430 2646 13550 2672
tri 13427 2629 13428 2633 se
rect 13428 2629 13550 2646
tri 13550 2629 13552 2672 sw
tri 17293 2671 17304 2672 se
rect 17304 2671 17556 2672
tri 17556 2671 17566 2672 sw
tri 17269 2666 17293 2671 se
rect 17293 2666 17566 2671
tri 17566 2666 17590 2671 sw
tri 17246 2660 17269 2666 se
rect 17269 2660 17590 2666
tri 17590 2660 17613 2666 sw
tri 17225 2654 17246 2660 se
rect 17246 2654 17613 2660
tri 17613 2654 17634 2660 sw
tri 17206 2647 17225 2654 se
rect 17225 2647 17634 2654
tri 17634 2647 17653 2654 sw
tri 17189 2639 17206 2647 se
rect 17206 2639 17653 2647
tri 17653 2639 17670 2647 sw
tri 17175 2631 17189 2639 se
rect 17189 2631 17670 2639
tri 17670 2631 17685 2639 sw
tri 17172 2629 17175 2631 se
rect 17175 2629 17685 2631
tri 17685 2629 17687 2631 sw
tri 13278 2601 13279 2629 ne
rect 13279 2601 13407 2629
rect 13279 2585 13406 2601
tri 13406 2585 13407 2601 nw
tri 13426 2602 13427 2629 se
rect 13427 2602 13552 2629
rect 13426 2585 13552 2602
tri 13552 2585 13554 2629 sw
tri 17163 2623 17172 2629 se
rect 17172 2623 17687 2629
tri 17687 2623 17697 2629 sw
tri 17153 2614 17163 2623 se
rect 17163 2614 17697 2623
tri 17697 2614 17707 2623 sw
tri 17146 2605 17153 2614 se
rect 17153 2605 17707 2614
tri 17707 2605 17713 2614 sw
tri 17142 2595 17146 2605 se
rect 17146 2595 17713 2605
tri 17713 2595 17718 2605 sw
tri 17141 2586 17142 2595 se
rect 17142 2586 17718 2595
tri 17718 2586 17719 2595 sw
rect 17141 2585 17718 2586
tri 13279 2556 13280 2585 ne
rect 13280 2584 13406 2585
rect 13280 2556 13405 2584
tri 13405 2556 13406 2584 nw
tri 13425 2556 13426 2585 se
rect 13426 2556 13554 2585
tri 13280 2544 13281 2556 ne
rect 13281 2541 13404 2556
tri 13404 2541 13405 2556 nw
rect 13425 2541 13554 2556
tri 13554 2541 13555 2585 sw
tri 17141 2576 17142 2585 ne
rect 17142 2576 17718 2585
tri 17718 2576 17719 2586 nw
tri 17142 2567 17146 2576 ne
rect 17146 2567 17713 2576
tri 17713 2567 17718 2576 nw
tri 17146 2558 17153 2567 ne
rect 17153 2558 17707 2567
tri 17707 2558 17713 2567 nw
tri 17153 2549 17163 2558 ne
rect 17163 2549 17697 2558
tri 17697 2549 17707 2558 nw
tri 17163 2541 17174 2549 ne
rect 17174 2541 17685 2549
tri 13281 2513 13283 2541 ne
rect 13283 2540 13404 2541
rect 13283 2513 13403 2540
tri 13403 2513 13404 2540 nw
tri 13283 2471 13285 2513 ne
rect 13285 2471 13400 2513
tri 13400 2471 13403 2513 nw
tri 13285 2452 13287 2471 ne
rect 13287 2450 13399 2471
tri 13399 2450 13400 2471 nw
rect 13425 2450 13555 2541
tri 17174 2540 17175 2541 ne
rect 17175 2540 17685 2541
tri 17685 2540 17697 2549 nw
tri 17175 2532 17189 2540 ne
rect 17189 2532 17670 2540
tri 17670 2532 17685 2540 nw
tri 17189 2525 17206 2532 ne
rect 17206 2525 17653 2532
tri 17653 2525 17670 2532 nw
tri 17206 2518 17225 2525 ne
rect 17225 2518 17634 2525
tri 17634 2518 17653 2525 nw
tri 17225 2511 17246 2518 ne
rect 17246 2511 17613 2518
tri 17613 2511 17634 2518 nw
tri 17246 2506 17269 2511 ne
rect 17269 2506 17590 2511
tri 17590 2506 17613 2511 nw
tri 17269 2501 17293 2506 ne
rect 17293 2501 17566 2506
tri 17566 2501 17590 2506 nw
tri 17293 2497 17319 2501 ne
rect 17319 2497 17540 2501
tri 17540 2497 17566 2501 nw
tri 17319 2494 17346 2497 ne
rect 17346 2494 17514 2497
tri 17514 2494 17540 2497 nw
tri 17346 2491 17373 2494 ne
rect 17373 2491 17486 2494
tri 17486 2491 17514 2494 nw
tri 17373 2490 17401 2491 ne
rect 17401 2490 17458 2491
tri 17458 2490 17486 2491 nw
tri 13287 2431 13289 2450 ne
rect 13289 2431 13397 2450
tri 13397 2431 13399 2450 nw
rect 13425 2431 13554 2450
tri 13289 2406 13291 2431 ne
rect 13291 2405 13394 2431
tri 13394 2406 13397 2431 nw
tri 13425 2417 13426 2431 ne
tri 13291 2394 13292 2405 ne
rect 13292 2394 13393 2405
tri 13393 2394 13394 2405 nw
rect 13426 2405 13554 2431
tri 13554 2405 13555 2450 nw
rect 13426 2394 13552 2405
tri 13292 2362 13296 2394 ne
rect 13296 2361 13389 2394
tri 13389 2362 13393 2394 nw
tri 13426 2367 13427 2394 ne
tri 13296 2360 13297 2361 ne
rect 13297 2360 13389 2361
tri 13297 2329 13301 2360 ne
rect 13301 2329 13384 2360
tri 13384 2329 13389 2360 nw
rect 13427 2361 13552 2394
tri 13552 2361 13554 2405 nw
rect 13427 2360 13550 2361
tri 13427 2330 13429 2360 ne
rect 13429 2329 13550 2360
tri 13301 2319 13303 2329 ne
rect 13303 2319 13382 2329
tri 13382 2319 13384 2329 nw
tri 13429 2319 13430 2329 ne
rect 13430 2319 13550 2329
tri 13550 2319 13552 2361 nw
tri 13303 2302 13307 2319 ne
rect 13307 2302 13379 2319
tri 13379 2302 13382 2319 nw
tri 13430 2303 13431 2319 ne
rect 13431 2302 13547 2319
tri 13307 2278 13312 2302 ne
rect 13312 2278 13374 2302
tri 13374 2278 13379 2302 nw
tri 13431 2281 13432 2302 ne
rect 13432 2278 13547 2302
tri 13547 2278 13550 2319 nw
tri 13312 2258 13318 2278 ne
rect 13318 2258 13368 2278
tri 13368 2258 13374 2278 nw
tri 13432 2259 13434 2278 ne
rect 13434 2258 13544 2278
tri 13318 2243 13324 2258 ne
rect 13324 2243 13362 2258
tri 13362 2243 13368 2258 nw
tri 13434 2243 13435 2258 ne
rect 13435 2243 13544 2258
tri 13324 2239 13326 2243 ne
rect 13326 2239 13360 2243
tri 13360 2239 13362 2243 nw
tri 13435 2239 13436 2243 ne
rect 13436 2239 13544 2243
tri 13544 2239 13547 2278 nw
tri 13326 2232 13330 2239 ne
rect 13330 2232 13356 2239
tri 13356 2232 13360 2239 nw
rect 13436 2232 13540 2239
tri 13330 2225 13336 2232 ne
rect 13336 2225 13349 2232
tri 13349 2225 13356 2232 nw
tri 13436 2225 13437 2232 ne
tri 13336 2223 13343 2225 ne
tri 13343 2223 13349 2225 nw
rect 13437 2223 13540 2232
tri 13437 2202 13439 2223 ne
rect 13439 2202 13540 2223
tri 13540 2202 13544 2239 nw
tri 13439 2169 13444 2202 ne
rect 13444 2169 13536 2202
tri 13536 2169 13540 2202 nw
tri 13444 2138 13448 2169 ne
rect 13448 2138 13531 2169
tri 13531 2138 13536 2169 nw
tri 13448 2111 13454 2138 ne
rect 13454 2111 13526 2138
tri 13526 2111 13531 2138 nw
tri 13454 2088 13459 2111 ne
rect 13459 2088 13521 2111
tri 13521 2088 13526 2111 nw
tri 13459 2069 13465 2088 ne
rect 13465 2069 13515 2088
tri 13515 2069 13521 2088 nw
tri 13465 2053 13471 2069 ne
rect 13471 2053 13509 2069
tri 13509 2053 13515 2069 nw
tri 13471 2042 13477 2053 ne
rect 13477 2042 13503 2053
tri 13503 2042 13509 2053 nw
tri 13477 2036 13483 2042 ne
rect 13483 2036 13496 2042
tri 13496 2036 13503 2042 nw
tri 13483 2034 13490 2036 ne
tri 13490 2034 13496 2036 nw
tri 24257 -37 24279 -36 se
rect 24279 -37 24323 -36
tri 24323 -37 24345 -36 sw
tri 24236 -38 24257 -37 se
rect 24257 -38 24345 -37
tri 24345 -38 24366 -37 sw
tri 24215 -39 24236 -38 se
rect 24236 -39 24366 -38
tri 24366 -39 24387 -38 sw
tri 24195 -40 24215 -39 se
rect 24215 -40 24387 -39
tri 24387 -40 24407 -39 sw
tri 24177 -42 24195 -40 se
rect 24195 -42 24407 -40
tri 24407 -42 24425 -40 sw
tri 24159 -44 24177 -42 se
rect 24177 -44 24425 -42
tri 24425 -44 24443 -42 sw
tri 24143 -47 24159 -44 se
rect 24159 -47 24443 -44
tri 24443 -47 24459 -44 sw
tri 24128 -49 24143 -47 se
rect 24143 -49 24459 -47
tri 24459 -49 24474 -47 sw
tri 24115 -52 24128 -49 se
rect 24128 -52 24474 -49
tri 24474 -52 24487 -49 sw
tri 24103 -55 24115 -52 se
rect 24115 -55 24487 -52
tri 24487 -55 24499 -52 sw
tri 24094 -58 24103 -55 se
rect 24103 -58 24499 -55
tri 24499 -58 24508 -55 sw
tri 24087 -62 24094 -58 se
rect 24094 -62 24508 -58
tri 24508 -62 24515 -58 sw
tri 24081 -65 24087 -62 se
rect 24087 -65 24515 -62
tri 24515 -65 24521 -62 sw
tri 24078 -68 24081 -65 se
rect 24081 -68 24521 -65
tri 24521 -68 24524 -65 sw
tri 24077 -72 24078 -68 se
tri 24077 -76 24078 -72 ne
rect 24078 -76 24524 -68
tri 24524 -72 24525 -68 sw
tri 24524 -76 24525 -72 nw
tri 24078 -79 24081 -76 ne
rect 24081 -79 24521 -76
tri 24521 -79 24524 -76 nw
tri 24081 -82 24087 -79 ne
rect 24087 -82 24515 -79
tri 24515 -82 24521 -79 nw
tri 24087 -86 24094 -82 ne
rect 24094 -86 24508 -82
tri 24508 -86 24515 -82 nw
tri 24094 -89 24103 -86 ne
rect 24103 -89 24499 -86
tri 24499 -89 24508 -86 nw
tri 24103 -92 24115 -89 ne
rect 24115 -92 24487 -89
tri 24487 -92 24499 -89 nw
tri 24115 -95 24128 -92 ne
rect 24128 -95 24474 -92
tri 24474 -95 24487 -92 nw
tri 24128 -97 24143 -95 ne
rect 24143 -97 24459 -95
tri 24459 -97 24474 -95 nw
tri 24143 -100 24159 -97 ne
rect 24159 -100 24443 -97
tri 24443 -100 24459 -97 nw
tri 24159 -102 24177 -100 ne
rect 24177 -102 24425 -100
tri 24425 -102 24443 -100 nw
tri 24177 -104 24195 -102 ne
rect 24195 -104 24407 -102
tri 24407 -104 24425 -102 nw
tri 24195 -105 24215 -104 ne
rect 24215 -105 24387 -104
tri 24387 -105 24407 -104 nw
tri 24215 -106 24236 -105 ne
rect 24236 -106 24366 -105
tri 24366 -106 24387 -105 nw
tri 24236 -107 24257 -106 ne
rect 24257 -107 24345 -106
tri 24345 -107 24366 -106 nw
tri 24257 -108 24279 -107 ne
rect 24279 -108 24323 -107
tri 24323 -108 24345 -107 nw
tri 24257 -322 24279 -321 se
rect 24279 -322 24323 -321
tri 24323 -322 24345 -321 sw
tri 24236 -323 24257 -322 se
rect 24257 -323 24345 -322
tri 24345 -323 24366 -322 sw
tri 24215 -325 24236 -323 se
rect 24236 -325 24366 -323
tri 24366 -325 24387 -323 sw
tri 24195 -327 24215 -325 se
rect 24215 -327 24387 -325
tri 24387 -327 24407 -325 sw
tri 24177 -329 24195 -327 se
rect 24195 -329 24407 -327
tri 24407 -329 24425 -327 sw
tri 24159 -332 24177 -329 se
rect 24177 -332 24425 -329
tri 24425 -332 24443 -329 sw
tri 24143 -335 24159 -332 se
rect 24159 -335 24443 -332
tri 24443 -335 24459 -332 sw
tri 24128 -339 24143 -335 se
rect 24143 -339 24459 -335
tri 24459 -339 24474 -335 sw
tri 24115 -343 24128 -339 se
rect 24128 -343 24474 -339
tri 24474 -343 24487 -339 sw
tri 24103 -347 24115 -343 se
rect 24115 -347 24487 -343
tri 24487 -347 24499 -343 sw
tri 24094 -351 24103 -347 se
rect 24103 -351 24499 -347
tri 24499 -351 24508 -347 sw
tri 24087 -356 24094 -351 se
rect 24094 -356 24508 -351
tri 24508 -356 24515 -351 sw
tri 24081 -361 24087 -356 se
rect 24087 -361 24515 -356
tri 24515 -361 24521 -356 sw
tri 24078 -366 24081 -361 se
rect 24081 -366 24521 -361
tri 24521 -366 24524 -361 sw
tri 24077 -370 24078 -366 se
tri 24077 -375 24078 -370 ne
rect 24078 -375 24524 -366
tri 24524 -370 24525 -366 sw
tri 24524 -375 24525 -370 nw
tri 24078 -380 24081 -375 ne
rect 24081 -380 24521 -375
tri 24521 -380 24524 -375 nw
tri 24081 -385 24087 -380 ne
rect 24087 -385 24515 -380
tri 24515 -385 24521 -380 nw
tri 24087 -389 24094 -385 ne
rect 24094 -389 24508 -385
tri 24508 -389 24515 -385 nw
tri 24094 -394 24103 -389 ne
rect 24103 -394 24499 -389
tri 24499 -394 24508 -389 nw
tri 24103 -398 24115 -394 ne
rect 24115 -398 24487 -394
tri 24487 -398 24499 -394 nw
tri 24115 -402 24128 -398 ne
rect 24128 -402 24474 -398
tri 24474 -402 24487 -398 nw
tri 24128 -405 24143 -402 ne
rect 24143 -405 24459 -402
tri 24459 -405 24474 -402 nw
tri 24143 -409 24159 -405 ne
rect 24159 -409 24443 -405
tri 24443 -409 24459 -405 nw
tri 24159 -411 24177 -409 ne
rect 24177 -411 24425 -409
tri 24425 -411 24443 -409 nw
tri 24177 -414 24195 -411 ne
rect 24195 -414 24407 -411
tri 24407 -414 24425 -411 nw
tri 24195 -416 24215 -414 ne
rect 24215 -416 24387 -414
tri 24387 -416 24407 -414 nw
tri 24215 -418 24236 -416 ne
rect 24236 -418 24366 -416
tri 24366 -418 24387 -416 nw
tri 24236 -419 24257 -418 ne
rect 24257 -419 24345 -418
tri 24345 -419 24366 -418 nw
tri 24257 -420 24279 -419 ne
rect 24279 -420 24323 -419
tri 24323 -420 24345 -419 nw
tri 25546 -530 25579 -529 se
tri 25579 -530 25611 -529 sw
tri 25481 -531 25513 -530 se
rect 25513 -531 25644 -530
tri 25644 -531 25676 -530 sw
tri 25450 -532 25481 -531 se
rect 25481 -532 25676 -531
tri 25676 -532 25707 -531 sw
tri 25421 -534 25450 -532 se
rect 25450 -534 25707 -532
tri 25707 -534 25737 -532 sw
tri 25392 -536 25421 -534 se
rect 25421 -536 25737 -534
tri 25737 -536 25765 -534 sw
tri 25366 -538 25392 -536 se
rect 25392 -538 25765 -536
tri 25765 -538 25791 -536 sw
tri 25342 -541 25366 -538 se
rect 25366 -541 25791 -538
tri 25791 -541 25816 -538 sw
tri 25319 -544 25342 -541 se
rect 25342 -544 25816 -541
tri 25816 -544 25838 -541 sw
tri 25300 -547 25319 -544 se
rect 25319 -547 25838 -544
tri 25838 -547 25857 -544 sw
tri 25283 -550 25300 -547 se
rect 25300 -550 25857 -547
tri 25857 -550 25874 -547 sw
tri 25269 -554 25283 -550 se
rect 25283 -554 25874 -550
tri 25874 -554 25888 -550 sw
tri 25258 -557 25269 -554 se
rect 25269 -557 25888 -554
tri 25888 -557 25899 -554 sw
tri 25250 -561 25258 -557 se
rect 25258 -561 25899 -557
tri 25899 -561 25907 -557 sw
tri 25245 -565 25250 -561 se
rect 25250 -565 25907 -561
tri 25907 -565 25912 -561 sw
tri 25243 -569 25245 -565 se
tri 25243 -572 25245 -569 ne
rect 25245 -572 25912 -565
tri 25912 -569 25914 -565 sw
tri 25912 -572 25914 -569 nw
tri 25245 -576 25250 -572 ne
rect 25250 -576 25907 -572
tri 25907 -576 25912 -572 nw
tri 25250 -580 25258 -576 ne
rect 25258 -580 25899 -576
tri 25899 -580 25907 -576 nw
tri 25258 -584 25269 -580 ne
rect 25269 -584 25888 -580
tri 25888 -584 25899 -580 nw
tri 25269 -587 25283 -584 ne
rect 25283 -587 25874 -584
tri 25874 -587 25888 -584 nw
tri 25283 -590 25300 -587 ne
rect 25300 -590 25857 -587
tri 25857 -590 25874 -587 nw
tri 25300 -593 25319 -590 ne
rect 25319 -593 25838 -590
tri 25838 -593 25857 -590 nw
tri 25319 -596 25342 -593 ne
rect 25342 -596 25816 -593
tri 25816 -596 25838 -593 nw
tri 25342 -599 25366 -596 ne
rect 25366 -599 25791 -596
tri 25791 -599 25816 -596 nw
tri 25366 -601 25392 -599 ne
rect 25392 -601 25765 -599
tri 25765 -601 25791 -599 nw
tri 25392 -603 25421 -601 ne
rect 25421 -603 25737 -601
tri 25737 -603 25765 -601 nw
tri 25421 -605 25450 -603 ne
rect 25450 -605 25707 -603
tri 25707 -605 25737 -603 nw
tri 25450 -606 25481 -605 ne
rect 25481 -606 25676 -605
tri 25676 -606 25707 -605 nw
tri 25481 -607 25513 -606 ne
rect 25513 -607 25644 -606
tri 25644 -607 25676 -606 nw
tri 25513 -608 25546 -607 ne
rect 25546 -608 25611 -607
tri 25611 -608 25644 -607 nw
tri 25691 -737 25722 -736 se
rect 25722 -737 25783 -736
tri 25783 -737 25814 -736 sw
tri 25661 -738 25691 -737 se
rect 25691 -738 25814 -737
tri 25814 -738 25843 -737 sw
tri 25633 -739 25661 -738 se
rect 25661 -739 25843 -738
tri 25843 -739 25872 -738 sw
tri 25605 -741 25633 -739 se
rect 25633 -741 25872 -739
tri 25872 -741 25900 -739 sw
tri 25578 -743 25605 -741 se
rect 25605 -743 25900 -741
tri 25900 -743 25926 -741 sw
tri 25554 -745 25578 -743 se
rect 25578 -745 25926 -743
tri 25926 -745 25951 -743 sw
tri 25531 -748 25554 -745 se
rect 25554 -748 25951 -745
tri 25951 -748 25974 -745 sw
tri 25510 -751 25531 -748 se
rect 25531 -751 25974 -748
tri 25974 -751 25995 -748 sw
tri 25492 -754 25510 -751 se
rect 25510 -754 25995 -751
tri 25995 -754 26013 -751 sw
tri 25476 -757 25492 -754 se
rect 25492 -757 26013 -754
tri 26013 -757 26029 -754 sw
tri 25463 -760 25476 -757 se
rect 25476 -760 26029 -757
tri 26029 -760 26042 -757 sw
tri 25453 -764 25463 -760 se
rect 25463 -764 26042 -760
tri 26042 -764 26052 -760 sw
tri 25445 -768 25453 -764 se
rect 25453 -768 26052 -764
tri 26052 -768 26060 -764 sw
tri 25441 -772 25445 -768 se
rect 25445 -772 26060 -768
tri 26060 -772 26064 -768 sw
tri 25439 -775 25441 -772 se
tri 25439 -779 25441 -775 ne
rect 25441 -779 26064 -772
tri 26064 -775 26066 -772 sw
tri 26064 -779 26066 -775 nw
tri 25441 -783 25445 -779 ne
rect 25445 -783 26060 -779
tri 26060 -783 26064 -779 nw
tri 25445 -787 25453 -783 ne
rect 25453 -787 26052 -783
tri 26052 -787 26060 -783 nw
tri 25453 -790 25463 -787 ne
rect 25463 -790 26042 -787
tri 26042 -790 26052 -787 nw
tri 25463 -794 25476 -790 ne
rect 25476 -794 26029 -790
tri 26029 -794 26042 -790 nw
tri 25476 -797 25492 -794 ne
rect 25492 -797 26013 -794
tri 26013 -797 26029 -794 nw
tri 25492 -800 25510 -797 ne
rect 25510 -800 25995 -797
tri 25995 -800 26013 -797 nw
tri 25510 -803 25531 -800 ne
rect 25531 -803 25974 -800
tri 25974 -803 25995 -800 nw
tri 25531 -806 25554 -803 ne
rect 25554 -806 25951 -803
tri 25951 -806 25974 -803 nw
tri 25554 -808 25578 -806 ne
rect 25578 -808 25926 -806
tri 25926 -808 25951 -806 nw
tri 25578 -810 25605 -808 ne
rect 25605 -810 25900 -808
tri 25900 -810 25926 -808 nw
tri 25605 -812 25633 -810 ne
rect 25633 -812 25872 -810
tri 25872 -812 25900 -810 nw
tri 25633 -813 25661 -812 ne
rect 25661 -813 25843 -812
tri 25843 -813 25872 -812 nw
tri 25661 -814 25691 -813 ne
rect 25691 -814 25814 -813
tri 25814 -814 25843 -813 nw
tri 25722 -815 25752 -814 ne
tri 25752 -815 25783 -814 nw
tri 23374 -1320 23400 -1319 se
rect 23400 -1320 23453 -1319
tri 23453 -1320 23479 -1319 sw
tri 23366 -1321 23374 -1320 se
rect 23374 -1321 23479 -1320
tri 21651 -1322 21677 -1321 se
rect 21677 -1322 21730 -1321
tri 21730 -1322 21751 -1321 sw
tri 23349 -1322 23360 -1321 se
rect 23360 -1322 23479 -1321
tri 23479 -1322 23504 -1320 sw
tri 21626 -1324 21651 -1322 se
rect 21651 -1324 21756 -1322
tri 21756 -1324 21781 -1322 sw
tri 23330 -1324 23347 -1322 se
rect 23347 -1324 23504 -1322
tri 21601 -1327 21626 -1324 se
rect 21626 -1325 21781 -1324
tri 21781 -1325 21787 -1324 sw
tri 23324 -1325 23330 -1324 se
rect 23330 -1325 23504 -1324
tri 23504 -1325 23529 -1322 sw
rect 21626 -1327 21787 -1325
tri 21787 -1327 21806 -1325 sw
tri 23308 -1327 23324 -1325 se
rect 23324 -1327 23529 -1325
tri 21577 -1330 21601 -1327 se
rect 21601 -1328 21806 -1327
tri 21806 -1328 21814 -1327 sw
tri 23300 -1328 23308 -1327 se
rect 23308 -1328 23529 -1327
tri 23529 -1328 23553 -1325 sw
rect 21601 -1330 21814 -1328
tri 21814 -1330 21830 -1328 sw
tri 23289 -1330 23300 -1328 se
rect 23300 -1330 23553 -1328
tri 21555 -1333 21577 -1330 se
rect 21577 -1331 21830 -1330
tri 21830 -1331 21840 -1330 sw
tri 23278 -1331 23289 -1330 se
rect 23289 -1331 23553 -1330
tri 23553 -1331 23575 -1328 sw
rect 21577 -1333 21840 -1331
tri 21840 -1333 21852 -1331 sw
tri 23268 -1333 23278 -1331 se
rect 23278 -1333 23575 -1331
tri 21534 -1338 21555 -1333 se
rect 21555 -1336 21852 -1333
tri 21852 -1336 21864 -1333 sw
tri 23257 -1336 23268 -1333 se
rect 23268 -1336 23575 -1333
tri 23575 -1336 23596 -1331 sw
rect 21555 -1338 21864 -1336
tri 21864 -1338 21873 -1336 sw
tri 23249 -1338 23257 -1336 se
rect 23257 -1338 23596 -1336
tri 21514 -1343 21534 -1338 se
rect 21534 -1341 21873 -1338
tri 21873 -1341 21885 -1338 sw
tri 23237 -1341 23249 -1338 se
rect 23249 -1341 23596 -1338
tri 23596 -1341 23616 -1336 sw
rect 21534 -1343 21885 -1341
tri 21885 -1343 21893 -1341 sw
tri 23231 -1343 23237 -1341 se
rect 23237 -1343 23616 -1341
tri 21497 -1348 21514 -1343 se
rect 21514 -1346 21893 -1343
tri 21893 -1346 21904 -1343 sw
tri 23220 -1346 23231 -1343 se
rect 23231 -1346 23616 -1343
tri 23616 -1346 23633 -1341 sw
rect 21514 -1348 21904 -1346
tri 21904 -1348 21910 -1346 sw
tri 23215 -1348 23220 -1346 se
rect 23220 -1348 23633 -1346
tri 21481 -1354 21497 -1348 se
rect 21497 -1352 21910 -1348
tri 21910 -1352 21921 -1348 sw
tri 23204 -1352 23215 -1348 se
rect 23215 -1352 23633 -1348
tri 23633 -1352 23649 -1346 sw
rect 21497 -1354 21921 -1352
tri 21921 -1354 21926 -1352 sw
tri 23200 -1354 23204 -1352 se
rect 23204 -1354 23649 -1352
tri 21468 -1360 21481 -1354 se
rect 21481 -1358 21926 -1354
tri 21926 -1358 21935 -1354 sw
tri 23191 -1358 23200 -1354 se
rect 23200 -1358 23649 -1354
tri 23649 -1358 23663 -1352 sw
rect 21481 -1360 21935 -1358
tri 21935 -1360 21940 -1358 sw
tri 23187 -1360 23191 -1358 se
rect 23191 -1360 23663 -1358
tri 21456 -1367 21468 -1360 se
rect 21468 -1365 21940 -1360
tri 21940 -1365 21947 -1360 sw
tri 23179 -1365 23187 -1360 se
rect 23187 -1365 23663 -1360
tri 23663 -1365 23674 -1358 sw
rect 21468 -1367 21947 -1365
tri 21947 -1367 21951 -1365 sw
tri 23177 -1367 23179 -1365 se
rect 23179 -1367 23674 -1365
tri 21448 -1374 21456 -1367 se
rect 21456 -1372 21951 -1367
tri 21951 -1372 21957 -1367 sw
tri 23171 -1372 23177 -1367 se
rect 23177 -1372 23674 -1367
tri 23674 -1372 23683 -1365 sw
rect 21456 -1374 21957 -1372
tri 21957 -1374 21960 -1372 sw
tri 23169 -1374 23171 -1372 se
rect 23171 -1374 23683 -1372
tri 21441 -1381 21448 -1374 se
rect 21448 -1379 21960 -1374
tri 21960 -1379 21964 -1374 sw
tri 23164 -1379 23169 -1374 se
rect 23169 -1379 23683 -1374
tri 23683 -1379 23689 -1372 sw
rect 21448 -1381 21964 -1379
tri 21964 -1381 21966 -1379 sw
tri 23163 -1381 23164 -1379 se
rect 23164 -1381 23689 -1379
tri 21437 -1388 21441 -1381 se
rect 21441 -1386 21966 -1381
tri 21966 -1386 21969 -1381 sw
tri 23160 -1386 23163 -1381 se
rect 23163 -1386 23689 -1381
tri 23689 -1386 23693 -1379 sw
rect 21441 -1388 21969 -1386
tri 21969 -1388 21970 -1386 sw
tri 21436 -1396 21437 -1388 se
tri 21436 -1401 21437 -1396 ne
rect 21437 -1403 21970 -1388
tri 21970 -1396 21971 -1388 sw
tri 21970 -1401 21971 -1396 nw
tri 23159 -1394 23160 -1389 se
tri 23159 -1400 23160 -1394 ne
rect 23160 -1401 23693 -1386
tri 23693 -1394 23694 -1386 sw
tri 23693 -1401 23694 -1394 nw
tri 23160 -1403 23161 -1401 ne
rect 23161 -1403 23689 -1401
tri 21437 -1408 21440 -1403 ne
rect 21440 -1408 21967 -1403
tri 21967 -1408 21970 -1403 nw
tri 23161 -1408 23164 -1403 ne
rect 23164 -1408 23689 -1403
tri 23689 -1408 23693 -1401 nw
tri 21440 -1410 21441 -1408 ne
rect 21441 -1410 21966 -1408
tri 21966 -1410 21967 -1408 nw
tri 23164 -1410 23166 -1408 ne
rect 23166 -1410 23683 -1408
tri 21441 -1416 21446 -1410 ne
rect 21446 -1416 21961 -1410
tri 21961 -1416 21966 -1410 nw
tri 23166 -1416 23171 -1410 ne
rect 23171 -1416 23683 -1410
tri 23683 -1416 23689 -1408 nw
tri 21446 -1418 21448 -1416 ne
rect 21448 -1418 21960 -1416
tri 21960 -1418 21961 -1416 nw
tri 23171 -1418 23173 -1416 ne
rect 23173 -1418 23674 -1416
tri 21448 -1423 21454 -1418 ne
rect 21454 -1423 21953 -1418
tri 21953 -1423 21960 -1418 nw
tri 23173 -1423 23179 -1418 ne
rect 23179 -1423 23674 -1418
tri 23674 -1423 23683 -1416 nw
tri 21454 -1425 21456 -1423 ne
rect 21456 -1425 21951 -1423
tri 21951 -1425 21953 -1423 nw
tri 23179 -1425 23183 -1423 ne
rect 23183 -1425 23663 -1423
tri 21456 -1429 21464 -1425 ne
rect 21464 -1429 21943 -1425
tri 21943 -1429 21951 -1425 nw
tri 23183 -1429 23191 -1425 ne
rect 23191 -1429 23663 -1425
tri 23663 -1429 23674 -1423 nw
tri 21464 -1431 21468 -1429 ne
rect 21468 -1431 21940 -1429
tri 21940 -1431 21943 -1429 nw
tri 23191 -1431 23195 -1429 ne
rect 23195 -1431 23649 -1429
tri 21468 -1435 21477 -1431 ne
rect 21477 -1435 21931 -1431
tri 21931 -1435 21940 -1431 nw
tri 23195 -1435 23204 -1431 ne
rect 23204 -1435 23649 -1431
tri 23649 -1435 23663 -1429 nw
tri 21477 -1437 21481 -1435 ne
rect 21481 -1437 21926 -1435
tri 21926 -1437 21931 -1435 nw
tri 23204 -1437 23209 -1435 ne
rect 23209 -1437 23633 -1435
tri 21481 -1441 21491 -1437 ne
rect 21491 -1441 21916 -1437
tri 21916 -1441 21926 -1437 nw
tri 23209 -1441 23220 -1437 ne
rect 23220 -1441 23633 -1437
tri 23633 -1441 23649 -1435 nw
tri 21491 -1443 21497 -1441 ne
rect 21497 -1443 21910 -1441
tri 21910 -1443 21916 -1441 nw
tri 23220 -1443 23226 -1441 ne
rect 23226 -1443 23616 -1441
tri 21497 -1447 21508 -1443 ne
rect 21508 -1447 21899 -1443
tri 21899 -1447 21910 -1443 nw
tri 23226 -1447 23237 -1443 ne
rect 23237 -1447 23616 -1443
tri 23616 -1447 23633 -1441 nw
tri 21508 -1449 21514 -1447 ne
rect 21514 -1449 21893 -1447
tri 21893 -1449 21899 -1447 nw
tri 23237 -1449 23245 -1447 ne
rect 23245 -1449 23596 -1447
tri 21514 -1452 21526 -1449 ne
rect 21526 -1452 21881 -1449
tri 21881 -1452 21893 -1449 nw
tri 23245 -1452 23257 -1449 ne
rect 23257 -1452 23596 -1449
tri 23596 -1452 23616 -1447 nw
tri 21526 -1454 21534 -1452 ne
rect 21534 -1454 21873 -1452
tri 21873 -1454 21881 -1452 nw
tri 23257 -1454 23266 -1452 ne
rect 23266 -1454 23575 -1452
tri 21534 -1456 21545 -1454 ne
rect 21545 -1456 21862 -1454
tri 21862 -1456 21873 -1454 nw
tri 23266 -1456 23278 -1454 ne
rect 23278 -1456 23575 -1454
tri 23575 -1456 23596 -1452 nw
tri 21545 -1458 21555 -1456 ne
rect 21555 -1458 21852 -1456
tri 21852 -1458 21862 -1456 nw
tri 23278 -1458 23290 -1456 ne
rect 23290 -1458 23553 -1456
tri 21555 -1460 21566 -1458 ne
rect 21566 -1460 21842 -1458
tri 21842 -1460 21852 -1458 nw
tri 23290 -1460 23300 -1458 ne
rect 23300 -1460 23553 -1458
tri 23553 -1460 23575 -1456 nw
tri 21566 -1462 21577 -1460 ne
rect 21577 -1462 21830 -1460
tri 21830 -1462 21842 -1460 nw
tri 23300 -1462 23316 -1460 ne
rect 23316 -1462 23529 -1460
tri 21577 -1463 21585 -1462 ne
rect 21585 -1463 21822 -1462
tri 21822 -1463 21830 -1462 nw
tri 23316 -1463 23324 -1462 ne
rect 23324 -1463 23529 -1462
tri 23529 -1463 23553 -1460 nw
tri 21585 -1465 21601 -1463 ne
rect 21601 -1465 21806 -1463
tri 21806 -1465 21822 -1463 nw
tri 23324 -1465 23343 -1463 ne
rect 23343 -1465 23504 -1463
tri 21601 -1466 21607 -1465 ne
rect 21607 -1466 21800 -1465
tri 21800 -1466 21806 -1465 nw
tri 23343 -1466 23349 -1465 ne
rect 23349 -1466 23504 -1465
tri 23504 -1466 23529 -1463 nw
tri 21607 -1467 21624 -1466 ne
rect 21624 -1467 21783 -1466
tri 21783 -1467 21800 -1466 nw
tri 23349 -1467 23374 -1466 ne
rect 23374 -1467 23479 -1466
tri 23479 -1467 23504 -1466 nw
tri 21624 -1468 21626 -1467 ne
rect 21626 -1468 21781 -1467
tri 21781 -1468 21783 -1467 nw
tri 23374 -1468 23380 -1467 ne
rect 23380 -1468 23453 -1467
tri 23453 -1468 23479 -1467 nw
tri 21637 -1469 21643 -1468 ne
rect 21643 -1469 21764 -1468
tri 21764 -1469 21770 -1468 nw
tri 23400 -1469 23427 -1468 ne
tri 23427 -1469 23453 -1468 nw
tri 21651 -1470 21677 -1469 ne
rect 21677 -1470 21730 -1469
tri 21730 -1470 21756 -1469 nw
tri 21677 -1471 21704 -1470 ne
tri 21704 -1471 21730 -1470 nw
tri 21651 -1755 21677 -1754 se
rect 21677 -1755 21730 -1754
tri 21730 -1755 21756 -1754 sw
tri 23374 -1755 23400 -1754 se
rect 23400 -1755 23453 -1754
tri 23453 -1755 23479 -1754 sw
tri 21626 -1757 21651 -1755 se
rect 21651 -1757 21756 -1755
tri 21756 -1757 21781 -1755 sw
tri 23349 -1757 23374 -1755 se
rect 23374 -1757 23479 -1755
tri 23479 -1757 23504 -1755 sw
tri 21601 -1760 21626 -1757 se
rect 21626 -1760 21781 -1757
tri 21781 -1760 21806 -1757 sw
tri 23324 -1760 23349 -1757 se
rect 23349 -1760 23504 -1757
tri 23504 -1760 23529 -1757 sw
tri 21577 -1763 21601 -1760 se
rect 21601 -1763 21806 -1760
tri 21806 -1763 21830 -1760 sw
tri 23300 -1763 23324 -1760 se
rect 23324 -1763 23529 -1760
tri 23529 -1763 23553 -1760 sw
tri 21555 -1766 21577 -1763 se
rect 21577 -1766 21830 -1763
tri 21830 -1766 21852 -1763 sw
tri 23278 -1766 23300 -1763 se
rect 23300 -1766 23553 -1763
tri 23553 -1766 23575 -1763 sw
tri 21534 -1771 21555 -1766 se
rect 21555 -1771 21852 -1766
tri 21852 -1771 21873 -1766 sw
tri 23257 -1771 23278 -1766 se
rect 23278 -1771 23575 -1766
tri 23575 -1771 23596 -1766 sw
tri 21514 -1776 21534 -1771 se
rect 21534 -1776 21873 -1771
tri 21873 -1776 21893 -1771 sw
tri 23237 -1776 23257 -1771 se
rect 23257 -1776 23596 -1771
tri 23596 -1776 23616 -1771 sw
tri 21497 -1781 21514 -1776 se
rect 21514 -1781 21893 -1776
tri 21893 -1781 21910 -1776 sw
tri 23220 -1781 23237 -1776 se
rect 23237 -1781 23616 -1776
tri 23616 -1781 23633 -1776 sw
tri 21481 -1787 21497 -1781 se
rect 21497 -1787 21910 -1781
tri 21910 -1787 21926 -1781 sw
tri 23204 -1787 23220 -1781 se
rect 23220 -1787 23633 -1781
tri 23633 -1787 23649 -1781 sw
tri 21468 -1793 21481 -1787 se
rect 21481 -1793 21926 -1787
tri 21926 -1793 21940 -1787 sw
tri 23191 -1793 23204 -1787 se
rect 23204 -1793 23649 -1787
tri 23649 -1793 23663 -1787 sw
tri 21456 -1800 21468 -1793 se
rect 21468 -1800 21940 -1793
tri 21940 -1800 21951 -1793 sw
tri 23179 -1800 23191 -1793 se
rect 23191 -1800 23663 -1793
tri 23663 -1800 23674 -1793 sw
tri 21448 -1807 21456 -1800 se
rect 21456 -1807 21951 -1800
tri 21951 -1807 21960 -1800 sw
tri 23171 -1807 23179 -1800 se
rect 23179 -1807 23674 -1800
tri 23674 -1807 23683 -1800 sw
tri 21441 -1814 21448 -1807 se
rect 21448 -1814 21960 -1807
tri 21960 -1814 21966 -1807 sw
tri 23164 -1814 23171 -1807 se
rect 23171 -1814 23683 -1807
tri 23683 -1814 23689 -1807 sw
tri 21437 -1821 21441 -1814 se
rect 21441 -1821 21966 -1814
tri 21966 -1821 21970 -1814 sw
tri 23160 -1821 23164 -1814 se
rect 23164 -1821 23689 -1814
tri 23689 -1821 23693 -1814 sw
tri 21436 -1829 21437 -1821 se
tri 21436 -1836 21437 -1829 ne
rect 21437 -1836 21970 -1821
tri 21970 -1829 21971 -1821 sw
tri 21970 -1836 21971 -1829 nw
tri 23159 -1829 23160 -1821 se
tri 23159 -1836 23160 -1829 ne
rect 23160 -1836 23693 -1821
tri 23693 -1829 23694 -1821 sw
tri 23693 -1836 23694 -1829 nw
tri 21437 -1843 21441 -1836 ne
rect 21441 -1843 21966 -1836
tri 21966 -1843 21970 -1836 nw
tri 23160 -1843 23164 -1836 ne
rect 23164 -1843 23689 -1836
tri 23689 -1843 23693 -1836 nw
tri 21441 -1851 21448 -1843 ne
rect 21448 -1851 21960 -1843
tri 21960 -1851 21966 -1843 nw
tri 23164 -1851 23171 -1843 ne
rect 23171 -1851 23683 -1843
tri 23683 -1851 23689 -1843 nw
tri 21448 -1858 21456 -1851 ne
rect 21456 -1858 21951 -1851
tri 21951 -1858 21960 -1851 nw
tri 23171 -1858 23179 -1851 ne
rect 23179 -1858 23674 -1851
tri 23674 -1858 23683 -1851 nw
tri 21456 -1864 21468 -1858 ne
rect 21468 -1864 21940 -1858
tri 21940 -1864 21951 -1858 nw
tri 23179 -1864 23191 -1858 ne
rect 23191 -1864 23663 -1858
tri 23663 -1864 23674 -1858 nw
tri 21468 -1870 21481 -1864 ne
rect 21481 -1870 21926 -1864
tri 21926 -1870 21940 -1864 nw
tri 23191 -1870 23204 -1864 ne
rect 23204 -1870 23649 -1864
tri 23649 -1870 23663 -1864 nw
tri 21481 -1876 21497 -1870 ne
rect 21497 -1876 21910 -1870
tri 21910 -1876 21926 -1870 nw
tri 23204 -1876 23220 -1870 ne
rect 23220 -1876 23633 -1870
tri 23633 -1876 23649 -1870 nw
tri 21497 -1882 21514 -1876 ne
rect 21514 -1882 21893 -1876
tri 21893 -1882 21910 -1876 nw
tri 23220 -1882 23237 -1876 ne
rect 23237 -1882 23616 -1876
tri 23616 -1882 23633 -1876 nw
tri 21514 -1887 21534 -1882 ne
rect 21534 -1887 21873 -1882
tri 21873 -1887 21893 -1882 nw
tri 23237 -1887 23257 -1882 ne
rect 23257 -1887 23596 -1882
tri 23596 -1887 23616 -1882 nw
tri 21534 -1891 21555 -1887 ne
rect 21555 -1891 21852 -1887
tri 21852 -1891 21873 -1887 nw
tri 23257 -1891 23278 -1887 ne
rect 23278 -1891 23575 -1887
tri 23575 -1891 23596 -1887 nw
tri 21555 -1895 21577 -1891 ne
rect 21577 -1895 21830 -1891
tri 21830 -1895 21852 -1891 nw
tri 23278 -1895 23300 -1891 ne
rect 23300 -1895 23553 -1891
tri 23553 -1895 23575 -1891 nw
tri 21577 -1898 21601 -1895 ne
rect 21601 -1898 21806 -1895
tri 21806 -1898 21830 -1895 nw
tri 23300 -1898 23324 -1895 ne
rect 23324 -1898 23529 -1895
tri 23529 -1898 23553 -1895 nw
tri 21601 -1901 21626 -1898 ne
rect 21626 -1901 21781 -1898
tri 21781 -1901 21806 -1898 nw
tri 23324 -1901 23349 -1898 ne
rect 23349 -1901 23504 -1898
tri 23504 -1901 23529 -1898 nw
tri 21626 -1902 21651 -1901 ne
rect 21651 -1902 21756 -1901
tri 21756 -1902 21781 -1901 nw
tri 23349 -1902 23374 -1901 ne
rect 23374 -1902 23479 -1901
tri 23479 -1902 23504 -1901 nw
tri 21651 -1903 21677 -1902 ne
rect 21677 -1903 21730 -1902
tri 21730 -1903 21756 -1902 nw
tri 23374 -1903 23400 -1902 ne
rect 23400 -1903 23453 -1902
tri 23453 -1903 23479 -1902 nw
tri 21677 -1904 21704 -1903 ne
tri 21704 -1904 21730 -1903 nw
tri 23400 -1904 23427 -1903 ne
tri 23427 -1904 23453 -1903 nw
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1707688321
transform 1 0 16973 0 1 4222
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1707688321
transform 1 0 3946 0 1 4026
box 0 0 1 1
use L1M1_CDNS_52468879185193  L1M1_CDNS_52468879185193_0
timestamp 1707688321
transform -1 0 21519 0 1 -1923
box 0 0 1 1
use L1M1_CDNS_524688791851191  L1M1_CDNS_524688791851191_0
timestamp 1707688321
transform -1 0 12475 0 1 2841
box -12 -6 766 112
use L1M1_CDNS_524688791851443  L1M1_CDNS_524688791851443_0
timestamp 1707688321
transform 1 0 11729 0 1 4102
box -12 -6 694 112
use L1M1_CDNS_524688791851444  L1M1_CDNS_524688791851444_0
timestamp 1707688321
transform 1 0 19124 0 1 4223
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1707688321
transform -1 0 17609 0 1 5375
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1707688321
transform -1 0 17020 0 1 4210
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1707688321
transform 0 -1 24281 1 0 10869
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1707688321
transform 0 -1 23795 1 0 13188
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1707688321
transform 1 0 16495 0 1 2465
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_5
timestamp 1707688321
transform 1 0 25505 0 1 9922
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_6
timestamp 1707688321
transform 1 0 25666 0 1 10812
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_7
timestamp 1707688321
transform 1 0 25294 0 1 10812
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_8
timestamp 1707688321
transform 1 0 25705 0 1 10504
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_9
timestamp 1707688321
transform 1 0 25402 0 1 10072
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_10
timestamp 1707688321
transform 1 0 25256 0 1 10504
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_11
timestamp 1707688321
transform 1 0 27434 0 1 10905
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_12
timestamp 1707688321
transform 1 0 24735 0 1 10905
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_13
timestamp 1707688321
transform 1 0 24189 0 1 10071
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_14
timestamp 1707688321
transform 1 0 28063 0 1 10072
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_15
timestamp 1707688321
transform 1 0 27499 0 1 10504
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_16
timestamp 1707688321
transform 1 0 25241 0 1 9727
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_17
timestamp 1707688321
transform 1 0 27658 0 1 9922
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_18
timestamp 1707688321
transform 1 0 27306 0 1 9728
box 0 0 1 1
use M1M2_CDNS_52468879185197  M1M2_CDNS_52468879185197_0
timestamp 1707688321
transform -1 0 27257 0 1 -2273
box 0 0 256 116
use M1M2_CDNS_52468879185197  M1M2_CDNS_52468879185197_1
timestamp 1707688321
transform 1 0 753 0 1 415
box 0 0 256 116
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_0
timestamp 1707688321
transform 0 -1 5978 -1 0 4139
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_1
timestamp 1707688321
transform -1 0 17391 0 -1 2632
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_2
timestamp 1707688321
transform 0 -1 5978 1 0 2209
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_3
timestamp 1707688321
transform 1 0 14334 0 1 2761
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_4
timestamp 1707688321
transform 1 0 14334 0 1 4269
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_0
timestamp 1707688321
transform 1 0 5338 0 1 3594
box 0 0 1 1
use M1M2_CDNS_52468879185204  M1M2_CDNS_52468879185204_0
timestamp 1707688321
transform 1 0 2098 0 1 1786
box 0 0 1 1
use M1M2_CDNS_52468879185204  M1M2_CDNS_52468879185204_1
timestamp 1707688321
transform 1 0 2098 0 1 2712
box 0 0 1 1
use M1M2_CDNS_52468879185204  M1M2_CDNS_52468879185204_2
timestamp 1707688321
transform 1 0 2098 0 1 3594
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_0
timestamp 1707688321
transform 0 -1 4488 1 0 1332
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_1
timestamp 1707688321
transform 0 -1 4488 1 0 3148
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_2
timestamp 1707688321
transform 0 -1 7846 1 0 2715
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_3
timestamp 1707688321
transform 0 -1 8262 1 0 1789
box 0 0 1 1
use M1M2_CDNS_52468879185371  M1M2_CDNS_52468879185371_0
timestamp 1707688321
transform 1 0 23699 0 -1 1213
box 0 0 1 1
use M1M2_CDNS_52468879185371  M1M2_CDNS_52468879185371_1
timestamp 1707688321
transform 1 0 15699 0 1 3877
box 0 0 1 1
use M1M2_CDNS_52468879185961  M1M2_CDNS_52468879185961_0
timestamp 1707688321
transform 0 1 22947 -1 0 4270
box 0 0 1 1
use M1M2_CDNS_52468879185961  M1M2_CDNS_52468879185961_1
timestamp 1707688321
transform 1 0 23635 0 -1 1213
box 0 0 1 1
use M1M2_CDNS_52468879185972  M1M2_CDNS_52468879185972_0
timestamp 1707688321
transform 1 0 23571 0 -1 1213
box 0 0 1 1
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_0
timestamp 1707688321
transform 1 0 16668 0 1 1673
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_1
timestamp 1707688321
transform 1 0 14251 0 1 413
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_2
timestamp 1707688321
transform 1 0 14251 0 1 1673
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_3
timestamp 1707688321
transform 1 0 13561 0 1 2835
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_4
timestamp 1707688321
transform 1 0 13561 0 1 1918
box 0 0 192 180
use M1M2_CDNS_524688791851084  M1M2_CDNS_524688791851084_0
timestamp 1707688321
transform 0 1 23161 -1 0 1852
box 0 0 512 52
use M1M2_CDNS_524688791851250  M1M2_CDNS_524688791851250_0
timestamp 1707688321
transform 0 -1 11889 1 0 3766
box 0 0 448 180
use M1M2_CDNS_524688791851445  M1M2_CDNS_524688791851445_0
timestamp 1707688321
transform 1 0 23967 0 -1 5614
box 0 0 128 3892
use M1M2_CDNS_524688791851446  M1M2_CDNS_524688791851446_0
timestamp 1707688321
transform 1 0 15699 0 1 2255
box 0 0 704 116
use M1M2_CDNS_524688791851446  M1M2_CDNS_524688791851446_1
timestamp 1707688321
transform 1 0 15699 0 1 4432
box 0 0 704 116
use M2M3_CDNS_524688791851447  M2M3_CDNS_524688791851447_0
timestamp 1707688321
transform 1 0 11700 0 1 3755
box -5 0 221 474
use M2short_CDNS_524688791851492  M2short_CDNS_524688791851492_0
timestamp 1707688321
transform 0 -1 25384 1 0 10669
box 0 0 1 1
use M2short_CDNS_524688791851493  M2short_CDNS_524688791851493_0
timestamp 1707688321
transform 1 0 13386 0 1 2433
box 0 0 1 1
use M2short_CDNS_524688791851494  M2short_CDNS_524688791851494_0
timestamp 1707688321
transform 0 -1 13408 1 0 2633
box 0 0 1 1
use M2short_CDNS_524688791851494  M2short_CDNS_524688791851494_1
timestamp 1707688321
transform 1 0 17398 0 1 2516
box 0 0 1 1
use M2short_CDNS_524688791851494  M2short_CDNS_524688791851494_2
timestamp 1707688321
transform 1 0 62 0 1 833
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_0
timestamp 1707688321
transform -1 0 4062 0 1 4010
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_1
timestamp 1707688321
transform -1 0 1920 0 1 4010
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_2
timestamp 1707688321
transform 1 0 16960 0 1 4207
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_3
timestamp 1707688321
transform 1 0 19102 0 1 4207
box 0 0 1 1
use PYres_CDNS_524688791856  PYres_CDNS_524688791856_0
timestamp 1707688321
transform -1 0 19118 0 1 4190
box -50 0 2090 100
use PYres_CDNS_524688791856  PYres_CDNS_524688791856_1
timestamp 1707688321
transform 1 0 1904 0 1 3993
box -50 0 2090 100
use s8_esd_res75only_noshorts_nometal  s8_esd_res75only_noshorts_nometal_0
timestamp 1707688321
transform 0 -1 12488 -1 0 4230
box 2 0 1466 804
use sky130_fd_io__sio_hotswap_bias  sky130_fd_io__sio_hotswap_bias_0
timestamp 1707688321
transform 1 0 16648 0 1 4745
box 15 0 6144 4780
use sky130_fd_io__sio_hotswap_nonoverlap  sky130_fd_io__sio_hotswap_nonoverlap_0
timestamp 1707688321
transform 1 0 26057 0 1 3516
box -603 -778 2953 6069
use sky130_fd_io__sio_hotswap_pghs  sky130_fd_io__sio_hotswap_pghs_0
timestamp 1707688321
transform 1 0 10049 0 1 -2365
box -91 -99 19259 17793
use sky130_fd_io__sio_hotswap_pug  sky130_fd_io__sio_hotswap_pug_0
timestamp 1707688321
transform 0 -1 8374 -1 0 2894
box -289 20 603 3310
use sky130_fd_io__sio_hotswap_pug  sky130_fd_io__sio_hotswap_pug_1
timestamp 1707688321
transform 0 1 1728 -1 0 2894
box -289 20 603 3310
use sky130_fd_io__sio_hotswap_pug  sky130_fd_io__sio_hotswap_pug_2
timestamp 1707688321
transform 0 1 5202 1 0 3464
box -289 20 603 3310
use sky130_fd_io__sio_hotswap_pug  sky130_fd_io__sio_hotswap_pug_3
timestamp 1707688321
transform 0 1 1728 1 0 1656
box -289 20 603 3310
use sky130_fd_io__sio_hotswap_pug  sky130_fd_io__sio_hotswap_pug_4
timestamp 1707688321
transform 0 1 1728 1 0 3464
box -289 20 603 3310
use sky130_fd_io__sio_hotswap_pug  sky130_fd_io__sio_hotswap_pug_5
timestamp 1707688321
transform 0 -1 8374 1 0 1656
box -289 20 603 3310
<< labels >>
flabel comment s 29502 6414 29502 6414 0 FreeSans 200 0 0 0 padlo
flabel comment s 21728 -1864 21728 -1864 0 FreeSans 600 180 0 0 ModB10X
flabel comment s 15189 4701 15189 4701 0 FreeSans 600 90 0 0 ModA1X
flabel comment s 13487 2492 13487 2492 0 FreeSans 600 90 0 0 ModA2X/ModB2Y
flabel comment s 17425 2592 17425 2592 0 FreeSans 400 0 0 0 ModA3X/ModB3Y
flabel comment s 21238 2629 21238 2629 0 FreeSans 1000 0 0 0 pghs_h_int
flabel comment s 26210 10922 26210 10922 0 FreeSans 400 0 0 0 ModA6
flabel comment s 20527 8597 20527 8597 0 FreeSans 400 0 0 0 MOdA3Y
flabel comment s 25752 -779 25752 -779 0 FreeSans 400 0 0 0 ModA4Y
flabel comment s 23451 -1864 23451 -1864 0 FreeSans 600 180 0 0 ModB10X
flabel comment s 14980 4701 14980 4701 0 FreeSans 600 90 0 0 ModA1Y
flabel comment s 13340 2696 13340 2696 0 FreeSans 600 90 0 0 ModA2Y/ModB2X
flabel comment s 20077 3157 20077 3157 0 FreeSans 400 270 0 0 ModB3X
flabel comment s 13309 5445 13309 5445 0 FreeSans 400 0 0 0 ModB4Y
flabel comment s 13397 5511 13397 5511 0 FreeSans 400 0 0 0 ModB4X
flabel comment s 25607 11591 25607 11591 0 FreeSans 600 90 0 0 ModB6X
flabel comment s 25632 10537 25632 10537 0 FreeSans 600 0 0 0 ModB6Y
flabel comment s 25489 10173 25489 10173 0 FreeSans 400 0 0 0 ModA5Y/ModB5X
flabel comment s 24298 -73 24298 -73 0 FreeSans 600 0 0 0 ModB7X
flabel comment s 24298 -380 24298 -380 0 FreeSans 600 0 0 0 ModB8X
flabel comment s 29506 6587 29506 6587 0 FreeSans 200 0 0 0 pu_h_n<0>
flabel comment s 29506 6500 29506 6500 0 FreeSans 200 0 0 0 vpb_drvr
flabel comment s 29506 6325 29506 6325 0 FreeSans 200 0 0 0 p2g
flabel comment s 29506 6240 29506 6240 0 FreeSans 200 0 0 0 n2
flabel comment s 29506 6150 29506 6150 0 FreeSans 200 0 0 0 p1g
flabel comment s 29506 6064 29506 6064 0 FreeSans 200 0 0 0 pghs_h_int
flabel comment s 23451 -1429 23451 -1429 0 FreeSans 600 180 0 0 ModB10X
flabel comment s 21728 -1429 21728 -1429 0 FreeSans 600 180 0 0 ModB10X
flabel comment s 26933 12450 26933 12450 0 FreeSans 600 180 0 0 ModB5Y
flabel comment s 25565 -588 25565 -588 0 FreeSans 400 180 0 0 ModA4X
flabel comment s 26456 10658 26456 10658 0 FreeSans 400 90 0 0 ModA6B
flabel comment s 23162 10053 23162 10053 0 FreeSans 600 180 0 0 padlo
flabel comment s 23168 10235 23168 10235 0 FreeSans 600 0 0 0 p2g
flabel comment s 23169 9955 23169 9955 0 FreeSans 600 0 0 0 p1g
flabel metal1 s 20975 6790 21921 6963 0 FreeSans 800 0 0 0 vcc_io
port 2 nsew
flabel metal1 s 7349 4078 7349 4078 0 FreeSans 400 0 0 0 tie_hi
flabel metal1 s 16510 4197 16510 4197 0 FreeSans 600 0 0 0 padlo
flabel metal1 s 20975 6526 21921 6699 0 FreeSans 800 0 0 0 vcc_io
port 2 nsew
flabel metal1 s 20975 6265 21921 6438 0 FreeSans 800 0 0 0 vcc_io
port 2 nsew
flabel metal1 s 20975 5999 21921 6172 0 FreeSans 800 0 0 0 vcc_io
port 2 nsew
flabel metal1 s 20975 5734 21921 5907 0 FreeSans 800 0 0 0 vcc_io
port 2 nsew
flabel metal1 s 20975 5470 21921 5643 0 FreeSans 800 0 0 0 vcc_io
port 2 nsew
flabel metal1 s 21199 -1929 21480 -1883 0 FreeSans 400 180 0 0 vpwr_ka
port 3 nsew
flabel metal1 s 22198 4819 22571 4905 0 FreeSans 400 0 0 0 vgnd
port 4 nsew
flabel metal1 s 14462 4624 14489 4676 0 FreeSans 600 270 0 0 p2g
port 5 nsew
flabel metal5 s 29810 56 29810 56 0 FreeSans 600 0 0 0 pghs_h_int
flabel metal5 s 29819 4682 29819 4682 0 FreeSans 800 0 0 0 vpb_drvr
flabel metal5 s 29810 2819 29810 2819 0 FreeSans 1200 0 0 0 p2g
flabel metal5 s 29810 1882 29810 1882 0 FreeSans 1200 0 0 0 n2
flabel metal5 s 29810 961 29810 961 0 FreeSans 1200 0 0 0 p1g
flabel metal5 s 29799 5606 29799 5606 0 FreeSans 600 0 0 0 pu_h_n<0>
flabel metal5 s 29813 3747 29813 3747 0 FreeSans 1200 0 0 0 padlo
flabel metal3 s 11695 3983 11921 4069 0 FreeSans 400 0 0 0 pad
port 6 nsew
flabel metal2 s 23583 -1899 23839 -1783 0 FreeSans 400 0 0 0 vgnd
port 4 nsew
flabel metal2 s 23037 -2275 23089 -2253 0 FreeSans 200 0 0 0 force_h<1>
port 7 nsew
flabel metal2 s 20884 -2464 20936 -2425 0 FreeSans 400 0 0 0 oe_hs_h
port 8 nsew
flabel metal2 s 28226 -2129 28278 -2077 0 FreeSans 400 180 0 0 od_h
port 9 nsew
flabel metal2 s 24908 -1953 25101 -1909 0 FreeSans 200 0 0 0 vcc_io
port 2 nsew
flabel metal2 s 23932 8641 24514 9132 0 FreeSans 600 0 0 0 vcc_io
port 2 nsew
flabel metal2 s 23867 -2273 24123 -2103 0 FreeSans 400 0 0 0 vgnd
port 4 nsew
flabel metal2 s 25993 10225 26429 10300 0 FreeSans 800 0 0 0 vpb_drvr
port 10 nsew
flabel metal2 s 24392 12365 24721 12603 0 FreeSans 600 0 0 0 vcc_io
port 2 nsew
flabel metal2 s -232 3962 -173 4014 3 FreeSans 400 0 0 0 pug_h<3>
port 11 nsew
flabel metal2 s -232 3594 -177 3646 3 FreeSans 400 0 0 0 pug_h<2>
port 12 nsew
flabel metal2 s -232 2712 -172 2764 3 FreeSans 400 0 0 0 pug_h<1>
port 13 nsew
flabel metal2 s -232 1786 -167 1838 3 FreeSans 400 0 0 0 pug_h<0>
port 14 nsew
flabel metal2 s 15699 4206 16439 4281 0 FreeSans 800 0 0 0 vpb_drvr
port 10 nsew
flabel metal2 s 7730 4624 7846 4660 0 FreeSans 400 0 0 0 pug_h<4>
port 15 nsew
flabel metal2 s 16964 4652 16964 4652 0 FreeSans 200 270 0 0 vcc_io_soft
flabel metal2 s -232 833 -121 949 3 FreeSans 1000 0 0 0 pghs_h
port 16 nsew
flabel metal2 s 8146 4626 8262 4660 0 FreeSans 400 0 0 0 pug_h<5>
port 17 nsew
<< properties >>
string GDS_END 90825434
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 89708954
string path 749.275 123.750 749.275 120.100 
<< end >>
