magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -89 -36 585 236
<< pmos >>
rect 0 0 36 200
rect 92 0 128 200
rect 184 0 220 200
rect 276 0 312 200
rect 368 0 404 200
rect 460 0 496 200
<< pdiff >>
rect -50 0 0 200
rect 496 0 546 200
<< poly >>
rect 0 200 36 226
rect 0 -26 36 0
rect 92 200 128 226
rect 92 -26 128 0
rect 184 200 220 226
rect 184 -26 220 0
rect 276 200 312 226
rect 276 -26 312 0
rect 368 200 404 226
rect 368 -26 404 0
rect 460 200 496 226
rect 460 -26 496 0
<< metal1 >>
rect -51 -16 -5 186
rect 41 -16 87 186
rect 133 -16 179 186
rect 225 -16 271 186
rect 317 -16 363 186
rect 409 -16 455 186
rect 501 -16 547 186
use DFM1sd2_CDNS_524688791851378  DFM1sd2_CDNS_524688791851378_0
timestamp 1707688321
transform 1 0 404 0 1 0
box -36 -36 92 236
use DFM1sd2_CDNS_524688791851378  DFM1sd2_CDNS_524688791851378_1
timestamp 1707688321
transform 1 0 312 0 1 0
box -36 -36 92 236
use DFM1sd2_CDNS_524688791851378  DFM1sd2_CDNS_524688791851378_2
timestamp 1707688321
transform 1 0 220 0 1 0
box -36 -36 92 236
use DFM1sd2_CDNS_524688791851378  DFM1sd2_CDNS_524688791851378_3
timestamp 1707688321
transform 1 0 128 0 1 0
box -36 -36 92 236
use DFM1sd2_CDNS_524688791851378  DFM1sd2_CDNS_524688791851378_4
timestamp 1707688321
transform 1 0 36 0 1 0
box -36 -36 92 236
use DFM1sd_CDNS_524688791851377  DFM1sd_CDNS_524688791851377_0
timestamp 1707688321
transform -1 0 0 0 1 0
box -36 -36 89 236
use DFM1sd_CDNS_524688791851377  DFM1sd_CDNS_524688791851377_1
timestamp 1707688321
transform 1 0 496 0 1 0
box -36 -36 89 236
<< labels >>
flabel comment s -28 85 -28 85 0 FreeSans 300 0 0 0 S
flabel comment s 64 85 64 85 0 FreeSans 300 0 0 0 D
flabel comment s 156 85 156 85 0 FreeSans 300 0 0 0 S
flabel comment s 248 85 248 85 0 FreeSans 300 0 0 0 D
flabel comment s 340 85 340 85 0 FreeSans 300 0 0 0 S
flabel comment s 432 85 432 85 0 FreeSans 300 0 0 0 D
flabel comment s 524 85 524 85 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 85971138
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85967758
<< end >>
