magic
tech sky130A
timestamp 1707688321
<< metal1 >>
rect 0 0 3 218
rect 125 0 128 218
<< via1 >>
rect 3 0 125 218
<< metal2 >>
rect 0 0 3 218
rect 125 0 128 218
<< properties >>
string GDS_END 86911404
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86909480
<< end >>
