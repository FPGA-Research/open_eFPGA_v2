magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< pwell >>
rect 1179 1269 1189 1279
rect 467 1202 491 1253
rect 1277 1202 1301 1253
rect 467 350 491 401
rect 1277 350 1301 401
<< obsli1 >>
rect 0 0 1686 1770
<< obsm1 >>
rect 0 1704 1686 1770
rect 0 918 66 1704
rect 113 1343 141 1676
rect 169 1371 197 1704
rect 225 1343 253 1676
rect 281 1371 309 1704
rect 337 1343 365 1676
rect 411 1343 465 1676
rect 511 1343 539 1676
rect 567 1371 595 1704
rect 623 1343 651 1676
rect 679 1371 707 1704
rect 735 1343 763 1676
rect 113 1279 763 1343
rect 113 946 141 1279
rect 169 918 197 1251
rect 225 946 253 1279
rect 281 918 309 1251
rect 337 946 365 1279
rect 411 946 465 1279
rect 511 946 539 1279
rect 567 918 595 1251
rect 623 946 651 1279
rect 679 918 707 1251
rect 735 946 763 1279
rect 810 918 876 1704
rect 923 1343 951 1676
rect 979 1371 1007 1704
rect 1035 1343 1063 1676
rect 1091 1371 1119 1704
rect 1147 1343 1175 1676
rect 1221 1343 1275 1676
rect 1321 1343 1349 1676
rect 1377 1371 1405 1704
rect 1433 1343 1461 1676
rect 1489 1371 1517 1704
rect 1545 1343 1573 1676
rect 923 1279 1573 1343
rect 923 946 951 1279
rect 979 918 1007 1251
rect 1035 946 1063 1279
rect 1091 918 1119 1251
rect 1147 946 1175 1279
rect 1221 946 1275 1279
rect 1321 946 1349 1279
rect 1377 918 1405 1251
rect 1433 946 1461 1279
rect 1489 918 1517 1251
rect 1545 946 1573 1279
rect 1620 918 1686 1704
rect 0 852 1686 918
rect 0 66 66 852
rect 113 491 141 824
rect 169 519 197 852
rect 225 491 253 824
rect 281 519 309 852
rect 337 491 365 824
rect 411 491 465 824
rect 511 491 539 824
rect 567 519 595 852
rect 623 491 651 824
rect 679 519 707 852
rect 735 491 763 824
rect 113 427 763 491
rect 113 94 141 427
rect 169 66 197 399
rect 225 94 253 427
rect 281 66 309 399
rect 337 94 365 427
rect 411 94 465 427
rect 511 94 539 427
rect 567 66 595 399
rect 623 94 651 427
rect 679 66 707 399
rect 735 94 763 427
rect 810 66 876 852
rect 923 491 951 824
rect 979 519 1007 852
rect 1035 491 1063 824
rect 1091 519 1119 852
rect 1147 491 1175 824
rect 1221 491 1275 824
rect 1321 491 1349 824
rect 1377 519 1405 852
rect 1433 491 1461 824
rect 1489 519 1517 852
rect 1545 491 1573 824
rect 923 427 1573 491
rect 923 94 951 427
rect 979 66 1007 399
rect 1035 94 1063 427
rect 1091 66 1119 399
rect 1147 94 1175 427
rect 1221 94 1275 427
rect 1321 94 1349 427
rect 1377 66 1405 399
rect 1433 94 1461 427
rect 1489 66 1517 399
rect 1545 94 1573 427
rect 1620 66 1686 852
rect 0 0 1686 66
<< obsm2 >>
rect 0 1704 383 1770
rect 0 1620 66 1704
rect 411 1676 465 1770
rect 493 1704 1193 1770
rect 94 1648 782 1676
rect 0 1592 382 1620
rect 0 1508 66 1592
rect 410 1564 466 1648
rect 810 1620 876 1704
rect 1221 1676 1275 1770
rect 1303 1704 1686 1770
rect 904 1648 1592 1676
rect 494 1592 1192 1620
rect 94 1536 782 1564
rect 0 1480 382 1508
rect 0 1396 66 1480
rect 410 1452 466 1536
rect 810 1508 876 1592
rect 1220 1564 1276 1648
rect 1620 1620 1686 1704
rect 1304 1592 1686 1620
rect 904 1536 1592 1564
rect 494 1480 1192 1508
rect 94 1424 782 1452
rect 0 1368 382 1396
rect 0 1366 66 1368
rect 410 1339 466 1424
rect 810 1396 876 1480
rect 1220 1452 1276 1536
rect 1620 1508 1686 1592
rect 1304 1480 1686 1508
rect 904 1424 1592 1452
rect 494 1368 1192 1396
rect 810 1366 876 1368
rect 1220 1339 1276 1424
rect 1620 1396 1686 1480
rect 1304 1368 1686 1396
rect 1620 1366 1686 1368
rect 74 1338 802 1339
rect 884 1338 1612 1339
rect 0 1284 1686 1338
rect 74 1283 802 1284
rect 884 1283 1612 1284
rect 0 1254 66 1256
rect 0 1226 382 1254
rect 0 1142 66 1226
rect 410 1198 466 1283
rect 810 1254 876 1256
rect 494 1226 1192 1254
rect 94 1170 782 1198
rect 0 1114 382 1142
rect 0 1030 66 1114
rect 410 1086 466 1170
rect 810 1142 876 1226
rect 1220 1198 1276 1283
rect 1620 1254 1686 1256
rect 1304 1226 1686 1254
rect 904 1170 1592 1198
rect 494 1114 1192 1142
rect 94 1058 782 1086
rect 0 1002 382 1030
rect 0 918 66 1002
rect 410 974 466 1058
rect 810 1030 876 1114
rect 1220 1086 1276 1170
rect 1620 1142 1686 1226
rect 1304 1114 1686 1142
rect 904 1058 1592 1086
rect 494 1002 1192 1030
rect 94 946 782 974
rect 0 852 383 918
rect 0 768 66 852
rect 411 824 465 946
rect 810 918 876 1002
rect 1220 974 1276 1058
rect 1620 1030 1686 1114
rect 1304 1002 1686 1030
rect 904 946 1592 974
rect 493 852 1193 918
rect 94 796 782 824
rect 0 740 382 768
rect 0 656 66 740
rect 410 712 466 796
rect 810 768 876 852
rect 1221 824 1275 946
rect 1620 918 1686 1002
rect 1303 852 1686 918
rect 904 796 1592 824
rect 494 740 1192 768
rect 94 684 782 712
rect 0 628 382 656
rect 0 544 66 628
rect 410 600 466 684
rect 810 656 876 740
rect 1220 712 1276 796
rect 1620 768 1686 852
rect 1304 740 1686 768
rect 904 684 1592 712
rect 494 628 1192 656
rect 94 572 782 600
rect 0 516 382 544
rect 0 514 66 516
rect 410 487 466 572
rect 810 544 876 628
rect 1220 600 1276 684
rect 1620 656 1686 740
rect 1304 628 1686 656
rect 904 572 1592 600
rect 494 516 1192 544
rect 810 514 876 516
rect 1220 487 1276 572
rect 1620 544 1686 628
rect 1304 516 1686 544
rect 1620 514 1686 516
rect 74 486 802 487
rect 884 486 1612 487
rect 0 432 1686 486
rect 74 431 802 432
rect 884 431 1612 432
rect 0 402 66 404
rect 0 374 382 402
rect 0 290 66 374
rect 410 346 466 431
rect 810 402 876 404
rect 494 374 1192 402
rect 94 318 782 346
rect 0 262 382 290
rect 0 178 66 262
rect 410 234 466 318
rect 810 290 876 374
rect 1220 346 1276 431
rect 1620 402 1686 404
rect 1304 374 1686 402
rect 904 318 1592 346
rect 494 262 1192 290
rect 94 206 782 234
rect 0 150 382 178
rect 0 66 66 150
rect 410 122 466 206
rect 810 178 876 262
rect 1220 234 1276 318
rect 1620 290 1686 374
rect 1304 262 1686 290
rect 904 206 1592 234
rect 494 150 1192 178
rect 94 94 782 122
rect 0 0 383 66
rect 411 0 465 94
rect 810 66 876 150
rect 1220 122 1276 206
rect 1620 178 1686 262
rect 1304 150 1686 178
rect 904 94 1592 122
rect 493 0 1193 66
rect 1221 0 1275 94
rect 1620 66 1686 150
rect 1303 0 1686 66
<< metal3 >>
rect 0 1704 1686 1770
rect 0 918 66 1704
rect 126 1344 186 1644
rect 246 1404 306 1704
rect 405 1344 471 1644
rect 570 1404 630 1704
rect 690 1344 750 1644
rect 126 1278 750 1344
rect 126 978 186 1278
rect 246 918 306 1218
rect 405 978 471 1278
rect 570 918 630 1218
rect 690 978 750 1278
rect 810 918 876 1704
rect 936 1344 996 1644
rect 1056 1404 1116 1704
rect 1215 1344 1281 1644
rect 1380 1404 1440 1704
rect 1500 1344 1560 1644
rect 936 1278 1560 1344
rect 936 978 996 1278
rect 1056 918 1116 1218
rect 1215 978 1281 1278
rect 1380 918 1440 1218
rect 1500 978 1560 1278
rect 1620 918 1686 1704
rect 0 852 1686 918
rect 0 66 66 852
rect 126 492 186 792
rect 246 552 306 852
rect 405 492 471 792
rect 570 552 630 852
rect 690 492 750 792
rect 126 426 750 492
rect 126 126 186 426
rect 246 66 306 366
rect 405 126 471 426
rect 570 66 630 366
rect 690 126 750 426
rect 810 66 876 852
rect 936 492 996 792
rect 1056 552 1116 852
rect 1215 492 1281 792
rect 1380 552 1440 852
rect 1500 492 1560 792
rect 936 426 1560 492
rect 936 126 996 426
rect 1056 66 1116 366
rect 1215 126 1281 426
rect 1380 66 1440 366
rect 1500 126 1560 426
rect 1620 66 1686 852
rect 0 0 1686 66
<< obsm4 >>
rect 74 1396 374 1696
rect 502 1396 802 1696
rect 884 1396 1184 1696
rect 1312 1396 1612 1696
rect 74 926 374 1226
rect 502 926 802 1226
rect 884 926 1184 1226
rect 1312 926 1612 1226
rect 74 544 374 844
rect 502 544 802 844
rect 884 544 1184 844
rect 1312 544 1612 844
rect 74 74 374 374
rect 502 74 802 374
rect 884 74 1184 374
rect 1312 74 1612 374
<< metal5 >>
rect 0 0 1686 1770
<< labels >>
rlabel metal3 s 1620 918 1686 1704 6 C0
port 1 nsew
rlabel metal3 s 1620 66 1686 852 6 C0
port 1 nsew
rlabel metal3 s 1380 1404 1440 1704 6 C0
port 1 nsew
rlabel metal3 s 1380 918 1440 1218 6 C0
port 1 nsew
rlabel metal3 s 1380 552 1440 852 6 C0
port 1 nsew
rlabel metal3 s 1380 66 1440 366 6 C0
port 1 nsew
rlabel metal3 s 1056 1404 1116 1704 6 C0
port 1 nsew
rlabel metal3 s 1056 918 1116 1218 6 C0
port 1 nsew
rlabel metal3 s 1056 552 1116 852 6 C0
port 1 nsew
rlabel metal3 s 1056 66 1116 366 6 C0
port 1 nsew
rlabel metal3 s 810 918 876 1704 6 C0
port 1 nsew
rlabel metal3 s 810 66 876 852 6 C0
port 1 nsew
rlabel metal3 s 570 1404 630 1704 6 C0
port 1 nsew
rlabel metal3 s 570 918 630 1218 6 C0
port 1 nsew
rlabel metal3 s 570 552 630 852 6 C0
port 1 nsew
rlabel metal3 s 570 66 630 366 6 C0
port 1 nsew
rlabel metal3 s 246 1404 306 1704 6 C0
port 1 nsew
rlabel metal3 s 246 918 306 1218 6 C0
port 1 nsew
rlabel metal3 s 246 552 306 852 6 C0
port 1 nsew
rlabel metal3 s 246 66 306 366 6 C0
port 1 nsew
rlabel metal3 s 0 1704 1686 1770 6 C0
port 1 nsew
rlabel metal3 s 0 918 66 1704 6 C0
port 1 nsew
rlabel metal3 s 0 852 1686 918 6 C0
port 1 nsew
rlabel metal3 s 0 66 66 852 6 C0
port 1 nsew
rlabel metal3 s 0 0 1686 66 6 C0
port 1 nsew
rlabel metal3 s 1500 1344 1560 1644 6 C1
port 2 nsew
rlabel metal3 s 1500 978 1560 1278 6 C1
port 2 nsew
rlabel metal3 s 1500 492 1560 792 6 C1
port 2 nsew
rlabel metal3 s 1500 126 1560 426 6 C1
port 2 nsew
rlabel metal3 s 1215 1344 1281 1644 6 C1
port 2 nsew
rlabel metal3 s 1215 978 1281 1278 6 C1
port 2 nsew
rlabel metal3 s 1215 492 1281 792 6 C1
port 2 nsew
rlabel metal3 s 1215 126 1281 426 6 C1
port 2 nsew
rlabel metal3 s 936 1344 996 1644 6 C1
port 2 nsew
rlabel metal3 s 936 1278 1560 1344 6 C1
port 2 nsew
rlabel metal3 s 936 978 996 1278 6 C1
port 2 nsew
rlabel metal3 s 936 492 996 792 6 C1
port 2 nsew
rlabel metal3 s 936 426 1560 492 6 C1
port 2 nsew
rlabel metal3 s 936 126 996 426 6 C1
port 2 nsew
rlabel metal3 s 690 1344 750 1644 6 C1
port 2 nsew
rlabel metal3 s 690 978 750 1278 6 C1
port 2 nsew
rlabel metal3 s 690 492 750 792 6 C1
port 2 nsew
rlabel metal3 s 690 126 750 426 6 C1
port 2 nsew
rlabel metal3 s 405 1344 471 1644 6 C1
port 2 nsew
rlabel metal3 s 405 978 471 1278 6 C1
port 2 nsew
rlabel metal3 s 405 492 471 792 6 C1
port 2 nsew
rlabel metal3 s 405 126 471 426 6 C1
port 2 nsew
rlabel metal3 s 126 1344 186 1644 6 C1
port 2 nsew
rlabel metal3 s 126 1278 750 1344 6 C1
port 2 nsew
rlabel metal3 s 126 978 186 1278 6 C1
port 2 nsew
rlabel metal3 s 126 492 186 792 6 C1
port 2 nsew
rlabel metal3 s 126 426 750 492 6 C1
port 2 nsew
rlabel metal3 s 126 126 186 426 6 C1
port 2 nsew
rlabel metal5 s 0 0 1686 1770 6 M5
port 3 nsew
rlabel pwell s 1179 1269 1189 1279 6 SUB
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 1686 1770
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 135652
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 135072
<< end >>
