magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -76 -26 532 626
<< mvnmos >>
rect 0 0 200 600
rect 256 0 456 600
<< mvndiff >>
rect -50 0 0 600
rect 456 0 506 600
<< poly >>
rect 0 600 200 632
rect 0 -32 200 0
rect 256 600 456 632
rect 256 -32 456 0
<< locali >>
rect -45 -4 -11 538
rect 211 -4 245 538
rect 467 -4 501 538
use hvDFL1sd2_CDNS_52468879185120  hvDFL1sd2_CDNS_52468879185120_0
timestamp 1707688321
transform -1 0 0 0 1 0
box -26 -26 82 626
use hvDFL1sd2_CDNS_52468879185120  hvDFL1sd2_CDNS_52468879185120_1
timestamp 1707688321
transform 1 0 456 0 1 0
box -26 -26 82 626
use hvDFL1sd2_CDNS_52468879185120  hvDFL1sd2_CDNS_52468879185120_2
timestamp 1707688321
transform 1 0 200 0 1 0
box -26 -26 82 626
<< labels >>
flabel comment s -28 267 -28 267 0 FreeSans 300 0 0 0 S
flabel comment s 228 267 228 267 0 FreeSans 300 0 0 0 D
flabel comment s 484 267 484 267 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 85635130
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85633736
<< end >>
