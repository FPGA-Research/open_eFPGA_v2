magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 1 21 827 203
rect 30 -17 64 21
<< locali >>
rect 119 151 157 493
rect 280 215 346 259
rect 400 199 467 325
rect 537 287 618 325
rect 537 199 571 287
rect 667 249 710 325
rect 617 215 710 249
rect 119 59 153 151
rect 667 149 710 215
rect 757 146 801 325
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 19 299 85 527
rect 19 17 85 161
rect 203 367 253 527
rect 291 333 357 485
rect 391 393 425 493
rect 467 435 517 527
rect 559 393 593 493
rect 667 435 717 527
rect 759 393 793 493
rect 391 359 793 393
rect 196 299 357 333
rect 196 161 230 299
rect 196 127 509 161
rect 187 17 253 93
rect 299 51 341 127
rect 475 93 509 127
rect 375 17 441 93
rect 475 59 809 93
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
rlabel locali s 757 146 801 325 6 A1
port 1 nsew signal input
rlabel locali s 667 149 710 215 6 A2
port 2 nsew signal input
rlabel locali s 617 215 710 249 6 A2
port 2 nsew signal input
rlabel locali s 667 249 710 325 6 A2
port 2 nsew signal input
rlabel locali s 537 199 571 287 6 A3
port 3 nsew signal input
rlabel locali s 537 287 618 325 6 A3
port 3 nsew signal input
rlabel locali s 400 199 467 325 6 A4
port 4 nsew signal input
rlabel locali s 280 215 346 259 6 B1
port 5 nsew signal input
rlabel metal1 s 0 -48 828 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1 21 827 203 6 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 866 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 828 592 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 119 59 153 151 6 X
port 10 nsew signal output
rlabel locali s 119 151 157 493 6 X
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 828 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3517434
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3509180
<< end >>
