magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -80 33103 15080 33442
rect -80 28738 290 33103
rect 14636 28738 15080 33103
rect -80 28380 15080 28738
rect -17 25533 15032 27476
<< obsli1 >>
rect 0 25445 14983 33379
rect -41 24648 14983 25445
rect 0 19884 14983 24648
rect -17 19879 14983 19884
rect -41 18589 14983 19879
rect 0 17855 14983 18589
<< obsm1 >>
rect 0 33391 15000 36050
rect -29 28431 15029 33391
rect 0 27189 15029 28431
rect 0 25052 15000 27189
rect -29 19864 15029 25052
rect -29 19560 15000 19864
rect 0 17881 15000 19560
<< obsm2 >>
rect 164 7916 14983 35764
<< metal3 >>
rect 7766 0 9562 2834
<< obsm3 >>
rect 198 2914 14784 39600
rect 198 2834 7686 2914
rect 9642 2834 14784 2914
<< metal4 >>
rect 0 34757 15000 39600
rect 0 13607 254 18600
rect 14746 13607 15000 18600
rect 0 12417 254 13307
rect 14746 12417 15000 13307
rect 0 11247 254 12137
rect 14746 11247 15000 12137
rect 0 10881 15000 10947
rect 0 10225 15000 10821
rect 0 9929 254 10165
rect 14746 9929 15000 10165
rect 0 9273 15000 9869
rect 0 9147 15000 9213
rect 0 7917 254 8847
rect 14746 7917 15000 8847
rect 0 6947 254 7637
rect 14746 6947 15000 7637
rect 0 5977 254 6667
rect 14746 5977 15000 6667
rect 0 4767 15000 5697
rect 0 3557 254 4487
rect 14746 3557 15000 4487
rect 0 2587 193 3277
rect 14807 2587 15000 3277
rect 0 1377 254 2307
rect 14746 1377 15000 2307
rect 0 7 254 1097
rect 14746 7 15000 1097
<< obsm4 >>
rect 193 18680 14807 34220
rect 334 13527 14666 18680
rect 193 13387 14807 13527
rect 334 12337 14666 13387
rect 193 12217 14807 12337
rect 334 11167 14666 12217
rect 193 11027 14807 11167
rect 334 9949 14666 10145
rect 193 8927 14807 9067
rect 334 7837 14666 8927
rect 193 7717 14807 7837
rect 334 6867 14666 7717
rect 193 6747 14807 6867
rect 334 5897 14666 6747
rect 193 5777 14807 5897
rect 193 4567 14807 4687
rect 334 3477 14666 4567
rect 193 3357 14807 3477
rect 273 2507 14727 3357
rect 193 2387 14807 2507
rect 334 1297 14666 2387
rect 193 1177 14807 1297
rect 334 7 14666 1177
<< metal5 >>
rect 0 34757 254 39600
rect 14746 34757 15000 39600
rect 1240 20435 13760 32925
rect 0 13607 254 18597
rect 0 12437 254 13287
rect 0 11267 254 12117
rect 0 9147 254 10947
rect 0 7937 254 8827
rect 0 6968 254 7617
rect 0 5997 254 6647
rect 0 4787 254 5677
rect 0 3577 254 4467
rect 14746 13607 15000 18597
rect 14746 12437 15000 13287
rect 14746 11267 15000 12117
rect 14746 9147 15000 10947
rect 14746 7937 15000 8827
rect 14746 6968 15000 7617
rect 14746 5997 15000 6647
rect 14746 4787 15000 5677
rect 14746 3577 15000 4467
rect 0 2607 193 3257
rect 14807 2607 15000 3257
rect 0 1397 254 2287
rect 0 27 254 1077
rect 14746 1397 15000 2287
rect 14746 27 15000 1077
<< obsm5 >>
rect 574 34437 14426 39600
rect 0 33245 15000 34437
rect 0 20115 920 33245
rect 14080 20115 15000 33245
rect 0 18917 15000 20115
rect 574 3257 14426 18917
rect 513 2607 14487 3257
rect 574 27 14426 2607
<< labels >>
rlabel metal5 s 14746 34757 15000 39600 6 vssio
port 1 nsew ground bidirectional
rlabel metal5 s 14746 4787 15000 5677 6 vssio
port 1 nsew ground bidirectional
rlabel metal5 s 0 34757 254 39600 6 vssio
port 1 nsew ground bidirectional
rlabel metal5 s 0 4787 254 5677 6 vssio
port 1 nsew ground bidirectional
rlabel metal4 s 14746 34757 15000 39600 6 vssio
port 1 nsew ground bidirectional
rlabel metal4 s 14746 4767 15000 5697 6 vssio
port 1 nsew ground bidirectional
rlabel metal4 s 0 34757 254 39600 6 vssio
port 1 nsew ground bidirectional
rlabel metal4 s 0 4767 254 5697 6 vssio
port 1 nsew ground bidirectional
rlabel metal5 s 14746 1397 15000 2287 6 vccd
port 2 nsew power bidirectional
rlabel metal5 s 0 1397 254 2287 6 vccd
port 2 nsew power bidirectional
rlabel metal4 s 14746 1377 15000 2307 6 vccd
port 2 nsew power bidirectional
rlabel metal4 s 0 1377 254 2307 6 vccd
port 2 nsew power bidirectional
rlabel metal5 s 14746 12437 15000 13287 6 vddio_q
port 3 nsew power bidirectional
rlabel metal5 s 0 12437 254 13287 6 vddio_q
port 3 nsew power bidirectional
rlabel metal4 s 14746 12417 15000 13307 6 vddio_q
port 3 nsew power bidirectional
rlabel metal4 s 0 12417 254 13307 6 vddio_q
port 3 nsew power bidirectional
rlabel metal5 s 14746 9147 15000 10947 6 vssa
port 4 nsew ground bidirectional
rlabel metal5 s 14746 6968 15000 7617 6 vssa
port 4 nsew ground bidirectional
rlabel metal5 s 0 9147 254 10947 6 vssa
port 4 nsew ground bidirectional
rlabel metal5 s 0 6968 254 7617 6 vssa
port 4 nsew ground bidirectional
rlabel metal4 s 14746 6947 15000 7637 6 vssa
port 4 nsew ground bidirectional
rlabel metal4 s 0 9147 15000 9213 6 vssa
port 4 nsew ground bidirectional
rlabel metal4 s 0 10881 15000 10947 6 vssa
port 4 nsew ground bidirectional
rlabel metal4 s 14746 9929 15000 10165 6 vssa
port 4 nsew ground bidirectional
rlabel metal4 s 0 9929 254 10165 6 vssa
port 4 nsew ground bidirectional
rlabel metal4 s 0 6947 254 7637 6 vssa
port 4 nsew ground bidirectional
rlabel metal5 s 14746 13607 15000 18597 6 vddio
port 5 nsew power bidirectional
rlabel metal5 s 14746 3577 15000 4467 6 vddio
port 5 nsew power bidirectional
rlabel metal5 s 0 13607 254 18597 6 vddio
port 5 nsew power bidirectional
rlabel metal5 s 0 3577 254 4467 6 vddio
port 5 nsew power bidirectional
rlabel metal4 s 14746 3557 15000 4487 6 vddio
port 5 nsew power bidirectional
rlabel metal4 s 14746 13607 15000 18600 6 vddio
port 5 nsew power bidirectional
rlabel metal4 s 0 3557 254 4487 6 vddio
port 5 nsew power bidirectional
rlabel metal4 s 0 13607 254 18600 6 vddio
port 5 nsew power bidirectional
rlabel metal5 s 14746 27 15000 1077 6 vcchib
port 6 nsew power bidirectional
rlabel metal5 s 0 27 254 1077 6 vcchib
port 6 nsew power bidirectional
rlabel metal4 s 14746 7 15000 1097 6 vcchib
port 6 nsew power bidirectional
rlabel metal4 s 0 7 254 1097 6 vcchib
port 6 nsew power bidirectional
rlabel metal5 s 14746 5997 15000 6647 6 vswitch
port 7 nsew power bidirectional
rlabel metal5 s 0 5997 254 6647 6 vswitch
port 7 nsew power bidirectional
rlabel metal4 s 14746 5977 15000 6667 6 vswitch
port 7 nsew power bidirectional
rlabel metal4 s 0 5977 254 6667 6 vswitch
port 7 nsew power bidirectional
rlabel metal5 s 14746 11267 15000 12117 6 vssio_q
port 8 nsew ground bidirectional
rlabel metal5 s 0 11267 254 12117 6 vssio_q
port 8 nsew ground bidirectional
rlabel metal4 s 14746 11247 15000 12137 6 vssio_q
port 8 nsew ground bidirectional
rlabel metal4 s 0 11247 254 12137 6 vssio_q
port 8 nsew ground bidirectional
rlabel metal5 s 14807 2607 15000 3257 6 vdda
port 9 nsew power bidirectional
rlabel metal5 s 0 2607 193 3257 6 vdda
port 9 nsew power bidirectional
rlabel metal4 s 14807 2587 15000 3277 6 vdda
port 9 nsew power bidirectional
rlabel metal4 s 0 2587 193 3277 6 vdda
port 9 nsew power bidirectional
rlabel metal5 s 14746 7937 15000 8827 6 vssd
port 10 nsew ground bidirectional
rlabel metal5 s 0 7937 254 8827 6 vssd
port 10 nsew ground bidirectional
rlabel metal4 s 14746 7917 15000 8847 6 vssd
port 10 nsew ground bidirectional
rlabel metal4 s 0 7917 254 8847 6 vssd
port 10 nsew ground bidirectional
rlabel metal5 s 1240 20435 13760 32925 6 pad
port 11 nsew signal bidirectional
rlabel metal4 s 0 9273 15000 9869 6 amuxbus_b
port 12 nsew signal bidirectional
rlabel metal4 s 0 10225 15000 10821 6 amuxbus_a
port 13 nsew signal bidirectional
rlabel metal3 s 7766 0 9562 2834 6 pad_core
port 14 nsew signal bidirectional
rlabel metal4 s 0 4767 15000 5697 6 vssio
port 15 nsew ground bidirectional
rlabel metal4 s 0 34757 15000 39600 6 vssio
port 16 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 39600
string LEFclass BLOCK
string LEFsymmetry R90
string LEFview TRUE
string GDS_END 16732744
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 14492232
<< end >>
