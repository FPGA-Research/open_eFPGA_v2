magic
tech sky130B
timestamp 1707688321
<< viali >>
rect 0 0 197 197
<< metal1 >>
rect -6 197 203 200
rect -6 0 0 197
rect 197 0 203 197
rect -6 -3 203 0
<< properties >>
string GDS_END 86922910
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86920474
<< end >>
