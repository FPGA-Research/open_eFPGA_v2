magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 107 157 527 203
rect 1 21 735 157
rect 30 -17 64 21
<< scnmos >>
rect 81 47 111 131
rect 191 47 227 177
rect 387 47 423 177
rect 518 47 548 131
rect 604 47 634 131
<< scpmoshvt >>
rect 81 297 111 497
rect 191 333 227 497
rect 387 333 423 497
rect 518 297 548 497
rect 604 297 634 497
<< ndiff >>
rect 133 131 191 177
rect 27 104 81 131
rect 27 70 36 104
rect 70 70 81 104
rect 27 47 81 70
rect 111 97 191 131
rect 111 63 133 97
rect 167 63 191 97
rect 111 47 191 63
rect 227 104 280 177
rect 227 70 238 104
rect 272 70 280 104
rect 227 47 280 70
rect 334 104 387 177
rect 334 70 342 104
rect 376 70 387 104
rect 334 47 387 70
rect 423 131 501 177
rect 423 97 518 131
rect 423 63 451 97
rect 485 63 518 97
rect 423 47 518 63
rect 548 104 604 131
rect 548 70 559 104
rect 593 70 604 104
rect 548 47 604 70
rect 634 104 709 131
rect 634 70 664 104
rect 698 70 709 104
rect 634 47 709 70
<< pdiff >>
rect 27 478 81 497
rect 27 444 36 478
rect 70 444 81 478
rect 27 410 81 444
rect 27 376 36 410
rect 70 376 81 410
rect 27 297 81 376
rect 111 478 191 497
rect 111 444 136 478
rect 170 444 191 478
rect 111 410 191 444
rect 111 376 136 410
rect 170 376 191 410
rect 111 333 191 376
rect 227 478 280 497
rect 227 444 238 478
rect 272 444 280 478
rect 227 410 280 444
rect 227 376 238 410
rect 272 376 280 410
rect 227 333 280 376
rect 334 478 387 497
rect 334 444 342 478
rect 376 444 387 478
rect 334 410 387 444
rect 334 376 342 410
rect 376 376 387 410
rect 334 333 387 376
rect 423 478 518 497
rect 423 444 453 478
rect 487 444 518 478
rect 423 410 518 444
rect 423 376 453 410
rect 487 376 518 410
rect 423 333 518 376
rect 111 297 161 333
rect 468 297 518 333
rect 548 478 604 497
rect 548 444 559 478
rect 593 444 604 478
rect 548 410 604 444
rect 548 376 559 410
rect 593 376 604 410
rect 548 297 604 376
rect 634 478 709 497
rect 634 444 664 478
rect 698 444 709 478
rect 634 410 709 444
rect 634 376 664 410
rect 698 376 709 410
rect 634 297 709 376
<< ndiffc >>
rect 36 70 70 104
rect 133 63 167 97
rect 238 70 272 104
rect 342 70 376 104
rect 451 63 485 97
rect 559 70 593 104
rect 664 70 698 104
<< pdiffc >>
rect 36 444 70 478
rect 36 376 70 410
rect 136 444 170 478
rect 136 376 170 410
rect 238 444 272 478
rect 238 376 272 410
rect 342 444 376 478
rect 342 376 376 410
rect 453 444 487 478
rect 453 376 487 410
rect 559 444 593 478
rect 559 376 593 410
rect 664 444 698 478
rect 664 376 698 410
<< poly >>
rect 81 497 111 523
rect 191 497 227 523
rect 387 497 423 523
rect 518 497 548 523
rect 604 497 634 523
rect 81 261 111 297
rect 46 259 111 261
rect 191 259 227 333
rect 387 259 423 333
rect 518 259 548 297
rect 604 259 634 297
rect 46 249 112 259
rect 46 215 62 249
rect 96 215 112 249
rect 46 205 112 215
rect 161 249 227 259
rect 161 215 177 249
rect 211 215 227 249
rect 161 205 227 215
rect 307 249 441 259
rect 307 215 323 249
rect 357 215 391 249
rect 425 215 441 249
rect 307 205 441 215
rect 502 249 634 259
rect 502 215 518 249
rect 552 215 634 249
rect 502 205 634 215
rect 46 203 111 205
rect 81 131 111 203
rect 191 177 227 205
rect 387 177 423 205
rect 518 131 548 205
rect 604 131 634 205
rect 81 21 111 47
rect 191 21 227 47
rect 387 21 423 47
rect 518 21 548 47
rect 604 21 634 47
<< polycont >>
rect 62 215 96 249
rect 177 215 211 249
rect 323 215 357 249
rect 391 215 425 249
rect 518 215 552 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 17 478 86 493
rect 17 444 36 478
rect 70 444 86 478
rect 17 410 86 444
rect 17 376 36 410
rect 70 376 86 410
rect 17 326 86 376
rect 120 478 186 527
rect 120 444 136 478
rect 170 444 186 478
rect 120 410 186 444
rect 120 376 136 410
rect 170 376 186 410
rect 120 360 186 376
rect 222 478 288 493
rect 222 444 238 478
rect 272 444 288 478
rect 222 410 288 444
rect 222 376 238 410
rect 272 376 288 410
rect 222 360 288 376
rect 17 292 211 326
rect 17 249 112 258
rect 17 215 62 249
rect 96 215 112 249
rect 146 249 211 292
rect 146 215 177 249
rect 146 181 211 215
rect 17 147 211 181
rect 254 251 288 360
rect 326 478 392 493
rect 326 444 342 478
rect 376 444 392 478
rect 326 410 392 444
rect 326 376 342 410
rect 376 376 392 410
rect 326 326 392 376
rect 426 478 509 527
rect 426 444 453 478
rect 487 444 509 478
rect 426 410 509 444
rect 426 376 453 410
rect 487 376 509 410
rect 426 360 509 376
rect 543 478 630 493
rect 543 444 559 478
rect 593 444 630 478
rect 543 410 630 444
rect 543 376 559 410
rect 593 376 630 410
rect 326 292 509 326
rect 254 249 441 251
rect 254 215 323 249
rect 357 215 391 249
rect 425 215 441 249
rect 475 249 509 292
rect 543 305 630 376
rect 664 478 719 527
rect 698 444 719 478
rect 664 410 719 444
rect 698 376 719 410
rect 664 325 719 376
rect 543 284 636 305
rect 475 215 518 249
rect 552 215 568 249
rect 17 104 83 147
rect 254 120 288 215
rect 475 181 509 215
rect 602 189 636 284
rect 17 70 36 104
rect 70 70 83 104
rect 17 54 83 70
rect 117 97 183 113
rect 117 63 133 97
rect 167 63 183 97
rect 117 17 183 63
rect 232 104 288 120
rect 232 70 238 104
rect 272 70 288 104
rect 232 54 288 70
rect 326 147 509 181
rect 593 156 636 189
rect 326 104 392 147
rect 593 128 630 156
rect 326 70 342 104
rect 376 70 392 104
rect 326 54 392 70
rect 433 97 507 113
rect 433 63 451 97
rect 485 63 507 97
rect 433 17 507 63
rect 541 104 630 128
rect 541 70 559 104
rect 593 70 630 104
rect 541 54 630 70
rect 664 104 719 129
rect 698 70 719 104
rect 664 17 719 70
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel locali s 30 221 64 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 586 85 620 119 0 FreeSans 400 0 0 0 X
port 6 nsew signal output
flabel locali s 586 425 620 459 0 FreeSans 400 0 0 0 X
port 6 nsew signal output
flabel locali s 586 357 620 391 0 FreeSans 400 0 0 0 X
port 6 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 clkdlybuf4s18_2
rlabel metal1 s 0 -48 736 48 1 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 496 736 592 1 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_END 3255508
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3249398
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 13.600 18.400 13.600 
<< end >>
