magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect 0 0 3132 494
<< mvpmos >>
rect 66 275 3066 375
rect 66 119 3066 219
<< mvpdiff >>
rect 66 420 3066 428
rect 66 386 78 420
rect 112 386 146 420
rect 180 386 214 420
rect 248 386 282 420
rect 316 386 350 420
rect 384 386 418 420
rect 452 386 486 420
rect 520 386 554 420
rect 588 386 622 420
rect 656 386 690 420
rect 724 386 758 420
rect 792 386 826 420
rect 860 386 894 420
rect 928 386 962 420
rect 996 386 1030 420
rect 1064 386 1098 420
rect 1132 386 1166 420
rect 1200 386 1234 420
rect 1268 386 1302 420
rect 1336 386 1370 420
rect 1404 386 1438 420
rect 1472 386 1506 420
rect 1540 386 1574 420
rect 1608 386 1642 420
rect 1676 386 1710 420
rect 1744 386 1778 420
rect 1812 386 1846 420
rect 1880 386 1914 420
rect 1948 386 1982 420
rect 2016 386 2050 420
rect 2084 386 2118 420
rect 2152 386 2186 420
rect 2220 386 2254 420
rect 2288 386 2322 420
rect 2356 386 2390 420
rect 2424 386 2458 420
rect 2492 386 2526 420
rect 2560 386 2594 420
rect 2628 386 2662 420
rect 2696 386 2730 420
rect 2764 386 2798 420
rect 2832 386 2866 420
rect 2900 386 2934 420
rect 2968 386 3002 420
rect 3036 386 3066 420
rect 66 375 3066 386
rect 66 264 3066 275
rect 66 230 78 264
rect 112 230 146 264
rect 180 230 214 264
rect 248 230 282 264
rect 316 230 350 264
rect 384 230 418 264
rect 452 230 486 264
rect 520 230 554 264
rect 588 230 622 264
rect 656 230 690 264
rect 724 230 758 264
rect 792 230 826 264
rect 860 230 894 264
rect 928 230 962 264
rect 996 230 1030 264
rect 1064 230 1098 264
rect 1132 230 1166 264
rect 1200 230 1234 264
rect 1268 230 1302 264
rect 1336 230 1370 264
rect 1404 230 1438 264
rect 1472 230 1506 264
rect 1540 230 1574 264
rect 1608 230 1642 264
rect 1676 230 1710 264
rect 1744 230 1778 264
rect 1812 230 1846 264
rect 1880 230 1914 264
rect 1948 230 1982 264
rect 2016 230 2050 264
rect 2084 230 2118 264
rect 2152 230 2186 264
rect 2220 230 2254 264
rect 2288 230 2322 264
rect 2356 230 2390 264
rect 2424 230 2458 264
rect 2492 230 2526 264
rect 2560 230 2594 264
rect 2628 230 2662 264
rect 2696 230 2730 264
rect 2764 230 2798 264
rect 2832 230 2866 264
rect 2900 230 2934 264
rect 2968 230 3002 264
rect 3036 230 3066 264
rect 66 219 3066 230
rect 66 108 3066 119
rect 66 74 78 108
rect 112 74 146 108
rect 180 74 214 108
rect 248 74 282 108
rect 316 74 350 108
rect 384 74 418 108
rect 452 74 486 108
rect 520 74 554 108
rect 588 74 622 108
rect 656 74 690 108
rect 724 74 758 108
rect 792 74 826 108
rect 860 74 894 108
rect 928 74 962 108
rect 996 74 1030 108
rect 1064 74 1098 108
rect 1132 74 1166 108
rect 1200 74 1234 108
rect 1268 74 1302 108
rect 1336 74 1370 108
rect 1404 74 1438 108
rect 1472 74 1506 108
rect 1540 74 1574 108
rect 1608 74 1642 108
rect 1676 74 1710 108
rect 1744 74 1778 108
rect 1812 74 1846 108
rect 1880 74 1914 108
rect 1948 74 1982 108
rect 2016 74 2050 108
rect 2084 74 2118 108
rect 2152 74 2186 108
rect 2220 74 2254 108
rect 2288 74 2322 108
rect 2356 74 2390 108
rect 2424 74 2458 108
rect 2492 74 2526 108
rect 2560 74 2594 108
rect 2628 74 2662 108
rect 2696 74 2730 108
rect 2764 74 2798 108
rect 2832 74 2866 108
rect 2900 74 2934 108
rect 2968 74 3002 108
rect 3036 74 3066 108
rect 66 66 3066 74
<< mvpdiffc >>
rect 78 386 112 420
rect 146 386 180 420
rect 214 386 248 420
rect 282 386 316 420
rect 350 386 384 420
rect 418 386 452 420
rect 486 386 520 420
rect 554 386 588 420
rect 622 386 656 420
rect 690 386 724 420
rect 758 386 792 420
rect 826 386 860 420
rect 894 386 928 420
rect 962 386 996 420
rect 1030 386 1064 420
rect 1098 386 1132 420
rect 1166 386 1200 420
rect 1234 386 1268 420
rect 1302 386 1336 420
rect 1370 386 1404 420
rect 1438 386 1472 420
rect 1506 386 1540 420
rect 1574 386 1608 420
rect 1642 386 1676 420
rect 1710 386 1744 420
rect 1778 386 1812 420
rect 1846 386 1880 420
rect 1914 386 1948 420
rect 1982 386 2016 420
rect 2050 386 2084 420
rect 2118 386 2152 420
rect 2186 386 2220 420
rect 2254 386 2288 420
rect 2322 386 2356 420
rect 2390 386 2424 420
rect 2458 386 2492 420
rect 2526 386 2560 420
rect 2594 386 2628 420
rect 2662 386 2696 420
rect 2730 386 2764 420
rect 2798 386 2832 420
rect 2866 386 2900 420
rect 2934 386 2968 420
rect 3002 386 3036 420
rect 78 230 112 264
rect 146 230 180 264
rect 214 230 248 264
rect 282 230 316 264
rect 350 230 384 264
rect 418 230 452 264
rect 486 230 520 264
rect 554 230 588 264
rect 622 230 656 264
rect 690 230 724 264
rect 758 230 792 264
rect 826 230 860 264
rect 894 230 928 264
rect 962 230 996 264
rect 1030 230 1064 264
rect 1098 230 1132 264
rect 1166 230 1200 264
rect 1234 230 1268 264
rect 1302 230 1336 264
rect 1370 230 1404 264
rect 1438 230 1472 264
rect 1506 230 1540 264
rect 1574 230 1608 264
rect 1642 230 1676 264
rect 1710 230 1744 264
rect 1778 230 1812 264
rect 1846 230 1880 264
rect 1914 230 1948 264
rect 1982 230 2016 264
rect 2050 230 2084 264
rect 2118 230 2152 264
rect 2186 230 2220 264
rect 2254 230 2288 264
rect 2322 230 2356 264
rect 2390 230 2424 264
rect 2458 230 2492 264
rect 2526 230 2560 264
rect 2594 230 2628 264
rect 2662 230 2696 264
rect 2730 230 2764 264
rect 2798 230 2832 264
rect 2866 230 2900 264
rect 2934 230 2968 264
rect 3002 230 3036 264
rect 78 74 112 108
rect 146 74 180 108
rect 214 74 248 108
rect 282 74 316 108
rect 350 74 384 108
rect 418 74 452 108
rect 486 74 520 108
rect 554 74 588 108
rect 622 74 656 108
rect 690 74 724 108
rect 758 74 792 108
rect 826 74 860 108
rect 894 74 928 108
rect 962 74 996 108
rect 1030 74 1064 108
rect 1098 74 1132 108
rect 1166 74 1200 108
rect 1234 74 1268 108
rect 1302 74 1336 108
rect 1370 74 1404 108
rect 1438 74 1472 108
rect 1506 74 1540 108
rect 1574 74 1608 108
rect 1642 74 1676 108
rect 1710 74 1744 108
rect 1778 74 1812 108
rect 1846 74 1880 108
rect 1914 74 1948 108
rect 1982 74 2016 108
rect 2050 74 2084 108
rect 2118 74 2152 108
rect 2186 74 2220 108
rect 2254 74 2288 108
rect 2322 74 2356 108
rect 2390 74 2424 108
rect 2458 74 2492 108
rect 2526 74 2560 108
rect 2594 74 2628 108
rect 2662 74 2696 108
rect 2730 74 2764 108
rect 2798 74 2832 108
rect 2866 74 2900 108
rect 2934 74 2968 108
rect 3002 74 3036 108
<< poly >>
rect 3092 410 3172 426
rect 3092 376 3115 410
rect 3149 376 3172 410
rect 3092 375 3172 376
rect 40 275 66 375
rect 3066 342 3172 375
rect 3066 308 3115 342
rect 3149 308 3172 342
rect 3066 275 3172 308
rect 40 119 66 219
rect 3066 187 3172 219
rect 3066 153 3115 187
rect 3149 153 3172 187
rect 3066 119 3172 153
rect 3092 85 3115 119
rect 3149 85 3172 119
rect 3092 69 3172 85
<< polycont >>
rect 3115 376 3149 410
rect 3115 308 3149 342
rect 3115 153 3149 187
rect 3115 85 3149 119
<< locali >>
rect 112 386 134 420
rect 180 386 206 420
rect 248 386 278 420
rect 316 386 350 420
rect 384 386 418 420
rect 456 386 486 420
rect 528 386 554 420
rect 600 386 622 420
rect 672 386 690 420
rect 744 386 758 420
rect 816 386 826 420
rect 888 386 894 420
rect 960 386 962 420
rect 996 386 998 420
rect 1064 386 1070 420
rect 1132 386 1142 420
rect 1200 386 1214 420
rect 1268 386 1286 420
rect 1336 386 1358 420
rect 1404 386 1430 420
rect 1472 386 1502 420
rect 1540 386 1574 420
rect 1608 386 1642 420
rect 1680 386 1710 420
rect 1752 386 1778 420
rect 1824 386 1846 420
rect 1896 386 1914 420
rect 1968 386 1982 420
rect 2040 386 2050 420
rect 2112 386 2118 420
rect 2184 386 2186 420
rect 2220 386 2222 420
rect 2288 386 2294 420
rect 2356 386 2366 420
rect 2424 386 2438 420
rect 2492 386 2510 420
rect 2560 386 2582 420
rect 2628 386 2654 420
rect 2696 386 2726 420
rect 2764 386 2798 420
rect 2832 386 2866 420
rect 2904 386 2934 420
rect 2976 386 3002 420
rect 3048 386 3052 420
rect 3108 410 3156 426
rect 3108 376 3115 410
rect 3149 376 3156 410
rect 3108 342 3156 376
rect 3108 338 3115 342
rect 3012 335 3115 338
rect 3046 301 3084 335
rect 3149 308 3156 342
rect 3118 301 3156 308
rect 3012 298 3156 301
rect 3108 292 3156 298
rect 62 230 78 264
rect 112 230 146 264
rect 185 230 214 264
rect 258 230 282 264
rect 331 230 350 264
rect 404 230 418 264
rect 477 230 486 264
rect 550 230 554 264
rect 588 230 589 264
rect 656 230 662 264
rect 724 230 735 264
rect 792 230 808 264
rect 860 230 881 264
rect 928 230 954 264
rect 996 230 1027 264
rect 1064 230 1098 264
rect 1134 230 1166 264
rect 1207 230 1234 264
rect 1280 230 1302 264
rect 1353 230 1370 264
rect 1426 230 1438 264
rect 1499 230 1506 264
rect 1572 230 1574 264
rect 1608 230 1610 264
rect 1676 230 1682 264
rect 1744 230 1754 264
rect 1812 230 1826 264
rect 1880 230 1898 264
rect 1948 230 1970 264
rect 2016 230 2042 264
rect 2084 230 2114 264
rect 2152 230 2186 264
rect 2220 230 2254 264
rect 2292 230 2322 264
rect 2364 230 2390 264
rect 2436 230 2458 264
rect 2508 230 2526 264
rect 2580 230 2594 264
rect 2652 230 2662 264
rect 2724 230 2730 264
rect 2796 230 2798 264
rect 2832 230 2834 264
rect 2900 230 2906 264
rect 2968 230 3002 264
rect 3036 230 3052 264
rect 3108 194 3156 203
rect 3026 187 3156 194
rect 3026 186 3115 187
rect 3026 152 3038 186
rect 3072 152 3110 186
rect 3149 153 3156 187
rect 3144 152 3156 153
rect 3026 143 3156 152
rect 3108 119 3156 143
rect 112 74 134 108
rect 180 74 206 108
rect 248 74 278 108
rect 316 74 350 108
rect 384 74 418 108
rect 456 74 486 108
rect 528 74 554 108
rect 600 74 622 108
rect 672 74 690 108
rect 744 74 758 108
rect 816 74 826 108
rect 888 74 894 108
rect 960 74 962 108
rect 996 74 998 108
rect 1064 74 1070 108
rect 1132 74 1142 108
rect 1200 74 1214 108
rect 1268 74 1286 108
rect 1336 74 1358 108
rect 1404 74 1430 108
rect 1472 74 1502 108
rect 1540 74 1574 108
rect 1608 74 1642 108
rect 1680 74 1710 108
rect 1752 74 1778 108
rect 1824 74 1846 108
rect 1896 74 1914 108
rect 1968 74 1982 108
rect 2040 74 2050 108
rect 2112 74 2118 108
rect 2184 74 2186 108
rect 2220 74 2222 108
rect 2288 74 2294 108
rect 2356 74 2366 108
rect 2424 74 2438 108
rect 2492 74 2510 108
rect 2560 74 2582 108
rect 2628 74 2654 108
rect 2696 74 2726 108
rect 2764 74 2798 108
rect 2832 74 2866 108
rect 2904 74 2934 108
rect 2976 74 3002 108
rect 3048 74 3052 108
rect 3108 85 3115 119
rect 3149 85 3156 119
rect 3108 69 3156 85
<< viali >>
rect 62 386 78 420
rect 78 386 96 420
rect 134 386 146 420
rect 146 386 168 420
rect 206 386 214 420
rect 214 386 240 420
rect 278 386 282 420
rect 282 386 312 420
rect 350 386 384 420
rect 422 386 452 420
rect 452 386 456 420
rect 494 386 520 420
rect 520 386 528 420
rect 566 386 588 420
rect 588 386 600 420
rect 638 386 656 420
rect 656 386 672 420
rect 710 386 724 420
rect 724 386 744 420
rect 782 386 792 420
rect 792 386 816 420
rect 854 386 860 420
rect 860 386 888 420
rect 926 386 928 420
rect 928 386 960 420
rect 998 386 1030 420
rect 1030 386 1032 420
rect 1070 386 1098 420
rect 1098 386 1104 420
rect 1142 386 1166 420
rect 1166 386 1176 420
rect 1214 386 1234 420
rect 1234 386 1248 420
rect 1286 386 1302 420
rect 1302 386 1320 420
rect 1358 386 1370 420
rect 1370 386 1392 420
rect 1430 386 1438 420
rect 1438 386 1464 420
rect 1502 386 1506 420
rect 1506 386 1536 420
rect 1574 386 1608 420
rect 1646 386 1676 420
rect 1676 386 1680 420
rect 1718 386 1744 420
rect 1744 386 1752 420
rect 1790 386 1812 420
rect 1812 386 1824 420
rect 1862 386 1880 420
rect 1880 386 1896 420
rect 1934 386 1948 420
rect 1948 386 1968 420
rect 2006 386 2016 420
rect 2016 386 2040 420
rect 2078 386 2084 420
rect 2084 386 2112 420
rect 2150 386 2152 420
rect 2152 386 2184 420
rect 2222 386 2254 420
rect 2254 386 2256 420
rect 2294 386 2322 420
rect 2322 386 2328 420
rect 2366 386 2390 420
rect 2390 386 2400 420
rect 2438 386 2458 420
rect 2458 386 2472 420
rect 2510 386 2526 420
rect 2526 386 2544 420
rect 2582 386 2594 420
rect 2594 386 2616 420
rect 2654 386 2662 420
rect 2662 386 2688 420
rect 2726 386 2730 420
rect 2730 386 2760 420
rect 2798 386 2832 420
rect 2870 386 2900 420
rect 2900 386 2904 420
rect 2942 386 2968 420
rect 2968 386 2976 420
rect 3014 386 3036 420
rect 3036 386 3048 420
rect 3012 301 3046 335
rect 3084 308 3115 335
rect 3115 308 3118 335
rect 3084 301 3118 308
rect 78 230 112 264
rect 151 230 180 264
rect 180 230 185 264
rect 224 230 248 264
rect 248 230 258 264
rect 297 230 316 264
rect 316 230 331 264
rect 370 230 384 264
rect 384 230 404 264
rect 443 230 452 264
rect 452 230 477 264
rect 516 230 520 264
rect 520 230 550 264
rect 589 230 622 264
rect 622 230 623 264
rect 662 230 690 264
rect 690 230 696 264
rect 735 230 758 264
rect 758 230 769 264
rect 808 230 826 264
rect 826 230 842 264
rect 881 230 894 264
rect 894 230 915 264
rect 954 230 962 264
rect 962 230 988 264
rect 1027 230 1030 264
rect 1030 230 1061 264
rect 1100 230 1132 264
rect 1132 230 1134 264
rect 1173 230 1200 264
rect 1200 230 1207 264
rect 1246 230 1268 264
rect 1268 230 1280 264
rect 1319 230 1336 264
rect 1336 230 1353 264
rect 1392 230 1404 264
rect 1404 230 1426 264
rect 1465 230 1472 264
rect 1472 230 1499 264
rect 1538 230 1540 264
rect 1540 230 1572 264
rect 1610 230 1642 264
rect 1642 230 1644 264
rect 1682 230 1710 264
rect 1710 230 1716 264
rect 1754 230 1778 264
rect 1778 230 1788 264
rect 1826 230 1846 264
rect 1846 230 1860 264
rect 1898 230 1914 264
rect 1914 230 1932 264
rect 1970 230 1982 264
rect 1982 230 2004 264
rect 2042 230 2050 264
rect 2050 230 2076 264
rect 2114 230 2118 264
rect 2118 230 2148 264
rect 2186 230 2220 264
rect 2258 230 2288 264
rect 2288 230 2292 264
rect 2330 230 2356 264
rect 2356 230 2364 264
rect 2402 230 2424 264
rect 2424 230 2436 264
rect 2474 230 2492 264
rect 2492 230 2508 264
rect 2546 230 2560 264
rect 2560 230 2580 264
rect 2618 230 2628 264
rect 2628 230 2652 264
rect 2690 230 2696 264
rect 2696 230 2724 264
rect 2762 230 2764 264
rect 2764 230 2796 264
rect 2834 230 2866 264
rect 2866 230 2868 264
rect 2906 230 2934 264
rect 2934 230 2940 264
rect 3038 152 3072 186
rect 3110 153 3115 186
rect 3115 153 3144 186
rect 3110 152 3144 153
rect 62 74 78 108
rect 78 74 96 108
rect 134 74 146 108
rect 146 74 168 108
rect 206 74 214 108
rect 214 74 240 108
rect 278 74 282 108
rect 282 74 312 108
rect 350 74 384 108
rect 422 74 452 108
rect 452 74 456 108
rect 494 74 520 108
rect 520 74 528 108
rect 566 74 588 108
rect 588 74 600 108
rect 638 74 656 108
rect 656 74 672 108
rect 710 74 724 108
rect 724 74 744 108
rect 782 74 792 108
rect 792 74 816 108
rect 854 74 860 108
rect 860 74 888 108
rect 926 74 928 108
rect 928 74 960 108
rect 998 74 1030 108
rect 1030 74 1032 108
rect 1070 74 1098 108
rect 1098 74 1104 108
rect 1142 74 1166 108
rect 1166 74 1176 108
rect 1214 74 1234 108
rect 1234 74 1248 108
rect 1286 74 1302 108
rect 1302 74 1320 108
rect 1358 74 1370 108
rect 1370 74 1392 108
rect 1430 74 1438 108
rect 1438 74 1464 108
rect 1502 74 1506 108
rect 1506 74 1536 108
rect 1574 74 1608 108
rect 1646 74 1676 108
rect 1676 74 1680 108
rect 1718 74 1744 108
rect 1744 74 1752 108
rect 1790 74 1812 108
rect 1812 74 1824 108
rect 1862 74 1880 108
rect 1880 74 1896 108
rect 1934 74 1948 108
rect 1948 74 1968 108
rect 2006 74 2016 108
rect 2016 74 2040 108
rect 2078 74 2084 108
rect 2084 74 2112 108
rect 2150 74 2152 108
rect 2152 74 2184 108
rect 2222 74 2254 108
rect 2254 74 2256 108
rect 2294 74 2322 108
rect 2322 74 2328 108
rect 2366 74 2390 108
rect 2390 74 2400 108
rect 2438 74 2458 108
rect 2458 74 2472 108
rect 2510 74 2526 108
rect 2526 74 2544 108
rect 2582 74 2594 108
rect 2594 74 2616 108
rect 2654 74 2662 108
rect 2662 74 2688 108
rect 2726 74 2730 108
rect 2730 74 2760 108
rect 2798 74 2832 108
rect 2870 74 2900 108
rect 2900 74 2904 108
rect 2942 74 2968 108
rect 2968 74 2976 108
rect 3014 74 3036 108
rect 3036 74 3048 108
<< metal1 >>
rect 44 461 3318 507
tri 3113 436 3138 461 ne
rect 50 420 3060 426
rect 50 386 62 420
rect 96 386 134 420
rect 168 386 206 420
rect 240 386 278 420
rect 312 386 350 420
rect 384 386 422 420
rect 456 386 494 420
rect 528 386 566 420
rect 600 386 638 420
rect 672 386 710 420
rect 744 386 782 420
rect 816 386 854 420
rect 888 386 926 420
rect 960 386 998 420
rect 1032 386 1070 420
rect 1104 386 1142 420
rect 1176 386 1214 420
rect 1248 386 1286 420
rect 1320 386 1358 420
rect 1392 386 1430 420
rect 1464 386 1502 420
rect 1536 386 1574 420
rect 1608 386 1646 420
rect 1680 386 1718 420
rect 1752 386 1790 420
rect 1824 386 1862 420
rect 1896 386 1934 420
rect 1968 386 2006 420
rect 2040 386 2078 420
rect 2112 386 2150 420
rect 2184 386 2222 420
rect 2256 386 2294 420
rect 2328 386 2366 420
rect 2400 386 2438 420
rect 2472 386 2510 420
rect 2544 386 2582 420
rect 2616 386 2654 420
rect 2688 386 2726 420
rect 2760 386 2798 420
rect 2832 386 2870 420
rect 2904 386 2942 420
rect 2976 386 3014 420
rect 3048 386 3060 420
rect 50 380 3060 386
tri 3112 344 3138 370 se
rect 3138 344 3190 461
tri 3190 436 3215 461 nw
rect 3000 335 3034 344
rect 3086 335 3098 344
rect 3000 301 3012 335
rect 3000 292 3034 301
rect 3086 292 3098 301
rect 3150 292 3190 344
rect 66 264 2952 270
rect 66 230 78 264
rect 112 230 151 264
rect 185 230 224 264
rect 258 230 297 264
rect 331 230 370 264
rect 404 230 443 264
rect 477 230 516 264
rect 550 230 589 264
rect 623 230 662 264
rect 696 230 735 264
rect 769 230 808 264
rect 842 230 881 264
rect 915 230 954 264
rect 988 230 1027 264
rect 1061 230 1100 264
rect 1134 230 1173 264
rect 1207 230 1246 264
rect 1280 230 1319 264
rect 1353 230 1392 264
rect 1426 230 1465 264
rect 1499 230 1538 264
rect 1572 230 1610 264
rect 1644 230 1682 264
rect 1716 230 1754 264
rect 1788 230 1826 264
rect 1860 230 1898 264
rect 1932 230 1970 264
rect 2004 230 2042 264
rect 2076 230 2114 264
rect 2148 230 2186 264
rect 2220 230 2258 264
rect 2292 230 2330 264
rect 2364 230 2402 264
rect 2436 230 2474 264
rect 2508 230 2546 264
rect 2580 230 2618 264
rect 2652 230 2690 264
rect 2724 230 2762 264
rect 2796 230 2834 264
rect 2868 230 2906 264
rect 2940 230 2952 264
rect 66 224 2952 230
rect 3026 143 3034 195
rect 3086 143 3098 195
rect 3150 143 3156 195
rect 50 108 3060 114
rect 50 74 62 108
rect 96 74 134 108
rect 168 74 206 108
rect 240 74 278 108
rect 312 74 350 108
rect 384 74 422 108
rect 456 74 494 108
rect 528 74 566 108
rect 600 74 638 108
rect 672 74 710 108
rect 744 74 782 108
rect 816 74 854 108
rect 888 74 926 108
rect 960 74 998 108
rect 1032 74 1070 108
rect 1104 74 1142 108
rect 1176 74 1214 108
rect 1248 74 1286 108
rect 1320 74 1358 108
rect 1392 74 1430 108
rect 1464 74 1502 108
rect 1536 74 1574 108
rect 1608 74 1646 108
rect 1680 74 1718 108
rect 1752 74 1790 108
rect 1824 74 1862 108
rect 1896 74 1934 108
rect 1968 74 2006 108
rect 2040 74 2078 108
rect 2112 74 2150 108
rect 2184 74 2222 108
rect 2256 74 2294 108
rect 2328 74 2366 108
rect 2400 74 2438 108
rect 2472 74 2510 108
rect 2544 74 2582 108
rect 2616 74 2654 108
rect 2688 74 2726 108
rect 2760 74 2798 108
rect 2832 74 2870 108
rect 2904 74 2942 108
rect 2976 74 3014 108
rect 3048 74 3060 108
rect 50 68 3060 74
<< via1 >>
rect 3034 335 3086 344
rect 3098 335 3150 344
rect 3034 301 3046 335
rect 3046 301 3084 335
rect 3084 301 3086 335
rect 3098 301 3118 335
rect 3118 301 3150 335
rect 3034 292 3086 301
rect 3098 292 3150 301
rect 3034 186 3086 195
rect 3034 152 3038 186
rect 3038 152 3072 186
rect 3072 152 3086 186
rect 3034 143 3086 152
rect 3098 186 3150 195
rect 3098 152 3110 186
rect 3110 152 3144 186
rect 3144 152 3150 186
rect 3098 143 3150 152
<< metal2 >>
rect 3028 292 3034 344
rect 3086 292 3098 344
rect 3150 292 3156 344
rect 3028 195 3156 292
rect 3028 143 3034 195
rect 3086 143 3098 195
rect 3150 143 3156 195
use sky130_fd_pr__pfet_01v8__example_55959141808177  sky130_fd_pr__pfet_01v8__example_55959141808177_0
timestamp 1707688321
transform 0 1 66 -1 0 375
box -1 0 257 1
<< labels >>
flabel metal1 s 3128 471 3174 500 3 FreeSans 520 0 0 0 PADLO
port 1 nsew
flabel metal1 s 2209 224 2342 270 3 FreeSans 520 0 0 0 TIE_HI
port 2 nsew
flabel metal1 s 2208 69 2338 108 3 FreeSans 520 0 0 0 PUG7_H
port 3 nsew
flabel metal1 s 2209 380 2343 426 3 FreeSans 520 0 0 0 PUG4_H
port 4 nsew
<< properties >>
string GDS_END 69205836
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 69200478
<< end >>
