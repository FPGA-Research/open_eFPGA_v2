magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< pwell >>
rect 8132 936 9681 1121
rect 7115 850 9681 936
rect 7115 380 7201 850
rect 7969 380 9681 850
rect 7115 294 9681 380
rect 8132 67 9681 294
<< mvpsubdiff >>
rect 8158 1087 9655 1095
rect 8158 1053 8182 1087
rect 8216 1053 8253 1087
rect 8287 1053 8324 1087
rect 8358 1053 8395 1087
rect 8429 1053 8466 1087
rect 8500 1053 8537 1087
rect 8571 1053 8608 1087
rect 8642 1053 8679 1087
rect 8713 1053 8750 1087
rect 8784 1053 8821 1087
rect 8855 1053 8892 1087
rect 8926 1053 8963 1087
rect 8997 1053 9034 1087
rect 9068 1053 9105 1087
rect 9139 1053 9176 1087
rect 9210 1053 9247 1087
rect 9281 1053 9317 1087
rect 9351 1053 9387 1087
rect 9421 1053 9457 1087
rect 9491 1053 9527 1087
rect 9561 1053 9597 1087
rect 9631 1053 9655 1087
rect 8158 1019 9655 1053
rect 8158 985 8182 1019
rect 8216 985 8253 1019
rect 8287 985 8324 1019
rect 8358 985 8395 1019
rect 8429 985 8466 1019
rect 8500 985 8537 1019
rect 8571 985 8608 1019
rect 8642 985 8679 1019
rect 8713 985 8750 1019
rect 8784 985 8821 1019
rect 8855 985 8892 1019
rect 8926 985 8963 1019
rect 8997 985 9034 1019
rect 9068 985 9105 1019
rect 9139 985 9176 1019
rect 9210 985 9247 1019
rect 9281 985 9317 1019
rect 9351 985 9387 1019
rect 9421 985 9457 1019
rect 9491 985 9527 1019
rect 9561 985 9597 1019
rect 9631 985 9655 1019
rect 8158 951 9655 985
rect 8158 917 8182 951
rect 8216 917 8253 951
rect 8287 917 8324 951
rect 8358 917 8395 951
rect 8429 917 8466 951
rect 8500 917 8537 951
rect 8571 917 8608 951
rect 8642 917 8679 951
rect 8713 917 8750 951
rect 8784 917 8821 951
rect 8855 917 8892 951
rect 8926 917 8963 951
rect 8997 917 9034 951
rect 9068 917 9105 951
rect 9139 917 9176 951
rect 9210 917 9247 951
rect 9281 917 9317 951
rect 9351 917 9387 951
rect 9421 917 9457 951
rect 9491 917 9527 951
rect 9561 917 9597 951
rect 9631 917 9655 951
rect 7141 876 7209 910
rect 7243 876 7277 910
rect 7311 876 7345 910
rect 7379 876 7413 910
rect 7447 876 7481 910
rect 7515 876 7549 910
rect 7583 876 7617 910
rect 7651 876 7685 910
rect 7719 876 7753 910
rect 7787 876 7821 910
rect 7855 876 7889 910
rect 7923 876 8029 910
rect 7141 830 7175 876
rect 7141 762 7175 796
rect 7995 842 8029 876
rect 7995 774 8029 808
rect 7141 694 7175 728
rect 7141 626 7175 660
rect 7141 558 7175 592
rect 7141 490 7175 524
rect 7995 706 8029 740
rect 7995 638 8029 672
rect 7995 570 8029 604
rect 7995 502 8029 536
rect 7141 422 7175 456
rect 7141 354 7175 388
rect 7995 434 8029 468
rect 7995 354 8029 400
rect 7141 320 7247 354
rect 7281 320 7315 354
rect 7349 320 7383 354
rect 7417 320 7451 354
rect 7485 320 7519 354
rect 7553 320 7587 354
rect 7621 320 7655 354
rect 7689 320 7723 354
rect 7757 320 7791 354
rect 7825 320 7859 354
rect 7893 320 7927 354
rect 7961 320 8029 354
rect 8158 883 9655 917
rect 8158 849 8182 883
rect 8216 849 8253 883
rect 8287 849 8324 883
rect 8358 849 8395 883
rect 8429 849 8466 883
rect 8500 849 8537 883
rect 8571 849 8608 883
rect 8642 849 8679 883
rect 8713 849 8750 883
rect 8784 849 8821 883
rect 8855 849 8892 883
rect 8926 849 8963 883
rect 8997 849 9034 883
rect 9068 849 9105 883
rect 9139 849 9176 883
rect 9210 849 9247 883
rect 9281 849 9317 883
rect 9351 849 9387 883
rect 9421 849 9457 883
rect 9491 849 9527 883
rect 9561 849 9597 883
rect 9631 849 9655 883
rect 8158 815 9655 849
rect 8158 781 8182 815
rect 8216 781 8253 815
rect 8287 781 8324 815
rect 8358 781 8395 815
rect 8429 781 8466 815
rect 8500 781 8537 815
rect 8571 781 8608 815
rect 8642 781 8679 815
rect 8713 781 8750 815
rect 8784 781 8821 815
rect 8855 781 8892 815
rect 8926 781 8963 815
rect 8997 781 9034 815
rect 9068 781 9105 815
rect 9139 781 9176 815
rect 9210 781 9247 815
rect 9281 781 9317 815
rect 9351 781 9387 815
rect 9421 781 9457 815
rect 9491 781 9527 815
rect 9561 781 9597 815
rect 9631 781 9655 815
rect 8158 747 9655 781
rect 8158 713 8182 747
rect 8216 713 8253 747
rect 8287 713 8324 747
rect 8358 713 8395 747
rect 8429 713 8466 747
rect 8500 713 8537 747
rect 8571 713 8608 747
rect 8642 713 8679 747
rect 8713 713 8750 747
rect 8784 713 8821 747
rect 8855 713 8892 747
rect 8926 713 8963 747
rect 8997 713 9034 747
rect 9068 713 9105 747
rect 9139 713 9176 747
rect 9210 713 9247 747
rect 9281 713 9317 747
rect 9351 713 9387 747
rect 9421 713 9457 747
rect 9491 713 9527 747
rect 9561 713 9597 747
rect 9631 713 9655 747
rect 8158 679 9655 713
rect 8158 645 8182 679
rect 8216 645 8253 679
rect 8287 645 8324 679
rect 8358 645 8395 679
rect 8429 645 8466 679
rect 8500 645 8537 679
rect 8571 645 8608 679
rect 8642 645 8679 679
rect 8713 645 8750 679
rect 8784 645 8821 679
rect 8855 645 8892 679
rect 8926 645 8963 679
rect 8997 645 9034 679
rect 9068 645 9105 679
rect 9139 645 9176 679
rect 9210 645 9247 679
rect 9281 645 9317 679
rect 9351 645 9387 679
rect 9421 645 9457 679
rect 9491 645 9527 679
rect 9561 645 9597 679
rect 9631 645 9655 679
rect 8158 611 9655 645
rect 8158 577 8182 611
rect 8216 577 8253 611
rect 8287 577 8324 611
rect 8358 577 8395 611
rect 8429 577 8466 611
rect 8500 577 8537 611
rect 8571 577 8608 611
rect 8642 577 8679 611
rect 8713 577 8750 611
rect 8784 577 8821 611
rect 8855 577 8892 611
rect 8926 577 8963 611
rect 8997 577 9034 611
rect 9068 577 9105 611
rect 9139 577 9176 611
rect 9210 577 9247 611
rect 9281 577 9317 611
rect 9351 577 9387 611
rect 9421 577 9457 611
rect 9491 577 9527 611
rect 9561 577 9597 611
rect 9631 577 9655 611
rect 8158 543 9655 577
rect 8158 509 8182 543
rect 8216 509 8253 543
rect 8287 509 8324 543
rect 8358 509 8395 543
rect 8429 509 8466 543
rect 8500 509 8537 543
rect 8571 509 8608 543
rect 8642 509 8679 543
rect 8713 509 8750 543
rect 8784 509 8821 543
rect 8855 509 8892 543
rect 8926 509 8963 543
rect 8997 509 9034 543
rect 9068 509 9105 543
rect 9139 509 9176 543
rect 9210 509 9247 543
rect 9281 509 9317 543
rect 9351 509 9387 543
rect 9421 509 9457 543
rect 9491 509 9527 543
rect 9561 509 9597 543
rect 9631 509 9655 543
rect 8158 475 9655 509
rect 8158 441 8182 475
rect 8216 441 8253 475
rect 8287 441 8324 475
rect 8358 441 8395 475
rect 8429 441 8466 475
rect 8500 441 8537 475
rect 8571 441 8608 475
rect 8642 441 8679 475
rect 8713 441 8750 475
rect 8784 441 8821 475
rect 8855 441 8892 475
rect 8926 441 8963 475
rect 8997 441 9034 475
rect 9068 441 9105 475
rect 9139 441 9176 475
rect 9210 441 9247 475
rect 9281 441 9317 475
rect 9351 441 9387 475
rect 9421 441 9457 475
rect 9491 441 9527 475
rect 9561 441 9597 475
rect 9631 441 9655 475
rect 8158 407 9655 441
rect 8158 373 8182 407
rect 8216 373 8253 407
rect 8287 373 8324 407
rect 8358 373 8395 407
rect 8429 373 8466 407
rect 8500 373 8537 407
rect 8571 373 8608 407
rect 8642 373 8679 407
rect 8713 373 8750 407
rect 8784 373 8821 407
rect 8855 373 8892 407
rect 8926 373 8963 407
rect 8997 373 9034 407
rect 9068 373 9105 407
rect 9139 373 9176 407
rect 9210 373 9247 407
rect 9281 373 9317 407
rect 9351 373 9387 407
rect 9421 373 9457 407
rect 9491 373 9527 407
rect 9561 373 9597 407
rect 9631 373 9655 407
rect 8158 339 9655 373
rect 8158 305 8182 339
rect 8216 305 8253 339
rect 8287 305 8324 339
rect 8358 305 8395 339
rect 8429 305 8466 339
rect 8500 305 8537 339
rect 8571 305 8608 339
rect 8642 305 8679 339
rect 8713 305 8750 339
rect 8784 305 8821 339
rect 8855 305 8892 339
rect 8926 305 8963 339
rect 8997 305 9034 339
rect 9068 305 9105 339
rect 9139 305 9176 339
rect 9210 305 9247 339
rect 9281 305 9317 339
rect 9351 305 9387 339
rect 9421 305 9457 339
rect 9491 305 9527 339
rect 9561 305 9597 339
rect 9631 305 9655 339
rect 8158 271 9655 305
rect 8158 237 8182 271
rect 8216 237 8253 271
rect 8287 237 8324 271
rect 8358 237 8395 271
rect 8429 237 8466 271
rect 8500 237 8537 271
rect 8571 237 8608 271
rect 8642 237 8679 271
rect 8713 237 8750 271
rect 8784 237 8821 271
rect 8855 237 8892 271
rect 8926 237 8963 271
rect 8997 237 9034 271
rect 9068 237 9105 271
rect 9139 237 9176 271
rect 9210 237 9247 271
rect 9281 237 9317 271
rect 9351 237 9387 271
rect 9421 237 9457 271
rect 9491 237 9527 271
rect 9561 237 9597 271
rect 9631 237 9655 271
rect 8158 203 9655 237
rect 8158 169 8182 203
rect 8216 169 8253 203
rect 8287 169 8324 203
rect 8358 169 8395 203
rect 8429 169 8466 203
rect 8500 169 8537 203
rect 8571 169 8608 203
rect 8642 169 8679 203
rect 8713 169 8750 203
rect 8784 169 8821 203
rect 8855 169 8892 203
rect 8926 169 8963 203
rect 8997 169 9034 203
rect 9068 169 9105 203
rect 9139 169 9176 203
rect 9210 169 9247 203
rect 9281 169 9317 203
rect 9351 169 9387 203
rect 9421 169 9457 203
rect 9491 169 9527 203
rect 9561 169 9597 203
rect 9631 169 9655 203
rect 8158 135 9655 169
rect 8158 101 8182 135
rect 8216 101 8253 135
rect 8287 101 8324 135
rect 8358 101 8395 135
rect 8429 101 8466 135
rect 8500 101 8537 135
rect 8571 101 8608 135
rect 8642 101 8679 135
rect 8713 101 8750 135
rect 8784 101 8821 135
rect 8855 101 8892 135
rect 8926 101 8963 135
rect 8997 101 9034 135
rect 9068 101 9105 135
rect 9139 101 9176 135
rect 9210 101 9247 135
rect 9281 101 9317 135
rect 9351 101 9387 135
rect 9421 101 9457 135
rect 9491 101 9527 135
rect 9561 101 9597 135
rect 9631 101 9655 135
rect 8158 93 9655 101
<< mvpsubdiffcont >>
rect 8182 1053 8216 1087
rect 8253 1053 8287 1087
rect 8324 1053 8358 1087
rect 8395 1053 8429 1087
rect 8466 1053 8500 1087
rect 8537 1053 8571 1087
rect 8608 1053 8642 1087
rect 8679 1053 8713 1087
rect 8750 1053 8784 1087
rect 8821 1053 8855 1087
rect 8892 1053 8926 1087
rect 8963 1053 8997 1087
rect 9034 1053 9068 1087
rect 9105 1053 9139 1087
rect 9176 1053 9210 1087
rect 9247 1053 9281 1087
rect 9317 1053 9351 1087
rect 9387 1053 9421 1087
rect 9457 1053 9491 1087
rect 9527 1053 9561 1087
rect 9597 1053 9631 1087
rect 8182 985 8216 1019
rect 8253 985 8287 1019
rect 8324 985 8358 1019
rect 8395 985 8429 1019
rect 8466 985 8500 1019
rect 8537 985 8571 1019
rect 8608 985 8642 1019
rect 8679 985 8713 1019
rect 8750 985 8784 1019
rect 8821 985 8855 1019
rect 8892 985 8926 1019
rect 8963 985 8997 1019
rect 9034 985 9068 1019
rect 9105 985 9139 1019
rect 9176 985 9210 1019
rect 9247 985 9281 1019
rect 9317 985 9351 1019
rect 9387 985 9421 1019
rect 9457 985 9491 1019
rect 9527 985 9561 1019
rect 9597 985 9631 1019
rect 8182 917 8216 951
rect 8253 917 8287 951
rect 8324 917 8358 951
rect 8395 917 8429 951
rect 8466 917 8500 951
rect 8537 917 8571 951
rect 8608 917 8642 951
rect 8679 917 8713 951
rect 8750 917 8784 951
rect 8821 917 8855 951
rect 8892 917 8926 951
rect 8963 917 8997 951
rect 9034 917 9068 951
rect 9105 917 9139 951
rect 9176 917 9210 951
rect 9247 917 9281 951
rect 9317 917 9351 951
rect 9387 917 9421 951
rect 9457 917 9491 951
rect 9527 917 9561 951
rect 9597 917 9631 951
rect 7209 876 7243 910
rect 7277 876 7311 910
rect 7345 876 7379 910
rect 7413 876 7447 910
rect 7481 876 7515 910
rect 7549 876 7583 910
rect 7617 876 7651 910
rect 7685 876 7719 910
rect 7753 876 7787 910
rect 7821 876 7855 910
rect 7889 876 7923 910
rect 7141 796 7175 830
rect 7141 728 7175 762
rect 7995 808 8029 842
rect 7141 660 7175 694
rect 7141 592 7175 626
rect 7141 524 7175 558
rect 7141 456 7175 490
rect 7995 740 8029 774
rect 7995 672 8029 706
rect 7995 604 8029 638
rect 7995 536 8029 570
rect 7141 388 7175 422
rect 7995 468 8029 502
rect 7995 400 8029 434
rect 7247 320 7281 354
rect 7315 320 7349 354
rect 7383 320 7417 354
rect 7451 320 7485 354
rect 7519 320 7553 354
rect 7587 320 7621 354
rect 7655 320 7689 354
rect 7723 320 7757 354
rect 7791 320 7825 354
rect 7859 320 7893 354
rect 7927 320 7961 354
rect 8182 849 8216 883
rect 8253 849 8287 883
rect 8324 849 8358 883
rect 8395 849 8429 883
rect 8466 849 8500 883
rect 8537 849 8571 883
rect 8608 849 8642 883
rect 8679 849 8713 883
rect 8750 849 8784 883
rect 8821 849 8855 883
rect 8892 849 8926 883
rect 8963 849 8997 883
rect 9034 849 9068 883
rect 9105 849 9139 883
rect 9176 849 9210 883
rect 9247 849 9281 883
rect 9317 849 9351 883
rect 9387 849 9421 883
rect 9457 849 9491 883
rect 9527 849 9561 883
rect 9597 849 9631 883
rect 8182 781 8216 815
rect 8253 781 8287 815
rect 8324 781 8358 815
rect 8395 781 8429 815
rect 8466 781 8500 815
rect 8537 781 8571 815
rect 8608 781 8642 815
rect 8679 781 8713 815
rect 8750 781 8784 815
rect 8821 781 8855 815
rect 8892 781 8926 815
rect 8963 781 8997 815
rect 9034 781 9068 815
rect 9105 781 9139 815
rect 9176 781 9210 815
rect 9247 781 9281 815
rect 9317 781 9351 815
rect 9387 781 9421 815
rect 9457 781 9491 815
rect 9527 781 9561 815
rect 9597 781 9631 815
rect 8182 713 8216 747
rect 8253 713 8287 747
rect 8324 713 8358 747
rect 8395 713 8429 747
rect 8466 713 8500 747
rect 8537 713 8571 747
rect 8608 713 8642 747
rect 8679 713 8713 747
rect 8750 713 8784 747
rect 8821 713 8855 747
rect 8892 713 8926 747
rect 8963 713 8997 747
rect 9034 713 9068 747
rect 9105 713 9139 747
rect 9176 713 9210 747
rect 9247 713 9281 747
rect 9317 713 9351 747
rect 9387 713 9421 747
rect 9457 713 9491 747
rect 9527 713 9561 747
rect 9597 713 9631 747
rect 8182 645 8216 679
rect 8253 645 8287 679
rect 8324 645 8358 679
rect 8395 645 8429 679
rect 8466 645 8500 679
rect 8537 645 8571 679
rect 8608 645 8642 679
rect 8679 645 8713 679
rect 8750 645 8784 679
rect 8821 645 8855 679
rect 8892 645 8926 679
rect 8963 645 8997 679
rect 9034 645 9068 679
rect 9105 645 9139 679
rect 9176 645 9210 679
rect 9247 645 9281 679
rect 9317 645 9351 679
rect 9387 645 9421 679
rect 9457 645 9491 679
rect 9527 645 9561 679
rect 9597 645 9631 679
rect 8182 577 8216 611
rect 8253 577 8287 611
rect 8324 577 8358 611
rect 8395 577 8429 611
rect 8466 577 8500 611
rect 8537 577 8571 611
rect 8608 577 8642 611
rect 8679 577 8713 611
rect 8750 577 8784 611
rect 8821 577 8855 611
rect 8892 577 8926 611
rect 8963 577 8997 611
rect 9034 577 9068 611
rect 9105 577 9139 611
rect 9176 577 9210 611
rect 9247 577 9281 611
rect 9317 577 9351 611
rect 9387 577 9421 611
rect 9457 577 9491 611
rect 9527 577 9561 611
rect 9597 577 9631 611
rect 8182 509 8216 543
rect 8253 509 8287 543
rect 8324 509 8358 543
rect 8395 509 8429 543
rect 8466 509 8500 543
rect 8537 509 8571 543
rect 8608 509 8642 543
rect 8679 509 8713 543
rect 8750 509 8784 543
rect 8821 509 8855 543
rect 8892 509 8926 543
rect 8963 509 8997 543
rect 9034 509 9068 543
rect 9105 509 9139 543
rect 9176 509 9210 543
rect 9247 509 9281 543
rect 9317 509 9351 543
rect 9387 509 9421 543
rect 9457 509 9491 543
rect 9527 509 9561 543
rect 9597 509 9631 543
rect 8182 441 8216 475
rect 8253 441 8287 475
rect 8324 441 8358 475
rect 8395 441 8429 475
rect 8466 441 8500 475
rect 8537 441 8571 475
rect 8608 441 8642 475
rect 8679 441 8713 475
rect 8750 441 8784 475
rect 8821 441 8855 475
rect 8892 441 8926 475
rect 8963 441 8997 475
rect 9034 441 9068 475
rect 9105 441 9139 475
rect 9176 441 9210 475
rect 9247 441 9281 475
rect 9317 441 9351 475
rect 9387 441 9421 475
rect 9457 441 9491 475
rect 9527 441 9561 475
rect 9597 441 9631 475
rect 8182 373 8216 407
rect 8253 373 8287 407
rect 8324 373 8358 407
rect 8395 373 8429 407
rect 8466 373 8500 407
rect 8537 373 8571 407
rect 8608 373 8642 407
rect 8679 373 8713 407
rect 8750 373 8784 407
rect 8821 373 8855 407
rect 8892 373 8926 407
rect 8963 373 8997 407
rect 9034 373 9068 407
rect 9105 373 9139 407
rect 9176 373 9210 407
rect 9247 373 9281 407
rect 9317 373 9351 407
rect 9387 373 9421 407
rect 9457 373 9491 407
rect 9527 373 9561 407
rect 9597 373 9631 407
rect 8182 305 8216 339
rect 8253 305 8287 339
rect 8324 305 8358 339
rect 8395 305 8429 339
rect 8466 305 8500 339
rect 8537 305 8571 339
rect 8608 305 8642 339
rect 8679 305 8713 339
rect 8750 305 8784 339
rect 8821 305 8855 339
rect 8892 305 8926 339
rect 8963 305 8997 339
rect 9034 305 9068 339
rect 9105 305 9139 339
rect 9176 305 9210 339
rect 9247 305 9281 339
rect 9317 305 9351 339
rect 9387 305 9421 339
rect 9457 305 9491 339
rect 9527 305 9561 339
rect 9597 305 9631 339
rect 8182 237 8216 271
rect 8253 237 8287 271
rect 8324 237 8358 271
rect 8395 237 8429 271
rect 8466 237 8500 271
rect 8537 237 8571 271
rect 8608 237 8642 271
rect 8679 237 8713 271
rect 8750 237 8784 271
rect 8821 237 8855 271
rect 8892 237 8926 271
rect 8963 237 8997 271
rect 9034 237 9068 271
rect 9105 237 9139 271
rect 9176 237 9210 271
rect 9247 237 9281 271
rect 9317 237 9351 271
rect 9387 237 9421 271
rect 9457 237 9491 271
rect 9527 237 9561 271
rect 9597 237 9631 271
rect 8182 169 8216 203
rect 8253 169 8287 203
rect 8324 169 8358 203
rect 8395 169 8429 203
rect 8466 169 8500 203
rect 8537 169 8571 203
rect 8608 169 8642 203
rect 8679 169 8713 203
rect 8750 169 8784 203
rect 8821 169 8855 203
rect 8892 169 8926 203
rect 8963 169 8997 203
rect 9034 169 9068 203
rect 9105 169 9139 203
rect 9176 169 9210 203
rect 9247 169 9281 203
rect 9317 169 9351 203
rect 9387 169 9421 203
rect 9457 169 9491 203
rect 9527 169 9561 203
rect 9597 169 9631 203
rect 8182 101 8216 135
rect 8253 101 8287 135
rect 8324 101 8358 135
rect 8395 101 8429 135
rect 8466 101 8500 135
rect 8537 101 8571 135
rect 8608 101 8642 135
rect 8679 101 8713 135
rect 8750 101 8784 135
rect 8821 101 8855 135
rect 8892 101 8926 135
rect 8963 101 8997 135
rect 9034 101 9068 135
rect 9105 101 9139 135
rect 9176 101 9210 135
rect 9247 101 9281 135
rect 9317 101 9351 135
rect 9387 101 9421 135
rect 9457 101 9491 135
rect 9527 101 9561 135
rect 9597 101 9631 135
<< poly >>
rect 7217 727 7283 743
rect 7217 693 7233 727
rect 7267 693 7283 727
rect 7217 632 7283 693
rect 7217 598 7233 632
rect 7267 598 7283 632
rect 7217 537 7283 598
rect 7217 503 7233 537
rect 7267 503 7283 537
rect 7217 487 7283 503
<< polycont >>
rect 7233 693 7267 727
rect 7233 598 7267 632
rect 7233 503 7267 537
<< locali >>
rect 8158 1087 9655 1095
rect 8158 1053 8182 1087
rect 8216 1053 8253 1087
rect 8287 1053 8324 1087
rect 8358 1053 8395 1087
rect 8429 1053 8466 1087
rect 8500 1053 8537 1087
rect 8571 1053 8608 1087
rect 8642 1053 8679 1087
rect 8713 1053 8750 1087
rect 8784 1053 8821 1087
rect 8855 1053 8892 1087
rect 8926 1053 8963 1087
rect 8997 1053 9034 1087
rect 9068 1053 9105 1087
rect 9139 1053 9176 1087
rect 9210 1053 9247 1087
rect 9281 1053 9317 1087
rect 9351 1053 9387 1087
rect 9421 1053 9457 1087
rect 9491 1053 9527 1087
rect 9561 1053 9597 1087
rect 9631 1053 9655 1087
rect 8158 1019 9655 1053
rect 8158 985 8182 1019
rect 8216 985 8253 1019
rect 8287 985 8324 1019
rect 8358 985 8395 1019
rect 8429 985 8466 1019
rect 8500 985 8537 1019
rect 8571 985 8608 1019
rect 8642 985 8679 1019
rect 8713 985 8750 1019
rect 8784 985 8821 1019
rect 8855 985 8892 1019
rect 8926 985 8963 1019
rect 8997 985 9034 1019
rect 9068 985 9105 1019
rect 9139 985 9176 1019
rect 9210 985 9247 1019
rect 9281 985 9317 1019
rect 9351 985 9387 1019
rect 9421 985 9457 1019
rect 9491 985 9527 1019
rect 9561 985 9597 1019
rect 9631 985 9655 1019
rect 8158 951 9655 985
rect 8158 917 8182 951
rect 8216 917 8253 951
rect 8287 917 8324 951
rect 8358 917 8395 951
rect 8429 917 8466 951
rect 8500 917 8537 951
rect 8571 917 8608 951
rect 8642 917 8679 951
rect 8713 917 8750 951
rect 8784 917 8821 951
rect 8855 917 8892 951
rect 8926 917 8963 951
rect 8997 917 9034 951
rect 9068 917 9105 951
rect 9139 917 9176 951
rect 9210 917 9247 951
rect 9281 917 9317 951
rect 9351 917 9387 951
rect 9421 917 9457 951
rect 9491 917 9527 951
rect 9561 917 9597 951
rect 9631 917 9655 951
rect 7135 910 8035 916
rect 7135 876 7209 910
rect 7253 876 7277 910
rect 7331 876 7345 910
rect 7409 876 7413 910
rect 7447 876 7453 910
rect 7515 876 7531 910
rect 7583 876 7609 910
rect 7651 876 7685 910
rect 7721 876 7753 910
rect 7799 876 7821 910
rect 7878 876 7889 910
rect 7957 876 8035 910
rect 7135 870 8035 876
rect 7135 838 7181 870
rect 7135 796 7141 838
rect 7175 796 7181 838
rect 7135 762 7181 796
rect 7989 842 8035 870
rect 7989 798 7995 842
rect 8029 798 8035 842
rect 7135 717 7141 762
rect 7175 717 7181 762
rect 7423 754 7469 788
rect 7503 754 7549 788
rect 7583 754 7629 788
rect 7663 754 7709 788
rect 7743 754 7789 788
rect 7823 754 7869 788
rect 7989 774 8035 798
rect 7135 694 7181 717
rect 7135 630 7141 694
rect 7175 630 7181 694
rect 7135 626 7181 630
rect 7135 592 7141 626
rect 7175 592 7181 626
rect 7135 577 7181 592
rect 7135 524 7141 577
rect 7175 524 7181 577
rect 7135 490 7181 524
rect 7135 456 7141 490
rect 7175 456 7181 490
rect 7233 727 7267 743
rect 7233 632 7267 688
rect 7989 720 7995 774
rect 8029 720 8035 774
rect 7989 706 8035 720
rect 7989 641 7995 706
rect 8029 641 8035 706
rect 7989 638 8035 641
rect 7361 598 7412 632
rect 7446 598 7497 632
rect 7531 598 7581 632
rect 7615 598 7665 632
rect 7699 598 7749 632
rect 7989 604 7995 638
rect 8029 604 8035 638
rect 7233 539 7267 597
rect 7233 487 7267 503
rect 7989 596 8035 604
rect 7989 536 7995 596
rect 8029 536 8035 596
rect 7989 517 8035 536
rect 7135 452 7181 456
rect 7135 388 7141 452
rect 7175 388 7181 452
rect 7423 442 7469 476
rect 7503 442 7549 476
rect 7583 442 7629 476
rect 7663 442 7709 476
rect 7743 442 7789 476
rect 7823 442 7869 476
rect 7989 468 7995 517
rect 8029 468 8035 517
rect 7135 360 7181 388
rect 7989 434 8035 468
rect 7989 400 7995 434
rect 8029 400 8035 434
rect 7989 360 8035 400
rect 7135 354 8035 360
rect 7135 320 7219 354
rect 7281 320 7297 354
rect 7349 320 7375 354
rect 7417 320 7451 354
rect 7487 320 7519 354
rect 7565 320 7587 354
rect 7643 320 7655 354
rect 7721 320 7723 354
rect 7757 320 7765 354
rect 7825 320 7844 354
rect 7893 320 7923 354
rect 7961 320 8035 354
rect 7135 314 8035 320
rect 8158 883 9655 917
rect 8158 849 8182 883
rect 8216 849 8253 883
rect 8287 863 8324 883
rect 8358 863 8395 883
rect 8287 849 8316 863
rect 8358 849 8393 863
rect 8429 849 8466 883
rect 8500 863 8537 883
rect 8571 863 8608 883
rect 8642 863 8679 883
rect 8713 863 8750 883
rect 8784 863 8821 883
rect 8855 863 8892 883
rect 8926 863 8963 883
rect 8503 849 8537 863
rect 8579 849 8608 863
rect 8655 849 8679 863
rect 8731 849 8750 863
rect 8807 849 8821 863
rect 8883 849 8892 863
rect 8959 849 8963 863
rect 8997 863 9034 883
rect 9068 863 9105 883
rect 9139 863 9176 883
rect 9210 863 9247 883
rect 9281 863 9317 883
rect 9351 863 9387 883
rect 8997 849 9001 863
rect 9068 849 9077 863
rect 9139 849 9153 863
rect 9210 849 9229 863
rect 9281 849 9305 863
rect 9351 849 9381 863
rect 9421 849 9457 883
rect 9491 849 9527 883
rect 9561 863 9597 883
rect 9631 863 9655 883
rect 9567 849 9597 863
rect 8158 829 8316 849
rect 8350 829 8393 849
rect 8427 829 8469 849
rect 8503 829 8545 849
rect 8579 829 8621 849
rect 8655 829 8697 849
rect 8731 829 8773 849
rect 8807 829 8849 849
rect 8883 829 8925 849
rect 8959 829 9001 849
rect 9035 829 9077 849
rect 9111 829 9153 849
rect 9187 829 9229 849
rect 9263 829 9305 849
rect 9339 829 9381 849
rect 9415 829 9457 849
rect 9491 829 9533 849
rect 9567 829 9609 849
rect 9643 829 9655 863
rect 8158 815 9655 829
rect 8158 781 8182 815
rect 8216 781 8253 815
rect 8287 785 8324 815
rect 8358 785 8395 815
rect 8287 781 8316 785
rect 8358 781 8393 785
rect 8429 781 8466 815
rect 8500 785 8537 815
rect 8571 785 8608 815
rect 8642 785 8679 815
rect 8713 785 8750 815
rect 8784 785 8821 815
rect 8855 785 8892 815
rect 8926 785 8963 815
rect 8503 781 8537 785
rect 8579 781 8608 785
rect 8655 781 8679 785
rect 8731 781 8750 785
rect 8807 781 8821 785
rect 8883 781 8892 785
rect 8959 781 8963 785
rect 8997 785 9034 815
rect 9068 785 9105 815
rect 9139 785 9176 815
rect 9210 785 9247 815
rect 9281 785 9317 815
rect 9351 785 9387 815
rect 8997 781 9001 785
rect 9068 781 9077 785
rect 9139 781 9153 785
rect 9210 781 9229 785
rect 9281 781 9305 785
rect 9351 781 9381 785
rect 9421 781 9457 815
rect 9491 781 9527 815
rect 9561 785 9597 815
rect 9631 785 9655 815
rect 9567 781 9597 785
rect 8158 751 8316 781
rect 8350 751 8393 781
rect 8427 751 8469 781
rect 8503 751 8545 781
rect 8579 751 8621 781
rect 8655 751 8697 781
rect 8731 751 8773 781
rect 8807 751 8849 781
rect 8883 751 8925 781
rect 8959 751 9001 781
rect 9035 751 9077 781
rect 9111 751 9153 781
rect 9187 751 9229 781
rect 9263 751 9305 781
rect 9339 751 9381 781
rect 9415 751 9457 781
rect 9491 751 9533 781
rect 9567 751 9609 781
rect 9643 751 9655 785
rect 8158 747 9655 751
rect 8158 713 8182 747
rect 8216 713 8253 747
rect 8287 713 8324 747
rect 8358 713 8395 747
rect 8429 713 8466 747
rect 8500 713 8537 747
rect 8571 713 8608 747
rect 8642 713 8679 747
rect 8713 713 8750 747
rect 8784 713 8821 747
rect 8855 713 8892 747
rect 8926 713 8963 747
rect 8997 713 9034 747
rect 9068 713 9105 747
rect 9139 713 9176 747
rect 9210 713 9247 747
rect 9281 713 9317 747
rect 9351 713 9387 747
rect 9421 713 9457 747
rect 9491 713 9527 747
rect 9561 713 9597 747
rect 9631 713 9655 747
rect 8158 707 9655 713
rect 8158 679 8316 707
rect 8350 679 8393 707
rect 8427 679 8469 707
rect 8503 679 8545 707
rect 8579 679 8621 707
rect 8655 679 8697 707
rect 8731 679 8773 707
rect 8807 679 8849 707
rect 8883 679 8925 707
rect 8959 679 9001 707
rect 9035 679 9077 707
rect 9111 679 9153 707
rect 9187 679 9229 707
rect 9263 679 9305 707
rect 9339 679 9381 707
rect 9415 679 9457 707
rect 9491 679 9533 707
rect 9567 679 9609 707
rect 8158 645 8182 679
rect 8216 645 8253 679
rect 8287 673 8316 679
rect 8358 673 8393 679
rect 8287 645 8324 673
rect 8358 645 8395 673
rect 8429 645 8466 679
rect 8503 673 8537 679
rect 8579 673 8608 679
rect 8655 673 8679 679
rect 8731 673 8750 679
rect 8807 673 8821 679
rect 8883 673 8892 679
rect 8959 673 8963 679
rect 8500 645 8537 673
rect 8571 645 8608 673
rect 8642 645 8679 673
rect 8713 645 8750 673
rect 8784 645 8821 673
rect 8855 645 8892 673
rect 8926 645 8963 673
rect 8997 673 9001 679
rect 9068 673 9077 679
rect 9139 673 9153 679
rect 9210 673 9229 679
rect 9281 673 9305 679
rect 9351 673 9381 679
rect 8997 645 9034 673
rect 9068 645 9105 673
rect 9139 645 9176 673
rect 9210 645 9247 673
rect 9281 645 9317 673
rect 9351 645 9387 673
rect 9421 645 9457 679
rect 9491 645 9527 679
rect 9567 673 9597 679
rect 9643 673 9655 707
rect 9561 645 9597 673
rect 9631 645 9655 673
rect 8158 629 9655 645
rect 8158 611 8316 629
rect 8350 611 8393 629
rect 8427 611 8469 629
rect 8503 611 8545 629
rect 8579 611 8621 629
rect 8655 611 8697 629
rect 8731 611 8773 629
rect 8807 611 8849 629
rect 8883 611 8925 629
rect 8959 611 9001 629
rect 9035 611 9077 629
rect 9111 611 9153 629
rect 9187 611 9229 629
rect 9263 611 9305 629
rect 9339 611 9381 629
rect 9415 611 9457 629
rect 9491 611 9533 629
rect 9567 611 9609 629
rect 8158 577 8182 611
rect 8216 577 8253 611
rect 8287 595 8316 611
rect 8358 595 8393 611
rect 8287 577 8324 595
rect 8358 577 8395 595
rect 8429 577 8466 611
rect 8503 595 8537 611
rect 8579 595 8608 611
rect 8655 595 8679 611
rect 8731 595 8750 611
rect 8807 595 8821 611
rect 8883 595 8892 611
rect 8959 595 8963 611
rect 8500 577 8537 595
rect 8571 577 8608 595
rect 8642 577 8679 595
rect 8713 577 8750 595
rect 8784 577 8821 595
rect 8855 577 8892 595
rect 8926 577 8963 595
rect 8997 595 9001 611
rect 9068 595 9077 611
rect 9139 595 9153 611
rect 9210 595 9229 611
rect 9281 595 9305 611
rect 9351 595 9381 611
rect 8997 577 9034 595
rect 9068 577 9105 595
rect 9139 577 9176 595
rect 9210 577 9247 595
rect 9281 577 9317 595
rect 9351 577 9387 595
rect 9421 577 9457 611
rect 9491 577 9527 611
rect 9567 595 9597 611
rect 9643 595 9655 629
rect 9561 577 9597 595
rect 9631 577 9655 595
rect 8158 551 9655 577
rect 8158 543 8316 551
rect 8350 543 8393 551
rect 8427 543 8469 551
rect 8503 543 8545 551
rect 8579 543 8621 551
rect 8655 543 8697 551
rect 8731 543 8773 551
rect 8807 543 8849 551
rect 8883 543 8925 551
rect 8959 543 9001 551
rect 9035 543 9077 551
rect 9111 543 9153 551
rect 9187 543 9229 551
rect 9263 543 9305 551
rect 9339 543 9381 551
rect 9415 543 9457 551
rect 9491 543 9533 551
rect 9567 543 9609 551
rect 8158 509 8182 543
rect 8216 509 8253 543
rect 8287 517 8316 543
rect 8358 517 8393 543
rect 8287 509 8324 517
rect 8358 509 8395 517
rect 8429 509 8466 543
rect 8503 517 8537 543
rect 8579 517 8608 543
rect 8655 517 8679 543
rect 8731 517 8750 543
rect 8807 517 8821 543
rect 8883 517 8892 543
rect 8959 517 8963 543
rect 8500 509 8537 517
rect 8571 509 8608 517
rect 8642 509 8679 517
rect 8713 509 8750 517
rect 8784 509 8821 517
rect 8855 509 8892 517
rect 8926 509 8963 517
rect 8997 517 9001 543
rect 9068 517 9077 543
rect 9139 517 9153 543
rect 9210 517 9229 543
rect 9281 517 9305 543
rect 9351 517 9381 543
rect 8997 509 9034 517
rect 9068 509 9105 517
rect 9139 509 9176 517
rect 9210 509 9247 517
rect 9281 509 9317 517
rect 9351 509 9387 517
rect 9421 509 9457 543
rect 9491 509 9527 543
rect 9567 517 9597 543
rect 9643 517 9655 551
rect 9561 509 9597 517
rect 9631 509 9655 517
rect 8158 475 9655 509
rect 8158 441 8182 475
rect 8216 441 8253 475
rect 8287 473 8324 475
rect 8358 473 8395 475
rect 8287 441 8316 473
rect 8358 441 8393 473
rect 8429 441 8466 475
rect 8500 473 8537 475
rect 8571 473 8608 475
rect 8642 473 8679 475
rect 8713 473 8750 475
rect 8784 473 8821 475
rect 8855 473 8892 475
rect 8926 473 8963 475
rect 8503 441 8537 473
rect 8579 441 8608 473
rect 8655 441 8679 473
rect 8731 441 8750 473
rect 8807 441 8821 473
rect 8883 441 8892 473
rect 8959 441 8963 473
rect 8997 473 9034 475
rect 9068 473 9105 475
rect 9139 473 9176 475
rect 9210 473 9247 475
rect 9281 473 9317 475
rect 9351 473 9387 475
rect 8997 441 9001 473
rect 9068 441 9077 473
rect 9139 441 9153 473
rect 9210 441 9229 473
rect 9281 441 9305 473
rect 9351 441 9381 473
rect 9421 441 9457 475
rect 9491 441 9527 475
rect 9561 473 9597 475
rect 9631 473 9655 475
rect 9567 441 9597 473
rect 8158 439 8316 441
rect 8350 439 8393 441
rect 8427 439 8469 441
rect 8503 439 8545 441
rect 8579 439 8621 441
rect 8655 439 8697 441
rect 8731 439 8773 441
rect 8807 439 8849 441
rect 8883 439 8925 441
rect 8959 439 9001 441
rect 9035 439 9077 441
rect 9111 439 9153 441
rect 9187 439 9229 441
rect 9263 439 9305 441
rect 9339 439 9381 441
rect 9415 439 9457 441
rect 9491 439 9533 441
rect 9567 439 9609 441
rect 9643 439 9655 473
rect 8158 407 9655 439
rect 8158 373 8182 407
rect 8216 373 8253 407
rect 8287 395 8324 407
rect 8358 395 8395 407
rect 8287 373 8316 395
rect 8358 373 8393 395
rect 8429 373 8466 407
rect 8500 395 8537 407
rect 8571 395 8608 407
rect 8642 395 8679 407
rect 8713 395 8750 407
rect 8784 395 8821 407
rect 8855 395 8892 407
rect 8926 395 8963 407
rect 8503 373 8537 395
rect 8579 373 8608 395
rect 8655 373 8679 395
rect 8731 373 8750 395
rect 8807 373 8821 395
rect 8883 373 8892 395
rect 8959 373 8963 395
rect 8997 395 9034 407
rect 9068 395 9105 407
rect 9139 395 9176 407
rect 9210 395 9247 407
rect 9281 395 9317 407
rect 9351 395 9387 407
rect 8997 373 9001 395
rect 9068 373 9077 395
rect 9139 373 9153 395
rect 9210 373 9229 395
rect 9281 373 9305 395
rect 9351 373 9381 395
rect 9421 373 9457 407
rect 9491 373 9527 407
rect 9561 395 9597 407
rect 9631 395 9655 407
rect 9567 373 9597 395
rect 8158 361 8316 373
rect 8350 361 8393 373
rect 8427 361 8469 373
rect 8503 361 8545 373
rect 8579 361 8621 373
rect 8655 361 8697 373
rect 8731 361 8773 373
rect 8807 361 8849 373
rect 8883 361 8925 373
rect 8959 361 9001 373
rect 9035 361 9077 373
rect 9111 361 9153 373
rect 9187 361 9229 373
rect 9263 361 9305 373
rect 9339 361 9381 373
rect 9415 361 9457 373
rect 9491 361 9533 373
rect 9567 361 9609 373
rect 9643 361 9655 395
rect 8158 339 9655 361
rect 8158 305 8182 339
rect 8216 305 8253 339
rect 8287 305 8324 339
rect 8358 305 8395 339
rect 8429 305 8466 339
rect 8500 305 8537 339
rect 8571 305 8608 339
rect 8642 305 8679 339
rect 8713 305 8750 339
rect 8784 305 8821 339
rect 8855 305 8892 339
rect 8926 305 8963 339
rect 8997 305 9034 339
rect 9068 305 9105 339
rect 9139 305 9176 339
rect 9210 305 9247 339
rect 9281 305 9317 339
rect 9351 305 9387 339
rect 9421 305 9457 339
rect 9491 305 9527 339
rect 9561 305 9597 339
rect 9631 305 9655 339
rect 8158 271 9655 305
rect 8158 237 8182 271
rect 8216 237 8253 271
rect 8287 237 8324 271
rect 8358 237 8395 271
rect 8429 237 8466 271
rect 8500 237 8537 271
rect 8571 237 8608 271
rect 8642 237 8679 271
rect 8713 237 8750 271
rect 8784 237 8821 271
rect 8855 237 8892 271
rect 8926 237 8963 271
rect 8997 237 9034 271
rect 9068 237 9105 271
rect 9139 237 9176 271
rect 9210 237 9247 271
rect 9281 237 9317 271
rect 9351 237 9387 271
rect 9421 237 9457 271
rect 9491 237 9527 271
rect 9561 237 9597 271
rect 9631 237 9655 271
rect 8158 203 9655 237
rect 8158 169 8182 203
rect 8216 169 8253 203
rect 8287 169 8324 203
rect 8358 169 8395 203
rect 8429 169 8466 203
rect 8500 169 8537 203
rect 8571 169 8608 203
rect 8642 169 8679 203
rect 8713 169 8750 203
rect 8784 169 8821 203
rect 8855 169 8892 203
rect 8926 169 8963 203
rect 8997 169 9034 203
rect 9068 169 9105 203
rect 9139 169 9176 203
rect 9210 169 9247 203
rect 9281 169 9317 203
rect 9351 169 9387 203
rect 9421 169 9457 203
rect 9491 169 9527 203
rect 9561 169 9597 203
rect 9631 169 9655 203
rect 8158 135 9655 169
rect 8158 101 8182 135
rect 8216 101 8253 135
rect 8287 101 8324 135
rect 8358 101 8395 135
rect 8429 101 8466 135
rect 8500 101 8537 135
rect 8571 101 8608 135
rect 8642 101 8679 135
rect 8713 101 8750 135
rect 8784 101 8821 135
rect 8855 101 8892 135
rect 8926 101 8963 135
rect 8997 101 9034 135
rect 9068 101 9105 135
rect 9139 101 9176 135
rect 9210 101 9247 135
rect 9281 101 9317 135
rect 9351 101 9387 135
rect 9421 101 9457 135
rect 9491 101 9527 135
rect 9561 101 9597 135
rect 9631 101 9655 135
rect 8158 93 9655 101
<< viali >>
rect 7219 876 7243 910
rect 7243 876 7253 910
rect 7297 876 7311 910
rect 7311 876 7331 910
rect 7375 876 7379 910
rect 7379 876 7409 910
rect 7453 876 7481 910
rect 7481 876 7487 910
rect 7531 876 7549 910
rect 7549 876 7565 910
rect 7609 876 7617 910
rect 7617 876 7643 910
rect 7687 876 7719 910
rect 7719 876 7721 910
rect 7765 876 7787 910
rect 7787 876 7799 910
rect 7844 876 7855 910
rect 7855 876 7878 910
rect 7923 876 7957 910
rect 7141 830 7175 838
rect 7141 804 7175 830
rect 7995 808 8029 832
rect 7995 798 8029 808
rect 7141 728 7175 751
rect 7141 717 7175 728
rect 7389 754 7423 788
rect 7469 754 7503 788
rect 7549 754 7583 788
rect 7629 754 7663 788
rect 7709 754 7743 788
rect 7789 754 7823 788
rect 7869 754 7903 788
rect 7141 660 7175 664
rect 7141 630 7175 660
rect 7141 558 7175 577
rect 7141 543 7175 558
rect 7233 693 7267 722
rect 7233 688 7267 693
rect 7995 740 8029 754
rect 7995 720 8029 740
rect 7995 672 8029 675
rect 7995 641 8029 672
rect 7233 598 7267 631
rect 7327 598 7361 632
rect 7412 598 7446 632
rect 7497 598 7531 632
rect 7581 598 7615 632
rect 7665 598 7699 632
rect 7749 598 7783 632
rect 7233 597 7267 598
rect 7233 537 7267 539
rect 7233 505 7267 537
rect 7995 570 8029 596
rect 7995 562 8029 570
rect 7141 422 7175 452
rect 7141 418 7175 422
rect 7389 442 7423 476
rect 7469 442 7503 476
rect 7549 442 7583 476
rect 7629 442 7663 476
rect 7709 442 7743 476
rect 7789 442 7823 476
rect 7869 442 7903 476
rect 7995 502 8029 517
rect 7995 483 8029 502
rect 7219 320 7247 354
rect 7247 320 7253 354
rect 7297 320 7315 354
rect 7315 320 7331 354
rect 7375 320 7383 354
rect 7383 320 7409 354
rect 7453 320 7485 354
rect 7485 320 7487 354
rect 7531 320 7553 354
rect 7553 320 7565 354
rect 7609 320 7621 354
rect 7621 320 7643 354
rect 7687 320 7689 354
rect 7689 320 7721 354
rect 7765 320 7791 354
rect 7791 320 7799 354
rect 7844 320 7859 354
rect 7859 320 7878 354
rect 7923 320 7927 354
rect 7927 320 7957 354
rect 8316 849 8324 863
rect 8324 849 8350 863
rect 8393 849 8395 863
rect 8395 849 8427 863
rect 8469 849 8500 863
rect 8500 849 8503 863
rect 8545 849 8571 863
rect 8571 849 8579 863
rect 8621 849 8642 863
rect 8642 849 8655 863
rect 8697 849 8713 863
rect 8713 849 8731 863
rect 8773 849 8784 863
rect 8784 849 8807 863
rect 8849 849 8855 863
rect 8855 849 8883 863
rect 8925 849 8926 863
rect 8926 849 8959 863
rect 9001 849 9034 863
rect 9034 849 9035 863
rect 9077 849 9105 863
rect 9105 849 9111 863
rect 9153 849 9176 863
rect 9176 849 9187 863
rect 9229 849 9247 863
rect 9247 849 9263 863
rect 9305 849 9317 863
rect 9317 849 9339 863
rect 9381 849 9387 863
rect 9387 849 9415 863
rect 9457 849 9491 863
rect 9533 849 9561 863
rect 9561 849 9567 863
rect 9609 849 9631 863
rect 9631 849 9643 863
rect 8316 829 8350 849
rect 8393 829 8427 849
rect 8469 829 8503 849
rect 8545 829 8579 849
rect 8621 829 8655 849
rect 8697 829 8731 849
rect 8773 829 8807 849
rect 8849 829 8883 849
rect 8925 829 8959 849
rect 9001 829 9035 849
rect 9077 829 9111 849
rect 9153 829 9187 849
rect 9229 829 9263 849
rect 9305 829 9339 849
rect 9381 829 9415 849
rect 9457 829 9491 849
rect 9533 829 9567 849
rect 9609 829 9643 849
rect 8316 781 8324 785
rect 8324 781 8350 785
rect 8393 781 8395 785
rect 8395 781 8427 785
rect 8469 781 8500 785
rect 8500 781 8503 785
rect 8545 781 8571 785
rect 8571 781 8579 785
rect 8621 781 8642 785
rect 8642 781 8655 785
rect 8697 781 8713 785
rect 8713 781 8731 785
rect 8773 781 8784 785
rect 8784 781 8807 785
rect 8849 781 8855 785
rect 8855 781 8883 785
rect 8925 781 8926 785
rect 8926 781 8959 785
rect 9001 781 9034 785
rect 9034 781 9035 785
rect 9077 781 9105 785
rect 9105 781 9111 785
rect 9153 781 9176 785
rect 9176 781 9187 785
rect 9229 781 9247 785
rect 9247 781 9263 785
rect 9305 781 9317 785
rect 9317 781 9339 785
rect 9381 781 9387 785
rect 9387 781 9415 785
rect 9457 781 9491 785
rect 9533 781 9561 785
rect 9561 781 9567 785
rect 9609 781 9631 785
rect 9631 781 9643 785
rect 8316 751 8350 781
rect 8393 751 8427 781
rect 8469 751 8503 781
rect 8545 751 8579 781
rect 8621 751 8655 781
rect 8697 751 8731 781
rect 8773 751 8807 781
rect 8849 751 8883 781
rect 8925 751 8959 781
rect 9001 751 9035 781
rect 9077 751 9111 781
rect 9153 751 9187 781
rect 9229 751 9263 781
rect 9305 751 9339 781
rect 9381 751 9415 781
rect 9457 751 9491 781
rect 9533 751 9567 781
rect 9609 751 9643 781
rect 8316 679 8350 707
rect 8393 679 8427 707
rect 8469 679 8503 707
rect 8545 679 8579 707
rect 8621 679 8655 707
rect 8697 679 8731 707
rect 8773 679 8807 707
rect 8849 679 8883 707
rect 8925 679 8959 707
rect 9001 679 9035 707
rect 9077 679 9111 707
rect 9153 679 9187 707
rect 9229 679 9263 707
rect 9305 679 9339 707
rect 9381 679 9415 707
rect 9457 679 9491 707
rect 9533 679 9567 707
rect 9609 679 9643 707
rect 8316 673 8324 679
rect 8324 673 8350 679
rect 8393 673 8395 679
rect 8395 673 8427 679
rect 8469 673 8500 679
rect 8500 673 8503 679
rect 8545 673 8571 679
rect 8571 673 8579 679
rect 8621 673 8642 679
rect 8642 673 8655 679
rect 8697 673 8713 679
rect 8713 673 8731 679
rect 8773 673 8784 679
rect 8784 673 8807 679
rect 8849 673 8855 679
rect 8855 673 8883 679
rect 8925 673 8926 679
rect 8926 673 8959 679
rect 9001 673 9034 679
rect 9034 673 9035 679
rect 9077 673 9105 679
rect 9105 673 9111 679
rect 9153 673 9176 679
rect 9176 673 9187 679
rect 9229 673 9247 679
rect 9247 673 9263 679
rect 9305 673 9317 679
rect 9317 673 9339 679
rect 9381 673 9387 679
rect 9387 673 9415 679
rect 9457 673 9491 679
rect 9533 673 9561 679
rect 9561 673 9567 679
rect 9609 673 9631 679
rect 9631 673 9643 679
rect 8316 611 8350 629
rect 8393 611 8427 629
rect 8469 611 8503 629
rect 8545 611 8579 629
rect 8621 611 8655 629
rect 8697 611 8731 629
rect 8773 611 8807 629
rect 8849 611 8883 629
rect 8925 611 8959 629
rect 9001 611 9035 629
rect 9077 611 9111 629
rect 9153 611 9187 629
rect 9229 611 9263 629
rect 9305 611 9339 629
rect 9381 611 9415 629
rect 9457 611 9491 629
rect 9533 611 9567 629
rect 9609 611 9643 629
rect 8316 595 8324 611
rect 8324 595 8350 611
rect 8393 595 8395 611
rect 8395 595 8427 611
rect 8469 595 8500 611
rect 8500 595 8503 611
rect 8545 595 8571 611
rect 8571 595 8579 611
rect 8621 595 8642 611
rect 8642 595 8655 611
rect 8697 595 8713 611
rect 8713 595 8731 611
rect 8773 595 8784 611
rect 8784 595 8807 611
rect 8849 595 8855 611
rect 8855 595 8883 611
rect 8925 595 8926 611
rect 8926 595 8959 611
rect 9001 595 9034 611
rect 9034 595 9035 611
rect 9077 595 9105 611
rect 9105 595 9111 611
rect 9153 595 9176 611
rect 9176 595 9187 611
rect 9229 595 9247 611
rect 9247 595 9263 611
rect 9305 595 9317 611
rect 9317 595 9339 611
rect 9381 595 9387 611
rect 9387 595 9415 611
rect 9457 595 9491 611
rect 9533 595 9561 611
rect 9561 595 9567 611
rect 9609 595 9631 611
rect 9631 595 9643 611
rect 8316 543 8350 551
rect 8393 543 8427 551
rect 8469 543 8503 551
rect 8545 543 8579 551
rect 8621 543 8655 551
rect 8697 543 8731 551
rect 8773 543 8807 551
rect 8849 543 8883 551
rect 8925 543 8959 551
rect 9001 543 9035 551
rect 9077 543 9111 551
rect 9153 543 9187 551
rect 9229 543 9263 551
rect 9305 543 9339 551
rect 9381 543 9415 551
rect 9457 543 9491 551
rect 9533 543 9567 551
rect 9609 543 9643 551
rect 8316 517 8324 543
rect 8324 517 8350 543
rect 8393 517 8395 543
rect 8395 517 8427 543
rect 8469 517 8500 543
rect 8500 517 8503 543
rect 8545 517 8571 543
rect 8571 517 8579 543
rect 8621 517 8642 543
rect 8642 517 8655 543
rect 8697 517 8713 543
rect 8713 517 8731 543
rect 8773 517 8784 543
rect 8784 517 8807 543
rect 8849 517 8855 543
rect 8855 517 8883 543
rect 8925 517 8926 543
rect 8926 517 8959 543
rect 9001 517 9034 543
rect 9034 517 9035 543
rect 9077 517 9105 543
rect 9105 517 9111 543
rect 9153 517 9176 543
rect 9176 517 9187 543
rect 9229 517 9247 543
rect 9247 517 9263 543
rect 9305 517 9317 543
rect 9317 517 9339 543
rect 9381 517 9387 543
rect 9387 517 9415 543
rect 9457 517 9491 543
rect 9533 517 9561 543
rect 9561 517 9567 543
rect 9609 517 9631 543
rect 9631 517 9643 543
rect 8316 441 8324 473
rect 8324 441 8350 473
rect 8393 441 8395 473
rect 8395 441 8427 473
rect 8469 441 8500 473
rect 8500 441 8503 473
rect 8545 441 8571 473
rect 8571 441 8579 473
rect 8621 441 8642 473
rect 8642 441 8655 473
rect 8697 441 8713 473
rect 8713 441 8731 473
rect 8773 441 8784 473
rect 8784 441 8807 473
rect 8849 441 8855 473
rect 8855 441 8883 473
rect 8925 441 8926 473
rect 8926 441 8959 473
rect 9001 441 9034 473
rect 9034 441 9035 473
rect 9077 441 9105 473
rect 9105 441 9111 473
rect 9153 441 9176 473
rect 9176 441 9187 473
rect 9229 441 9247 473
rect 9247 441 9263 473
rect 9305 441 9317 473
rect 9317 441 9339 473
rect 9381 441 9387 473
rect 9387 441 9415 473
rect 9457 441 9491 473
rect 9533 441 9561 473
rect 9561 441 9567 473
rect 9609 441 9631 473
rect 9631 441 9643 473
rect 8316 439 8350 441
rect 8393 439 8427 441
rect 8469 439 8503 441
rect 8545 439 8579 441
rect 8621 439 8655 441
rect 8697 439 8731 441
rect 8773 439 8807 441
rect 8849 439 8883 441
rect 8925 439 8959 441
rect 9001 439 9035 441
rect 9077 439 9111 441
rect 9153 439 9187 441
rect 9229 439 9263 441
rect 9305 439 9339 441
rect 9381 439 9415 441
rect 9457 439 9491 441
rect 9533 439 9567 441
rect 9609 439 9643 441
rect 8316 373 8324 395
rect 8324 373 8350 395
rect 8393 373 8395 395
rect 8395 373 8427 395
rect 8469 373 8500 395
rect 8500 373 8503 395
rect 8545 373 8571 395
rect 8571 373 8579 395
rect 8621 373 8642 395
rect 8642 373 8655 395
rect 8697 373 8713 395
rect 8713 373 8731 395
rect 8773 373 8784 395
rect 8784 373 8807 395
rect 8849 373 8855 395
rect 8855 373 8883 395
rect 8925 373 8926 395
rect 8926 373 8959 395
rect 9001 373 9034 395
rect 9034 373 9035 395
rect 9077 373 9105 395
rect 9105 373 9111 395
rect 9153 373 9176 395
rect 9176 373 9187 395
rect 9229 373 9247 395
rect 9247 373 9263 395
rect 9305 373 9317 395
rect 9317 373 9339 395
rect 9381 373 9387 395
rect 9387 373 9415 395
rect 9457 373 9491 395
rect 9533 373 9561 395
rect 9561 373 9567 395
rect 9609 373 9631 395
rect 9631 373 9643 395
rect 8316 361 8350 373
rect 8393 361 8427 373
rect 8469 361 8503 373
rect 8545 361 8579 373
rect 8621 361 8655 373
rect 8697 361 8731 373
rect 8773 361 8807 373
rect 8849 361 8883 373
rect 8925 361 8959 373
rect 9001 361 9035 373
rect 9077 361 9111 373
rect 9153 361 9187 373
rect 9229 361 9263 373
rect 9305 361 9339 373
rect 9381 361 9415 373
rect 9457 361 9491 373
rect 9533 361 9567 373
rect 9609 361 9643 373
<< metal1 >>
tri 6795 39966 6829 40000 se
rect 385 38879 437 39966
tri 437 39886 471 39920 nw
tri 2430 39886 2464 39920 ne
rect 385 38811 437 38827
rect 385 38743 437 38759
rect 385 36155 437 38691
rect 2464 38879 2516 39966
tri 2516 39886 2550 39920 nw
tri 4572 39886 4606 39920 ne
rect 2464 38811 2516 38827
rect 2464 38743 2516 38759
rect 385 36087 437 36103
rect 385 36019 437 36035
rect 385 34047 437 35967
rect 385 33979 437 33995
rect 385 33911 437 33927
rect 385 31323 437 33859
rect 385 31255 437 31271
rect 385 31187 437 31203
rect 385 29215 437 31135
rect 385 29147 437 29163
rect 385 29079 437 29095
rect 385 26491 437 29027
rect 385 26423 437 26439
rect 385 26355 437 26371
rect 385 24383 437 26303
rect 385 24315 437 24331
rect 385 24247 437 24263
rect 385 21659 437 24195
rect 385 21591 437 21607
rect 385 21523 437 21539
rect 385 19551 437 21471
rect 385 19483 437 19499
rect 385 19415 437 19431
rect 385 16827 437 19363
rect 385 16759 437 16775
rect 385 16691 437 16707
rect 385 14719 437 16639
rect 385 14651 437 14667
rect 385 14583 437 14599
rect 385 11995 437 14531
rect 385 11927 437 11943
rect 385 11859 437 11875
rect 385 9887 437 11807
rect 385 9819 437 9835
rect 385 9751 437 9767
rect 385 4376 437 9699
rect 626 38055 678 38061
rect 626 37991 678 38003
rect 626 4684 678 37939
rect 862 37087 914 37093
rect 862 37023 914 37035
tri 678 4701 712 4735 sw
rect 862 4684 914 36971
rect 2464 36155 2516 38691
rect 2464 36087 2516 36103
rect 2464 36019 2516 36035
rect 2464 34047 2516 35967
rect 2464 33979 2516 33995
rect 2464 33911 2516 33927
rect 1098 33223 1150 33229
rect 1098 33159 1150 33171
tri 914 4701 948 4735 sw
rect 1098 4684 1150 33107
rect 1337 32255 1389 32261
rect 1337 32191 1389 32203
tri 1150 4701 1184 4735 sw
rect 1337 4684 1389 32139
rect 2464 31323 2516 33859
rect 2464 31255 2516 31271
rect 2464 31187 2516 31203
rect 2464 29215 2516 31135
rect 2464 29147 2516 29163
rect 2464 29079 2516 29095
rect 1573 28391 1625 28397
rect 1573 28327 1625 28339
tri 1389 4701 1423 4735 sw
rect 1573 4684 1625 28275
rect 1809 27423 1861 27429
rect 1809 27359 1861 27371
tri 1625 4701 1659 4735 sw
rect 1809 4684 1861 27307
rect 2464 26491 2516 29027
rect 2464 26423 2516 26439
rect 2464 26355 2516 26371
rect 2464 24383 2516 26303
rect 2464 24315 2516 24331
rect 2464 24247 2516 24263
rect 2045 23559 2097 23565
rect 2045 23495 2097 23507
tri 1861 4701 1895 4735 sw
rect 2045 4684 2097 23443
rect 2278 22591 2330 22597
rect 2278 22527 2330 22539
tri 2097 4701 2131 4735 sw
rect 2278 4684 2330 22475
rect 2464 21659 2516 24195
rect 2464 21591 2516 21607
rect 2464 21523 2516 21539
rect 2464 19551 2516 21471
rect 2464 19483 2516 19499
rect 2464 19415 2516 19431
rect 2464 16827 2516 19363
rect 4606 38879 4658 39966
tri 4658 39886 4692 39920 nw
tri 6711 39886 6745 39920 ne
rect 4606 38811 4658 38827
rect 4606 38743 4658 38759
rect 4606 36155 4658 38691
rect 6745 38879 6829 39966
rect 9725 39919 9777 39965
rect 10860 39920 10912 39965
tri 10826 39919 10827 39920 ne
rect 10827 39919 10912 39920
rect 9725 39886 9778 39919
tri 9778 39886 9811 39919 nw
tri 10827 39886 10860 39919 ne
rect 6797 38827 6829 38879
rect 6745 38811 6829 38827
rect 6797 38759 6829 38811
rect 6745 38743 6829 38759
rect 6797 38691 6829 38743
rect 4606 36087 4658 36103
rect 4606 36019 4658 36035
rect 4606 34047 4658 35967
rect 4606 33979 4658 33995
rect 4606 33911 4658 33927
rect 4606 31323 4658 33859
rect 4606 31255 4658 31271
rect 4606 31187 4658 31203
rect 4606 29215 4658 31135
rect 4606 29147 4658 29163
rect 4606 29079 4658 29095
rect 4606 26491 4658 29027
rect 4606 26423 4658 26439
rect 4606 26355 4658 26371
rect 4606 24383 4658 26303
rect 4606 24315 4658 24331
rect 4606 24247 4658 24263
rect 4606 21659 4658 24195
rect 4606 21591 4658 21607
rect 4606 21523 4658 21539
rect 4606 19551 4658 21471
rect 4606 19483 4658 19499
rect 4606 19415 4658 19431
rect 2464 16759 2516 16775
rect 2464 16691 2516 16707
rect 2464 14719 2516 16639
rect 2464 14651 2516 14667
rect 2464 14583 2516 14599
rect 2464 11995 2516 14531
rect 2464 11927 2516 11943
rect 2464 11859 2516 11875
rect 2464 9887 2516 11807
rect 2464 9819 2516 9835
rect 2464 9751 2516 9767
tri 437 4422 471 4456 sw
tri 2430 4422 2464 4456 se
rect 2464 4376 2516 9699
rect 2771 18727 2823 18733
rect 2771 18663 2823 18675
rect 2771 4684 2823 18611
rect 3007 17759 3059 17765
rect 3007 17695 3059 17707
tri 2823 4701 2857 4735 sw
rect 3007 4684 3059 17643
rect 4606 16827 4658 19363
rect 4606 16759 4658 16775
rect 4606 16691 4658 16707
rect 4606 14719 4658 16639
rect 4606 14651 4658 14667
rect 4606 14583 4658 14599
rect 3243 13895 3295 13901
rect 3243 13831 3295 13843
tri 3059 4701 3093 4735 sw
rect 3243 4684 3295 13779
rect 3479 12927 3531 12933
rect 3479 12863 3531 12875
tri 3295 4701 3329 4735 sw
rect 3479 4684 3531 12811
rect 4606 11995 4658 14531
rect 4606 11927 4658 11943
rect 4606 11859 4658 11875
rect 4606 9887 4658 11807
rect 4606 9819 4658 9835
rect 4606 9751 4658 9767
rect 3715 9063 3767 9069
rect 3715 8999 3767 9011
tri 3531 4701 3565 4735 sw
rect 3715 4684 3767 8947
rect 3951 8095 4003 8101
rect 3951 8031 4003 8043
tri 3767 4701 3801 4735 sw
rect 3951 4684 4003 7979
tri 4003 4701 4037 4735 sw
rect 4299 4695 4351 4701
rect 4299 4631 4351 4643
rect 4299 4573 4351 4579
tri 2516 4422 2550 4456 sw
tri 4572 4422 4606 4456 se
rect 4606 4376 4658 9699
rect 4910 38432 4962 38438
rect 4910 38368 4962 38380
rect 4910 4684 4962 38316
rect 5146 36710 5198 36716
rect 5146 36646 5198 36658
tri 4962 4702 4996 4736 sw
rect 5146 4684 5198 36594
rect 6745 36155 6829 38691
rect 9633 38879 9685 38885
rect 9633 38811 9685 38827
rect 9633 38743 9685 38759
rect 9633 38685 9685 38691
rect 9725 38879 9777 39886
tri 9777 39885 9778 39886 nw
rect 9725 38811 9777 38827
rect 9725 38743 9777 38759
rect 6797 36103 6829 36155
rect 6745 36087 6829 36103
rect 6797 36035 6829 36087
rect 6745 36019 6829 36035
rect 6797 35967 6829 36019
rect 6745 34047 6829 35967
rect 9633 36155 9685 36161
rect 9633 36087 9685 36103
rect 9633 36019 9685 36035
rect 9633 35961 9685 35967
rect 9725 36155 9777 38691
rect 9725 36087 9777 36103
rect 9725 36019 9777 36035
rect 6797 33995 6829 34047
rect 6745 33979 6829 33995
rect 6797 33927 6829 33979
rect 6745 33911 6829 33927
rect 6797 33859 6829 33911
rect 5382 33600 5434 33606
rect 5382 33536 5434 33548
tri 5198 4702 5232 4736 sw
rect 5382 4684 5434 33484
rect 5618 31878 5670 31884
rect 5618 31814 5670 31826
tri 5434 4702 5468 4736 sw
rect 5618 4684 5670 31762
rect 6745 31323 6829 33859
rect 9633 34047 9685 34053
rect 9633 33979 9685 33995
rect 9633 33911 9685 33927
rect 9633 33853 9685 33859
rect 9725 34047 9777 35967
rect 9725 33979 9777 33995
rect 9725 33911 9777 33927
rect 6797 31271 6829 31323
rect 6745 31255 6829 31271
rect 6797 31203 6829 31255
rect 6745 31187 6829 31203
rect 6797 31135 6829 31187
rect 6745 29215 6829 31135
rect 9633 31323 9685 31329
rect 9633 31255 9685 31271
rect 9633 31187 9685 31203
rect 9633 31129 9685 31135
rect 9725 31323 9777 33859
rect 9725 31255 9777 31271
rect 9725 31187 9777 31203
rect 6797 29163 6829 29215
rect 6745 29147 6829 29163
rect 6797 29095 6829 29147
rect 6745 29079 6829 29095
rect 6797 29027 6829 29079
rect 5854 28768 5906 28774
rect 5854 28704 5906 28716
tri 5670 4702 5704 4736 sw
rect 5854 4684 5906 28652
rect 6090 27046 6142 27052
rect 6090 26982 6142 26994
tri 5906 4702 5940 4736 sw
rect 6090 4684 6142 26930
rect 6745 26491 6829 29027
rect 9633 29215 9685 29221
rect 9633 29147 9685 29163
rect 9633 29079 9685 29095
rect 9633 29021 9685 29027
rect 9725 29215 9777 31135
rect 9725 29147 9777 29163
rect 9725 29079 9777 29095
rect 6797 26439 6829 26491
rect 6745 26423 6829 26439
rect 6797 26371 6829 26423
rect 6745 26355 6829 26371
rect 6797 26303 6829 26355
rect 6745 24383 6829 26303
rect 9633 26491 9685 26497
rect 9633 26423 9685 26439
rect 9633 26355 9685 26371
rect 9633 26297 9685 26303
rect 9725 26491 9777 29027
rect 9725 26423 9777 26439
rect 9725 26355 9777 26371
rect 6797 24331 6829 24383
rect 6745 24315 6829 24331
rect 6797 24263 6829 24315
rect 6745 24247 6829 24263
rect 6797 24195 6829 24247
rect 6326 24012 6378 24018
rect 6326 23948 6378 23960
tri 6142 4702 6176 4736 sw
rect 6326 4684 6378 23896
rect 6562 22214 6614 22220
rect 6562 22150 6614 22162
tri 6378 4702 6412 4736 sw
rect 6562 4684 6614 22098
rect 6745 21659 6829 24195
rect 9633 24383 9685 24389
rect 9633 24315 9685 24331
rect 9633 24247 9685 24263
rect 9633 24189 9685 24195
rect 9725 24383 9777 26303
rect 9725 24315 9777 24331
rect 9725 24247 9777 24263
rect 6797 21607 6829 21659
rect 6745 21591 6829 21607
rect 6797 21539 6829 21591
rect 6745 21523 6829 21539
rect 6797 21471 6829 21523
rect 6745 19551 6829 21471
rect 9633 21659 9685 21665
rect 9633 21591 9685 21607
rect 9633 21523 9685 21539
rect 9633 21465 9685 21471
rect 9725 21659 9777 24195
rect 9725 21591 9777 21607
rect 9725 21523 9777 21539
rect 6797 19499 6829 19551
rect 6745 19483 6829 19499
rect 6797 19431 6829 19483
rect 6745 19415 6829 19431
rect 6797 19363 6829 19415
rect 6745 16827 6829 19363
rect 6797 16775 6829 16827
rect 6745 16759 6829 16775
rect 6797 16707 6829 16759
rect 6745 16691 6829 16707
rect 6797 16639 6829 16691
rect 6745 14719 6829 16639
rect 9633 16827 9685 16833
rect 9633 16759 9685 16775
rect 9633 16691 9685 16707
rect 9633 16633 9685 16639
rect 9725 16827 9777 21471
rect 10860 38879 10912 39919
tri 10912 39886 10946 39920 nw
tri 12024 39886 12058 39920 ne
rect 10860 38811 10912 38827
rect 10860 38743 10912 38759
rect 10860 36155 10912 38691
rect 10860 36087 10912 36103
rect 10860 36019 10912 36035
rect 10860 34047 10912 35967
rect 10860 33979 10912 33995
rect 10860 33911 10912 33927
rect 10860 31323 10912 33859
rect 10860 31255 10912 31271
rect 10860 31187 10912 31203
rect 10860 29215 10912 31135
rect 10860 29147 10912 29163
rect 10860 29079 10912 29095
rect 10860 26491 10912 29027
rect 10860 26423 10912 26439
rect 10860 26355 10912 26371
rect 10860 24383 10912 26303
rect 10860 24315 10912 24331
rect 10860 24247 10912 24263
rect 10860 21659 10912 24195
rect 10860 21591 10912 21607
rect 10860 21523 10912 21539
rect 9725 16759 9777 16775
rect 9725 16691 9777 16707
rect 6797 14667 6829 14719
rect 6745 14651 6829 14667
rect 6797 14599 6829 14651
rect 6745 14583 6829 14599
rect 6797 14531 6829 14583
rect 6745 11995 6829 14531
rect 9633 14719 9685 14725
rect 9633 14651 9685 14667
rect 9633 14583 9685 14599
rect 9633 14525 9685 14531
rect 9725 14719 9777 16639
rect 9725 14651 9777 14667
rect 9725 14583 9777 14599
rect 6797 11943 6829 11995
rect 6745 11927 6829 11943
rect 6797 11875 6829 11927
rect 6745 11859 6829 11875
rect 6797 11807 6829 11859
rect 6745 9887 6829 11807
rect 9633 11995 9685 12001
rect 9633 11927 9685 11943
rect 9633 11859 9685 11875
rect 9633 11801 9685 11807
rect 9725 11995 9777 14531
rect 9725 11927 9777 11943
rect 9725 11859 9777 11875
rect 6797 9835 6829 9887
rect 6745 9819 6829 9835
rect 6797 9767 6829 9819
rect 6745 9751 6829 9767
rect 6797 9699 6829 9751
tri 4658 4422 4692 4456 sw
tri 6711 4422 6745 4456 se
rect 6745 4376 6829 9699
rect 9633 9887 9685 9893
rect 9633 9819 9685 9835
rect 9633 9751 9685 9767
rect 9633 9693 9685 9699
rect 9725 9887 9777 11807
rect 9725 9819 9777 9835
rect 9725 9751 9777 9767
rect 9633 7163 9685 7169
rect 9633 7095 9685 7111
rect 9633 7027 9685 7043
rect 9633 6969 9685 6975
rect 7887 6188 7939 6194
rect 7887 6124 7939 6136
rect 7887 6066 7939 6072
rect 8287 5303 8339 5309
rect 8287 5239 8339 5251
rect 8287 5181 8339 5187
rect 8367 5147 8419 5153
rect 8367 5083 8419 5095
rect 7967 5067 8019 5073
rect 8367 5025 8419 5031
rect 7967 5003 8019 5015
rect 7967 4945 8019 4951
rect 8447 4987 8499 4993
rect 8447 4923 8499 4935
rect 8447 4865 8499 4871
rect 8047 4824 8099 4830
rect 8047 4760 8099 4772
rect 8047 4702 8099 4708
tri 6795 4375 6796 4376 ne
rect 6796 4375 6829 4376
rect 9725 4375 9777 9699
rect 9966 18727 10018 18733
rect 9966 18663 10018 18675
rect 9966 4684 10018 18611
rect 10202 17759 10254 17765
rect 10202 17695 10254 17707
tri 10018 4702 10052 4736 sw
rect 10202 4684 10254 17643
rect 10860 16827 10912 21471
rect 10860 16759 10912 16775
rect 10860 16691 10912 16707
rect 10860 14719 10912 16639
rect 10860 14651 10912 14667
rect 10860 14583 10912 14599
rect 10438 13895 10490 13901
rect 10438 13831 10490 13843
tri 10254 4702 10288 4736 sw
rect 10438 4684 10490 13779
rect 10674 12927 10726 12933
rect 10674 12863 10726 12875
tri 10490 4702 10524 4736 sw
rect 10674 4684 10726 12811
rect 10860 11995 10912 14531
rect 10860 11927 10912 11943
rect 10860 11859 10912 11875
rect 10860 9887 10912 11807
rect 10860 9819 10912 9835
rect 10860 9751 10912 9767
tri 9777 4421 9811 4455 sw
tri 10826 4421 10860 4455 se
rect 10860 4376 10912 9699
rect 12058 38879 12110 39965
tri 12110 39886 12144 39920 nw
tri 13812 39886 13846 39920 ne
rect 12058 38811 12110 38827
rect 12058 38743 12110 38759
rect 12058 36155 12110 38691
rect 12058 36087 12110 36103
rect 12058 36019 12110 36035
rect 12058 34047 12110 35967
rect 12058 33979 12110 33995
rect 12058 33911 12110 33927
rect 12058 31323 12110 33859
rect 12058 31255 12110 31271
rect 12058 31187 12110 31203
rect 12058 29215 12110 31135
rect 12058 29147 12110 29163
rect 12058 29079 12110 29095
rect 12058 26491 12110 29027
rect 12058 26423 12110 26439
rect 12058 26355 12110 26371
rect 12058 24383 12110 26303
rect 12058 24315 12110 24331
rect 12058 24247 12110 24263
rect 12058 21659 12110 24195
rect 12058 21591 12110 21607
rect 12058 21523 12110 21539
rect 12058 16827 12110 21471
rect 12058 16759 12110 16775
rect 12058 16691 12110 16707
rect 12058 14719 12110 16639
rect 12058 14651 12110 14667
rect 12058 14583 12110 14599
rect 12058 11995 12110 14531
rect 12058 11927 12110 11943
rect 12058 11859 12110 11875
rect 12058 9887 12110 11807
rect 12058 9819 12110 9835
rect 12058 9751 12110 9767
rect 11164 9063 11216 9069
rect 11164 8999 11216 9011
rect 11164 4684 11216 8947
rect 11400 8095 11452 8101
rect 11400 8031 11452 8043
tri 11216 4702 11250 4736 sw
rect 11400 4684 11452 7979
tri 11452 4702 11486 4736 sw
rect 11694 4694 11746 4700
rect 11694 4630 11746 4642
rect 11694 4572 11746 4578
tri 10912 4421 10946 4455 sw
tri 12024 4421 12058 4455 se
rect 12058 4375 12110 9699
rect 13846 38879 13898 39965
tri 13898 39886 13932 39920 nw
tri 15537 39886 15571 39920 ne
rect 13846 38811 13898 38827
rect 13846 38743 13898 38759
rect 13846 36155 13898 38691
rect 13846 36087 13898 36103
rect 13846 36019 13898 36035
rect 13846 34047 13898 35967
rect 13846 33979 13898 33995
rect 13846 33911 13898 33927
rect 13846 31323 13898 33859
rect 13846 31255 13898 31271
rect 13846 31187 13898 31203
rect 13846 29215 13898 31135
rect 13846 29147 13898 29163
rect 13846 29079 13898 29095
rect 13846 26491 13898 29027
rect 13846 26423 13898 26439
rect 13846 26355 13898 26371
rect 13846 24383 13898 26303
rect 13846 24315 13898 24331
rect 13846 24247 13898 24263
rect 13846 21659 13898 24195
rect 13846 21591 13898 21607
rect 13846 21523 13898 21539
rect 13846 16827 13898 21471
rect 13846 16759 13898 16775
rect 13846 16691 13898 16707
rect 13846 14719 13898 16639
rect 13846 14651 13898 14667
rect 13846 14583 13898 14599
rect 13846 11995 13898 14531
rect 13846 11927 13898 11943
rect 13846 11859 13898 11875
rect 13846 9887 13898 11807
rect 13846 9819 13898 9835
rect 13846 9751 13898 9767
tri 6796 4342 6829 4375 ne
tri 12024 4342 12057 4375 ne
rect 12057 4342 12110 4375
tri 12057 4341 12058 4342 ne
rect 9847 4268 9853 4320
rect 9905 4268 9917 4320
rect 9969 4268 9975 4320
rect 6669 4187 6675 4239
rect 6727 4187 6739 4239
rect 6791 4187 6797 4239
tri 6711 4153 6745 4187 ne
rect 5336 3964 5574 3965
rect 5336 3912 5342 3964
rect 5394 3912 5429 3964
rect 5481 3912 5516 3964
rect 5568 3912 5574 3964
rect 5336 3890 5574 3912
rect 5336 3838 5342 3890
rect 5394 3838 5429 3890
rect 5481 3838 5516 3890
rect 5568 3838 5574 3890
rect 6484 3958 6684 3964
rect 6536 3906 6558 3958
rect 6610 3906 6632 3958
rect 6484 3890 6684 3906
rect 6536 3838 6558 3890
rect 6610 3838 6632 3890
rect 5336 3816 5574 3838
rect 5336 3764 5342 3816
rect 5394 3764 5429 3816
rect 5481 3764 5516 3816
rect 5568 3764 5574 3816
tri 6450 3804 6484 3838 se
rect 6484 3821 6684 3838
rect 6536 3769 6558 3821
rect 6610 3769 6632 3821
rect 5336 3763 5574 3764
rect 547 3683 553 3735
rect 605 3683 621 3735
rect 673 3683 688 3735
rect 740 3683 755 3735
rect 807 3683 822 3735
rect 874 3683 889 3735
rect 941 3683 1420 3735
rect 547 3657 1420 3683
rect 547 3605 553 3657
rect 605 3605 621 3657
rect 673 3605 688 3657
rect 740 3605 755 3657
rect 807 3605 822 3657
rect 874 3605 889 3657
rect 941 3605 1420 3657
rect 979 3410 1481 3416
rect 1031 3364 1481 3410
rect 3016 3397 3341 3449
rect 3393 3397 3405 3449
rect 3457 3397 3463 3449
rect 3531 3397 3856 3449
rect 3908 3397 3920 3449
rect 3972 3397 3978 3449
rect 5417 3364 5423 3416
rect 5475 3364 5487 3416
rect 5539 3364 5545 3416
rect 979 3346 1031 3358
tri 1031 3330 1065 3364 nw
rect 979 3288 1031 3294
rect 3243 3080 3249 3132
rect 3301 3080 3313 3132
rect 3365 3080 3371 3132
rect 3531 3080 3537 3132
rect 3589 3080 3601 3132
rect 3653 3080 3659 3132
rect 5416 2961 5574 2967
rect 5468 2909 5522 2961
rect 5416 2894 5574 2909
rect 5468 2842 5522 2894
rect 5416 2826 5574 2842
rect 5468 2774 5522 2826
rect 5416 2768 5574 2774
rect 547 2219 553 2271
rect 605 2219 621 2271
rect 673 2219 688 2271
rect 740 2219 755 2271
rect 807 2219 822 2271
rect 874 2219 889 2271
rect 941 2219 1420 2271
rect 547 2197 1420 2219
rect 547 2145 553 2197
rect 605 2145 621 2197
rect 673 2145 688 2197
rect 740 2145 755 2197
rect 807 2145 822 2197
rect 874 2145 889 2197
rect 941 2145 1420 2197
rect 547 2123 1420 2145
rect 547 2071 553 2123
rect 605 2071 621 2123
rect 673 2071 688 2123
rect 740 2071 755 2123
rect 807 2071 822 2123
rect 874 2071 889 2123
rect 941 2071 1420 2123
rect 547 2070 1420 2071
rect 547 1962 553 2014
rect 605 1962 621 2014
rect 673 1962 688 2014
rect 740 1962 755 2014
rect 807 1962 822 2014
rect 874 1962 889 2014
rect 941 1962 1420 2014
rect 547 1940 1420 1962
rect 547 1888 553 1940
rect 605 1888 621 1940
rect 673 1888 688 1940
rect 740 1888 755 1940
rect 807 1888 822 1940
rect 874 1888 889 1940
rect 941 1888 1420 1940
rect 547 1866 1420 1888
rect 5818 1937 5870 3764
rect 6484 3763 6684 3769
rect 6745 3339 6797 4187
tri 9793 3999 9847 4053 se
rect 9847 4031 9899 4268
tri 9899 4234 9933 4268 nw
rect 9847 3999 9867 4031
tri 9867 3999 9899 4031 nw
rect 8127 3525 8179 3531
rect 8127 3461 8179 3473
rect 8127 3403 8179 3409
rect 6745 3275 6797 3287
rect 6745 3217 6797 3223
rect 9793 3339 9845 3999
tri 9845 3977 9867 3999 nw
rect 11899 3486 11951 3492
rect 9917 3403 9923 3455
rect 9975 3403 9987 3455
rect 10039 3403 10364 3455
tri 11865 3416 11899 3450 se
rect 11899 3422 11951 3434
rect 11899 3364 11951 3370
rect 9793 3275 9845 3287
rect 9793 3217 9845 3223
rect 9917 3080 9923 3132
rect 9975 3080 9987 3132
rect 10039 3080 10045 3132
rect 6745 3001 6797 3007
rect 6745 2937 6797 2949
rect 6484 2587 6684 2593
rect 6536 2535 6558 2587
rect 6610 2535 6632 2587
rect 6484 2519 6684 2535
rect 6536 2467 6558 2519
rect 6610 2467 6632 2519
rect 6484 2451 6684 2467
rect 6536 2399 6558 2451
rect 6610 2399 6632 2451
rect 6484 2393 6684 2399
tri 6450 2164 6484 2198 ne
tri 5870 1937 5946 2013 sw
rect 5818 1885 5824 1937
rect 5876 1885 5888 1937
rect 5940 1885 5946 1937
rect 547 1814 553 1866
rect 605 1814 621 1866
rect 673 1814 688 1866
rect 740 1814 755 1866
rect 807 1814 822 1866
rect 874 1814 889 1866
rect 941 1814 1420 1866
rect 547 1813 1420 1814
tri 6420 1813 6484 1877 se
rect 6484 1813 6684 2204
tri 6280 1673 6420 1813 se
rect 6420 1673 6684 1813
tri 6684 1673 6714 1703 sw
rect 6484 1470 6684 1673
rect 6347 1056 6399 1064
rect 3151 952 3157 1004
rect 3209 952 3221 1004
rect 3273 952 3279 1004
rect 3707 952 3713 1004
rect 3765 952 3777 1004
rect 3829 952 3835 1004
rect 6347 992 6399 1004
rect 6347 934 6399 940
rect 6547 1056 6599 1062
rect 6547 992 6599 1004
rect 6547 931 6599 940
rect 1231 668 1237 720
rect 1289 668 1301 720
rect 1353 668 1513 720
rect 3068 680 3074 681
rect 3016 629 3074 680
rect 3126 629 3138 681
rect 3190 680 3196 681
rect 3190 629 3463 680
rect 3531 635 3856 687
rect 3908 635 3920 687
rect 3972 635 3978 687
rect 5476 668 5528 720
tri 5442 664 5446 668 ne
rect 5446 664 5528 668
tri 5446 635 5475 664 ne
rect 5475 635 5528 664
tri 5475 634 5476 635 ne
rect 5476 630 5528 635
tri 5528 630 5531 633 sw
rect 5476 599 5531 630
tri 5531 599 5562 630 sw
rect 5476 547 5482 599
rect 5534 547 5546 599
rect 5598 547 5604 599
rect 5983 547 5989 599
rect 6041 547 6053 599
rect 6105 547 6111 599
tri 6025 513 6059 547 ne
rect 547 427 553 479
rect 605 427 621 479
rect 673 427 688 479
rect 740 427 755 479
rect 807 427 822 479
rect 874 427 889 479
rect 941 427 1420 479
rect 547 401 1420 427
rect 547 349 553 401
rect 605 349 621 401
rect 673 349 688 401
rect 740 349 755 401
rect 807 349 822 401
rect 874 349 889 401
rect 941 349 1420 401
rect 979 122 1031 128
rect 979 58 1031 70
rect 979 0 1031 6
rect 1231 122 1283 128
rect 1231 58 1283 70
rect 1231 0 1283 6
rect 6059 122 6111 547
rect 6059 58 6111 70
rect 6059 0 6111 6
rect 6347 459 6399 465
rect 6347 395 6399 407
rect 6347 122 6399 343
rect 6347 58 6399 70
rect 6347 0 6399 6
rect 6547 459 6599 465
rect 6547 395 6599 407
rect 6547 122 6599 343
rect 6547 58 6599 70
rect 6547 0 6599 6
rect 6745 122 6797 2885
rect 8527 2870 8579 2876
rect 8527 2806 8579 2818
rect 8527 2748 8579 2754
rect 6840 1305 6847 1326
tri 7171 1309 7172 1310 se
tri 7172 1309 7173 1310 sw
rect 6829 1002 6857 1278
rect 6885 1158 6937 1282
rect 7021 1252 7185 1303
tri 6937 1158 6971 1192 sw
rect 6885 1134 7014 1158
rect 6885 1082 6891 1134
rect 6943 1082 6956 1134
rect 7008 1082 7014 1134
rect 6885 1058 7014 1082
rect 7393 1024 7445 1030
tri 7359 916 7393 950 se
rect 7393 928 7445 972
rect 7135 910 7393 916
tri 7445 916 7479 950 sw
rect 7445 910 8035 916
rect 7135 876 7219 910
rect 7253 876 7297 910
rect 7331 876 7375 910
rect 7445 876 7453 910
rect 7487 876 7531 910
rect 7565 876 7609 910
rect 7643 876 7687 910
rect 7721 876 7765 910
rect 7799 876 7835 910
rect 7135 870 7835 876
rect 7135 863 7208 870
tri 7208 863 7215 870 nw
tri 7343 863 7350 870 ne
rect 7350 863 7835 870
rect 7135 838 7181 863
rect 7135 804 7141 838
rect 7175 804 7181 838
tri 7181 836 7208 863 nw
tri 7350 836 7377 863 ne
rect 7377 858 7835 863
rect 7887 858 7909 910
rect 7961 858 7983 910
rect 7135 751 7181 804
rect 7135 717 7141 751
rect 7175 717 7181 751
rect 7377 832 8035 858
rect 7377 803 7995 832
rect 8029 803 8035 832
rect 7377 788 7835 803
rect 7887 788 7909 803
rect 7377 754 7389 788
rect 7423 754 7469 788
rect 7503 754 7549 788
rect 7583 754 7629 788
rect 7663 754 7709 788
rect 7743 754 7789 788
rect 7823 754 7835 788
rect 7903 754 7909 788
rect 7377 751 7835 754
rect 7887 751 7909 754
rect 7961 751 7983 803
rect 7377 748 7995 751
tri 7801 734 7815 748 ne
rect 7815 734 7995 748
rect 7135 664 7181 717
rect 7135 630 7141 664
rect 7175 630 7181 664
rect 7135 577 7181 630
rect 7135 543 7141 577
rect 7175 543 7181 577
rect 7135 452 7181 543
rect 7224 722 7276 734
rect 7224 688 7233 722
rect 7267 688 7276 722
tri 7815 720 7829 734 ne
rect 7829 720 7995 734
rect 8029 720 8035 751
tri 7829 714 7835 720 ne
rect 7224 631 7276 688
rect 7835 696 8035 720
rect 7887 644 7909 696
rect 7961 644 7983 696
rect 7835 641 7995 644
rect 8029 641 8035 644
rect 7224 601 7233 631
rect 7267 601 7276 631
rect 7315 632 7503 641
rect 7315 598 7327 632
rect 7361 598 7412 632
rect 7446 598 7497 632
rect 7315 589 7503 598
rect 7555 589 7567 641
rect 7619 632 7795 641
rect 7619 598 7665 632
rect 7699 598 7749 632
rect 7783 598 7795 632
rect 7619 589 7795 598
rect 7835 596 8035 641
rect 8207 757 8259 1278
rect 8607 1002 8659 1278
tri 9519 1158 9553 1192 se
rect 9553 1158 9605 1285
rect 9476 1134 9605 1158
rect 9476 1082 9482 1134
rect 9534 1082 9547 1134
rect 9599 1082 9605 1134
rect 9476 1058 9605 1082
rect 9633 1237 9685 1281
tri 9685 1237 9700 1252 sw
rect 12058 1237 12110 4342
rect 12636 7727 12836 7746
rect 12636 7675 12642 7727
rect 12694 7675 12710 7727
rect 12762 7675 12778 7727
rect 12830 7675 12836 7727
rect 12636 2961 12836 7675
rect 12636 2909 12637 2961
rect 12689 2909 12709 2961
rect 12761 2909 12781 2961
rect 12833 2909 12836 2961
rect 12636 2894 12836 2909
rect 12636 2842 12637 2894
rect 12689 2842 12709 2894
rect 12761 2842 12781 2894
rect 12833 2842 12836 2894
rect 12636 2826 12836 2842
rect 12636 2774 12637 2826
rect 12689 2774 12709 2826
rect 12761 2774 12781 2826
rect 12833 2774 12836 2826
rect 12636 1795 12836 2774
rect 12636 1743 12642 1795
rect 12694 1743 12710 1795
rect 12762 1743 12778 1795
rect 12830 1743 12836 1795
rect 12636 1723 12836 1743
rect 12636 1671 12642 1723
rect 12694 1671 12710 1723
rect 12762 1671 12778 1723
rect 12830 1671 12836 1723
rect 12636 1651 12836 1671
rect 12636 1599 12642 1651
rect 12694 1599 12710 1651
rect 12762 1599 12778 1651
rect 12830 1599 12836 1651
rect 12636 1598 12836 1599
tri 12110 1283 12144 1317 sw
tri 13812 1283 13846 1317 se
rect 13846 1237 13898 9699
rect 15571 38879 15623 39965
rect 15571 38811 15623 38827
rect 15571 38743 15623 38759
rect 15571 36155 15623 38691
rect 15571 36087 15623 36103
rect 15571 36019 15623 36035
rect 15571 34047 15623 35967
rect 15571 33979 15623 33995
rect 15571 33911 15623 33927
rect 15571 31323 15623 33859
rect 15571 31255 15623 31271
rect 15571 31187 15623 31203
rect 15571 29215 15623 31135
rect 15571 29147 15623 29163
rect 15571 29079 15623 29095
rect 15571 26491 15623 29027
rect 15571 26423 15623 26439
rect 15571 26355 15623 26371
rect 15571 24383 15623 26303
rect 15571 24315 15623 24331
rect 15571 24247 15623 24263
rect 15571 21659 15623 24195
rect 15571 21591 15623 21607
rect 15571 21523 15623 21539
rect 15571 16827 15623 21471
rect 15571 16759 15623 16775
rect 15571 16691 15623 16707
rect 15571 14719 15623 16639
rect 15571 14651 15623 14667
rect 15571 14583 15623 14599
rect 15571 11995 15623 14531
rect 15571 11927 15623 11943
rect 15571 11859 15623 11875
rect 15571 9887 15623 11807
rect 15571 9819 15623 9835
rect 15571 9751 15623 9767
tri 13898 1283 13932 1317 sw
tri 15537 1283 15571 1317 se
rect 15571 1237 15623 9699
rect 9633 1218 9700 1237
tri 9700 1218 9719 1237 sw
rect 9633 1212 9737 1218
rect 9633 1160 9685 1212
rect 9633 1136 9737 1160
rect 9633 1084 9685 1136
rect 9633 1060 9737 1084
rect 9633 1008 9685 1060
tri 8659 1002 8661 1004 sw
rect 9633 1002 9737 1008
rect 13301 1022 13307 1074
rect 13359 1022 13375 1074
rect 13427 1022 13442 1074
rect 13494 1022 13509 1074
rect 13561 1022 13576 1074
rect 13628 1022 13643 1074
rect 13695 1022 13701 1074
rect 8607 970 8661 1002
tri 8661 970 8693 1002 sw
rect 8607 918 8613 970
rect 8665 918 8677 970
rect 8729 918 8735 970
rect 9917 952 9923 1004
rect 9975 952 9987 1004
rect 10039 952 10045 1004
rect 13301 988 13701 1022
rect 13301 936 13307 988
rect 13359 936 13375 988
rect 13427 936 13442 988
rect 13494 936 13509 988
rect 13561 936 13576 988
rect 13628 936 13643 988
rect 13695 936 13701 988
rect 13301 902 13701 936
rect 8207 693 8259 705
rect 8207 635 8259 641
rect 8304 863 8859 870
rect 8911 863 8927 870
rect 8304 829 8316 863
rect 8350 829 8393 863
rect 8427 829 8469 863
rect 8503 829 8545 863
rect 8579 829 8621 863
rect 8655 829 8697 863
rect 8731 829 8773 863
rect 8807 829 8849 863
rect 8911 829 8925 863
rect 8304 818 8859 829
rect 8911 818 8927 829
rect 8979 818 8994 870
rect 9046 818 9061 870
rect 9113 818 9128 870
rect 9180 863 9195 870
rect 9247 863 9262 870
rect 9314 863 9329 870
rect 9381 863 9396 870
rect 9448 863 9463 870
rect 9187 829 9195 863
rect 9448 829 9457 863
rect 9180 818 9195 829
rect 9247 818 9262 829
rect 9314 818 9329 829
rect 9381 818 9396 829
rect 9448 818 9463 829
rect 9515 818 9530 870
rect 9582 818 9597 870
rect 9649 818 9655 870
rect 13301 850 13307 902
rect 13359 850 13375 902
rect 13427 850 13442 902
rect 13494 850 13509 902
rect 13561 850 13576 902
rect 13628 850 13643 902
rect 13695 850 13701 902
rect 13301 849 13701 850
rect 8304 806 9655 818
rect 8304 785 8859 806
rect 8911 785 8927 806
rect 8304 751 8316 785
rect 8350 751 8393 785
rect 8427 751 8469 785
rect 8503 751 8545 785
rect 8579 751 8621 785
rect 8655 751 8697 785
rect 8731 751 8773 785
rect 8807 751 8849 785
rect 8911 754 8925 785
rect 8979 754 8994 806
rect 9046 754 9061 806
rect 9113 754 9128 806
rect 9180 785 9195 806
rect 9247 785 9262 806
rect 9314 785 9329 806
rect 9381 785 9396 806
rect 9448 785 9463 806
rect 9187 754 9195 785
rect 9448 754 9457 785
rect 9515 754 9530 806
rect 9582 754 9597 806
rect 9649 754 9655 806
rect 8883 751 8925 754
rect 8959 751 9001 754
rect 9035 751 9077 754
rect 9111 751 9153 754
rect 9187 751 9229 754
rect 9263 751 9305 754
rect 9339 751 9381 754
rect 9415 751 9457 754
rect 9491 751 9533 754
rect 9567 751 9609 754
rect 9643 751 9655 754
rect 8304 707 9655 751
rect 8304 673 8316 707
rect 8350 673 8393 707
rect 8427 673 8469 707
rect 8503 673 8545 707
rect 8579 673 8621 707
rect 8655 673 8697 707
rect 8731 673 8773 707
rect 8807 673 8849 707
rect 8883 673 8925 707
rect 8959 673 9001 707
rect 9035 673 9077 707
rect 9111 673 9153 707
rect 9187 673 9229 707
rect 9263 673 9305 707
rect 9339 673 9381 707
rect 9415 673 9457 707
rect 9491 673 9533 707
rect 9567 673 9609 707
rect 9643 673 9655 707
rect 7224 539 7276 549
rect 7224 537 7233 539
rect 7267 537 7276 539
rect 7835 588 7995 596
rect 8029 588 8035 596
rect 7887 536 7909 588
rect 7961 536 7983 588
rect 7835 517 8035 536
rect 7224 479 7276 485
tri 7802 483 7835 516 se
rect 7835 483 7995 517
rect 8029 483 8035 517
tri 7801 482 7802 483 se
rect 7802 482 8035 483
rect 7377 480 8035 482
rect 7135 418 7141 452
rect 7175 418 7181 452
rect 7135 361 7181 418
rect 7377 476 7835 480
rect 7887 476 7909 480
rect 7377 442 7389 476
rect 7423 442 7469 476
rect 7503 442 7549 476
rect 7583 442 7629 476
rect 7663 442 7709 476
rect 7743 442 7789 476
rect 7823 442 7835 476
rect 7903 442 7909 476
rect 7377 428 7835 442
rect 7887 428 7909 442
rect 7961 428 7983 480
tri 7181 361 7214 394 sw
tri 7344 361 7377 394 se
rect 7377 372 8035 428
rect 7377 361 7835 372
rect 7135 360 7214 361
tri 7214 360 7215 361 sw
tri 7343 360 7344 361 se
rect 7344 360 7835 361
rect 7135 354 7835 360
rect 7135 320 7219 354
rect 7253 320 7297 354
rect 7331 320 7375 354
rect 7409 320 7453 354
rect 7487 320 7531 354
rect 7565 320 7609 354
rect 7643 320 7687 354
rect 7721 320 7765 354
rect 7799 320 7835 354
rect 7887 320 7909 372
rect 7961 320 7983 372
rect 8304 629 9655 673
rect 9917 635 9923 687
rect 9975 635 9987 687
rect 10039 635 10364 687
rect 11899 668 12080 720
tri 12058 667 12059 668 ne
rect 12059 667 12080 668
tri 12059 658 12068 667 ne
rect 12068 658 12080 667
tri 12068 646 12080 658 ne
tri 12080 649 12151 720 sw
rect 12080 646 12151 649
rect 8304 595 8316 629
rect 8350 595 8393 629
rect 8427 595 8469 629
rect 8503 595 8545 629
rect 8579 595 8621 629
rect 8655 595 8697 629
rect 8731 595 8773 629
rect 8807 595 8849 629
rect 8883 595 8925 629
rect 8959 595 9001 629
rect 9035 595 9077 629
rect 9111 595 9153 629
rect 9187 595 9229 629
rect 9263 595 9305 629
rect 9339 595 9381 629
rect 9415 595 9457 629
rect 9491 595 9533 629
rect 9567 595 9609 629
rect 9643 595 9655 629
tri 12080 627 12099 646 ne
rect 8304 551 9655 595
rect 8304 517 8316 551
rect 8350 517 8393 551
rect 8427 517 8469 551
rect 8503 517 8545 551
rect 8579 517 8621 551
rect 8655 517 8697 551
rect 8731 517 8773 551
rect 8807 517 8849 551
rect 8883 517 8925 551
rect 8959 517 9001 551
rect 9035 517 9077 551
rect 9111 517 9153 551
rect 9187 517 9229 551
rect 9263 517 9305 551
rect 9339 517 9381 551
rect 9415 517 9457 551
rect 9491 517 9533 551
rect 9567 517 9609 551
rect 9643 517 9655 551
rect 8304 473 9655 517
rect 8304 439 8316 473
rect 8350 439 8393 473
rect 8427 439 8469 473
rect 8503 439 8545 473
rect 8579 439 8621 473
rect 8655 439 8697 473
rect 8731 439 8773 473
rect 8807 439 8849 473
rect 8883 439 8925 473
rect 8959 439 9001 473
rect 9035 439 9077 473
rect 9111 439 9153 473
rect 9187 439 9229 473
rect 9263 439 9305 473
rect 9339 439 9381 473
rect 9415 439 9457 473
rect 9491 439 9533 473
rect 9567 439 9609 473
rect 9643 439 9655 473
rect 8304 395 9655 439
rect 8304 361 8316 395
rect 8350 361 8393 395
rect 8427 361 8469 395
rect 8503 361 8545 395
rect 8579 361 8621 395
rect 8655 361 8697 395
rect 8731 361 8773 395
rect 8807 361 8849 395
rect 8883 361 8925 395
rect 8959 361 9001 395
rect 9035 361 9077 395
rect 9111 361 9153 395
rect 9187 361 9229 395
rect 9263 361 9305 395
rect 9339 361 9381 395
rect 9415 361 9457 395
rect 9491 361 9533 395
rect 9567 361 9609 395
rect 9643 361 9655 395
rect 8304 354 9655 361
rect 7135 314 8035 320
rect 8333 320 9883 321
rect 8333 268 8339 320
rect 8391 268 8407 320
rect 8459 268 8474 320
rect 8526 268 8541 320
rect 8593 268 8608 320
rect 8660 268 8675 320
rect 8727 268 9883 320
rect 8333 246 9883 268
rect 6874 161 6880 213
rect 6932 161 6944 213
rect 6996 161 8044 213
rect 8096 161 8108 213
rect 8160 161 8166 213
rect 8333 194 8339 246
rect 8391 194 8407 246
rect 8459 194 8474 246
rect 8526 194 8541 246
rect 8593 194 8608 246
rect 8660 194 8675 246
rect 8727 194 9883 246
rect 8333 172 9883 194
rect 6745 58 6797 70
rect 6745 0 6797 6
rect 7497 76 7503 128
rect 7555 76 7567 128
rect 7619 76 7625 128
rect 8333 120 8339 172
rect 8391 120 8407 172
rect 8459 120 8474 172
rect 8526 120 8541 172
rect 8593 120 8608 172
rect 8660 120 8675 172
rect 8727 120 9883 172
rect 8333 119 9883 120
rect 12099 122 12151 646
rect 12321 240 12327 292
rect 12379 240 12403 292
rect 12455 240 12479 292
rect 12531 240 12555 292
rect 12607 240 12631 292
rect 12683 240 12706 292
rect 12758 240 15367 292
rect 7497 52 7625 76
rect 7497 0 7503 52
rect 7555 0 7567 52
rect 7619 0 7625 52
rect 12099 58 12151 70
rect 12099 0 12151 6
rect 13080 122 13132 128
rect 13080 58 13132 70
rect 13080 0 13132 6
<< via1 >>
rect 385 38827 437 38879
rect 385 38759 437 38811
rect 385 38691 437 38743
rect 2464 38827 2516 38879
rect 2464 38759 2516 38811
rect 2464 38691 2516 38743
rect 385 36103 437 36155
rect 385 36035 437 36087
rect 385 35967 437 36019
rect 385 33995 437 34047
rect 385 33927 437 33979
rect 385 33859 437 33911
rect 385 31271 437 31323
rect 385 31203 437 31255
rect 385 31135 437 31187
rect 385 29163 437 29215
rect 385 29095 437 29147
rect 385 29027 437 29079
rect 385 26439 437 26491
rect 385 26371 437 26423
rect 385 26303 437 26355
rect 385 24331 437 24383
rect 385 24263 437 24315
rect 385 24195 437 24247
rect 385 21607 437 21659
rect 385 21539 437 21591
rect 385 21471 437 21523
rect 385 19499 437 19551
rect 385 19431 437 19483
rect 385 19363 437 19415
rect 385 16775 437 16827
rect 385 16707 437 16759
rect 385 16639 437 16691
rect 385 14667 437 14719
rect 385 14599 437 14651
rect 385 14531 437 14583
rect 385 11943 437 11995
rect 385 11875 437 11927
rect 385 11807 437 11859
rect 385 9835 437 9887
rect 385 9767 437 9819
rect 385 9699 437 9751
rect 626 38003 678 38055
rect 626 37939 678 37991
rect 862 37035 914 37087
rect 862 36971 914 37023
rect 2464 36103 2516 36155
rect 2464 36035 2516 36087
rect 2464 35967 2516 36019
rect 2464 33995 2516 34047
rect 2464 33927 2516 33979
rect 2464 33859 2516 33911
rect 1098 33171 1150 33223
rect 1098 33107 1150 33159
rect 1337 32203 1389 32255
rect 1337 32139 1389 32191
rect 2464 31271 2516 31323
rect 2464 31203 2516 31255
rect 2464 31135 2516 31187
rect 2464 29163 2516 29215
rect 2464 29095 2516 29147
rect 2464 29027 2516 29079
rect 1573 28339 1625 28391
rect 1573 28275 1625 28327
rect 1809 27371 1861 27423
rect 1809 27307 1861 27359
rect 2464 26439 2516 26491
rect 2464 26371 2516 26423
rect 2464 26303 2516 26355
rect 2464 24331 2516 24383
rect 2464 24263 2516 24315
rect 2464 24195 2516 24247
rect 2045 23507 2097 23559
rect 2045 23443 2097 23495
rect 2278 22539 2330 22591
rect 2278 22475 2330 22527
rect 2464 21607 2516 21659
rect 2464 21539 2516 21591
rect 2464 21471 2516 21523
rect 2464 19499 2516 19551
rect 2464 19431 2516 19483
rect 2464 19363 2516 19415
rect 4606 38827 4658 38879
rect 4606 38759 4658 38811
rect 4606 38691 4658 38743
rect 6745 38827 6797 38879
rect 6745 38759 6797 38811
rect 6745 38691 6797 38743
rect 4606 36103 4658 36155
rect 4606 36035 4658 36087
rect 4606 35967 4658 36019
rect 4606 33995 4658 34047
rect 4606 33927 4658 33979
rect 4606 33859 4658 33911
rect 4606 31271 4658 31323
rect 4606 31203 4658 31255
rect 4606 31135 4658 31187
rect 4606 29163 4658 29215
rect 4606 29095 4658 29147
rect 4606 29027 4658 29079
rect 4606 26439 4658 26491
rect 4606 26371 4658 26423
rect 4606 26303 4658 26355
rect 4606 24331 4658 24383
rect 4606 24263 4658 24315
rect 4606 24195 4658 24247
rect 4606 21607 4658 21659
rect 4606 21539 4658 21591
rect 4606 21471 4658 21523
rect 4606 19499 4658 19551
rect 4606 19431 4658 19483
rect 4606 19363 4658 19415
rect 2464 16775 2516 16827
rect 2464 16707 2516 16759
rect 2464 16639 2516 16691
rect 2464 14667 2516 14719
rect 2464 14599 2516 14651
rect 2464 14531 2516 14583
rect 2464 11943 2516 11995
rect 2464 11875 2516 11927
rect 2464 11807 2516 11859
rect 2464 9835 2516 9887
rect 2464 9767 2516 9819
rect 2464 9699 2516 9751
rect 2771 18675 2823 18727
rect 2771 18611 2823 18663
rect 3007 17707 3059 17759
rect 3007 17643 3059 17695
rect 4606 16775 4658 16827
rect 4606 16707 4658 16759
rect 4606 16639 4658 16691
rect 4606 14667 4658 14719
rect 4606 14599 4658 14651
rect 4606 14531 4658 14583
rect 3243 13843 3295 13895
rect 3243 13779 3295 13831
rect 3479 12875 3531 12927
rect 3479 12811 3531 12863
rect 4606 11943 4658 11995
rect 4606 11875 4658 11927
rect 4606 11807 4658 11859
rect 4606 9835 4658 9887
rect 4606 9767 4658 9819
rect 4606 9699 4658 9751
rect 3715 9011 3767 9063
rect 3715 8947 3767 8999
rect 3951 8043 4003 8095
rect 3951 7979 4003 8031
rect 4299 4643 4351 4695
rect 4299 4579 4351 4631
rect 4910 38380 4962 38432
rect 4910 38316 4962 38368
rect 5146 36658 5198 36710
rect 5146 36594 5198 36646
rect 9633 38827 9685 38879
rect 9633 38759 9685 38811
rect 9633 38691 9685 38743
rect 9725 38827 9777 38879
rect 9725 38759 9777 38811
rect 9725 38691 9777 38743
rect 6745 36103 6797 36155
rect 6745 36035 6797 36087
rect 6745 35967 6797 36019
rect 9633 36103 9685 36155
rect 9633 36035 9685 36087
rect 9633 35967 9685 36019
rect 9725 36103 9777 36155
rect 9725 36035 9777 36087
rect 9725 35967 9777 36019
rect 6745 33995 6797 34047
rect 6745 33927 6797 33979
rect 6745 33859 6797 33911
rect 5382 33548 5434 33600
rect 5382 33484 5434 33536
rect 5618 31826 5670 31878
rect 5618 31762 5670 31814
rect 9633 33995 9685 34047
rect 9633 33927 9685 33979
rect 9633 33859 9685 33911
rect 9725 33995 9777 34047
rect 9725 33927 9777 33979
rect 9725 33859 9777 33911
rect 6745 31271 6797 31323
rect 6745 31203 6797 31255
rect 6745 31135 6797 31187
rect 9633 31271 9685 31323
rect 9633 31203 9685 31255
rect 9633 31135 9685 31187
rect 9725 31271 9777 31323
rect 9725 31203 9777 31255
rect 9725 31135 9777 31187
rect 6745 29163 6797 29215
rect 6745 29095 6797 29147
rect 6745 29027 6797 29079
rect 5854 28716 5906 28768
rect 5854 28652 5906 28704
rect 6090 26994 6142 27046
rect 6090 26930 6142 26982
rect 9633 29163 9685 29215
rect 9633 29095 9685 29147
rect 9633 29027 9685 29079
rect 9725 29163 9777 29215
rect 9725 29095 9777 29147
rect 9725 29027 9777 29079
rect 6745 26439 6797 26491
rect 6745 26371 6797 26423
rect 6745 26303 6797 26355
rect 9633 26439 9685 26491
rect 9633 26371 9685 26423
rect 9633 26303 9685 26355
rect 9725 26439 9777 26491
rect 9725 26371 9777 26423
rect 9725 26303 9777 26355
rect 6745 24331 6797 24383
rect 6745 24263 6797 24315
rect 6745 24195 6797 24247
rect 6326 23960 6378 24012
rect 6326 23896 6378 23948
rect 6562 22162 6614 22214
rect 6562 22098 6614 22150
rect 9633 24331 9685 24383
rect 9633 24263 9685 24315
rect 9633 24195 9685 24247
rect 9725 24331 9777 24383
rect 9725 24263 9777 24315
rect 9725 24195 9777 24247
rect 6745 21607 6797 21659
rect 6745 21539 6797 21591
rect 6745 21471 6797 21523
rect 9633 21607 9685 21659
rect 9633 21539 9685 21591
rect 9633 21471 9685 21523
rect 9725 21607 9777 21659
rect 9725 21539 9777 21591
rect 9725 21471 9777 21523
rect 6745 19499 6797 19551
rect 6745 19431 6797 19483
rect 6745 19363 6797 19415
rect 6745 16775 6797 16827
rect 6745 16707 6797 16759
rect 6745 16639 6797 16691
rect 9633 16775 9685 16827
rect 9633 16707 9685 16759
rect 9633 16639 9685 16691
rect 10860 38827 10912 38879
rect 10860 38759 10912 38811
rect 10860 38691 10912 38743
rect 10860 36103 10912 36155
rect 10860 36035 10912 36087
rect 10860 35967 10912 36019
rect 10860 33995 10912 34047
rect 10860 33927 10912 33979
rect 10860 33859 10912 33911
rect 10860 31271 10912 31323
rect 10860 31203 10912 31255
rect 10860 31135 10912 31187
rect 10860 29163 10912 29215
rect 10860 29095 10912 29147
rect 10860 29027 10912 29079
rect 10860 26439 10912 26491
rect 10860 26371 10912 26423
rect 10860 26303 10912 26355
rect 10860 24331 10912 24383
rect 10860 24263 10912 24315
rect 10860 24195 10912 24247
rect 10860 21607 10912 21659
rect 10860 21539 10912 21591
rect 10860 21471 10912 21523
rect 9725 16775 9777 16827
rect 9725 16707 9777 16759
rect 9725 16639 9777 16691
rect 6745 14667 6797 14719
rect 6745 14599 6797 14651
rect 6745 14531 6797 14583
rect 9633 14667 9685 14719
rect 9633 14599 9685 14651
rect 9633 14531 9685 14583
rect 9725 14667 9777 14719
rect 9725 14599 9777 14651
rect 9725 14531 9777 14583
rect 6745 11943 6797 11995
rect 6745 11875 6797 11927
rect 6745 11807 6797 11859
rect 9633 11943 9685 11995
rect 9633 11875 9685 11927
rect 9633 11807 9685 11859
rect 9725 11943 9777 11995
rect 9725 11875 9777 11927
rect 9725 11807 9777 11859
rect 6745 9835 6797 9887
rect 6745 9767 6797 9819
rect 6745 9699 6797 9751
rect 9633 9835 9685 9887
rect 9633 9767 9685 9819
rect 9633 9699 9685 9751
rect 9725 9835 9777 9887
rect 9725 9767 9777 9819
rect 9725 9699 9777 9751
rect 9633 7111 9685 7163
rect 9633 7043 9685 7095
rect 9633 6975 9685 7027
rect 7887 6136 7939 6188
rect 7887 6072 7939 6124
rect 8287 5251 8339 5303
rect 8287 5187 8339 5239
rect 8367 5095 8419 5147
rect 7967 5015 8019 5067
rect 8367 5031 8419 5083
rect 7967 4951 8019 5003
rect 8447 4935 8499 4987
rect 8447 4871 8499 4923
rect 8047 4772 8099 4824
rect 8047 4708 8099 4760
rect 9966 18675 10018 18727
rect 9966 18611 10018 18663
rect 10202 17707 10254 17759
rect 10202 17643 10254 17695
rect 10860 16775 10912 16827
rect 10860 16707 10912 16759
rect 10860 16639 10912 16691
rect 10860 14667 10912 14719
rect 10860 14599 10912 14651
rect 10860 14531 10912 14583
rect 10438 13843 10490 13895
rect 10438 13779 10490 13831
rect 10674 12875 10726 12927
rect 10674 12811 10726 12863
rect 10860 11943 10912 11995
rect 10860 11875 10912 11927
rect 10860 11807 10912 11859
rect 10860 9835 10912 9887
rect 10860 9767 10912 9819
rect 10860 9699 10912 9751
rect 12058 38827 12110 38879
rect 12058 38759 12110 38811
rect 12058 38691 12110 38743
rect 12058 36103 12110 36155
rect 12058 36035 12110 36087
rect 12058 35967 12110 36019
rect 12058 33995 12110 34047
rect 12058 33927 12110 33979
rect 12058 33859 12110 33911
rect 12058 31271 12110 31323
rect 12058 31203 12110 31255
rect 12058 31135 12110 31187
rect 12058 29163 12110 29215
rect 12058 29095 12110 29147
rect 12058 29027 12110 29079
rect 12058 26439 12110 26491
rect 12058 26371 12110 26423
rect 12058 26303 12110 26355
rect 12058 24331 12110 24383
rect 12058 24263 12110 24315
rect 12058 24195 12110 24247
rect 12058 21607 12110 21659
rect 12058 21539 12110 21591
rect 12058 21471 12110 21523
rect 12058 16775 12110 16827
rect 12058 16707 12110 16759
rect 12058 16639 12110 16691
rect 12058 14667 12110 14719
rect 12058 14599 12110 14651
rect 12058 14531 12110 14583
rect 12058 11943 12110 11995
rect 12058 11875 12110 11927
rect 12058 11807 12110 11859
rect 12058 9835 12110 9887
rect 12058 9767 12110 9819
rect 12058 9699 12110 9751
rect 11164 9011 11216 9063
rect 11164 8947 11216 8999
rect 11400 8043 11452 8095
rect 11400 7979 11452 8031
rect 11694 4642 11746 4694
rect 11694 4578 11746 4630
rect 13846 38827 13898 38879
rect 13846 38759 13898 38811
rect 13846 38691 13898 38743
rect 13846 36103 13898 36155
rect 13846 36035 13898 36087
rect 13846 35967 13898 36019
rect 13846 33995 13898 34047
rect 13846 33927 13898 33979
rect 13846 33859 13898 33911
rect 13846 31271 13898 31323
rect 13846 31203 13898 31255
rect 13846 31135 13898 31187
rect 13846 29163 13898 29215
rect 13846 29095 13898 29147
rect 13846 29027 13898 29079
rect 13846 26439 13898 26491
rect 13846 26371 13898 26423
rect 13846 26303 13898 26355
rect 13846 24331 13898 24383
rect 13846 24263 13898 24315
rect 13846 24195 13898 24247
rect 13846 21607 13898 21659
rect 13846 21539 13898 21591
rect 13846 21471 13898 21523
rect 13846 16775 13898 16827
rect 13846 16707 13898 16759
rect 13846 16639 13898 16691
rect 13846 14667 13898 14719
rect 13846 14599 13898 14651
rect 13846 14531 13898 14583
rect 13846 11943 13898 11995
rect 13846 11875 13898 11927
rect 13846 11807 13898 11859
rect 13846 9835 13898 9887
rect 13846 9767 13898 9819
rect 13846 9699 13898 9751
rect 9853 4268 9905 4320
rect 9917 4268 9969 4320
rect 6675 4187 6727 4239
rect 6739 4187 6791 4239
rect 5342 3912 5394 3964
rect 5429 3912 5481 3964
rect 5516 3912 5568 3964
rect 5342 3838 5394 3890
rect 5429 3838 5481 3890
rect 5516 3838 5568 3890
rect 6484 3906 6536 3958
rect 6558 3906 6610 3958
rect 6632 3906 6684 3958
rect 6484 3838 6536 3890
rect 6558 3838 6610 3890
rect 6632 3838 6684 3890
rect 5342 3764 5394 3816
rect 5429 3764 5481 3816
rect 5516 3764 5568 3816
rect 6484 3769 6536 3821
rect 6558 3769 6610 3821
rect 6632 3769 6684 3821
rect 553 3683 605 3735
rect 621 3683 673 3735
rect 688 3683 740 3735
rect 755 3683 807 3735
rect 822 3683 874 3735
rect 889 3683 941 3735
rect 553 3605 605 3657
rect 621 3605 673 3657
rect 688 3605 740 3657
rect 755 3605 807 3657
rect 822 3605 874 3657
rect 889 3605 941 3657
rect 979 3358 1031 3410
rect 3341 3397 3393 3449
rect 3405 3397 3457 3449
rect 3856 3397 3908 3449
rect 3920 3397 3972 3449
rect 5423 3364 5475 3416
rect 5487 3364 5539 3416
rect 979 3294 1031 3346
rect 3249 3080 3301 3132
rect 3313 3080 3365 3132
rect 3537 3080 3589 3132
rect 3601 3080 3653 3132
rect 5416 2909 5468 2961
rect 5522 2909 5574 2961
rect 5416 2842 5468 2894
rect 5522 2842 5574 2894
rect 5416 2774 5468 2826
rect 5522 2774 5574 2826
rect 553 2219 605 2271
rect 621 2219 673 2271
rect 688 2219 740 2271
rect 755 2219 807 2271
rect 822 2219 874 2271
rect 889 2219 941 2271
rect 553 2145 605 2197
rect 621 2145 673 2197
rect 688 2145 740 2197
rect 755 2145 807 2197
rect 822 2145 874 2197
rect 889 2145 941 2197
rect 553 2071 605 2123
rect 621 2071 673 2123
rect 688 2071 740 2123
rect 755 2071 807 2123
rect 822 2071 874 2123
rect 889 2071 941 2123
rect 553 1962 605 2014
rect 621 1962 673 2014
rect 688 1962 740 2014
rect 755 1962 807 2014
rect 822 1962 874 2014
rect 889 1962 941 2014
rect 553 1888 605 1940
rect 621 1888 673 1940
rect 688 1888 740 1940
rect 755 1888 807 1940
rect 822 1888 874 1940
rect 889 1888 941 1940
rect 8127 3473 8179 3525
rect 8127 3409 8179 3461
rect 6745 3287 6797 3339
rect 6745 3223 6797 3275
rect 9923 3403 9975 3455
rect 9987 3403 10039 3455
rect 11899 3434 11951 3486
rect 11899 3370 11951 3422
rect 9793 3287 9845 3339
rect 9793 3223 9845 3275
rect 9923 3080 9975 3132
rect 9987 3080 10039 3132
rect 6745 2949 6797 3001
rect 6745 2885 6797 2937
rect 6484 2535 6536 2587
rect 6558 2535 6610 2587
rect 6632 2535 6684 2587
rect 6484 2467 6536 2519
rect 6558 2467 6610 2519
rect 6632 2467 6684 2519
rect 6484 2399 6536 2451
rect 6558 2399 6610 2451
rect 6632 2399 6684 2451
rect 5824 1885 5876 1937
rect 5888 1885 5940 1937
rect 553 1814 605 1866
rect 621 1814 673 1866
rect 688 1814 740 1866
rect 755 1814 807 1866
rect 822 1814 874 1866
rect 889 1814 941 1866
rect 6347 1004 6399 1056
rect 3157 952 3209 1004
rect 3221 952 3273 1004
rect 3713 952 3765 1004
rect 3777 952 3829 1004
rect 6347 940 6399 992
rect 6547 1004 6599 1056
rect 6547 940 6599 992
rect 1237 668 1289 720
rect 1301 668 1353 720
rect 3074 629 3126 681
rect 3138 629 3190 681
rect 3856 635 3908 687
rect 3920 635 3972 687
rect 5482 547 5534 599
rect 5546 547 5598 599
rect 5989 547 6041 599
rect 6053 547 6105 599
rect 553 427 605 479
rect 621 427 673 479
rect 688 427 740 479
rect 755 427 807 479
rect 822 427 874 479
rect 889 427 941 479
rect 553 349 605 401
rect 621 349 673 401
rect 688 349 740 401
rect 755 349 807 401
rect 822 349 874 401
rect 889 349 941 401
rect 979 70 1031 122
rect 979 6 1031 58
rect 1231 70 1283 122
rect 1231 6 1283 58
rect 6059 70 6111 122
rect 6059 6 6111 58
rect 6347 407 6399 459
rect 6347 343 6399 395
rect 6347 70 6399 122
rect 6347 6 6399 58
rect 6547 407 6599 459
rect 6547 343 6599 395
rect 6547 70 6599 122
rect 6547 6 6599 58
rect 8527 2818 8579 2870
rect 8527 2754 8579 2806
rect 6891 1082 6943 1134
rect 6956 1082 7008 1134
rect 7393 972 7445 1024
rect 7393 910 7445 928
rect 7393 876 7409 910
rect 7409 876 7445 910
rect 7835 876 7844 910
rect 7844 876 7878 910
rect 7878 876 7887 910
rect 7835 858 7887 876
rect 7909 876 7923 910
rect 7923 876 7957 910
rect 7957 876 7961 910
rect 7909 858 7961 876
rect 7983 858 8035 910
rect 7835 788 7887 803
rect 7835 754 7869 788
rect 7869 754 7887 788
rect 7835 751 7887 754
rect 7909 751 7961 803
rect 7983 798 7995 803
rect 7995 798 8029 803
rect 8029 798 8035 803
rect 7983 754 8035 798
rect 7983 751 7995 754
rect 7995 751 8029 754
rect 8029 751 8035 754
rect 7835 644 7887 696
rect 7909 644 7961 696
rect 7983 675 8035 696
rect 7983 644 7995 675
rect 7995 644 8029 675
rect 8029 644 8035 675
rect 7224 597 7233 601
rect 7233 597 7267 601
rect 7267 597 7276 601
rect 7224 549 7276 597
rect 7503 632 7555 641
rect 7503 598 7531 632
rect 7531 598 7555 632
rect 7503 589 7555 598
rect 7567 632 7619 641
rect 7567 598 7581 632
rect 7581 598 7615 632
rect 7615 598 7619 632
rect 7567 589 7619 598
rect 9482 1082 9534 1134
rect 9547 1082 9599 1134
rect 12642 7675 12694 7727
rect 12710 7675 12762 7727
rect 12778 7675 12830 7727
rect 12637 2909 12689 2961
rect 12709 2909 12761 2961
rect 12781 2909 12833 2961
rect 12637 2842 12689 2894
rect 12709 2842 12761 2894
rect 12781 2842 12833 2894
rect 12637 2774 12689 2826
rect 12709 2774 12761 2826
rect 12781 2774 12833 2826
rect 12642 1743 12694 1795
rect 12710 1743 12762 1795
rect 12778 1743 12830 1795
rect 12642 1671 12694 1723
rect 12710 1671 12762 1723
rect 12778 1671 12830 1723
rect 12642 1599 12694 1651
rect 12710 1599 12762 1651
rect 12778 1599 12830 1651
rect 15571 38827 15623 38879
rect 15571 38759 15623 38811
rect 15571 38691 15623 38743
rect 15571 36103 15623 36155
rect 15571 36035 15623 36087
rect 15571 35967 15623 36019
rect 15571 33995 15623 34047
rect 15571 33927 15623 33979
rect 15571 33859 15623 33911
rect 15571 31271 15623 31323
rect 15571 31203 15623 31255
rect 15571 31135 15623 31187
rect 15571 29163 15623 29215
rect 15571 29095 15623 29147
rect 15571 29027 15623 29079
rect 15571 26439 15623 26491
rect 15571 26371 15623 26423
rect 15571 26303 15623 26355
rect 15571 24331 15623 24383
rect 15571 24263 15623 24315
rect 15571 24195 15623 24247
rect 15571 21607 15623 21659
rect 15571 21539 15623 21591
rect 15571 21471 15623 21523
rect 15571 16775 15623 16827
rect 15571 16707 15623 16759
rect 15571 16639 15623 16691
rect 15571 14667 15623 14719
rect 15571 14599 15623 14651
rect 15571 14531 15623 14583
rect 15571 11943 15623 11995
rect 15571 11875 15623 11927
rect 15571 11807 15623 11859
rect 15571 9835 15623 9887
rect 15571 9767 15623 9819
rect 15571 9699 15623 9751
rect 9685 1160 9737 1212
rect 9685 1084 9737 1136
rect 9685 1008 9737 1060
rect 13307 1022 13359 1074
rect 13375 1022 13427 1074
rect 13442 1022 13494 1074
rect 13509 1022 13561 1074
rect 13576 1022 13628 1074
rect 13643 1022 13695 1074
rect 8613 918 8665 970
rect 8677 918 8729 970
rect 9923 952 9975 1004
rect 9987 952 10039 1004
rect 13307 936 13359 988
rect 13375 936 13427 988
rect 13442 936 13494 988
rect 13509 936 13561 988
rect 13576 936 13628 988
rect 13643 936 13695 988
rect 8207 705 8259 757
rect 8207 641 8259 693
rect 8859 863 8911 870
rect 8927 863 8979 870
rect 8859 829 8883 863
rect 8883 829 8911 863
rect 8927 829 8959 863
rect 8959 829 8979 863
rect 8859 818 8911 829
rect 8927 818 8979 829
rect 8994 863 9046 870
rect 8994 829 9001 863
rect 9001 829 9035 863
rect 9035 829 9046 863
rect 8994 818 9046 829
rect 9061 863 9113 870
rect 9061 829 9077 863
rect 9077 829 9111 863
rect 9111 829 9113 863
rect 9061 818 9113 829
rect 9128 863 9180 870
rect 9195 863 9247 870
rect 9262 863 9314 870
rect 9329 863 9381 870
rect 9396 863 9448 870
rect 9463 863 9515 870
rect 9128 829 9153 863
rect 9153 829 9180 863
rect 9195 829 9229 863
rect 9229 829 9247 863
rect 9262 829 9263 863
rect 9263 829 9305 863
rect 9305 829 9314 863
rect 9329 829 9339 863
rect 9339 829 9381 863
rect 9396 829 9415 863
rect 9415 829 9448 863
rect 9463 829 9491 863
rect 9491 829 9515 863
rect 9128 818 9180 829
rect 9195 818 9247 829
rect 9262 818 9314 829
rect 9329 818 9381 829
rect 9396 818 9448 829
rect 9463 818 9515 829
rect 9530 863 9582 870
rect 9530 829 9533 863
rect 9533 829 9567 863
rect 9567 829 9582 863
rect 9530 818 9582 829
rect 9597 863 9649 870
rect 9597 829 9609 863
rect 9609 829 9643 863
rect 9643 829 9649 863
rect 9597 818 9649 829
rect 13307 850 13359 902
rect 13375 850 13427 902
rect 13442 850 13494 902
rect 13509 850 13561 902
rect 13576 850 13628 902
rect 13643 850 13695 902
rect 8859 785 8911 806
rect 8927 785 8979 806
rect 8859 754 8883 785
rect 8883 754 8911 785
rect 8927 754 8959 785
rect 8959 754 8979 785
rect 8994 785 9046 806
rect 8994 754 9001 785
rect 9001 754 9035 785
rect 9035 754 9046 785
rect 9061 785 9113 806
rect 9061 754 9077 785
rect 9077 754 9111 785
rect 9111 754 9113 785
rect 9128 785 9180 806
rect 9195 785 9247 806
rect 9262 785 9314 806
rect 9329 785 9381 806
rect 9396 785 9448 806
rect 9463 785 9515 806
rect 9128 754 9153 785
rect 9153 754 9180 785
rect 9195 754 9229 785
rect 9229 754 9247 785
rect 9262 754 9263 785
rect 9263 754 9305 785
rect 9305 754 9314 785
rect 9329 754 9339 785
rect 9339 754 9381 785
rect 9396 754 9415 785
rect 9415 754 9448 785
rect 9463 754 9491 785
rect 9491 754 9515 785
rect 9530 785 9582 806
rect 9530 754 9533 785
rect 9533 754 9567 785
rect 9567 754 9582 785
rect 9597 785 9649 806
rect 9597 754 9609 785
rect 9609 754 9643 785
rect 9643 754 9649 785
rect 7224 505 7233 537
rect 7233 505 7267 537
rect 7267 505 7276 537
rect 7835 536 7887 588
rect 7909 536 7961 588
rect 7983 562 7995 588
rect 7995 562 8029 588
rect 8029 562 8035 588
rect 7983 536 8035 562
rect 7224 485 7276 505
rect 7835 476 7887 480
rect 7835 442 7869 476
rect 7869 442 7887 476
rect 7835 428 7887 442
rect 7909 428 7961 480
rect 7983 428 8035 480
rect 7835 354 7887 372
rect 7835 320 7844 354
rect 7844 320 7878 354
rect 7878 320 7887 354
rect 7909 354 7961 372
rect 7909 320 7923 354
rect 7923 320 7957 354
rect 7957 320 7961 354
rect 7983 320 8035 372
rect 9923 635 9975 687
rect 9987 635 10039 687
rect 8339 268 8391 320
rect 8407 268 8459 320
rect 8474 268 8526 320
rect 8541 268 8593 320
rect 8608 268 8660 320
rect 8675 268 8727 320
rect 6880 161 6932 213
rect 6944 161 6996 213
rect 8044 161 8096 213
rect 8108 161 8160 213
rect 8339 194 8391 246
rect 8407 194 8459 246
rect 8474 194 8526 246
rect 8541 194 8593 246
rect 8608 194 8660 246
rect 8675 194 8727 246
rect 6745 70 6797 122
rect 6745 6 6797 58
rect 7503 76 7555 128
rect 7567 76 7619 128
rect 8339 120 8391 172
rect 8407 120 8459 172
rect 8474 120 8526 172
rect 8541 120 8593 172
rect 8608 120 8660 172
rect 8675 120 8727 172
rect 12327 240 12379 292
rect 12403 240 12455 292
rect 12479 240 12531 292
rect 12555 240 12607 292
rect 12631 240 12683 292
rect 12706 240 12758 292
rect 7503 0 7555 52
rect 7567 0 7619 52
rect 12099 70 12151 122
rect 12099 6 12151 58
rect 13080 70 13132 122
rect 13080 6 13132 58
<< metal2 >>
rect 8333 39085 8342 39141
rect 8398 39085 8424 39141
rect 8480 39085 8506 39141
rect 8562 39085 8587 39141
rect 8643 39085 8668 39141
rect 8724 39085 8733 39141
rect 8333 38997 8733 39085
rect 8333 38941 8342 38997
rect 8398 38941 8424 38997
rect 8480 38941 8506 38997
rect 8562 38941 8587 38997
rect 8643 38941 8668 38997
rect 8724 38941 8733 38997
rect 385 38879 7020 38885
rect 437 38827 2464 38879
rect 2516 38827 4606 38879
rect 4658 38827 6745 38879
rect 6797 38827 7020 38879
rect 385 38811 7020 38827
rect 437 38759 2464 38811
rect 2516 38759 4606 38811
rect 4658 38759 6745 38811
rect 6797 38759 7020 38811
rect 385 38743 7020 38759
rect 437 38691 2464 38743
rect 2516 38691 4606 38743
rect 4658 38691 6745 38743
rect 6797 38691 7020 38743
rect 385 38685 7020 38691
rect 7813 38829 7822 38885
rect 7878 38829 7904 38885
rect 7960 38829 7986 38885
rect 8042 38829 8067 38885
rect 8123 38829 8148 38885
rect 8204 38829 8213 38885
rect 7813 38741 8213 38829
rect 7813 38685 7822 38741
rect 7878 38685 7904 38741
rect 7960 38685 7986 38741
rect 8042 38685 8067 38741
rect 8123 38685 8148 38741
rect 8204 38685 8213 38741
rect 9525 38879 15623 38885
rect 9525 38827 9633 38879
rect 9685 38827 9725 38879
rect 9777 38827 10860 38879
rect 10912 38827 12058 38879
rect 12110 38827 13846 38879
rect 13898 38827 15571 38879
rect 9525 38811 15623 38827
rect 9525 38759 9633 38811
rect 9685 38759 9725 38811
rect 9777 38759 10860 38811
rect 10912 38759 12058 38811
rect 12110 38759 13846 38811
rect 13898 38759 15571 38811
rect 9525 38743 15623 38759
rect 9525 38691 9633 38743
rect 9685 38691 9725 38743
rect 9777 38691 10860 38743
rect 10912 38691 12058 38743
rect 12110 38691 13846 38743
rect 13898 38691 15571 38743
rect 9525 38685 15623 38691
rect 4910 38432 7890 38438
rect 4962 38431 7890 38432
tri 7890 38431 7897 38438 sw
rect 4962 38386 7897 38431
rect 4962 38380 4967 38386
rect 4910 38368 4967 38380
rect 4962 38357 4967 38368
tri 4967 38357 4996 38386 nw
tri 7868 38357 7897 38386 ne
tri 7897 38357 7971 38431 sw
tri 4962 38352 4967 38357 nw
tri 7897 38352 7902 38357 ne
rect 7902 38352 7971 38357
rect 4910 38310 4962 38316
tri 7902 38310 7944 38352 ne
rect 7944 38310 7971 38352
tri 7944 38283 7971 38310 ne
tri 7971 38283 8045 38357 sw
tri 7971 38209 8045 38283 ne
tri 8045 38209 8119 38283 sw
tri 8045 38135 8119 38209 ne
tri 8119 38135 8193 38209 sw
tri 8119 38061 8193 38135 ne
tri 8193 38061 8267 38135 sw
rect 626 38055 7245 38061
rect 678 38009 7245 38055
tri 8193 38009 8245 38061 ne
rect 8245 38009 8785 38061
rect 626 37991 678 38003
tri 678 37975 712 38009 nw
tri 7210 37975 7244 38009 ne
tri 8751 37975 8785 38009 ne
rect 626 37933 678 37939
tri 7210 37093 7244 37127 se
tri 8751 37093 8785 37127 se
rect 862 37087 7245 37093
rect 914 37041 7245 37087
tri 8193 37041 8245 37093 se
rect 8245 37041 8785 37093
rect 914 37035 926 37041
rect 862 37023 926 37035
rect 914 37019 926 37023
tri 926 37019 948 37041 nw
tri 8171 37019 8193 37041 se
rect 8193 37019 8245 37041
tri 8245 37019 8267 37041 nw
tri 914 37007 926 37019 nw
tri 8159 37007 8171 37019 se
rect 862 36965 914 36971
tri 8117 36965 8159 37007 se
rect 8159 36965 8171 37007
tri 8097 36945 8117 36965 se
rect 8117 36945 8171 36965
tri 8171 36945 8245 37019 nw
tri 8023 36871 8097 36945 se
tri 8097 36871 8171 36945 nw
tri 7949 36797 8023 36871 se
tri 8023 36797 8097 36871 nw
tri 7875 36723 7949 36797 se
tri 7949 36723 8023 36797 nw
tri 7868 36716 7875 36723 se
rect 7875 36716 7942 36723
tri 7942 36716 7949 36723 nw
rect 5146 36710 7890 36716
rect 5198 36664 7890 36710
tri 7890 36664 7942 36716 nw
rect 5146 36646 5198 36658
tri 5198 36630 5232 36664 nw
rect 5146 36588 5198 36594
rect 8333 36361 8342 36417
rect 8398 36361 8424 36417
rect 8480 36361 8506 36417
rect 8562 36361 8587 36417
rect 8643 36361 8668 36417
rect 8724 36361 8733 36417
rect 8333 36273 8733 36361
rect 8333 36217 8342 36273
rect 8398 36217 8424 36273
rect 8480 36217 8506 36273
rect 8562 36217 8587 36273
rect 8643 36217 8668 36273
rect 8724 36217 8733 36273
rect 385 36155 7026 36161
rect 437 36103 2464 36155
rect 2516 36103 4606 36155
rect 4658 36103 6745 36155
rect 6797 36103 7026 36155
rect 385 36087 7026 36103
rect 437 36035 2464 36087
rect 2516 36035 4606 36087
rect 4658 36035 6745 36087
rect 6797 36035 7026 36087
rect 385 36019 7026 36035
rect 437 35967 2464 36019
rect 2516 35967 4606 36019
rect 4658 35967 6745 36019
rect 6797 35967 7026 36019
rect 385 35961 7026 35967
rect 7813 36105 7822 36161
rect 7878 36105 7904 36161
rect 7960 36105 7986 36161
rect 8042 36105 8067 36161
rect 8123 36105 8148 36161
rect 8204 36105 8213 36161
rect 7813 36017 8213 36105
rect 7813 35961 7822 36017
rect 7878 35961 7904 36017
rect 7960 35961 7986 36017
rect 8042 35961 8067 36017
rect 8123 35961 8148 36017
rect 8204 35961 8213 36017
rect 9498 36155 15623 36161
rect 9498 36103 9633 36155
rect 9685 36103 9725 36155
rect 9777 36103 10860 36155
rect 10912 36103 12058 36155
rect 12110 36103 13846 36155
rect 13898 36103 15571 36155
rect 9498 36087 15623 36103
rect 9498 36035 9633 36087
rect 9685 36035 9725 36087
rect 9777 36035 10860 36087
rect 10912 36035 12058 36087
rect 12110 36035 13846 36087
rect 13898 36035 15571 36087
rect 9498 36019 15623 36035
rect 9498 35967 9633 36019
rect 9685 35967 9725 36019
rect 9777 35967 10860 36019
rect 10912 35967 12058 36019
rect 12110 35967 13846 36019
rect 13898 35967 15571 36019
rect 9498 35961 15623 35967
rect 8333 34253 8342 34309
rect 8398 34253 8424 34309
rect 8480 34253 8506 34309
rect 8562 34253 8587 34309
rect 8643 34253 8668 34309
rect 8724 34253 8733 34309
rect 8333 34165 8733 34253
rect 8333 34109 8342 34165
rect 8398 34109 8424 34165
rect 8480 34109 8506 34165
rect 8562 34109 8587 34165
rect 8643 34109 8668 34165
rect 8724 34109 8733 34165
rect 385 34047 7026 34053
rect 437 33995 2464 34047
rect 2516 33995 4606 34047
rect 4658 33995 6745 34047
rect 6797 33995 7026 34047
rect 385 33979 7026 33995
rect 437 33927 2464 33979
rect 2516 33927 4606 33979
rect 4658 33927 6745 33979
rect 6797 33927 7026 33979
rect 385 33911 7026 33927
rect 437 33859 2464 33911
rect 2516 33859 4606 33911
rect 4658 33859 6745 33911
rect 6797 33859 7026 33911
rect 385 33853 7026 33859
rect 7813 33997 7822 34053
rect 7878 33997 7904 34053
rect 7960 33997 7986 34053
rect 8042 33997 8067 34053
rect 8123 33997 8148 34053
rect 8204 33997 8213 34053
rect 7813 33909 8213 33997
rect 7813 33853 7822 33909
rect 7878 33853 7904 33909
rect 7960 33853 7986 33909
rect 8042 33853 8067 33909
rect 8123 33853 8148 33909
rect 8204 33853 8213 33909
rect 9498 34047 15623 34053
rect 9498 33995 9633 34047
rect 9685 33995 9725 34047
rect 9777 33995 10860 34047
rect 10912 33995 12058 34047
rect 12110 33995 13846 34047
rect 13898 33995 15571 34047
rect 9498 33979 15623 33995
rect 9498 33927 9633 33979
rect 9685 33927 9725 33979
rect 9777 33927 10860 33979
rect 10912 33927 12058 33979
rect 12110 33927 13846 33979
rect 13898 33927 15571 33979
rect 9498 33911 15623 33927
rect 9498 33859 9633 33911
rect 9685 33859 9725 33911
rect 9777 33859 10860 33911
rect 10912 33859 12058 33911
rect 12110 33859 13846 33911
rect 13898 33859 15571 33911
rect 9498 33853 15623 33859
rect 5382 33600 7890 33606
rect 5434 33599 7890 33600
tri 7890 33599 7897 33606 sw
rect 5434 33554 7897 33599
rect 5434 33548 5439 33554
rect 5382 33536 5439 33548
rect 5434 33525 5439 33536
tri 5439 33525 5468 33554 nw
tri 7868 33525 7897 33554 ne
tri 7897 33525 7971 33599 sw
tri 5434 33520 5439 33525 nw
tri 7897 33520 7902 33525 ne
rect 7902 33520 7971 33525
rect 5382 33478 5434 33484
tri 7902 33478 7944 33520 ne
rect 7944 33478 7971 33520
tri 7944 33451 7971 33478 ne
tri 7971 33451 8045 33525 sw
tri 7971 33377 8045 33451 ne
tri 8045 33377 8119 33451 sw
tri 8045 33303 8119 33377 ne
tri 8119 33303 8193 33377 sw
tri 8119 33229 8193 33303 ne
tri 8193 33229 8267 33303 sw
rect 1098 33223 7245 33229
rect 1150 33177 7245 33223
tri 8193 33177 8245 33229 ne
rect 8245 33177 8785 33229
rect 1098 33159 1150 33171
tri 1150 33143 1184 33177 nw
tri 7210 33143 7244 33177 ne
tri 8751 33143 8785 33177 ne
rect 1098 33101 1150 33107
tri 7210 32261 7244 32295 se
tri 8751 32261 8785 32295 se
rect 1337 32255 7245 32261
rect 1389 32209 7245 32255
tri 8193 32209 8245 32261 se
rect 8245 32209 8785 32261
rect 1389 32203 1401 32209
rect 1337 32191 1401 32203
rect 1389 32187 1401 32191
tri 1401 32187 1423 32209 nw
tri 8171 32187 8193 32209 se
rect 8193 32187 8245 32209
tri 8245 32187 8267 32209 nw
tri 1389 32175 1401 32187 nw
tri 8159 32175 8171 32187 se
rect 1337 32133 1389 32139
tri 8117 32133 8159 32175 se
rect 8159 32133 8171 32175
tri 8097 32113 8117 32133 se
rect 8117 32113 8171 32133
tri 8171 32113 8245 32187 nw
tri 8023 32039 8097 32113 se
tri 8097 32039 8171 32113 nw
tri 7949 31965 8023 32039 se
tri 8023 31965 8097 32039 nw
tri 7875 31891 7949 31965 se
tri 7949 31891 8023 31965 nw
tri 7868 31884 7875 31891 se
rect 7875 31884 7942 31891
tri 7942 31884 7949 31891 nw
rect 5618 31878 7890 31884
rect 5670 31832 7890 31878
tri 7890 31832 7942 31884 nw
rect 5618 31814 5670 31826
tri 5670 31798 5704 31832 nw
rect 5618 31756 5670 31762
rect 8333 31529 8342 31585
rect 8398 31529 8424 31585
rect 8480 31529 8506 31585
rect 8562 31529 8587 31585
rect 8643 31529 8668 31585
rect 8724 31529 8733 31585
rect 8333 31441 8733 31529
rect 8333 31385 8342 31441
rect 8398 31385 8424 31441
rect 8480 31385 8506 31441
rect 8562 31385 8587 31441
rect 8643 31385 8668 31441
rect 8724 31385 8733 31441
rect 385 31323 7026 31329
rect 437 31271 2464 31323
rect 2516 31271 4606 31323
rect 4658 31271 6745 31323
rect 6797 31271 7026 31323
rect 385 31255 7026 31271
rect 437 31203 2464 31255
rect 2516 31203 4606 31255
rect 4658 31203 6745 31255
rect 6797 31203 7026 31255
rect 385 31187 7026 31203
rect 437 31135 2464 31187
rect 2516 31135 4606 31187
rect 4658 31135 6745 31187
rect 6797 31135 7026 31187
rect 385 31129 7026 31135
rect 7813 31273 7822 31329
rect 7878 31273 7904 31329
rect 7960 31273 7986 31329
rect 8042 31273 8067 31329
rect 8123 31273 8148 31329
rect 8204 31273 8213 31329
rect 7813 31185 8213 31273
rect 7813 31129 7822 31185
rect 7878 31129 7904 31185
rect 7960 31129 7986 31185
rect 8042 31129 8067 31185
rect 8123 31129 8148 31185
rect 8204 31129 8213 31185
rect 9498 31323 15623 31329
rect 9498 31271 9633 31323
rect 9685 31271 9725 31323
rect 9777 31271 10860 31323
rect 10912 31271 12058 31323
rect 12110 31271 13846 31323
rect 13898 31271 15571 31323
rect 9498 31255 15623 31271
rect 9498 31203 9633 31255
rect 9685 31203 9725 31255
rect 9777 31203 10860 31255
rect 10912 31203 12058 31255
rect 12110 31203 13846 31255
rect 13898 31203 15571 31255
rect 9498 31187 15623 31203
rect 9498 31135 9633 31187
rect 9685 31135 9725 31187
rect 9777 31135 10860 31187
rect 10912 31135 12058 31187
rect 12110 31135 13846 31187
rect 13898 31135 15571 31187
rect 9498 31129 15623 31135
rect 8333 29421 8342 29477
rect 8398 29421 8424 29477
rect 8480 29421 8506 29477
rect 8562 29421 8587 29477
rect 8643 29421 8668 29477
rect 8724 29421 8733 29477
rect 8333 29333 8733 29421
rect 8333 29277 8342 29333
rect 8398 29277 8424 29333
rect 8480 29277 8506 29333
rect 8562 29277 8587 29333
rect 8643 29277 8668 29333
rect 8724 29277 8733 29333
rect 385 29215 7020 29221
rect 437 29163 2464 29215
rect 2516 29163 4606 29215
rect 4658 29163 6745 29215
rect 6797 29163 7020 29215
rect 385 29147 7020 29163
rect 437 29095 2464 29147
rect 2516 29095 4606 29147
rect 4658 29095 6745 29147
rect 6797 29095 7020 29147
rect 385 29079 7020 29095
rect 437 29027 2464 29079
rect 2516 29027 4606 29079
rect 4658 29027 6745 29079
rect 6797 29027 7020 29079
rect 385 29021 7020 29027
rect 7813 29165 7822 29221
rect 7878 29165 7904 29221
rect 7960 29165 7986 29221
rect 8042 29165 8067 29221
rect 8123 29165 8148 29221
rect 8204 29165 8213 29221
rect 7813 29077 8213 29165
rect 7813 29021 7822 29077
rect 7878 29021 7904 29077
rect 7960 29021 7986 29077
rect 8042 29021 8067 29077
rect 8123 29021 8148 29077
rect 8204 29021 8213 29077
rect 9525 29215 15623 29221
rect 9525 29163 9633 29215
rect 9685 29163 9725 29215
rect 9777 29163 10860 29215
rect 10912 29163 12058 29215
rect 12110 29163 13846 29215
rect 13898 29163 15571 29215
rect 9525 29147 15623 29163
rect 9525 29095 9633 29147
rect 9685 29095 9725 29147
rect 9777 29095 10860 29147
rect 10912 29095 12058 29147
rect 12110 29095 13846 29147
rect 13898 29095 15571 29147
rect 9525 29079 15623 29095
rect 9525 29027 9633 29079
rect 9685 29027 9725 29079
rect 9777 29027 10860 29079
rect 10912 29027 12058 29079
rect 12110 29027 13846 29079
rect 13898 29027 15571 29079
rect 9525 29021 15623 29027
rect 5854 28768 7890 28774
rect 5906 28767 7890 28768
tri 7890 28767 7897 28774 sw
rect 5906 28722 7897 28767
rect 5906 28716 5911 28722
rect 5854 28704 5911 28716
rect 5906 28693 5911 28704
tri 5911 28693 5940 28722 nw
tri 7868 28693 7897 28722 ne
tri 7897 28693 7971 28767 sw
tri 5906 28688 5911 28693 nw
tri 7897 28688 7902 28693 ne
rect 7902 28688 7971 28693
rect 5854 28646 5906 28652
tri 7902 28646 7944 28688 ne
rect 7944 28646 7971 28688
tri 7944 28619 7971 28646 ne
tri 7971 28619 8045 28693 sw
tri 7971 28545 8045 28619 ne
tri 8045 28545 8119 28619 sw
tri 8045 28471 8119 28545 ne
tri 8119 28471 8193 28545 sw
tri 8119 28397 8193 28471 ne
tri 8193 28397 8267 28471 sw
rect 1573 28391 7245 28397
rect 1625 28345 7245 28391
tri 8193 28345 8245 28397 ne
rect 8245 28345 8785 28397
rect 1573 28327 1625 28339
tri 1625 28311 1659 28345 nw
tri 7210 28311 7244 28345 ne
tri 8751 28311 8785 28345 ne
rect 1573 28269 1625 28275
tri 7210 27429 7244 27463 se
tri 8751 27429 8785 27463 se
rect 1809 27423 7245 27429
rect 1861 27377 7245 27423
tri 8193 27377 8245 27429 se
rect 8245 27377 8785 27429
rect 1861 27371 1873 27377
rect 1809 27359 1873 27371
rect 1861 27355 1873 27359
tri 1873 27355 1895 27377 nw
tri 8171 27355 8193 27377 se
rect 8193 27355 8245 27377
tri 8245 27355 8267 27377 nw
tri 1861 27343 1873 27355 nw
tri 8159 27343 8171 27355 se
rect 1809 27301 1861 27307
tri 8117 27301 8159 27343 se
rect 8159 27301 8171 27343
tri 8097 27281 8117 27301 se
rect 8117 27281 8171 27301
tri 8171 27281 8245 27355 nw
tri 8023 27207 8097 27281 se
tri 8097 27207 8171 27281 nw
tri 7949 27133 8023 27207 se
tri 8023 27133 8097 27207 nw
tri 7875 27059 7949 27133 se
tri 7949 27059 8023 27133 nw
tri 7868 27052 7875 27059 se
rect 7875 27052 7942 27059
tri 7942 27052 7949 27059 nw
rect 6090 27046 7890 27052
rect 6142 27000 7890 27046
tri 7890 27000 7942 27052 nw
rect 6090 26982 6142 26994
tri 6142 26966 6176 27000 nw
rect 6090 26924 6142 26930
rect 8333 26697 8342 26753
rect 8398 26697 8424 26753
rect 8480 26697 8506 26753
rect 8562 26697 8587 26753
rect 8643 26697 8668 26753
rect 8724 26697 8733 26753
rect 8333 26609 8733 26697
rect 8333 26553 8342 26609
rect 8398 26553 8424 26609
rect 8480 26553 8506 26609
rect 8562 26553 8587 26609
rect 8643 26553 8668 26609
rect 8724 26553 8733 26609
rect 385 26491 7026 26497
rect 437 26439 2464 26491
rect 2516 26439 4606 26491
rect 4658 26439 6745 26491
rect 6797 26439 7026 26491
rect 385 26423 7026 26439
rect 437 26371 2464 26423
rect 2516 26371 4606 26423
rect 4658 26371 6745 26423
rect 6797 26371 7026 26423
rect 385 26355 7026 26371
rect 437 26303 2464 26355
rect 2516 26303 4606 26355
rect 4658 26303 6745 26355
rect 6797 26303 7026 26355
rect 385 26297 7026 26303
rect 7813 26441 7822 26497
rect 7878 26441 7904 26497
rect 7960 26441 7986 26497
rect 8042 26441 8067 26497
rect 8123 26441 8148 26497
rect 8204 26441 8213 26497
rect 7813 26353 8213 26441
rect 7813 26297 7822 26353
rect 7878 26297 7904 26353
rect 7960 26297 7986 26353
rect 8042 26297 8067 26353
rect 8123 26297 8148 26353
rect 8204 26297 8213 26353
rect 9498 26491 15623 26497
rect 9498 26439 9633 26491
rect 9685 26439 9725 26491
rect 9777 26439 10860 26491
rect 10912 26439 12058 26491
rect 12110 26439 13846 26491
rect 13898 26439 15571 26491
rect 9498 26423 15623 26439
rect 9498 26371 9633 26423
rect 9685 26371 9725 26423
rect 9777 26371 10860 26423
rect 10912 26371 12058 26423
rect 12110 26371 13846 26423
rect 13898 26371 15571 26423
rect 9498 26355 15623 26371
rect 9498 26303 9633 26355
rect 9685 26303 9725 26355
rect 9777 26303 10860 26355
rect 10912 26303 12058 26355
rect 12110 26303 13846 26355
rect 13898 26303 15571 26355
rect 9498 26297 15623 26303
rect 8333 24589 8342 24645
rect 8398 24589 8424 24645
rect 8480 24589 8506 24645
rect 8562 24589 8587 24645
rect 8643 24589 8668 24645
rect 8724 24589 8733 24645
rect 8333 24501 8733 24589
rect 8333 24445 8342 24501
rect 8398 24445 8424 24501
rect 8480 24445 8506 24501
rect 8562 24445 8587 24501
rect 8643 24445 8668 24501
rect 8724 24445 8733 24501
rect 385 24383 7026 24389
rect 437 24331 2464 24383
rect 2516 24331 4606 24383
rect 4658 24331 6745 24383
rect 6797 24331 7026 24383
rect 385 24315 7026 24331
rect 437 24263 2464 24315
rect 2516 24263 4606 24315
rect 4658 24263 6745 24315
rect 6797 24263 7026 24315
rect 385 24247 7026 24263
rect 437 24195 2464 24247
rect 2516 24195 4606 24247
rect 4658 24195 6745 24247
rect 6797 24195 7026 24247
rect 385 24189 7026 24195
rect 7813 24333 7822 24389
rect 7878 24333 7904 24389
rect 7960 24333 7986 24389
rect 8042 24333 8067 24389
rect 8123 24333 8148 24389
rect 8204 24333 8213 24389
rect 7813 24245 8213 24333
rect 7813 24189 7822 24245
rect 7878 24189 7904 24245
rect 7960 24189 7986 24245
rect 8042 24189 8067 24245
rect 8123 24189 8148 24245
rect 8204 24189 8213 24245
rect 9498 24383 15623 24389
rect 9498 24331 9633 24383
rect 9685 24331 9725 24383
rect 9777 24331 10860 24383
rect 10912 24331 12058 24383
rect 12110 24331 13846 24383
rect 13898 24331 15571 24383
rect 9498 24315 15623 24331
rect 9498 24263 9633 24315
rect 9685 24263 9725 24315
rect 9777 24263 10860 24315
rect 10912 24263 12058 24315
rect 12110 24263 13846 24315
rect 13898 24263 15571 24315
rect 9498 24247 15623 24263
rect 9498 24195 9633 24247
rect 9685 24195 9725 24247
rect 9777 24195 10860 24247
rect 10912 24195 12058 24247
rect 12110 24195 13846 24247
rect 13898 24195 15571 24247
rect 9498 24189 15623 24195
rect 6326 24012 6378 24018
rect 6326 23948 6378 23960
tri 6378 23942 6412 23976 sw
rect 6378 23935 7890 23942
tri 7890 23935 7897 23942 sw
rect 6378 23896 7897 23935
rect 6326 23890 7897 23896
tri 7868 23861 7897 23890 ne
tri 7897 23861 7971 23935 sw
tri 7897 23787 7971 23861 ne
tri 7971 23787 8045 23861 sw
tri 7971 23713 8045 23787 ne
tri 8045 23713 8119 23787 sw
tri 8045 23639 8119 23713 ne
tri 8119 23639 8193 23713 sw
tri 8119 23565 8193 23639 ne
tri 8193 23565 8267 23639 sw
rect 2045 23559 7245 23565
rect 2097 23513 7245 23559
tri 8193 23513 8245 23565 ne
rect 8245 23513 8785 23565
rect 2045 23495 2097 23507
tri 2097 23479 2131 23513 nw
tri 7210 23479 7244 23513 ne
tri 8751 23479 8785 23513 ne
rect 2045 23437 2097 23443
tri 7210 22597 7244 22631 se
tri 8751 22597 8785 22631 se
rect 2278 22591 7245 22597
rect 2330 22545 7245 22591
tri 8193 22545 8245 22597 se
rect 8245 22545 8785 22597
rect 2330 22539 2342 22545
rect 2278 22527 2342 22539
rect 2330 22523 2342 22527
tri 2342 22523 2364 22545 nw
tri 8171 22523 8193 22545 se
rect 8193 22523 8245 22545
tri 8245 22523 8267 22545 nw
tri 2330 22511 2342 22523 nw
tri 8159 22511 8171 22523 se
rect 2278 22469 2330 22475
tri 8117 22469 8159 22511 se
rect 8159 22469 8171 22511
tri 8097 22449 8117 22469 se
rect 8117 22449 8171 22469
tri 8171 22449 8245 22523 nw
tri 8023 22375 8097 22449 se
tri 8097 22375 8171 22449 nw
tri 7949 22301 8023 22375 se
tri 8023 22301 8097 22375 nw
tri 7875 22227 7949 22301 se
tri 7949 22227 8023 22301 nw
tri 7868 22220 7875 22227 se
rect 7875 22220 7942 22227
tri 7942 22220 7949 22227 nw
rect 6562 22214 7890 22220
rect 6614 22168 7890 22214
tri 7890 22168 7942 22220 nw
rect 6562 22150 6614 22162
tri 6614 22134 6648 22168 nw
rect 6562 22092 6614 22098
rect 8333 21865 8342 21921
rect 8398 21865 8424 21921
rect 8480 21865 8506 21921
rect 8562 21865 8587 21921
rect 8643 21865 8668 21921
rect 8724 21865 8733 21921
rect 8333 21777 8733 21865
rect 8333 21721 8342 21777
rect 8398 21721 8424 21777
rect 8480 21721 8506 21777
rect 8562 21721 8587 21777
rect 8643 21721 8668 21777
rect 8724 21721 8733 21777
rect 385 21659 7026 21665
rect 437 21607 2464 21659
rect 2516 21607 4606 21659
rect 4658 21607 6745 21659
rect 6797 21607 7026 21659
rect 385 21591 7026 21607
rect 437 21539 2464 21591
rect 2516 21539 4606 21591
rect 4658 21539 6745 21591
rect 6797 21539 7026 21591
rect 385 21523 7026 21539
rect 437 21471 2464 21523
rect 2516 21471 4606 21523
rect 4658 21471 6745 21523
rect 6797 21471 7026 21523
rect 385 21465 7026 21471
rect 7813 21609 7822 21665
rect 7878 21609 7904 21665
rect 7960 21609 7986 21665
rect 8042 21609 8067 21665
rect 8123 21609 8148 21665
rect 8204 21609 8213 21665
rect 7813 21521 8213 21609
rect 7813 21465 7822 21521
rect 7878 21465 7904 21521
rect 7960 21465 7986 21521
rect 8042 21465 8067 21521
rect 8123 21465 8148 21521
rect 8204 21465 8213 21521
rect 9498 21659 15623 21665
rect 9498 21607 9633 21659
rect 9685 21607 9725 21659
rect 9777 21607 10860 21659
rect 10912 21607 12058 21659
rect 12110 21607 13846 21659
rect 13898 21607 15571 21659
rect 9498 21591 15623 21607
rect 9498 21539 9633 21591
rect 9685 21539 9725 21591
rect 9777 21539 10860 21591
rect 10912 21539 12058 21591
rect 12110 21539 13846 21591
rect 13898 21539 15571 21591
rect 9498 21523 15623 21539
rect 9498 21471 9633 21523
rect 9685 21471 9725 21523
rect 9777 21471 10860 21523
rect 10912 21471 12058 21523
rect 12110 21471 13846 21523
rect 13898 21471 15571 21523
rect 9498 21465 15623 21471
rect 8333 19757 8342 19813
rect 8398 19757 8424 19813
rect 8480 19757 8506 19813
rect 8562 19757 8587 19813
rect 8643 19757 8668 19813
rect 8724 19757 8733 19813
rect 8333 19669 8733 19757
rect 8333 19613 8342 19669
rect 8398 19613 8424 19669
rect 8480 19613 8506 19669
rect 8562 19613 8587 19669
rect 8643 19613 8668 19669
rect 8724 19613 8733 19669
rect 385 19551 7026 19557
rect 437 19499 2464 19551
rect 2516 19499 4606 19551
rect 4658 19499 6745 19551
rect 6797 19499 7026 19551
rect 385 19483 7026 19499
rect 437 19431 2464 19483
rect 2516 19431 4606 19483
rect 4658 19431 6745 19483
rect 6797 19431 7026 19483
rect 385 19415 7026 19431
rect 437 19363 2464 19415
rect 2516 19363 4606 19415
rect 4658 19363 6745 19415
rect 6797 19363 7026 19415
rect 385 19357 7026 19363
rect 7813 19501 7822 19557
rect 7878 19501 7904 19557
rect 7960 19501 7986 19557
rect 8042 19501 8067 19557
rect 8123 19501 8148 19557
rect 8204 19501 8213 19557
rect 7813 19413 8213 19501
rect 7813 19357 7822 19413
rect 7878 19357 7904 19413
rect 7960 19357 7986 19413
rect 8042 19357 8067 19413
rect 8123 19357 8148 19413
rect 8204 19357 8213 19413
rect 2771 18727 7245 18733
rect 2823 18681 7245 18727
rect 9294 18727 10018 18733
rect 9294 18681 9966 18727
rect 2823 18675 2851 18681
tri 2851 18675 2857 18681 nw
tri 7210 18675 7216 18681 ne
rect 7216 18675 7244 18681
rect 2771 18663 2839 18675
tri 2839 18663 2851 18675 nw
tri 7216 18663 7228 18675 ne
rect 7228 18663 7244 18675
tri 2823 18647 2839 18663 nw
tri 7228 18647 7244 18663 ne
rect 9302 18675 9330 18681
tri 9330 18675 9336 18681 nw
tri 9932 18675 9938 18681 ne
rect 9938 18675 9966 18681
rect 9302 18663 9318 18675
tri 9318 18663 9330 18675 nw
tri 9938 18663 9950 18675 ne
rect 9950 18663 10018 18675
tri 9302 18647 9318 18663 nw
tri 9950 18647 9966 18663 ne
rect 2771 18605 2823 18611
rect 9966 18605 10018 18611
tri 7210 17765 7244 17799 se
tri 9302 17765 9336 17799 sw
rect 3007 17759 7245 17765
rect 3059 17713 7245 17759
rect 9271 17759 10254 17765
rect 9271 17713 10202 17759
rect 3059 17707 3087 17713
tri 3087 17707 3093 17713 nw
tri 10168 17707 10174 17713 ne
rect 10174 17707 10202 17713
rect 3007 17695 3075 17707
tri 3075 17695 3087 17707 nw
tri 10174 17695 10186 17707 ne
rect 10186 17695 10254 17707
tri 3059 17679 3075 17695 nw
tri 10186 17679 10202 17695 ne
rect 3007 17637 3059 17643
rect 10202 17637 10254 17643
rect 8333 17033 8342 17089
rect 8398 17033 8424 17089
rect 8480 17033 8506 17089
rect 8562 17033 8587 17089
rect 8643 17033 8668 17089
rect 8724 17033 8733 17089
rect 8333 16945 8733 17033
rect 8333 16889 8342 16945
rect 8398 16889 8424 16945
rect 8480 16889 8506 16945
rect 8562 16889 8587 16945
rect 8643 16889 8668 16945
rect 8724 16889 8733 16945
rect 385 16827 7027 16833
rect 437 16775 2464 16827
rect 2516 16775 4606 16827
rect 4658 16775 6745 16827
rect 6797 16775 7027 16827
rect 385 16759 7027 16775
rect 437 16707 2464 16759
rect 2516 16707 4606 16759
rect 4658 16707 6745 16759
rect 6797 16707 7027 16759
rect 385 16691 7027 16707
rect 437 16639 2464 16691
rect 2516 16639 4606 16691
rect 4658 16639 6745 16691
rect 6797 16639 7027 16691
rect 385 16633 7027 16639
rect 7813 16777 7822 16833
rect 7878 16777 7904 16833
rect 7960 16777 7986 16833
rect 8042 16777 8067 16833
rect 8123 16777 8148 16833
rect 8204 16777 8213 16833
rect 7813 16689 8213 16777
rect 7813 16633 7822 16689
rect 7878 16633 7904 16689
rect 7960 16633 7986 16689
rect 8042 16633 8067 16689
rect 8123 16633 8148 16689
rect 8204 16633 8213 16689
rect 9525 16827 15623 16833
rect 9525 16775 9633 16827
rect 9685 16775 9725 16827
rect 9777 16775 10860 16827
rect 10912 16775 12058 16827
rect 12110 16775 13846 16827
rect 13898 16775 15571 16827
rect 9525 16759 15623 16775
rect 9525 16707 9633 16759
rect 9685 16707 9725 16759
rect 9777 16707 10860 16759
rect 10912 16707 12058 16759
rect 12110 16707 13846 16759
rect 13898 16707 15571 16759
rect 9525 16691 15623 16707
rect 9525 16639 9633 16691
rect 9685 16639 9725 16691
rect 9777 16639 10860 16691
rect 10912 16639 12058 16691
rect 12110 16639 13846 16691
rect 13898 16639 15571 16691
rect 9525 16633 15623 16639
rect 8333 14925 8342 14981
rect 8398 14925 8424 14981
rect 8480 14925 8506 14981
rect 8562 14925 8587 14981
rect 8643 14925 8668 14981
rect 8724 14925 8733 14981
rect 8333 14837 8733 14925
rect 8333 14781 8342 14837
rect 8398 14781 8424 14837
rect 8480 14781 8506 14837
rect 8562 14781 8587 14837
rect 8643 14781 8668 14837
rect 8724 14781 8733 14837
rect 385 14719 7026 14725
rect 437 14667 2464 14719
rect 2516 14667 4606 14719
rect 4658 14667 6745 14719
rect 6797 14667 7026 14719
rect 385 14651 7026 14667
rect 437 14599 2464 14651
rect 2516 14599 4606 14651
rect 4658 14599 6745 14651
rect 6797 14599 7026 14651
rect 385 14583 7026 14599
rect 437 14531 2464 14583
rect 2516 14531 4606 14583
rect 4658 14531 6745 14583
rect 6797 14531 7026 14583
rect 385 14525 7026 14531
rect 7813 14669 7822 14725
rect 7878 14669 7904 14725
rect 7960 14669 7986 14725
rect 8042 14669 8067 14725
rect 8123 14669 8148 14725
rect 8204 14669 8213 14725
rect 7813 14581 8213 14669
rect 7813 14525 7822 14581
rect 7878 14525 7904 14581
rect 7960 14525 7986 14581
rect 8042 14525 8067 14581
rect 8123 14525 8148 14581
rect 8204 14525 8213 14581
rect 9498 14719 15623 14725
rect 9498 14667 9633 14719
rect 9685 14667 9725 14719
rect 9777 14667 10860 14719
rect 10912 14667 12058 14719
rect 12110 14667 13846 14719
rect 13898 14667 15571 14719
rect 9498 14651 15623 14667
rect 9498 14599 9633 14651
rect 9685 14599 9725 14651
rect 9777 14599 10860 14651
rect 10912 14599 12058 14651
rect 12110 14599 13846 14651
rect 13898 14599 15571 14651
rect 9498 14583 15623 14599
rect 9498 14531 9633 14583
rect 9685 14531 9725 14583
rect 9777 14531 10860 14583
rect 10912 14531 12058 14583
rect 12110 14531 13846 14583
rect 13898 14531 15571 14583
rect 9498 14525 15623 14531
rect 3243 13895 7245 13901
rect 3295 13849 7245 13895
rect 9294 13895 10490 13901
rect 9294 13849 10438 13895
rect 3295 13843 3323 13849
tri 3323 13843 3329 13849 nw
tri 7210 13843 7216 13849 ne
rect 7216 13843 7244 13849
rect 3243 13831 3311 13843
tri 3311 13831 3323 13843 nw
tri 7216 13831 7228 13843 ne
rect 7228 13831 7244 13843
tri 3295 13815 3311 13831 nw
tri 7228 13815 7244 13831 ne
rect 9302 13843 9330 13849
tri 9330 13843 9336 13849 nw
tri 10404 13843 10410 13849 ne
rect 10410 13843 10438 13849
rect 9302 13831 9318 13843
tri 9318 13831 9330 13843 nw
tri 10410 13831 10422 13843 ne
rect 10422 13831 10490 13843
tri 9302 13815 9318 13831 nw
tri 10422 13815 10438 13831 ne
rect 3243 13773 3295 13779
rect 10438 13773 10490 13779
tri 7210 12933 7244 12967 se
tri 9302 12933 9336 12967 sw
rect 3479 12927 7245 12933
rect 3531 12881 7245 12927
rect 9271 12927 10726 12933
rect 9271 12881 10674 12927
rect 3531 12875 3559 12881
tri 3559 12875 3565 12881 nw
tri 10640 12875 10646 12881 ne
rect 10646 12875 10674 12881
rect 3479 12863 3547 12875
tri 3547 12863 3559 12875 nw
tri 10646 12863 10658 12875 ne
rect 10658 12863 10726 12875
tri 3531 12847 3547 12863 nw
tri 10658 12847 10674 12863 ne
rect 3479 12805 3531 12811
rect 10674 12805 10726 12811
rect 8333 12201 8342 12257
rect 8398 12201 8424 12257
rect 8480 12201 8506 12257
rect 8562 12201 8587 12257
rect 8643 12201 8668 12257
rect 8724 12201 8733 12257
rect 8333 12113 8733 12201
rect 8333 12057 8342 12113
rect 8398 12057 8424 12113
rect 8480 12057 8506 12113
rect 8562 12057 8587 12113
rect 8643 12057 8668 12113
rect 8724 12057 8733 12113
rect 385 11995 7026 12001
rect 437 11943 2464 11995
rect 2516 11943 4606 11995
rect 4658 11943 6745 11995
rect 6797 11943 7026 11995
rect 385 11927 7026 11943
rect 437 11875 2464 11927
rect 2516 11875 4606 11927
rect 4658 11875 6745 11927
rect 6797 11875 7026 11927
rect 385 11859 7026 11875
rect 437 11807 2464 11859
rect 2516 11807 4606 11859
rect 4658 11807 6745 11859
rect 6797 11807 7026 11859
rect 385 11801 7026 11807
rect 7813 11945 7822 12001
rect 7878 11945 7904 12001
rect 7960 11945 7986 12001
rect 8042 11945 8067 12001
rect 8123 11945 8148 12001
rect 8204 11945 8213 12001
rect 7813 11857 8213 11945
rect 7813 11801 7822 11857
rect 7878 11801 7904 11857
rect 7960 11801 7986 11857
rect 8042 11801 8067 11857
rect 8123 11801 8148 11857
rect 8204 11801 8213 11857
rect 9498 11995 15623 12001
rect 9498 11943 9633 11995
rect 9685 11943 9725 11995
rect 9777 11943 10860 11995
rect 10912 11943 12058 11995
rect 12110 11943 13846 11995
rect 13898 11943 15571 11995
rect 9498 11927 15623 11943
rect 9498 11875 9633 11927
rect 9685 11875 9725 11927
rect 9777 11875 10860 11927
rect 10912 11875 12058 11927
rect 12110 11875 13846 11927
rect 13898 11875 15571 11927
rect 9498 11859 15623 11875
rect 9498 11807 9633 11859
rect 9685 11807 9725 11859
rect 9777 11807 10860 11859
rect 10912 11807 12058 11859
rect 12110 11807 13846 11859
rect 13898 11807 15571 11859
rect 9498 11801 15623 11807
rect 8333 10093 8342 10149
rect 8398 10093 8424 10149
rect 8480 10093 8506 10149
rect 8562 10093 8587 10149
rect 8643 10093 8668 10149
rect 8724 10093 8733 10149
rect 8333 10005 8733 10093
rect 8333 9949 8342 10005
rect 8398 9949 8424 10005
rect 8480 9949 8506 10005
rect 8562 9949 8587 10005
rect 8643 9949 8668 10005
rect 8724 9949 8733 10005
rect 385 9887 7026 9893
rect 437 9835 2464 9887
rect 2516 9835 4606 9887
rect 4658 9835 6745 9887
rect 6797 9835 7026 9887
rect 385 9819 7026 9835
rect 437 9767 2464 9819
rect 2516 9767 4606 9819
rect 4658 9767 6745 9819
rect 6797 9767 7026 9819
rect 385 9751 7026 9767
rect 437 9699 2464 9751
rect 2516 9699 4606 9751
rect 4658 9699 6745 9751
rect 6797 9699 7026 9751
rect 385 9693 7026 9699
rect 7813 9837 7822 9893
rect 7878 9837 7904 9893
rect 7960 9837 7986 9893
rect 8042 9837 8067 9893
rect 8123 9837 8148 9893
rect 8204 9837 8213 9893
rect 7813 9749 8213 9837
rect 7813 9693 7822 9749
rect 7878 9693 7904 9749
rect 7960 9693 7986 9749
rect 8042 9693 8067 9749
rect 8123 9693 8148 9749
rect 8204 9693 8213 9749
rect 9498 9887 15623 9893
rect 9498 9835 9633 9887
rect 9685 9835 9725 9887
rect 9777 9835 10860 9887
rect 10912 9835 12058 9887
rect 12110 9835 13846 9887
rect 13898 9835 15571 9887
rect 9498 9819 15623 9835
rect 9498 9767 9633 9819
rect 9685 9767 9725 9819
rect 9777 9767 10860 9819
rect 10912 9767 12058 9819
rect 12110 9767 13846 9819
rect 13898 9767 15571 9819
rect 9498 9751 15623 9767
rect 9498 9699 9633 9751
rect 9685 9699 9725 9751
rect 9777 9699 10860 9751
rect 10912 9699 12058 9751
rect 12110 9699 13846 9751
rect 13898 9699 15571 9751
rect 9498 9693 15623 9699
rect 3715 9063 7245 9069
rect 3767 9017 7245 9063
rect 9294 9063 11216 9069
rect 9294 9017 11164 9063
rect 3767 9011 3795 9017
tri 3795 9011 3801 9017 nw
tri 7210 9011 7216 9017 ne
rect 7216 9011 7244 9017
rect 3715 8999 3783 9011
tri 3783 8999 3795 9011 nw
tri 7216 8999 7228 9011 ne
rect 7228 8999 7244 9011
tri 3767 8983 3783 8999 nw
tri 7228 8983 7244 8999 ne
rect 9302 9011 9330 9017
tri 9330 9011 9336 9017 nw
tri 11130 9011 11136 9017 ne
rect 11136 9011 11164 9017
rect 9302 8999 9318 9011
tri 9318 8999 9330 9011 nw
tri 11136 8999 11148 9011 ne
rect 11148 8999 11216 9011
tri 9302 8983 9318 8999 nw
tri 11148 8983 11164 8999 ne
rect 3715 8941 3767 8947
rect 11164 8941 11216 8947
tri 7210 8101 7244 8135 se
tri 9302 8101 9336 8135 sw
rect 3951 8095 7245 8101
rect 4003 8049 7245 8095
rect 9271 8095 11452 8101
rect 9271 8049 11400 8095
rect 4003 8043 4031 8049
tri 4031 8043 4037 8049 nw
tri 11366 8043 11372 8049 ne
rect 11372 8043 11400 8049
rect 3951 8031 4019 8043
tri 4019 8031 4031 8043 nw
tri 11372 8031 11384 8043 ne
rect 11384 8031 11452 8043
tri 4003 8015 4019 8031 nw
tri 11384 8015 11400 8031 ne
rect 3951 7973 4003 7979
rect 11400 7973 11452 7979
rect 7814 7729 12836 7746
rect 7814 7673 7823 7729
rect 7879 7673 7932 7729
rect 7988 7673 8040 7729
rect 8096 7673 8148 7729
rect 8204 7727 12836 7729
rect 8204 7675 12642 7727
rect 12694 7675 12710 7727
rect 12762 7675 12778 7727
rect 12830 7675 12836 7727
rect 8204 7673 12836 7675
rect 7814 7656 12836 7673
tri 3502 7225 3702 7425 se
rect 3702 7225 7021 7425
rect 8333 7369 8342 7425
rect 8398 7369 8424 7425
rect 8480 7369 8506 7425
rect 8562 7369 8587 7425
rect 8643 7369 8668 7425
rect 8724 7369 8733 7425
rect 8333 7281 8733 7369
rect 8333 7225 8342 7281
rect 8398 7225 8424 7281
rect 8480 7225 8506 7281
rect 8562 7225 8587 7281
rect 8643 7225 8668 7281
rect 8724 7225 8733 7281
tri 3446 7169 3502 7225 se
rect 3502 7169 3728 7225
tri 3728 7169 3784 7225 nw
tri 3440 7163 3446 7169 se
rect 3446 7163 3722 7169
tri 3722 7163 3728 7169 nw
tri 3420 7143 3440 7163 se
rect 3440 7143 3702 7163
tri 3702 7143 3722 7163 nw
tri 3388 7111 3420 7143 se
rect 3420 7111 3670 7143
tri 3670 7111 3702 7143 nw
rect 7813 7113 7822 7169
rect 7878 7113 7904 7169
rect 7960 7113 7986 7169
rect 8042 7113 8067 7169
rect 8123 7113 8148 7169
rect 8204 7113 8213 7169
tri 3372 7095 3388 7111 se
rect 3388 7095 3654 7111
tri 3654 7095 3670 7111 nw
tri 3320 7043 3372 7095 se
rect 3372 7043 3602 7095
tri 3602 7043 3654 7095 nw
tri 3304 7027 3320 7043 se
rect 3320 7027 3586 7043
tri 3586 7027 3602 7043 nw
tri 3252 6975 3304 7027 se
rect 3304 6975 3534 7027
tri 3534 6975 3586 7027 nw
rect 7813 7025 8213 7113
tri 3246 6969 3252 6975 se
rect 3252 6969 3528 6975
tri 3528 6969 3534 6975 nw
rect 7813 6969 7822 7025
rect 7878 6969 7904 7025
rect 7960 6969 7986 7025
rect 8042 6969 8067 7025
rect 8123 6969 8148 7025
rect 8204 6969 8213 7025
rect 9487 7163 13701 7169
rect 9487 7111 9633 7163
rect 9685 7111 13701 7163
rect 9487 7095 13701 7111
rect 9487 7043 9633 7095
rect 9685 7043 13701 7095
rect 9487 7027 13701 7043
rect 9487 6975 9633 7027
rect 9685 6975 13701 7027
rect 9487 6969 13701 6975
tri 3138 6861 3246 6969 se
rect 3246 6861 3420 6969
tri 3420 6861 3528 6969 nw
tri 13087 6861 13195 6969 ne
rect 13195 6861 13701 6969
tri 3032 6755 3138 6861 se
rect 3138 6755 3314 6861
tri 3314 6755 3420 6861 nw
tri 13195 6755 13301 6861 ne
tri 2856 6579 3032 6755 se
rect 3032 6579 3138 6755
tri 3138 6579 3314 6755 nw
tri 2832 6555 2856 6579 se
rect 2856 6555 3114 6579
tri 3114 6555 3138 6579 nw
rect 2832 3933 3032 6555
tri 3032 6473 3114 6555 nw
rect 3068 6188 7939 6194
rect 3068 6142 7887 6188
rect 3068 6136 3148 6142
tri 3148 6136 3154 6142 nw
tri 7853 6136 7859 6142 ne
rect 7859 6136 7887 6142
rect 3068 6124 3136 6136
tri 3136 6124 3148 6136 nw
tri 7859 6124 7871 6136 ne
rect 7871 6124 7939 6136
rect 547 3683 553 3735
rect 605 3683 621 3735
rect 673 3683 688 3735
rect 740 3683 755 3735
rect 807 3683 822 3735
rect 874 3683 889 3735
rect 941 3683 947 3735
rect 547 3657 947 3683
rect 547 3605 553 3657
rect 605 3605 621 3657
rect 673 3605 688 3657
rect 740 3605 755 3657
rect 807 3605 822 3657
rect 874 3605 889 3657
rect 941 3605 947 3657
rect 547 2698 947 3605
rect 547 2642 548 2698
rect 604 2642 662 2698
rect 718 2642 776 2698
rect 832 2642 890 2698
rect 946 2642 947 2698
rect 547 2576 947 2642
rect 547 2520 548 2576
rect 604 2520 662 2576
rect 718 2520 776 2576
rect 832 2520 890 2576
rect 946 2520 947 2576
rect 547 2454 947 2520
rect 547 2398 548 2454
rect 604 2398 662 2454
rect 718 2398 776 2454
rect 832 2398 890 2454
rect 946 2398 947 2454
rect 547 2332 947 2398
rect 547 2276 548 2332
rect 604 2276 662 2332
rect 718 2276 776 2332
rect 832 2276 890 2332
rect 946 2276 947 2332
rect 547 2271 947 2276
rect 547 2219 553 2271
rect 605 2219 621 2271
rect 673 2219 688 2271
rect 740 2219 755 2271
rect 807 2219 822 2271
rect 874 2219 889 2271
rect 941 2219 947 2271
rect 547 2210 947 2219
rect 547 2154 548 2210
rect 604 2197 662 2210
rect 718 2197 776 2210
rect 832 2197 890 2210
rect 547 2145 553 2154
rect 605 2145 621 2197
rect 673 2145 688 2154
rect 740 2145 755 2197
rect 807 2145 822 2154
rect 874 2145 889 2197
rect 946 2154 947 2210
rect 941 2145 947 2154
rect 547 2123 947 2145
rect 547 2088 553 2123
rect 547 2032 548 2088
rect 605 2071 621 2123
rect 673 2088 688 2123
rect 740 2071 755 2123
rect 807 2088 822 2123
rect 874 2071 889 2123
rect 941 2088 947 2123
rect 604 2032 662 2071
rect 718 2032 776 2071
rect 832 2032 890 2071
rect 946 2032 947 2088
rect 547 2014 947 2032
rect 547 1965 553 2014
rect 547 1909 548 1965
rect 605 1962 621 2014
rect 673 1965 688 2014
rect 740 1962 755 2014
rect 807 1965 822 2014
rect 874 1962 889 2014
rect 941 1965 947 2014
rect 604 1940 662 1962
rect 718 1940 776 1962
rect 832 1940 890 1962
rect 547 1888 553 1909
rect 605 1888 621 1940
rect 673 1888 688 1909
rect 740 1888 755 1940
rect 807 1888 822 1909
rect 874 1888 889 1940
rect 946 1909 947 1965
rect 941 1888 947 1909
rect 547 1866 947 1888
rect 547 1842 553 1866
rect 547 1786 548 1842
rect 605 1814 621 1866
rect 673 1842 688 1866
rect 740 1814 755 1866
rect 807 1842 822 1866
rect 874 1814 889 1866
rect 941 1842 947 1866
rect 604 1786 662 1814
rect 718 1786 776 1814
rect 832 1786 890 1814
rect 946 1786 947 1842
rect 547 479 947 1786
rect 547 427 553 479
rect 605 427 621 479
rect 673 427 688 479
rect 740 427 755 479
rect 807 427 822 479
rect 874 427 889 479
rect 941 427 947 479
rect 547 401 947 427
rect 547 349 553 401
rect 605 349 621 401
rect 673 349 688 401
rect 740 349 755 401
rect 807 349 822 401
rect 874 349 889 401
rect 941 349 947 401
rect 979 3410 1031 3416
rect 979 3346 1031 3358
rect 979 122 1031 3294
rect 979 58 1031 70
rect 979 0 1031 6
rect 1231 668 1237 720
rect 1289 668 1301 720
rect 1353 668 1359 720
rect 3068 705 3120 6124
tri 3120 6108 3136 6124 nw
tri 7871 6108 7887 6124 ne
rect 7887 6066 7939 6072
rect 3151 5303 8339 5309
rect 3151 5257 8287 5303
rect 3151 5251 3231 5257
tri 3231 5251 3237 5257 nw
tri 8253 5251 8259 5257 ne
rect 8259 5251 8287 5257
rect 3151 5239 3219 5251
tri 3219 5239 3231 5251 nw
tri 8259 5239 8271 5251 ne
rect 8271 5239 8339 5251
rect 3151 1004 3203 5239
tri 3203 5223 3219 5239 nw
tri 8271 5223 8287 5239 ne
rect 8287 5181 8339 5187
rect 3243 5147 8419 5153
rect 3243 5101 8367 5147
rect 3243 5095 3323 5101
tri 3323 5095 3329 5101 nw
tri 8333 5095 8339 5101 ne
rect 8339 5095 8367 5101
rect 3243 5083 3311 5095
tri 3311 5083 3323 5095 nw
tri 8339 5083 8351 5095 ne
rect 8351 5083 8419 5095
rect 3243 3132 3295 5083
tri 3295 5067 3311 5083 nw
tri 8351 5073 8361 5083 ne
rect 8361 5073 8367 5083
rect 3411 5067 8019 5073
tri 8361 5067 8367 5073 ne
rect 3411 5021 7967 5067
rect 3411 5015 3491 5021
tri 3491 5015 3497 5021 nw
tri 7933 5015 7939 5021 ne
rect 7939 5015 7967 5021
rect 8367 5025 8419 5031
rect 3411 5003 3479 5015
tri 3479 5003 3491 5015 nw
tri 7939 5003 7951 5015 ne
rect 7951 5003 8019 5015
rect 3411 4993 3469 5003
tri 3469 4993 3479 5003 nw
tri 7951 4993 7961 5003 ne
rect 7961 4993 7967 5003
tri 3401 3473 3411 3483 se
rect 3411 3473 3463 4993
tri 3463 4987 3469 4993 nw
rect 3531 4989 7799 4993
tri 7799 4989 7803 4993 sw
tri 7961 4989 7965 4993 ne
rect 7965 4989 7967 4993
tri 3389 3461 3401 3473 se
rect 3401 3461 3463 3473
tri 3377 3449 3389 3461 se
rect 3389 3449 3463 3461
rect 3335 3397 3341 3449
rect 3393 3397 3405 3449
rect 3457 3397 3463 3449
rect 3531 4951 7803 4989
tri 7803 4951 7841 4989 sw
tri 7965 4987 7967 4989 ne
rect 3531 4949 7841 4951
tri 7841 4949 7843 4951 sw
rect 3531 4941 7843 4949
rect 3531 4935 3611 4941
tri 3611 4935 3617 4941 nw
tri 7777 4935 7783 4941 ne
rect 7783 4935 7843 4941
tri 7843 4935 7857 4949 sw
rect 7967 4945 8019 4951
rect 8447 4987 8499 4993
tri 8443 4945 8447 4949 se
tri 8433 4935 8443 4945 se
rect 8443 4935 8447 4945
rect 3531 4923 3599 4935
tri 3599 4923 3611 4935 nw
tri 7783 4923 7795 4935 ne
rect 7795 4923 7857 4935
tri 7857 4923 7869 4935 sw
tri 8421 4923 8433 4935 se
rect 8433 4923 8499 4935
rect 3531 4915 3591 4923
tri 3591 4915 3599 4923 nw
tri 7795 4915 7803 4923 ne
rect 7803 4915 7869 4923
tri 7869 4915 7877 4923 sw
tri 8413 4915 8421 4923 se
rect 8421 4915 8447 4923
tri 3295 3132 3329 3166 sw
rect 3531 3132 3583 4915
tri 3583 4907 3591 4915 nw
tri 7803 4913 7805 4915 ne
rect 7805 4913 8447 4915
rect 3926 4907 7689 4913
tri 7689 4907 7695 4913 sw
tri 7805 4907 7811 4913 ne
rect 7811 4907 8447 4913
rect 3926 4902 7695 4907
tri 7695 4902 7700 4907 sw
tri 7811 4902 7816 4907 ne
rect 7816 4902 8447 4907
rect 3926 4871 7700 4902
tri 7700 4871 7731 4902 sw
tri 7816 4871 7847 4902 ne
rect 7847 4871 8447 4902
rect 3926 4863 7731 4871
tri 7731 4863 7739 4871 sw
tri 7847 4863 7855 4871 ne
rect 7855 4863 8499 4871
rect 3926 4861 7739 4863
rect 3926 4828 3979 4861
tri 3979 4828 4012 4861 nw
tri 7667 4828 7700 4861 ne
rect 7700 4828 7739 4861
tri 7739 4828 7774 4863 sw
tri 3916 3473 3926 3483 se
rect 3926 3473 3978 4828
tri 3978 4827 3979 4828 nw
tri 7700 4827 7701 4828 ne
rect 7701 4827 7774 4828
tri 7701 4824 7704 4827 ne
rect 7704 4824 7774 4827
tri 7774 4824 7778 4828 sw
rect 8047 4824 8099 4830
tri 7704 4793 7735 4824 ne
rect 7735 4793 7778 4824
tri 4341 4772 4362 4793 se
rect 4362 4772 5051 4793
tri 5051 4772 5072 4793 sw
tri 7735 4772 7756 4793 ne
rect 7756 4788 7778 4793
tri 7778 4788 7814 4824 sw
rect 7756 4772 7814 4788
tri 7814 4772 7830 4788 sw
tri 8031 4772 8047 4788 se
tri 4329 4760 4341 4772 se
rect 4341 4760 5072 4772
tri 5072 4760 5084 4772 sw
tri 7756 4760 7768 4772 ne
rect 7768 4760 7830 4772
tri 7830 4760 7842 4772 sw
tri 8019 4760 8031 4772 se
rect 8031 4760 8099 4772
tri 4322 4753 4329 4760 se
rect 4329 4754 5084 4760
tri 5084 4754 5090 4760 sw
tri 7768 4754 7774 4760 ne
rect 7774 4754 7842 4760
tri 7842 4754 7848 4760 sw
tri 8013 4754 8019 4760 se
rect 8019 4754 8047 4760
rect 4329 4753 5090 4754
tri 5090 4753 5091 4754 sw
tri 7774 4753 7775 4754 ne
rect 7775 4753 8047 4754
tri 4299 4730 4322 4753 se
rect 4322 4741 5091 4753
rect 4322 4730 4373 4741
tri 4373 4730 4384 4741 nw
tri 5029 4730 5040 4741 ne
rect 5040 4730 5091 4741
rect 4299 4695 4351 4730
tri 4351 4708 4373 4730 nw
tri 5040 4708 5062 4730 ne
rect 5062 4708 5091 4730
tri 5091 4708 5136 4753 sw
tri 7775 4708 7820 4753 ne
rect 7820 4708 8047 4753
tri 5062 4694 5076 4708 ne
rect 5076 4702 5136 4708
tri 5136 4702 5142 4708 sw
tri 7820 4702 7826 4708 ne
rect 7826 4702 8099 4708
rect 5076 4694 5142 4702
tri 5142 4694 5150 4702 sw
rect 11694 4694 11746 4700
tri 5076 4679 5091 4694 ne
rect 5091 4679 5150 4694
tri 5150 4679 5165 4694 sw
tri 5091 4669 5101 4679 ne
rect 5101 4669 5165 4679
tri 5101 4657 5113 4669 ne
rect 4299 4631 4351 4643
rect 4299 4573 4351 4579
tri 4758 4539 4792 4573 ne
rect 4792 4299 4844 4590
rect 5113 4380 5165 4669
rect 11694 4630 11746 4642
tri 11632 4447 11694 4509 se
rect 11694 4487 11746 4578
rect 11694 4447 11706 4487
tri 11706 4447 11746 4487 nw
tri 9713 4402 9758 4447 se
rect 9758 4402 11654 4447
tri 5113 4333 5160 4380 ne
rect 5160 4373 5165 4380
tri 5165 4373 5194 4402 sw
tri 9684 4373 9713 4402 se
rect 9713 4395 11654 4402
tri 11654 4395 11706 4447 nw
rect 9713 4373 9758 4395
tri 9758 4373 9780 4395 nw
rect 5160 4354 5194 4373
tri 5194 4354 5213 4373 sw
tri 9665 4354 9684 4373 se
rect 9684 4354 9739 4373
tri 9739 4354 9758 4373 nw
rect 5160 4333 5213 4354
tri 5213 4333 5234 4354 sw
tri 9644 4333 9665 4354 se
rect 9665 4333 9705 4354
tri 5160 4328 5165 4333 ne
rect 5165 4328 7296 4333
tri 5165 4320 5173 4328 ne
rect 5173 4320 7296 4328
tri 9631 4320 9644 4333 se
rect 9644 4320 9705 4333
tri 9705 4320 9739 4354 nw
tri 11838 4320 11872 4354 se
rect 11872 4320 11924 4584
tri 11924 4540 11958 4574 nw
tri 5173 4313 5180 4320 ne
rect 5180 4313 7296 4320
tri 4844 4299 4858 4313 sw
tri 5180 4299 5194 4313 ne
rect 5194 4299 7296 4313
tri 9610 4299 9631 4320 se
rect 9631 4299 9684 4320
tri 9684 4299 9705 4320 nw
rect 4792 4291 4858 4299
tri 4792 4268 4815 4291 ne
rect 4815 4281 4858 4291
tri 4858 4281 4876 4299 sw
tri 5194 4281 5212 4299 ne
rect 5212 4281 7296 4299
rect 4815 4271 4876 4281
tri 4876 4271 4886 4281 sw
tri 7210 4271 7220 4281 ne
rect 7220 4271 7296 4281
tri 9582 4271 9610 4299 se
rect 9610 4271 9653 4299
rect 4815 4268 4886 4271
tri 4886 4268 4889 4271 sw
tri 7220 4268 7223 4271 ne
rect 7223 4268 7296 4271
tri 7296 4268 7299 4271 sw
tri 9579 4268 9582 4271 se
rect 9582 4268 9653 4271
tri 9653 4268 9684 4299 nw
rect 9847 4268 9853 4320
rect 9905 4268 9917 4320
rect 9969 4268 11924 4320
tri 4815 4239 4844 4268 ne
rect 4844 4247 4889 4268
tri 4889 4247 4910 4268 sw
tri 7223 4247 7244 4268 ne
rect 4844 4239 4910 4247
tri 4910 4239 4918 4247 sw
tri 4844 4187 4896 4239 ne
rect 4896 4187 6675 4239
rect 6727 4187 6739 4239
rect 6791 4187 6797 4239
rect 7244 4237 7299 4268
tri 7299 4237 7330 4268 sw
tri 9548 4237 9579 4268 se
rect 9579 4237 9622 4268
tri 9622 4237 9653 4268 nw
rect 7244 4226 7296 4237
rect 9302 4185 9570 4237
tri 9570 4185 9622 4237 nw
tri 9302 4151 9336 4185 nw
rect 5336 3964 6684 3965
rect 5336 3912 5342 3964
rect 5394 3912 5429 3964
rect 5481 3912 5516 3964
rect 5568 3958 6684 3964
rect 5568 3912 6484 3958
rect 5336 3906 6484 3912
rect 6536 3906 6558 3958
rect 6610 3906 6632 3958
rect 5336 3890 6684 3906
rect 5336 3838 5342 3890
rect 5394 3838 5429 3890
rect 5481 3838 5516 3890
rect 5568 3838 6484 3890
rect 6536 3838 6558 3890
rect 6610 3838 6632 3890
rect 5336 3821 6684 3838
rect 5336 3816 6484 3821
rect 5336 3764 5342 3816
rect 5394 3764 5429 3816
rect 5481 3764 5516 3816
rect 5568 3769 6484 3816
rect 6536 3769 6558 3821
rect 6610 3769 6632 3821
rect 5568 3764 6684 3769
rect 5336 3763 6684 3764
tri 3904 3461 3916 3473 se
rect 3916 3461 3978 3473
tri 3898 3455 3904 3461 se
rect 3904 3455 3978 3461
tri 3892 3449 3898 3455 se
rect 3898 3449 3978 3455
rect 3850 3397 3856 3449
rect 3908 3397 3920 3449
rect 3972 3397 3978 3449
rect 8127 3525 8179 3531
tri 8179 3486 8182 3489 sw
rect 11899 3486 11951 3492
rect 8179 3473 8182 3486
rect 8127 3461 8182 3473
rect 5417 3364 5423 3416
rect 5475 3364 5487 3416
rect 5539 3409 5799 3416
tri 5799 3409 5806 3416 sw
rect 8179 3455 8182 3461
tri 8182 3455 8213 3486 sw
rect 8179 3409 9923 3455
rect 5539 3403 5806 3409
tri 5806 3403 5812 3409 sw
rect 8127 3403 9923 3409
rect 9975 3403 9987 3455
rect 10039 3403 10045 3455
rect 11899 3422 11951 3434
rect 5539 3397 5812 3403
tri 5812 3397 5818 3403 sw
rect 5539 3377 5818 3397
tri 5818 3377 5838 3397 sw
rect 5539 3370 5838 3377
tri 5838 3370 5845 3377 sw
tri 11951 3416 11985 3450 sw
rect 11951 3370 13132 3416
rect 5539 3364 5845 3370
tri 5845 3364 5851 3370 sw
rect 11899 3364 13132 3370
tri 5777 3339 5802 3364 ne
rect 5802 3345 5851 3364
tri 5851 3345 5870 3364 sw
tri 13046 3345 13065 3364 ne
rect 13065 3345 13132 3364
rect 5802 3339 5870 3345
tri 5870 3339 5876 3345 sw
rect 6745 3339 6797 3345
tri 5802 3303 5838 3339 ne
rect 5838 3303 5876 3339
tri 5876 3303 5912 3339 sw
tri 5838 3287 5854 3303 ne
rect 5854 3287 5912 3303
tri 5912 3287 5928 3303 sw
rect 9793 3339 9845 3345
tri 6797 3287 6813 3303 sw
tri 7228 3287 7244 3303 se
tri 5854 3275 5866 3287 ne
rect 5866 3275 5928 3287
tri 5928 3275 5940 3287 sw
rect 6745 3275 6813 3287
tri 6813 3275 6825 3287 sw
tri 7216 3275 7228 3287 se
rect 7228 3275 7244 3287
tri 5866 3229 5912 3275 ne
rect 5912 3229 5940 3275
tri 5940 3229 5986 3275 sw
tri 5912 3223 5918 3229 ne
rect 5918 3223 5986 3229
tri 5986 3223 5992 3229 sw
rect 6797 3269 6825 3275
tri 6825 3269 6831 3275 sw
tri 7210 3269 7216 3275 se
rect 7216 3269 7244 3275
tri 9302 3287 9318 3303 sw
tri 9777 3287 9793 3303 se
tri 13065 3330 13080 3345 ne
rect 9302 3275 9318 3287
tri 9318 3275 9330 3287 sw
tri 9765 3275 9777 3287 se
rect 9777 3275 9845 3287
rect 9302 3269 9330 3275
tri 9330 3269 9336 3275 sw
tri 9759 3269 9765 3275 se
rect 9765 3269 9793 3275
rect 6797 3223 7253 3269
tri 5918 3166 5975 3223 ne
rect 5975 3217 5992 3223
tri 5992 3217 5998 3223 sw
rect 6745 3217 7253 3223
rect 9295 3223 9793 3269
rect 9295 3217 9845 3223
rect 5975 3166 5998 3217
tri 5998 3166 6049 3217 sw
tri 3583 3132 3617 3166 sw
tri 5975 3155 5986 3166 ne
rect 5986 3155 6049 3166
tri 6049 3155 6060 3166 sw
tri 5986 3132 6009 3155 ne
rect 6009 3132 6060 3155
tri 6060 3132 6083 3155 sw
rect 3243 3080 3249 3132
rect 3301 3080 3313 3132
rect 3365 3080 3371 3132
rect 3531 3080 3537 3132
rect 3589 3080 3601 3132
rect 3653 3080 3659 3132
tri 6009 3093 6048 3132 ne
rect 6048 3093 6083 3132
tri 6083 3093 6122 3132 sw
tri 9813 3093 9852 3132 se
rect 9852 3093 9923 3132
tri 6048 3081 6060 3093 ne
rect 6060 3081 6122 3093
tri 6122 3081 6134 3093 sw
tri 9801 3081 9813 3093 se
rect 9813 3081 9923 3093
tri 6060 3080 6061 3081 ne
rect 6061 3080 6134 3081
tri 6134 3080 6135 3081 sw
tri 9800 3080 9801 3081 se
rect 9801 3080 9923 3081
rect 9975 3080 9987 3132
rect 10039 3080 10045 3132
tri 6061 3007 6134 3080 ne
rect 6134 3058 6135 3080
tri 6135 3058 6157 3080 sw
tri 9778 3058 9800 3080 se
rect 9800 3058 9852 3080
tri 9852 3058 9874 3080 nw
rect 6134 3007 6157 3058
tri 6157 3007 6208 3058 sw
tri 9727 3007 9778 3058 se
tri 6134 3001 6140 3007 ne
rect 6140 3001 6797 3007
tri 6140 2967 6174 3001 ne
rect 6174 2967 6745 3001
rect 5416 2961 5574 2967
rect 5468 2909 5522 2961
tri 6174 2955 6186 2967 ne
rect 6186 2955 6745 2967
tri 6711 2949 6717 2955 ne
rect 6717 2949 6745 2955
tri 9704 2984 9727 3007 se
rect 9727 2984 9778 3007
tri 9778 2984 9852 3058 nw
tri 9687 2967 9704 2984 se
rect 9704 2967 9761 2984
tri 9761 2967 9778 2984 nw
tri 9681 2961 9687 2967 se
rect 9687 2961 9755 2967
tri 9755 2961 9761 2967 nw
rect 11988 2961 12834 2967
tri 6717 2937 6729 2949 ne
rect 6729 2937 6797 2949
tri 6729 2921 6745 2937 ne
rect 5416 2894 5574 2909
rect 5468 2842 5522 2894
tri 9630 2910 9681 2961 se
rect 9681 2910 9704 2961
tri 9704 2910 9755 2961 nw
tri 9629 2909 9630 2910 se
rect 9630 2909 9703 2910
tri 9703 2909 9704 2910 nw
rect 11988 2909 12637 2961
rect 12689 2909 12709 2961
rect 12761 2909 12781 2961
rect 12833 2909 12834 2961
tri 9614 2894 9629 2909 se
rect 9629 2894 9688 2909
tri 9688 2894 9703 2909 nw
rect 11988 2894 12834 2909
rect 6745 2879 6797 2885
tri 9599 2879 9614 2894 se
rect 9614 2879 9670 2894
tri 9596 2876 9599 2879 se
rect 9599 2876 9670 2879
tri 9670 2876 9688 2894 nw
rect 5416 2826 5574 2842
rect 5468 2774 5522 2826
rect 5416 2467 5574 2774
rect 8527 2870 9636 2876
rect 8579 2842 9636 2870
tri 9636 2842 9670 2876 nw
rect 11988 2842 12637 2894
rect 12689 2842 12709 2894
rect 12761 2842 12781 2894
rect 12833 2842 12834 2894
rect 8579 2826 9620 2842
tri 9620 2826 9636 2842 nw
rect 11988 2826 12834 2842
rect 8579 2824 9618 2826
tri 9618 2824 9620 2826 nw
rect 8527 2806 8579 2818
tri 8579 2790 8613 2824 nw
rect 11988 2774 12637 2826
rect 12689 2774 12709 2826
rect 12761 2774 12781 2826
rect 12833 2774 12834 2826
rect 11988 2768 12834 2774
rect 8527 2748 8579 2754
rect 11994 2748 12028 2768
tri 12028 2748 12048 2768 nw
tri 11994 2714 12028 2748 nw
rect 11642 2698 11770 2707
rect 11642 2642 11678 2698
rect 11734 2642 11770 2698
rect 6484 2587 7040 2593
rect 6536 2535 6558 2587
rect 6610 2535 6632 2587
rect 6684 2535 7040 2587
rect 6484 2519 7040 2535
tri 5574 2467 5599 2492 sw
rect 6536 2467 6558 2519
rect 6610 2467 6632 2519
rect 6684 2467 7040 2519
rect 5416 2451 5599 2467
tri 5599 2451 5615 2467 sw
rect 6484 2451 7040 2467
rect 5416 2399 5615 2451
tri 5615 2399 5667 2451 sw
rect 6536 2399 6558 2451
rect 6610 2399 6632 2451
rect 6684 2399 7040 2451
rect 5416 2393 5667 2399
tri 5667 2393 5673 2399 sw
rect 6484 2393 7040 2399
rect 8333 2537 8342 2593
rect 8398 2537 8424 2593
rect 8480 2537 8506 2593
rect 8562 2537 8587 2593
rect 8643 2537 8668 2593
rect 8724 2537 8733 2593
rect 8333 2449 8733 2537
rect 8333 2393 8342 2449
rect 8398 2393 8424 2449
rect 8480 2393 8506 2449
rect 8562 2393 8587 2449
rect 8643 2393 8668 2449
rect 8724 2393 8733 2449
rect 9459 2408 9758 2593
tri 9758 2408 9943 2593 sw
rect 9459 2393 9943 2408
rect 5416 2368 5673 2393
tri 5416 2337 5447 2368 ne
rect 5447 2337 5673 2368
tri 5673 2337 5729 2393 sw
tri 9676 2337 9732 2393 ne
rect 9732 2337 9943 2393
tri 5447 2210 5574 2337 ne
rect 5574 2210 7122 2337
tri 5574 2137 5647 2210 ne
rect 5647 2137 7122 2210
rect 7813 2281 7822 2337
rect 7878 2281 7904 2337
rect 7960 2281 7986 2337
rect 8042 2281 8067 2337
rect 8123 2281 8148 2337
rect 8204 2281 8213 2337
tri 9732 2326 9743 2337 ne
rect 7813 2193 8213 2281
rect 7813 2137 7822 2193
rect 7878 2137 7904 2193
rect 7960 2137 7986 2193
rect 8042 2137 8067 2193
rect 8123 2137 8148 2193
rect 8204 2137 8213 2193
rect 9743 2119 9943 2337
rect 11642 2576 11770 2642
rect 11642 2520 11678 2576
rect 11734 2520 11770 2576
rect 11642 2454 11770 2520
rect 11642 2398 11678 2454
rect 11734 2398 11770 2454
rect 11642 2332 11770 2398
rect 11642 2276 11678 2332
rect 11734 2276 11770 2332
tri 10288 2156 10376 2244 se
tri 9943 2119 9980 2156 sw
tri 10251 2119 10288 2156 se
rect 10288 2119 10376 2156
rect 9743 2074 9980 2119
tri 9980 2074 10025 2119 sw
tri 10206 2074 10251 2119 se
rect 10251 2074 10376 2119
tri 9743 2037 9780 2074 ne
rect 9780 2037 10025 2074
tri 10025 2037 10062 2074 sw
tri 10169 2037 10206 2074 se
rect 10206 2037 10376 2074
tri 9780 1937 9880 2037 ne
rect 9880 1937 10376 2037
rect 5818 1885 5824 1937
rect 5876 1885 5888 1937
rect 5940 1885 6110 1937
tri 6088 1877 6096 1885 ne
rect 6096 1877 6110 1885
tri 6110 1877 6170 1937 sw
tri 9880 1877 9940 1937 ne
rect 9940 1877 10376 1937
tri 6096 1863 6110 1877 ne
rect 6110 1863 6170 1877
tri 6110 1803 6170 1863 ne
tri 6170 1837 6210 1877 sw
tri 9940 1837 9980 1877 ne
rect 9980 1837 10376 1877
rect 6170 1803 6210 1837
tri 6210 1803 6244 1837 sw
tri 6170 1796 6177 1803 ne
rect 6177 1796 6244 1803
tri 10169 1796 10210 1837 ne
rect 10210 1796 10376 1837
tri 6177 1795 6178 1796 ne
rect 6178 1795 6244 1796
tri 10210 1795 10211 1796 ne
rect 10211 1795 10376 1796
tri 6178 1781 6192 1795 ne
rect 3783 1540 4730 1592
rect 3783 1507 3836 1540
tri 3836 1507 3869 1540 nw
tri 4644 1507 4677 1540 ne
rect 4677 1507 4730 1540
tri 3203 1004 3237 1038 sw
tri 3749 1004 3783 1038 se
rect 3783 1004 3835 1507
tri 3835 1506 3836 1507 nw
tri 4677 1506 4678 1507 ne
rect 3151 952 3157 1004
rect 3209 952 3221 1004
rect 3273 952 3279 1004
rect 3707 952 3713 1004
rect 3765 952 3777 1004
rect 3829 952 3835 1004
rect 3926 1385 4631 1437
tri 3920 715 3926 721 se
rect 3926 715 3978 1385
tri 3978 1351 4012 1385 nw
tri 4545 1351 4579 1385 ne
tri 3120 705 3130 715 sw
tri 3910 705 3920 715 se
rect 3920 705 3978 715
rect 3068 696 3130 705
tri 3130 696 3139 705 sw
tri 3901 696 3910 705 se
rect 3910 696 3978 705
rect 3068 687 3139 696
tri 3139 687 3148 696 sw
tri 3892 687 3901 696 se
rect 3901 687 3978 696
rect 3068 681 3148 687
tri 3148 681 3154 687 sw
rect 1231 635 1284 668
tri 1284 635 1317 668 nw
rect 1231 122 1283 635
tri 1283 634 1284 635 nw
rect 3068 629 3074 681
rect 3126 629 3138 681
rect 3190 629 3196 681
rect 3850 635 3856 687
rect 3908 635 3920 687
rect 3972 635 3978 687
rect 4579 343 4631 1385
rect 4678 410 4730 1507
rect 5476 547 5482 599
rect 5534 547 5546 599
rect 5598 547 5989 599
rect 6041 547 6053 599
rect 6105 547 6111 599
tri 4678 407 4681 410 ne
rect 4681 407 4730 410
tri 4730 407 4755 432 sw
tri 4681 395 4693 407 ne
rect 4693 395 4755 407
tri 4755 395 4767 407 sw
tri 4693 371 4717 395 ne
rect 4717 371 4767 395
tri 4767 371 4791 395 sw
tri 4717 358 4730 371 ne
rect 4730 358 4791 371
tri 4730 348 4740 358 ne
rect 4740 348 4791 358
tri 4631 343 4636 348 sw
tri 4740 343 4745 348 ne
rect 4745 343 4791 348
tri 4791 343 4819 371 sw
rect 4579 326 4636 343
tri 4579 320 4585 326 ne
rect 4585 320 4636 326
tri 4636 320 4659 343 sw
tri 4745 320 4768 343 ne
rect 4768 337 4819 343
tri 4819 337 4825 343 sw
rect 4768 331 4825 337
tri 4825 331 4831 337 sw
rect 4768 320 4831 331
tri 4831 320 4842 331 sw
tri 6181 320 6192 331 se
rect 6192 320 6244 1795
tri 10211 1743 10263 1795 ne
rect 10263 1743 10376 1795
rect 11642 2210 11770 2276
rect 11642 2154 11678 2210
rect 11734 2154 11770 2210
rect 11642 2088 11770 2154
rect 11642 2032 11678 2088
rect 11734 2032 11770 2088
rect 11642 1965 11770 2032
rect 11642 1909 11678 1965
rect 11734 1909 11770 1965
rect 11642 1842 11770 1909
rect 11642 1786 11678 1842
rect 11734 1786 11770 1842
rect 11642 1777 11770 1786
rect 12636 1795 12836 1796
tri 10263 1723 10283 1743 ne
rect 10283 1723 10376 1743
tri 10283 1671 10335 1723 ne
rect 10335 1671 10376 1723
tri 10335 1651 10355 1671 ne
rect 10355 1651 10376 1671
tri 10355 1630 10376 1651 ne
rect 12636 1743 12642 1795
rect 12694 1743 12710 1795
rect 12762 1743 12778 1795
rect 12830 1743 12836 1795
rect 12636 1723 12836 1743
rect 12636 1671 12642 1723
rect 12694 1671 12710 1723
rect 12762 1671 12778 1723
rect 12830 1671 12836 1723
rect 12636 1651 12836 1671
rect 12636 1599 12642 1651
rect 12694 1599 12710 1651
rect 12762 1599 12778 1651
rect 12830 1599 12836 1651
rect 10768 1455 11100 1507
rect 10768 1428 10827 1455
tri 10827 1428 10854 1455 nw
tri 11014 1428 11041 1455 ne
rect 11041 1428 11100 1455
rect 6829 1212 9737 1218
rect 6829 1190 9685 1212
tri 9651 1160 9681 1190 ne
rect 9681 1160 9685 1190
tri 9681 1158 9683 1160 ne
rect 9683 1158 9737 1160
rect 6885 1134 9605 1158
tri 9683 1156 9685 1158 ne
rect 6885 1082 6891 1134
rect 6943 1082 6956 1134
rect 7008 1082 9482 1134
rect 9534 1082 9547 1134
rect 9599 1082 9605 1134
rect 6347 1056 6399 1062
rect 6347 992 6399 1004
rect 6347 459 6399 940
rect 6347 395 6399 407
rect 6347 337 6399 343
rect 6547 1056 6599 1062
rect 6885 1058 9605 1082
rect 9685 1136 9737 1158
tri 9683 1062 9685 1064 se
rect 9685 1062 9737 1084
tri 9681 1060 9683 1062 se
rect 9683 1060 9737 1062
tri 9679 1058 9681 1060 se
rect 9681 1058 9685 1060
tri 7463 1030 7491 1058 ne
rect 7491 1030 7631 1058
tri 7631 1030 7659 1058 nw
tri 9651 1030 9679 1058 se
rect 9679 1030 9685 1058
rect 6547 992 6599 1004
rect 6829 1024 7445 1030
tri 7491 1024 7497 1030 ne
rect 6829 1002 7393 1024
tri 7359 972 7389 1002 ne
rect 7389 972 7393 1002
tri 7389 970 7391 972 ne
rect 7391 970 7445 972
tri 7391 968 7393 970 ne
rect 6547 459 6599 940
rect 7393 928 7445 970
rect 6547 395 6599 407
rect 6547 337 6599 343
rect 7224 601 7276 607
rect 7224 537 7276 549
tri 6244 320 6255 331 sw
tri 7213 320 7224 331 se
rect 7224 320 7276 485
tri 4585 287 4618 320 ne
rect 4618 297 4659 320
tri 4659 297 4682 320 sw
tri 4768 297 4791 320 ne
rect 4791 297 4842 320
tri 4842 297 4865 320 sw
tri 6158 297 6181 320 se
rect 6181 297 6255 320
tri 6255 297 6278 320 sw
tri 7190 297 7213 320 se
rect 7213 297 7276 320
rect 4618 287 4682 297
tri 4682 287 4692 297 sw
tri 4791 287 4801 297 ne
rect 4801 287 7276 297
tri 4618 274 4631 287 ne
rect 4631 274 4692 287
tri 4631 268 4637 274 ne
rect 4637 268 4692 274
tri 4692 268 4711 287 sw
tri 4801 268 4820 287 ne
rect 4820 268 7276 287
tri 4637 246 4659 268 ne
rect 4659 246 4711 268
tri 4711 246 4733 268 sw
tri 4820 246 4842 268 ne
rect 4842 246 7276 268
tri 4659 213 4692 246 ne
rect 4692 245 4733 246
tri 4733 245 4734 246 sw
tri 4842 245 4843 246 ne
rect 4843 245 7276 246
rect 4692 213 4734 245
tri 4734 213 4766 245 sw
tri 4692 161 4744 213 ne
rect 4744 161 6880 213
rect 6932 161 6944 213
rect 6996 161 7002 213
rect 1231 58 1283 70
rect 1231 0 1283 6
rect 6059 122 6111 128
rect 6059 58 6111 70
rect 6059 0 6111 6
rect 6347 122 6399 128
rect 6347 58 6399 70
rect 6347 0 6399 6
rect 6547 122 6599 128
rect 6547 58 6599 70
rect 6547 0 6599 6
rect 6745 122 6797 128
rect 6745 58 6797 70
rect 6745 0 6797 6
rect 7393 0 7445 876
rect 7497 641 7625 1030
tri 7625 1024 7631 1030 nw
rect 7497 589 7503 641
rect 7555 589 7567 641
rect 7619 589 7625 641
rect 7497 128 7625 589
rect 7497 76 7503 128
rect 7555 76 7567 128
rect 7619 76 7625 128
rect 7497 52 7625 76
rect 7497 0 7503 52
rect 7555 0 7567 52
rect 7619 0 7625 52
rect 7677 1008 9685 1030
rect 7677 1002 9737 1008
tri 9823 1002 9825 1004 se
rect 9825 1002 9923 1004
rect 7677 970 7731 1002
tri 7731 970 7763 1002 nw
tri 9791 970 9823 1002 se
rect 9823 970 9923 1002
rect 7677 0 7729 970
tri 7729 968 7731 970 nw
rect 8607 918 8613 970
rect 8665 918 8677 970
rect 8729 952 9923 970
rect 9975 952 9987 1004
rect 10039 952 10045 1004
rect 8729 936 9831 952
tri 9831 936 9847 952 nw
rect 8729 918 9813 936
tri 9813 918 9831 936 nw
rect 7835 910 8035 916
rect 7887 907 7909 910
rect 7891 858 7909 907
rect 7961 907 7983 910
rect 7961 858 7979 907
rect 7891 851 7979 858
rect 7835 803 8035 851
rect 7887 802 7909 803
rect 7891 751 7909 802
rect 7961 802 7983 803
rect 7961 751 7979 802
rect 8853 818 8859 870
rect 8911 840 8927 870
rect 8979 840 8994 870
rect 9046 840 9061 870
rect 9113 840 9128 870
rect 9180 840 9195 870
rect 8919 818 8927 840
rect 9180 818 9187 840
rect 9247 818 9262 870
rect 9314 840 9329 870
rect 9381 840 9396 870
rect 9448 840 9463 870
rect 9515 840 9530 870
rect 9582 840 9597 870
rect 9324 818 9329 840
rect 9582 818 9590 840
rect 9649 818 9655 870
rect 8853 806 8863 818
rect 8919 806 8944 818
rect 9000 806 9025 818
rect 9081 806 9106 818
rect 9162 806 9187 818
rect 9243 806 9268 818
rect 9324 806 9349 818
rect 9405 806 9430 818
rect 9486 806 9510 818
rect 9566 806 9590 818
rect 9646 806 9655 818
rect 7891 746 7979 751
rect 7835 697 8035 746
rect 7891 696 7979 697
rect 7891 644 7909 696
rect 7961 644 7979 696
rect 7891 641 7979 644
rect 7835 591 8035 641
rect 8207 757 8259 763
rect 8853 754 8859 806
rect 8919 784 8927 806
rect 9180 784 9187 806
rect 8911 754 8927 784
rect 8979 754 8994 784
rect 9046 754 9061 784
rect 9113 754 9128 784
rect 9180 754 9195 784
rect 9247 754 9262 806
rect 9324 784 9329 806
rect 9582 784 9590 806
rect 9314 754 9329 784
rect 9381 754 9396 784
rect 9448 754 9463 784
rect 9515 754 9530 784
rect 9582 754 9597 784
rect 9649 754 9655 806
rect 8207 693 8259 705
tri 8259 687 8293 721 sw
rect 8259 641 9923 687
rect 8207 635 9923 641
rect 9975 635 9987 687
rect 10039 635 10045 687
rect 7891 588 7979 591
rect 7891 536 7909 588
rect 7961 536 7979 588
rect 7891 535 7979 536
rect 7835 485 8035 535
rect 7891 480 7979 485
rect 7891 429 7909 480
rect 7887 428 7909 429
rect 7961 429 7979 480
rect 7961 428 7983 429
rect 7835 379 8035 428
rect 7891 372 7979 379
rect 7891 323 7909 372
rect 7887 320 7909 323
rect 7961 323 7979 372
rect 7961 320 7983 323
rect 7835 314 8035 320
rect 8114 555 9589 607
rect 8114 533 8178 555
tri 8178 533 8200 555 nw
tri 9567 533 9589 555 ne
tri 9589 533 9663 607 sw
tri 8113 246 8114 247 se
rect 8114 246 8166 533
tri 8166 521 8178 533 nw
tri 9589 521 9601 533 ne
rect 9601 521 9663 533
tri 9601 459 9663 521 ne
tri 9663 459 9737 533 sw
tri 9663 385 9737 459 ne
tri 9737 385 9811 459 sw
tri 9737 337 9785 385 ne
rect 9785 358 9811 385
tri 9811 358 9838 385 sw
rect 9785 337 9838 358
tri 9838 337 9859 358 sw
tri 10747 337 10768 358 se
rect 10768 337 10820 1428
tri 10820 1421 10827 1428 nw
tri 11041 1421 11048 1428 ne
tri 9785 321 9801 337 ne
rect 9801 326 9859 337
tri 9859 326 9870 337 sw
tri 10736 326 10747 337 se
rect 10747 336 10820 337
rect 10747 326 10810 336
tri 10810 326 10820 336 nw
rect 9801 321 9870 326
tri 8104 237 8113 246 se
rect 8113 237 8166 246
tri 8080 213 8104 237 se
rect 8104 213 8166 237
rect 8038 161 8044 213
rect 8096 161 8108 213
rect 8160 161 8166 213
rect 8333 320 8342 321
rect 8398 320 8424 321
rect 8480 320 8506 321
rect 8562 320 8587 321
rect 8643 320 8668 321
rect 8724 320 8733 321
rect 8333 268 8339 320
rect 8398 268 8407 320
rect 8660 268 8668 320
rect 8727 268 8733 320
tri 9801 311 9811 321 ne
rect 9811 311 9870 321
tri 9870 311 9885 326 sw
tri 10721 311 10736 326 se
rect 10736 311 10776 326
tri 9811 292 9830 311 ne
rect 9830 292 9885 311
tri 9885 292 9904 311 sw
tri 10702 292 10721 311 se
rect 10721 292 10776 311
tri 10776 292 10810 326 nw
rect 11048 292 11100 1428
tri 11994 1316 12106 1428 sw
tri 12524 1316 12636 1428 se
rect 12636 1316 12836 1599
rect 11986 1117 12836 1316
tri 11100 292 11134 326 sw
rect 8333 265 8342 268
rect 8398 265 8424 268
rect 8480 265 8506 268
rect 8562 265 8587 268
rect 8643 265 8668 268
rect 8724 265 8733 268
rect 8333 246 8733 265
tri 9830 247 9875 292 ne
rect 9875 284 9904 292
tri 9904 284 9912 292 sw
tri 10694 284 10702 292 se
rect 10702 284 10768 292
tri 10768 284 10776 292 nw
rect 9875 247 9912 284
rect 8333 194 8339 246
rect 8391 194 8407 246
rect 8459 194 8474 246
rect 8526 194 8541 246
rect 8593 194 8608 246
rect 8660 194 8675 246
rect 8727 194 8733 246
tri 9875 240 9882 247 ne
rect 9882 243 9912 247
tri 9912 243 9953 284 sw
tri 10653 243 10694 284 se
rect 10694 243 10727 284
tri 10727 243 10768 284 nw
rect 9882 240 9953 243
tri 9953 240 9956 243 sw
rect 10653 240 10724 243
tri 10724 240 10727 243 nw
rect 11048 240 12327 292
rect 12379 240 12403 292
rect 12455 240 12479 292
rect 12531 240 12555 292
rect 12607 240 12631 292
rect 12683 240 12706 292
rect 12758 240 12769 292
tri 9882 237 9885 240 ne
rect 9885 237 9956 240
tri 9956 237 9959 240 sw
rect 10653 237 10721 240
tri 10721 237 10724 240 nw
tri 9885 213 9909 237 ne
rect 9909 213 9959 237
rect 8333 175 8733 194
rect 8333 172 8342 175
rect 8398 172 8424 175
rect 8480 172 8506 175
rect 8562 172 8587 175
rect 8643 172 8668 175
rect 8724 172 8733 175
rect 8333 120 8339 172
rect 8398 120 8407 172
rect 8660 120 8668 172
rect 8727 120 8733 172
tri 9909 163 9959 213 ne
tri 9959 163 10033 237 sw
tri 9959 122 10000 163 ne
rect 10000 123 10033 163
tri 10033 123 10073 163 sw
rect 10000 122 10073 123
tri 10073 122 10074 123 sw
tri 10652 122 10653 123 se
rect 10653 122 10705 237
tri 10705 221 10721 237 nw
rect 8333 119 8342 120
rect 8398 119 8424 120
rect 8480 119 8506 120
rect 8562 119 8587 120
rect 8643 119 8668 120
rect 8724 119 8733 120
tri 10000 119 10003 122 ne
rect 10003 119 10074 122
tri 10003 89 10033 119 ne
rect 10033 89 10074 119
tri 10074 89 10107 122 sw
tri 10619 89 10652 122 se
rect 10652 89 10705 122
tri 10033 70 10052 89 ne
rect 10052 70 10705 89
tri 10052 58 10064 70 ne
rect 10064 58 10705 70
tri 10064 37 10085 58 ne
rect 10085 37 10705 58
rect 12099 122 12151 128
rect 12099 58 12151 70
rect 12099 0 12151 6
rect 13080 122 13132 3345
rect 13301 1074 13701 6861
rect 13301 1022 13307 1074
rect 13359 1022 13375 1074
rect 13427 1022 13442 1074
rect 13494 1022 13509 1074
rect 13561 1022 13576 1074
rect 13628 1022 13643 1074
rect 13695 1022 13701 1074
rect 13301 988 13701 1022
rect 13301 936 13307 988
rect 13359 936 13375 988
rect 13427 936 13442 988
rect 13494 936 13509 988
rect 13561 936 13576 988
rect 13628 936 13643 988
rect 13695 936 13701 988
rect 13301 902 13701 936
rect 13301 850 13307 902
rect 13359 850 13375 902
rect 13427 850 13442 902
rect 13494 850 13509 902
rect 13561 850 13576 902
rect 13628 850 13643 902
rect 13695 850 13701 902
rect 13301 849 13701 850
rect 13080 58 13132 70
rect 13080 0 13132 6
<< via2 >>
rect 8342 39085 8398 39141
rect 8424 39085 8480 39141
rect 8506 39085 8562 39141
rect 8587 39085 8643 39141
rect 8668 39085 8724 39141
rect 8342 38941 8398 38997
rect 8424 38941 8480 38997
rect 8506 38941 8562 38997
rect 8587 38941 8643 38997
rect 8668 38941 8724 38997
rect 7822 38829 7878 38885
rect 7904 38829 7960 38885
rect 7986 38829 8042 38885
rect 8067 38829 8123 38885
rect 8148 38829 8204 38885
rect 7822 38685 7878 38741
rect 7904 38685 7960 38741
rect 7986 38685 8042 38741
rect 8067 38685 8123 38741
rect 8148 38685 8204 38741
rect 8342 36361 8398 36417
rect 8424 36361 8480 36417
rect 8506 36361 8562 36417
rect 8587 36361 8643 36417
rect 8668 36361 8724 36417
rect 8342 36217 8398 36273
rect 8424 36217 8480 36273
rect 8506 36217 8562 36273
rect 8587 36217 8643 36273
rect 8668 36217 8724 36273
rect 7822 36105 7878 36161
rect 7904 36105 7960 36161
rect 7986 36105 8042 36161
rect 8067 36105 8123 36161
rect 8148 36105 8204 36161
rect 7822 35961 7878 36017
rect 7904 35961 7960 36017
rect 7986 35961 8042 36017
rect 8067 35961 8123 36017
rect 8148 35961 8204 36017
rect 8342 34253 8398 34309
rect 8424 34253 8480 34309
rect 8506 34253 8562 34309
rect 8587 34253 8643 34309
rect 8668 34253 8724 34309
rect 8342 34109 8398 34165
rect 8424 34109 8480 34165
rect 8506 34109 8562 34165
rect 8587 34109 8643 34165
rect 8668 34109 8724 34165
rect 7822 33997 7878 34053
rect 7904 33997 7960 34053
rect 7986 33997 8042 34053
rect 8067 33997 8123 34053
rect 8148 33997 8204 34053
rect 7822 33853 7878 33909
rect 7904 33853 7960 33909
rect 7986 33853 8042 33909
rect 8067 33853 8123 33909
rect 8148 33853 8204 33909
rect 8342 31529 8398 31585
rect 8424 31529 8480 31585
rect 8506 31529 8562 31585
rect 8587 31529 8643 31585
rect 8668 31529 8724 31585
rect 8342 31385 8398 31441
rect 8424 31385 8480 31441
rect 8506 31385 8562 31441
rect 8587 31385 8643 31441
rect 8668 31385 8724 31441
rect 7822 31273 7878 31329
rect 7904 31273 7960 31329
rect 7986 31273 8042 31329
rect 8067 31273 8123 31329
rect 8148 31273 8204 31329
rect 7822 31129 7878 31185
rect 7904 31129 7960 31185
rect 7986 31129 8042 31185
rect 8067 31129 8123 31185
rect 8148 31129 8204 31185
rect 8342 29421 8398 29477
rect 8424 29421 8480 29477
rect 8506 29421 8562 29477
rect 8587 29421 8643 29477
rect 8668 29421 8724 29477
rect 8342 29277 8398 29333
rect 8424 29277 8480 29333
rect 8506 29277 8562 29333
rect 8587 29277 8643 29333
rect 8668 29277 8724 29333
rect 7822 29165 7878 29221
rect 7904 29165 7960 29221
rect 7986 29165 8042 29221
rect 8067 29165 8123 29221
rect 8148 29165 8204 29221
rect 7822 29021 7878 29077
rect 7904 29021 7960 29077
rect 7986 29021 8042 29077
rect 8067 29021 8123 29077
rect 8148 29021 8204 29077
rect 8342 26697 8398 26753
rect 8424 26697 8480 26753
rect 8506 26697 8562 26753
rect 8587 26697 8643 26753
rect 8668 26697 8724 26753
rect 8342 26553 8398 26609
rect 8424 26553 8480 26609
rect 8506 26553 8562 26609
rect 8587 26553 8643 26609
rect 8668 26553 8724 26609
rect 7822 26441 7878 26497
rect 7904 26441 7960 26497
rect 7986 26441 8042 26497
rect 8067 26441 8123 26497
rect 8148 26441 8204 26497
rect 7822 26297 7878 26353
rect 7904 26297 7960 26353
rect 7986 26297 8042 26353
rect 8067 26297 8123 26353
rect 8148 26297 8204 26353
rect 8342 24589 8398 24645
rect 8424 24589 8480 24645
rect 8506 24589 8562 24645
rect 8587 24589 8643 24645
rect 8668 24589 8724 24645
rect 8342 24445 8398 24501
rect 8424 24445 8480 24501
rect 8506 24445 8562 24501
rect 8587 24445 8643 24501
rect 8668 24445 8724 24501
rect 7822 24333 7878 24389
rect 7904 24333 7960 24389
rect 7986 24333 8042 24389
rect 8067 24333 8123 24389
rect 8148 24333 8204 24389
rect 7822 24189 7878 24245
rect 7904 24189 7960 24245
rect 7986 24189 8042 24245
rect 8067 24189 8123 24245
rect 8148 24189 8204 24245
rect 8342 21865 8398 21921
rect 8424 21865 8480 21921
rect 8506 21865 8562 21921
rect 8587 21865 8643 21921
rect 8668 21865 8724 21921
rect 8342 21721 8398 21777
rect 8424 21721 8480 21777
rect 8506 21721 8562 21777
rect 8587 21721 8643 21777
rect 8668 21721 8724 21777
rect 7822 21609 7878 21665
rect 7904 21609 7960 21665
rect 7986 21609 8042 21665
rect 8067 21609 8123 21665
rect 8148 21609 8204 21665
rect 7822 21465 7878 21521
rect 7904 21465 7960 21521
rect 7986 21465 8042 21521
rect 8067 21465 8123 21521
rect 8148 21465 8204 21521
rect 8342 19757 8398 19813
rect 8424 19757 8480 19813
rect 8506 19757 8562 19813
rect 8587 19757 8643 19813
rect 8668 19757 8724 19813
rect 8342 19613 8398 19669
rect 8424 19613 8480 19669
rect 8506 19613 8562 19669
rect 8587 19613 8643 19669
rect 8668 19613 8724 19669
rect 7822 19501 7878 19557
rect 7904 19501 7960 19557
rect 7986 19501 8042 19557
rect 8067 19501 8123 19557
rect 8148 19501 8204 19557
rect 7822 19357 7878 19413
rect 7904 19357 7960 19413
rect 7986 19357 8042 19413
rect 8067 19357 8123 19413
rect 8148 19357 8204 19413
rect 8342 17033 8398 17089
rect 8424 17033 8480 17089
rect 8506 17033 8562 17089
rect 8587 17033 8643 17089
rect 8668 17033 8724 17089
rect 8342 16889 8398 16945
rect 8424 16889 8480 16945
rect 8506 16889 8562 16945
rect 8587 16889 8643 16945
rect 8668 16889 8724 16945
rect 7822 16777 7878 16833
rect 7904 16777 7960 16833
rect 7986 16777 8042 16833
rect 8067 16777 8123 16833
rect 8148 16777 8204 16833
rect 7822 16633 7878 16689
rect 7904 16633 7960 16689
rect 7986 16633 8042 16689
rect 8067 16633 8123 16689
rect 8148 16633 8204 16689
rect 8342 14925 8398 14981
rect 8424 14925 8480 14981
rect 8506 14925 8562 14981
rect 8587 14925 8643 14981
rect 8668 14925 8724 14981
rect 8342 14781 8398 14837
rect 8424 14781 8480 14837
rect 8506 14781 8562 14837
rect 8587 14781 8643 14837
rect 8668 14781 8724 14837
rect 7822 14669 7878 14725
rect 7904 14669 7960 14725
rect 7986 14669 8042 14725
rect 8067 14669 8123 14725
rect 8148 14669 8204 14725
rect 7822 14525 7878 14581
rect 7904 14525 7960 14581
rect 7986 14525 8042 14581
rect 8067 14525 8123 14581
rect 8148 14525 8204 14581
rect 8342 12201 8398 12257
rect 8424 12201 8480 12257
rect 8506 12201 8562 12257
rect 8587 12201 8643 12257
rect 8668 12201 8724 12257
rect 8342 12057 8398 12113
rect 8424 12057 8480 12113
rect 8506 12057 8562 12113
rect 8587 12057 8643 12113
rect 8668 12057 8724 12113
rect 7822 11945 7878 12001
rect 7904 11945 7960 12001
rect 7986 11945 8042 12001
rect 8067 11945 8123 12001
rect 8148 11945 8204 12001
rect 7822 11801 7878 11857
rect 7904 11801 7960 11857
rect 7986 11801 8042 11857
rect 8067 11801 8123 11857
rect 8148 11801 8204 11857
rect 8342 10093 8398 10149
rect 8424 10093 8480 10149
rect 8506 10093 8562 10149
rect 8587 10093 8643 10149
rect 8668 10093 8724 10149
rect 8342 9949 8398 10005
rect 8424 9949 8480 10005
rect 8506 9949 8562 10005
rect 8587 9949 8643 10005
rect 8668 9949 8724 10005
rect 7822 9837 7878 9893
rect 7904 9837 7960 9893
rect 7986 9837 8042 9893
rect 8067 9837 8123 9893
rect 8148 9837 8204 9893
rect 7822 9693 7878 9749
rect 7904 9693 7960 9749
rect 7986 9693 8042 9749
rect 8067 9693 8123 9749
rect 8148 9693 8204 9749
rect 7823 7673 7879 7729
rect 7932 7673 7988 7729
rect 8040 7673 8096 7729
rect 8148 7673 8204 7729
rect 8342 7369 8398 7425
rect 8424 7369 8480 7425
rect 8506 7369 8562 7425
rect 8587 7369 8643 7425
rect 8668 7369 8724 7425
rect 8342 7225 8398 7281
rect 8424 7225 8480 7281
rect 8506 7225 8562 7281
rect 8587 7225 8643 7281
rect 8668 7225 8724 7281
rect 7822 7113 7878 7169
rect 7904 7113 7960 7169
rect 7986 7113 8042 7169
rect 8067 7113 8123 7169
rect 8148 7113 8204 7169
rect 7822 6969 7878 7025
rect 7904 6969 7960 7025
rect 7986 6969 8042 7025
rect 8067 6969 8123 7025
rect 8148 6969 8204 7025
rect 548 2642 604 2698
rect 662 2642 718 2698
rect 776 2642 832 2698
rect 890 2642 946 2698
rect 548 2520 604 2576
rect 662 2520 718 2576
rect 776 2520 832 2576
rect 890 2520 946 2576
rect 548 2398 604 2454
rect 662 2398 718 2454
rect 776 2398 832 2454
rect 890 2398 946 2454
rect 548 2276 604 2332
rect 662 2276 718 2332
rect 776 2276 832 2332
rect 890 2276 946 2332
rect 548 2197 604 2210
rect 662 2197 718 2210
rect 776 2197 832 2210
rect 890 2197 946 2210
rect 548 2154 553 2197
rect 553 2154 604 2197
rect 662 2154 673 2197
rect 673 2154 688 2197
rect 688 2154 718 2197
rect 776 2154 807 2197
rect 807 2154 822 2197
rect 822 2154 832 2197
rect 890 2154 941 2197
rect 941 2154 946 2197
rect 548 2071 553 2088
rect 553 2071 604 2088
rect 662 2071 673 2088
rect 673 2071 688 2088
rect 688 2071 718 2088
rect 776 2071 807 2088
rect 807 2071 822 2088
rect 822 2071 832 2088
rect 890 2071 941 2088
rect 941 2071 946 2088
rect 548 2032 604 2071
rect 662 2032 718 2071
rect 776 2032 832 2071
rect 890 2032 946 2071
rect 548 1962 553 1965
rect 553 1962 604 1965
rect 662 1962 673 1965
rect 673 1962 688 1965
rect 688 1962 718 1965
rect 776 1962 807 1965
rect 807 1962 822 1965
rect 822 1962 832 1965
rect 890 1962 941 1965
rect 941 1962 946 1965
rect 548 1940 604 1962
rect 662 1940 718 1962
rect 776 1940 832 1962
rect 890 1940 946 1962
rect 548 1909 553 1940
rect 553 1909 604 1940
rect 662 1909 673 1940
rect 673 1909 688 1940
rect 688 1909 718 1940
rect 776 1909 807 1940
rect 807 1909 822 1940
rect 822 1909 832 1940
rect 890 1909 941 1940
rect 941 1909 946 1940
rect 548 1814 553 1842
rect 553 1814 604 1842
rect 662 1814 673 1842
rect 673 1814 688 1842
rect 688 1814 718 1842
rect 776 1814 807 1842
rect 807 1814 822 1842
rect 822 1814 832 1842
rect 890 1814 941 1842
rect 941 1814 946 1842
rect 548 1786 604 1814
rect 662 1786 718 1814
rect 776 1786 832 1814
rect 890 1786 946 1814
rect 11678 2642 11734 2698
rect 8342 2537 8398 2593
rect 8424 2537 8480 2593
rect 8506 2537 8562 2593
rect 8587 2537 8643 2593
rect 8668 2537 8724 2593
rect 8342 2393 8398 2449
rect 8424 2393 8480 2449
rect 8506 2393 8562 2449
rect 8587 2393 8643 2449
rect 8668 2393 8724 2449
rect 7822 2281 7878 2337
rect 7904 2281 7960 2337
rect 7986 2281 8042 2337
rect 8067 2281 8123 2337
rect 8148 2281 8204 2337
rect 7822 2137 7878 2193
rect 7904 2137 7960 2193
rect 7986 2137 8042 2193
rect 8067 2137 8123 2193
rect 8148 2137 8204 2193
rect 11678 2520 11734 2576
rect 11678 2398 11734 2454
rect 11678 2276 11734 2332
rect 11678 2154 11734 2210
rect 11678 2032 11734 2088
rect 11678 1909 11734 1965
rect 11678 1786 11734 1842
rect 7835 858 7887 907
rect 7887 858 7891 907
rect 7979 858 7983 907
rect 7983 858 8035 907
rect 7835 851 7891 858
rect 7979 851 8035 858
rect 7835 751 7887 802
rect 7887 751 7891 802
rect 7979 751 7983 802
rect 7983 751 8035 802
rect 8863 818 8911 840
rect 8911 818 8919 840
rect 8944 818 8979 840
rect 8979 818 8994 840
rect 8994 818 9000 840
rect 9025 818 9046 840
rect 9046 818 9061 840
rect 9061 818 9081 840
rect 9106 818 9113 840
rect 9113 818 9128 840
rect 9128 818 9162 840
rect 9187 818 9195 840
rect 9195 818 9243 840
rect 9268 818 9314 840
rect 9314 818 9324 840
rect 9349 818 9381 840
rect 9381 818 9396 840
rect 9396 818 9405 840
rect 9430 818 9448 840
rect 9448 818 9463 840
rect 9463 818 9486 840
rect 9510 818 9515 840
rect 9515 818 9530 840
rect 9530 818 9566 840
rect 9590 818 9597 840
rect 9597 818 9646 840
rect 8863 806 8919 818
rect 8944 806 9000 818
rect 9025 806 9081 818
rect 9106 806 9162 818
rect 9187 806 9243 818
rect 9268 806 9324 818
rect 9349 806 9405 818
rect 9430 806 9486 818
rect 9510 806 9566 818
rect 9590 806 9646 818
rect 7835 746 7891 751
rect 7979 746 8035 751
rect 7835 696 7891 697
rect 7979 696 8035 697
rect 7835 644 7887 696
rect 7887 644 7891 696
rect 7979 644 7983 696
rect 7983 644 8035 696
rect 7835 641 7891 644
rect 7979 641 8035 644
rect 8863 784 8911 806
rect 8911 784 8919 806
rect 8944 784 8979 806
rect 8979 784 8994 806
rect 8994 784 9000 806
rect 9025 784 9046 806
rect 9046 784 9061 806
rect 9061 784 9081 806
rect 9106 784 9113 806
rect 9113 784 9128 806
rect 9128 784 9162 806
rect 9187 784 9195 806
rect 9195 784 9243 806
rect 9268 784 9314 806
rect 9314 784 9324 806
rect 9349 784 9381 806
rect 9381 784 9396 806
rect 9396 784 9405 806
rect 9430 784 9448 806
rect 9448 784 9463 806
rect 9463 784 9486 806
rect 9510 784 9515 806
rect 9515 784 9530 806
rect 9530 784 9566 806
rect 9590 784 9597 806
rect 9597 784 9646 806
rect 7835 588 7891 591
rect 7979 588 8035 591
rect 7835 536 7887 588
rect 7887 536 7891 588
rect 7979 536 7983 588
rect 7983 536 8035 588
rect 7835 535 7891 536
rect 7979 535 8035 536
rect 7835 480 7891 485
rect 7979 480 8035 485
rect 7835 429 7887 480
rect 7887 429 7891 480
rect 7979 429 7983 480
rect 7983 429 8035 480
rect 7835 372 7891 379
rect 7979 372 8035 379
rect 7835 323 7887 372
rect 7887 323 7891 372
rect 7979 323 7983 372
rect 7983 323 8035 372
rect 8342 320 8398 321
rect 8424 320 8480 321
rect 8506 320 8562 321
rect 8587 320 8643 321
rect 8668 320 8724 321
rect 8342 268 8391 320
rect 8391 268 8398 320
rect 8424 268 8459 320
rect 8459 268 8474 320
rect 8474 268 8480 320
rect 8506 268 8526 320
rect 8526 268 8541 320
rect 8541 268 8562 320
rect 8587 268 8593 320
rect 8593 268 8608 320
rect 8608 268 8643 320
rect 8668 268 8675 320
rect 8675 268 8724 320
rect 8342 265 8398 268
rect 8424 265 8480 268
rect 8506 265 8562 268
rect 8587 265 8643 268
rect 8668 265 8724 268
rect 8342 172 8398 175
rect 8424 172 8480 175
rect 8506 172 8562 175
rect 8587 172 8643 175
rect 8668 172 8724 175
rect 8342 120 8391 172
rect 8391 120 8398 172
rect 8424 120 8459 172
rect 8459 120 8474 172
rect 8474 120 8480 172
rect 8506 120 8526 172
rect 8526 120 8541 172
rect 8541 120 8562 172
rect 8587 120 8593 172
rect 8593 120 8608 172
rect 8608 120 8643 172
rect 8668 120 8675 172
rect 8675 120 8724 172
rect 8342 119 8398 120
rect 8424 119 8480 120
rect 8506 119 8562 120
rect 8587 119 8643 120
rect 8668 119 8724 120
<< metal3 >>
rect 391 9244 2433 40000
rect 391 9180 397 9244
rect 461 9180 479 9244
rect 543 9180 561 9244
rect 625 9180 643 9244
rect 707 9180 725 9244
rect 789 9180 807 9244
rect 871 9180 889 9244
rect 953 9180 971 9244
rect 1035 9180 1053 9244
rect 1117 9180 1135 9244
rect 1199 9180 1217 9244
rect 1281 9180 1299 9244
rect 1363 9180 1381 9244
rect 1445 9180 1463 9244
rect 1527 9180 1545 9244
rect 1609 9180 1627 9244
rect 1691 9180 1709 9244
rect 1773 9180 1791 9244
rect 1855 9180 1873 9244
rect 1937 9180 1955 9244
rect 2019 9180 2037 9244
rect 2101 9180 2119 9244
rect 2183 9180 2201 9244
rect 2265 9180 2282 9244
rect 2346 9180 2363 9244
rect 2427 9180 2433 9244
rect 391 9158 2433 9180
rect 391 9094 397 9158
rect 461 9094 479 9158
rect 543 9094 561 9158
rect 625 9094 643 9158
rect 707 9094 725 9158
rect 789 9094 807 9158
rect 871 9094 889 9158
rect 953 9094 971 9158
rect 1035 9094 1053 9158
rect 1117 9094 1135 9158
rect 1199 9094 1217 9158
rect 1281 9094 1299 9158
rect 1363 9094 1381 9158
rect 1445 9094 1463 9158
rect 1527 9094 1545 9158
rect 1609 9094 1627 9158
rect 1691 9094 1709 9158
rect 1773 9094 1791 9158
rect 1855 9094 1873 9158
rect 1937 9094 1955 9158
rect 2019 9094 2037 9158
rect 2101 9094 2119 9158
rect 2183 9094 2201 9158
rect 2265 9094 2282 9158
rect 2346 9094 2363 9158
rect 2427 9094 2433 9158
rect 391 9072 2433 9094
rect 391 9008 397 9072
rect 461 9008 479 9072
rect 543 9008 561 9072
rect 625 9008 643 9072
rect 707 9008 725 9072
rect 789 9008 807 9072
rect 871 9008 889 9072
rect 953 9008 971 9072
rect 1035 9008 1053 9072
rect 1117 9008 1135 9072
rect 1199 9008 1217 9072
rect 1281 9008 1299 9072
rect 1363 9008 1381 9072
rect 1445 9008 1463 9072
rect 1527 9008 1545 9072
rect 1609 9008 1627 9072
rect 1691 9008 1709 9072
rect 1773 9008 1791 9072
rect 1855 9008 1873 9072
rect 1937 9008 1955 9072
rect 2019 9008 2037 9072
rect 2101 9008 2119 9072
rect 2183 9008 2201 9072
rect 2265 9008 2282 9072
rect 2346 9008 2363 9072
rect 2427 9008 2433 9072
rect 391 8986 2433 9008
rect 391 8922 397 8986
rect 461 8922 479 8986
rect 543 8922 561 8986
rect 625 8922 643 8986
rect 707 8922 725 8986
rect 789 8922 807 8986
rect 871 8922 889 8986
rect 953 8922 971 8986
rect 1035 8922 1053 8986
rect 1117 8922 1135 8986
rect 1199 8922 1217 8986
rect 1281 8922 1299 8986
rect 1363 8922 1381 8986
rect 1445 8922 1463 8986
rect 1527 8922 1545 8986
rect 1609 8922 1627 8986
rect 1691 8922 1709 8986
rect 1773 8922 1791 8986
rect 1855 8922 1873 8986
rect 1937 8922 1955 8986
rect 2019 8922 2037 8986
rect 2101 8922 2119 8986
rect 2183 8922 2201 8986
rect 2265 8922 2282 8986
rect 2346 8922 2363 8986
rect 2427 8922 2433 8986
rect 391 8900 2433 8922
rect 391 8836 397 8900
rect 461 8836 479 8900
rect 543 8836 561 8900
rect 625 8836 643 8900
rect 707 8836 725 8900
rect 789 8836 807 8900
rect 871 8836 889 8900
rect 953 8836 971 8900
rect 1035 8836 1053 8900
rect 1117 8836 1135 8900
rect 1199 8836 1217 8900
rect 1281 8836 1299 8900
rect 1363 8836 1381 8900
rect 1445 8836 1463 8900
rect 1527 8836 1545 8900
rect 1609 8836 1627 8900
rect 1691 8836 1709 8900
rect 1773 8836 1791 8900
rect 1855 8836 1873 8900
rect 1937 8836 1955 8900
rect 2019 8836 2037 8900
rect 2101 8836 2119 8900
rect 2183 8836 2201 8900
rect 2265 8836 2282 8900
rect 2346 8836 2363 8900
rect 2427 8836 2433 8900
rect 391 8814 2433 8836
rect 391 8750 397 8814
rect 461 8750 479 8814
rect 543 8750 561 8814
rect 625 8750 643 8814
rect 707 8750 725 8814
rect 789 8750 807 8814
rect 871 8750 889 8814
rect 953 8750 971 8814
rect 1035 8750 1053 8814
rect 1117 8750 1135 8814
rect 1199 8750 1217 8814
rect 1281 8750 1299 8814
rect 1363 8750 1381 8814
rect 1445 8750 1463 8814
rect 1527 8750 1545 8814
rect 1609 8750 1627 8814
rect 1691 8750 1709 8814
rect 1773 8750 1791 8814
rect 1855 8750 1873 8814
rect 1937 8750 1955 8814
rect 2019 8750 2037 8814
rect 2101 8750 2119 8814
rect 2183 8750 2201 8814
rect 2265 8750 2282 8814
rect 2346 8750 2363 8814
rect 2427 8750 2433 8814
rect 391 8728 2433 8750
rect 391 8664 397 8728
rect 461 8664 479 8728
rect 543 8664 561 8728
rect 625 8664 643 8728
rect 707 8664 725 8728
rect 789 8664 807 8728
rect 871 8664 889 8728
rect 953 8664 971 8728
rect 1035 8664 1053 8728
rect 1117 8664 1135 8728
rect 1199 8664 1217 8728
rect 1281 8664 1299 8728
rect 1363 8664 1381 8728
rect 1445 8664 1463 8728
rect 1527 8664 1545 8728
rect 1609 8664 1627 8728
rect 1691 8664 1709 8728
rect 1773 8664 1791 8728
rect 1855 8664 1873 8728
rect 1937 8664 1955 8728
rect 2019 8664 2037 8728
rect 2101 8664 2119 8728
rect 2183 8664 2201 8728
rect 2265 8664 2282 8728
rect 2346 8664 2363 8728
rect 2427 8664 2433 8728
rect 391 8642 2433 8664
rect 391 8578 397 8642
rect 461 8578 479 8642
rect 543 8578 561 8642
rect 625 8578 643 8642
rect 707 8578 725 8642
rect 789 8578 807 8642
rect 871 8578 889 8642
rect 953 8578 971 8642
rect 1035 8578 1053 8642
rect 1117 8578 1135 8642
rect 1199 8578 1217 8642
rect 1281 8578 1299 8642
rect 1363 8578 1381 8642
rect 1445 8578 1463 8642
rect 1527 8578 1545 8642
rect 1609 8578 1627 8642
rect 1691 8578 1709 8642
rect 1773 8578 1791 8642
rect 1855 8578 1873 8642
rect 1937 8578 1955 8642
rect 2019 8578 2037 8642
rect 2101 8578 2119 8642
rect 2183 8578 2201 8642
rect 2265 8578 2282 8642
rect 2346 8578 2363 8642
rect 2427 8578 2433 8642
rect 391 8556 2433 8578
rect 391 8492 397 8556
rect 461 8492 479 8556
rect 543 8492 561 8556
rect 625 8492 643 8556
rect 707 8492 725 8556
rect 789 8492 807 8556
rect 871 8492 889 8556
rect 953 8492 971 8556
rect 1035 8492 1053 8556
rect 1117 8492 1135 8556
rect 1199 8492 1217 8556
rect 1281 8492 1299 8556
rect 1363 8492 1381 8556
rect 1445 8492 1463 8556
rect 1527 8492 1545 8556
rect 1609 8492 1627 8556
rect 1691 8492 1709 8556
rect 1773 8492 1791 8556
rect 1855 8492 1873 8556
rect 1937 8492 1955 8556
rect 2019 8492 2037 8556
rect 2101 8492 2119 8556
rect 2183 8492 2201 8556
rect 2265 8492 2282 8556
rect 2346 8492 2363 8556
rect 2427 8492 2433 8556
rect 391 8470 2433 8492
rect 391 8406 397 8470
rect 461 8406 479 8470
rect 543 8406 561 8470
rect 625 8406 643 8470
rect 707 8406 725 8470
rect 789 8406 807 8470
rect 871 8406 889 8470
rect 953 8406 971 8470
rect 1035 8406 1053 8470
rect 1117 8406 1135 8470
rect 1199 8406 1217 8470
rect 1281 8406 1299 8470
rect 1363 8406 1381 8470
rect 1445 8406 1463 8470
rect 1527 8406 1545 8470
rect 1609 8406 1627 8470
rect 1691 8406 1709 8470
rect 1773 8406 1791 8470
rect 1855 8406 1873 8470
rect 1937 8406 1955 8470
rect 2019 8406 2037 8470
rect 2101 8406 2119 8470
rect 2183 8406 2201 8470
rect 2265 8406 2282 8470
rect 2346 8406 2363 8470
rect 2427 8406 2433 8470
rect 391 8384 2433 8406
rect 391 8320 397 8384
rect 461 8320 479 8384
rect 543 8320 561 8384
rect 625 8320 643 8384
rect 707 8320 725 8384
rect 789 8320 807 8384
rect 871 8320 889 8384
rect 953 8320 971 8384
rect 1035 8320 1053 8384
rect 1117 8320 1135 8384
rect 1199 8320 1217 8384
rect 1281 8320 1299 8384
rect 1363 8320 1381 8384
rect 1445 8320 1463 8384
rect 1527 8320 1545 8384
rect 1609 8320 1627 8384
rect 1691 8320 1709 8384
rect 1773 8320 1791 8384
rect 1855 8320 1873 8384
rect 1937 8320 1955 8384
rect 2019 8320 2037 8384
rect 2101 8320 2119 8384
rect 2183 8320 2201 8384
rect 2265 8320 2282 8384
rect 2346 8320 2363 8384
rect 2427 8320 2433 8384
rect 391 2962 2433 8320
tri 1322 2707 1577 2962 ne
rect 1577 2707 2433 2962
rect 542 2701 952 2707
rect 542 2637 547 2701
rect 611 2637 659 2701
rect 723 2637 771 2701
rect 835 2637 883 2701
rect 947 2637 952 2701
tri 1577 2698 1586 2707 ne
rect 1586 2698 2433 2707
tri 1586 2651 1633 2698 ne
rect 542 2579 952 2637
rect 542 2515 547 2579
rect 611 2515 659 2579
rect 723 2515 771 2579
rect 835 2515 883 2579
rect 947 2515 952 2579
rect 542 2457 952 2515
rect 542 2393 547 2457
rect 611 2393 659 2457
rect 723 2393 771 2457
rect 835 2393 883 2457
rect 947 2393 952 2457
rect 542 2335 952 2393
rect 542 2271 547 2335
rect 611 2271 659 2335
rect 723 2271 771 2335
rect 835 2271 883 2335
rect 947 2271 952 2335
rect 542 2213 952 2271
rect 542 2149 547 2213
rect 611 2149 659 2213
rect 723 2149 771 2213
rect 835 2149 883 2213
rect 947 2149 952 2213
rect 542 2091 952 2149
rect 542 2027 547 2091
rect 611 2027 659 2091
rect 723 2027 771 2091
rect 835 2027 883 2091
rect 947 2027 952 2091
rect 542 1969 952 2027
rect 542 1905 547 1969
rect 611 1905 659 1969
rect 723 1905 771 1969
rect 835 1905 883 1969
rect 947 1905 952 1969
rect 542 1847 952 1905
rect 542 1783 547 1847
rect 611 1783 659 1847
rect 723 1783 771 1847
rect 835 1783 883 1847
rect 947 1783 952 1847
rect 542 1777 952 1783
rect 1633 0 2433 2698
rect 2547 9244 4575 40000
rect 2547 9180 2553 9244
rect 2617 9180 2635 9244
rect 2699 9180 2717 9244
rect 2781 9180 2799 9244
rect 2863 9180 2881 9244
rect 2945 9180 2963 9244
rect 3027 9180 3045 9244
rect 3109 9180 3127 9244
rect 3191 9180 3209 9244
rect 3273 9180 3290 9244
rect 3354 9180 3371 9244
rect 3435 9180 3452 9244
rect 3516 9180 3533 9244
rect 3597 9180 3614 9244
rect 3678 9180 3695 9244
rect 3759 9180 3776 9244
rect 3840 9180 3857 9244
rect 3921 9180 3938 9244
rect 4002 9180 4019 9244
rect 4083 9180 4100 9244
rect 4164 9180 4181 9244
rect 4245 9180 4262 9244
rect 4326 9180 4343 9244
rect 4407 9180 4424 9244
rect 4488 9180 4505 9244
rect 4569 9180 4575 9244
rect 2547 9158 4575 9180
rect 2547 9094 2553 9158
rect 2617 9094 2635 9158
rect 2699 9094 2717 9158
rect 2781 9094 2799 9158
rect 2863 9094 2881 9158
rect 2945 9094 2963 9158
rect 3027 9094 3045 9158
rect 3109 9094 3127 9158
rect 3191 9094 3209 9158
rect 3273 9094 3290 9158
rect 3354 9094 3371 9158
rect 3435 9094 3452 9158
rect 3516 9094 3533 9158
rect 3597 9094 3614 9158
rect 3678 9094 3695 9158
rect 3759 9094 3776 9158
rect 3840 9094 3857 9158
rect 3921 9094 3938 9158
rect 4002 9094 4019 9158
rect 4083 9094 4100 9158
rect 4164 9094 4181 9158
rect 4245 9094 4262 9158
rect 4326 9094 4343 9158
rect 4407 9094 4424 9158
rect 4488 9094 4505 9158
rect 4569 9094 4575 9158
rect 2547 9072 4575 9094
rect 2547 9008 2553 9072
rect 2617 9008 2635 9072
rect 2699 9008 2717 9072
rect 2781 9008 2799 9072
rect 2863 9008 2881 9072
rect 2945 9008 2963 9072
rect 3027 9008 3045 9072
rect 3109 9008 3127 9072
rect 3191 9008 3209 9072
rect 3273 9008 3290 9072
rect 3354 9008 3371 9072
rect 3435 9008 3452 9072
rect 3516 9008 3533 9072
rect 3597 9008 3614 9072
rect 3678 9008 3695 9072
rect 3759 9008 3776 9072
rect 3840 9008 3857 9072
rect 3921 9008 3938 9072
rect 4002 9008 4019 9072
rect 4083 9008 4100 9072
rect 4164 9008 4181 9072
rect 4245 9008 4262 9072
rect 4326 9008 4343 9072
rect 4407 9008 4424 9072
rect 4488 9008 4505 9072
rect 4569 9008 4575 9072
rect 2547 8986 4575 9008
rect 2547 8922 2553 8986
rect 2617 8922 2635 8986
rect 2699 8922 2717 8986
rect 2781 8922 2799 8986
rect 2863 8922 2881 8986
rect 2945 8922 2963 8986
rect 3027 8922 3045 8986
rect 3109 8922 3127 8986
rect 3191 8922 3209 8986
rect 3273 8922 3290 8986
rect 3354 8922 3371 8986
rect 3435 8922 3452 8986
rect 3516 8922 3533 8986
rect 3597 8922 3614 8986
rect 3678 8922 3695 8986
rect 3759 8922 3776 8986
rect 3840 8922 3857 8986
rect 3921 8922 3938 8986
rect 4002 8922 4019 8986
rect 4083 8922 4100 8986
rect 4164 8922 4181 8986
rect 4245 8922 4262 8986
rect 4326 8922 4343 8986
rect 4407 8922 4424 8986
rect 4488 8922 4505 8986
rect 4569 8922 4575 8986
rect 2547 8900 4575 8922
rect 2547 8836 2553 8900
rect 2617 8836 2635 8900
rect 2699 8836 2717 8900
rect 2781 8836 2799 8900
rect 2863 8836 2881 8900
rect 2945 8836 2963 8900
rect 3027 8836 3045 8900
rect 3109 8836 3127 8900
rect 3191 8836 3209 8900
rect 3273 8836 3290 8900
rect 3354 8836 3371 8900
rect 3435 8836 3452 8900
rect 3516 8836 3533 8900
rect 3597 8836 3614 8900
rect 3678 8836 3695 8900
rect 3759 8836 3776 8900
rect 3840 8836 3857 8900
rect 3921 8836 3938 8900
rect 4002 8836 4019 8900
rect 4083 8836 4100 8900
rect 4164 8836 4181 8900
rect 4245 8836 4262 8900
rect 4326 8836 4343 8900
rect 4407 8836 4424 8900
rect 4488 8836 4505 8900
rect 4569 8836 4575 8900
rect 2547 8814 4575 8836
rect 2547 8750 2553 8814
rect 2617 8750 2635 8814
rect 2699 8750 2717 8814
rect 2781 8750 2799 8814
rect 2863 8750 2881 8814
rect 2945 8750 2963 8814
rect 3027 8750 3045 8814
rect 3109 8750 3127 8814
rect 3191 8750 3209 8814
rect 3273 8750 3290 8814
rect 3354 8750 3371 8814
rect 3435 8750 3452 8814
rect 3516 8750 3533 8814
rect 3597 8750 3614 8814
rect 3678 8750 3695 8814
rect 3759 8750 3776 8814
rect 3840 8750 3857 8814
rect 3921 8750 3938 8814
rect 4002 8750 4019 8814
rect 4083 8750 4100 8814
rect 4164 8750 4181 8814
rect 4245 8750 4262 8814
rect 4326 8750 4343 8814
rect 4407 8750 4424 8814
rect 4488 8750 4505 8814
rect 4569 8750 4575 8814
rect 2547 8728 4575 8750
rect 2547 8664 2553 8728
rect 2617 8664 2635 8728
rect 2699 8664 2717 8728
rect 2781 8664 2799 8728
rect 2863 8664 2881 8728
rect 2945 8664 2963 8728
rect 3027 8664 3045 8728
rect 3109 8664 3127 8728
rect 3191 8664 3209 8728
rect 3273 8664 3290 8728
rect 3354 8664 3371 8728
rect 3435 8664 3452 8728
rect 3516 8664 3533 8728
rect 3597 8664 3614 8728
rect 3678 8664 3695 8728
rect 3759 8664 3776 8728
rect 3840 8664 3857 8728
rect 3921 8664 3938 8728
rect 4002 8664 4019 8728
rect 4083 8664 4100 8728
rect 4164 8664 4181 8728
rect 4245 8664 4262 8728
rect 4326 8664 4343 8728
rect 4407 8664 4424 8728
rect 4488 8664 4505 8728
rect 4569 8664 4575 8728
rect 2547 8642 4575 8664
rect 2547 8578 2553 8642
rect 2617 8578 2635 8642
rect 2699 8578 2717 8642
rect 2781 8578 2799 8642
rect 2863 8578 2881 8642
rect 2945 8578 2963 8642
rect 3027 8578 3045 8642
rect 3109 8578 3127 8642
rect 3191 8578 3209 8642
rect 3273 8578 3290 8642
rect 3354 8578 3371 8642
rect 3435 8578 3452 8642
rect 3516 8578 3533 8642
rect 3597 8578 3614 8642
rect 3678 8578 3695 8642
rect 3759 8578 3776 8642
rect 3840 8578 3857 8642
rect 3921 8578 3938 8642
rect 4002 8578 4019 8642
rect 4083 8578 4100 8642
rect 4164 8578 4181 8642
rect 4245 8578 4262 8642
rect 4326 8578 4343 8642
rect 4407 8578 4424 8642
rect 4488 8578 4505 8642
rect 4569 8578 4575 8642
rect 2547 8556 4575 8578
rect 2547 8492 2553 8556
rect 2617 8492 2635 8556
rect 2699 8492 2717 8556
rect 2781 8492 2799 8556
rect 2863 8492 2881 8556
rect 2945 8492 2963 8556
rect 3027 8492 3045 8556
rect 3109 8492 3127 8556
rect 3191 8492 3209 8556
rect 3273 8492 3290 8556
rect 3354 8492 3371 8556
rect 3435 8492 3452 8556
rect 3516 8492 3533 8556
rect 3597 8492 3614 8556
rect 3678 8492 3695 8556
rect 3759 8492 3776 8556
rect 3840 8492 3857 8556
rect 3921 8492 3938 8556
rect 4002 8492 4019 8556
rect 4083 8492 4100 8556
rect 4164 8492 4181 8556
rect 4245 8492 4262 8556
rect 4326 8492 4343 8556
rect 4407 8492 4424 8556
rect 4488 8492 4505 8556
rect 4569 8492 4575 8556
rect 2547 8470 4575 8492
rect 2547 8406 2553 8470
rect 2617 8406 2635 8470
rect 2699 8406 2717 8470
rect 2781 8406 2799 8470
rect 2863 8406 2881 8470
rect 2945 8406 2963 8470
rect 3027 8406 3045 8470
rect 3109 8406 3127 8470
rect 3191 8406 3209 8470
rect 3273 8406 3290 8470
rect 3354 8406 3371 8470
rect 3435 8406 3452 8470
rect 3516 8406 3533 8470
rect 3597 8406 3614 8470
rect 3678 8406 3695 8470
rect 3759 8406 3776 8470
rect 3840 8406 3857 8470
rect 3921 8406 3938 8470
rect 4002 8406 4019 8470
rect 4083 8406 4100 8470
rect 4164 8406 4181 8470
rect 4245 8406 4262 8470
rect 4326 8406 4343 8470
rect 4407 8406 4424 8470
rect 4488 8406 4505 8470
rect 4569 8406 4575 8470
rect 2547 8384 4575 8406
rect 2547 8320 2553 8384
rect 2617 8320 2635 8384
rect 2699 8320 2717 8384
rect 2781 8320 2799 8384
rect 2863 8320 2881 8384
rect 2945 8320 2963 8384
rect 3027 8320 3045 8384
rect 3109 8320 3127 8384
rect 3191 8320 3209 8384
rect 3273 8320 3290 8384
rect 3354 8320 3371 8384
rect 3435 8320 3452 8384
rect 3516 8320 3533 8384
rect 3597 8320 3614 8384
rect 3678 8320 3695 8384
rect 3759 8320 3776 8384
rect 3840 8320 3857 8384
rect 3921 8320 3938 8384
rect 4002 8320 4019 8384
rect 4083 8320 4100 8384
rect 4164 8320 4181 8384
rect 4245 8320 4262 8384
rect 4326 8320 4343 8384
rect 4407 8320 4424 8384
rect 4488 8320 4505 8384
rect 4569 8320 4575 8384
rect 2547 0 4575 8320
rect 4689 9244 7693 40000
rect 4689 9180 4695 9244
rect 4759 9180 4777 9244
rect 4841 9180 4859 9244
rect 4923 9180 4941 9244
rect 5005 9180 5023 9244
rect 5087 9180 5105 9244
rect 5169 9180 5187 9244
rect 5251 9180 5269 9244
rect 5333 9180 5351 9244
rect 5415 9180 5433 9244
rect 5497 9180 5515 9244
rect 5579 9180 5597 9244
rect 5661 9180 5679 9244
rect 5743 9180 5760 9244
rect 5824 9180 5841 9244
rect 5905 9180 5922 9244
rect 5986 9180 6003 9244
rect 6067 9180 6084 9244
rect 6148 9180 6165 9244
rect 6229 9180 6246 9244
rect 6310 9180 6327 9244
rect 6391 9180 6408 9244
rect 6472 9180 6489 9244
rect 6553 9180 6570 9244
rect 6634 9180 6651 9244
rect 6715 9180 6732 9244
rect 6796 9180 6813 9244
rect 6877 9180 6894 9244
rect 6958 9180 6975 9244
rect 7039 9180 7056 9244
rect 7120 9180 7137 9244
rect 7201 9180 7218 9244
rect 7282 9180 7299 9244
rect 7363 9180 7380 9244
rect 7444 9180 7461 9244
rect 7525 9180 7542 9244
rect 7606 9180 7623 9244
rect 7687 9180 7693 9244
rect 4689 9158 7693 9180
rect 4689 9094 4695 9158
rect 4759 9094 4777 9158
rect 4841 9094 4859 9158
rect 4923 9094 4941 9158
rect 5005 9094 5023 9158
rect 5087 9094 5105 9158
rect 5169 9094 5187 9158
rect 5251 9094 5269 9158
rect 5333 9094 5351 9158
rect 5415 9094 5433 9158
rect 5497 9094 5515 9158
rect 5579 9094 5597 9158
rect 5661 9094 5679 9158
rect 5743 9094 5760 9158
rect 5824 9094 5841 9158
rect 5905 9094 5922 9158
rect 5986 9094 6003 9158
rect 6067 9094 6084 9158
rect 6148 9094 6165 9158
rect 6229 9094 6246 9158
rect 6310 9094 6327 9158
rect 6391 9094 6408 9158
rect 6472 9094 6489 9158
rect 6553 9094 6570 9158
rect 6634 9094 6651 9158
rect 6715 9094 6732 9158
rect 6796 9094 6813 9158
rect 6877 9094 6894 9158
rect 6958 9094 6975 9158
rect 7039 9094 7056 9158
rect 7120 9094 7137 9158
rect 7201 9094 7218 9158
rect 7282 9094 7299 9158
rect 7363 9094 7380 9158
rect 7444 9094 7461 9158
rect 7525 9094 7542 9158
rect 7606 9094 7623 9158
rect 7687 9094 7693 9158
rect 4689 9072 7693 9094
rect 4689 9008 4695 9072
rect 4759 9008 4777 9072
rect 4841 9008 4859 9072
rect 4923 9008 4941 9072
rect 5005 9008 5023 9072
rect 5087 9008 5105 9072
rect 5169 9008 5187 9072
rect 5251 9008 5269 9072
rect 5333 9008 5351 9072
rect 5415 9008 5433 9072
rect 5497 9008 5515 9072
rect 5579 9008 5597 9072
rect 5661 9008 5679 9072
rect 5743 9008 5760 9072
rect 5824 9008 5841 9072
rect 5905 9008 5922 9072
rect 5986 9008 6003 9072
rect 6067 9008 6084 9072
rect 6148 9008 6165 9072
rect 6229 9008 6246 9072
rect 6310 9008 6327 9072
rect 6391 9008 6408 9072
rect 6472 9008 6489 9072
rect 6553 9008 6570 9072
rect 6634 9008 6651 9072
rect 6715 9008 6732 9072
rect 6796 9008 6813 9072
rect 6877 9008 6894 9072
rect 6958 9008 6975 9072
rect 7039 9008 7056 9072
rect 7120 9008 7137 9072
rect 7201 9008 7218 9072
rect 7282 9008 7299 9072
rect 7363 9008 7380 9072
rect 7444 9008 7461 9072
rect 7525 9008 7542 9072
rect 7606 9008 7623 9072
rect 7687 9008 7693 9072
rect 4689 8986 7693 9008
rect 4689 8922 4695 8986
rect 4759 8922 4777 8986
rect 4841 8922 4859 8986
rect 4923 8922 4941 8986
rect 5005 8922 5023 8986
rect 5087 8922 5105 8986
rect 5169 8922 5187 8986
rect 5251 8922 5269 8986
rect 5333 8922 5351 8986
rect 5415 8922 5433 8986
rect 5497 8922 5515 8986
rect 5579 8922 5597 8986
rect 5661 8922 5679 8986
rect 5743 8922 5760 8986
rect 5824 8922 5841 8986
rect 5905 8922 5922 8986
rect 5986 8922 6003 8986
rect 6067 8922 6084 8986
rect 6148 8922 6165 8986
rect 6229 8922 6246 8986
rect 6310 8922 6327 8986
rect 6391 8922 6408 8986
rect 6472 8922 6489 8986
rect 6553 8922 6570 8986
rect 6634 8922 6651 8986
rect 6715 8922 6732 8986
rect 6796 8922 6813 8986
rect 6877 8922 6894 8986
rect 6958 8922 6975 8986
rect 7039 8922 7056 8986
rect 7120 8922 7137 8986
rect 7201 8922 7218 8986
rect 7282 8922 7299 8986
rect 7363 8922 7380 8986
rect 7444 8922 7461 8986
rect 7525 8922 7542 8986
rect 7606 8922 7623 8986
rect 7687 8922 7693 8986
rect 4689 8900 7693 8922
rect 4689 8836 4695 8900
rect 4759 8836 4777 8900
rect 4841 8836 4859 8900
rect 4923 8836 4941 8900
rect 5005 8836 5023 8900
rect 5087 8836 5105 8900
rect 5169 8836 5187 8900
rect 5251 8836 5269 8900
rect 5333 8836 5351 8900
rect 5415 8836 5433 8900
rect 5497 8836 5515 8900
rect 5579 8836 5597 8900
rect 5661 8836 5679 8900
rect 5743 8836 5760 8900
rect 5824 8836 5841 8900
rect 5905 8836 5922 8900
rect 5986 8836 6003 8900
rect 6067 8836 6084 8900
rect 6148 8836 6165 8900
rect 6229 8836 6246 8900
rect 6310 8836 6327 8900
rect 6391 8836 6408 8900
rect 6472 8836 6489 8900
rect 6553 8836 6570 8900
rect 6634 8836 6651 8900
rect 6715 8836 6732 8900
rect 6796 8836 6813 8900
rect 6877 8836 6894 8900
rect 6958 8836 6975 8900
rect 7039 8836 7056 8900
rect 7120 8836 7137 8900
rect 7201 8836 7218 8900
rect 7282 8836 7299 8900
rect 7363 8836 7380 8900
rect 7444 8836 7461 8900
rect 7525 8836 7542 8900
rect 7606 8836 7623 8900
rect 7687 8836 7693 8900
rect 4689 8814 7693 8836
rect 4689 8750 4695 8814
rect 4759 8750 4777 8814
rect 4841 8750 4859 8814
rect 4923 8750 4941 8814
rect 5005 8750 5023 8814
rect 5087 8750 5105 8814
rect 5169 8750 5187 8814
rect 5251 8750 5269 8814
rect 5333 8750 5351 8814
rect 5415 8750 5433 8814
rect 5497 8750 5515 8814
rect 5579 8750 5597 8814
rect 5661 8750 5679 8814
rect 5743 8750 5760 8814
rect 5824 8750 5841 8814
rect 5905 8750 5922 8814
rect 5986 8750 6003 8814
rect 6067 8750 6084 8814
rect 6148 8750 6165 8814
rect 6229 8750 6246 8814
rect 6310 8750 6327 8814
rect 6391 8750 6408 8814
rect 6472 8750 6489 8814
rect 6553 8750 6570 8814
rect 6634 8750 6651 8814
rect 6715 8750 6732 8814
rect 6796 8750 6813 8814
rect 6877 8750 6894 8814
rect 6958 8750 6975 8814
rect 7039 8750 7056 8814
rect 7120 8750 7137 8814
rect 7201 8750 7218 8814
rect 7282 8750 7299 8814
rect 7363 8750 7380 8814
rect 7444 8750 7461 8814
rect 7525 8750 7542 8814
rect 7606 8750 7623 8814
rect 7687 8750 7693 8814
rect 4689 8728 7693 8750
rect 4689 8664 4695 8728
rect 4759 8664 4777 8728
rect 4841 8664 4859 8728
rect 4923 8664 4941 8728
rect 5005 8664 5023 8728
rect 5087 8664 5105 8728
rect 5169 8664 5187 8728
rect 5251 8664 5269 8728
rect 5333 8664 5351 8728
rect 5415 8664 5433 8728
rect 5497 8664 5515 8728
rect 5579 8664 5597 8728
rect 5661 8664 5679 8728
rect 5743 8664 5760 8728
rect 5824 8664 5841 8728
rect 5905 8664 5922 8728
rect 5986 8664 6003 8728
rect 6067 8664 6084 8728
rect 6148 8664 6165 8728
rect 6229 8664 6246 8728
rect 6310 8664 6327 8728
rect 6391 8664 6408 8728
rect 6472 8664 6489 8728
rect 6553 8664 6570 8728
rect 6634 8664 6651 8728
rect 6715 8664 6732 8728
rect 6796 8664 6813 8728
rect 6877 8664 6894 8728
rect 6958 8664 6975 8728
rect 7039 8664 7056 8728
rect 7120 8664 7137 8728
rect 7201 8664 7218 8728
rect 7282 8664 7299 8728
rect 7363 8664 7380 8728
rect 7444 8664 7461 8728
rect 7525 8664 7542 8728
rect 7606 8664 7623 8728
rect 7687 8664 7693 8728
rect 4689 8642 7693 8664
rect 4689 8578 4695 8642
rect 4759 8578 4777 8642
rect 4841 8578 4859 8642
rect 4923 8578 4941 8642
rect 5005 8578 5023 8642
rect 5087 8578 5105 8642
rect 5169 8578 5187 8642
rect 5251 8578 5269 8642
rect 5333 8578 5351 8642
rect 5415 8578 5433 8642
rect 5497 8578 5515 8642
rect 5579 8578 5597 8642
rect 5661 8578 5679 8642
rect 5743 8578 5760 8642
rect 5824 8578 5841 8642
rect 5905 8578 5922 8642
rect 5986 8578 6003 8642
rect 6067 8578 6084 8642
rect 6148 8578 6165 8642
rect 6229 8578 6246 8642
rect 6310 8578 6327 8642
rect 6391 8578 6408 8642
rect 6472 8578 6489 8642
rect 6553 8578 6570 8642
rect 6634 8578 6651 8642
rect 6715 8578 6732 8642
rect 6796 8578 6813 8642
rect 6877 8578 6894 8642
rect 6958 8578 6975 8642
rect 7039 8578 7056 8642
rect 7120 8578 7137 8642
rect 7201 8578 7218 8642
rect 7282 8578 7299 8642
rect 7363 8578 7380 8642
rect 7444 8578 7461 8642
rect 7525 8578 7542 8642
rect 7606 8578 7623 8642
rect 7687 8578 7693 8642
rect 4689 8556 7693 8578
rect 4689 8492 4695 8556
rect 4759 8492 4777 8556
rect 4841 8492 4859 8556
rect 4923 8492 4941 8556
rect 5005 8492 5023 8556
rect 5087 8492 5105 8556
rect 5169 8492 5187 8556
rect 5251 8492 5269 8556
rect 5333 8492 5351 8556
rect 5415 8492 5433 8556
rect 5497 8492 5515 8556
rect 5579 8492 5597 8556
rect 5661 8492 5679 8556
rect 5743 8492 5760 8556
rect 5824 8492 5841 8556
rect 5905 8492 5922 8556
rect 5986 8492 6003 8556
rect 6067 8492 6084 8556
rect 6148 8492 6165 8556
rect 6229 8492 6246 8556
rect 6310 8492 6327 8556
rect 6391 8492 6408 8556
rect 6472 8492 6489 8556
rect 6553 8492 6570 8556
rect 6634 8492 6651 8556
rect 6715 8492 6732 8556
rect 6796 8492 6813 8556
rect 6877 8492 6894 8556
rect 6958 8492 6975 8556
rect 7039 8492 7056 8556
rect 7120 8492 7137 8556
rect 7201 8492 7218 8556
rect 7282 8492 7299 8556
rect 7363 8492 7380 8556
rect 7444 8492 7461 8556
rect 7525 8492 7542 8556
rect 7606 8492 7623 8556
rect 7687 8492 7693 8556
rect 4689 8470 7693 8492
rect 4689 8406 4695 8470
rect 4759 8406 4777 8470
rect 4841 8406 4859 8470
rect 4923 8406 4941 8470
rect 5005 8406 5023 8470
rect 5087 8406 5105 8470
rect 5169 8406 5187 8470
rect 5251 8406 5269 8470
rect 5333 8406 5351 8470
rect 5415 8406 5433 8470
rect 5497 8406 5515 8470
rect 5579 8406 5597 8470
rect 5661 8406 5679 8470
rect 5743 8406 5760 8470
rect 5824 8406 5841 8470
rect 5905 8406 5922 8470
rect 5986 8406 6003 8470
rect 6067 8406 6084 8470
rect 6148 8406 6165 8470
rect 6229 8406 6246 8470
rect 6310 8406 6327 8470
rect 6391 8406 6408 8470
rect 6472 8406 6489 8470
rect 6553 8406 6570 8470
rect 6634 8406 6651 8470
rect 6715 8406 6732 8470
rect 6796 8406 6813 8470
rect 6877 8406 6894 8470
rect 6958 8406 6975 8470
rect 7039 8406 7056 8470
rect 7120 8406 7137 8470
rect 7201 8406 7218 8470
rect 7282 8406 7299 8470
rect 7363 8406 7380 8470
rect 7444 8406 7461 8470
rect 7525 8406 7542 8470
rect 7606 8406 7623 8470
rect 7687 8406 7693 8470
rect 4689 8384 7693 8406
rect 4689 8320 4695 8384
rect 4759 8320 4777 8384
rect 4841 8320 4859 8384
rect 4923 8320 4941 8384
rect 5005 8320 5023 8384
rect 5087 8320 5105 8384
rect 5169 8320 5187 8384
rect 5251 8320 5269 8384
rect 5333 8320 5351 8384
rect 5415 8320 5433 8384
rect 5497 8320 5515 8384
rect 5579 8320 5597 8384
rect 5661 8320 5679 8384
rect 5743 8320 5760 8384
rect 5824 8320 5841 8384
rect 5905 8320 5922 8384
rect 5986 8320 6003 8384
rect 6067 8320 6084 8384
rect 6148 8320 6165 8384
rect 6229 8320 6246 8384
rect 6310 8320 6327 8384
rect 6391 8320 6408 8384
rect 6472 8320 6489 8384
rect 6553 8320 6570 8384
rect 6634 8320 6651 8384
rect 6715 8320 6732 8384
rect 6796 8320 6813 8384
rect 6877 8320 6894 8384
rect 6958 8320 6975 8384
rect 7039 8320 7056 8384
rect 7120 8320 7137 8384
rect 7201 8320 7218 8384
rect 7282 8320 7299 8384
rect 7363 8320 7380 8384
rect 7444 8320 7461 8384
rect 7525 8320 7542 8384
rect 7606 8320 7623 8384
rect 7687 8320 7693 8384
rect 4689 0 7693 8320
rect 7813 38885 8213 40000
rect 7813 38829 7822 38885
rect 7878 38829 7904 38885
rect 7960 38829 7986 38885
rect 8042 38829 8067 38885
rect 8123 38829 8148 38885
rect 8204 38829 8213 38885
rect 7813 38741 8213 38829
rect 7813 38685 7822 38741
rect 7878 38685 7904 38741
rect 7960 38685 7986 38741
rect 8042 38685 8067 38741
rect 8123 38685 8148 38741
rect 8204 38685 8213 38741
rect 7813 36161 8213 38685
rect 7813 36105 7822 36161
rect 7878 36105 7904 36161
rect 7960 36105 7986 36161
rect 8042 36105 8067 36161
rect 8123 36105 8148 36161
rect 8204 36105 8213 36161
rect 7813 36017 8213 36105
rect 7813 35961 7822 36017
rect 7878 35961 7904 36017
rect 7960 35961 7986 36017
rect 8042 35961 8067 36017
rect 8123 35961 8148 36017
rect 8204 35961 8213 36017
rect 7813 34053 8213 35961
rect 7813 33997 7822 34053
rect 7878 33997 7904 34053
rect 7960 33997 7986 34053
rect 8042 33997 8067 34053
rect 8123 33997 8148 34053
rect 8204 33997 8213 34053
rect 7813 33909 8213 33997
rect 7813 33853 7822 33909
rect 7878 33853 7904 33909
rect 7960 33853 7986 33909
rect 8042 33853 8067 33909
rect 8123 33853 8148 33909
rect 8204 33853 8213 33909
rect 7813 31329 8213 33853
rect 7813 31273 7822 31329
rect 7878 31273 7904 31329
rect 7960 31273 7986 31329
rect 8042 31273 8067 31329
rect 8123 31273 8148 31329
rect 8204 31273 8213 31329
rect 7813 31185 8213 31273
rect 7813 31129 7822 31185
rect 7878 31129 7904 31185
rect 7960 31129 7986 31185
rect 8042 31129 8067 31185
rect 8123 31129 8148 31185
rect 8204 31129 8213 31185
rect 7813 29221 8213 31129
rect 7813 29165 7822 29221
rect 7878 29165 7904 29221
rect 7960 29165 7986 29221
rect 8042 29165 8067 29221
rect 8123 29165 8148 29221
rect 8204 29165 8213 29221
rect 7813 29077 8213 29165
rect 7813 29021 7822 29077
rect 7878 29021 7904 29077
rect 7960 29021 7986 29077
rect 8042 29021 8067 29077
rect 8123 29021 8148 29077
rect 8204 29021 8213 29077
rect 7813 26497 8213 29021
rect 7813 26441 7822 26497
rect 7878 26441 7904 26497
rect 7960 26441 7986 26497
rect 8042 26441 8067 26497
rect 8123 26441 8148 26497
rect 8204 26441 8213 26497
rect 7813 26353 8213 26441
rect 7813 26297 7822 26353
rect 7878 26297 7904 26353
rect 7960 26297 7986 26353
rect 8042 26297 8067 26353
rect 8123 26297 8148 26353
rect 8204 26297 8213 26353
rect 7813 24389 8213 26297
rect 7813 24333 7822 24389
rect 7878 24333 7904 24389
rect 7960 24333 7986 24389
rect 8042 24333 8067 24389
rect 8123 24333 8148 24389
rect 8204 24333 8213 24389
rect 7813 24245 8213 24333
rect 7813 24189 7822 24245
rect 7878 24189 7904 24245
rect 7960 24189 7986 24245
rect 8042 24189 8067 24245
rect 8123 24189 8148 24245
rect 8204 24189 8213 24245
rect 7813 21665 8213 24189
rect 7813 21609 7822 21665
rect 7878 21609 7904 21665
rect 7960 21609 7986 21665
rect 8042 21609 8067 21665
rect 8123 21609 8148 21665
rect 8204 21609 8213 21665
rect 7813 21521 8213 21609
rect 7813 21465 7822 21521
rect 7878 21465 7904 21521
rect 7960 21465 7986 21521
rect 8042 21465 8067 21521
rect 8123 21465 8148 21521
rect 8204 21465 8213 21521
rect 7813 19557 8213 21465
rect 7813 19501 7822 19557
rect 7878 19501 7904 19557
rect 7960 19501 7986 19557
rect 8042 19501 8067 19557
rect 8123 19501 8148 19557
rect 8204 19501 8213 19557
rect 7813 19413 8213 19501
rect 7813 19357 7822 19413
rect 7878 19357 7904 19413
rect 7960 19357 7986 19413
rect 8042 19357 8067 19413
rect 8123 19357 8148 19413
rect 8204 19357 8213 19413
rect 7813 16833 8213 19357
rect 7813 16777 7822 16833
rect 7878 16777 7904 16833
rect 7960 16777 7986 16833
rect 8042 16777 8067 16833
rect 8123 16777 8148 16833
rect 8204 16777 8213 16833
rect 7813 16689 8213 16777
rect 7813 16633 7822 16689
rect 7878 16633 7904 16689
rect 7960 16633 7986 16689
rect 8042 16633 8067 16689
rect 8123 16633 8148 16689
rect 8204 16633 8213 16689
rect 7813 14725 8213 16633
rect 7813 14669 7822 14725
rect 7878 14669 7904 14725
rect 7960 14669 7986 14725
rect 8042 14669 8067 14725
rect 8123 14669 8148 14725
rect 8204 14669 8213 14725
rect 7813 14581 8213 14669
rect 7813 14525 7822 14581
rect 7878 14525 7904 14581
rect 7960 14525 7986 14581
rect 8042 14525 8067 14581
rect 8123 14525 8148 14581
rect 8204 14525 8213 14581
rect 7813 12001 8213 14525
rect 7813 11945 7822 12001
rect 7878 11945 7904 12001
rect 7960 11945 7986 12001
rect 8042 11945 8067 12001
rect 8123 11945 8148 12001
rect 8204 11945 8213 12001
rect 7813 11857 8213 11945
rect 7813 11801 7822 11857
rect 7878 11801 7904 11857
rect 7960 11801 7986 11857
rect 8042 11801 8067 11857
rect 8123 11801 8148 11857
rect 8204 11801 8213 11857
rect 7813 9893 8213 11801
rect 7813 9837 7822 9893
rect 7878 9837 7904 9893
rect 7960 9837 7986 9893
rect 8042 9837 8067 9893
rect 8123 9837 8148 9893
rect 8204 9837 8213 9893
rect 7813 9749 8213 9837
rect 7813 9693 7822 9749
rect 7878 9693 7904 9749
rect 7960 9693 7986 9749
rect 8042 9693 8067 9749
rect 8123 9693 8148 9749
rect 8204 9693 8213 9749
rect 7813 9241 8213 9693
rect 7877 9177 7897 9241
rect 7961 9177 7981 9241
rect 8045 9177 8065 9241
rect 8129 9177 8149 9241
rect 7813 9156 8213 9177
rect 7877 9092 7897 9156
rect 7961 9092 7981 9156
rect 8045 9092 8065 9156
rect 8129 9092 8149 9156
rect 7813 9071 8213 9092
rect 7877 9007 7897 9071
rect 7961 9007 7981 9071
rect 8045 9007 8065 9071
rect 8129 9007 8149 9071
rect 7813 8986 8213 9007
rect 7877 8922 7897 8986
rect 7961 8922 7981 8986
rect 8045 8922 8065 8986
rect 8129 8922 8149 8986
rect 7813 8901 8213 8922
rect 7877 8837 7897 8901
rect 7961 8837 7981 8901
rect 8045 8837 8065 8901
rect 8129 8837 8149 8901
rect 7813 8816 8213 8837
rect 7877 8752 7897 8816
rect 7961 8752 7981 8816
rect 8045 8752 8065 8816
rect 8129 8752 8149 8816
rect 7813 8731 8213 8752
rect 7877 8667 7897 8731
rect 7961 8667 7981 8731
rect 8045 8667 8065 8731
rect 8129 8667 8149 8731
rect 7813 8645 8213 8667
rect 7877 8581 7897 8645
rect 7961 8581 7981 8645
rect 8045 8581 8065 8645
rect 8129 8581 8149 8645
rect 7813 8559 8213 8581
rect 7877 8495 7897 8559
rect 7961 8495 7981 8559
rect 8045 8495 8065 8559
rect 8129 8495 8149 8559
rect 7813 8473 8213 8495
rect 7877 8409 7897 8473
rect 7961 8409 7981 8473
rect 8045 8409 8065 8473
rect 8129 8409 8149 8473
rect 7813 8387 8213 8409
rect 7877 8323 7897 8387
rect 7961 8323 7981 8387
rect 8045 8323 8065 8387
rect 8129 8323 8149 8387
rect 7813 7729 8213 8323
rect 7813 7673 7823 7729
rect 7879 7673 7932 7729
rect 7988 7673 8040 7729
rect 8096 7673 8148 7729
rect 8204 7673 8213 7729
rect 7813 7169 8213 7673
rect 7813 7113 7822 7169
rect 7878 7113 7904 7169
rect 7960 7113 7986 7169
rect 8042 7113 8067 7169
rect 8123 7113 8148 7169
rect 8204 7113 8213 7169
rect 7813 7025 8213 7113
rect 7813 6969 7822 7025
rect 7878 6969 7904 7025
rect 7960 6969 7986 7025
rect 8042 6969 8067 7025
rect 8123 6969 8148 7025
rect 8204 6969 8213 7025
rect 7813 2337 8213 6969
rect 7813 2281 7822 2337
rect 7878 2281 7904 2337
rect 7960 2281 7986 2337
rect 8042 2281 8067 2337
rect 8123 2281 8148 2337
rect 8204 2281 8213 2337
rect 7813 2193 8213 2281
rect 7813 2137 7822 2193
rect 7878 2137 7904 2193
rect 7960 2137 7986 2193
rect 8042 2137 8067 2193
rect 8123 2137 8148 2193
rect 8204 2137 8213 2193
rect 7813 907 8213 2137
rect 7813 851 7835 907
rect 7891 851 7979 907
rect 8035 851 8213 907
rect 7813 802 8213 851
rect 7813 746 7835 802
rect 7891 746 7979 802
rect 8035 746 8213 802
rect 7813 697 8213 746
rect 7813 641 7835 697
rect 7891 641 7979 697
rect 8035 641 8213 697
rect 7813 591 8213 641
rect 7813 535 7835 591
rect 7891 535 7979 591
rect 8035 535 8213 591
rect 7813 485 8213 535
rect 7813 429 7835 485
rect 7891 429 7979 485
rect 8035 429 8213 485
rect 7813 379 8213 429
rect 7813 323 7835 379
rect 7891 323 7979 379
rect 8035 323 8213 379
rect 7813 0 8213 323
rect 8333 39141 8733 40000
rect 8333 39085 8342 39141
rect 8398 39085 8424 39141
rect 8480 39085 8506 39141
rect 8562 39085 8587 39141
rect 8643 39085 8668 39141
rect 8724 39085 8733 39141
rect 8333 38997 8733 39085
rect 8333 38941 8342 38997
rect 8398 38941 8424 38997
rect 8480 38941 8506 38997
rect 8562 38941 8587 38997
rect 8643 38941 8668 38997
rect 8724 38941 8733 38997
rect 8333 36417 8733 38941
rect 8333 36361 8342 36417
rect 8398 36361 8424 36417
rect 8480 36361 8506 36417
rect 8562 36361 8587 36417
rect 8643 36361 8668 36417
rect 8724 36361 8733 36417
rect 8333 36273 8733 36361
rect 8333 36217 8342 36273
rect 8398 36217 8424 36273
rect 8480 36217 8506 36273
rect 8562 36217 8587 36273
rect 8643 36217 8668 36273
rect 8724 36217 8733 36273
rect 8333 34309 8733 36217
rect 8333 34253 8342 34309
rect 8398 34253 8424 34309
rect 8480 34253 8506 34309
rect 8562 34253 8587 34309
rect 8643 34253 8668 34309
rect 8724 34253 8733 34309
rect 8333 34165 8733 34253
rect 8333 34109 8342 34165
rect 8398 34109 8424 34165
rect 8480 34109 8506 34165
rect 8562 34109 8587 34165
rect 8643 34109 8668 34165
rect 8724 34109 8733 34165
rect 8333 31585 8733 34109
rect 8333 31529 8342 31585
rect 8398 31529 8424 31585
rect 8480 31529 8506 31585
rect 8562 31529 8587 31585
rect 8643 31529 8668 31585
rect 8724 31529 8733 31585
rect 8333 31441 8733 31529
rect 8333 31385 8342 31441
rect 8398 31385 8424 31441
rect 8480 31385 8506 31441
rect 8562 31385 8587 31441
rect 8643 31385 8668 31441
rect 8724 31385 8733 31441
rect 8333 29477 8733 31385
rect 8333 29421 8342 29477
rect 8398 29421 8424 29477
rect 8480 29421 8506 29477
rect 8562 29421 8587 29477
rect 8643 29421 8668 29477
rect 8724 29421 8733 29477
rect 8333 29333 8733 29421
rect 8333 29277 8342 29333
rect 8398 29277 8424 29333
rect 8480 29277 8506 29333
rect 8562 29277 8587 29333
rect 8643 29277 8668 29333
rect 8724 29277 8733 29333
rect 8333 26753 8733 29277
rect 8333 26697 8342 26753
rect 8398 26697 8424 26753
rect 8480 26697 8506 26753
rect 8562 26697 8587 26753
rect 8643 26697 8668 26753
rect 8724 26697 8733 26753
rect 8333 26609 8733 26697
rect 8333 26553 8342 26609
rect 8398 26553 8424 26609
rect 8480 26553 8506 26609
rect 8562 26553 8587 26609
rect 8643 26553 8668 26609
rect 8724 26553 8733 26609
rect 8333 24645 8733 26553
rect 8333 24589 8342 24645
rect 8398 24589 8424 24645
rect 8480 24589 8506 24645
rect 8562 24589 8587 24645
rect 8643 24589 8668 24645
rect 8724 24589 8733 24645
rect 8333 24501 8733 24589
rect 8333 24445 8342 24501
rect 8398 24445 8424 24501
rect 8480 24445 8506 24501
rect 8562 24445 8587 24501
rect 8643 24445 8668 24501
rect 8724 24445 8733 24501
rect 8333 21921 8733 24445
rect 8333 21865 8342 21921
rect 8398 21865 8424 21921
rect 8480 21865 8506 21921
rect 8562 21865 8587 21921
rect 8643 21865 8668 21921
rect 8724 21865 8733 21921
rect 8333 21777 8733 21865
rect 8333 21721 8342 21777
rect 8398 21721 8424 21777
rect 8480 21721 8506 21777
rect 8562 21721 8587 21777
rect 8643 21721 8668 21777
rect 8724 21721 8733 21777
rect 8333 19813 8733 21721
rect 8333 19757 8342 19813
rect 8398 19757 8424 19813
rect 8480 19757 8506 19813
rect 8562 19757 8587 19813
rect 8643 19757 8668 19813
rect 8724 19757 8733 19813
rect 8333 19669 8733 19757
rect 8333 19613 8342 19669
rect 8398 19613 8424 19669
rect 8480 19613 8506 19669
rect 8562 19613 8587 19669
rect 8643 19613 8668 19669
rect 8724 19613 8733 19669
rect 8333 17089 8733 19613
rect 8333 17033 8342 17089
rect 8398 17033 8424 17089
rect 8480 17033 8506 17089
rect 8562 17033 8587 17089
rect 8643 17033 8668 17089
rect 8724 17033 8733 17089
rect 8333 16945 8733 17033
rect 8333 16889 8342 16945
rect 8398 16889 8424 16945
rect 8480 16889 8506 16945
rect 8562 16889 8587 16945
rect 8643 16889 8668 16945
rect 8724 16889 8733 16945
rect 8333 14981 8733 16889
rect 8333 14925 8342 14981
rect 8398 14925 8424 14981
rect 8480 14925 8506 14981
rect 8562 14925 8587 14981
rect 8643 14925 8668 14981
rect 8724 14925 8733 14981
rect 8333 14837 8733 14925
rect 8333 14781 8342 14837
rect 8398 14781 8424 14837
rect 8480 14781 8506 14837
rect 8562 14781 8587 14837
rect 8643 14781 8668 14837
rect 8724 14781 8733 14837
rect 8333 13701 8733 14781
rect 8397 13637 8417 13701
rect 8481 13637 8501 13701
rect 8565 13637 8585 13701
rect 8649 13637 8669 13701
rect 8333 13620 8733 13637
rect 8397 13556 8417 13620
rect 8481 13556 8501 13620
rect 8565 13556 8585 13620
rect 8649 13556 8669 13620
rect 8333 13539 8733 13556
rect 8397 13475 8417 13539
rect 8481 13475 8501 13539
rect 8565 13475 8585 13539
rect 8649 13475 8669 13539
rect 8333 13458 8733 13475
rect 8397 13394 8417 13458
rect 8481 13394 8501 13458
rect 8565 13394 8585 13458
rect 8649 13394 8669 13458
rect 8333 13377 8733 13394
rect 8397 13313 8417 13377
rect 8481 13313 8501 13377
rect 8565 13313 8585 13377
rect 8649 13313 8669 13377
rect 8333 13296 8733 13313
rect 8397 13232 8417 13296
rect 8481 13232 8501 13296
rect 8565 13232 8585 13296
rect 8649 13232 8669 13296
rect 8333 13215 8733 13232
rect 8397 13151 8417 13215
rect 8481 13151 8501 13215
rect 8565 13151 8585 13215
rect 8649 13151 8669 13215
rect 8333 13133 8733 13151
rect 8397 13069 8417 13133
rect 8481 13069 8501 13133
rect 8565 13069 8585 13133
rect 8649 13069 8669 13133
rect 8333 13051 8733 13069
rect 8397 12987 8417 13051
rect 8481 12987 8501 13051
rect 8565 12987 8585 13051
rect 8649 12987 8669 13051
rect 8333 12969 8733 12987
rect 8397 12905 8417 12969
rect 8481 12905 8501 12969
rect 8565 12905 8585 12969
rect 8649 12905 8669 12969
rect 8333 12887 8733 12905
rect 8397 12823 8417 12887
rect 8481 12823 8501 12887
rect 8565 12823 8585 12887
rect 8649 12823 8669 12887
rect 8333 12257 8733 12823
rect 8333 12201 8342 12257
rect 8398 12201 8424 12257
rect 8480 12201 8506 12257
rect 8562 12201 8587 12257
rect 8643 12201 8668 12257
rect 8724 12201 8733 12257
rect 8333 12113 8733 12201
rect 8333 12057 8342 12113
rect 8398 12057 8424 12113
rect 8480 12057 8506 12113
rect 8562 12057 8587 12113
rect 8643 12057 8668 12113
rect 8724 12057 8733 12113
rect 8333 10149 8733 12057
rect 8333 10093 8342 10149
rect 8398 10093 8424 10149
rect 8480 10093 8506 10149
rect 8562 10093 8587 10149
rect 8643 10093 8668 10149
rect 8724 10093 8733 10149
rect 8333 10005 8733 10093
rect 8333 9949 8342 10005
rect 8398 9949 8424 10005
rect 8480 9949 8506 10005
rect 8562 9949 8587 10005
rect 8643 9949 8668 10005
rect 8724 9949 8733 10005
rect 8333 7425 8733 9949
rect 8333 7369 8342 7425
rect 8398 7369 8424 7425
rect 8480 7369 8506 7425
rect 8562 7369 8587 7425
rect 8643 7369 8668 7425
rect 8724 7369 8733 7425
rect 8333 7281 8733 7369
rect 8333 7225 8342 7281
rect 8398 7225 8424 7281
rect 8480 7225 8506 7281
rect 8562 7225 8587 7281
rect 8643 7225 8668 7281
rect 8724 7225 8733 7281
rect 8333 2593 8733 7225
rect 8333 2537 8342 2593
rect 8398 2537 8424 2593
rect 8480 2537 8506 2593
rect 8562 2537 8587 2593
rect 8643 2537 8668 2593
rect 8724 2537 8733 2593
rect 8333 2449 8733 2537
rect 8333 2393 8342 2449
rect 8398 2393 8424 2449
rect 8480 2393 8506 2449
rect 8562 2393 8587 2449
rect 8643 2393 8668 2449
rect 8724 2393 8733 2449
rect 8333 321 8733 2393
rect 8333 265 8342 321
rect 8398 265 8424 321
rect 8480 265 8506 321
rect 8562 265 8587 321
rect 8643 265 8668 321
rect 8724 265 8733 321
rect 8333 175 8733 265
rect 8333 119 8342 175
rect 8398 119 8424 175
rect 8480 119 8506 175
rect 8562 119 8587 175
rect 8643 119 8668 175
rect 8724 119 8733 175
rect 8333 0 8733 119
rect 8853 9244 11983 40000
rect 8853 9180 8859 9244
rect 8923 9180 8940 9244
rect 9004 9180 9021 9244
rect 9085 9180 9102 9244
rect 9166 9180 9183 9244
rect 9247 9180 9264 9244
rect 9328 9180 9345 9244
rect 9409 9180 9426 9244
rect 9490 9180 9507 9244
rect 9571 9180 9588 9244
rect 9652 9180 9669 9244
rect 9733 9180 9750 9244
rect 9814 9180 9831 9244
rect 9895 9180 9912 9244
rect 9976 9180 9993 9244
rect 10057 9180 10073 9244
rect 10137 9180 10153 9244
rect 10217 9180 10233 9244
rect 10297 9180 10313 9244
rect 10377 9180 10393 9244
rect 10457 9180 10473 9244
rect 10537 9180 10553 9244
rect 10617 9180 10633 9244
rect 10697 9180 10713 9244
rect 10777 9180 10793 9244
rect 10857 9180 10873 9244
rect 10937 9180 10953 9244
rect 11017 9180 11033 9244
rect 11097 9180 11113 9244
rect 11177 9180 11193 9244
rect 11257 9180 11273 9244
rect 11337 9180 11353 9244
rect 11417 9180 11433 9244
rect 11497 9180 11513 9244
rect 11577 9180 11593 9244
rect 11657 9180 11673 9244
rect 11737 9180 11753 9244
rect 11817 9180 11833 9244
rect 11897 9180 11913 9244
rect 11977 9180 11983 9244
rect 8853 9158 11983 9180
rect 8853 9094 8859 9158
rect 8923 9094 8940 9158
rect 9004 9094 9021 9158
rect 9085 9094 9102 9158
rect 9166 9094 9183 9158
rect 9247 9094 9264 9158
rect 9328 9094 9345 9158
rect 9409 9094 9426 9158
rect 9490 9094 9507 9158
rect 9571 9094 9588 9158
rect 9652 9094 9669 9158
rect 9733 9094 9750 9158
rect 9814 9094 9831 9158
rect 9895 9094 9912 9158
rect 9976 9094 9993 9158
rect 10057 9094 10073 9158
rect 10137 9094 10153 9158
rect 10217 9094 10233 9158
rect 10297 9094 10313 9158
rect 10377 9094 10393 9158
rect 10457 9094 10473 9158
rect 10537 9094 10553 9158
rect 10617 9094 10633 9158
rect 10697 9094 10713 9158
rect 10777 9094 10793 9158
rect 10857 9094 10873 9158
rect 10937 9094 10953 9158
rect 11017 9094 11033 9158
rect 11097 9094 11113 9158
rect 11177 9094 11193 9158
rect 11257 9094 11273 9158
rect 11337 9094 11353 9158
rect 11417 9094 11433 9158
rect 11497 9094 11513 9158
rect 11577 9094 11593 9158
rect 11657 9094 11673 9158
rect 11737 9094 11753 9158
rect 11817 9094 11833 9158
rect 11897 9094 11913 9158
rect 11977 9094 11983 9158
rect 8853 9072 11983 9094
rect 8853 9008 8859 9072
rect 8923 9008 8940 9072
rect 9004 9008 9021 9072
rect 9085 9008 9102 9072
rect 9166 9008 9183 9072
rect 9247 9008 9264 9072
rect 9328 9008 9345 9072
rect 9409 9008 9426 9072
rect 9490 9008 9507 9072
rect 9571 9008 9588 9072
rect 9652 9008 9669 9072
rect 9733 9008 9750 9072
rect 9814 9008 9831 9072
rect 9895 9008 9912 9072
rect 9976 9008 9993 9072
rect 10057 9008 10073 9072
rect 10137 9008 10153 9072
rect 10217 9008 10233 9072
rect 10297 9008 10313 9072
rect 10377 9008 10393 9072
rect 10457 9008 10473 9072
rect 10537 9008 10553 9072
rect 10617 9008 10633 9072
rect 10697 9008 10713 9072
rect 10777 9008 10793 9072
rect 10857 9008 10873 9072
rect 10937 9008 10953 9072
rect 11017 9008 11033 9072
rect 11097 9008 11113 9072
rect 11177 9008 11193 9072
rect 11257 9008 11273 9072
rect 11337 9008 11353 9072
rect 11417 9008 11433 9072
rect 11497 9008 11513 9072
rect 11577 9008 11593 9072
rect 11657 9008 11673 9072
rect 11737 9008 11753 9072
rect 11817 9008 11833 9072
rect 11897 9008 11913 9072
rect 11977 9008 11983 9072
rect 8853 8986 11983 9008
rect 8853 8922 8859 8986
rect 8923 8922 8940 8986
rect 9004 8922 9021 8986
rect 9085 8922 9102 8986
rect 9166 8922 9183 8986
rect 9247 8922 9264 8986
rect 9328 8922 9345 8986
rect 9409 8922 9426 8986
rect 9490 8922 9507 8986
rect 9571 8922 9588 8986
rect 9652 8922 9669 8986
rect 9733 8922 9750 8986
rect 9814 8922 9831 8986
rect 9895 8922 9912 8986
rect 9976 8922 9993 8986
rect 10057 8922 10073 8986
rect 10137 8922 10153 8986
rect 10217 8922 10233 8986
rect 10297 8922 10313 8986
rect 10377 8922 10393 8986
rect 10457 8922 10473 8986
rect 10537 8922 10553 8986
rect 10617 8922 10633 8986
rect 10697 8922 10713 8986
rect 10777 8922 10793 8986
rect 10857 8922 10873 8986
rect 10937 8922 10953 8986
rect 11017 8922 11033 8986
rect 11097 8922 11113 8986
rect 11177 8922 11193 8986
rect 11257 8922 11273 8986
rect 11337 8922 11353 8986
rect 11417 8922 11433 8986
rect 11497 8922 11513 8986
rect 11577 8922 11593 8986
rect 11657 8922 11673 8986
rect 11737 8922 11753 8986
rect 11817 8922 11833 8986
rect 11897 8922 11913 8986
rect 11977 8922 11983 8986
rect 8853 8900 11983 8922
rect 8853 8836 8859 8900
rect 8923 8836 8940 8900
rect 9004 8836 9021 8900
rect 9085 8836 9102 8900
rect 9166 8836 9183 8900
rect 9247 8836 9264 8900
rect 9328 8836 9345 8900
rect 9409 8836 9426 8900
rect 9490 8836 9507 8900
rect 9571 8836 9588 8900
rect 9652 8836 9669 8900
rect 9733 8836 9750 8900
rect 9814 8836 9831 8900
rect 9895 8836 9912 8900
rect 9976 8836 9993 8900
rect 10057 8836 10073 8900
rect 10137 8836 10153 8900
rect 10217 8836 10233 8900
rect 10297 8836 10313 8900
rect 10377 8836 10393 8900
rect 10457 8836 10473 8900
rect 10537 8836 10553 8900
rect 10617 8836 10633 8900
rect 10697 8836 10713 8900
rect 10777 8836 10793 8900
rect 10857 8836 10873 8900
rect 10937 8836 10953 8900
rect 11017 8836 11033 8900
rect 11097 8836 11113 8900
rect 11177 8836 11193 8900
rect 11257 8836 11273 8900
rect 11337 8836 11353 8900
rect 11417 8836 11433 8900
rect 11497 8836 11513 8900
rect 11577 8836 11593 8900
rect 11657 8836 11673 8900
rect 11737 8836 11753 8900
rect 11817 8836 11833 8900
rect 11897 8836 11913 8900
rect 11977 8836 11983 8900
rect 8853 8814 11983 8836
rect 8853 8750 8859 8814
rect 8923 8750 8940 8814
rect 9004 8750 9021 8814
rect 9085 8750 9102 8814
rect 9166 8750 9183 8814
rect 9247 8750 9264 8814
rect 9328 8750 9345 8814
rect 9409 8750 9426 8814
rect 9490 8750 9507 8814
rect 9571 8750 9588 8814
rect 9652 8750 9669 8814
rect 9733 8750 9750 8814
rect 9814 8750 9831 8814
rect 9895 8750 9912 8814
rect 9976 8750 9993 8814
rect 10057 8750 10073 8814
rect 10137 8750 10153 8814
rect 10217 8750 10233 8814
rect 10297 8750 10313 8814
rect 10377 8750 10393 8814
rect 10457 8750 10473 8814
rect 10537 8750 10553 8814
rect 10617 8750 10633 8814
rect 10697 8750 10713 8814
rect 10777 8750 10793 8814
rect 10857 8750 10873 8814
rect 10937 8750 10953 8814
rect 11017 8750 11033 8814
rect 11097 8750 11113 8814
rect 11177 8750 11193 8814
rect 11257 8750 11273 8814
rect 11337 8750 11353 8814
rect 11417 8750 11433 8814
rect 11497 8750 11513 8814
rect 11577 8750 11593 8814
rect 11657 8750 11673 8814
rect 11737 8750 11753 8814
rect 11817 8750 11833 8814
rect 11897 8750 11913 8814
rect 11977 8750 11983 8814
rect 8853 8728 11983 8750
rect 8853 8664 8859 8728
rect 8923 8664 8940 8728
rect 9004 8664 9021 8728
rect 9085 8664 9102 8728
rect 9166 8664 9183 8728
rect 9247 8664 9264 8728
rect 9328 8664 9345 8728
rect 9409 8664 9426 8728
rect 9490 8664 9507 8728
rect 9571 8664 9588 8728
rect 9652 8664 9669 8728
rect 9733 8664 9750 8728
rect 9814 8664 9831 8728
rect 9895 8664 9912 8728
rect 9976 8664 9993 8728
rect 10057 8664 10073 8728
rect 10137 8664 10153 8728
rect 10217 8664 10233 8728
rect 10297 8664 10313 8728
rect 10377 8664 10393 8728
rect 10457 8664 10473 8728
rect 10537 8664 10553 8728
rect 10617 8664 10633 8728
rect 10697 8664 10713 8728
rect 10777 8664 10793 8728
rect 10857 8664 10873 8728
rect 10937 8664 10953 8728
rect 11017 8664 11033 8728
rect 11097 8664 11113 8728
rect 11177 8664 11193 8728
rect 11257 8664 11273 8728
rect 11337 8664 11353 8728
rect 11417 8664 11433 8728
rect 11497 8664 11513 8728
rect 11577 8664 11593 8728
rect 11657 8664 11673 8728
rect 11737 8664 11753 8728
rect 11817 8664 11833 8728
rect 11897 8664 11913 8728
rect 11977 8664 11983 8728
rect 8853 8642 11983 8664
rect 8853 8578 8859 8642
rect 8923 8578 8940 8642
rect 9004 8578 9021 8642
rect 9085 8578 9102 8642
rect 9166 8578 9183 8642
rect 9247 8578 9264 8642
rect 9328 8578 9345 8642
rect 9409 8578 9426 8642
rect 9490 8578 9507 8642
rect 9571 8578 9588 8642
rect 9652 8578 9669 8642
rect 9733 8578 9750 8642
rect 9814 8578 9831 8642
rect 9895 8578 9912 8642
rect 9976 8578 9993 8642
rect 10057 8578 10073 8642
rect 10137 8578 10153 8642
rect 10217 8578 10233 8642
rect 10297 8578 10313 8642
rect 10377 8578 10393 8642
rect 10457 8578 10473 8642
rect 10537 8578 10553 8642
rect 10617 8578 10633 8642
rect 10697 8578 10713 8642
rect 10777 8578 10793 8642
rect 10857 8578 10873 8642
rect 10937 8578 10953 8642
rect 11017 8578 11033 8642
rect 11097 8578 11113 8642
rect 11177 8578 11193 8642
rect 11257 8578 11273 8642
rect 11337 8578 11353 8642
rect 11417 8578 11433 8642
rect 11497 8578 11513 8642
rect 11577 8578 11593 8642
rect 11657 8578 11673 8642
rect 11737 8578 11753 8642
rect 11817 8578 11833 8642
rect 11897 8578 11913 8642
rect 11977 8578 11983 8642
rect 8853 8556 11983 8578
rect 8853 8492 8859 8556
rect 8923 8492 8940 8556
rect 9004 8492 9021 8556
rect 9085 8492 9102 8556
rect 9166 8492 9183 8556
rect 9247 8492 9264 8556
rect 9328 8492 9345 8556
rect 9409 8492 9426 8556
rect 9490 8492 9507 8556
rect 9571 8492 9588 8556
rect 9652 8492 9669 8556
rect 9733 8492 9750 8556
rect 9814 8492 9831 8556
rect 9895 8492 9912 8556
rect 9976 8492 9993 8556
rect 10057 8492 10073 8556
rect 10137 8492 10153 8556
rect 10217 8492 10233 8556
rect 10297 8492 10313 8556
rect 10377 8492 10393 8556
rect 10457 8492 10473 8556
rect 10537 8492 10553 8556
rect 10617 8492 10633 8556
rect 10697 8492 10713 8556
rect 10777 8492 10793 8556
rect 10857 8492 10873 8556
rect 10937 8492 10953 8556
rect 11017 8492 11033 8556
rect 11097 8492 11113 8556
rect 11177 8492 11193 8556
rect 11257 8492 11273 8556
rect 11337 8492 11353 8556
rect 11417 8492 11433 8556
rect 11497 8492 11513 8556
rect 11577 8492 11593 8556
rect 11657 8492 11673 8556
rect 11737 8492 11753 8556
rect 11817 8492 11833 8556
rect 11897 8492 11913 8556
rect 11977 8492 11983 8556
rect 8853 8470 11983 8492
rect 8853 8406 8859 8470
rect 8923 8406 8940 8470
rect 9004 8406 9021 8470
rect 9085 8406 9102 8470
rect 9166 8406 9183 8470
rect 9247 8406 9264 8470
rect 9328 8406 9345 8470
rect 9409 8406 9426 8470
rect 9490 8406 9507 8470
rect 9571 8406 9588 8470
rect 9652 8406 9669 8470
rect 9733 8406 9750 8470
rect 9814 8406 9831 8470
rect 9895 8406 9912 8470
rect 9976 8406 9993 8470
rect 10057 8406 10073 8470
rect 10137 8406 10153 8470
rect 10217 8406 10233 8470
rect 10297 8406 10313 8470
rect 10377 8406 10393 8470
rect 10457 8406 10473 8470
rect 10537 8406 10553 8470
rect 10617 8406 10633 8470
rect 10697 8406 10713 8470
rect 10777 8406 10793 8470
rect 10857 8406 10873 8470
rect 10937 8406 10953 8470
rect 11017 8406 11033 8470
rect 11097 8406 11113 8470
rect 11177 8406 11193 8470
rect 11257 8406 11273 8470
rect 11337 8406 11353 8470
rect 11417 8406 11433 8470
rect 11497 8406 11513 8470
rect 11577 8406 11593 8470
rect 11657 8406 11673 8470
rect 11737 8406 11753 8470
rect 11817 8406 11833 8470
rect 11897 8406 11913 8470
rect 11977 8406 11983 8470
rect 8853 8384 11983 8406
rect 8853 8320 8859 8384
rect 8923 8320 8940 8384
rect 9004 8320 9021 8384
rect 9085 8320 9102 8384
rect 9166 8320 9183 8384
rect 9247 8320 9264 8384
rect 9328 8320 9345 8384
rect 9409 8320 9426 8384
rect 9490 8320 9507 8384
rect 9571 8320 9588 8384
rect 9652 8320 9669 8384
rect 9733 8320 9750 8384
rect 9814 8320 9831 8384
rect 9895 8320 9912 8384
rect 9976 8320 9993 8384
rect 10057 8320 10073 8384
rect 10137 8320 10153 8384
rect 10217 8320 10233 8384
rect 10297 8320 10313 8384
rect 10377 8320 10393 8384
rect 10457 8320 10473 8384
rect 10537 8320 10553 8384
rect 10617 8320 10633 8384
rect 10697 8320 10713 8384
rect 10777 8320 10793 8384
rect 10857 8320 10873 8384
rect 10937 8320 10953 8384
rect 11017 8320 11033 8384
rect 11097 8320 11113 8384
rect 11177 8320 11193 8384
rect 11257 8320 11273 8384
rect 11337 8320 11353 8384
rect 11417 8320 11433 8384
rect 11497 8320 11513 8384
rect 11577 8320 11593 8384
rect 11657 8320 11673 8384
rect 11737 8320 11753 8384
rect 11817 8320 11833 8384
rect 11897 8320 11913 8384
rect 11977 8320 11983 8384
rect 8853 3725 11983 8320
rect 8853 840 11082 3725
tri 11082 2824 11983 3725 nw
rect 12159 9244 15623 40000
rect 12159 9180 12165 9244
rect 12229 9180 12246 9244
rect 12310 9180 12327 9244
rect 12391 9180 12408 9244
rect 12472 9180 12489 9244
rect 12553 9180 12570 9244
rect 12634 9180 12651 9244
rect 12715 9180 12732 9244
rect 12796 9180 12813 9244
rect 12877 9180 12894 9244
rect 12958 9180 12975 9244
rect 13039 9180 13056 9244
rect 13120 9180 13137 9244
rect 13201 9180 13218 9244
rect 13282 9180 13299 9244
rect 13363 9180 13380 9244
rect 13444 9180 13461 9244
rect 13525 9180 13542 9244
rect 13606 9180 13623 9244
rect 13687 9180 13704 9244
rect 13768 9180 13785 9244
rect 13849 9180 13866 9244
rect 13930 9180 13947 9244
rect 14011 9180 14028 9244
rect 14092 9180 14109 9244
rect 14173 9180 14190 9244
rect 14254 9180 14271 9244
rect 14335 9180 14352 9244
rect 14416 9180 14433 9244
rect 14497 9180 14513 9244
rect 14577 9180 14593 9244
rect 14657 9180 14673 9244
rect 14737 9180 14753 9244
rect 14817 9180 14833 9244
rect 14897 9180 14913 9244
rect 14977 9180 14993 9244
rect 15057 9180 15073 9244
rect 15137 9180 15153 9244
rect 15217 9180 15233 9244
rect 15297 9180 15313 9244
rect 15377 9180 15393 9244
rect 15457 9180 15473 9244
rect 15537 9180 15553 9244
rect 15617 9180 15623 9244
rect 12159 9158 15623 9180
rect 12159 9094 12165 9158
rect 12229 9094 12246 9158
rect 12310 9094 12327 9158
rect 12391 9094 12408 9158
rect 12472 9094 12489 9158
rect 12553 9094 12570 9158
rect 12634 9094 12651 9158
rect 12715 9094 12732 9158
rect 12796 9094 12813 9158
rect 12877 9094 12894 9158
rect 12958 9094 12975 9158
rect 13039 9094 13056 9158
rect 13120 9094 13137 9158
rect 13201 9094 13218 9158
rect 13282 9094 13299 9158
rect 13363 9094 13380 9158
rect 13444 9094 13461 9158
rect 13525 9094 13542 9158
rect 13606 9094 13623 9158
rect 13687 9094 13704 9158
rect 13768 9094 13785 9158
rect 13849 9094 13866 9158
rect 13930 9094 13947 9158
rect 14011 9094 14028 9158
rect 14092 9094 14109 9158
rect 14173 9094 14190 9158
rect 14254 9094 14271 9158
rect 14335 9094 14352 9158
rect 14416 9094 14433 9158
rect 14497 9094 14513 9158
rect 14577 9094 14593 9158
rect 14657 9094 14673 9158
rect 14737 9094 14753 9158
rect 14817 9094 14833 9158
rect 14897 9094 14913 9158
rect 14977 9094 14993 9158
rect 15057 9094 15073 9158
rect 15137 9094 15153 9158
rect 15217 9094 15233 9158
rect 15297 9094 15313 9158
rect 15377 9094 15393 9158
rect 15457 9094 15473 9158
rect 15537 9094 15553 9158
rect 15617 9094 15623 9158
rect 12159 9072 15623 9094
rect 12159 9008 12165 9072
rect 12229 9008 12246 9072
rect 12310 9008 12327 9072
rect 12391 9008 12408 9072
rect 12472 9008 12489 9072
rect 12553 9008 12570 9072
rect 12634 9008 12651 9072
rect 12715 9008 12732 9072
rect 12796 9008 12813 9072
rect 12877 9008 12894 9072
rect 12958 9008 12975 9072
rect 13039 9008 13056 9072
rect 13120 9008 13137 9072
rect 13201 9008 13218 9072
rect 13282 9008 13299 9072
rect 13363 9008 13380 9072
rect 13444 9008 13461 9072
rect 13525 9008 13542 9072
rect 13606 9008 13623 9072
rect 13687 9008 13704 9072
rect 13768 9008 13785 9072
rect 13849 9008 13866 9072
rect 13930 9008 13947 9072
rect 14011 9008 14028 9072
rect 14092 9008 14109 9072
rect 14173 9008 14190 9072
rect 14254 9008 14271 9072
rect 14335 9008 14352 9072
rect 14416 9008 14433 9072
rect 14497 9008 14513 9072
rect 14577 9008 14593 9072
rect 14657 9008 14673 9072
rect 14737 9008 14753 9072
rect 14817 9008 14833 9072
rect 14897 9008 14913 9072
rect 14977 9008 14993 9072
rect 15057 9008 15073 9072
rect 15137 9008 15153 9072
rect 15217 9008 15233 9072
rect 15297 9008 15313 9072
rect 15377 9008 15393 9072
rect 15457 9008 15473 9072
rect 15537 9008 15553 9072
rect 15617 9008 15623 9072
rect 12159 8986 15623 9008
rect 12159 8922 12165 8986
rect 12229 8922 12246 8986
rect 12310 8922 12327 8986
rect 12391 8922 12408 8986
rect 12472 8922 12489 8986
rect 12553 8922 12570 8986
rect 12634 8922 12651 8986
rect 12715 8922 12732 8986
rect 12796 8922 12813 8986
rect 12877 8922 12894 8986
rect 12958 8922 12975 8986
rect 13039 8922 13056 8986
rect 13120 8922 13137 8986
rect 13201 8922 13218 8986
rect 13282 8922 13299 8986
rect 13363 8922 13380 8986
rect 13444 8922 13461 8986
rect 13525 8922 13542 8986
rect 13606 8922 13623 8986
rect 13687 8922 13704 8986
rect 13768 8922 13785 8986
rect 13849 8922 13866 8986
rect 13930 8922 13947 8986
rect 14011 8922 14028 8986
rect 14092 8922 14109 8986
rect 14173 8922 14190 8986
rect 14254 8922 14271 8986
rect 14335 8922 14352 8986
rect 14416 8922 14433 8986
rect 14497 8922 14513 8986
rect 14577 8922 14593 8986
rect 14657 8922 14673 8986
rect 14737 8922 14753 8986
rect 14817 8922 14833 8986
rect 14897 8922 14913 8986
rect 14977 8922 14993 8986
rect 15057 8922 15073 8986
rect 15137 8922 15153 8986
rect 15217 8922 15233 8986
rect 15297 8922 15313 8986
rect 15377 8922 15393 8986
rect 15457 8922 15473 8986
rect 15537 8922 15553 8986
rect 15617 8922 15623 8986
rect 12159 8900 15623 8922
rect 12159 8836 12165 8900
rect 12229 8836 12246 8900
rect 12310 8836 12327 8900
rect 12391 8836 12408 8900
rect 12472 8836 12489 8900
rect 12553 8836 12570 8900
rect 12634 8836 12651 8900
rect 12715 8836 12732 8900
rect 12796 8836 12813 8900
rect 12877 8836 12894 8900
rect 12958 8836 12975 8900
rect 13039 8836 13056 8900
rect 13120 8836 13137 8900
rect 13201 8836 13218 8900
rect 13282 8836 13299 8900
rect 13363 8836 13380 8900
rect 13444 8836 13461 8900
rect 13525 8836 13542 8900
rect 13606 8836 13623 8900
rect 13687 8836 13704 8900
rect 13768 8836 13785 8900
rect 13849 8836 13866 8900
rect 13930 8836 13947 8900
rect 14011 8836 14028 8900
rect 14092 8836 14109 8900
rect 14173 8836 14190 8900
rect 14254 8836 14271 8900
rect 14335 8836 14352 8900
rect 14416 8836 14433 8900
rect 14497 8836 14513 8900
rect 14577 8836 14593 8900
rect 14657 8836 14673 8900
rect 14737 8836 14753 8900
rect 14817 8836 14833 8900
rect 14897 8836 14913 8900
rect 14977 8836 14993 8900
rect 15057 8836 15073 8900
rect 15137 8836 15153 8900
rect 15217 8836 15233 8900
rect 15297 8836 15313 8900
rect 15377 8836 15393 8900
rect 15457 8836 15473 8900
rect 15537 8836 15553 8900
rect 15617 8836 15623 8900
rect 12159 8814 15623 8836
rect 12159 8750 12165 8814
rect 12229 8750 12246 8814
rect 12310 8750 12327 8814
rect 12391 8750 12408 8814
rect 12472 8750 12489 8814
rect 12553 8750 12570 8814
rect 12634 8750 12651 8814
rect 12715 8750 12732 8814
rect 12796 8750 12813 8814
rect 12877 8750 12894 8814
rect 12958 8750 12975 8814
rect 13039 8750 13056 8814
rect 13120 8750 13137 8814
rect 13201 8750 13218 8814
rect 13282 8750 13299 8814
rect 13363 8750 13380 8814
rect 13444 8750 13461 8814
rect 13525 8750 13542 8814
rect 13606 8750 13623 8814
rect 13687 8750 13704 8814
rect 13768 8750 13785 8814
rect 13849 8750 13866 8814
rect 13930 8750 13947 8814
rect 14011 8750 14028 8814
rect 14092 8750 14109 8814
rect 14173 8750 14190 8814
rect 14254 8750 14271 8814
rect 14335 8750 14352 8814
rect 14416 8750 14433 8814
rect 14497 8750 14513 8814
rect 14577 8750 14593 8814
rect 14657 8750 14673 8814
rect 14737 8750 14753 8814
rect 14817 8750 14833 8814
rect 14897 8750 14913 8814
rect 14977 8750 14993 8814
rect 15057 8750 15073 8814
rect 15137 8750 15153 8814
rect 15217 8750 15233 8814
rect 15297 8750 15313 8814
rect 15377 8750 15393 8814
rect 15457 8750 15473 8814
rect 15537 8750 15553 8814
rect 15617 8750 15623 8814
rect 12159 8728 15623 8750
rect 12159 8664 12165 8728
rect 12229 8664 12246 8728
rect 12310 8664 12327 8728
rect 12391 8664 12408 8728
rect 12472 8664 12489 8728
rect 12553 8664 12570 8728
rect 12634 8664 12651 8728
rect 12715 8664 12732 8728
rect 12796 8664 12813 8728
rect 12877 8664 12894 8728
rect 12958 8664 12975 8728
rect 13039 8664 13056 8728
rect 13120 8664 13137 8728
rect 13201 8664 13218 8728
rect 13282 8664 13299 8728
rect 13363 8664 13380 8728
rect 13444 8664 13461 8728
rect 13525 8664 13542 8728
rect 13606 8664 13623 8728
rect 13687 8664 13704 8728
rect 13768 8664 13785 8728
rect 13849 8664 13866 8728
rect 13930 8664 13947 8728
rect 14011 8664 14028 8728
rect 14092 8664 14109 8728
rect 14173 8664 14190 8728
rect 14254 8664 14271 8728
rect 14335 8664 14352 8728
rect 14416 8664 14433 8728
rect 14497 8664 14513 8728
rect 14577 8664 14593 8728
rect 14657 8664 14673 8728
rect 14737 8664 14753 8728
rect 14817 8664 14833 8728
rect 14897 8664 14913 8728
rect 14977 8664 14993 8728
rect 15057 8664 15073 8728
rect 15137 8664 15153 8728
rect 15217 8664 15233 8728
rect 15297 8664 15313 8728
rect 15377 8664 15393 8728
rect 15457 8664 15473 8728
rect 15537 8664 15553 8728
rect 15617 8664 15623 8728
rect 12159 8642 15623 8664
rect 12159 8578 12165 8642
rect 12229 8578 12246 8642
rect 12310 8578 12327 8642
rect 12391 8578 12408 8642
rect 12472 8578 12489 8642
rect 12553 8578 12570 8642
rect 12634 8578 12651 8642
rect 12715 8578 12732 8642
rect 12796 8578 12813 8642
rect 12877 8578 12894 8642
rect 12958 8578 12975 8642
rect 13039 8578 13056 8642
rect 13120 8578 13137 8642
rect 13201 8578 13218 8642
rect 13282 8578 13299 8642
rect 13363 8578 13380 8642
rect 13444 8578 13461 8642
rect 13525 8578 13542 8642
rect 13606 8578 13623 8642
rect 13687 8578 13704 8642
rect 13768 8578 13785 8642
rect 13849 8578 13866 8642
rect 13930 8578 13947 8642
rect 14011 8578 14028 8642
rect 14092 8578 14109 8642
rect 14173 8578 14190 8642
rect 14254 8578 14271 8642
rect 14335 8578 14352 8642
rect 14416 8578 14433 8642
rect 14497 8578 14513 8642
rect 14577 8578 14593 8642
rect 14657 8578 14673 8642
rect 14737 8578 14753 8642
rect 14817 8578 14833 8642
rect 14897 8578 14913 8642
rect 14977 8578 14993 8642
rect 15057 8578 15073 8642
rect 15137 8578 15153 8642
rect 15217 8578 15233 8642
rect 15297 8578 15313 8642
rect 15377 8578 15393 8642
rect 15457 8578 15473 8642
rect 15537 8578 15553 8642
rect 15617 8578 15623 8642
rect 12159 8556 15623 8578
rect 12159 8492 12165 8556
rect 12229 8492 12246 8556
rect 12310 8492 12327 8556
rect 12391 8492 12408 8556
rect 12472 8492 12489 8556
rect 12553 8492 12570 8556
rect 12634 8492 12651 8556
rect 12715 8492 12732 8556
rect 12796 8492 12813 8556
rect 12877 8492 12894 8556
rect 12958 8492 12975 8556
rect 13039 8492 13056 8556
rect 13120 8492 13137 8556
rect 13201 8492 13218 8556
rect 13282 8492 13299 8556
rect 13363 8492 13380 8556
rect 13444 8492 13461 8556
rect 13525 8492 13542 8556
rect 13606 8492 13623 8556
rect 13687 8492 13704 8556
rect 13768 8492 13785 8556
rect 13849 8492 13866 8556
rect 13930 8492 13947 8556
rect 14011 8492 14028 8556
rect 14092 8492 14109 8556
rect 14173 8492 14190 8556
rect 14254 8492 14271 8556
rect 14335 8492 14352 8556
rect 14416 8492 14433 8556
rect 14497 8492 14513 8556
rect 14577 8492 14593 8556
rect 14657 8492 14673 8556
rect 14737 8492 14753 8556
rect 14817 8492 14833 8556
rect 14897 8492 14913 8556
rect 14977 8492 14993 8556
rect 15057 8492 15073 8556
rect 15137 8492 15153 8556
rect 15217 8492 15233 8556
rect 15297 8492 15313 8556
rect 15377 8492 15393 8556
rect 15457 8492 15473 8556
rect 15537 8492 15553 8556
rect 15617 8492 15623 8556
rect 12159 8470 15623 8492
rect 12159 8406 12165 8470
rect 12229 8406 12246 8470
rect 12310 8406 12327 8470
rect 12391 8406 12408 8470
rect 12472 8406 12489 8470
rect 12553 8406 12570 8470
rect 12634 8406 12651 8470
rect 12715 8406 12732 8470
rect 12796 8406 12813 8470
rect 12877 8406 12894 8470
rect 12958 8406 12975 8470
rect 13039 8406 13056 8470
rect 13120 8406 13137 8470
rect 13201 8406 13218 8470
rect 13282 8406 13299 8470
rect 13363 8406 13380 8470
rect 13444 8406 13461 8470
rect 13525 8406 13542 8470
rect 13606 8406 13623 8470
rect 13687 8406 13704 8470
rect 13768 8406 13785 8470
rect 13849 8406 13866 8470
rect 13930 8406 13947 8470
rect 14011 8406 14028 8470
rect 14092 8406 14109 8470
rect 14173 8406 14190 8470
rect 14254 8406 14271 8470
rect 14335 8406 14352 8470
rect 14416 8406 14433 8470
rect 14497 8406 14513 8470
rect 14577 8406 14593 8470
rect 14657 8406 14673 8470
rect 14737 8406 14753 8470
rect 14817 8406 14833 8470
rect 14897 8406 14913 8470
rect 14977 8406 14993 8470
rect 15057 8406 15073 8470
rect 15137 8406 15153 8470
rect 15217 8406 15233 8470
rect 15297 8406 15313 8470
rect 15377 8406 15393 8470
rect 15457 8406 15473 8470
rect 15537 8406 15553 8470
rect 15617 8406 15623 8470
rect 12159 8384 15623 8406
rect 12159 8320 12165 8384
rect 12229 8320 12246 8384
rect 12310 8320 12327 8384
rect 12391 8320 12408 8384
rect 12472 8320 12489 8384
rect 12553 8320 12570 8384
rect 12634 8320 12651 8384
rect 12715 8320 12732 8384
rect 12796 8320 12813 8384
rect 12877 8320 12894 8384
rect 12958 8320 12975 8384
rect 13039 8320 13056 8384
rect 13120 8320 13137 8384
rect 13201 8320 13218 8384
rect 13282 8320 13299 8384
rect 13363 8320 13380 8384
rect 13444 8320 13461 8384
rect 13525 8320 13542 8384
rect 13606 8320 13623 8384
rect 13687 8320 13704 8384
rect 13768 8320 13785 8384
rect 13849 8320 13866 8384
rect 13930 8320 13947 8384
rect 14011 8320 14028 8384
rect 14092 8320 14109 8384
rect 14173 8320 14190 8384
rect 14254 8320 14271 8384
rect 14335 8320 14352 8384
rect 14416 8320 14433 8384
rect 14497 8320 14513 8384
rect 14577 8320 14593 8384
rect 14657 8320 14673 8384
rect 14737 8320 14753 8384
rect 14817 8320 14833 8384
rect 14897 8320 14913 8384
rect 14977 8320 14993 8384
rect 15057 8320 15073 8384
rect 15137 8320 15153 8384
rect 15217 8320 15233 8384
rect 15297 8320 15313 8384
rect 15377 8320 15393 8384
rect 15457 8320 15473 8384
rect 15537 8320 15553 8384
rect 15617 8320 15623 8384
rect 11637 2701 11775 2707
rect 11637 2637 11674 2701
rect 11738 2637 11775 2701
rect 11637 2579 11775 2637
rect 11637 2515 11674 2579
rect 11738 2515 11775 2579
rect 11637 2457 11775 2515
rect 11637 2393 11674 2457
rect 11738 2393 11775 2457
rect 11637 2335 11775 2393
rect 11637 2271 11674 2335
rect 11738 2271 11775 2335
rect 11637 2213 11775 2271
rect 11637 2149 11674 2213
rect 11738 2149 11775 2213
rect 11637 2091 11775 2149
rect 11637 2027 11674 2091
rect 11738 2027 11775 2091
rect 11637 1969 11775 2027
rect 11637 1905 11674 1969
rect 11738 1905 11775 1969
rect 11637 1847 11775 1905
rect 11637 1783 11674 1847
rect 11738 1783 11775 1847
rect 11637 1777 11775 1783
rect 8853 784 8863 840
rect 8919 784 8944 840
rect 9000 784 9025 840
rect 9081 784 9106 840
rect 9162 784 9187 840
rect 9243 784 9268 840
rect 9324 784 9349 840
rect 9405 784 9430 840
rect 9486 784 9510 840
rect 9566 784 9590 840
rect 9646 784 11082 840
rect 8853 0 11082 784
rect 12159 0 15623 8320
<< via3 >>
rect 397 9180 461 9244
rect 479 9180 543 9244
rect 561 9180 625 9244
rect 643 9180 707 9244
rect 725 9180 789 9244
rect 807 9180 871 9244
rect 889 9180 953 9244
rect 971 9180 1035 9244
rect 1053 9180 1117 9244
rect 1135 9180 1199 9244
rect 1217 9180 1281 9244
rect 1299 9180 1363 9244
rect 1381 9180 1445 9244
rect 1463 9180 1527 9244
rect 1545 9180 1609 9244
rect 1627 9180 1691 9244
rect 1709 9180 1773 9244
rect 1791 9180 1855 9244
rect 1873 9180 1937 9244
rect 1955 9180 2019 9244
rect 2037 9180 2101 9244
rect 2119 9180 2183 9244
rect 2201 9180 2265 9244
rect 2282 9180 2346 9244
rect 2363 9180 2427 9244
rect 397 9094 461 9158
rect 479 9094 543 9158
rect 561 9094 625 9158
rect 643 9094 707 9158
rect 725 9094 789 9158
rect 807 9094 871 9158
rect 889 9094 953 9158
rect 971 9094 1035 9158
rect 1053 9094 1117 9158
rect 1135 9094 1199 9158
rect 1217 9094 1281 9158
rect 1299 9094 1363 9158
rect 1381 9094 1445 9158
rect 1463 9094 1527 9158
rect 1545 9094 1609 9158
rect 1627 9094 1691 9158
rect 1709 9094 1773 9158
rect 1791 9094 1855 9158
rect 1873 9094 1937 9158
rect 1955 9094 2019 9158
rect 2037 9094 2101 9158
rect 2119 9094 2183 9158
rect 2201 9094 2265 9158
rect 2282 9094 2346 9158
rect 2363 9094 2427 9158
rect 397 9008 461 9072
rect 479 9008 543 9072
rect 561 9008 625 9072
rect 643 9008 707 9072
rect 725 9008 789 9072
rect 807 9008 871 9072
rect 889 9008 953 9072
rect 971 9008 1035 9072
rect 1053 9008 1117 9072
rect 1135 9008 1199 9072
rect 1217 9008 1281 9072
rect 1299 9008 1363 9072
rect 1381 9008 1445 9072
rect 1463 9008 1527 9072
rect 1545 9008 1609 9072
rect 1627 9008 1691 9072
rect 1709 9008 1773 9072
rect 1791 9008 1855 9072
rect 1873 9008 1937 9072
rect 1955 9008 2019 9072
rect 2037 9008 2101 9072
rect 2119 9008 2183 9072
rect 2201 9008 2265 9072
rect 2282 9008 2346 9072
rect 2363 9008 2427 9072
rect 397 8922 461 8986
rect 479 8922 543 8986
rect 561 8922 625 8986
rect 643 8922 707 8986
rect 725 8922 789 8986
rect 807 8922 871 8986
rect 889 8922 953 8986
rect 971 8922 1035 8986
rect 1053 8922 1117 8986
rect 1135 8922 1199 8986
rect 1217 8922 1281 8986
rect 1299 8922 1363 8986
rect 1381 8922 1445 8986
rect 1463 8922 1527 8986
rect 1545 8922 1609 8986
rect 1627 8922 1691 8986
rect 1709 8922 1773 8986
rect 1791 8922 1855 8986
rect 1873 8922 1937 8986
rect 1955 8922 2019 8986
rect 2037 8922 2101 8986
rect 2119 8922 2183 8986
rect 2201 8922 2265 8986
rect 2282 8922 2346 8986
rect 2363 8922 2427 8986
rect 397 8836 461 8900
rect 479 8836 543 8900
rect 561 8836 625 8900
rect 643 8836 707 8900
rect 725 8836 789 8900
rect 807 8836 871 8900
rect 889 8836 953 8900
rect 971 8836 1035 8900
rect 1053 8836 1117 8900
rect 1135 8836 1199 8900
rect 1217 8836 1281 8900
rect 1299 8836 1363 8900
rect 1381 8836 1445 8900
rect 1463 8836 1527 8900
rect 1545 8836 1609 8900
rect 1627 8836 1691 8900
rect 1709 8836 1773 8900
rect 1791 8836 1855 8900
rect 1873 8836 1937 8900
rect 1955 8836 2019 8900
rect 2037 8836 2101 8900
rect 2119 8836 2183 8900
rect 2201 8836 2265 8900
rect 2282 8836 2346 8900
rect 2363 8836 2427 8900
rect 397 8750 461 8814
rect 479 8750 543 8814
rect 561 8750 625 8814
rect 643 8750 707 8814
rect 725 8750 789 8814
rect 807 8750 871 8814
rect 889 8750 953 8814
rect 971 8750 1035 8814
rect 1053 8750 1117 8814
rect 1135 8750 1199 8814
rect 1217 8750 1281 8814
rect 1299 8750 1363 8814
rect 1381 8750 1445 8814
rect 1463 8750 1527 8814
rect 1545 8750 1609 8814
rect 1627 8750 1691 8814
rect 1709 8750 1773 8814
rect 1791 8750 1855 8814
rect 1873 8750 1937 8814
rect 1955 8750 2019 8814
rect 2037 8750 2101 8814
rect 2119 8750 2183 8814
rect 2201 8750 2265 8814
rect 2282 8750 2346 8814
rect 2363 8750 2427 8814
rect 397 8664 461 8728
rect 479 8664 543 8728
rect 561 8664 625 8728
rect 643 8664 707 8728
rect 725 8664 789 8728
rect 807 8664 871 8728
rect 889 8664 953 8728
rect 971 8664 1035 8728
rect 1053 8664 1117 8728
rect 1135 8664 1199 8728
rect 1217 8664 1281 8728
rect 1299 8664 1363 8728
rect 1381 8664 1445 8728
rect 1463 8664 1527 8728
rect 1545 8664 1609 8728
rect 1627 8664 1691 8728
rect 1709 8664 1773 8728
rect 1791 8664 1855 8728
rect 1873 8664 1937 8728
rect 1955 8664 2019 8728
rect 2037 8664 2101 8728
rect 2119 8664 2183 8728
rect 2201 8664 2265 8728
rect 2282 8664 2346 8728
rect 2363 8664 2427 8728
rect 397 8578 461 8642
rect 479 8578 543 8642
rect 561 8578 625 8642
rect 643 8578 707 8642
rect 725 8578 789 8642
rect 807 8578 871 8642
rect 889 8578 953 8642
rect 971 8578 1035 8642
rect 1053 8578 1117 8642
rect 1135 8578 1199 8642
rect 1217 8578 1281 8642
rect 1299 8578 1363 8642
rect 1381 8578 1445 8642
rect 1463 8578 1527 8642
rect 1545 8578 1609 8642
rect 1627 8578 1691 8642
rect 1709 8578 1773 8642
rect 1791 8578 1855 8642
rect 1873 8578 1937 8642
rect 1955 8578 2019 8642
rect 2037 8578 2101 8642
rect 2119 8578 2183 8642
rect 2201 8578 2265 8642
rect 2282 8578 2346 8642
rect 2363 8578 2427 8642
rect 397 8492 461 8556
rect 479 8492 543 8556
rect 561 8492 625 8556
rect 643 8492 707 8556
rect 725 8492 789 8556
rect 807 8492 871 8556
rect 889 8492 953 8556
rect 971 8492 1035 8556
rect 1053 8492 1117 8556
rect 1135 8492 1199 8556
rect 1217 8492 1281 8556
rect 1299 8492 1363 8556
rect 1381 8492 1445 8556
rect 1463 8492 1527 8556
rect 1545 8492 1609 8556
rect 1627 8492 1691 8556
rect 1709 8492 1773 8556
rect 1791 8492 1855 8556
rect 1873 8492 1937 8556
rect 1955 8492 2019 8556
rect 2037 8492 2101 8556
rect 2119 8492 2183 8556
rect 2201 8492 2265 8556
rect 2282 8492 2346 8556
rect 2363 8492 2427 8556
rect 397 8406 461 8470
rect 479 8406 543 8470
rect 561 8406 625 8470
rect 643 8406 707 8470
rect 725 8406 789 8470
rect 807 8406 871 8470
rect 889 8406 953 8470
rect 971 8406 1035 8470
rect 1053 8406 1117 8470
rect 1135 8406 1199 8470
rect 1217 8406 1281 8470
rect 1299 8406 1363 8470
rect 1381 8406 1445 8470
rect 1463 8406 1527 8470
rect 1545 8406 1609 8470
rect 1627 8406 1691 8470
rect 1709 8406 1773 8470
rect 1791 8406 1855 8470
rect 1873 8406 1937 8470
rect 1955 8406 2019 8470
rect 2037 8406 2101 8470
rect 2119 8406 2183 8470
rect 2201 8406 2265 8470
rect 2282 8406 2346 8470
rect 2363 8406 2427 8470
rect 397 8320 461 8384
rect 479 8320 543 8384
rect 561 8320 625 8384
rect 643 8320 707 8384
rect 725 8320 789 8384
rect 807 8320 871 8384
rect 889 8320 953 8384
rect 971 8320 1035 8384
rect 1053 8320 1117 8384
rect 1135 8320 1199 8384
rect 1217 8320 1281 8384
rect 1299 8320 1363 8384
rect 1381 8320 1445 8384
rect 1463 8320 1527 8384
rect 1545 8320 1609 8384
rect 1627 8320 1691 8384
rect 1709 8320 1773 8384
rect 1791 8320 1855 8384
rect 1873 8320 1937 8384
rect 1955 8320 2019 8384
rect 2037 8320 2101 8384
rect 2119 8320 2183 8384
rect 2201 8320 2265 8384
rect 2282 8320 2346 8384
rect 2363 8320 2427 8384
rect 547 2698 611 2701
rect 547 2642 548 2698
rect 548 2642 604 2698
rect 604 2642 611 2698
rect 547 2637 611 2642
rect 659 2698 723 2701
rect 659 2642 662 2698
rect 662 2642 718 2698
rect 718 2642 723 2698
rect 659 2637 723 2642
rect 771 2698 835 2701
rect 771 2642 776 2698
rect 776 2642 832 2698
rect 832 2642 835 2698
rect 771 2637 835 2642
rect 883 2698 947 2701
rect 883 2642 890 2698
rect 890 2642 946 2698
rect 946 2642 947 2698
rect 883 2637 947 2642
rect 547 2576 611 2579
rect 547 2520 548 2576
rect 548 2520 604 2576
rect 604 2520 611 2576
rect 547 2515 611 2520
rect 659 2576 723 2579
rect 659 2520 662 2576
rect 662 2520 718 2576
rect 718 2520 723 2576
rect 659 2515 723 2520
rect 771 2576 835 2579
rect 771 2520 776 2576
rect 776 2520 832 2576
rect 832 2520 835 2576
rect 771 2515 835 2520
rect 883 2576 947 2579
rect 883 2520 890 2576
rect 890 2520 946 2576
rect 946 2520 947 2576
rect 883 2515 947 2520
rect 547 2454 611 2457
rect 547 2398 548 2454
rect 548 2398 604 2454
rect 604 2398 611 2454
rect 547 2393 611 2398
rect 659 2454 723 2457
rect 659 2398 662 2454
rect 662 2398 718 2454
rect 718 2398 723 2454
rect 659 2393 723 2398
rect 771 2454 835 2457
rect 771 2398 776 2454
rect 776 2398 832 2454
rect 832 2398 835 2454
rect 771 2393 835 2398
rect 883 2454 947 2457
rect 883 2398 890 2454
rect 890 2398 946 2454
rect 946 2398 947 2454
rect 883 2393 947 2398
rect 547 2332 611 2335
rect 547 2276 548 2332
rect 548 2276 604 2332
rect 604 2276 611 2332
rect 547 2271 611 2276
rect 659 2332 723 2335
rect 659 2276 662 2332
rect 662 2276 718 2332
rect 718 2276 723 2332
rect 659 2271 723 2276
rect 771 2332 835 2335
rect 771 2276 776 2332
rect 776 2276 832 2332
rect 832 2276 835 2332
rect 771 2271 835 2276
rect 883 2332 947 2335
rect 883 2276 890 2332
rect 890 2276 946 2332
rect 946 2276 947 2332
rect 883 2271 947 2276
rect 547 2210 611 2213
rect 547 2154 548 2210
rect 548 2154 604 2210
rect 604 2154 611 2210
rect 547 2149 611 2154
rect 659 2210 723 2213
rect 659 2154 662 2210
rect 662 2154 718 2210
rect 718 2154 723 2210
rect 659 2149 723 2154
rect 771 2210 835 2213
rect 771 2154 776 2210
rect 776 2154 832 2210
rect 832 2154 835 2210
rect 771 2149 835 2154
rect 883 2210 947 2213
rect 883 2154 890 2210
rect 890 2154 946 2210
rect 946 2154 947 2210
rect 883 2149 947 2154
rect 547 2088 611 2091
rect 547 2032 548 2088
rect 548 2032 604 2088
rect 604 2032 611 2088
rect 547 2027 611 2032
rect 659 2088 723 2091
rect 659 2032 662 2088
rect 662 2032 718 2088
rect 718 2032 723 2088
rect 659 2027 723 2032
rect 771 2088 835 2091
rect 771 2032 776 2088
rect 776 2032 832 2088
rect 832 2032 835 2088
rect 771 2027 835 2032
rect 883 2088 947 2091
rect 883 2032 890 2088
rect 890 2032 946 2088
rect 946 2032 947 2088
rect 883 2027 947 2032
rect 547 1965 611 1969
rect 547 1909 548 1965
rect 548 1909 604 1965
rect 604 1909 611 1965
rect 547 1905 611 1909
rect 659 1965 723 1969
rect 659 1909 662 1965
rect 662 1909 718 1965
rect 718 1909 723 1965
rect 659 1905 723 1909
rect 771 1965 835 1969
rect 771 1909 776 1965
rect 776 1909 832 1965
rect 832 1909 835 1965
rect 771 1905 835 1909
rect 883 1965 947 1969
rect 883 1909 890 1965
rect 890 1909 946 1965
rect 946 1909 947 1965
rect 883 1905 947 1909
rect 547 1842 611 1847
rect 547 1786 548 1842
rect 548 1786 604 1842
rect 604 1786 611 1842
rect 547 1783 611 1786
rect 659 1842 723 1847
rect 659 1786 662 1842
rect 662 1786 718 1842
rect 718 1786 723 1842
rect 659 1783 723 1786
rect 771 1842 835 1847
rect 771 1786 776 1842
rect 776 1786 832 1842
rect 832 1786 835 1842
rect 771 1783 835 1786
rect 883 1842 947 1847
rect 883 1786 890 1842
rect 890 1786 946 1842
rect 946 1786 947 1842
rect 883 1783 947 1786
rect 2553 9180 2617 9244
rect 2635 9180 2699 9244
rect 2717 9180 2781 9244
rect 2799 9180 2863 9244
rect 2881 9180 2945 9244
rect 2963 9180 3027 9244
rect 3045 9180 3109 9244
rect 3127 9180 3191 9244
rect 3209 9180 3273 9244
rect 3290 9180 3354 9244
rect 3371 9180 3435 9244
rect 3452 9180 3516 9244
rect 3533 9180 3597 9244
rect 3614 9180 3678 9244
rect 3695 9180 3759 9244
rect 3776 9180 3840 9244
rect 3857 9180 3921 9244
rect 3938 9180 4002 9244
rect 4019 9180 4083 9244
rect 4100 9180 4164 9244
rect 4181 9180 4245 9244
rect 4262 9180 4326 9244
rect 4343 9180 4407 9244
rect 4424 9180 4488 9244
rect 4505 9180 4569 9244
rect 2553 9094 2617 9158
rect 2635 9094 2699 9158
rect 2717 9094 2781 9158
rect 2799 9094 2863 9158
rect 2881 9094 2945 9158
rect 2963 9094 3027 9158
rect 3045 9094 3109 9158
rect 3127 9094 3191 9158
rect 3209 9094 3273 9158
rect 3290 9094 3354 9158
rect 3371 9094 3435 9158
rect 3452 9094 3516 9158
rect 3533 9094 3597 9158
rect 3614 9094 3678 9158
rect 3695 9094 3759 9158
rect 3776 9094 3840 9158
rect 3857 9094 3921 9158
rect 3938 9094 4002 9158
rect 4019 9094 4083 9158
rect 4100 9094 4164 9158
rect 4181 9094 4245 9158
rect 4262 9094 4326 9158
rect 4343 9094 4407 9158
rect 4424 9094 4488 9158
rect 4505 9094 4569 9158
rect 2553 9008 2617 9072
rect 2635 9008 2699 9072
rect 2717 9008 2781 9072
rect 2799 9008 2863 9072
rect 2881 9008 2945 9072
rect 2963 9008 3027 9072
rect 3045 9008 3109 9072
rect 3127 9008 3191 9072
rect 3209 9008 3273 9072
rect 3290 9008 3354 9072
rect 3371 9008 3435 9072
rect 3452 9008 3516 9072
rect 3533 9008 3597 9072
rect 3614 9008 3678 9072
rect 3695 9008 3759 9072
rect 3776 9008 3840 9072
rect 3857 9008 3921 9072
rect 3938 9008 4002 9072
rect 4019 9008 4083 9072
rect 4100 9008 4164 9072
rect 4181 9008 4245 9072
rect 4262 9008 4326 9072
rect 4343 9008 4407 9072
rect 4424 9008 4488 9072
rect 4505 9008 4569 9072
rect 2553 8922 2617 8986
rect 2635 8922 2699 8986
rect 2717 8922 2781 8986
rect 2799 8922 2863 8986
rect 2881 8922 2945 8986
rect 2963 8922 3027 8986
rect 3045 8922 3109 8986
rect 3127 8922 3191 8986
rect 3209 8922 3273 8986
rect 3290 8922 3354 8986
rect 3371 8922 3435 8986
rect 3452 8922 3516 8986
rect 3533 8922 3597 8986
rect 3614 8922 3678 8986
rect 3695 8922 3759 8986
rect 3776 8922 3840 8986
rect 3857 8922 3921 8986
rect 3938 8922 4002 8986
rect 4019 8922 4083 8986
rect 4100 8922 4164 8986
rect 4181 8922 4245 8986
rect 4262 8922 4326 8986
rect 4343 8922 4407 8986
rect 4424 8922 4488 8986
rect 4505 8922 4569 8986
rect 2553 8836 2617 8900
rect 2635 8836 2699 8900
rect 2717 8836 2781 8900
rect 2799 8836 2863 8900
rect 2881 8836 2945 8900
rect 2963 8836 3027 8900
rect 3045 8836 3109 8900
rect 3127 8836 3191 8900
rect 3209 8836 3273 8900
rect 3290 8836 3354 8900
rect 3371 8836 3435 8900
rect 3452 8836 3516 8900
rect 3533 8836 3597 8900
rect 3614 8836 3678 8900
rect 3695 8836 3759 8900
rect 3776 8836 3840 8900
rect 3857 8836 3921 8900
rect 3938 8836 4002 8900
rect 4019 8836 4083 8900
rect 4100 8836 4164 8900
rect 4181 8836 4245 8900
rect 4262 8836 4326 8900
rect 4343 8836 4407 8900
rect 4424 8836 4488 8900
rect 4505 8836 4569 8900
rect 2553 8750 2617 8814
rect 2635 8750 2699 8814
rect 2717 8750 2781 8814
rect 2799 8750 2863 8814
rect 2881 8750 2945 8814
rect 2963 8750 3027 8814
rect 3045 8750 3109 8814
rect 3127 8750 3191 8814
rect 3209 8750 3273 8814
rect 3290 8750 3354 8814
rect 3371 8750 3435 8814
rect 3452 8750 3516 8814
rect 3533 8750 3597 8814
rect 3614 8750 3678 8814
rect 3695 8750 3759 8814
rect 3776 8750 3840 8814
rect 3857 8750 3921 8814
rect 3938 8750 4002 8814
rect 4019 8750 4083 8814
rect 4100 8750 4164 8814
rect 4181 8750 4245 8814
rect 4262 8750 4326 8814
rect 4343 8750 4407 8814
rect 4424 8750 4488 8814
rect 4505 8750 4569 8814
rect 2553 8664 2617 8728
rect 2635 8664 2699 8728
rect 2717 8664 2781 8728
rect 2799 8664 2863 8728
rect 2881 8664 2945 8728
rect 2963 8664 3027 8728
rect 3045 8664 3109 8728
rect 3127 8664 3191 8728
rect 3209 8664 3273 8728
rect 3290 8664 3354 8728
rect 3371 8664 3435 8728
rect 3452 8664 3516 8728
rect 3533 8664 3597 8728
rect 3614 8664 3678 8728
rect 3695 8664 3759 8728
rect 3776 8664 3840 8728
rect 3857 8664 3921 8728
rect 3938 8664 4002 8728
rect 4019 8664 4083 8728
rect 4100 8664 4164 8728
rect 4181 8664 4245 8728
rect 4262 8664 4326 8728
rect 4343 8664 4407 8728
rect 4424 8664 4488 8728
rect 4505 8664 4569 8728
rect 2553 8578 2617 8642
rect 2635 8578 2699 8642
rect 2717 8578 2781 8642
rect 2799 8578 2863 8642
rect 2881 8578 2945 8642
rect 2963 8578 3027 8642
rect 3045 8578 3109 8642
rect 3127 8578 3191 8642
rect 3209 8578 3273 8642
rect 3290 8578 3354 8642
rect 3371 8578 3435 8642
rect 3452 8578 3516 8642
rect 3533 8578 3597 8642
rect 3614 8578 3678 8642
rect 3695 8578 3759 8642
rect 3776 8578 3840 8642
rect 3857 8578 3921 8642
rect 3938 8578 4002 8642
rect 4019 8578 4083 8642
rect 4100 8578 4164 8642
rect 4181 8578 4245 8642
rect 4262 8578 4326 8642
rect 4343 8578 4407 8642
rect 4424 8578 4488 8642
rect 4505 8578 4569 8642
rect 2553 8492 2617 8556
rect 2635 8492 2699 8556
rect 2717 8492 2781 8556
rect 2799 8492 2863 8556
rect 2881 8492 2945 8556
rect 2963 8492 3027 8556
rect 3045 8492 3109 8556
rect 3127 8492 3191 8556
rect 3209 8492 3273 8556
rect 3290 8492 3354 8556
rect 3371 8492 3435 8556
rect 3452 8492 3516 8556
rect 3533 8492 3597 8556
rect 3614 8492 3678 8556
rect 3695 8492 3759 8556
rect 3776 8492 3840 8556
rect 3857 8492 3921 8556
rect 3938 8492 4002 8556
rect 4019 8492 4083 8556
rect 4100 8492 4164 8556
rect 4181 8492 4245 8556
rect 4262 8492 4326 8556
rect 4343 8492 4407 8556
rect 4424 8492 4488 8556
rect 4505 8492 4569 8556
rect 2553 8406 2617 8470
rect 2635 8406 2699 8470
rect 2717 8406 2781 8470
rect 2799 8406 2863 8470
rect 2881 8406 2945 8470
rect 2963 8406 3027 8470
rect 3045 8406 3109 8470
rect 3127 8406 3191 8470
rect 3209 8406 3273 8470
rect 3290 8406 3354 8470
rect 3371 8406 3435 8470
rect 3452 8406 3516 8470
rect 3533 8406 3597 8470
rect 3614 8406 3678 8470
rect 3695 8406 3759 8470
rect 3776 8406 3840 8470
rect 3857 8406 3921 8470
rect 3938 8406 4002 8470
rect 4019 8406 4083 8470
rect 4100 8406 4164 8470
rect 4181 8406 4245 8470
rect 4262 8406 4326 8470
rect 4343 8406 4407 8470
rect 4424 8406 4488 8470
rect 4505 8406 4569 8470
rect 2553 8320 2617 8384
rect 2635 8320 2699 8384
rect 2717 8320 2781 8384
rect 2799 8320 2863 8384
rect 2881 8320 2945 8384
rect 2963 8320 3027 8384
rect 3045 8320 3109 8384
rect 3127 8320 3191 8384
rect 3209 8320 3273 8384
rect 3290 8320 3354 8384
rect 3371 8320 3435 8384
rect 3452 8320 3516 8384
rect 3533 8320 3597 8384
rect 3614 8320 3678 8384
rect 3695 8320 3759 8384
rect 3776 8320 3840 8384
rect 3857 8320 3921 8384
rect 3938 8320 4002 8384
rect 4019 8320 4083 8384
rect 4100 8320 4164 8384
rect 4181 8320 4245 8384
rect 4262 8320 4326 8384
rect 4343 8320 4407 8384
rect 4424 8320 4488 8384
rect 4505 8320 4569 8384
rect 4695 9180 4759 9244
rect 4777 9180 4841 9244
rect 4859 9180 4923 9244
rect 4941 9180 5005 9244
rect 5023 9180 5087 9244
rect 5105 9180 5169 9244
rect 5187 9180 5251 9244
rect 5269 9180 5333 9244
rect 5351 9180 5415 9244
rect 5433 9180 5497 9244
rect 5515 9180 5579 9244
rect 5597 9180 5661 9244
rect 5679 9180 5743 9244
rect 5760 9180 5824 9244
rect 5841 9180 5905 9244
rect 5922 9180 5986 9244
rect 6003 9180 6067 9244
rect 6084 9180 6148 9244
rect 6165 9180 6229 9244
rect 6246 9180 6310 9244
rect 6327 9180 6391 9244
rect 6408 9180 6472 9244
rect 6489 9180 6553 9244
rect 6570 9180 6634 9244
rect 6651 9180 6715 9244
rect 6732 9180 6796 9244
rect 6813 9180 6877 9244
rect 6894 9180 6958 9244
rect 6975 9180 7039 9244
rect 7056 9180 7120 9244
rect 7137 9180 7201 9244
rect 7218 9180 7282 9244
rect 7299 9180 7363 9244
rect 7380 9180 7444 9244
rect 7461 9180 7525 9244
rect 7542 9180 7606 9244
rect 7623 9180 7687 9244
rect 4695 9094 4759 9158
rect 4777 9094 4841 9158
rect 4859 9094 4923 9158
rect 4941 9094 5005 9158
rect 5023 9094 5087 9158
rect 5105 9094 5169 9158
rect 5187 9094 5251 9158
rect 5269 9094 5333 9158
rect 5351 9094 5415 9158
rect 5433 9094 5497 9158
rect 5515 9094 5579 9158
rect 5597 9094 5661 9158
rect 5679 9094 5743 9158
rect 5760 9094 5824 9158
rect 5841 9094 5905 9158
rect 5922 9094 5986 9158
rect 6003 9094 6067 9158
rect 6084 9094 6148 9158
rect 6165 9094 6229 9158
rect 6246 9094 6310 9158
rect 6327 9094 6391 9158
rect 6408 9094 6472 9158
rect 6489 9094 6553 9158
rect 6570 9094 6634 9158
rect 6651 9094 6715 9158
rect 6732 9094 6796 9158
rect 6813 9094 6877 9158
rect 6894 9094 6958 9158
rect 6975 9094 7039 9158
rect 7056 9094 7120 9158
rect 7137 9094 7201 9158
rect 7218 9094 7282 9158
rect 7299 9094 7363 9158
rect 7380 9094 7444 9158
rect 7461 9094 7525 9158
rect 7542 9094 7606 9158
rect 7623 9094 7687 9158
rect 4695 9008 4759 9072
rect 4777 9008 4841 9072
rect 4859 9008 4923 9072
rect 4941 9008 5005 9072
rect 5023 9008 5087 9072
rect 5105 9008 5169 9072
rect 5187 9008 5251 9072
rect 5269 9008 5333 9072
rect 5351 9008 5415 9072
rect 5433 9008 5497 9072
rect 5515 9008 5579 9072
rect 5597 9008 5661 9072
rect 5679 9008 5743 9072
rect 5760 9008 5824 9072
rect 5841 9008 5905 9072
rect 5922 9008 5986 9072
rect 6003 9008 6067 9072
rect 6084 9008 6148 9072
rect 6165 9008 6229 9072
rect 6246 9008 6310 9072
rect 6327 9008 6391 9072
rect 6408 9008 6472 9072
rect 6489 9008 6553 9072
rect 6570 9008 6634 9072
rect 6651 9008 6715 9072
rect 6732 9008 6796 9072
rect 6813 9008 6877 9072
rect 6894 9008 6958 9072
rect 6975 9008 7039 9072
rect 7056 9008 7120 9072
rect 7137 9008 7201 9072
rect 7218 9008 7282 9072
rect 7299 9008 7363 9072
rect 7380 9008 7444 9072
rect 7461 9008 7525 9072
rect 7542 9008 7606 9072
rect 7623 9008 7687 9072
rect 4695 8922 4759 8986
rect 4777 8922 4841 8986
rect 4859 8922 4923 8986
rect 4941 8922 5005 8986
rect 5023 8922 5087 8986
rect 5105 8922 5169 8986
rect 5187 8922 5251 8986
rect 5269 8922 5333 8986
rect 5351 8922 5415 8986
rect 5433 8922 5497 8986
rect 5515 8922 5579 8986
rect 5597 8922 5661 8986
rect 5679 8922 5743 8986
rect 5760 8922 5824 8986
rect 5841 8922 5905 8986
rect 5922 8922 5986 8986
rect 6003 8922 6067 8986
rect 6084 8922 6148 8986
rect 6165 8922 6229 8986
rect 6246 8922 6310 8986
rect 6327 8922 6391 8986
rect 6408 8922 6472 8986
rect 6489 8922 6553 8986
rect 6570 8922 6634 8986
rect 6651 8922 6715 8986
rect 6732 8922 6796 8986
rect 6813 8922 6877 8986
rect 6894 8922 6958 8986
rect 6975 8922 7039 8986
rect 7056 8922 7120 8986
rect 7137 8922 7201 8986
rect 7218 8922 7282 8986
rect 7299 8922 7363 8986
rect 7380 8922 7444 8986
rect 7461 8922 7525 8986
rect 7542 8922 7606 8986
rect 7623 8922 7687 8986
rect 4695 8836 4759 8900
rect 4777 8836 4841 8900
rect 4859 8836 4923 8900
rect 4941 8836 5005 8900
rect 5023 8836 5087 8900
rect 5105 8836 5169 8900
rect 5187 8836 5251 8900
rect 5269 8836 5333 8900
rect 5351 8836 5415 8900
rect 5433 8836 5497 8900
rect 5515 8836 5579 8900
rect 5597 8836 5661 8900
rect 5679 8836 5743 8900
rect 5760 8836 5824 8900
rect 5841 8836 5905 8900
rect 5922 8836 5986 8900
rect 6003 8836 6067 8900
rect 6084 8836 6148 8900
rect 6165 8836 6229 8900
rect 6246 8836 6310 8900
rect 6327 8836 6391 8900
rect 6408 8836 6472 8900
rect 6489 8836 6553 8900
rect 6570 8836 6634 8900
rect 6651 8836 6715 8900
rect 6732 8836 6796 8900
rect 6813 8836 6877 8900
rect 6894 8836 6958 8900
rect 6975 8836 7039 8900
rect 7056 8836 7120 8900
rect 7137 8836 7201 8900
rect 7218 8836 7282 8900
rect 7299 8836 7363 8900
rect 7380 8836 7444 8900
rect 7461 8836 7525 8900
rect 7542 8836 7606 8900
rect 7623 8836 7687 8900
rect 4695 8750 4759 8814
rect 4777 8750 4841 8814
rect 4859 8750 4923 8814
rect 4941 8750 5005 8814
rect 5023 8750 5087 8814
rect 5105 8750 5169 8814
rect 5187 8750 5251 8814
rect 5269 8750 5333 8814
rect 5351 8750 5415 8814
rect 5433 8750 5497 8814
rect 5515 8750 5579 8814
rect 5597 8750 5661 8814
rect 5679 8750 5743 8814
rect 5760 8750 5824 8814
rect 5841 8750 5905 8814
rect 5922 8750 5986 8814
rect 6003 8750 6067 8814
rect 6084 8750 6148 8814
rect 6165 8750 6229 8814
rect 6246 8750 6310 8814
rect 6327 8750 6391 8814
rect 6408 8750 6472 8814
rect 6489 8750 6553 8814
rect 6570 8750 6634 8814
rect 6651 8750 6715 8814
rect 6732 8750 6796 8814
rect 6813 8750 6877 8814
rect 6894 8750 6958 8814
rect 6975 8750 7039 8814
rect 7056 8750 7120 8814
rect 7137 8750 7201 8814
rect 7218 8750 7282 8814
rect 7299 8750 7363 8814
rect 7380 8750 7444 8814
rect 7461 8750 7525 8814
rect 7542 8750 7606 8814
rect 7623 8750 7687 8814
rect 4695 8664 4759 8728
rect 4777 8664 4841 8728
rect 4859 8664 4923 8728
rect 4941 8664 5005 8728
rect 5023 8664 5087 8728
rect 5105 8664 5169 8728
rect 5187 8664 5251 8728
rect 5269 8664 5333 8728
rect 5351 8664 5415 8728
rect 5433 8664 5497 8728
rect 5515 8664 5579 8728
rect 5597 8664 5661 8728
rect 5679 8664 5743 8728
rect 5760 8664 5824 8728
rect 5841 8664 5905 8728
rect 5922 8664 5986 8728
rect 6003 8664 6067 8728
rect 6084 8664 6148 8728
rect 6165 8664 6229 8728
rect 6246 8664 6310 8728
rect 6327 8664 6391 8728
rect 6408 8664 6472 8728
rect 6489 8664 6553 8728
rect 6570 8664 6634 8728
rect 6651 8664 6715 8728
rect 6732 8664 6796 8728
rect 6813 8664 6877 8728
rect 6894 8664 6958 8728
rect 6975 8664 7039 8728
rect 7056 8664 7120 8728
rect 7137 8664 7201 8728
rect 7218 8664 7282 8728
rect 7299 8664 7363 8728
rect 7380 8664 7444 8728
rect 7461 8664 7525 8728
rect 7542 8664 7606 8728
rect 7623 8664 7687 8728
rect 4695 8578 4759 8642
rect 4777 8578 4841 8642
rect 4859 8578 4923 8642
rect 4941 8578 5005 8642
rect 5023 8578 5087 8642
rect 5105 8578 5169 8642
rect 5187 8578 5251 8642
rect 5269 8578 5333 8642
rect 5351 8578 5415 8642
rect 5433 8578 5497 8642
rect 5515 8578 5579 8642
rect 5597 8578 5661 8642
rect 5679 8578 5743 8642
rect 5760 8578 5824 8642
rect 5841 8578 5905 8642
rect 5922 8578 5986 8642
rect 6003 8578 6067 8642
rect 6084 8578 6148 8642
rect 6165 8578 6229 8642
rect 6246 8578 6310 8642
rect 6327 8578 6391 8642
rect 6408 8578 6472 8642
rect 6489 8578 6553 8642
rect 6570 8578 6634 8642
rect 6651 8578 6715 8642
rect 6732 8578 6796 8642
rect 6813 8578 6877 8642
rect 6894 8578 6958 8642
rect 6975 8578 7039 8642
rect 7056 8578 7120 8642
rect 7137 8578 7201 8642
rect 7218 8578 7282 8642
rect 7299 8578 7363 8642
rect 7380 8578 7444 8642
rect 7461 8578 7525 8642
rect 7542 8578 7606 8642
rect 7623 8578 7687 8642
rect 4695 8492 4759 8556
rect 4777 8492 4841 8556
rect 4859 8492 4923 8556
rect 4941 8492 5005 8556
rect 5023 8492 5087 8556
rect 5105 8492 5169 8556
rect 5187 8492 5251 8556
rect 5269 8492 5333 8556
rect 5351 8492 5415 8556
rect 5433 8492 5497 8556
rect 5515 8492 5579 8556
rect 5597 8492 5661 8556
rect 5679 8492 5743 8556
rect 5760 8492 5824 8556
rect 5841 8492 5905 8556
rect 5922 8492 5986 8556
rect 6003 8492 6067 8556
rect 6084 8492 6148 8556
rect 6165 8492 6229 8556
rect 6246 8492 6310 8556
rect 6327 8492 6391 8556
rect 6408 8492 6472 8556
rect 6489 8492 6553 8556
rect 6570 8492 6634 8556
rect 6651 8492 6715 8556
rect 6732 8492 6796 8556
rect 6813 8492 6877 8556
rect 6894 8492 6958 8556
rect 6975 8492 7039 8556
rect 7056 8492 7120 8556
rect 7137 8492 7201 8556
rect 7218 8492 7282 8556
rect 7299 8492 7363 8556
rect 7380 8492 7444 8556
rect 7461 8492 7525 8556
rect 7542 8492 7606 8556
rect 7623 8492 7687 8556
rect 4695 8406 4759 8470
rect 4777 8406 4841 8470
rect 4859 8406 4923 8470
rect 4941 8406 5005 8470
rect 5023 8406 5087 8470
rect 5105 8406 5169 8470
rect 5187 8406 5251 8470
rect 5269 8406 5333 8470
rect 5351 8406 5415 8470
rect 5433 8406 5497 8470
rect 5515 8406 5579 8470
rect 5597 8406 5661 8470
rect 5679 8406 5743 8470
rect 5760 8406 5824 8470
rect 5841 8406 5905 8470
rect 5922 8406 5986 8470
rect 6003 8406 6067 8470
rect 6084 8406 6148 8470
rect 6165 8406 6229 8470
rect 6246 8406 6310 8470
rect 6327 8406 6391 8470
rect 6408 8406 6472 8470
rect 6489 8406 6553 8470
rect 6570 8406 6634 8470
rect 6651 8406 6715 8470
rect 6732 8406 6796 8470
rect 6813 8406 6877 8470
rect 6894 8406 6958 8470
rect 6975 8406 7039 8470
rect 7056 8406 7120 8470
rect 7137 8406 7201 8470
rect 7218 8406 7282 8470
rect 7299 8406 7363 8470
rect 7380 8406 7444 8470
rect 7461 8406 7525 8470
rect 7542 8406 7606 8470
rect 7623 8406 7687 8470
rect 4695 8320 4759 8384
rect 4777 8320 4841 8384
rect 4859 8320 4923 8384
rect 4941 8320 5005 8384
rect 5023 8320 5087 8384
rect 5105 8320 5169 8384
rect 5187 8320 5251 8384
rect 5269 8320 5333 8384
rect 5351 8320 5415 8384
rect 5433 8320 5497 8384
rect 5515 8320 5579 8384
rect 5597 8320 5661 8384
rect 5679 8320 5743 8384
rect 5760 8320 5824 8384
rect 5841 8320 5905 8384
rect 5922 8320 5986 8384
rect 6003 8320 6067 8384
rect 6084 8320 6148 8384
rect 6165 8320 6229 8384
rect 6246 8320 6310 8384
rect 6327 8320 6391 8384
rect 6408 8320 6472 8384
rect 6489 8320 6553 8384
rect 6570 8320 6634 8384
rect 6651 8320 6715 8384
rect 6732 8320 6796 8384
rect 6813 8320 6877 8384
rect 6894 8320 6958 8384
rect 6975 8320 7039 8384
rect 7056 8320 7120 8384
rect 7137 8320 7201 8384
rect 7218 8320 7282 8384
rect 7299 8320 7363 8384
rect 7380 8320 7444 8384
rect 7461 8320 7525 8384
rect 7542 8320 7606 8384
rect 7623 8320 7687 8384
rect 7813 9177 7877 9241
rect 7897 9177 7961 9241
rect 7981 9177 8045 9241
rect 8065 9177 8129 9241
rect 8149 9177 8213 9241
rect 7813 9092 7877 9156
rect 7897 9092 7961 9156
rect 7981 9092 8045 9156
rect 8065 9092 8129 9156
rect 8149 9092 8213 9156
rect 7813 9007 7877 9071
rect 7897 9007 7961 9071
rect 7981 9007 8045 9071
rect 8065 9007 8129 9071
rect 8149 9007 8213 9071
rect 7813 8922 7877 8986
rect 7897 8922 7961 8986
rect 7981 8922 8045 8986
rect 8065 8922 8129 8986
rect 8149 8922 8213 8986
rect 7813 8837 7877 8901
rect 7897 8837 7961 8901
rect 7981 8837 8045 8901
rect 8065 8837 8129 8901
rect 8149 8837 8213 8901
rect 7813 8752 7877 8816
rect 7897 8752 7961 8816
rect 7981 8752 8045 8816
rect 8065 8752 8129 8816
rect 8149 8752 8213 8816
rect 7813 8667 7877 8731
rect 7897 8667 7961 8731
rect 7981 8667 8045 8731
rect 8065 8667 8129 8731
rect 8149 8667 8213 8731
rect 7813 8581 7877 8645
rect 7897 8581 7961 8645
rect 7981 8581 8045 8645
rect 8065 8581 8129 8645
rect 8149 8581 8213 8645
rect 7813 8495 7877 8559
rect 7897 8495 7961 8559
rect 7981 8495 8045 8559
rect 8065 8495 8129 8559
rect 8149 8495 8213 8559
rect 7813 8409 7877 8473
rect 7897 8409 7961 8473
rect 7981 8409 8045 8473
rect 8065 8409 8129 8473
rect 8149 8409 8213 8473
rect 7813 8323 7877 8387
rect 7897 8323 7961 8387
rect 7981 8323 8045 8387
rect 8065 8323 8129 8387
rect 8149 8323 8213 8387
rect 8333 13637 8397 13701
rect 8417 13637 8481 13701
rect 8501 13637 8565 13701
rect 8585 13637 8649 13701
rect 8669 13637 8733 13701
rect 8333 13556 8397 13620
rect 8417 13556 8481 13620
rect 8501 13556 8565 13620
rect 8585 13556 8649 13620
rect 8669 13556 8733 13620
rect 8333 13475 8397 13539
rect 8417 13475 8481 13539
rect 8501 13475 8565 13539
rect 8585 13475 8649 13539
rect 8669 13475 8733 13539
rect 8333 13394 8397 13458
rect 8417 13394 8481 13458
rect 8501 13394 8565 13458
rect 8585 13394 8649 13458
rect 8669 13394 8733 13458
rect 8333 13313 8397 13377
rect 8417 13313 8481 13377
rect 8501 13313 8565 13377
rect 8585 13313 8649 13377
rect 8669 13313 8733 13377
rect 8333 13232 8397 13296
rect 8417 13232 8481 13296
rect 8501 13232 8565 13296
rect 8585 13232 8649 13296
rect 8669 13232 8733 13296
rect 8333 13151 8397 13215
rect 8417 13151 8481 13215
rect 8501 13151 8565 13215
rect 8585 13151 8649 13215
rect 8669 13151 8733 13215
rect 8333 13069 8397 13133
rect 8417 13069 8481 13133
rect 8501 13069 8565 13133
rect 8585 13069 8649 13133
rect 8669 13069 8733 13133
rect 8333 12987 8397 13051
rect 8417 12987 8481 13051
rect 8501 12987 8565 13051
rect 8585 12987 8649 13051
rect 8669 12987 8733 13051
rect 8333 12905 8397 12969
rect 8417 12905 8481 12969
rect 8501 12905 8565 12969
rect 8585 12905 8649 12969
rect 8669 12905 8733 12969
rect 8333 12823 8397 12887
rect 8417 12823 8481 12887
rect 8501 12823 8565 12887
rect 8585 12823 8649 12887
rect 8669 12823 8733 12887
rect 8859 9180 8923 9244
rect 8940 9180 9004 9244
rect 9021 9180 9085 9244
rect 9102 9180 9166 9244
rect 9183 9180 9247 9244
rect 9264 9180 9328 9244
rect 9345 9180 9409 9244
rect 9426 9180 9490 9244
rect 9507 9180 9571 9244
rect 9588 9180 9652 9244
rect 9669 9180 9733 9244
rect 9750 9180 9814 9244
rect 9831 9180 9895 9244
rect 9912 9180 9976 9244
rect 9993 9180 10057 9244
rect 10073 9180 10137 9244
rect 10153 9180 10217 9244
rect 10233 9180 10297 9244
rect 10313 9180 10377 9244
rect 10393 9180 10457 9244
rect 10473 9180 10537 9244
rect 10553 9180 10617 9244
rect 10633 9180 10697 9244
rect 10713 9180 10777 9244
rect 10793 9180 10857 9244
rect 10873 9180 10937 9244
rect 10953 9180 11017 9244
rect 11033 9180 11097 9244
rect 11113 9180 11177 9244
rect 11193 9180 11257 9244
rect 11273 9180 11337 9244
rect 11353 9180 11417 9244
rect 11433 9180 11497 9244
rect 11513 9180 11577 9244
rect 11593 9180 11657 9244
rect 11673 9180 11737 9244
rect 11753 9180 11817 9244
rect 11833 9180 11897 9244
rect 11913 9180 11977 9244
rect 8859 9094 8923 9158
rect 8940 9094 9004 9158
rect 9021 9094 9085 9158
rect 9102 9094 9166 9158
rect 9183 9094 9247 9158
rect 9264 9094 9328 9158
rect 9345 9094 9409 9158
rect 9426 9094 9490 9158
rect 9507 9094 9571 9158
rect 9588 9094 9652 9158
rect 9669 9094 9733 9158
rect 9750 9094 9814 9158
rect 9831 9094 9895 9158
rect 9912 9094 9976 9158
rect 9993 9094 10057 9158
rect 10073 9094 10137 9158
rect 10153 9094 10217 9158
rect 10233 9094 10297 9158
rect 10313 9094 10377 9158
rect 10393 9094 10457 9158
rect 10473 9094 10537 9158
rect 10553 9094 10617 9158
rect 10633 9094 10697 9158
rect 10713 9094 10777 9158
rect 10793 9094 10857 9158
rect 10873 9094 10937 9158
rect 10953 9094 11017 9158
rect 11033 9094 11097 9158
rect 11113 9094 11177 9158
rect 11193 9094 11257 9158
rect 11273 9094 11337 9158
rect 11353 9094 11417 9158
rect 11433 9094 11497 9158
rect 11513 9094 11577 9158
rect 11593 9094 11657 9158
rect 11673 9094 11737 9158
rect 11753 9094 11817 9158
rect 11833 9094 11897 9158
rect 11913 9094 11977 9158
rect 8859 9008 8923 9072
rect 8940 9008 9004 9072
rect 9021 9008 9085 9072
rect 9102 9008 9166 9072
rect 9183 9008 9247 9072
rect 9264 9008 9328 9072
rect 9345 9008 9409 9072
rect 9426 9008 9490 9072
rect 9507 9008 9571 9072
rect 9588 9008 9652 9072
rect 9669 9008 9733 9072
rect 9750 9008 9814 9072
rect 9831 9008 9895 9072
rect 9912 9008 9976 9072
rect 9993 9008 10057 9072
rect 10073 9008 10137 9072
rect 10153 9008 10217 9072
rect 10233 9008 10297 9072
rect 10313 9008 10377 9072
rect 10393 9008 10457 9072
rect 10473 9008 10537 9072
rect 10553 9008 10617 9072
rect 10633 9008 10697 9072
rect 10713 9008 10777 9072
rect 10793 9008 10857 9072
rect 10873 9008 10937 9072
rect 10953 9008 11017 9072
rect 11033 9008 11097 9072
rect 11113 9008 11177 9072
rect 11193 9008 11257 9072
rect 11273 9008 11337 9072
rect 11353 9008 11417 9072
rect 11433 9008 11497 9072
rect 11513 9008 11577 9072
rect 11593 9008 11657 9072
rect 11673 9008 11737 9072
rect 11753 9008 11817 9072
rect 11833 9008 11897 9072
rect 11913 9008 11977 9072
rect 8859 8922 8923 8986
rect 8940 8922 9004 8986
rect 9021 8922 9085 8986
rect 9102 8922 9166 8986
rect 9183 8922 9247 8986
rect 9264 8922 9328 8986
rect 9345 8922 9409 8986
rect 9426 8922 9490 8986
rect 9507 8922 9571 8986
rect 9588 8922 9652 8986
rect 9669 8922 9733 8986
rect 9750 8922 9814 8986
rect 9831 8922 9895 8986
rect 9912 8922 9976 8986
rect 9993 8922 10057 8986
rect 10073 8922 10137 8986
rect 10153 8922 10217 8986
rect 10233 8922 10297 8986
rect 10313 8922 10377 8986
rect 10393 8922 10457 8986
rect 10473 8922 10537 8986
rect 10553 8922 10617 8986
rect 10633 8922 10697 8986
rect 10713 8922 10777 8986
rect 10793 8922 10857 8986
rect 10873 8922 10937 8986
rect 10953 8922 11017 8986
rect 11033 8922 11097 8986
rect 11113 8922 11177 8986
rect 11193 8922 11257 8986
rect 11273 8922 11337 8986
rect 11353 8922 11417 8986
rect 11433 8922 11497 8986
rect 11513 8922 11577 8986
rect 11593 8922 11657 8986
rect 11673 8922 11737 8986
rect 11753 8922 11817 8986
rect 11833 8922 11897 8986
rect 11913 8922 11977 8986
rect 8859 8836 8923 8900
rect 8940 8836 9004 8900
rect 9021 8836 9085 8900
rect 9102 8836 9166 8900
rect 9183 8836 9247 8900
rect 9264 8836 9328 8900
rect 9345 8836 9409 8900
rect 9426 8836 9490 8900
rect 9507 8836 9571 8900
rect 9588 8836 9652 8900
rect 9669 8836 9733 8900
rect 9750 8836 9814 8900
rect 9831 8836 9895 8900
rect 9912 8836 9976 8900
rect 9993 8836 10057 8900
rect 10073 8836 10137 8900
rect 10153 8836 10217 8900
rect 10233 8836 10297 8900
rect 10313 8836 10377 8900
rect 10393 8836 10457 8900
rect 10473 8836 10537 8900
rect 10553 8836 10617 8900
rect 10633 8836 10697 8900
rect 10713 8836 10777 8900
rect 10793 8836 10857 8900
rect 10873 8836 10937 8900
rect 10953 8836 11017 8900
rect 11033 8836 11097 8900
rect 11113 8836 11177 8900
rect 11193 8836 11257 8900
rect 11273 8836 11337 8900
rect 11353 8836 11417 8900
rect 11433 8836 11497 8900
rect 11513 8836 11577 8900
rect 11593 8836 11657 8900
rect 11673 8836 11737 8900
rect 11753 8836 11817 8900
rect 11833 8836 11897 8900
rect 11913 8836 11977 8900
rect 8859 8750 8923 8814
rect 8940 8750 9004 8814
rect 9021 8750 9085 8814
rect 9102 8750 9166 8814
rect 9183 8750 9247 8814
rect 9264 8750 9328 8814
rect 9345 8750 9409 8814
rect 9426 8750 9490 8814
rect 9507 8750 9571 8814
rect 9588 8750 9652 8814
rect 9669 8750 9733 8814
rect 9750 8750 9814 8814
rect 9831 8750 9895 8814
rect 9912 8750 9976 8814
rect 9993 8750 10057 8814
rect 10073 8750 10137 8814
rect 10153 8750 10217 8814
rect 10233 8750 10297 8814
rect 10313 8750 10377 8814
rect 10393 8750 10457 8814
rect 10473 8750 10537 8814
rect 10553 8750 10617 8814
rect 10633 8750 10697 8814
rect 10713 8750 10777 8814
rect 10793 8750 10857 8814
rect 10873 8750 10937 8814
rect 10953 8750 11017 8814
rect 11033 8750 11097 8814
rect 11113 8750 11177 8814
rect 11193 8750 11257 8814
rect 11273 8750 11337 8814
rect 11353 8750 11417 8814
rect 11433 8750 11497 8814
rect 11513 8750 11577 8814
rect 11593 8750 11657 8814
rect 11673 8750 11737 8814
rect 11753 8750 11817 8814
rect 11833 8750 11897 8814
rect 11913 8750 11977 8814
rect 8859 8664 8923 8728
rect 8940 8664 9004 8728
rect 9021 8664 9085 8728
rect 9102 8664 9166 8728
rect 9183 8664 9247 8728
rect 9264 8664 9328 8728
rect 9345 8664 9409 8728
rect 9426 8664 9490 8728
rect 9507 8664 9571 8728
rect 9588 8664 9652 8728
rect 9669 8664 9733 8728
rect 9750 8664 9814 8728
rect 9831 8664 9895 8728
rect 9912 8664 9976 8728
rect 9993 8664 10057 8728
rect 10073 8664 10137 8728
rect 10153 8664 10217 8728
rect 10233 8664 10297 8728
rect 10313 8664 10377 8728
rect 10393 8664 10457 8728
rect 10473 8664 10537 8728
rect 10553 8664 10617 8728
rect 10633 8664 10697 8728
rect 10713 8664 10777 8728
rect 10793 8664 10857 8728
rect 10873 8664 10937 8728
rect 10953 8664 11017 8728
rect 11033 8664 11097 8728
rect 11113 8664 11177 8728
rect 11193 8664 11257 8728
rect 11273 8664 11337 8728
rect 11353 8664 11417 8728
rect 11433 8664 11497 8728
rect 11513 8664 11577 8728
rect 11593 8664 11657 8728
rect 11673 8664 11737 8728
rect 11753 8664 11817 8728
rect 11833 8664 11897 8728
rect 11913 8664 11977 8728
rect 8859 8578 8923 8642
rect 8940 8578 9004 8642
rect 9021 8578 9085 8642
rect 9102 8578 9166 8642
rect 9183 8578 9247 8642
rect 9264 8578 9328 8642
rect 9345 8578 9409 8642
rect 9426 8578 9490 8642
rect 9507 8578 9571 8642
rect 9588 8578 9652 8642
rect 9669 8578 9733 8642
rect 9750 8578 9814 8642
rect 9831 8578 9895 8642
rect 9912 8578 9976 8642
rect 9993 8578 10057 8642
rect 10073 8578 10137 8642
rect 10153 8578 10217 8642
rect 10233 8578 10297 8642
rect 10313 8578 10377 8642
rect 10393 8578 10457 8642
rect 10473 8578 10537 8642
rect 10553 8578 10617 8642
rect 10633 8578 10697 8642
rect 10713 8578 10777 8642
rect 10793 8578 10857 8642
rect 10873 8578 10937 8642
rect 10953 8578 11017 8642
rect 11033 8578 11097 8642
rect 11113 8578 11177 8642
rect 11193 8578 11257 8642
rect 11273 8578 11337 8642
rect 11353 8578 11417 8642
rect 11433 8578 11497 8642
rect 11513 8578 11577 8642
rect 11593 8578 11657 8642
rect 11673 8578 11737 8642
rect 11753 8578 11817 8642
rect 11833 8578 11897 8642
rect 11913 8578 11977 8642
rect 8859 8492 8923 8556
rect 8940 8492 9004 8556
rect 9021 8492 9085 8556
rect 9102 8492 9166 8556
rect 9183 8492 9247 8556
rect 9264 8492 9328 8556
rect 9345 8492 9409 8556
rect 9426 8492 9490 8556
rect 9507 8492 9571 8556
rect 9588 8492 9652 8556
rect 9669 8492 9733 8556
rect 9750 8492 9814 8556
rect 9831 8492 9895 8556
rect 9912 8492 9976 8556
rect 9993 8492 10057 8556
rect 10073 8492 10137 8556
rect 10153 8492 10217 8556
rect 10233 8492 10297 8556
rect 10313 8492 10377 8556
rect 10393 8492 10457 8556
rect 10473 8492 10537 8556
rect 10553 8492 10617 8556
rect 10633 8492 10697 8556
rect 10713 8492 10777 8556
rect 10793 8492 10857 8556
rect 10873 8492 10937 8556
rect 10953 8492 11017 8556
rect 11033 8492 11097 8556
rect 11113 8492 11177 8556
rect 11193 8492 11257 8556
rect 11273 8492 11337 8556
rect 11353 8492 11417 8556
rect 11433 8492 11497 8556
rect 11513 8492 11577 8556
rect 11593 8492 11657 8556
rect 11673 8492 11737 8556
rect 11753 8492 11817 8556
rect 11833 8492 11897 8556
rect 11913 8492 11977 8556
rect 8859 8406 8923 8470
rect 8940 8406 9004 8470
rect 9021 8406 9085 8470
rect 9102 8406 9166 8470
rect 9183 8406 9247 8470
rect 9264 8406 9328 8470
rect 9345 8406 9409 8470
rect 9426 8406 9490 8470
rect 9507 8406 9571 8470
rect 9588 8406 9652 8470
rect 9669 8406 9733 8470
rect 9750 8406 9814 8470
rect 9831 8406 9895 8470
rect 9912 8406 9976 8470
rect 9993 8406 10057 8470
rect 10073 8406 10137 8470
rect 10153 8406 10217 8470
rect 10233 8406 10297 8470
rect 10313 8406 10377 8470
rect 10393 8406 10457 8470
rect 10473 8406 10537 8470
rect 10553 8406 10617 8470
rect 10633 8406 10697 8470
rect 10713 8406 10777 8470
rect 10793 8406 10857 8470
rect 10873 8406 10937 8470
rect 10953 8406 11017 8470
rect 11033 8406 11097 8470
rect 11113 8406 11177 8470
rect 11193 8406 11257 8470
rect 11273 8406 11337 8470
rect 11353 8406 11417 8470
rect 11433 8406 11497 8470
rect 11513 8406 11577 8470
rect 11593 8406 11657 8470
rect 11673 8406 11737 8470
rect 11753 8406 11817 8470
rect 11833 8406 11897 8470
rect 11913 8406 11977 8470
rect 8859 8320 8923 8384
rect 8940 8320 9004 8384
rect 9021 8320 9085 8384
rect 9102 8320 9166 8384
rect 9183 8320 9247 8384
rect 9264 8320 9328 8384
rect 9345 8320 9409 8384
rect 9426 8320 9490 8384
rect 9507 8320 9571 8384
rect 9588 8320 9652 8384
rect 9669 8320 9733 8384
rect 9750 8320 9814 8384
rect 9831 8320 9895 8384
rect 9912 8320 9976 8384
rect 9993 8320 10057 8384
rect 10073 8320 10137 8384
rect 10153 8320 10217 8384
rect 10233 8320 10297 8384
rect 10313 8320 10377 8384
rect 10393 8320 10457 8384
rect 10473 8320 10537 8384
rect 10553 8320 10617 8384
rect 10633 8320 10697 8384
rect 10713 8320 10777 8384
rect 10793 8320 10857 8384
rect 10873 8320 10937 8384
rect 10953 8320 11017 8384
rect 11033 8320 11097 8384
rect 11113 8320 11177 8384
rect 11193 8320 11257 8384
rect 11273 8320 11337 8384
rect 11353 8320 11417 8384
rect 11433 8320 11497 8384
rect 11513 8320 11577 8384
rect 11593 8320 11657 8384
rect 11673 8320 11737 8384
rect 11753 8320 11817 8384
rect 11833 8320 11897 8384
rect 11913 8320 11977 8384
rect 12165 9180 12229 9244
rect 12246 9180 12310 9244
rect 12327 9180 12391 9244
rect 12408 9180 12472 9244
rect 12489 9180 12553 9244
rect 12570 9180 12634 9244
rect 12651 9180 12715 9244
rect 12732 9180 12796 9244
rect 12813 9180 12877 9244
rect 12894 9180 12958 9244
rect 12975 9180 13039 9244
rect 13056 9180 13120 9244
rect 13137 9180 13201 9244
rect 13218 9180 13282 9244
rect 13299 9180 13363 9244
rect 13380 9180 13444 9244
rect 13461 9180 13525 9244
rect 13542 9180 13606 9244
rect 13623 9180 13687 9244
rect 13704 9180 13768 9244
rect 13785 9180 13849 9244
rect 13866 9180 13930 9244
rect 13947 9180 14011 9244
rect 14028 9180 14092 9244
rect 14109 9180 14173 9244
rect 14190 9180 14254 9244
rect 14271 9180 14335 9244
rect 14352 9180 14416 9244
rect 14433 9180 14497 9244
rect 14513 9180 14577 9244
rect 14593 9180 14657 9244
rect 14673 9180 14737 9244
rect 14753 9180 14817 9244
rect 14833 9180 14897 9244
rect 14913 9180 14977 9244
rect 14993 9180 15057 9244
rect 15073 9180 15137 9244
rect 15153 9180 15217 9244
rect 15233 9180 15297 9244
rect 15313 9180 15377 9244
rect 15393 9180 15457 9244
rect 15473 9180 15537 9244
rect 15553 9180 15617 9244
rect 12165 9094 12229 9158
rect 12246 9094 12310 9158
rect 12327 9094 12391 9158
rect 12408 9094 12472 9158
rect 12489 9094 12553 9158
rect 12570 9094 12634 9158
rect 12651 9094 12715 9158
rect 12732 9094 12796 9158
rect 12813 9094 12877 9158
rect 12894 9094 12958 9158
rect 12975 9094 13039 9158
rect 13056 9094 13120 9158
rect 13137 9094 13201 9158
rect 13218 9094 13282 9158
rect 13299 9094 13363 9158
rect 13380 9094 13444 9158
rect 13461 9094 13525 9158
rect 13542 9094 13606 9158
rect 13623 9094 13687 9158
rect 13704 9094 13768 9158
rect 13785 9094 13849 9158
rect 13866 9094 13930 9158
rect 13947 9094 14011 9158
rect 14028 9094 14092 9158
rect 14109 9094 14173 9158
rect 14190 9094 14254 9158
rect 14271 9094 14335 9158
rect 14352 9094 14416 9158
rect 14433 9094 14497 9158
rect 14513 9094 14577 9158
rect 14593 9094 14657 9158
rect 14673 9094 14737 9158
rect 14753 9094 14817 9158
rect 14833 9094 14897 9158
rect 14913 9094 14977 9158
rect 14993 9094 15057 9158
rect 15073 9094 15137 9158
rect 15153 9094 15217 9158
rect 15233 9094 15297 9158
rect 15313 9094 15377 9158
rect 15393 9094 15457 9158
rect 15473 9094 15537 9158
rect 15553 9094 15617 9158
rect 12165 9008 12229 9072
rect 12246 9008 12310 9072
rect 12327 9008 12391 9072
rect 12408 9008 12472 9072
rect 12489 9008 12553 9072
rect 12570 9008 12634 9072
rect 12651 9008 12715 9072
rect 12732 9008 12796 9072
rect 12813 9008 12877 9072
rect 12894 9008 12958 9072
rect 12975 9008 13039 9072
rect 13056 9008 13120 9072
rect 13137 9008 13201 9072
rect 13218 9008 13282 9072
rect 13299 9008 13363 9072
rect 13380 9008 13444 9072
rect 13461 9008 13525 9072
rect 13542 9008 13606 9072
rect 13623 9008 13687 9072
rect 13704 9008 13768 9072
rect 13785 9008 13849 9072
rect 13866 9008 13930 9072
rect 13947 9008 14011 9072
rect 14028 9008 14092 9072
rect 14109 9008 14173 9072
rect 14190 9008 14254 9072
rect 14271 9008 14335 9072
rect 14352 9008 14416 9072
rect 14433 9008 14497 9072
rect 14513 9008 14577 9072
rect 14593 9008 14657 9072
rect 14673 9008 14737 9072
rect 14753 9008 14817 9072
rect 14833 9008 14897 9072
rect 14913 9008 14977 9072
rect 14993 9008 15057 9072
rect 15073 9008 15137 9072
rect 15153 9008 15217 9072
rect 15233 9008 15297 9072
rect 15313 9008 15377 9072
rect 15393 9008 15457 9072
rect 15473 9008 15537 9072
rect 15553 9008 15617 9072
rect 12165 8922 12229 8986
rect 12246 8922 12310 8986
rect 12327 8922 12391 8986
rect 12408 8922 12472 8986
rect 12489 8922 12553 8986
rect 12570 8922 12634 8986
rect 12651 8922 12715 8986
rect 12732 8922 12796 8986
rect 12813 8922 12877 8986
rect 12894 8922 12958 8986
rect 12975 8922 13039 8986
rect 13056 8922 13120 8986
rect 13137 8922 13201 8986
rect 13218 8922 13282 8986
rect 13299 8922 13363 8986
rect 13380 8922 13444 8986
rect 13461 8922 13525 8986
rect 13542 8922 13606 8986
rect 13623 8922 13687 8986
rect 13704 8922 13768 8986
rect 13785 8922 13849 8986
rect 13866 8922 13930 8986
rect 13947 8922 14011 8986
rect 14028 8922 14092 8986
rect 14109 8922 14173 8986
rect 14190 8922 14254 8986
rect 14271 8922 14335 8986
rect 14352 8922 14416 8986
rect 14433 8922 14497 8986
rect 14513 8922 14577 8986
rect 14593 8922 14657 8986
rect 14673 8922 14737 8986
rect 14753 8922 14817 8986
rect 14833 8922 14897 8986
rect 14913 8922 14977 8986
rect 14993 8922 15057 8986
rect 15073 8922 15137 8986
rect 15153 8922 15217 8986
rect 15233 8922 15297 8986
rect 15313 8922 15377 8986
rect 15393 8922 15457 8986
rect 15473 8922 15537 8986
rect 15553 8922 15617 8986
rect 12165 8836 12229 8900
rect 12246 8836 12310 8900
rect 12327 8836 12391 8900
rect 12408 8836 12472 8900
rect 12489 8836 12553 8900
rect 12570 8836 12634 8900
rect 12651 8836 12715 8900
rect 12732 8836 12796 8900
rect 12813 8836 12877 8900
rect 12894 8836 12958 8900
rect 12975 8836 13039 8900
rect 13056 8836 13120 8900
rect 13137 8836 13201 8900
rect 13218 8836 13282 8900
rect 13299 8836 13363 8900
rect 13380 8836 13444 8900
rect 13461 8836 13525 8900
rect 13542 8836 13606 8900
rect 13623 8836 13687 8900
rect 13704 8836 13768 8900
rect 13785 8836 13849 8900
rect 13866 8836 13930 8900
rect 13947 8836 14011 8900
rect 14028 8836 14092 8900
rect 14109 8836 14173 8900
rect 14190 8836 14254 8900
rect 14271 8836 14335 8900
rect 14352 8836 14416 8900
rect 14433 8836 14497 8900
rect 14513 8836 14577 8900
rect 14593 8836 14657 8900
rect 14673 8836 14737 8900
rect 14753 8836 14817 8900
rect 14833 8836 14897 8900
rect 14913 8836 14977 8900
rect 14993 8836 15057 8900
rect 15073 8836 15137 8900
rect 15153 8836 15217 8900
rect 15233 8836 15297 8900
rect 15313 8836 15377 8900
rect 15393 8836 15457 8900
rect 15473 8836 15537 8900
rect 15553 8836 15617 8900
rect 12165 8750 12229 8814
rect 12246 8750 12310 8814
rect 12327 8750 12391 8814
rect 12408 8750 12472 8814
rect 12489 8750 12553 8814
rect 12570 8750 12634 8814
rect 12651 8750 12715 8814
rect 12732 8750 12796 8814
rect 12813 8750 12877 8814
rect 12894 8750 12958 8814
rect 12975 8750 13039 8814
rect 13056 8750 13120 8814
rect 13137 8750 13201 8814
rect 13218 8750 13282 8814
rect 13299 8750 13363 8814
rect 13380 8750 13444 8814
rect 13461 8750 13525 8814
rect 13542 8750 13606 8814
rect 13623 8750 13687 8814
rect 13704 8750 13768 8814
rect 13785 8750 13849 8814
rect 13866 8750 13930 8814
rect 13947 8750 14011 8814
rect 14028 8750 14092 8814
rect 14109 8750 14173 8814
rect 14190 8750 14254 8814
rect 14271 8750 14335 8814
rect 14352 8750 14416 8814
rect 14433 8750 14497 8814
rect 14513 8750 14577 8814
rect 14593 8750 14657 8814
rect 14673 8750 14737 8814
rect 14753 8750 14817 8814
rect 14833 8750 14897 8814
rect 14913 8750 14977 8814
rect 14993 8750 15057 8814
rect 15073 8750 15137 8814
rect 15153 8750 15217 8814
rect 15233 8750 15297 8814
rect 15313 8750 15377 8814
rect 15393 8750 15457 8814
rect 15473 8750 15537 8814
rect 15553 8750 15617 8814
rect 12165 8664 12229 8728
rect 12246 8664 12310 8728
rect 12327 8664 12391 8728
rect 12408 8664 12472 8728
rect 12489 8664 12553 8728
rect 12570 8664 12634 8728
rect 12651 8664 12715 8728
rect 12732 8664 12796 8728
rect 12813 8664 12877 8728
rect 12894 8664 12958 8728
rect 12975 8664 13039 8728
rect 13056 8664 13120 8728
rect 13137 8664 13201 8728
rect 13218 8664 13282 8728
rect 13299 8664 13363 8728
rect 13380 8664 13444 8728
rect 13461 8664 13525 8728
rect 13542 8664 13606 8728
rect 13623 8664 13687 8728
rect 13704 8664 13768 8728
rect 13785 8664 13849 8728
rect 13866 8664 13930 8728
rect 13947 8664 14011 8728
rect 14028 8664 14092 8728
rect 14109 8664 14173 8728
rect 14190 8664 14254 8728
rect 14271 8664 14335 8728
rect 14352 8664 14416 8728
rect 14433 8664 14497 8728
rect 14513 8664 14577 8728
rect 14593 8664 14657 8728
rect 14673 8664 14737 8728
rect 14753 8664 14817 8728
rect 14833 8664 14897 8728
rect 14913 8664 14977 8728
rect 14993 8664 15057 8728
rect 15073 8664 15137 8728
rect 15153 8664 15217 8728
rect 15233 8664 15297 8728
rect 15313 8664 15377 8728
rect 15393 8664 15457 8728
rect 15473 8664 15537 8728
rect 15553 8664 15617 8728
rect 12165 8578 12229 8642
rect 12246 8578 12310 8642
rect 12327 8578 12391 8642
rect 12408 8578 12472 8642
rect 12489 8578 12553 8642
rect 12570 8578 12634 8642
rect 12651 8578 12715 8642
rect 12732 8578 12796 8642
rect 12813 8578 12877 8642
rect 12894 8578 12958 8642
rect 12975 8578 13039 8642
rect 13056 8578 13120 8642
rect 13137 8578 13201 8642
rect 13218 8578 13282 8642
rect 13299 8578 13363 8642
rect 13380 8578 13444 8642
rect 13461 8578 13525 8642
rect 13542 8578 13606 8642
rect 13623 8578 13687 8642
rect 13704 8578 13768 8642
rect 13785 8578 13849 8642
rect 13866 8578 13930 8642
rect 13947 8578 14011 8642
rect 14028 8578 14092 8642
rect 14109 8578 14173 8642
rect 14190 8578 14254 8642
rect 14271 8578 14335 8642
rect 14352 8578 14416 8642
rect 14433 8578 14497 8642
rect 14513 8578 14577 8642
rect 14593 8578 14657 8642
rect 14673 8578 14737 8642
rect 14753 8578 14817 8642
rect 14833 8578 14897 8642
rect 14913 8578 14977 8642
rect 14993 8578 15057 8642
rect 15073 8578 15137 8642
rect 15153 8578 15217 8642
rect 15233 8578 15297 8642
rect 15313 8578 15377 8642
rect 15393 8578 15457 8642
rect 15473 8578 15537 8642
rect 15553 8578 15617 8642
rect 12165 8492 12229 8556
rect 12246 8492 12310 8556
rect 12327 8492 12391 8556
rect 12408 8492 12472 8556
rect 12489 8492 12553 8556
rect 12570 8492 12634 8556
rect 12651 8492 12715 8556
rect 12732 8492 12796 8556
rect 12813 8492 12877 8556
rect 12894 8492 12958 8556
rect 12975 8492 13039 8556
rect 13056 8492 13120 8556
rect 13137 8492 13201 8556
rect 13218 8492 13282 8556
rect 13299 8492 13363 8556
rect 13380 8492 13444 8556
rect 13461 8492 13525 8556
rect 13542 8492 13606 8556
rect 13623 8492 13687 8556
rect 13704 8492 13768 8556
rect 13785 8492 13849 8556
rect 13866 8492 13930 8556
rect 13947 8492 14011 8556
rect 14028 8492 14092 8556
rect 14109 8492 14173 8556
rect 14190 8492 14254 8556
rect 14271 8492 14335 8556
rect 14352 8492 14416 8556
rect 14433 8492 14497 8556
rect 14513 8492 14577 8556
rect 14593 8492 14657 8556
rect 14673 8492 14737 8556
rect 14753 8492 14817 8556
rect 14833 8492 14897 8556
rect 14913 8492 14977 8556
rect 14993 8492 15057 8556
rect 15073 8492 15137 8556
rect 15153 8492 15217 8556
rect 15233 8492 15297 8556
rect 15313 8492 15377 8556
rect 15393 8492 15457 8556
rect 15473 8492 15537 8556
rect 15553 8492 15617 8556
rect 12165 8406 12229 8470
rect 12246 8406 12310 8470
rect 12327 8406 12391 8470
rect 12408 8406 12472 8470
rect 12489 8406 12553 8470
rect 12570 8406 12634 8470
rect 12651 8406 12715 8470
rect 12732 8406 12796 8470
rect 12813 8406 12877 8470
rect 12894 8406 12958 8470
rect 12975 8406 13039 8470
rect 13056 8406 13120 8470
rect 13137 8406 13201 8470
rect 13218 8406 13282 8470
rect 13299 8406 13363 8470
rect 13380 8406 13444 8470
rect 13461 8406 13525 8470
rect 13542 8406 13606 8470
rect 13623 8406 13687 8470
rect 13704 8406 13768 8470
rect 13785 8406 13849 8470
rect 13866 8406 13930 8470
rect 13947 8406 14011 8470
rect 14028 8406 14092 8470
rect 14109 8406 14173 8470
rect 14190 8406 14254 8470
rect 14271 8406 14335 8470
rect 14352 8406 14416 8470
rect 14433 8406 14497 8470
rect 14513 8406 14577 8470
rect 14593 8406 14657 8470
rect 14673 8406 14737 8470
rect 14753 8406 14817 8470
rect 14833 8406 14897 8470
rect 14913 8406 14977 8470
rect 14993 8406 15057 8470
rect 15073 8406 15137 8470
rect 15153 8406 15217 8470
rect 15233 8406 15297 8470
rect 15313 8406 15377 8470
rect 15393 8406 15457 8470
rect 15473 8406 15537 8470
rect 15553 8406 15617 8470
rect 12165 8320 12229 8384
rect 12246 8320 12310 8384
rect 12327 8320 12391 8384
rect 12408 8320 12472 8384
rect 12489 8320 12553 8384
rect 12570 8320 12634 8384
rect 12651 8320 12715 8384
rect 12732 8320 12796 8384
rect 12813 8320 12877 8384
rect 12894 8320 12958 8384
rect 12975 8320 13039 8384
rect 13056 8320 13120 8384
rect 13137 8320 13201 8384
rect 13218 8320 13282 8384
rect 13299 8320 13363 8384
rect 13380 8320 13444 8384
rect 13461 8320 13525 8384
rect 13542 8320 13606 8384
rect 13623 8320 13687 8384
rect 13704 8320 13768 8384
rect 13785 8320 13849 8384
rect 13866 8320 13930 8384
rect 13947 8320 14011 8384
rect 14028 8320 14092 8384
rect 14109 8320 14173 8384
rect 14190 8320 14254 8384
rect 14271 8320 14335 8384
rect 14352 8320 14416 8384
rect 14433 8320 14497 8384
rect 14513 8320 14577 8384
rect 14593 8320 14657 8384
rect 14673 8320 14737 8384
rect 14753 8320 14817 8384
rect 14833 8320 14897 8384
rect 14913 8320 14977 8384
rect 14993 8320 15057 8384
rect 15073 8320 15137 8384
rect 15153 8320 15217 8384
rect 15233 8320 15297 8384
rect 15313 8320 15377 8384
rect 15393 8320 15457 8384
rect 15473 8320 15537 8384
rect 15553 8320 15617 8384
rect 11674 2698 11738 2701
rect 11674 2642 11678 2698
rect 11678 2642 11734 2698
rect 11734 2642 11738 2698
rect 11674 2637 11738 2642
rect 11674 2576 11738 2579
rect 11674 2520 11678 2576
rect 11678 2520 11734 2576
rect 11734 2520 11738 2576
rect 11674 2515 11738 2520
rect 11674 2454 11738 2457
rect 11674 2398 11678 2454
rect 11678 2398 11734 2454
rect 11734 2398 11738 2454
rect 11674 2393 11738 2398
rect 11674 2332 11738 2335
rect 11674 2276 11678 2332
rect 11678 2276 11734 2332
rect 11734 2276 11738 2332
rect 11674 2271 11738 2276
rect 11674 2210 11738 2213
rect 11674 2154 11678 2210
rect 11678 2154 11734 2210
rect 11734 2154 11738 2210
rect 11674 2149 11738 2154
rect 11674 2088 11738 2091
rect 11674 2032 11678 2088
rect 11678 2032 11734 2088
rect 11734 2032 11738 2088
rect 11674 2027 11738 2032
rect 11674 1965 11738 1969
rect 11674 1909 11678 1965
rect 11678 1909 11734 1965
rect 11734 1909 11738 1965
rect 11674 1905 11738 1909
rect 11674 1842 11738 1847
rect 11674 1786 11678 1842
rect 11678 1786 11734 1842
rect 11734 1786 11738 1842
rect 11674 1783 11738 1786
<< metal4 >>
rect 0 39964 16000 40000
rect 0 39728 215 39964
rect 451 39728 537 39964
rect 773 39728 859 39964
rect 1095 39728 1181 39964
rect 1417 39728 1503 39964
rect 1739 39728 1825 39964
rect 2061 39728 2147 39964
rect 2383 39728 2469 39964
rect 2705 39728 2791 39964
rect 3027 39728 3113 39964
rect 3349 39728 3435 39964
rect 3671 39728 3757 39964
rect 3993 39728 4079 39964
rect 4315 39728 4401 39964
rect 4637 39728 4723 39964
rect 4959 39728 5045 39964
rect 5281 39728 5367 39964
rect 5603 39728 5689 39964
rect 5925 39728 6011 39964
rect 6247 39728 6332 39964
rect 6568 39728 6653 39964
rect 6889 39728 6974 39964
rect 7210 39728 7295 39964
rect 7531 39728 7616 39964
rect 7852 39728 7937 39964
rect 8173 39728 8258 39964
rect 8494 39728 8579 39964
rect 8815 39728 8900 39964
rect 9136 39728 9221 39964
rect 9457 39728 9542 39964
rect 9778 39728 9863 39964
rect 10099 39728 10184 39964
rect 10420 39728 10505 39964
rect 10741 39728 10826 39964
rect 11062 39728 11147 39964
rect 11383 39728 11468 39964
rect 11704 39728 11789 39964
rect 12025 39728 12110 39964
rect 12346 39728 12431 39964
rect 12667 39728 12752 39964
rect 12988 39728 13073 39964
rect 13309 39728 13394 39964
rect 13630 39728 13715 39964
rect 13951 39728 14036 39964
rect 14272 39728 14357 39964
rect 14593 39728 14678 39964
rect 14914 39728 14999 39964
rect 15235 39728 15320 39964
rect 15556 39728 16000 39964
rect 0 39640 16000 39728
rect 0 39404 215 39640
rect 451 39404 537 39640
rect 773 39404 859 39640
rect 1095 39404 1181 39640
rect 1417 39404 1503 39640
rect 1739 39404 1825 39640
rect 2061 39404 2147 39640
rect 2383 39404 2469 39640
rect 2705 39404 2791 39640
rect 3027 39404 3113 39640
rect 3349 39404 3435 39640
rect 3671 39404 3757 39640
rect 3993 39404 4079 39640
rect 4315 39404 4401 39640
rect 4637 39404 4723 39640
rect 4959 39404 5045 39640
rect 5281 39404 5367 39640
rect 5603 39404 5689 39640
rect 5925 39404 6011 39640
rect 6247 39404 6332 39640
rect 6568 39404 6653 39640
rect 6889 39404 6974 39640
rect 7210 39404 7295 39640
rect 7531 39404 7616 39640
rect 7852 39404 7937 39640
rect 8173 39404 8258 39640
rect 8494 39404 8579 39640
rect 8815 39404 8900 39640
rect 9136 39404 9221 39640
rect 9457 39404 9542 39640
rect 9778 39404 9863 39640
rect 10099 39404 10184 39640
rect 10420 39404 10505 39640
rect 10741 39404 10826 39640
rect 11062 39404 11147 39640
rect 11383 39404 11468 39640
rect 11704 39404 11789 39640
rect 12025 39404 12110 39640
rect 12346 39404 12431 39640
rect 12667 39404 12752 39640
rect 12988 39404 13073 39640
rect 13309 39404 13394 39640
rect 13630 39404 13715 39640
rect 13951 39404 14036 39640
rect 14272 39404 14357 39640
rect 14593 39404 14678 39640
rect 14914 39404 14999 39640
rect 15235 39404 15320 39640
rect 15556 39404 16000 39640
rect 0 39316 16000 39404
rect 0 39080 215 39316
rect 451 39080 537 39316
rect 773 39080 859 39316
rect 1095 39080 1181 39316
rect 1417 39080 1503 39316
rect 1739 39080 1825 39316
rect 2061 39080 2147 39316
rect 2383 39080 2469 39316
rect 2705 39080 2791 39316
rect 3027 39080 3113 39316
rect 3349 39080 3435 39316
rect 3671 39080 3757 39316
rect 3993 39080 4079 39316
rect 4315 39080 4401 39316
rect 4637 39080 4723 39316
rect 4959 39080 5045 39316
rect 5281 39080 5367 39316
rect 5603 39080 5689 39316
rect 5925 39080 6011 39316
rect 6247 39080 6332 39316
rect 6568 39080 6653 39316
rect 6889 39080 6974 39316
rect 7210 39080 7295 39316
rect 7531 39080 7616 39316
rect 7852 39080 7937 39316
rect 8173 39080 8258 39316
rect 8494 39080 8579 39316
rect 8815 39080 8900 39316
rect 9136 39080 9221 39316
rect 9457 39080 9542 39316
rect 9778 39080 9863 39316
rect 10099 39080 10184 39316
rect 10420 39080 10505 39316
rect 10741 39080 10826 39316
rect 11062 39080 11147 39316
rect 11383 39080 11468 39316
rect 11704 39080 11789 39316
rect 12025 39080 12110 39316
rect 12346 39080 12431 39316
rect 12667 39080 12752 39316
rect 12988 39080 13073 39316
rect 13309 39080 13394 39316
rect 13630 39080 13715 39316
rect 13951 39080 14036 39316
rect 14272 39080 14357 39316
rect 14593 39080 14678 39316
rect 14914 39080 14999 39316
rect 15235 39080 15320 39316
rect 15556 39080 16000 39316
rect 0 38992 16000 39080
rect 0 38756 215 38992
rect 451 38756 537 38992
rect 773 38756 859 38992
rect 1095 38756 1181 38992
rect 1417 38756 1503 38992
rect 1739 38756 1825 38992
rect 2061 38756 2147 38992
rect 2383 38756 2469 38992
rect 2705 38756 2791 38992
rect 3027 38756 3113 38992
rect 3349 38756 3435 38992
rect 3671 38756 3757 38992
rect 3993 38756 4079 38992
rect 4315 38756 4401 38992
rect 4637 38756 4723 38992
rect 4959 38756 5045 38992
rect 5281 38756 5367 38992
rect 5603 38756 5689 38992
rect 5925 38756 6011 38992
rect 6247 38756 6332 38992
rect 6568 38756 6653 38992
rect 6889 38756 6974 38992
rect 7210 38756 7295 38992
rect 7531 38756 7616 38992
rect 7852 38756 7937 38992
rect 8173 38756 8258 38992
rect 8494 38756 8579 38992
rect 8815 38756 8900 38992
rect 9136 38756 9221 38992
rect 9457 38756 9542 38992
rect 9778 38756 9863 38992
rect 10099 38756 10184 38992
rect 10420 38756 10505 38992
rect 10741 38756 10826 38992
rect 11062 38756 11147 38992
rect 11383 38756 11468 38992
rect 11704 38756 11789 38992
rect 12025 38756 12110 38992
rect 12346 38756 12431 38992
rect 12667 38756 12752 38992
rect 12988 38756 13073 38992
rect 13309 38756 13394 38992
rect 13630 38756 13715 38992
rect 13951 38756 14036 38992
rect 14272 38756 14357 38992
rect 14593 38756 14678 38992
rect 14914 38756 14999 38992
rect 15235 38756 15320 38992
rect 15556 38756 16000 38992
rect 0 38668 16000 38756
rect 0 38432 215 38668
rect 451 38432 537 38668
rect 773 38432 859 38668
rect 1095 38432 1181 38668
rect 1417 38432 1503 38668
rect 1739 38432 1825 38668
rect 2061 38432 2147 38668
rect 2383 38432 2469 38668
rect 2705 38432 2791 38668
rect 3027 38432 3113 38668
rect 3349 38432 3435 38668
rect 3671 38432 3757 38668
rect 3993 38432 4079 38668
rect 4315 38432 4401 38668
rect 4637 38432 4723 38668
rect 4959 38432 5045 38668
rect 5281 38432 5367 38668
rect 5603 38432 5689 38668
rect 5925 38432 6011 38668
rect 6247 38432 6332 38668
rect 6568 38432 6653 38668
rect 6889 38432 6974 38668
rect 7210 38432 7295 38668
rect 7531 38432 7616 38668
rect 7852 38432 7937 38668
rect 8173 38432 8258 38668
rect 8494 38432 8579 38668
rect 8815 38432 8900 38668
rect 9136 38432 9221 38668
rect 9457 38432 9542 38668
rect 9778 38432 9863 38668
rect 10099 38432 10184 38668
rect 10420 38432 10505 38668
rect 10741 38432 10826 38668
rect 11062 38432 11147 38668
rect 11383 38432 11468 38668
rect 11704 38432 11789 38668
rect 12025 38432 12110 38668
rect 12346 38432 12431 38668
rect 12667 38432 12752 38668
rect 12988 38432 13073 38668
rect 13309 38432 13394 38668
rect 13630 38432 13715 38668
rect 13951 38432 14036 38668
rect 14272 38432 14357 38668
rect 14593 38432 14678 38668
rect 14914 38432 14999 38668
rect 15235 38432 15320 38668
rect 15556 38432 16000 38668
rect 0 38344 16000 38432
rect 0 38108 215 38344
rect 451 38108 537 38344
rect 773 38108 859 38344
rect 1095 38108 1181 38344
rect 1417 38108 1503 38344
rect 1739 38108 1825 38344
rect 2061 38108 2147 38344
rect 2383 38108 2469 38344
rect 2705 38108 2791 38344
rect 3027 38108 3113 38344
rect 3349 38108 3435 38344
rect 3671 38108 3757 38344
rect 3993 38108 4079 38344
rect 4315 38108 4401 38344
rect 4637 38108 4723 38344
rect 4959 38108 5045 38344
rect 5281 38108 5367 38344
rect 5603 38108 5689 38344
rect 5925 38108 6011 38344
rect 6247 38108 6332 38344
rect 6568 38108 6653 38344
rect 6889 38108 6974 38344
rect 7210 38108 7295 38344
rect 7531 38108 7616 38344
rect 7852 38108 7937 38344
rect 8173 38108 8258 38344
rect 8494 38108 8579 38344
rect 8815 38108 8900 38344
rect 9136 38108 9221 38344
rect 9457 38108 9542 38344
rect 9778 38108 9863 38344
rect 10099 38108 10184 38344
rect 10420 38108 10505 38344
rect 10741 38108 10826 38344
rect 11062 38108 11147 38344
rect 11383 38108 11468 38344
rect 11704 38108 11789 38344
rect 12025 38108 12110 38344
rect 12346 38108 12431 38344
rect 12667 38108 12752 38344
rect 12988 38108 13073 38344
rect 13309 38108 13394 38344
rect 13630 38108 13715 38344
rect 13951 38108 14036 38344
rect 14272 38108 14357 38344
rect 14593 38108 14678 38344
rect 14914 38108 14999 38344
rect 15235 38108 15320 38344
rect 15556 38108 16000 38344
rect 0 38020 16000 38108
rect 0 37784 215 38020
rect 451 37784 537 38020
rect 773 37784 859 38020
rect 1095 37784 1181 38020
rect 1417 37784 1503 38020
rect 1739 37784 1825 38020
rect 2061 37784 2147 38020
rect 2383 37784 2469 38020
rect 2705 37784 2791 38020
rect 3027 37784 3113 38020
rect 3349 37784 3435 38020
rect 3671 37784 3757 38020
rect 3993 37784 4079 38020
rect 4315 37784 4401 38020
rect 4637 37784 4723 38020
rect 4959 37784 5045 38020
rect 5281 37784 5367 38020
rect 5603 37784 5689 38020
rect 5925 37784 6011 38020
rect 6247 37784 6332 38020
rect 6568 37784 6653 38020
rect 6889 37784 6974 38020
rect 7210 37784 7295 38020
rect 7531 37784 7616 38020
rect 7852 37784 7937 38020
rect 8173 37784 8258 38020
rect 8494 37784 8579 38020
rect 8815 37784 8900 38020
rect 9136 37784 9221 38020
rect 9457 37784 9542 38020
rect 9778 37784 9863 38020
rect 10099 37784 10184 38020
rect 10420 37784 10505 38020
rect 10741 37784 10826 38020
rect 11062 37784 11147 38020
rect 11383 37784 11468 38020
rect 11704 37784 11789 38020
rect 12025 37784 12110 38020
rect 12346 37784 12431 38020
rect 12667 37784 12752 38020
rect 12988 37784 13073 38020
rect 13309 37784 13394 38020
rect 13630 37784 13715 38020
rect 13951 37784 14036 38020
rect 14272 37784 14357 38020
rect 14593 37784 14678 38020
rect 14914 37784 14999 38020
rect 15235 37784 15320 38020
rect 15556 37784 16000 38020
rect 0 37696 16000 37784
rect 0 37460 215 37696
rect 451 37460 537 37696
rect 773 37460 859 37696
rect 1095 37460 1181 37696
rect 1417 37460 1503 37696
rect 1739 37460 1825 37696
rect 2061 37460 2147 37696
rect 2383 37460 2469 37696
rect 2705 37460 2791 37696
rect 3027 37460 3113 37696
rect 3349 37460 3435 37696
rect 3671 37460 3757 37696
rect 3993 37460 4079 37696
rect 4315 37460 4401 37696
rect 4637 37460 4723 37696
rect 4959 37460 5045 37696
rect 5281 37460 5367 37696
rect 5603 37460 5689 37696
rect 5925 37460 6011 37696
rect 6247 37460 6332 37696
rect 6568 37460 6653 37696
rect 6889 37460 6974 37696
rect 7210 37460 7295 37696
rect 7531 37460 7616 37696
rect 7852 37460 7937 37696
rect 8173 37460 8258 37696
rect 8494 37460 8579 37696
rect 8815 37460 8900 37696
rect 9136 37460 9221 37696
rect 9457 37460 9542 37696
rect 9778 37460 9863 37696
rect 10099 37460 10184 37696
rect 10420 37460 10505 37696
rect 10741 37460 10826 37696
rect 11062 37460 11147 37696
rect 11383 37460 11468 37696
rect 11704 37460 11789 37696
rect 12025 37460 12110 37696
rect 12346 37460 12431 37696
rect 12667 37460 12752 37696
rect 12988 37460 13073 37696
rect 13309 37460 13394 37696
rect 13630 37460 13715 37696
rect 13951 37460 14036 37696
rect 14272 37460 14357 37696
rect 14593 37460 14678 37696
rect 14914 37460 14999 37696
rect 15235 37460 15320 37696
rect 15556 37460 16000 37696
rect 0 37372 16000 37460
rect 0 37136 215 37372
rect 451 37136 537 37372
rect 773 37136 859 37372
rect 1095 37136 1181 37372
rect 1417 37136 1503 37372
rect 1739 37136 1825 37372
rect 2061 37136 2147 37372
rect 2383 37136 2469 37372
rect 2705 37136 2791 37372
rect 3027 37136 3113 37372
rect 3349 37136 3435 37372
rect 3671 37136 3757 37372
rect 3993 37136 4079 37372
rect 4315 37136 4401 37372
rect 4637 37136 4723 37372
rect 4959 37136 5045 37372
rect 5281 37136 5367 37372
rect 5603 37136 5689 37372
rect 5925 37136 6011 37372
rect 6247 37136 6332 37372
rect 6568 37136 6653 37372
rect 6889 37136 6974 37372
rect 7210 37136 7295 37372
rect 7531 37136 7616 37372
rect 7852 37136 7937 37372
rect 8173 37136 8258 37372
rect 8494 37136 8579 37372
rect 8815 37136 8900 37372
rect 9136 37136 9221 37372
rect 9457 37136 9542 37372
rect 9778 37136 9863 37372
rect 10099 37136 10184 37372
rect 10420 37136 10505 37372
rect 10741 37136 10826 37372
rect 11062 37136 11147 37372
rect 11383 37136 11468 37372
rect 11704 37136 11789 37372
rect 12025 37136 12110 37372
rect 12346 37136 12431 37372
rect 12667 37136 12752 37372
rect 12988 37136 13073 37372
rect 13309 37136 13394 37372
rect 13630 37136 13715 37372
rect 13951 37136 14036 37372
rect 14272 37136 14357 37372
rect 14593 37136 14678 37372
rect 14914 37136 14999 37372
rect 15235 37136 15320 37372
rect 15556 37136 16000 37372
rect 0 37048 16000 37136
rect 0 36812 215 37048
rect 451 36812 537 37048
rect 773 36812 859 37048
rect 1095 36812 1181 37048
rect 1417 36812 1503 37048
rect 1739 36812 1825 37048
rect 2061 36812 2147 37048
rect 2383 36812 2469 37048
rect 2705 36812 2791 37048
rect 3027 36812 3113 37048
rect 3349 36812 3435 37048
rect 3671 36812 3757 37048
rect 3993 36812 4079 37048
rect 4315 36812 4401 37048
rect 4637 36812 4723 37048
rect 4959 36812 5045 37048
rect 5281 36812 5367 37048
rect 5603 36812 5689 37048
rect 5925 36812 6011 37048
rect 6247 36812 6332 37048
rect 6568 36812 6653 37048
rect 6889 36812 6974 37048
rect 7210 36812 7295 37048
rect 7531 36812 7616 37048
rect 7852 36812 7937 37048
rect 8173 36812 8258 37048
rect 8494 36812 8579 37048
rect 8815 36812 8900 37048
rect 9136 36812 9221 37048
rect 9457 36812 9542 37048
rect 9778 36812 9863 37048
rect 10099 36812 10184 37048
rect 10420 36812 10505 37048
rect 10741 36812 10826 37048
rect 11062 36812 11147 37048
rect 11383 36812 11468 37048
rect 11704 36812 11789 37048
rect 12025 36812 12110 37048
rect 12346 36812 12431 37048
rect 12667 36812 12752 37048
rect 12988 36812 13073 37048
rect 13309 36812 13394 37048
rect 13630 36812 13715 37048
rect 13951 36812 14036 37048
rect 14272 36812 14357 37048
rect 14593 36812 14678 37048
rect 14914 36812 14999 37048
rect 15235 36812 15320 37048
rect 15556 36812 16000 37048
rect 0 36724 16000 36812
rect 0 36488 215 36724
rect 451 36488 537 36724
rect 773 36488 859 36724
rect 1095 36488 1181 36724
rect 1417 36488 1503 36724
rect 1739 36488 1825 36724
rect 2061 36488 2147 36724
rect 2383 36488 2469 36724
rect 2705 36488 2791 36724
rect 3027 36488 3113 36724
rect 3349 36488 3435 36724
rect 3671 36488 3757 36724
rect 3993 36488 4079 36724
rect 4315 36488 4401 36724
rect 4637 36488 4723 36724
rect 4959 36488 5045 36724
rect 5281 36488 5367 36724
rect 5603 36488 5689 36724
rect 5925 36488 6011 36724
rect 6247 36488 6332 36724
rect 6568 36488 6653 36724
rect 6889 36488 6974 36724
rect 7210 36488 7295 36724
rect 7531 36488 7616 36724
rect 7852 36488 7937 36724
rect 8173 36488 8258 36724
rect 8494 36488 8579 36724
rect 8815 36488 8900 36724
rect 9136 36488 9221 36724
rect 9457 36488 9542 36724
rect 9778 36488 9863 36724
rect 10099 36488 10184 36724
rect 10420 36488 10505 36724
rect 10741 36488 10826 36724
rect 11062 36488 11147 36724
rect 11383 36488 11468 36724
rect 11704 36488 11789 36724
rect 12025 36488 12110 36724
rect 12346 36488 12431 36724
rect 12667 36488 12752 36724
rect 12988 36488 13073 36724
rect 13309 36488 13394 36724
rect 13630 36488 13715 36724
rect 13951 36488 14036 36724
rect 14272 36488 14357 36724
rect 14593 36488 14678 36724
rect 14914 36488 14999 36724
rect 15235 36488 15320 36724
rect 15556 36488 16000 36724
rect 0 36400 16000 36488
rect 0 36164 215 36400
rect 451 36164 537 36400
rect 773 36164 859 36400
rect 1095 36164 1181 36400
rect 1417 36164 1503 36400
rect 1739 36164 1825 36400
rect 2061 36164 2147 36400
rect 2383 36164 2469 36400
rect 2705 36164 2791 36400
rect 3027 36164 3113 36400
rect 3349 36164 3435 36400
rect 3671 36164 3757 36400
rect 3993 36164 4079 36400
rect 4315 36164 4401 36400
rect 4637 36164 4723 36400
rect 4959 36164 5045 36400
rect 5281 36164 5367 36400
rect 5603 36164 5689 36400
rect 5925 36164 6011 36400
rect 6247 36164 6332 36400
rect 6568 36164 6653 36400
rect 6889 36164 6974 36400
rect 7210 36164 7295 36400
rect 7531 36164 7616 36400
rect 7852 36164 7937 36400
rect 8173 36164 8258 36400
rect 8494 36164 8579 36400
rect 8815 36164 8900 36400
rect 9136 36164 9221 36400
rect 9457 36164 9542 36400
rect 9778 36164 9863 36400
rect 10099 36164 10184 36400
rect 10420 36164 10505 36400
rect 10741 36164 10826 36400
rect 11062 36164 11147 36400
rect 11383 36164 11468 36400
rect 11704 36164 11789 36400
rect 12025 36164 12110 36400
rect 12346 36164 12431 36400
rect 12667 36164 12752 36400
rect 12988 36164 13073 36400
rect 13309 36164 13394 36400
rect 13630 36164 13715 36400
rect 13951 36164 14036 36400
rect 14272 36164 14357 36400
rect 14593 36164 14678 36400
rect 14914 36164 14999 36400
rect 15235 36164 15320 36400
rect 15556 36164 16000 36400
rect 0 36076 16000 36164
rect 0 35840 215 36076
rect 451 35840 537 36076
rect 773 35840 859 36076
rect 1095 35840 1181 36076
rect 1417 35840 1503 36076
rect 1739 35840 1825 36076
rect 2061 35840 2147 36076
rect 2383 35840 2469 36076
rect 2705 35840 2791 36076
rect 3027 35840 3113 36076
rect 3349 35840 3435 36076
rect 3671 35840 3757 36076
rect 3993 35840 4079 36076
rect 4315 35840 4401 36076
rect 4637 35840 4723 36076
rect 4959 35840 5045 36076
rect 5281 35840 5367 36076
rect 5603 35840 5689 36076
rect 5925 35840 6011 36076
rect 6247 35840 6332 36076
rect 6568 35840 6653 36076
rect 6889 35840 6974 36076
rect 7210 35840 7295 36076
rect 7531 35840 7616 36076
rect 7852 35840 7937 36076
rect 8173 35840 8258 36076
rect 8494 35840 8579 36076
rect 8815 35840 8900 36076
rect 9136 35840 9221 36076
rect 9457 35840 9542 36076
rect 9778 35840 9863 36076
rect 10099 35840 10184 36076
rect 10420 35840 10505 36076
rect 10741 35840 10826 36076
rect 11062 35840 11147 36076
rect 11383 35840 11468 36076
rect 11704 35840 11789 36076
rect 12025 35840 12110 36076
rect 12346 35840 12431 36076
rect 12667 35840 12752 36076
rect 12988 35840 13073 36076
rect 13309 35840 13394 36076
rect 13630 35840 13715 36076
rect 13951 35840 14036 36076
rect 14272 35840 14357 36076
rect 14593 35840 14678 36076
rect 14914 35840 14999 36076
rect 15235 35840 15320 36076
rect 15556 35840 16000 36076
rect 0 35752 16000 35840
rect 0 35516 215 35752
rect 451 35516 537 35752
rect 773 35516 859 35752
rect 1095 35516 1181 35752
rect 1417 35516 1503 35752
rect 1739 35516 1825 35752
rect 2061 35516 2147 35752
rect 2383 35516 2469 35752
rect 2705 35516 2791 35752
rect 3027 35516 3113 35752
rect 3349 35516 3435 35752
rect 3671 35516 3757 35752
rect 3993 35516 4079 35752
rect 4315 35516 4401 35752
rect 4637 35516 4723 35752
rect 4959 35516 5045 35752
rect 5281 35516 5367 35752
rect 5603 35516 5689 35752
rect 5925 35516 6011 35752
rect 6247 35516 6332 35752
rect 6568 35516 6653 35752
rect 6889 35516 6974 35752
rect 7210 35516 7295 35752
rect 7531 35516 7616 35752
rect 7852 35516 7937 35752
rect 8173 35516 8258 35752
rect 8494 35516 8579 35752
rect 8815 35516 8900 35752
rect 9136 35516 9221 35752
rect 9457 35516 9542 35752
rect 9778 35516 9863 35752
rect 10099 35516 10184 35752
rect 10420 35516 10505 35752
rect 10741 35516 10826 35752
rect 11062 35516 11147 35752
rect 11383 35516 11468 35752
rect 11704 35516 11789 35752
rect 12025 35516 12110 35752
rect 12346 35516 12431 35752
rect 12667 35516 12752 35752
rect 12988 35516 13073 35752
rect 13309 35516 13394 35752
rect 13630 35516 13715 35752
rect 13951 35516 14036 35752
rect 14272 35516 14357 35752
rect 14593 35516 14678 35752
rect 14914 35516 14999 35752
rect 15235 35516 15320 35752
rect 15556 35516 16000 35752
rect 0 35428 16000 35516
rect 0 35192 215 35428
rect 451 35192 537 35428
rect 773 35192 859 35428
rect 1095 35192 1181 35428
rect 1417 35192 1503 35428
rect 1739 35192 1825 35428
rect 2061 35192 2147 35428
rect 2383 35192 2469 35428
rect 2705 35192 2791 35428
rect 3027 35192 3113 35428
rect 3349 35192 3435 35428
rect 3671 35192 3757 35428
rect 3993 35192 4079 35428
rect 4315 35192 4401 35428
rect 4637 35192 4723 35428
rect 4959 35192 5045 35428
rect 5281 35192 5367 35428
rect 5603 35192 5689 35428
rect 5925 35192 6011 35428
rect 6247 35192 6332 35428
rect 6568 35192 6653 35428
rect 6889 35192 6974 35428
rect 7210 35192 7295 35428
rect 7531 35192 7616 35428
rect 7852 35192 7937 35428
rect 8173 35192 8258 35428
rect 8494 35192 8579 35428
rect 8815 35192 8900 35428
rect 9136 35192 9221 35428
rect 9457 35192 9542 35428
rect 9778 35192 9863 35428
rect 10099 35192 10184 35428
rect 10420 35192 10505 35428
rect 10741 35192 10826 35428
rect 11062 35192 11147 35428
rect 11383 35192 11468 35428
rect 11704 35192 11789 35428
rect 12025 35192 12110 35428
rect 12346 35192 12431 35428
rect 12667 35192 12752 35428
rect 12988 35192 13073 35428
rect 13309 35192 13394 35428
rect 13630 35192 13715 35428
rect 13951 35192 14036 35428
rect 14272 35192 14357 35428
rect 14593 35192 14678 35428
rect 14914 35192 14999 35428
rect 15235 35192 15320 35428
rect 15556 35192 16000 35428
rect 0 35157 16000 35192
rect 0 18972 16000 19000
rect 0 18736 215 18972
rect 451 18736 538 18972
rect 774 18736 861 18972
rect 1097 18736 1184 18972
rect 1420 18736 1507 18972
rect 1743 18736 1830 18972
rect 2066 18736 2153 18972
rect 2389 18736 2476 18972
rect 2712 18736 2799 18972
rect 3035 18736 3122 18972
rect 3358 18736 3445 18972
rect 3681 18736 3768 18972
rect 4004 18736 4091 18972
rect 4327 18736 4414 18972
rect 4650 18736 4737 18972
rect 4973 18736 5060 18972
rect 5296 18736 5383 18972
rect 5619 18736 5706 18972
rect 5942 18736 6029 18972
rect 6265 18736 6351 18972
rect 6587 18736 6673 18972
rect 6909 18736 6995 18972
rect 7231 18736 7317 18972
rect 7553 18736 7639 18972
rect 7875 18736 7961 18972
rect 8197 18736 8283 18972
rect 8519 18736 8605 18972
rect 8841 18736 8927 18972
rect 9163 18736 9249 18972
rect 9485 18736 9571 18972
rect 9807 18736 9893 18972
rect 10129 18736 10215 18972
rect 10451 18736 10537 18972
rect 10773 18736 10859 18972
rect 11095 18736 11181 18972
rect 11417 18736 11503 18972
rect 11739 18736 11825 18972
rect 12061 18736 12147 18972
rect 12383 18736 12469 18972
rect 12705 18736 12791 18972
rect 13027 18736 13113 18972
rect 13349 18736 13435 18972
rect 13671 18736 13757 18972
rect 13993 18736 14079 18972
rect 14315 18736 14401 18972
rect 14637 18736 14723 18972
rect 14959 18736 15045 18972
rect 15281 18736 15367 18972
rect 15603 18736 16000 18972
rect 0 18636 16000 18736
rect 0 18400 215 18636
rect 451 18400 538 18636
rect 774 18400 861 18636
rect 1097 18400 1184 18636
rect 1420 18400 1507 18636
rect 1743 18400 1830 18636
rect 2066 18400 2153 18636
rect 2389 18400 2476 18636
rect 2712 18400 2799 18636
rect 3035 18400 3122 18636
rect 3358 18400 3445 18636
rect 3681 18400 3768 18636
rect 4004 18400 4091 18636
rect 4327 18400 4414 18636
rect 4650 18400 4737 18636
rect 4973 18400 5060 18636
rect 5296 18400 5383 18636
rect 5619 18400 5706 18636
rect 5942 18400 6029 18636
rect 6265 18400 6351 18636
rect 6587 18400 6673 18636
rect 6909 18400 6995 18636
rect 7231 18400 7317 18636
rect 7553 18400 7639 18636
rect 7875 18400 7961 18636
rect 8197 18400 8283 18636
rect 8519 18400 8605 18636
rect 8841 18400 8927 18636
rect 9163 18400 9249 18636
rect 9485 18400 9571 18636
rect 9807 18400 9893 18636
rect 10129 18400 10215 18636
rect 10451 18400 10537 18636
rect 10773 18400 10859 18636
rect 11095 18400 11181 18636
rect 11417 18400 11503 18636
rect 11739 18400 11825 18636
rect 12061 18400 12147 18636
rect 12383 18400 12469 18636
rect 12705 18400 12791 18636
rect 13027 18400 13113 18636
rect 13349 18400 13435 18636
rect 13671 18400 13757 18636
rect 13993 18400 14079 18636
rect 14315 18400 14401 18636
rect 14637 18400 14723 18636
rect 14959 18400 15045 18636
rect 15281 18400 15367 18636
rect 15603 18400 16000 18636
rect 0 18300 16000 18400
rect 0 18064 215 18300
rect 451 18064 538 18300
rect 774 18064 861 18300
rect 1097 18064 1184 18300
rect 1420 18064 1507 18300
rect 1743 18064 1830 18300
rect 2066 18064 2153 18300
rect 2389 18064 2476 18300
rect 2712 18064 2799 18300
rect 3035 18064 3122 18300
rect 3358 18064 3445 18300
rect 3681 18064 3768 18300
rect 4004 18064 4091 18300
rect 4327 18064 4414 18300
rect 4650 18064 4737 18300
rect 4973 18064 5060 18300
rect 5296 18064 5383 18300
rect 5619 18064 5706 18300
rect 5942 18064 6029 18300
rect 6265 18064 6351 18300
rect 6587 18064 6673 18300
rect 6909 18064 6995 18300
rect 7231 18064 7317 18300
rect 7553 18064 7639 18300
rect 7875 18064 7961 18300
rect 8197 18064 8283 18300
rect 8519 18064 8605 18300
rect 8841 18064 8927 18300
rect 9163 18064 9249 18300
rect 9485 18064 9571 18300
rect 9807 18064 9893 18300
rect 10129 18064 10215 18300
rect 10451 18064 10537 18300
rect 10773 18064 10859 18300
rect 11095 18064 11181 18300
rect 11417 18064 11503 18300
rect 11739 18064 11825 18300
rect 12061 18064 12147 18300
rect 12383 18064 12469 18300
rect 12705 18064 12791 18300
rect 13027 18064 13113 18300
rect 13349 18064 13435 18300
rect 13671 18064 13757 18300
rect 13993 18064 14079 18300
rect 14315 18064 14401 18300
rect 14637 18064 14723 18300
rect 14959 18064 15045 18300
rect 15281 18064 15367 18300
rect 15603 18064 16000 18300
rect 0 17964 16000 18064
rect 0 17728 215 17964
rect 451 17728 538 17964
rect 774 17728 861 17964
rect 1097 17728 1184 17964
rect 1420 17728 1507 17964
rect 1743 17728 1830 17964
rect 2066 17728 2153 17964
rect 2389 17728 2476 17964
rect 2712 17728 2799 17964
rect 3035 17728 3122 17964
rect 3358 17728 3445 17964
rect 3681 17728 3768 17964
rect 4004 17728 4091 17964
rect 4327 17728 4414 17964
rect 4650 17728 4737 17964
rect 4973 17728 5060 17964
rect 5296 17728 5383 17964
rect 5619 17728 5706 17964
rect 5942 17728 6029 17964
rect 6265 17728 6351 17964
rect 6587 17728 6673 17964
rect 6909 17728 6995 17964
rect 7231 17728 7317 17964
rect 7553 17728 7639 17964
rect 7875 17728 7961 17964
rect 8197 17728 8283 17964
rect 8519 17728 8605 17964
rect 8841 17728 8927 17964
rect 9163 17728 9249 17964
rect 9485 17728 9571 17964
rect 9807 17728 9893 17964
rect 10129 17728 10215 17964
rect 10451 17728 10537 17964
rect 10773 17728 10859 17964
rect 11095 17728 11181 17964
rect 11417 17728 11503 17964
rect 11739 17728 11825 17964
rect 12061 17728 12147 17964
rect 12383 17728 12469 17964
rect 12705 17728 12791 17964
rect 13027 17728 13113 17964
rect 13349 17728 13435 17964
rect 13671 17728 13757 17964
rect 13993 17728 14079 17964
rect 14315 17728 14401 17964
rect 14637 17728 14723 17964
rect 14959 17728 15045 17964
rect 15281 17728 15367 17964
rect 15603 17728 16000 17964
rect 0 17628 16000 17728
rect 0 17392 215 17628
rect 451 17392 538 17628
rect 774 17392 861 17628
rect 1097 17392 1184 17628
rect 1420 17392 1507 17628
rect 1743 17392 1830 17628
rect 2066 17392 2153 17628
rect 2389 17392 2476 17628
rect 2712 17392 2799 17628
rect 3035 17392 3122 17628
rect 3358 17392 3445 17628
rect 3681 17392 3768 17628
rect 4004 17392 4091 17628
rect 4327 17392 4414 17628
rect 4650 17392 4737 17628
rect 4973 17392 5060 17628
rect 5296 17392 5383 17628
rect 5619 17392 5706 17628
rect 5942 17392 6029 17628
rect 6265 17392 6351 17628
rect 6587 17392 6673 17628
rect 6909 17392 6995 17628
rect 7231 17392 7317 17628
rect 7553 17392 7639 17628
rect 7875 17392 7961 17628
rect 8197 17392 8283 17628
rect 8519 17392 8605 17628
rect 8841 17392 8927 17628
rect 9163 17392 9249 17628
rect 9485 17392 9571 17628
rect 9807 17392 9893 17628
rect 10129 17392 10215 17628
rect 10451 17392 10537 17628
rect 10773 17392 10859 17628
rect 11095 17392 11181 17628
rect 11417 17392 11503 17628
rect 11739 17392 11825 17628
rect 12061 17392 12147 17628
rect 12383 17392 12469 17628
rect 12705 17392 12791 17628
rect 13027 17392 13113 17628
rect 13349 17392 13435 17628
rect 13671 17392 13757 17628
rect 13993 17392 14079 17628
rect 14315 17392 14401 17628
rect 14637 17392 14723 17628
rect 14959 17392 15045 17628
rect 15281 17392 15367 17628
rect 15603 17392 16000 17628
rect 0 17292 16000 17392
rect 0 17056 215 17292
rect 451 17056 538 17292
rect 774 17056 861 17292
rect 1097 17056 1184 17292
rect 1420 17056 1507 17292
rect 1743 17056 1830 17292
rect 2066 17056 2153 17292
rect 2389 17056 2476 17292
rect 2712 17056 2799 17292
rect 3035 17056 3122 17292
rect 3358 17056 3445 17292
rect 3681 17056 3768 17292
rect 4004 17056 4091 17292
rect 4327 17056 4414 17292
rect 4650 17056 4737 17292
rect 4973 17056 5060 17292
rect 5296 17056 5383 17292
rect 5619 17056 5706 17292
rect 5942 17056 6029 17292
rect 6265 17056 6351 17292
rect 6587 17056 6673 17292
rect 6909 17056 6995 17292
rect 7231 17056 7317 17292
rect 7553 17056 7639 17292
rect 7875 17056 7961 17292
rect 8197 17056 8283 17292
rect 8519 17056 8605 17292
rect 8841 17056 8927 17292
rect 9163 17056 9249 17292
rect 9485 17056 9571 17292
rect 9807 17056 9893 17292
rect 10129 17056 10215 17292
rect 10451 17056 10537 17292
rect 10773 17056 10859 17292
rect 11095 17056 11181 17292
rect 11417 17056 11503 17292
rect 11739 17056 11825 17292
rect 12061 17056 12147 17292
rect 12383 17056 12469 17292
rect 12705 17056 12791 17292
rect 13027 17056 13113 17292
rect 13349 17056 13435 17292
rect 13671 17056 13757 17292
rect 13993 17056 14079 17292
rect 14315 17056 14401 17292
rect 14637 17056 14723 17292
rect 14959 17056 15045 17292
rect 15281 17056 15367 17292
rect 15603 17056 16000 17292
rect 0 16956 16000 17056
rect 0 16720 215 16956
rect 451 16720 538 16956
rect 774 16720 861 16956
rect 1097 16720 1184 16956
rect 1420 16720 1507 16956
rect 1743 16720 1830 16956
rect 2066 16720 2153 16956
rect 2389 16720 2476 16956
rect 2712 16720 2799 16956
rect 3035 16720 3122 16956
rect 3358 16720 3445 16956
rect 3681 16720 3768 16956
rect 4004 16720 4091 16956
rect 4327 16720 4414 16956
rect 4650 16720 4737 16956
rect 4973 16720 5060 16956
rect 5296 16720 5383 16956
rect 5619 16720 5706 16956
rect 5942 16720 6029 16956
rect 6265 16720 6351 16956
rect 6587 16720 6673 16956
rect 6909 16720 6995 16956
rect 7231 16720 7317 16956
rect 7553 16720 7639 16956
rect 7875 16720 7961 16956
rect 8197 16720 8283 16956
rect 8519 16720 8605 16956
rect 8841 16720 8927 16956
rect 9163 16720 9249 16956
rect 9485 16720 9571 16956
rect 9807 16720 9893 16956
rect 10129 16720 10215 16956
rect 10451 16720 10537 16956
rect 10773 16720 10859 16956
rect 11095 16720 11181 16956
rect 11417 16720 11503 16956
rect 11739 16720 11825 16956
rect 12061 16720 12147 16956
rect 12383 16720 12469 16956
rect 12705 16720 12791 16956
rect 13027 16720 13113 16956
rect 13349 16720 13435 16956
rect 13671 16720 13757 16956
rect 13993 16720 14079 16956
rect 14315 16720 14401 16956
rect 14637 16720 14723 16956
rect 14959 16720 15045 16956
rect 15281 16720 15367 16956
rect 15603 16720 16000 16956
rect 0 16620 16000 16720
rect 0 16384 215 16620
rect 451 16384 538 16620
rect 774 16384 861 16620
rect 1097 16384 1184 16620
rect 1420 16384 1507 16620
rect 1743 16384 1830 16620
rect 2066 16384 2153 16620
rect 2389 16384 2476 16620
rect 2712 16384 2799 16620
rect 3035 16384 3122 16620
rect 3358 16384 3445 16620
rect 3681 16384 3768 16620
rect 4004 16384 4091 16620
rect 4327 16384 4414 16620
rect 4650 16384 4737 16620
rect 4973 16384 5060 16620
rect 5296 16384 5383 16620
rect 5619 16384 5706 16620
rect 5942 16384 6029 16620
rect 6265 16384 6351 16620
rect 6587 16384 6673 16620
rect 6909 16384 6995 16620
rect 7231 16384 7317 16620
rect 7553 16384 7639 16620
rect 7875 16384 7961 16620
rect 8197 16384 8283 16620
rect 8519 16384 8605 16620
rect 8841 16384 8927 16620
rect 9163 16384 9249 16620
rect 9485 16384 9571 16620
rect 9807 16384 9893 16620
rect 10129 16384 10215 16620
rect 10451 16384 10537 16620
rect 10773 16384 10859 16620
rect 11095 16384 11181 16620
rect 11417 16384 11503 16620
rect 11739 16384 11825 16620
rect 12061 16384 12147 16620
rect 12383 16384 12469 16620
rect 12705 16384 12791 16620
rect 13027 16384 13113 16620
rect 13349 16384 13435 16620
rect 13671 16384 13757 16620
rect 13993 16384 14079 16620
rect 14315 16384 14401 16620
rect 14637 16384 14723 16620
rect 14959 16384 15045 16620
rect 15281 16384 15367 16620
rect 15603 16384 16000 16620
rect 0 16284 16000 16384
rect 0 16048 215 16284
rect 451 16048 538 16284
rect 774 16048 861 16284
rect 1097 16048 1184 16284
rect 1420 16048 1507 16284
rect 1743 16048 1830 16284
rect 2066 16048 2153 16284
rect 2389 16048 2476 16284
rect 2712 16048 2799 16284
rect 3035 16048 3122 16284
rect 3358 16048 3445 16284
rect 3681 16048 3768 16284
rect 4004 16048 4091 16284
rect 4327 16048 4414 16284
rect 4650 16048 4737 16284
rect 4973 16048 5060 16284
rect 5296 16048 5383 16284
rect 5619 16048 5706 16284
rect 5942 16048 6029 16284
rect 6265 16048 6351 16284
rect 6587 16048 6673 16284
rect 6909 16048 6995 16284
rect 7231 16048 7317 16284
rect 7553 16048 7639 16284
rect 7875 16048 7961 16284
rect 8197 16048 8283 16284
rect 8519 16048 8605 16284
rect 8841 16048 8927 16284
rect 9163 16048 9249 16284
rect 9485 16048 9571 16284
rect 9807 16048 9893 16284
rect 10129 16048 10215 16284
rect 10451 16048 10537 16284
rect 10773 16048 10859 16284
rect 11095 16048 11181 16284
rect 11417 16048 11503 16284
rect 11739 16048 11825 16284
rect 12061 16048 12147 16284
rect 12383 16048 12469 16284
rect 12705 16048 12791 16284
rect 13027 16048 13113 16284
rect 13349 16048 13435 16284
rect 13671 16048 13757 16284
rect 13993 16048 14079 16284
rect 14315 16048 14401 16284
rect 14637 16048 14723 16284
rect 14959 16048 15045 16284
rect 15281 16048 15367 16284
rect 15603 16048 16000 16284
rect 0 15948 16000 16048
rect 0 15712 215 15948
rect 451 15712 538 15948
rect 774 15712 861 15948
rect 1097 15712 1184 15948
rect 1420 15712 1507 15948
rect 1743 15712 1830 15948
rect 2066 15712 2153 15948
rect 2389 15712 2476 15948
rect 2712 15712 2799 15948
rect 3035 15712 3122 15948
rect 3358 15712 3445 15948
rect 3681 15712 3768 15948
rect 4004 15712 4091 15948
rect 4327 15712 4414 15948
rect 4650 15712 4737 15948
rect 4973 15712 5060 15948
rect 5296 15712 5383 15948
rect 5619 15712 5706 15948
rect 5942 15712 6029 15948
rect 6265 15712 6351 15948
rect 6587 15712 6673 15948
rect 6909 15712 6995 15948
rect 7231 15712 7317 15948
rect 7553 15712 7639 15948
rect 7875 15712 7961 15948
rect 8197 15712 8283 15948
rect 8519 15712 8605 15948
rect 8841 15712 8927 15948
rect 9163 15712 9249 15948
rect 9485 15712 9571 15948
rect 9807 15712 9893 15948
rect 10129 15712 10215 15948
rect 10451 15712 10537 15948
rect 10773 15712 10859 15948
rect 11095 15712 11181 15948
rect 11417 15712 11503 15948
rect 11739 15712 11825 15948
rect 12061 15712 12147 15948
rect 12383 15712 12469 15948
rect 12705 15712 12791 15948
rect 13027 15712 13113 15948
rect 13349 15712 13435 15948
rect 13671 15712 13757 15948
rect 13993 15712 14079 15948
rect 14315 15712 14401 15948
rect 14637 15712 14723 15948
rect 14959 15712 15045 15948
rect 15281 15712 15367 15948
rect 15603 15712 16000 15948
rect 0 15612 16000 15712
rect 0 15376 215 15612
rect 451 15376 538 15612
rect 774 15376 861 15612
rect 1097 15376 1184 15612
rect 1420 15376 1507 15612
rect 1743 15376 1830 15612
rect 2066 15376 2153 15612
rect 2389 15376 2476 15612
rect 2712 15376 2799 15612
rect 3035 15376 3122 15612
rect 3358 15376 3445 15612
rect 3681 15376 3768 15612
rect 4004 15376 4091 15612
rect 4327 15376 4414 15612
rect 4650 15376 4737 15612
rect 4973 15376 5060 15612
rect 5296 15376 5383 15612
rect 5619 15376 5706 15612
rect 5942 15376 6029 15612
rect 6265 15376 6351 15612
rect 6587 15376 6673 15612
rect 6909 15376 6995 15612
rect 7231 15376 7317 15612
rect 7553 15376 7639 15612
rect 7875 15376 7961 15612
rect 8197 15376 8283 15612
rect 8519 15376 8605 15612
rect 8841 15376 8927 15612
rect 9163 15376 9249 15612
rect 9485 15376 9571 15612
rect 9807 15376 9893 15612
rect 10129 15376 10215 15612
rect 10451 15376 10537 15612
rect 10773 15376 10859 15612
rect 11095 15376 11181 15612
rect 11417 15376 11503 15612
rect 11739 15376 11825 15612
rect 12061 15376 12147 15612
rect 12383 15376 12469 15612
rect 12705 15376 12791 15612
rect 13027 15376 13113 15612
rect 13349 15376 13435 15612
rect 13671 15376 13757 15612
rect 13993 15376 14079 15612
rect 14315 15376 14401 15612
rect 14637 15376 14723 15612
rect 14959 15376 15045 15612
rect 15281 15376 15367 15612
rect 15603 15376 16000 15612
rect 0 15276 16000 15376
rect 0 15040 215 15276
rect 451 15040 538 15276
rect 774 15040 861 15276
rect 1097 15040 1184 15276
rect 1420 15040 1507 15276
rect 1743 15040 1830 15276
rect 2066 15040 2153 15276
rect 2389 15040 2476 15276
rect 2712 15040 2799 15276
rect 3035 15040 3122 15276
rect 3358 15040 3445 15276
rect 3681 15040 3768 15276
rect 4004 15040 4091 15276
rect 4327 15040 4414 15276
rect 4650 15040 4737 15276
rect 4973 15040 5060 15276
rect 5296 15040 5383 15276
rect 5619 15040 5706 15276
rect 5942 15040 6029 15276
rect 6265 15040 6351 15276
rect 6587 15040 6673 15276
rect 6909 15040 6995 15276
rect 7231 15040 7317 15276
rect 7553 15040 7639 15276
rect 7875 15040 7961 15276
rect 8197 15040 8283 15276
rect 8519 15040 8605 15276
rect 8841 15040 8927 15276
rect 9163 15040 9249 15276
rect 9485 15040 9571 15276
rect 9807 15040 9893 15276
rect 10129 15040 10215 15276
rect 10451 15040 10537 15276
rect 10773 15040 10859 15276
rect 11095 15040 11181 15276
rect 11417 15040 11503 15276
rect 11739 15040 11825 15276
rect 12061 15040 12147 15276
rect 12383 15040 12469 15276
rect 12705 15040 12791 15276
rect 13027 15040 13113 15276
rect 13349 15040 13435 15276
rect 13671 15040 13757 15276
rect 13993 15040 14079 15276
rect 14315 15040 14401 15276
rect 14637 15040 14723 15276
rect 14959 15040 15045 15276
rect 15281 15040 15367 15276
rect 15603 15040 16000 15276
rect 0 14940 16000 15040
rect 0 14704 215 14940
rect 451 14704 538 14940
rect 774 14704 861 14940
rect 1097 14704 1184 14940
rect 1420 14704 1507 14940
rect 1743 14704 1830 14940
rect 2066 14704 2153 14940
rect 2389 14704 2476 14940
rect 2712 14704 2799 14940
rect 3035 14704 3122 14940
rect 3358 14704 3445 14940
rect 3681 14704 3768 14940
rect 4004 14704 4091 14940
rect 4327 14704 4414 14940
rect 4650 14704 4737 14940
rect 4973 14704 5060 14940
rect 5296 14704 5383 14940
rect 5619 14704 5706 14940
rect 5942 14704 6029 14940
rect 6265 14704 6351 14940
rect 6587 14704 6673 14940
rect 6909 14704 6995 14940
rect 7231 14704 7317 14940
rect 7553 14704 7639 14940
rect 7875 14704 7961 14940
rect 8197 14704 8283 14940
rect 8519 14704 8605 14940
rect 8841 14704 8927 14940
rect 9163 14704 9249 14940
rect 9485 14704 9571 14940
rect 9807 14704 9893 14940
rect 10129 14704 10215 14940
rect 10451 14704 10537 14940
rect 10773 14704 10859 14940
rect 11095 14704 11181 14940
rect 11417 14704 11503 14940
rect 11739 14704 11825 14940
rect 12061 14704 12147 14940
rect 12383 14704 12469 14940
rect 12705 14704 12791 14940
rect 13027 14704 13113 14940
rect 13349 14704 13435 14940
rect 13671 14704 13757 14940
rect 13993 14704 14079 14940
rect 14315 14704 14401 14940
rect 14637 14704 14723 14940
rect 14959 14704 15045 14940
rect 15281 14704 15367 14940
rect 15603 14704 16000 14940
rect 0 14604 16000 14704
rect 0 14368 215 14604
rect 451 14368 538 14604
rect 774 14368 861 14604
rect 1097 14368 1184 14604
rect 1420 14368 1507 14604
rect 1743 14368 1830 14604
rect 2066 14368 2153 14604
rect 2389 14368 2476 14604
rect 2712 14368 2799 14604
rect 3035 14368 3122 14604
rect 3358 14368 3445 14604
rect 3681 14368 3768 14604
rect 4004 14368 4091 14604
rect 4327 14368 4414 14604
rect 4650 14368 4737 14604
rect 4973 14368 5060 14604
rect 5296 14368 5383 14604
rect 5619 14368 5706 14604
rect 5942 14368 6029 14604
rect 6265 14368 6351 14604
rect 6587 14368 6673 14604
rect 6909 14368 6995 14604
rect 7231 14368 7317 14604
rect 7553 14368 7639 14604
rect 7875 14368 7961 14604
rect 8197 14368 8283 14604
rect 8519 14368 8605 14604
rect 8841 14368 8927 14604
rect 9163 14368 9249 14604
rect 9485 14368 9571 14604
rect 9807 14368 9893 14604
rect 10129 14368 10215 14604
rect 10451 14368 10537 14604
rect 10773 14368 10859 14604
rect 11095 14368 11181 14604
rect 11417 14368 11503 14604
rect 11739 14368 11825 14604
rect 12061 14368 12147 14604
rect 12383 14368 12469 14604
rect 12705 14368 12791 14604
rect 13027 14368 13113 14604
rect 13349 14368 13435 14604
rect 13671 14368 13757 14604
rect 13993 14368 14079 14604
rect 14315 14368 14401 14604
rect 14637 14368 14723 14604
rect 14959 14368 15045 14604
rect 15281 14368 15367 14604
rect 15603 14368 16000 14604
rect 0 14268 16000 14368
rect 0 14032 215 14268
rect 451 14032 538 14268
rect 774 14032 861 14268
rect 1097 14032 1184 14268
rect 1420 14032 1507 14268
rect 1743 14032 1830 14268
rect 2066 14032 2153 14268
rect 2389 14032 2476 14268
rect 2712 14032 2799 14268
rect 3035 14032 3122 14268
rect 3358 14032 3445 14268
rect 3681 14032 3768 14268
rect 4004 14032 4091 14268
rect 4327 14032 4414 14268
rect 4650 14032 4737 14268
rect 4973 14032 5060 14268
rect 5296 14032 5383 14268
rect 5619 14032 5706 14268
rect 5942 14032 6029 14268
rect 6265 14032 6351 14268
rect 6587 14032 6673 14268
rect 6909 14032 6995 14268
rect 7231 14032 7317 14268
rect 7553 14032 7639 14268
rect 7875 14032 7961 14268
rect 8197 14032 8283 14268
rect 8519 14032 8605 14268
rect 8841 14032 8927 14268
rect 9163 14032 9249 14268
rect 9485 14032 9571 14268
rect 9807 14032 9893 14268
rect 10129 14032 10215 14268
rect 10451 14032 10537 14268
rect 10773 14032 10859 14268
rect 11095 14032 11181 14268
rect 11417 14032 11503 14268
rect 11739 14032 11825 14268
rect 12061 14032 12147 14268
rect 12383 14032 12469 14268
rect 12705 14032 12791 14268
rect 13027 14032 13113 14268
rect 13349 14032 13435 14268
rect 13671 14032 13757 14268
rect 13993 14032 14079 14268
rect 14315 14032 14401 14268
rect 14637 14032 14723 14268
rect 14959 14032 15045 14268
rect 15281 14032 15367 14268
rect 15603 14032 16000 14268
rect 0 14007 16000 14032
rect 0 13701 16000 13707
rect 0 13663 8333 13701
rect 8397 13663 8417 13701
rect 8481 13663 8501 13701
rect 0 13427 216 13663
rect 452 13427 538 13663
rect 774 13427 860 13663
rect 1096 13427 1182 13663
rect 1418 13427 1504 13663
rect 1740 13427 1826 13663
rect 2062 13427 2148 13663
rect 2384 13427 2470 13663
rect 2706 13427 2792 13663
rect 3028 13427 3114 13663
rect 3350 13427 3436 13663
rect 3672 13427 3758 13663
rect 3994 13427 4080 13663
rect 4316 13427 4402 13663
rect 4638 13427 4724 13663
rect 4960 13427 5046 13663
rect 5282 13427 5368 13663
rect 5604 13427 5690 13663
rect 5926 13427 6012 13663
rect 6248 13427 6333 13663
rect 6569 13427 6654 13663
rect 6890 13427 6975 13663
rect 7211 13427 7296 13663
rect 7532 13427 7617 13663
rect 7853 13427 7938 13663
rect 8174 13427 8259 13663
rect 8495 13637 8501 13663
rect 8565 13663 8585 13701
rect 8649 13663 8669 13701
rect 8733 13663 16000 13701
rect 8565 13637 8580 13663
rect 8495 13620 8580 13637
rect 8495 13556 8501 13620
rect 8565 13556 8580 13620
rect 8495 13539 8580 13556
rect 8495 13475 8501 13539
rect 8565 13475 8580 13539
rect 8495 13458 8580 13475
rect 8495 13427 8501 13458
rect 0 13394 8333 13427
rect 8397 13394 8417 13427
rect 8481 13394 8501 13427
rect 8565 13427 8580 13458
rect 8816 13427 8901 13663
rect 9137 13427 9222 13663
rect 9458 13427 9543 13663
rect 9779 13427 9864 13663
rect 10100 13427 10185 13663
rect 10421 13427 10506 13663
rect 10742 13427 10827 13663
rect 11063 13427 11148 13663
rect 11384 13427 11469 13663
rect 11705 13427 11790 13663
rect 12026 13427 12111 13663
rect 12347 13427 12432 13663
rect 12668 13427 12753 13663
rect 12989 13427 13074 13663
rect 13310 13427 13395 13663
rect 13631 13427 13716 13663
rect 13952 13427 14037 13663
rect 14273 13427 14358 13663
rect 14594 13427 14679 13663
rect 14915 13427 15000 13663
rect 15236 13427 15321 13663
rect 15557 13427 16000 13663
rect 8565 13394 8585 13427
rect 8649 13394 8669 13427
rect 8733 13394 16000 13427
rect 0 13377 16000 13394
rect 0 13313 8333 13377
rect 8397 13313 8417 13377
rect 8481 13313 8501 13377
rect 8565 13313 8585 13377
rect 8649 13313 8669 13377
rect 8733 13313 16000 13377
rect 0 13296 16000 13313
rect 0 13232 8333 13296
rect 8397 13232 8417 13296
rect 8481 13232 8501 13296
rect 8565 13232 8585 13296
rect 8649 13232 8669 13296
rect 8733 13232 16000 13296
rect 0 13215 16000 13232
rect 0 13151 8333 13215
rect 8397 13151 8417 13215
rect 8481 13151 8501 13215
rect 8565 13151 8585 13215
rect 8649 13151 8669 13215
rect 8733 13151 16000 13215
rect 0 13133 16000 13151
rect 0 13097 8333 13133
rect 8397 13097 8417 13133
rect 8481 13097 8501 13133
rect 0 12861 216 13097
rect 452 12861 538 13097
rect 774 12861 860 13097
rect 1096 12861 1182 13097
rect 1418 12861 1504 13097
rect 1740 12861 1826 13097
rect 2062 12861 2148 13097
rect 2384 12861 2470 13097
rect 2706 12861 2792 13097
rect 3028 12861 3114 13097
rect 3350 12861 3436 13097
rect 3672 12861 3758 13097
rect 3994 12861 4080 13097
rect 4316 12861 4402 13097
rect 4638 12861 4724 13097
rect 4960 12861 5046 13097
rect 5282 12861 5368 13097
rect 5604 12861 5690 13097
rect 5926 12861 6012 13097
rect 6248 12861 6333 13097
rect 6569 12861 6654 13097
rect 6890 12861 6975 13097
rect 7211 12861 7296 13097
rect 7532 12861 7617 13097
rect 7853 12861 7938 13097
rect 8174 12861 8259 13097
rect 8495 13069 8501 13097
rect 8565 13097 8585 13133
rect 8649 13097 8669 13133
rect 8733 13097 16000 13133
rect 8565 13069 8580 13097
rect 8495 13051 8580 13069
rect 8495 12987 8501 13051
rect 8565 12987 8580 13051
rect 8495 12969 8580 12987
rect 8495 12905 8501 12969
rect 8565 12905 8580 12969
rect 8495 12887 8580 12905
rect 8495 12861 8501 12887
rect 0 12823 8333 12861
rect 8397 12823 8417 12861
rect 8481 12823 8501 12861
rect 8565 12861 8580 12887
rect 8816 12861 8901 13097
rect 9137 12861 9222 13097
rect 9458 12861 9543 13097
rect 9779 12861 9864 13097
rect 10100 12861 10185 13097
rect 10421 12861 10506 13097
rect 10742 12861 10827 13097
rect 11063 12861 11148 13097
rect 11384 12861 11469 13097
rect 11705 12861 11790 13097
rect 12026 12861 12111 13097
rect 12347 12861 12432 13097
rect 12668 12861 12753 13097
rect 12989 12861 13074 13097
rect 13310 12861 13395 13097
rect 13631 12861 13716 13097
rect 13952 12861 14037 13097
rect 14273 12861 14358 13097
rect 14594 12861 14679 13097
rect 14915 12861 15000 13097
rect 15236 12861 15321 13097
rect 15557 12861 16000 13097
rect 8565 12823 8585 12861
rect 8649 12823 8669 12861
rect 8733 12823 16000 12861
rect 0 12817 16000 12823
rect 0 12493 16000 12537
rect 0 12257 215 12493
rect 451 12257 537 12493
rect 773 12257 859 12493
rect 1095 12257 1181 12493
rect 1417 12257 1503 12493
rect 1739 12257 1825 12493
rect 2061 12257 2147 12493
rect 2383 12257 2469 12493
rect 2705 12257 2791 12493
rect 3027 12257 3113 12493
rect 3349 12257 3435 12493
rect 3671 12257 3757 12493
rect 3993 12257 4079 12493
rect 4315 12257 4401 12493
rect 4637 12257 4723 12493
rect 4959 12257 5045 12493
rect 5281 12257 5367 12493
rect 5603 12257 5689 12493
rect 5925 12257 6011 12493
rect 6247 12257 6332 12493
rect 6568 12257 6653 12493
rect 6889 12257 6974 12493
rect 7210 12257 7295 12493
rect 7531 12257 7616 12493
rect 7852 12257 7937 12493
rect 8173 12257 8258 12493
rect 8494 12257 8579 12493
rect 8815 12257 8900 12493
rect 9136 12257 9221 12493
rect 9457 12257 9542 12493
rect 9778 12257 9863 12493
rect 10099 12257 10184 12493
rect 10420 12257 10505 12493
rect 10741 12257 10826 12493
rect 11062 12257 11147 12493
rect 11383 12257 11468 12493
rect 11704 12257 11789 12493
rect 12025 12257 12110 12493
rect 12346 12257 12431 12493
rect 12667 12257 12752 12493
rect 12988 12257 13073 12493
rect 13309 12257 13394 12493
rect 13630 12257 13715 12493
rect 13951 12257 14036 12493
rect 14272 12257 14357 12493
rect 14593 12257 14678 12493
rect 14914 12257 14999 12493
rect 15235 12257 15320 12493
rect 15556 12257 16000 12493
rect 0 11927 16000 12257
rect 0 11691 215 11927
rect 451 11691 537 11927
rect 773 11691 859 11927
rect 1095 11691 1181 11927
rect 1417 11691 1503 11927
rect 1739 11691 1825 11927
rect 2061 11691 2147 11927
rect 2383 11691 2469 11927
rect 2705 11691 2791 11927
rect 3027 11691 3113 11927
rect 3349 11691 3435 11927
rect 3671 11691 3757 11927
rect 3993 11691 4079 11927
rect 4315 11691 4401 11927
rect 4637 11691 4723 11927
rect 4959 11691 5045 11927
rect 5281 11691 5367 11927
rect 5603 11691 5689 11927
rect 5925 11691 6011 11927
rect 6247 11691 6332 11927
rect 6568 11691 6653 11927
rect 6889 11691 6974 11927
rect 7210 11691 7295 11927
rect 7531 11691 7616 11927
rect 7852 11691 7937 11927
rect 8173 11691 8258 11927
rect 8494 11691 8579 11927
rect 8815 11691 8900 11927
rect 9136 11691 9221 11927
rect 9457 11691 9542 11927
rect 9778 11691 9863 11927
rect 10099 11691 10184 11927
rect 10420 11691 10505 11927
rect 10741 11691 10826 11927
rect 11062 11691 11147 11927
rect 11383 11691 11468 11927
rect 11704 11691 11789 11927
rect 12025 11691 12110 11927
rect 12346 11691 12431 11927
rect 12667 11691 12752 11927
rect 12988 11691 13073 11927
rect 13309 11691 13394 11927
rect 13630 11691 13715 11927
rect 13951 11691 14036 11927
rect 14272 11691 14357 11927
rect 14593 11691 14678 11927
rect 14914 11691 14999 11927
rect 15235 11691 15320 11927
rect 15556 11691 16000 11927
rect 0 11647 16000 11691
rect 0 11281 16000 11347
rect 0 10625 16000 11221
rect 0 10329 215 10565
rect 451 10329 537 10565
rect 773 10329 859 10565
rect 1095 10329 1181 10565
rect 1417 10329 1503 10565
rect 1739 10329 1825 10565
rect 2061 10329 2147 10565
rect 2383 10329 2469 10565
rect 2705 10329 2791 10565
rect 3027 10329 3113 10565
rect 3349 10329 3435 10565
rect 3671 10329 3757 10565
rect 3993 10329 4079 10565
rect 4315 10329 4401 10565
rect 4637 10329 4723 10565
rect 4959 10329 5045 10565
rect 5281 10329 5367 10565
rect 5603 10329 5689 10565
rect 5925 10329 6011 10565
rect 6247 10329 6332 10565
rect 6568 10329 6653 10565
rect 6889 10329 6974 10565
rect 7210 10329 7295 10565
rect 7531 10329 7616 10565
rect 7852 10329 7937 10565
rect 8173 10329 8258 10565
rect 8494 10329 8579 10565
rect 8815 10329 8900 10565
rect 9136 10329 9221 10565
rect 9457 10329 9542 10565
rect 9778 10329 9863 10565
rect 10099 10329 10184 10565
rect 10420 10329 10505 10565
rect 10741 10329 10826 10565
rect 11062 10329 11147 10565
rect 11383 10329 11468 10565
rect 11704 10329 11789 10565
rect 12025 10329 12110 10565
rect 12346 10329 12431 10565
rect 12667 10329 12752 10565
rect 12988 10329 13073 10565
rect 13309 10329 13394 10565
rect 13630 10329 13715 10565
rect 13951 10329 14036 10565
rect 14272 10329 14357 10565
rect 14593 10329 14678 10565
rect 14914 10329 14999 10565
rect 15235 10329 15320 10565
rect 15556 10329 16000 10565
rect 0 9673 16000 10269
rect 0 9547 16000 9613
rect 0 9244 16000 9247
rect 0 9203 397 9244
rect 0 8967 216 9203
rect 461 9180 479 9244
rect 543 9203 561 9244
rect 625 9203 643 9244
rect 707 9203 725 9244
rect 789 9180 807 9244
rect 871 9203 889 9244
rect 953 9203 971 9244
rect 1035 9203 1053 9244
rect 1117 9180 1135 9244
rect 1199 9203 1217 9244
rect 1281 9203 1299 9244
rect 1363 9203 1381 9244
rect 1445 9180 1463 9244
rect 1527 9203 1545 9244
rect 1609 9203 1627 9244
rect 1691 9203 1709 9244
rect 1773 9180 1791 9244
rect 1855 9203 1873 9244
rect 1937 9203 1955 9244
rect 2019 9203 2037 9244
rect 2101 9180 2119 9244
rect 2183 9203 2201 9244
rect 2265 9203 2282 9244
rect 2346 9203 2363 9244
rect 2427 9203 2553 9244
rect 2617 9203 2635 9244
rect 2699 9203 2717 9244
rect 2427 9180 2470 9203
rect 2706 9180 2717 9203
rect 2781 9203 2799 9244
rect 2863 9203 2881 9244
rect 2945 9203 2963 9244
rect 3027 9203 3045 9244
rect 2781 9180 2792 9203
rect 3028 9180 3045 9203
rect 3109 9203 3127 9244
rect 3191 9203 3209 9244
rect 3273 9203 3290 9244
rect 3109 9180 3114 9203
rect 3354 9180 3371 9244
rect 3435 9203 3452 9244
rect 3516 9203 3533 9244
rect 3597 9203 3614 9244
rect 3435 9180 3436 9203
rect 3678 9180 3695 9244
rect 3759 9203 3776 9244
rect 3840 9203 3857 9244
rect 3921 9203 3938 9244
rect 4002 9180 4019 9244
rect 4083 9203 4100 9244
rect 4164 9203 4181 9244
rect 4245 9203 4262 9244
rect 4326 9180 4343 9244
rect 4407 9203 4424 9244
rect 4488 9203 4505 9244
rect 4569 9203 4695 9244
rect 4759 9203 4777 9244
rect 4841 9203 4859 9244
rect 4923 9203 4941 9244
rect 4638 9180 4695 9203
rect 5005 9180 5023 9244
rect 5087 9203 5105 9244
rect 5169 9203 5187 9244
rect 5251 9203 5269 9244
rect 5333 9180 5351 9244
rect 5415 9203 5433 9244
rect 5497 9203 5515 9244
rect 5579 9203 5597 9244
rect 5661 9180 5679 9244
rect 5743 9203 5760 9244
rect 5824 9203 5841 9244
rect 5905 9203 5922 9244
rect 5986 9180 6003 9244
rect 6067 9203 6084 9244
rect 6148 9203 6165 9244
rect 6229 9203 6246 9244
rect 6310 9180 6327 9244
rect 6391 9203 6408 9244
rect 6472 9203 6489 9244
rect 6553 9203 6570 9244
rect 6569 9180 6570 9203
rect 6634 9180 6651 9244
rect 6715 9203 6732 9244
rect 6796 9203 6813 9244
rect 6877 9203 6894 9244
rect 6890 9180 6894 9203
rect 6958 9180 6975 9244
rect 7039 9203 7056 9244
rect 7120 9203 7137 9244
rect 7201 9203 7218 9244
rect 7211 9180 7218 9203
rect 7282 9203 7299 9244
rect 7363 9203 7380 9244
rect 7444 9203 7461 9244
rect 7525 9203 7542 9244
rect 7282 9180 7296 9203
rect 7532 9180 7542 9203
rect 7606 9203 7623 9244
rect 7687 9241 8859 9244
rect 7687 9203 7813 9241
rect 7606 9180 7617 9203
rect 452 9158 538 9180
rect 774 9158 860 9180
rect 1096 9158 1182 9180
rect 1418 9158 1504 9180
rect 1740 9158 1826 9180
rect 2062 9158 2148 9180
rect 2384 9158 2470 9180
rect 2706 9158 2792 9180
rect 3028 9158 3114 9180
rect 3350 9158 3436 9180
rect 3672 9158 3758 9180
rect 3994 9158 4080 9180
rect 4316 9158 4402 9180
rect 4638 9158 4724 9180
rect 4960 9158 5046 9180
rect 5282 9158 5368 9180
rect 5604 9158 5690 9180
rect 5926 9158 6012 9180
rect 6248 9158 6333 9180
rect 6569 9158 6654 9180
rect 6890 9158 6975 9180
rect 7211 9158 7296 9180
rect 7532 9158 7617 9180
rect 7877 9177 7897 9241
rect 7961 9203 7981 9241
rect 8045 9203 8065 9241
rect 8129 9203 8149 9241
rect 8213 9203 8859 9241
rect 8923 9203 8940 9244
rect 9004 9203 9021 9244
rect 9085 9203 9102 9244
rect 8213 9177 8259 9203
rect 461 9094 479 9158
rect 789 9094 807 9158
rect 1117 9094 1135 9158
rect 1445 9094 1463 9158
rect 1773 9094 1791 9158
rect 2101 9094 2119 9158
rect 2427 9094 2470 9158
rect 2706 9094 2717 9158
rect 2781 9094 2792 9158
rect 3028 9094 3045 9158
rect 3109 9094 3114 9158
rect 3354 9094 3371 9158
rect 3435 9094 3436 9158
rect 3678 9094 3695 9158
rect 4002 9094 4019 9158
rect 4326 9094 4343 9158
rect 4638 9094 4695 9158
rect 5005 9094 5023 9158
rect 5333 9094 5351 9158
rect 5661 9094 5679 9158
rect 5986 9094 6003 9158
rect 6310 9094 6327 9158
rect 6569 9094 6570 9158
rect 6634 9094 6651 9158
rect 6890 9094 6894 9158
rect 6958 9094 6975 9158
rect 7211 9094 7218 9158
rect 7282 9094 7296 9158
rect 7532 9094 7542 9158
rect 7606 9094 7617 9158
rect 7853 9156 7938 9177
rect 8174 9156 8259 9177
rect 452 9072 538 9094
rect 774 9072 860 9094
rect 1096 9072 1182 9094
rect 1418 9072 1504 9094
rect 1740 9072 1826 9094
rect 2062 9072 2148 9094
rect 2384 9072 2470 9094
rect 2706 9072 2792 9094
rect 3028 9072 3114 9094
rect 3350 9072 3436 9094
rect 3672 9072 3758 9094
rect 3994 9072 4080 9094
rect 4316 9072 4402 9094
rect 4638 9072 4724 9094
rect 4960 9072 5046 9094
rect 5282 9072 5368 9094
rect 5604 9072 5690 9094
rect 5926 9072 6012 9094
rect 6248 9072 6333 9094
rect 6569 9072 6654 9094
rect 6890 9072 6975 9094
rect 7211 9072 7296 9094
rect 7532 9072 7617 9094
rect 7877 9092 7897 9156
rect 8213 9092 8259 9156
rect 461 9008 479 9072
rect 789 9008 807 9072
rect 1117 9008 1135 9072
rect 1445 9008 1463 9072
rect 1773 9008 1791 9072
rect 2101 9008 2119 9072
rect 2427 9008 2470 9072
rect 2706 9008 2717 9072
rect 2781 9008 2792 9072
rect 3028 9008 3045 9072
rect 3109 9008 3114 9072
rect 3354 9008 3371 9072
rect 3435 9008 3436 9072
rect 3678 9008 3695 9072
rect 4002 9008 4019 9072
rect 4326 9008 4343 9072
rect 4638 9008 4695 9072
rect 5005 9008 5023 9072
rect 5333 9008 5351 9072
rect 5661 9008 5679 9072
rect 5986 9008 6003 9072
rect 6310 9008 6327 9072
rect 6569 9008 6570 9072
rect 6634 9008 6651 9072
rect 6890 9008 6894 9072
rect 6958 9008 6975 9072
rect 7211 9008 7218 9072
rect 7282 9008 7296 9072
rect 7532 9008 7542 9072
rect 7606 9008 7617 9072
rect 7853 9071 7938 9092
rect 8174 9071 8259 9092
rect 452 8986 538 9008
rect 774 8986 860 9008
rect 1096 8986 1182 9008
rect 1418 8986 1504 9008
rect 1740 8986 1826 9008
rect 2062 8986 2148 9008
rect 2384 8986 2470 9008
rect 2706 8986 2792 9008
rect 3028 8986 3114 9008
rect 3350 8986 3436 9008
rect 3672 8986 3758 9008
rect 3994 8986 4080 9008
rect 4316 8986 4402 9008
rect 4638 8986 4724 9008
rect 4960 8986 5046 9008
rect 5282 8986 5368 9008
rect 5604 8986 5690 9008
rect 5926 8986 6012 9008
rect 6248 8986 6333 9008
rect 6569 8986 6654 9008
rect 6890 8986 6975 9008
rect 7211 8986 7296 9008
rect 7532 8986 7617 9008
rect 7877 9007 7897 9071
rect 8213 9007 8259 9071
rect 7853 8986 7938 9007
rect 8174 8986 8259 9007
rect 0 8922 397 8967
rect 461 8922 479 8986
rect 543 8922 561 8967
rect 625 8922 643 8967
rect 707 8922 725 8967
rect 789 8922 807 8986
rect 871 8922 889 8967
rect 953 8922 971 8967
rect 1035 8922 1053 8967
rect 1117 8922 1135 8986
rect 1199 8922 1217 8967
rect 1281 8922 1299 8967
rect 1363 8922 1381 8967
rect 1445 8922 1463 8986
rect 1527 8922 1545 8967
rect 1609 8922 1627 8967
rect 1691 8922 1709 8967
rect 1773 8922 1791 8986
rect 1855 8922 1873 8967
rect 1937 8922 1955 8967
rect 2019 8922 2037 8967
rect 2101 8922 2119 8986
rect 2427 8967 2470 8986
rect 2706 8967 2717 8986
rect 2183 8922 2201 8967
rect 2265 8922 2282 8967
rect 2346 8922 2363 8967
rect 2427 8922 2553 8967
rect 2617 8922 2635 8967
rect 2699 8922 2717 8967
rect 2781 8967 2792 8986
rect 3028 8967 3045 8986
rect 2781 8922 2799 8967
rect 2863 8922 2881 8967
rect 2945 8922 2963 8967
rect 3027 8922 3045 8967
rect 3109 8967 3114 8986
rect 3109 8922 3127 8967
rect 3191 8922 3209 8967
rect 3273 8922 3290 8967
rect 3354 8922 3371 8986
rect 3435 8967 3436 8986
rect 3435 8922 3452 8967
rect 3516 8922 3533 8967
rect 3597 8922 3614 8967
rect 3678 8922 3695 8986
rect 3759 8922 3776 8967
rect 3840 8922 3857 8967
rect 3921 8922 3938 8967
rect 4002 8922 4019 8986
rect 4083 8922 4100 8967
rect 4164 8922 4181 8967
rect 4245 8922 4262 8967
rect 4326 8922 4343 8986
rect 4638 8967 4695 8986
rect 4407 8922 4424 8967
rect 4488 8922 4505 8967
rect 4569 8922 4695 8967
rect 4759 8922 4777 8967
rect 4841 8922 4859 8967
rect 4923 8922 4941 8967
rect 5005 8922 5023 8986
rect 5087 8922 5105 8967
rect 5169 8922 5187 8967
rect 5251 8922 5269 8967
rect 5333 8922 5351 8986
rect 5415 8922 5433 8967
rect 5497 8922 5515 8967
rect 5579 8922 5597 8967
rect 5661 8922 5679 8986
rect 5743 8922 5760 8967
rect 5824 8922 5841 8967
rect 5905 8922 5922 8967
rect 5986 8922 6003 8986
rect 6067 8922 6084 8967
rect 6148 8922 6165 8967
rect 6229 8922 6246 8967
rect 6310 8922 6327 8986
rect 6569 8967 6570 8986
rect 6391 8922 6408 8967
rect 6472 8922 6489 8967
rect 6553 8922 6570 8967
rect 6634 8922 6651 8986
rect 6890 8967 6894 8986
rect 6715 8922 6732 8967
rect 6796 8922 6813 8967
rect 6877 8922 6894 8967
rect 6958 8922 6975 8986
rect 7211 8967 7218 8986
rect 7039 8922 7056 8967
rect 7120 8922 7137 8967
rect 7201 8922 7218 8967
rect 7282 8967 7296 8986
rect 7532 8967 7542 8986
rect 7282 8922 7299 8967
rect 7363 8922 7380 8967
rect 7444 8922 7461 8967
rect 7525 8922 7542 8967
rect 7606 8967 7617 8986
rect 7606 8922 7623 8967
rect 7687 8922 7813 8967
rect 7877 8922 7897 8986
rect 8213 8967 8259 8986
rect 8495 8967 8580 9203
rect 8816 9180 8859 9203
rect 9166 9180 9183 9244
rect 9247 9203 9264 9244
rect 9328 9203 9345 9244
rect 9409 9203 9426 9244
rect 9490 9180 9507 9244
rect 9571 9203 9588 9244
rect 9652 9203 9669 9244
rect 9733 9203 9750 9244
rect 9814 9180 9831 9244
rect 9895 9203 9912 9244
rect 9976 9203 9993 9244
rect 10057 9203 10073 9244
rect 10137 9180 10153 9244
rect 10217 9203 10233 9244
rect 10297 9203 10313 9244
rect 10377 9203 10393 9244
rect 10457 9180 10473 9244
rect 10537 9203 10553 9244
rect 10617 9203 10633 9244
rect 10697 9203 10713 9244
rect 10777 9180 10793 9244
rect 10857 9203 10873 9244
rect 10937 9203 10953 9244
rect 11017 9203 11033 9244
rect 11097 9180 11113 9244
rect 11177 9203 11193 9244
rect 11257 9203 11273 9244
rect 11337 9203 11353 9244
rect 11417 9180 11433 9244
rect 11497 9203 11513 9244
rect 11577 9203 11593 9244
rect 11657 9203 11673 9244
rect 11737 9180 11753 9244
rect 11817 9203 11833 9244
rect 11897 9203 11913 9244
rect 11977 9203 12165 9244
rect 12229 9203 12246 9244
rect 12310 9203 12327 9244
rect 8816 9158 8901 9180
rect 9137 9158 9222 9180
rect 9458 9158 9543 9180
rect 9779 9158 9864 9180
rect 10100 9158 10185 9180
rect 10421 9158 10506 9180
rect 10742 9158 10827 9180
rect 11063 9158 11148 9180
rect 11384 9158 11469 9180
rect 11705 9158 11790 9180
rect 8816 9094 8859 9158
rect 9166 9094 9183 9158
rect 9490 9094 9507 9158
rect 9814 9094 9831 9158
rect 10137 9094 10153 9158
rect 10457 9094 10473 9158
rect 10777 9094 10793 9158
rect 11097 9094 11113 9158
rect 11417 9094 11433 9158
rect 11737 9094 11753 9158
rect 8816 9072 8901 9094
rect 9137 9072 9222 9094
rect 9458 9072 9543 9094
rect 9779 9072 9864 9094
rect 10100 9072 10185 9094
rect 10421 9072 10506 9094
rect 10742 9072 10827 9094
rect 11063 9072 11148 9094
rect 11384 9072 11469 9094
rect 11705 9072 11790 9094
rect 8816 9008 8859 9072
rect 9166 9008 9183 9072
rect 9490 9008 9507 9072
rect 9814 9008 9831 9072
rect 10137 9008 10153 9072
rect 10457 9008 10473 9072
rect 10777 9008 10793 9072
rect 11097 9008 11113 9072
rect 11417 9008 11433 9072
rect 11737 9008 11753 9072
rect 8816 8986 8901 9008
rect 9137 8986 9222 9008
rect 9458 8986 9543 9008
rect 9779 8986 9864 9008
rect 10100 8986 10185 9008
rect 10421 8986 10506 9008
rect 10742 8986 10827 9008
rect 11063 8986 11148 9008
rect 11384 8986 11469 9008
rect 11705 8986 11790 9008
rect 8816 8967 8859 8986
rect 7961 8922 7981 8967
rect 8045 8922 8065 8967
rect 8129 8922 8149 8967
rect 8213 8922 8859 8967
rect 8923 8922 8940 8967
rect 9004 8922 9021 8967
rect 9085 8922 9102 8967
rect 9166 8922 9183 8986
rect 9247 8922 9264 8967
rect 9328 8922 9345 8967
rect 9409 8922 9426 8967
rect 9490 8922 9507 8986
rect 9571 8922 9588 8967
rect 9652 8922 9669 8967
rect 9733 8922 9750 8967
rect 9814 8922 9831 8986
rect 9895 8922 9912 8967
rect 9976 8922 9993 8967
rect 10057 8922 10073 8967
rect 10137 8922 10153 8986
rect 10217 8922 10233 8967
rect 10297 8922 10313 8967
rect 10377 8922 10393 8967
rect 10457 8922 10473 8986
rect 10537 8922 10553 8967
rect 10617 8922 10633 8967
rect 10697 8922 10713 8967
rect 10777 8922 10793 8986
rect 10857 8922 10873 8967
rect 10937 8922 10953 8967
rect 11017 8922 11033 8967
rect 11097 8922 11113 8986
rect 11177 8922 11193 8967
rect 11257 8922 11273 8967
rect 11337 8922 11353 8967
rect 11417 8922 11433 8986
rect 11497 8922 11513 8967
rect 11577 8922 11593 8967
rect 11657 8922 11673 8967
rect 11737 8922 11753 8986
rect 12026 8967 12111 9203
rect 12391 9180 12408 9244
rect 12472 9203 12489 9244
rect 12553 9203 12570 9244
rect 12634 9203 12651 9244
rect 12715 9180 12732 9244
rect 12796 9203 12813 9244
rect 12877 9203 12894 9244
rect 12958 9203 12975 9244
rect 13039 9180 13056 9244
rect 13120 9203 13137 9244
rect 13201 9203 13218 9244
rect 13282 9203 13299 9244
rect 13363 9180 13380 9244
rect 13444 9203 13461 9244
rect 13525 9203 13542 9244
rect 13606 9203 13623 9244
rect 13687 9180 13704 9244
rect 13768 9203 13785 9244
rect 13849 9203 13866 9244
rect 13930 9203 13947 9244
rect 14011 9180 14028 9244
rect 14092 9203 14109 9244
rect 14173 9203 14190 9244
rect 14254 9203 14271 9244
rect 14335 9180 14352 9244
rect 14416 9203 14433 9244
rect 14497 9203 14513 9244
rect 14577 9203 14593 9244
rect 14657 9180 14673 9244
rect 14737 9203 14753 9244
rect 14817 9203 14833 9244
rect 14897 9203 14913 9244
rect 14977 9180 14993 9244
rect 15057 9203 15073 9244
rect 15137 9203 15153 9244
rect 15217 9203 15233 9244
rect 15297 9180 15313 9244
rect 15377 9203 15393 9244
rect 15457 9203 15473 9244
rect 15537 9203 15553 9244
rect 15617 9180 16000 9244
rect 12347 9158 12432 9180
rect 12668 9158 12753 9180
rect 12989 9158 13074 9180
rect 13310 9158 13395 9180
rect 13631 9158 13716 9180
rect 13952 9158 14037 9180
rect 14273 9158 14358 9180
rect 14594 9158 14679 9180
rect 14915 9158 15000 9180
rect 15236 9158 15321 9180
rect 15557 9158 16000 9180
rect 12391 9094 12408 9158
rect 12715 9094 12732 9158
rect 13039 9094 13056 9158
rect 13363 9094 13380 9158
rect 13687 9094 13704 9158
rect 14011 9094 14028 9158
rect 14335 9094 14352 9158
rect 14657 9094 14673 9158
rect 14977 9094 14993 9158
rect 15297 9094 15313 9158
rect 15617 9094 16000 9158
rect 12347 9072 12432 9094
rect 12668 9072 12753 9094
rect 12989 9072 13074 9094
rect 13310 9072 13395 9094
rect 13631 9072 13716 9094
rect 13952 9072 14037 9094
rect 14273 9072 14358 9094
rect 14594 9072 14679 9094
rect 14915 9072 15000 9094
rect 15236 9072 15321 9094
rect 15557 9072 16000 9094
rect 12391 9008 12408 9072
rect 12715 9008 12732 9072
rect 13039 9008 13056 9072
rect 13363 9008 13380 9072
rect 13687 9008 13704 9072
rect 14011 9008 14028 9072
rect 14335 9008 14352 9072
rect 14657 9008 14673 9072
rect 14977 9008 14993 9072
rect 15297 9008 15313 9072
rect 15617 9008 16000 9072
rect 12347 8986 12432 9008
rect 12668 8986 12753 9008
rect 12989 8986 13074 9008
rect 13310 8986 13395 9008
rect 13631 8986 13716 9008
rect 13952 8986 14037 9008
rect 14273 8986 14358 9008
rect 14594 8986 14679 9008
rect 14915 8986 15000 9008
rect 15236 8986 15321 9008
rect 15557 8986 16000 9008
rect 11817 8922 11833 8967
rect 11897 8922 11913 8967
rect 11977 8922 12165 8967
rect 12229 8922 12246 8967
rect 12310 8922 12327 8967
rect 12391 8922 12408 8986
rect 12472 8922 12489 8967
rect 12553 8922 12570 8967
rect 12634 8922 12651 8967
rect 12715 8922 12732 8986
rect 12796 8922 12813 8967
rect 12877 8922 12894 8967
rect 12958 8922 12975 8967
rect 13039 8922 13056 8986
rect 13120 8922 13137 8967
rect 13201 8922 13218 8967
rect 13282 8922 13299 8967
rect 13363 8922 13380 8986
rect 13444 8922 13461 8967
rect 13525 8922 13542 8967
rect 13606 8922 13623 8967
rect 13687 8922 13704 8986
rect 13768 8922 13785 8967
rect 13849 8922 13866 8967
rect 13930 8922 13947 8967
rect 14011 8922 14028 8986
rect 14092 8922 14109 8967
rect 14173 8922 14190 8967
rect 14254 8922 14271 8967
rect 14335 8922 14352 8986
rect 14416 8922 14433 8967
rect 14497 8922 14513 8967
rect 14577 8922 14593 8967
rect 14657 8922 14673 8986
rect 14737 8922 14753 8967
rect 14817 8922 14833 8967
rect 14897 8922 14913 8967
rect 14977 8922 14993 8986
rect 15057 8922 15073 8967
rect 15137 8922 15153 8967
rect 15217 8922 15233 8967
rect 15297 8922 15313 8986
rect 15377 8922 15393 8967
rect 15457 8922 15473 8967
rect 15537 8922 15553 8967
rect 15617 8922 16000 8986
rect 0 8901 16000 8922
rect 0 8900 7813 8901
rect 0 8836 397 8900
rect 461 8836 479 8900
rect 543 8836 561 8900
rect 625 8836 643 8900
rect 707 8836 725 8900
rect 789 8836 807 8900
rect 871 8836 889 8900
rect 953 8836 971 8900
rect 1035 8836 1053 8900
rect 1117 8836 1135 8900
rect 1199 8836 1217 8900
rect 1281 8836 1299 8900
rect 1363 8836 1381 8900
rect 1445 8836 1463 8900
rect 1527 8836 1545 8900
rect 1609 8836 1627 8900
rect 1691 8836 1709 8900
rect 1773 8836 1791 8900
rect 1855 8836 1873 8900
rect 1937 8836 1955 8900
rect 2019 8836 2037 8900
rect 2101 8836 2119 8900
rect 2183 8836 2201 8900
rect 2265 8836 2282 8900
rect 2346 8836 2363 8900
rect 2427 8836 2553 8900
rect 2617 8836 2635 8900
rect 2699 8836 2717 8900
rect 2781 8836 2799 8900
rect 2863 8836 2881 8900
rect 2945 8836 2963 8900
rect 3027 8836 3045 8900
rect 3109 8836 3127 8900
rect 3191 8836 3209 8900
rect 3273 8836 3290 8900
rect 3354 8836 3371 8900
rect 3435 8836 3452 8900
rect 3516 8836 3533 8900
rect 3597 8836 3614 8900
rect 3678 8836 3695 8900
rect 3759 8836 3776 8900
rect 3840 8836 3857 8900
rect 3921 8836 3938 8900
rect 4002 8836 4019 8900
rect 4083 8836 4100 8900
rect 4164 8836 4181 8900
rect 4245 8836 4262 8900
rect 4326 8836 4343 8900
rect 4407 8836 4424 8900
rect 4488 8836 4505 8900
rect 4569 8836 4695 8900
rect 4759 8836 4777 8900
rect 4841 8836 4859 8900
rect 4923 8836 4941 8900
rect 5005 8836 5023 8900
rect 5087 8836 5105 8900
rect 5169 8836 5187 8900
rect 5251 8836 5269 8900
rect 5333 8836 5351 8900
rect 5415 8836 5433 8900
rect 5497 8836 5515 8900
rect 5579 8836 5597 8900
rect 5661 8836 5679 8900
rect 5743 8836 5760 8900
rect 5824 8836 5841 8900
rect 5905 8836 5922 8900
rect 5986 8836 6003 8900
rect 6067 8836 6084 8900
rect 6148 8836 6165 8900
rect 6229 8836 6246 8900
rect 6310 8836 6327 8900
rect 6391 8836 6408 8900
rect 6472 8836 6489 8900
rect 6553 8836 6570 8900
rect 6634 8836 6651 8900
rect 6715 8836 6732 8900
rect 6796 8836 6813 8900
rect 6877 8836 6894 8900
rect 6958 8836 6975 8900
rect 7039 8836 7056 8900
rect 7120 8836 7137 8900
rect 7201 8836 7218 8900
rect 7282 8836 7299 8900
rect 7363 8836 7380 8900
rect 7444 8836 7461 8900
rect 7525 8836 7542 8900
rect 7606 8836 7623 8900
rect 7687 8837 7813 8900
rect 7877 8837 7897 8901
rect 7961 8837 7981 8901
rect 8045 8837 8065 8901
rect 8129 8837 8149 8901
rect 8213 8900 16000 8901
rect 8213 8837 8859 8900
rect 7687 8836 8859 8837
rect 8923 8836 8940 8900
rect 9004 8836 9021 8900
rect 9085 8836 9102 8900
rect 9166 8836 9183 8900
rect 9247 8836 9264 8900
rect 9328 8836 9345 8900
rect 9409 8836 9426 8900
rect 9490 8836 9507 8900
rect 9571 8836 9588 8900
rect 9652 8836 9669 8900
rect 9733 8836 9750 8900
rect 9814 8836 9831 8900
rect 9895 8836 9912 8900
rect 9976 8836 9993 8900
rect 10057 8836 10073 8900
rect 10137 8836 10153 8900
rect 10217 8836 10233 8900
rect 10297 8836 10313 8900
rect 10377 8836 10393 8900
rect 10457 8836 10473 8900
rect 10537 8836 10553 8900
rect 10617 8836 10633 8900
rect 10697 8836 10713 8900
rect 10777 8836 10793 8900
rect 10857 8836 10873 8900
rect 10937 8836 10953 8900
rect 11017 8836 11033 8900
rect 11097 8836 11113 8900
rect 11177 8836 11193 8900
rect 11257 8836 11273 8900
rect 11337 8836 11353 8900
rect 11417 8836 11433 8900
rect 11497 8836 11513 8900
rect 11577 8836 11593 8900
rect 11657 8836 11673 8900
rect 11737 8836 11753 8900
rect 11817 8836 11833 8900
rect 11897 8836 11913 8900
rect 11977 8836 12165 8900
rect 12229 8836 12246 8900
rect 12310 8836 12327 8900
rect 12391 8836 12408 8900
rect 12472 8836 12489 8900
rect 12553 8836 12570 8900
rect 12634 8836 12651 8900
rect 12715 8836 12732 8900
rect 12796 8836 12813 8900
rect 12877 8836 12894 8900
rect 12958 8836 12975 8900
rect 13039 8836 13056 8900
rect 13120 8836 13137 8900
rect 13201 8836 13218 8900
rect 13282 8836 13299 8900
rect 13363 8836 13380 8900
rect 13444 8836 13461 8900
rect 13525 8836 13542 8900
rect 13606 8836 13623 8900
rect 13687 8836 13704 8900
rect 13768 8836 13785 8900
rect 13849 8836 13866 8900
rect 13930 8836 13947 8900
rect 14011 8836 14028 8900
rect 14092 8836 14109 8900
rect 14173 8836 14190 8900
rect 14254 8836 14271 8900
rect 14335 8836 14352 8900
rect 14416 8836 14433 8900
rect 14497 8836 14513 8900
rect 14577 8836 14593 8900
rect 14657 8836 14673 8900
rect 14737 8836 14753 8900
rect 14817 8836 14833 8900
rect 14897 8836 14913 8900
rect 14977 8836 14993 8900
rect 15057 8836 15073 8900
rect 15137 8836 15153 8900
rect 15217 8836 15233 8900
rect 15297 8836 15313 8900
rect 15377 8836 15393 8900
rect 15457 8836 15473 8900
rect 15537 8836 15553 8900
rect 15617 8836 16000 8900
rect 0 8816 16000 8836
rect 0 8814 7813 8816
rect 0 8750 397 8814
rect 461 8750 479 8814
rect 543 8750 561 8814
rect 625 8750 643 8814
rect 707 8750 725 8814
rect 789 8750 807 8814
rect 871 8750 889 8814
rect 953 8750 971 8814
rect 1035 8750 1053 8814
rect 1117 8750 1135 8814
rect 1199 8750 1217 8814
rect 1281 8750 1299 8814
rect 1363 8750 1381 8814
rect 1445 8750 1463 8814
rect 1527 8750 1545 8814
rect 1609 8750 1627 8814
rect 1691 8750 1709 8814
rect 1773 8750 1791 8814
rect 1855 8750 1873 8814
rect 1937 8750 1955 8814
rect 2019 8750 2037 8814
rect 2101 8750 2119 8814
rect 2183 8750 2201 8814
rect 2265 8750 2282 8814
rect 2346 8750 2363 8814
rect 2427 8750 2553 8814
rect 2617 8750 2635 8814
rect 2699 8750 2717 8814
rect 2781 8750 2799 8814
rect 2863 8750 2881 8814
rect 2945 8750 2963 8814
rect 3027 8750 3045 8814
rect 3109 8750 3127 8814
rect 3191 8750 3209 8814
rect 3273 8750 3290 8814
rect 3354 8750 3371 8814
rect 3435 8750 3452 8814
rect 3516 8750 3533 8814
rect 3597 8750 3614 8814
rect 3678 8750 3695 8814
rect 3759 8750 3776 8814
rect 3840 8750 3857 8814
rect 3921 8750 3938 8814
rect 4002 8750 4019 8814
rect 4083 8750 4100 8814
rect 4164 8750 4181 8814
rect 4245 8750 4262 8814
rect 4326 8750 4343 8814
rect 4407 8750 4424 8814
rect 4488 8750 4505 8814
rect 4569 8750 4695 8814
rect 4759 8750 4777 8814
rect 4841 8750 4859 8814
rect 4923 8750 4941 8814
rect 5005 8750 5023 8814
rect 5087 8750 5105 8814
rect 5169 8750 5187 8814
rect 5251 8750 5269 8814
rect 5333 8750 5351 8814
rect 5415 8750 5433 8814
rect 5497 8750 5515 8814
rect 5579 8750 5597 8814
rect 5661 8750 5679 8814
rect 5743 8750 5760 8814
rect 5824 8750 5841 8814
rect 5905 8750 5922 8814
rect 5986 8750 6003 8814
rect 6067 8750 6084 8814
rect 6148 8750 6165 8814
rect 6229 8750 6246 8814
rect 6310 8750 6327 8814
rect 6391 8750 6408 8814
rect 6472 8750 6489 8814
rect 6553 8750 6570 8814
rect 6634 8750 6651 8814
rect 6715 8750 6732 8814
rect 6796 8750 6813 8814
rect 6877 8750 6894 8814
rect 6958 8750 6975 8814
rect 7039 8750 7056 8814
rect 7120 8750 7137 8814
rect 7201 8750 7218 8814
rect 7282 8750 7299 8814
rect 7363 8750 7380 8814
rect 7444 8750 7461 8814
rect 7525 8750 7542 8814
rect 7606 8750 7623 8814
rect 7687 8752 7813 8814
rect 7877 8752 7897 8816
rect 7961 8752 7981 8816
rect 8045 8752 8065 8816
rect 8129 8752 8149 8816
rect 8213 8814 16000 8816
rect 8213 8752 8859 8814
rect 7687 8750 8859 8752
rect 8923 8750 8940 8814
rect 9004 8750 9021 8814
rect 9085 8750 9102 8814
rect 9166 8750 9183 8814
rect 9247 8750 9264 8814
rect 9328 8750 9345 8814
rect 9409 8750 9426 8814
rect 9490 8750 9507 8814
rect 9571 8750 9588 8814
rect 9652 8750 9669 8814
rect 9733 8750 9750 8814
rect 9814 8750 9831 8814
rect 9895 8750 9912 8814
rect 9976 8750 9993 8814
rect 10057 8750 10073 8814
rect 10137 8750 10153 8814
rect 10217 8750 10233 8814
rect 10297 8750 10313 8814
rect 10377 8750 10393 8814
rect 10457 8750 10473 8814
rect 10537 8750 10553 8814
rect 10617 8750 10633 8814
rect 10697 8750 10713 8814
rect 10777 8750 10793 8814
rect 10857 8750 10873 8814
rect 10937 8750 10953 8814
rect 11017 8750 11033 8814
rect 11097 8750 11113 8814
rect 11177 8750 11193 8814
rect 11257 8750 11273 8814
rect 11337 8750 11353 8814
rect 11417 8750 11433 8814
rect 11497 8750 11513 8814
rect 11577 8750 11593 8814
rect 11657 8750 11673 8814
rect 11737 8750 11753 8814
rect 11817 8750 11833 8814
rect 11897 8750 11913 8814
rect 11977 8750 12165 8814
rect 12229 8750 12246 8814
rect 12310 8750 12327 8814
rect 12391 8750 12408 8814
rect 12472 8750 12489 8814
rect 12553 8750 12570 8814
rect 12634 8750 12651 8814
rect 12715 8750 12732 8814
rect 12796 8750 12813 8814
rect 12877 8750 12894 8814
rect 12958 8750 12975 8814
rect 13039 8750 13056 8814
rect 13120 8750 13137 8814
rect 13201 8750 13218 8814
rect 13282 8750 13299 8814
rect 13363 8750 13380 8814
rect 13444 8750 13461 8814
rect 13525 8750 13542 8814
rect 13606 8750 13623 8814
rect 13687 8750 13704 8814
rect 13768 8750 13785 8814
rect 13849 8750 13866 8814
rect 13930 8750 13947 8814
rect 14011 8750 14028 8814
rect 14092 8750 14109 8814
rect 14173 8750 14190 8814
rect 14254 8750 14271 8814
rect 14335 8750 14352 8814
rect 14416 8750 14433 8814
rect 14497 8750 14513 8814
rect 14577 8750 14593 8814
rect 14657 8750 14673 8814
rect 14737 8750 14753 8814
rect 14817 8750 14833 8814
rect 14897 8750 14913 8814
rect 14977 8750 14993 8814
rect 15057 8750 15073 8814
rect 15137 8750 15153 8814
rect 15217 8750 15233 8814
rect 15297 8750 15313 8814
rect 15377 8750 15393 8814
rect 15457 8750 15473 8814
rect 15537 8750 15553 8814
rect 15617 8750 16000 8814
rect 0 8731 16000 8750
rect 0 8728 7813 8731
rect 0 8664 397 8728
rect 461 8664 479 8728
rect 543 8664 561 8728
rect 625 8664 643 8728
rect 707 8664 725 8728
rect 789 8664 807 8728
rect 871 8664 889 8728
rect 953 8664 971 8728
rect 1035 8664 1053 8728
rect 1117 8664 1135 8728
rect 1199 8664 1217 8728
rect 1281 8664 1299 8728
rect 1363 8664 1381 8728
rect 1445 8664 1463 8728
rect 1527 8664 1545 8728
rect 1609 8664 1627 8728
rect 1691 8664 1709 8728
rect 1773 8664 1791 8728
rect 1855 8664 1873 8728
rect 1937 8664 1955 8728
rect 2019 8664 2037 8728
rect 2101 8664 2119 8728
rect 2183 8664 2201 8728
rect 2265 8664 2282 8728
rect 2346 8664 2363 8728
rect 2427 8664 2553 8728
rect 2617 8664 2635 8728
rect 2699 8664 2717 8728
rect 2781 8664 2799 8728
rect 2863 8664 2881 8728
rect 2945 8664 2963 8728
rect 3027 8664 3045 8728
rect 3109 8664 3127 8728
rect 3191 8664 3209 8728
rect 3273 8664 3290 8728
rect 3354 8664 3371 8728
rect 3435 8664 3452 8728
rect 3516 8664 3533 8728
rect 3597 8664 3614 8728
rect 3678 8664 3695 8728
rect 3759 8664 3776 8728
rect 3840 8664 3857 8728
rect 3921 8664 3938 8728
rect 4002 8664 4019 8728
rect 4083 8664 4100 8728
rect 4164 8664 4181 8728
rect 4245 8664 4262 8728
rect 4326 8664 4343 8728
rect 4407 8664 4424 8728
rect 4488 8664 4505 8728
rect 4569 8664 4695 8728
rect 4759 8664 4777 8728
rect 4841 8664 4859 8728
rect 4923 8664 4941 8728
rect 5005 8664 5023 8728
rect 5087 8664 5105 8728
rect 5169 8664 5187 8728
rect 5251 8664 5269 8728
rect 5333 8664 5351 8728
rect 5415 8664 5433 8728
rect 5497 8664 5515 8728
rect 5579 8664 5597 8728
rect 5661 8664 5679 8728
rect 5743 8664 5760 8728
rect 5824 8664 5841 8728
rect 5905 8664 5922 8728
rect 5986 8664 6003 8728
rect 6067 8664 6084 8728
rect 6148 8664 6165 8728
rect 6229 8664 6246 8728
rect 6310 8664 6327 8728
rect 6391 8664 6408 8728
rect 6472 8664 6489 8728
rect 6553 8664 6570 8728
rect 6634 8664 6651 8728
rect 6715 8664 6732 8728
rect 6796 8664 6813 8728
rect 6877 8664 6894 8728
rect 6958 8664 6975 8728
rect 7039 8664 7056 8728
rect 7120 8664 7137 8728
rect 7201 8664 7218 8728
rect 7282 8664 7299 8728
rect 7363 8664 7380 8728
rect 7444 8664 7461 8728
rect 7525 8664 7542 8728
rect 7606 8664 7623 8728
rect 7687 8667 7813 8728
rect 7877 8667 7897 8731
rect 7961 8667 7981 8731
rect 8045 8667 8065 8731
rect 8129 8667 8149 8731
rect 8213 8728 16000 8731
rect 8213 8667 8859 8728
rect 7687 8664 8859 8667
rect 8923 8664 8940 8728
rect 9004 8664 9021 8728
rect 9085 8664 9102 8728
rect 9166 8664 9183 8728
rect 9247 8664 9264 8728
rect 9328 8664 9345 8728
rect 9409 8664 9426 8728
rect 9490 8664 9507 8728
rect 9571 8664 9588 8728
rect 9652 8664 9669 8728
rect 9733 8664 9750 8728
rect 9814 8664 9831 8728
rect 9895 8664 9912 8728
rect 9976 8664 9993 8728
rect 10057 8664 10073 8728
rect 10137 8664 10153 8728
rect 10217 8664 10233 8728
rect 10297 8664 10313 8728
rect 10377 8664 10393 8728
rect 10457 8664 10473 8728
rect 10537 8664 10553 8728
rect 10617 8664 10633 8728
rect 10697 8664 10713 8728
rect 10777 8664 10793 8728
rect 10857 8664 10873 8728
rect 10937 8664 10953 8728
rect 11017 8664 11033 8728
rect 11097 8664 11113 8728
rect 11177 8664 11193 8728
rect 11257 8664 11273 8728
rect 11337 8664 11353 8728
rect 11417 8664 11433 8728
rect 11497 8664 11513 8728
rect 11577 8664 11593 8728
rect 11657 8664 11673 8728
rect 11737 8664 11753 8728
rect 11817 8664 11833 8728
rect 11897 8664 11913 8728
rect 11977 8664 12165 8728
rect 12229 8664 12246 8728
rect 12310 8664 12327 8728
rect 12391 8664 12408 8728
rect 12472 8664 12489 8728
rect 12553 8664 12570 8728
rect 12634 8664 12651 8728
rect 12715 8664 12732 8728
rect 12796 8664 12813 8728
rect 12877 8664 12894 8728
rect 12958 8664 12975 8728
rect 13039 8664 13056 8728
rect 13120 8664 13137 8728
rect 13201 8664 13218 8728
rect 13282 8664 13299 8728
rect 13363 8664 13380 8728
rect 13444 8664 13461 8728
rect 13525 8664 13542 8728
rect 13606 8664 13623 8728
rect 13687 8664 13704 8728
rect 13768 8664 13785 8728
rect 13849 8664 13866 8728
rect 13930 8664 13947 8728
rect 14011 8664 14028 8728
rect 14092 8664 14109 8728
rect 14173 8664 14190 8728
rect 14254 8664 14271 8728
rect 14335 8664 14352 8728
rect 14416 8664 14433 8728
rect 14497 8664 14513 8728
rect 14577 8664 14593 8728
rect 14657 8664 14673 8728
rect 14737 8664 14753 8728
rect 14817 8664 14833 8728
rect 14897 8664 14913 8728
rect 14977 8664 14993 8728
rect 15057 8664 15073 8728
rect 15137 8664 15153 8728
rect 15217 8664 15233 8728
rect 15297 8664 15313 8728
rect 15377 8664 15393 8728
rect 15457 8664 15473 8728
rect 15537 8664 15553 8728
rect 15617 8664 16000 8728
rect 0 8645 16000 8664
rect 0 8642 7813 8645
rect 0 8597 397 8642
rect 0 8361 216 8597
rect 461 8578 479 8642
rect 543 8597 561 8642
rect 625 8597 643 8642
rect 707 8597 725 8642
rect 789 8578 807 8642
rect 871 8597 889 8642
rect 953 8597 971 8642
rect 1035 8597 1053 8642
rect 1117 8578 1135 8642
rect 1199 8597 1217 8642
rect 1281 8597 1299 8642
rect 1363 8597 1381 8642
rect 1445 8578 1463 8642
rect 1527 8597 1545 8642
rect 1609 8597 1627 8642
rect 1691 8597 1709 8642
rect 1773 8578 1791 8642
rect 1855 8597 1873 8642
rect 1937 8597 1955 8642
rect 2019 8597 2037 8642
rect 2101 8578 2119 8642
rect 2183 8597 2201 8642
rect 2265 8597 2282 8642
rect 2346 8597 2363 8642
rect 2427 8597 2553 8642
rect 2617 8597 2635 8642
rect 2699 8597 2717 8642
rect 2427 8578 2470 8597
rect 2706 8578 2717 8597
rect 2781 8597 2799 8642
rect 2863 8597 2881 8642
rect 2945 8597 2963 8642
rect 3027 8597 3045 8642
rect 2781 8578 2792 8597
rect 3028 8578 3045 8597
rect 3109 8597 3127 8642
rect 3191 8597 3209 8642
rect 3273 8597 3290 8642
rect 3109 8578 3114 8597
rect 3354 8578 3371 8642
rect 3435 8597 3452 8642
rect 3516 8597 3533 8642
rect 3597 8597 3614 8642
rect 3435 8578 3436 8597
rect 3678 8578 3695 8642
rect 3759 8597 3776 8642
rect 3840 8597 3857 8642
rect 3921 8597 3938 8642
rect 4002 8578 4019 8642
rect 4083 8597 4100 8642
rect 4164 8597 4181 8642
rect 4245 8597 4262 8642
rect 4326 8578 4343 8642
rect 4407 8597 4424 8642
rect 4488 8597 4505 8642
rect 4569 8597 4695 8642
rect 4759 8597 4777 8642
rect 4841 8597 4859 8642
rect 4923 8597 4941 8642
rect 4638 8578 4695 8597
rect 5005 8578 5023 8642
rect 5087 8597 5105 8642
rect 5169 8597 5187 8642
rect 5251 8597 5269 8642
rect 5333 8578 5351 8642
rect 5415 8597 5433 8642
rect 5497 8597 5515 8642
rect 5579 8597 5597 8642
rect 5661 8578 5679 8642
rect 5743 8597 5760 8642
rect 5824 8597 5841 8642
rect 5905 8597 5922 8642
rect 5986 8578 6003 8642
rect 6067 8597 6084 8642
rect 6148 8597 6165 8642
rect 6229 8597 6246 8642
rect 6310 8578 6327 8642
rect 6391 8597 6408 8642
rect 6472 8597 6489 8642
rect 6553 8597 6570 8642
rect 6569 8578 6570 8597
rect 6634 8578 6651 8642
rect 6715 8597 6732 8642
rect 6796 8597 6813 8642
rect 6877 8597 6894 8642
rect 6890 8578 6894 8597
rect 6958 8578 6975 8642
rect 7039 8597 7056 8642
rect 7120 8597 7137 8642
rect 7201 8597 7218 8642
rect 7211 8578 7218 8597
rect 7282 8597 7299 8642
rect 7363 8597 7380 8642
rect 7444 8597 7461 8642
rect 7525 8597 7542 8642
rect 7282 8578 7296 8597
rect 7532 8578 7542 8597
rect 7606 8597 7623 8642
rect 7687 8597 7813 8642
rect 7606 8578 7617 8597
rect 7877 8581 7897 8645
rect 7961 8597 7981 8645
rect 8045 8597 8065 8645
rect 8129 8597 8149 8645
rect 8213 8642 16000 8645
rect 8213 8597 8859 8642
rect 8923 8597 8940 8642
rect 9004 8597 9021 8642
rect 9085 8597 9102 8642
rect 8213 8581 8259 8597
rect 452 8556 538 8578
rect 774 8556 860 8578
rect 1096 8556 1182 8578
rect 1418 8556 1504 8578
rect 1740 8556 1826 8578
rect 2062 8556 2148 8578
rect 2384 8556 2470 8578
rect 2706 8556 2792 8578
rect 3028 8556 3114 8578
rect 3350 8556 3436 8578
rect 3672 8556 3758 8578
rect 3994 8556 4080 8578
rect 4316 8556 4402 8578
rect 4638 8556 4724 8578
rect 4960 8556 5046 8578
rect 5282 8556 5368 8578
rect 5604 8556 5690 8578
rect 5926 8556 6012 8578
rect 6248 8556 6333 8578
rect 6569 8556 6654 8578
rect 6890 8556 6975 8578
rect 7211 8556 7296 8578
rect 7532 8556 7617 8578
rect 7853 8559 7938 8581
rect 8174 8559 8259 8581
rect 461 8492 479 8556
rect 789 8492 807 8556
rect 1117 8492 1135 8556
rect 1445 8492 1463 8556
rect 1773 8492 1791 8556
rect 2101 8492 2119 8556
rect 2427 8492 2470 8556
rect 2706 8492 2717 8556
rect 2781 8492 2792 8556
rect 3028 8492 3045 8556
rect 3109 8492 3114 8556
rect 3354 8492 3371 8556
rect 3435 8492 3436 8556
rect 3678 8492 3695 8556
rect 4002 8492 4019 8556
rect 4326 8492 4343 8556
rect 4638 8492 4695 8556
rect 5005 8492 5023 8556
rect 5333 8492 5351 8556
rect 5661 8492 5679 8556
rect 5986 8492 6003 8556
rect 6310 8492 6327 8556
rect 6569 8492 6570 8556
rect 6634 8492 6651 8556
rect 6890 8492 6894 8556
rect 6958 8492 6975 8556
rect 7211 8492 7218 8556
rect 7282 8492 7296 8556
rect 7532 8492 7542 8556
rect 7606 8492 7617 8556
rect 7877 8495 7897 8559
rect 8213 8495 8259 8559
rect 452 8470 538 8492
rect 774 8470 860 8492
rect 1096 8470 1182 8492
rect 1418 8470 1504 8492
rect 1740 8470 1826 8492
rect 2062 8470 2148 8492
rect 2384 8470 2470 8492
rect 2706 8470 2792 8492
rect 3028 8470 3114 8492
rect 3350 8470 3436 8492
rect 3672 8470 3758 8492
rect 3994 8470 4080 8492
rect 4316 8470 4402 8492
rect 4638 8470 4724 8492
rect 4960 8470 5046 8492
rect 5282 8470 5368 8492
rect 5604 8470 5690 8492
rect 5926 8470 6012 8492
rect 6248 8470 6333 8492
rect 6569 8470 6654 8492
rect 6890 8470 6975 8492
rect 7211 8470 7296 8492
rect 7532 8470 7617 8492
rect 7853 8473 7938 8495
rect 8174 8473 8259 8495
rect 461 8406 479 8470
rect 789 8406 807 8470
rect 1117 8406 1135 8470
rect 1445 8406 1463 8470
rect 1773 8406 1791 8470
rect 2101 8406 2119 8470
rect 2427 8406 2470 8470
rect 2706 8406 2717 8470
rect 2781 8406 2792 8470
rect 3028 8406 3045 8470
rect 3109 8406 3114 8470
rect 3354 8406 3371 8470
rect 3435 8406 3436 8470
rect 3678 8406 3695 8470
rect 4002 8406 4019 8470
rect 4326 8406 4343 8470
rect 4638 8406 4695 8470
rect 5005 8406 5023 8470
rect 5333 8406 5351 8470
rect 5661 8406 5679 8470
rect 5986 8406 6003 8470
rect 6310 8406 6327 8470
rect 6569 8406 6570 8470
rect 6634 8406 6651 8470
rect 6890 8406 6894 8470
rect 6958 8406 6975 8470
rect 7211 8406 7218 8470
rect 7282 8406 7296 8470
rect 7532 8406 7542 8470
rect 7606 8406 7617 8470
rect 7877 8409 7897 8473
rect 8213 8409 8259 8473
rect 452 8384 538 8406
rect 774 8384 860 8406
rect 1096 8384 1182 8406
rect 1418 8384 1504 8406
rect 1740 8384 1826 8406
rect 2062 8384 2148 8406
rect 2384 8384 2470 8406
rect 2706 8384 2792 8406
rect 3028 8384 3114 8406
rect 3350 8384 3436 8406
rect 3672 8384 3758 8406
rect 3994 8384 4080 8406
rect 4316 8384 4402 8406
rect 4638 8384 4724 8406
rect 4960 8384 5046 8406
rect 5282 8384 5368 8406
rect 5604 8384 5690 8406
rect 5926 8384 6012 8406
rect 6248 8384 6333 8406
rect 6569 8384 6654 8406
rect 6890 8384 6975 8406
rect 7211 8384 7296 8406
rect 7532 8384 7617 8406
rect 7853 8387 7938 8409
rect 8174 8387 8259 8409
rect 0 8320 397 8361
rect 461 8320 479 8384
rect 543 8320 561 8361
rect 625 8320 643 8361
rect 707 8320 725 8361
rect 789 8320 807 8384
rect 871 8320 889 8361
rect 953 8320 971 8361
rect 1035 8320 1053 8361
rect 1117 8320 1135 8384
rect 1199 8320 1217 8361
rect 1281 8320 1299 8361
rect 1363 8320 1381 8361
rect 1445 8320 1463 8384
rect 1527 8320 1545 8361
rect 1609 8320 1627 8361
rect 1691 8320 1709 8361
rect 1773 8320 1791 8384
rect 1855 8320 1873 8361
rect 1937 8320 1955 8361
rect 2019 8320 2037 8361
rect 2101 8320 2119 8384
rect 2427 8361 2470 8384
rect 2706 8361 2717 8384
rect 2183 8320 2201 8361
rect 2265 8320 2282 8361
rect 2346 8320 2363 8361
rect 2427 8320 2553 8361
rect 2617 8320 2635 8361
rect 2699 8320 2717 8361
rect 2781 8361 2792 8384
rect 3028 8361 3045 8384
rect 2781 8320 2799 8361
rect 2863 8320 2881 8361
rect 2945 8320 2963 8361
rect 3027 8320 3045 8361
rect 3109 8361 3114 8384
rect 3109 8320 3127 8361
rect 3191 8320 3209 8361
rect 3273 8320 3290 8361
rect 3354 8320 3371 8384
rect 3435 8361 3436 8384
rect 3435 8320 3452 8361
rect 3516 8320 3533 8361
rect 3597 8320 3614 8361
rect 3678 8320 3695 8384
rect 3759 8320 3776 8361
rect 3840 8320 3857 8361
rect 3921 8320 3938 8361
rect 4002 8320 4019 8384
rect 4083 8320 4100 8361
rect 4164 8320 4181 8361
rect 4245 8320 4262 8361
rect 4326 8320 4343 8384
rect 4638 8361 4695 8384
rect 4407 8320 4424 8361
rect 4488 8320 4505 8361
rect 4569 8320 4695 8361
rect 4759 8320 4777 8361
rect 4841 8320 4859 8361
rect 4923 8320 4941 8361
rect 5005 8320 5023 8384
rect 5087 8320 5105 8361
rect 5169 8320 5187 8361
rect 5251 8320 5269 8361
rect 5333 8320 5351 8384
rect 5415 8320 5433 8361
rect 5497 8320 5515 8361
rect 5579 8320 5597 8361
rect 5661 8320 5679 8384
rect 5743 8320 5760 8361
rect 5824 8320 5841 8361
rect 5905 8320 5922 8361
rect 5986 8320 6003 8384
rect 6067 8320 6084 8361
rect 6148 8320 6165 8361
rect 6229 8320 6246 8361
rect 6310 8320 6327 8384
rect 6569 8361 6570 8384
rect 6391 8320 6408 8361
rect 6472 8320 6489 8361
rect 6553 8320 6570 8361
rect 6634 8320 6651 8384
rect 6890 8361 6894 8384
rect 6715 8320 6732 8361
rect 6796 8320 6813 8361
rect 6877 8320 6894 8361
rect 6958 8320 6975 8384
rect 7211 8361 7218 8384
rect 7039 8320 7056 8361
rect 7120 8320 7137 8361
rect 7201 8320 7218 8361
rect 7282 8361 7296 8384
rect 7532 8361 7542 8384
rect 7282 8320 7299 8361
rect 7363 8320 7380 8361
rect 7444 8320 7461 8361
rect 7525 8320 7542 8361
rect 7606 8361 7617 8384
rect 7606 8320 7623 8361
rect 7687 8323 7813 8361
rect 7877 8323 7897 8387
rect 8213 8361 8259 8387
rect 8495 8361 8580 8597
rect 8816 8578 8859 8597
rect 9166 8578 9183 8642
rect 9247 8597 9264 8642
rect 9328 8597 9345 8642
rect 9409 8597 9426 8642
rect 9490 8578 9507 8642
rect 9571 8597 9588 8642
rect 9652 8597 9669 8642
rect 9733 8597 9750 8642
rect 9814 8578 9831 8642
rect 9895 8597 9912 8642
rect 9976 8597 9993 8642
rect 10057 8597 10073 8642
rect 10137 8578 10153 8642
rect 10217 8597 10233 8642
rect 10297 8597 10313 8642
rect 10377 8597 10393 8642
rect 10457 8578 10473 8642
rect 10537 8597 10553 8642
rect 10617 8597 10633 8642
rect 10697 8597 10713 8642
rect 10777 8578 10793 8642
rect 10857 8597 10873 8642
rect 10937 8597 10953 8642
rect 11017 8597 11033 8642
rect 11097 8578 11113 8642
rect 11177 8597 11193 8642
rect 11257 8597 11273 8642
rect 11337 8597 11353 8642
rect 11417 8578 11433 8642
rect 11497 8597 11513 8642
rect 11577 8597 11593 8642
rect 11657 8597 11673 8642
rect 11737 8578 11753 8642
rect 11817 8597 11833 8642
rect 11897 8597 11913 8642
rect 11977 8597 12165 8642
rect 12229 8597 12246 8642
rect 12310 8597 12327 8642
rect 8816 8556 8901 8578
rect 9137 8556 9222 8578
rect 9458 8556 9543 8578
rect 9779 8556 9864 8578
rect 10100 8556 10185 8578
rect 10421 8556 10506 8578
rect 10742 8556 10827 8578
rect 11063 8556 11148 8578
rect 11384 8556 11469 8578
rect 11705 8556 11790 8578
rect 8816 8492 8859 8556
rect 9166 8492 9183 8556
rect 9490 8492 9507 8556
rect 9814 8492 9831 8556
rect 10137 8492 10153 8556
rect 10457 8492 10473 8556
rect 10777 8492 10793 8556
rect 11097 8492 11113 8556
rect 11417 8492 11433 8556
rect 11737 8492 11753 8556
rect 8816 8470 8901 8492
rect 9137 8470 9222 8492
rect 9458 8470 9543 8492
rect 9779 8470 9864 8492
rect 10100 8470 10185 8492
rect 10421 8470 10506 8492
rect 10742 8470 10827 8492
rect 11063 8470 11148 8492
rect 11384 8470 11469 8492
rect 11705 8470 11790 8492
rect 8816 8406 8859 8470
rect 9166 8406 9183 8470
rect 9490 8406 9507 8470
rect 9814 8406 9831 8470
rect 10137 8406 10153 8470
rect 10457 8406 10473 8470
rect 10777 8406 10793 8470
rect 11097 8406 11113 8470
rect 11417 8406 11433 8470
rect 11737 8406 11753 8470
rect 8816 8384 8901 8406
rect 9137 8384 9222 8406
rect 9458 8384 9543 8406
rect 9779 8384 9864 8406
rect 10100 8384 10185 8406
rect 10421 8384 10506 8406
rect 10742 8384 10827 8406
rect 11063 8384 11148 8406
rect 11384 8384 11469 8406
rect 11705 8384 11790 8406
rect 8816 8361 8859 8384
rect 7961 8323 7981 8361
rect 8045 8323 8065 8361
rect 8129 8323 8149 8361
rect 8213 8323 8859 8361
rect 7687 8320 8859 8323
rect 8923 8320 8940 8361
rect 9004 8320 9021 8361
rect 9085 8320 9102 8361
rect 9166 8320 9183 8384
rect 9247 8320 9264 8361
rect 9328 8320 9345 8361
rect 9409 8320 9426 8361
rect 9490 8320 9507 8384
rect 9571 8320 9588 8361
rect 9652 8320 9669 8361
rect 9733 8320 9750 8361
rect 9814 8320 9831 8384
rect 9895 8320 9912 8361
rect 9976 8320 9993 8361
rect 10057 8320 10073 8361
rect 10137 8320 10153 8384
rect 10217 8320 10233 8361
rect 10297 8320 10313 8361
rect 10377 8320 10393 8361
rect 10457 8320 10473 8384
rect 10537 8320 10553 8361
rect 10617 8320 10633 8361
rect 10697 8320 10713 8361
rect 10777 8320 10793 8384
rect 10857 8320 10873 8361
rect 10937 8320 10953 8361
rect 11017 8320 11033 8361
rect 11097 8320 11113 8384
rect 11177 8320 11193 8361
rect 11257 8320 11273 8361
rect 11337 8320 11353 8361
rect 11417 8320 11433 8384
rect 11497 8320 11513 8361
rect 11577 8320 11593 8361
rect 11657 8320 11673 8361
rect 11737 8320 11753 8384
rect 12026 8361 12111 8597
rect 12391 8578 12408 8642
rect 12472 8597 12489 8642
rect 12553 8597 12570 8642
rect 12634 8597 12651 8642
rect 12715 8578 12732 8642
rect 12796 8597 12813 8642
rect 12877 8597 12894 8642
rect 12958 8597 12975 8642
rect 13039 8578 13056 8642
rect 13120 8597 13137 8642
rect 13201 8597 13218 8642
rect 13282 8597 13299 8642
rect 13363 8578 13380 8642
rect 13444 8597 13461 8642
rect 13525 8597 13542 8642
rect 13606 8597 13623 8642
rect 13687 8578 13704 8642
rect 13768 8597 13785 8642
rect 13849 8597 13866 8642
rect 13930 8597 13947 8642
rect 14011 8578 14028 8642
rect 14092 8597 14109 8642
rect 14173 8597 14190 8642
rect 14254 8597 14271 8642
rect 14335 8578 14352 8642
rect 14416 8597 14433 8642
rect 14497 8597 14513 8642
rect 14577 8597 14593 8642
rect 14657 8578 14673 8642
rect 14737 8597 14753 8642
rect 14817 8597 14833 8642
rect 14897 8597 14913 8642
rect 14977 8578 14993 8642
rect 15057 8597 15073 8642
rect 15137 8597 15153 8642
rect 15217 8597 15233 8642
rect 15297 8578 15313 8642
rect 15377 8597 15393 8642
rect 15457 8597 15473 8642
rect 15537 8597 15553 8642
rect 15617 8578 16000 8642
rect 12347 8556 12432 8578
rect 12668 8556 12753 8578
rect 12989 8556 13074 8578
rect 13310 8556 13395 8578
rect 13631 8556 13716 8578
rect 13952 8556 14037 8578
rect 14273 8556 14358 8578
rect 14594 8556 14679 8578
rect 14915 8556 15000 8578
rect 15236 8556 15321 8578
rect 15557 8556 16000 8578
rect 12391 8492 12408 8556
rect 12715 8492 12732 8556
rect 13039 8492 13056 8556
rect 13363 8492 13380 8556
rect 13687 8492 13704 8556
rect 14011 8492 14028 8556
rect 14335 8492 14352 8556
rect 14657 8492 14673 8556
rect 14977 8492 14993 8556
rect 15297 8492 15313 8556
rect 15617 8492 16000 8556
rect 12347 8470 12432 8492
rect 12668 8470 12753 8492
rect 12989 8470 13074 8492
rect 13310 8470 13395 8492
rect 13631 8470 13716 8492
rect 13952 8470 14037 8492
rect 14273 8470 14358 8492
rect 14594 8470 14679 8492
rect 14915 8470 15000 8492
rect 15236 8470 15321 8492
rect 15557 8470 16000 8492
rect 12391 8406 12408 8470
rect 12715 8406 12732 8470
rect 13039 8406 13056 8470
rect 13363 8406 13380 8470
rect 13687 8406 13704 8470
rect 14011 8406 14028 8470
rect 14335 8406 14352 8470
rect 14657 8406 14673 8470
rect 14977 8406 14993 8470
rect 15297 8406 15313 8470
rect 15617 8406 16000 8470
rect 12347 8384 12432 8406
rect 12668 8384 12753 8406
rect 12989 8384 13074 8406
rect 13310 8384 13395 8406
rect 13631 8384 13716 8406
rect 13952 8384 14037 8406
rect 14273 8384 14358 8406
rect 14594 8384 14679 8406
rect 14915 8384 15000 8406
rect 15236 8384 15321 8406
rect 15557 8384 16000 8406
rect 11817 8320 11833 8361
rect 11897 8320 11913 8361
rect 11977 8320 12165 8361
rect 12229 8320 12246 8361
rect 12310 8320 12327 8361
rect 12391 8320 12408 8384
rect 12472 8320 12489 8361
rect 12553 8320 12570 8361
rect 12634 8320 12651 8361
rect 12715 8320 12732 8384
rect 12796 8320 12813 8361
rect 12877 8320 12894 8361
rect 12958 8320 12975 8361
rect 13039 8320 13056 8384
rect 13120 8320 13137 8361
rect 13201 8320 13218 8361
rect 13282 8320 13299 8361
rect 13363 8320 13380 8384
rect 13444 8320 13461 8361
rect 13525 8320 13542 8361
rect 13606 8320 13623 8361
rect 13687 8320 13704 8384
rect 13768 8320 13785 8361
rect 13849 8320 13866 8361
rect 13930 8320 13947 8361
rect 14011 8320 14028 8384
rect 14092 8320 14109 8361
rect 14173 8320 14190 8361
rect 14254 8320 14271 8361
rect 14335 8320 14352 8384
rect 14416 8320 14433 8361
rect 14497 8320 14513 8361
rect 14577 8320 14593 8361
rect 14657 8320 14673 8384
rect 14737 8320 14753 8361
rect 14817 8320 14833 8361
rect 14897 8320 14913 8361
rect 14977 8320 14993 8384
rect 15057 8320 15073 8361
rect 15137 8320 15153 8361
rect 15217 8320 15233 8361
rect 15297 8320 15313 8384
rect 15377 8320 15393 8361
rect 15457 8320 15473 8361
rect 15537 8320 15553 8361
rect 15617 8320 16000 8384
rect 0 8317 16000 8320
rect 0 7993 16000 8037
rect 0 7757 215 7993
rect 451 7757 537 7993
rect 773 7757 859 7993
rect 1095 7757 1181 7993
rect 1417 7757 1503 7993
rect 1739 7757 1825 7993
rect 2061 7757 2147 7993
rect 2383 7757 2469 7993
rect 2705 7757 2791 7993
rect 3027 7757 3113 7993
rect 3349 7757 3435 7993
rect 3671 7757 3757 7993
rect 3993 7757 4079 7993
rect 4315 7757 4401 7993
rect 4637 7757 4723 7993
rect 4959 7757 5045 7993
rect 5281 7757 5367 7993
rect 5603 7757 5689 7993
rect 5925 7757 6011 7993
rect 6247 7757 6332 7993
rect 6568 7757 6653 7993
rect 6889 7757 6974 7993
rect 7210 7757 7295 7993
rect 7531 7757 7616 7993
rect 7852 7757 7937 7993
rect 8173 7757 8258 7993
rect 8494 7757 8579 7993
rect 8815 7757 8900 7993
rect 9136 7757 9221 7993
rect 9457 7757 9542 7993
rect 9778 7757 9863 7993
rect 10099 7757 10184 7993
rect 10420 7757 10505 7993
rect 10741 7757 10826 7993
rect 11062 7757 11147 7993
rect 11383 7757 11468 7993
rect 11704 7757 11789 7993
rect 12025 7757 12110 7993
rect 12346 7757 12431 7993
rect 12667 7757 12752 7993
rect 12988 7757 13073 7993
rect 13309 7757 13394 7993
rect 13630 7757 13715 7993
rect 13951 7757 14036 7993
rect 14272 7757 14357 7993
rect 14593 7757 14678 7993
rect 14914 7757 14999 7993
rect 15235 7757 15320 7993
rect 15556 7757 16000 7993
rect 0 7627 16000 7757
rect 0 7391 215 7627
rect 451 7391 537 7627
rect 773 7391 859 7627
rect 1095 7391 1181 7627
rect 1417 7391 1503 7627
rect 1739 7391 1825 7627
rect 2061 7391 2147 7627
rect 2383 7391 2469 7627
rect 2705 7391 2791 7627
rect 3027 7391 3113 7627
rect 3349 7391 3435 7627
rect 3671 7391 3757 7627
rect 3993 7391 4079 7627
rect 4315 7391 4401 7627
rect 4637 7391 4723 7627
rect 4959 7391 5045 7627
rect 5281 7391 5367 7627
rect 5603 7391 5689 7627
rect 5925 7391 6011 7627
rect 6247 7391 6332 7627
rect 6568 7391 6653 7627
rect 6889 7391 6974 7627
rect 7210 7391 7295 7627
rect 7531 7391 7616 7627
rect 7852 7391 7937 7627
rect 8173 7391 8258 7627
rect 8494 7391 8579 7627
rect 8815 7391 8900 7627
rect 9136 7391 9221 7627
rect 9457 7391 9542 7627
rect 9778 7391 9863 7627
rect 10099 7391 10184 7627
rect 10420 7391 10505 7627
rect 10741 7391 10826 7627
rect 11062 7391 11147 7627
rect 11383 7391 11468 7627
rect 11704 7391 11789 7627
rect 12025 7391 12110 7627
rect 12346 7391 12431 7627
rect 12667 7391 12752 7627
rect 12988 7391 13073 7627
rect 13309 7391 13394 7627
rect 13630 7391 13715 7627
rect 13951 7391 14036 7627
rect 14272 7391 14357 7627
rect 14593 7391 14678 7627
rect 14914 7391 14999 7627
rect 15235 7391 15320 7627
rect 15556 7391 16000 7627
rect 0 7347 16000 7391
rect 0 7023 16000 7067
rect 0 6787 215 7023
rect 451 6787 537 7023
rect 773 6787 859 7023
rect 1095 6787 1181 7023
rect 1417 6787 1503 7023
rect 1739 6787 1825 7023
rect 2061 6787 2147 7023
rect 2383 6787 2469 7023
rect 2705 6787 2791 7023
rect 3027 6787 3113 7023
rect 3349 6787 3435 7023
rect 3671 6787 3757 7023
rect 3993 6787 4079 7023
rect 4315 6787 4401 7023
rect 4637 6787 4723 7023
rect 4959 6787 5045 7023
rect 5281 6787 5367 7023
rect 5603 6787 5689 7023
rect 5925 6787 6011 7023
rect 6247 6787 6332 7023
rect 6568 6787 6653 7023
rect 6889 6787 6974 7023
rect 7210 6787 7295 7023
rect 7531 6787 7616 7023
rect 7852 6787 7937 7023
rect 8173 6787 8258 7023
rect 8494 6787 8579 7023
rect 8815 6787 8900 7023
rect 9136 6787 9221 7023
rect 9457 6787 9542 7023
rect 9778 6787 9863 7023
rect 10099 6787 10184 7023
rect 10420 6787 10505 7023
rect 10741 6787 10826 7023
rect 11062 6787 11147 7023
rect 11383 6787 11468 7023
rect 11704 6787 11789 7023
rect 12025 6787 12110 7023
rect 12346 6787 12431 7023
rect 12667 6787 12752 7023
rect 12988 6787 13073 7023
rect 13309 6787 13394 7023
rect 13630 6787 13715 7023
rect 13951 6787 14036 7023
rect 14272 6787 14357 7023
rect 14593 6787 14678 7023
rect 14914 6787 14999 7023
rect 15235 6787 15320 7023
rect 15556 6787 16000 7023
rect 0 6657 16000 6787
rect 0 6421 215 6657
rect 451 6421 537 6657
rect 773 6421 859 6657
rect 1095 6421 1181 6657
rect 1417 6421 1503 6657
rect 1739 6421 1825 6657
rect 2061 6421 2147 6657
rect 2383 6421 2469 6657
rect 2705 6421 2791 6657
rect 3027 6421 3113 6657
rect 3349 6421 3435 6657
rect 3671 6421 3757 6657
rect 3993 6421 4079 6657
rect 4315 6421 4401 6657
rect 4637 6421 4723 6657
rect 4959 6421 5045 6657
rect 5281 6421 5367 6657
rect 5603 6421 5689 6657
rect 5925 6421 6011 6657
rect 6247 6421 6332 6657
rect 6568 6421 6653 6657
rect 6889 6421 6974 6657
rect 7210 6421 7295 6657
rect 7531 6421 7616 6657
rect 7852 6421 7937 6657
rect 8173 6421 8258 6657
rect 8494 6421 8579 6657
rect 8815 6421 8900 6657
rect 9136 6421 9221 6657
rect 9457 6421 9542 6657
rect 9778 6421 9863 6657
rect 10099 6421 10184 6657
rect 10420 6421 10505 6657
rect 10741 6421 10826 6657
rect 11062 6421 11147 6657
rect 11383 6421 11468 6657
rect 11704 6421 11789 6657
rect 12025 6421 12110 6657
rect 12346 6421 12431 6657
rect 12667 6421 12752 6657
rect 12988 6421 13073 6657
rect 13309 6421 13394 6657
rect 13630 6421 13715 6657
rect 13951 6421 14036 6657
rect 14272 6421 14357 6657
rect 14593 6421 14678 6657
rect 14914 6421 14999 6657
rect 15235 6421 15320 6657
rect 15556 6421 16000 6657
rect 0 6377 16000 6421
rect 0 6053 16000 6097
rect 0 5817 215 6053
rect 451 5817 537 6053
rect 773 5817 859 6053
rect 1095 5817 1181 6053
rect 1417 5817 1503 6053
rect 1739 5817 1825 6053
rect 2061 5817 2147 6053
rect 2383 5817 2469 6053
rect 2705 5817 2791 6053
rect 3027 5817 3113 6053
rect 3349 5817 3435 6053
rect 3671 5817 3757 6053
rect 3993 5817 4079 6053
rect 4315 5817 4401 6053
rect 4637 5817 4723 6053
rect 4959 5817 5045 6053
rect 5281 5817 5367 6053
rect 5603 5817 5689 6053
rect 5925 5817 6011 6053
rect 6247 5817 6332 6053
rect 6568 5817 6653 6053
rect 6889 5817 6974 6053
rect 7210 5817 7295 6053
rect 7531 5817 7616 6053
rect 7852 5817 7937 6053
rect 8173 5817 8258 6053
rect 8494 5817 8579 6053
rect 8815 5817 8900 6053
rect 9136 5817 9221 6053
rect 9457 5817 9542 6053
rect 9778 5817 9863 6053
rect 10099 5817 10184 6053
rect 10420 5817 10505 6053
rect 10741 5817 10826 6053
rect 11062 5817 11147 6053
rect 11383 5817 11468 6053
rect 11704 5817 11789 6053
rect 12025 5817 12110 6053
rect 12346 5817 12431 6053
rect 12667 5817 12752 6053
rect 12988 5817 13073 6053
rect 13309 5817 13394 6053
rect 13630 5817 13715 6053
rect 13951 5817 14036 6053
rect 14272 5817 14357 6053
rect 14593 5817 14678 6053
rect 14914 5817 14999 6053
rect 15235 5817 15320 6053
rect 15556 5817 16000 6053
rect 0 5447 16000 5817
rect 0 5211 215 5447
rect 451 5211 537 5447
rect 773 5211 859 5447
rect 1095 5211 1181 5447
rect 1417 5211 1503 5447
rect 1739 5211 1825 5447
rect 2061 5211 2147 5447
rect 2383 5211 2469 5447
rect 2705 5211 2791 5447
rect 3027 5211 3113 5447
rect 3349 5211 3435 5447
rect 3671 5211 3757 5447
rect 3993 5211 4079 5447
rect 4315 5211 4401 5447
rect 4637 5211 4723 5447
rect 4959 5211 5045 5447
rect 5281 5211 5367 5447
rect 5603 5211 5689 5447
rect 5925 5211 6011 5447
rect 6247 5211 6332 5447
rect 6568 5211 6653 5447
rect 6889 5211 6974 5447
rect 7210 5211 7295 5447
rect 7531 5211 7616 5447
rect 7852 5211 7937 5447
rect 8173 5211 8258 5447
rect 8494 5211 8579 5447
rect 8815 5211 8900 5447
rect 9136 5211 9221 5447
rect 9457 5211 9542 5447
rect 9778 5211 9863 5447
rect 10099 5211 10184 5447
rect 10420 5211 10505 5447
rect 10741 5211 10826 5447
rect 11062 5211 11147 5447
rect 11383 5211 11468 5447
rect 11704 5211 11789 5447
rect 12025 5211 12110 5447
rect 12346 5211 12431 5447
rect 12667 5211 12752 5447
rect 12988 5211 13073 5447
rect 13309 5211 13394 5447
rect 13630 5211 13715 5447
rect 13951 5211 14036 5447
rect 14272 5211 14357 5447
rect 14593 5211 14678 5447
rect 14914 5211 14999 5447
rect 15235 5211 15320 5447
rect 15556 5211 16000 5447
rect 0 5167 16000 5211
rect 0 4843 16000 4887
rect 0 4607 215 4843
rect 451 4607 537 4843
rect 773 4607 859 4843
rect 1095 4607 1181 4843
rect 1417 4607 1503 4843
rect 1739 4607 1825 4843
rect 2061 4607 2147 4843
rect 2383 4607 2469 4843
rect 2705 4607 2791 4843
rect 3027 4607 3113 4843
rect 3349 4607 3435 4843
rect 3671 4607 3757 4843
rect 3993 4607 4079 4843
rect 4315 4607 4401 4843
rect 4637 4607 4723 4843
rect 4959 4607 5045 4843
rect 5281 4607 5367 4843
rect 5603 4607 5689 4843
rect 5925 4607 6011 4843
rect 6247 4607 6332 4843
rect 6568 4607 6653 4843
rect 6889 4607 6974 4843
rect 7210 4607 7295 4843
rect 7531 4607 7616 4843
rect 7852 4607 7937 4843
rect 8173 4607 8258 4843
rect 8494 4607 8579 4843
rect 8815 4607 8900 4843
rect 9136 4607 9221 4843
rect 9457 4607 9542 4843
rect 9778 4607 9863 4843
rect 10099 4607 10184 4843
rect 10420 4607 10505 4843
rect 10741 4607 10826 4843
rect 11062 4607 11147 4843
rect 11383 4607 11468 4843
rect 11704 4607 11789 4843
rect 12025 4607 12110 4843
rect 12346 4607 12431 4843
rect 12667 4607 12752 4843
rect 12988 4607 13073 4843
rect 13309 4607 13394 4843
rect 13630 4607 13715 4843
rect 13951 4607 14036 4843
rect 14272 4607 14357 4843
rect 14593 4607 14678 4843
rect 14914 4607 14999 4843
rect 15235 4607 15320 4843
rect 15556 4607 16000 4843
rect 0 4237 16000 4607
rect 0 4001 215 4237
rect 451 4001 537 4237
rect 773 4001 859 4237
rect 1095 4001 1181 4237
rect 1417 4001 1503 4237
rect 1739 4001 1825 4237
rect 2061 4001 2147 4237
rect 2383 4001 2469 4237
rect 2705 4001 2791 4237
rect 3027 4001 3113 4237
rect 3349 4001 3435 4237
rect 3671 4001 3757 4237
rect 3993 4001 4079 4237
rect 4315 4001 4401 4237
rect 4637 4001 4723 4237
rect 4959 4001 5045 4237
rect 5281 4001 5367 4237
rect 5603 4001 5689 4237
rect 5925 4001 6011 4237
rect 6247 4001 6332 4237
rect 6568 4001 6653 4237
rect 6889 4001 6974 4237
rect 7210 4001 7295 4237
rect 7531 4001 7616 4237
rect 7852 4001 7937 4237
rect 8173 4001 8258 4237
rect 8494 4001 8579 4237
rect 8815 4001 8900 4237
rect 9136 4001 9221 4237
rect 9457 4001 9542 4237
rect 9778 4001 9863 4237
rect 10099 4001 10184 4237
rect 10420 4001 10505 4237
rect 10741 4001 10826 4237
rect 11062 4001 11147 4237
rect 11383 4001 11468 4237
rect 11704 4001 11789 4237
rect 12025 4001 12110 4237
rect 12346 4001 12431 4237
rect 12667 4001 12752 4237
rect 12988 4001 13073 4237
rect 13309 4001 13394 4237
rect 13630 4001 13715 4237
rect 13951 4001 14036 4237
rect 14272 4001 14357 4237
rect 14593 4001 14678 4237
rect 14914 4001 14999 4237
rect 15235 4001 15320 4237
rect 15556 4001 16000 4237
rect 0 3957 16000 4001
rect 0 3633 16000 3677
rect 0 3397 215 3633
rect 451 3397 537 3633
rect 773 3397 859 3633
rect 1095 3397 1181 3633
rect 1417 3397 1503 3633
rect 1739 3397 1825 3633
rect 2061 3397 2147 3633
rect 2383 3397 2469 3633
rect 2705 3397 2791 3633
rect 3027 3397 3113 3633
rect 3349 3397 3435 3633
rect 3671 3397 3757 3633
rect 3993 3397 4079 3633
rect 4315 3397 4401 3633
rect 4637 3397 4723 3633
rect 4959 3397 5045 3633
rect 5281 3397 5367 3633
rect 5603 3397 5689 3633
rect 5925 3397 6011 3633
rect 6247 3397 6332 3633
rect 6568 3397 6653 3633
rect 6889 3397 6974 3633
rect 7210 3397 7295 3633
rect 7531 3397 7616 3633
rect 7852 3397 7937 3633
rect 8173 3397 8258 3633
rect 8494 3397 8579 3633
rect 8815 3397 8900 3633
rect 9136 3397 9221 3633
rect 9457 3397 9542 3633
rect 9778 3397 9863 3633
rect 10099 3397 10184 3633
rect 10420 3397 10505 3633
rect 10741 3397 10826 3633
rect 11062 3397 11147 3633
rect 11383 3397 11468 3633
rect 11704 3397 11789 3633
rect 12025 3397 12110 3633
rect 12346 3397 12431 3633
rect 12667 3397 12752 3633
rect 12988 3397 13073 3633
rect 13309 3397 13394 3633
rect 13630 3397 13715 3633
rect 13951 3397 14036 3633
rect 14272 3397 14357 3633
rect 14593 3397 14678 3633
rect 14914 3397 14999 3633
rect 15235 3397 15320 3633
rect 15556 3397 16000 3633
rect 0 3267 16000 3397
rect 0 3031 215 3267
rect 451 3031 537 3267
rect 773 3031 859 3267
rect 1095 3031 1181 3267
rect 1417 3031 1503 3267
rect 1739 3031 1825 3267
rect 2061 3031 2147 3267
rect 2383 3031 2469 3267
rect 2705 3031 2791 3267
rect 3027 3031 3113 3267
rect 3349 3031 3435 3267
rect 3671 3031 3757 3267
rect 3993 3031 4079 3267
rect 4315 3031 4401 3267
rect 4637 3031 4723 3267
rect 4959 3031 5045 3267
rect 5281 3031 5367 3267
rect 5603 3031 5689 3267
rect 5925 3031 6011 3267
rect 6247 3031 6332 3267
rect 6568 3031 6653 3267
rect 6889 3031 6974 3267
rect 7210 3031 7295 3267
rect 7531 3031 7616 3267
rect 7852 3031 7937 3267
rect 8173 3031 8258 3267
rect 8494 3031 8579 3267
rect 8815 3031 8900 3267
rect 9136 3031 9221 3267
rect 9457 3031 9542 3267
rect 9778 3031 9863 3267
rect 10099 3031 10184 3267
rect 10420 3031 10505 3267
rect 10741 3031 10826 3267
rect 11062 3031 11147 3267
rect 11383 3031 11468 3267
rect 11704 3031 11789 3267
rect 12025 3031 12110 3267
rect 12346 3031 12431 3267
rect 12667 3031 12752 3267
rect 12988 3031 13073 3267
rect 13309 3031 13394 3267
rect 13630 3031 13715 3267
rect 13951 3031 14036 3267
rect 14272 3031 14357 3267
rect 14593 3031 14678 3267
rect 14914 3031 14999 3267
rect 15235 3031 15320 3267
rect 15556 3031 16000 3267
rect 0 2987 16000 3031
rect 0 2701 16000 2707
rect 0 2663 547 2701
rect 611 2663 659 2701
rect 723 2663 771 2701
rect 835 2663 883 2701
rect 947 2663 11674 2701
rect 11738 2663 16000 2701
rect 0 2427 215 2663
rect 451 2427 537 2663
rect 835 2637 859 2663
rect 773 2579 859 2637
rect 835 2515 859 2579
rect 773 2457 859 2515
rect 835 2427 859 2457
rect 1095 2427 1181 2663
rect 1417 2427 1503 2663
rect 1739 2427 1825 2663
rect 2061 2427 2147 2663
rect 2383 2427 2469 2663
rect 2705 2427 2791 2663
rect 3027 2427 3113 2663
rect 3349 2427 3435 2663
rect 3671 2427 3757 2663
rect 3993 2427 4079 2663
rect 4315 2427 4401 2663
rect 4637 2427 4723 2663
rect 4959 2427 5045 2663
rect 5281 2427 5367 2663
rect 5603 2427 5689 2663
rect 5925 2427 6011 2663
rect 6247 2427 6332 2663
rect 6568 2427 6653 2663
rect 6889 2427 6974 2663
rect 7210 2427 7295 2663
rect 7531 2427 7616 2663
rect 7852 2427 7937 2663
rect 8173 2427 8258 2663
rect 8494 2427 8579 2663
rect 8815 2427 8900 2663
rect 9136 2427 9221 2663
rect 9457 2427 9542 2663
rect 9778 2427 9863 2663
rect 10099 2427 10184 2663
rect 10420 2427 10505 2663
rect 10741 2427 10826 2663
rect 11062 2427 11147 2663
rect 11383 2427 11468 2663
rect 11738 2637 11789 2663
rect 11704 2579 11789 2637
rect 11738 2515 11789 2579
rect 11704 2457 11789 2515
rect 11738 2427 11789 2457
rect 12025 2427 12110 2663
rect 12346 2427 12431 2663
rect 12667 2427 12752 2663
rect 12988 2427 13073 2663
rect 13309 2427 13394 2663
rect 13630 2427 13715 2663
rect 13951 2427 14036 2663
rect 14272 2427 14357 2663
rect 14593 2427 14678 2663
rect 14914 2427 14999 2663
rect 15235 2427 15320 2663
rect 15556 2427 16000 2663
rect 0 2393 547 2427
rect 611 2393 659 2427
rect 723 2393 771 2427
rect 835 2393 883 2427
rect 947 2393 11674 2427
rect 11738 2393 16000 2427
rect 0 2335 16000 2393
rect 0 2271 547 2335
rect 611 2271 659 2335
rect 723 2271 771 2335
rect 835 2271 883 2335
rect 947 2271 11674 2335
rect 11738 2271 16000 2335
rect 0 2213 16000 2271
rect 0 2149 547 2213
rect 611 2149 659 2213
rect 723 2149 771 2213
rect 835 2149 883 2213
rect 947 2149 11674 2213
rect 11738 2149 16000 2213
rect 0 2091 16000 2149
rect 0 2057 547 2091
rect 611 2057 659 2091
rect 723 2057 771 2091
rect 835 2057 883 2091
rect 947 2057 11674 2091
rect 11738 2057 16000 2091
rect 0 1821 215 2057
rect 451 1821 537 2057
rect 835 2027 859 2057
rect 773 1969 859 2027
rect 835 1905 859 1969
rect 773 1847 859 1905
rect 835 1821 859 1847
rect 1095 1821 1181 2057
rect 1417 1821 1503 2057
rect 1739 1821 1825 2057
rect 2061 1821 2147 2057
rect 2383 1821 2469 2057
rect 2705 1821 2791 2057
rect 3027 1821 3113 2057
rect 3349 1821 3435 2057
rect 3671 1821 3757 2057
rect 3993 1821 4079 2057
rect 4315 1821 4401 2057
rect 4637 1821 4723 2057
rect 4959 1821 5045 2057
rect 5281 1821 5367 2057
rect 5603 1821 5689 2057
rect 5925 1821 6011 2057
rect 6247 1821 6332 2057
rect 6568 1821 6653 2057
rect 6889 1821 6974 2057
rect 7210 1821 7295 2057
rect 7531 1821 7616 2057
rect 7852 1821 7937 2057
rect 8173 1821 8258 2057
rect 8494 1821 8579 2057
rect 8815 1821 8900 2057
rect 9136 1821 9221 2057
rect 9457 1821 9542 2057
rect 9778 1821 9863 2057
rect 10099 1821 10184 2057
rect 10420 1821 10505 2057
rect 10741 1821 10826 2057
rect 11062 1821 11147 2057
rect 11383 1821 11468 2057
rect 11738 2027 11789 2057
rect 11704 1969 11789 2027
rect 11738 1905 11789 1969
rect 11704 1847 11789 1905
rect 11738 1821 11789 1847
rect 12025 1821 12110 2057
rect 12346 1821 12431 2057
rect 12667 1821 12752 2057
rect 12988 1821 13073 2057
rect 13309 1821 13394 2057
rect 13630 1821 13715 2057
rect 13951 1821 14036 2057
rect 14272 1821 14357 2057
rect 14593 1821 14678 2057
rect 14914 1821 14999 2057
rect 15235 1821 15320 2057
rect 15556 1821 16000 2057
rect 0 1783 547 1821
rect 611 1783 659 1821
rect 723 1783 771 1821
rect 835 1783 883 1821
rect 947 1783 11674 1821
rect 11738 1783 16000 1821
rect 0 1777 16000 1783
rect 0 1452 16000 1497
rect 0 1216 215 1452
rect 451 1216 537 1452
rect 773 1216 859 1452
rect 1095 1216 1181 1452
rect 1417 1216 1503 1452
rect 1739 1216 1825 1452
rect 2061 1216 2147 1452
rect 2383 1216 2469 1452
rect 2705 1216 2791 1452
rect 3027 1216 3113 1452
rect 3349 1216 3435 1452
rect 3671 1216 3757 1452
rect 3993 1216 4079 1452
rect 4315 1216 4401 1452
rect 4637 1216 4723 1452
rect 4959 1216 5045 1452
rect 5281 1216 5367 1452
rect 5603 1216 5689 1452
rect 5925 1216 6011 1452
rect 6247 1216 6332 1452
rect 6568 1216 6653 1452
rect 6889 1216 6974 1452
rect 7210 1216 7295 1452
rect 7531 1216 7616 1452
rect 7852 1216 7937 1452
rect 8173 1216 8258 1452
rect 8494 1216 8579 1452
rect 8815 1216 8900 1452
rect 9136 1216 9221 1452
rect 9457 1216 9542 1452
rect 9778 1216 9863 1452
rect 10099 1216 10184 1452
rect 10420 1216 10505 1452
rect 10741 1216 10826 1452
rect 11062 1216 11147 1452
rect 11383 1216 11468 1452
rect 11704 1216 11789 1452
rect 12025 1216 12110 1452
rect 12346 1216 12431 1452
rect 12667 1216 12752 1452
rect 12988 1216 13073 1452
rect 13309 1216 13394 1452
rect 13630 1216 13715 1452
rect 13951 1216 14036 1452
rect 14272 1216 14357 1452
rect 14593 1216 14678 1452
rect 14914 1216 14999 1452
rect 15235 1216 15320 1452
rect 15556 1216 16000 1452
rect 0 1070 16000 1216
rect 0 834 215 1070
rect 451 834 537 1070
rect 773 834 859 1070
rect 1095 834 1181 1070
rect 1417 834 1503 1070
rect 1739 834 1825 1070
rect 2061 834 2147 1070
rect 2383 834 2469 1070
rect 2705 834 2791 1070
rect 3027 834 3113 1070
rect 3349 834 3435 1070
rect 3671 834 3757 1070
rect 3993 834 4079 1070
rect 4315 834 4401 1070
rect 4637 834 4723 1070
rect 4959 834 5045 1070
rect 5281 834 5367 1070
rect 5603 834 5689 1070
rect 5925 834 6011 1070
rect 6247 834 6332 1070
rect 6568 834 6653 1070
rect 6889 834 6974 1070
rect 7210 834 7295 1070
rect 7531 834 7616 1070
rect 7852 834 7937 1070
rect 8173 834 8258 1070
rect 8494 834 8579 1070
rect 8815 834 8900 1070
rect 9136 834 9221 1070
rect 9457 834 9542 1070
rect 9778 834 9863 1070
rect 10099 834 10184 1070
rect 10420 834 10505 1070
rect 10741 834 10826 1070
rect 11062 834 11147 1070
rect 11383 834 11468 1070
rect 11704 834 11789 1070
rect 12025 834 12110 1070
rect 12346 834 12431 1070
rect 12667 834 12752 1070
rect 12988 834 13073 1070
rect 13309 834 13394 1070
rect 13630 834 13715 1070
rect 13951 834 14036 1070
rect 14272 834 14357 1070
rect 14593 834 14678 1070
rect 14914 834 14999 1070
rect 15235 834 15320 1070
rect 15556 834 16000 1070
rect 0 688 16000 834
rect 0 452 215 688
rect 451 452 537 688
rect 773 452 859 688
rect 1095 452 1181 688
rect 1417 452 1503 688
rect 1739 452 1825 688
rect 2061 452 2147 688
rect 2383 452 2469 688
rect 2705 452 2791 688
rect 3027 452 3113 688
rect 3349 452 3435 688
rect 3671 452 3757 688
rect 3993 452 4079 688
rect 4315 452 4401 688
rect 4637 452 4723 688
rect 4959 452 5045 688
rect 5281 452 5367 688
rect 5603 452 5689 688
rect 5925 452 6011 688
rect 6247 452 6332 688
rect 6568 452 6653 688
rect 6889 452 6974 688
rect 7210 452 7295 688
rect 7531 452 7616 688
rect 7852 452 7937 688
rect 8173 452 8258 688
rect 8494 452 8579 688
rect 8815 452 8900 688
rect 9136 452 9221 688
rect 9457 452 9542 688
rect 9778 452 9863 688
rect 10099 452 10184 688
rect 10420 452 10505 688
rect 10741 452 10826 688
rect 11062 452 11147 688
rect 11383 452 11468 688
rect 11704 452 11789 688
rect 12025 452 12110 688
rect 12346 452 12431 688
rect 12667 452 12752 688
rect 12988 452 13073 688
rect 13309 452 13394 688
rect 13630 452 13715 688
rect 13951 452 14036 688
rect 14272 452 14357 688
rect 14593 452 14678 688
rect 14914 452 14999 688
rect 15235 452 15320 688
rect 15556 452 16000 688
rect 0 407 16000 452
<< via4 >>
rect 215 39728 451 39964
rect 537 39728 773 39964
rect 859 39728 1095 39964
rect 1181 39728 1417 39964
rect 1503 39728 1739 39964
rect 1825 39728 2061 39964
rect 2147 39728 2383 39964
rect 2469 39728 2705 39964
rect 2791 39728 3027 39964
rect 3113 39728 3349 39964
rect 3435 39728 3671 39964
rect 3757 39728 3993 39964
rect 4079 39728 4315 39964
rect 4401 39728 4637 39964
rect 4723 39728 4959 39964
rect 5045 39728 5281 39964
rect 5367 39728 5603 39964
rect 5689 39728 5925 39964
rect 6011 39728 6247 39964
rect 6332 39728 6568 39964
rect 6653 39728 6889 39964
rect 6974 39728 7210 39964
rect 7295 39728 7531 39964
rect 7616 39728 7852 39964
rect 7937 39728 8173 39964
rect 8258 39728 8494 39964
rect 8579 39728 8815 39964
rect 8900 39728 9136 39964
rect 9221 39728 9457 39964
rect 9542 39728 9778 39964
rect 9863 39728 10099 39964
rect 10184 39728 10420 39964
rect 10505 39728 10741 39964
rect 10826 39728 11062 39964
rect 11147 39728 11383 39964
rect 11468 39728 11704 39964
rect 11789 39728 12025 39964
rect 12110 39728 12346 39964
rect 12431 39728 12667 39964
rect 12752 39728 12988 39964
rect 13073 39728 13309 39964
rect 13394 39728 13630 39964
rect 13715 39728 13951 39964
rect 14036 39728 14272 39964
rect 14357 39728 14593 39964
rect 14678 39728 14914 39964
rect 14999 39728 15235 39964
rect 15320 39728 15556 39964
rect 215 39404 451 39640
rect 537 39404 773 39640
rect 859 39404 1095 39640
rect 1181 39404 1417 39640
rect 1503 39404 1739 39640
rect 1825 39404 2061 39640
rect 2147 39404 2383 39640
rect 2469 39404 2705 39640
rect 2791 39404 3027 39640
rect 3113 39404 3349 39640
rect 3435 39404 3671 39640
rect 3757 39404 3993 39640
rect 4079 39404 4315 39640
rect 4401 39404 4637 39640
rect 4723 39404 4959 39640
rect 5045 39404 5281 39640
rect 5367 39404 5603 39640
rect 5689 39404 5925 39640
rect 6011 39404 6247 39640
rect 6332 39404 6568 39640
rect 6653 39404 6889 39640
rect 6974 39404 7210 39640
rect 7295 39404 7531 39640
rect 7616 39404 7852 39640
rect 7937 39404 8173 39640
rect 8258 39404 8494 39640
rect 8579 39404 8815 39640
rect 8900 39404 9136 39640
rect 9221 39404 9457 39640
rect 9542 39404 9778 39640
rect 9863 39404 10099 39640
rect 10184 39404 10420 39640
rect 10505 39404 10741 39640
rect 10826 39404 11062 39640
rect 11147 39404 11383 39640
rect 11468 39404 11704 39640
rect 11789 39404 12025 39640
rect 12110 39404 12346 39640
rect 12431 39404 12667 39640
rect 12752 39404 12988 39640
rect 13073 39404 13309 39640
rect 13394 39404 13630 39640
rect 13715 39404 13951 39640
rect 14036 39404 14272 39640
rect 14357 39404 14593 39640
rect 14678 39404 14914 39640
rect 14999 39404 15235 39640
rect 15320 39404 15556 39640
rect 215 39080 451 39316
rect 537 39080 773 39316
rect 859 39080 1095 39316
rect 1181 39080 1417 39316
rect 1503 39080 1739 39316
rect 1825 39080 2061 39316
rect 2147 39080 2383 39316
rect 2469 39080 2705 39316
rect 2791 39080 3027 39316
rect 3113 39080 3349 39316
rect 3435 39080 3671 39316
rect 3757 39080 3993 39316
rect 4079 39080 4315 39316
rect 4401 39080 4637 39316
rect 4723 39080 4959 39316
rect 5045 39080 5281 39316
rect 5367 39080 5603 39316
rect 5689 39080 5925 39316
rect 6011 39080 6247 39316
rect 6332 39080 6568 39316
rect 6653 39080 6889 39316
rect 6974 39080 7210 39316
rect 7295 39080 7531 39316
rect 7616 39080 7852 39316
rect 7937 39080 8173 39316
rect 8258 39080 8494 39316
rect 8579 39080 8815 39316
rect 8900 39080 9136 39316
rect 9221 39080 9457 39316
rect 9542 39080 9778 39316
rect 9863 39080 10099 39316
rect 10184 39080 10420 39316
rect 10505 39080 10741 39316
rect 10826 39080 11062 39316
rect 11147 39080 11383 39316
rect 11468 39080 11704 39316
rect 11789 39080 12025 39316
rect 12110 39080 12346 39316
rect 12431 39080 12667 39316
rect 12752 39080 12988 39316
rect 13073 39080 13309 39316
rect 13394 39080 13630 39316
rect 13715 39080 13951 39316
rect 14036 39080 14272 39316
rect 14357 39080 14593 39316
rect 14678 39080 14914 39316
rect 14999 39080 15235 39316
rect 15320 39080 15556 39316
rect 215 38756 451 38992
rect 537 38756 773 38992
rect 859 38756 1095 38992
rect 1181 38756 1417 38992
rect 1503 38756 1739 38992
rect 1825 38756 2061 38992
rect 2147 38756 2383 38992
rect 2469 38756 2705 38992
rect 2791 38756 3027 38992
rect 3113 38756 3349 38992
rect 3435 38756 3671 38992
rect 3757 38756 3993 38992
rect 4079 38756 4315 38992
rect 4401 38756 4637 38992
rect 4723 38756 4959 38992
rect 5045 38756 5281 38992
rect 5367 38756 5603 38992
rect 5689 38756 5925 38992
rect 6011 38756 6247 38992
rect 6332 38756 6568 38992
rect 6653 38756 6889 38992
rect 6974 38756 7210 38992
rect 7295 38756 7531 38992
rect 7616 38756 7852 38992
rect 7937 38756 8173 38992
rect 8258 38756 8494 38992
rect 8579 38756 8815 38992
rect 8900 38756 9136 38992
rect 9221 38756 9457 38992
rect 9542 38756 9778 38992
rect 9863 38756 10099 38992
rect 10184 38756 10420 38992
rect 10505 38756 10741 38992
rect 10826 38756 11062 38992
rect 11147 38756 11383 38992
rect 11468 38756 11704 38992
rect 11789 38756 12025 38992
rect 12110 38756 12346 38992
rect 12431 38756 12667 38992
rect 12752 38756 12988 38992
rect 13073 38756 13309 38992
rect 13394 38756 13630 38992
rect 13715 38756 13951 38992
rect 14036 38756 14272 38992
rect 14357 38756 14593 38992
rect 14678 38756 14914 38992
rect 14999 38756 15235 38992
rect 15320 38756 15556 38992
rect 215 38432 451 38668
rect 537 38432 773 38668
rect 859 38432 1095 38668
rect 1181 38432 1417 38668
rect 1503 38432 1739 38668
rect 1825 38432 2061 38668
rect 2147 38432 2383 38668
rect 2469 38432 2705 38668
rect 2791 38432 3027 38668
rect 3113 38432 3349 38668
rect 3435 38432 3671 38668
rect 3757 38432 3993 38668
rect 4079 38432 4315 38668
rect 4401 38432 4637 38668
rect 4723 38432 4959 38668
rect 5045 38432 5281 38668
rect 5367 38432 5603 38668
rect 5689 38432 5925 38668
rect 6011 38432 6247 38668
rect 6332 38432 6568 38668
rect 6653 38432 6889 38668
rect 6974 38432 7210 38668
rect 7295 38432 7531 38668
rect 7616 38432 7852 38668
rect 7937 38432 8173 38668
rect 8258 38432 8494 38668
rect 8579 38432 8815 38668
rect 8900 38432 9136 38668
rect 9221 38432 9457 38668
rect 9542 38432 9778 38668
rect 9863 38432 10099 38668
rect 10184 38432 10420 38668
rect 10505 38432 10741 38668
rect 10826 38432 11062 38668
rect 11147 38432 11383 38668
rect 11468 38432 11704 38668
rect 11789 38432 12025 38668
rect 12110 38432 12346 38668
rect 12431 38432 12667 38668
rect 12752 38432 12988 38668
rect 13073 38432 13309 38668
rect 13394 38432 13630 38668
rect 13715 38432 13951 38668
rect 14036 38432 14272 38668
rect 14357 38432 14593 38668
rect 14678 38432 14914 38668
rect 14999 38432 15235 38668
rect 15320 38432 15556 38668
rect 215 38108 451 38344
rect 537 38108 773 38344
rect 859 38108 1095 38344
rect 1181 38108 1417 38344
rect 1503 38108 1739 38344
rect 1825 38108 2061 38344
rect 2147 38108 2383 38344
rect 2469 38108 2705 38344
rect 2791 38108 3027 38344
rect 3113 38108 3349 38344
rect 3435 38108 3671 38344
rect 3757 38108 3993 38344
rect 4079 38108 4315 38344
rect 4401 38108 4637 38344
rect 4723 38108 4959 38344
rect 5045 38108 5281 38344
rect 5367 38108 5603 38344
rect 5689 38108 5925 38344
rect 6011 38108 6247 38344
rect 6332 38108 6568 38344
rect 6653 38108 6889 38344
rect 6974 38108 7210 38344
rect 7295 38108 7531 38344
rect 7616 38108 7852 38344
rect 7937 38108 8173 38344
rect 8258 38108 8494 38344
rect 8579 38108 8815 38344
rect 8900 38108 9136 38344
rect 9221 38108 9457 38344
rect 9542 38108 9778 38344
rect 9863 38108 10099 38344
rect 10184 38108 10420 38344
rect 10505 38108 10741 38344
rect 10826 38108 11062 38344
rect 11147 38108 11383 38344
rect 11468 38108 11704 38344
rect 11789 38108 12025 38344
rect 12110 38108 12346 38344
rect 12431 38108 12667 38344
rect 12752 38108 12988 38344
rect 13073 38108 13309 38344
rect 13394 38108 13630 38344
rect 13715 38108 13951 38344
rect 14036 38108 14272 38344
rect 14357 38108 14593 38344
rect 14678 38108 14914 38344
rect 14999 38108 15235 38344
rect 15320 38108 15556 38344
rect 215 37784 451 38020
rect 537 37784 773 38020
rect 859 37784 1095 38020
rect 1181 37784 1417 38020
rect 1503 37784 1739 38020
rect 1825 37784 2061 38020
rect 2147 37784 2383 38020
rect 2469 37784 2705 38020
rect 2791 37784 3027 38020
rect 3113 37784 3349 38020
rect 3435 37784 3671 38020
rect 3757 37784 3993 38020
rect 4079 37784 4315 38020
rect 4401 37784 4637 38020
rect 4723 37784 4959 38020
rect 5045 37784 5281 38020
rect 5367 37784 5603 38020
rect 5689 37784 5925 38020
rect 6011 37784 6247 38020
rect 6332 37784 6568 38020
rect 6653 37784 6889 38020
rect 6974 37784 7210 38020
rect 7295 37784 7531 38020
rect 7616 37784 7852 38020
rect 7937 37784 8173 38020
rect 8258 37784 8494 38020
rect 8579 37784 8815 38020
rect 8900 37784 9136 38020
rect 9221 37784 9457 38020
rect 9542 37784 9778 38020
rect 9863 37784 10099 38020
rect 10184 37784 10420 38020
rect 10505 37784 10741 38020
rect 10826 37784 11062 38020
rect 11147 37784 11383 38020
rect 11468 37784 11704 38020
rect 11789 37784 12025 38020
rect 12110 37784 12346 38020
rect 12431 37784 12667 38020
rect 12752 37784 12988 38020
rect 13073 37784 13309 38020
rect 13394 37784 13630 38020
rect 13715 37784 13951 38020
rect 14036 37784 14272 38020
rect 14357 37784 14593 38020
rect 14678 37784 14914 38020
rect 14999 37784 15235 38020
rect 15320 37784 15556 38020
rect 215 37460 451 37696
rect 537 37460 773 37696
rect 859 37460 1095 37696
rect 1181 37460 1417 37696
rect 1503 37460 1739 37696
rect 1825 37460 2061 37696
rect 2147 37460 2383 37696
rect 2469 37460 2705 37696
rect 2791 37460 3027 37696
rect 3113 37460 3349 37696
rect 3435 37460 3671 37696
rect 3757 37460 3993 37696
rect 4079 37460 4315 37696
rect 4401 37460 4637 37696
rect 4723 37460 4959 37696
rect 5045 37460 5281 37696
rect 5367 37460 5603 37696
rect 5689 37460 5925 37696
rect 6011 37460 6247 37696
rect 6332 37460 6568 37696
rect 6653 37460 6889 37696
rect 6974 37460 7210 37696
rect 7295 37460 7531 37696
rect 7616 37460 7852 37696
rect 7937 37460 8173 37696
rect 8258 37460 8494 37696
rect 8579 37460 8815 37696
rect 8900 37460 9136 37696
rect 9221 37460 9457 37696
rect 9542 37460 9778 37696
rect 9863 37460 10099 37696
rect 10184 37460 10420 37696
rect 10505 37460 10741 37696
rect 10826 37460 11062 37696
rect 11147 37460 11383 37696
rect 11468 37460 11704 37696
rect 11789 37460 12025 37696
rect 12110 37460 12346 37696
rect 12431 37460 12667 37696
rect 12752 37460 12988 37696
rect 13073 37460 13309 37696
rect 13394 37460 13630 37696
rect 13715 37460 13951 37696
rect 14036 37460 14272 37696
rect 14357 37460 14593 37696
rect 14678 37460 14914 37696
rect 14999 37460 15235 37696
rect 15320 37460 15556 37696
rect 215 37136 451 37372
rect 537 37136 773 37372
rect 859 37136 1095 37372
rect 1181 37136 1417 37372
rect 1503 37136 1739 37372
rect 1825 37136 2061 37372
rect 2147 37136 2383 37372
rect 2469 37136 2705 37372
rect 2791 37136 3027 37372
rect 3113 37136 3349 37372
rect 3435 37136 3671 37372
rect 3757 37136 3993 37372
rect 4079 37136 4315 37372
rect 4401 37136 4637 37372
rect 4723 37136 4959 37372
rect 5045 37136 5281 37372
rect 5367 37136 5603 37372
rect 5689 37136 5925 37372
rect 6011 37136 6247 37372
rect 6332 37136 6568 37372
rect 6653 37136 6889 37372
rect 6974 37136 7210 37372
rect 7295 37136 7531 37372
rect 7616 37136 7852 37372
rect 7937 37136 8173 37372
rect 8258 37136 8494 37372
rect 8579 37136 8815 37372
rect 8900 37136 9136 37372
rect 9221 37136 9457 37372
rect 9542 37136 9778 37372
rect 9863 37136 10099 37372
rect 10184 37136 10420 37372
rect 10505 37136 10741 37372
rect 10826 37136 11062 37372
rect 11147 37136 11383 37372
rect 11468 37136 11704 37372
rect 11789 37136 12025 37372
rect 12110 37136 12346 37372
rect 12431 37136 12667 37372
rect 12752 37136 12988 37372
rect 13073 37136 13309 37372
rect 13394 37136 13630 37372
rect 13715 37136 13951 37372
rect 14036 37136 14272 37372
rect 14357 37136 14593 37372
rect 14678 37136 14914 37372
rect 14999 37136 15235 37372
rect 15320 37136 15556 37372
rect 215 36812 451 37048
rect 537 36812 773 37048
rect 859 36812 1095 37048
rect 1181 36812 1417 37048
rect 1503 36812 1739 37048
rect 1825 36812 2061 37048
rect 2147 36812 2383 37048
rect 2469 36812 2705 37048
rect 2791 36812 3027 37048
rect 3113 36812 3349 37048
rect 3435 36812 3671 37048
rect 3757 36812 3993 37048
rect 4079 36812 4315 37048
rect 4401 36812 4637 37048
rect 4723 36812 4959 37048
rect 5045 36812 5281 37048
rect 5367 36812 5603 37048
rect 5689 36812 5925 37048
rect 6011 36812 6247 37048
rect 6332 36812 6568 37048
rect 6653 36812 6889 37048
rect 6974 36812 7210 37048
rect 7295 36812 7531 37048
rect 7616 36812 7852 37048
rect 7937 36812 8173 37048
rect 8258 36812 8494 37048
rect 8579 36812 8815 37048
rect 8900 36812 9136 37048
rect 9221 36812 9457 37048
rect 9542 36812 9778 37048
rect 9863 36812 10099 37048
rect 10184 36812 10420 37048
rect 10505 36812 10741 37048
rect 10826 36812 11062 37048
rect 11147 36812 11383 37048
rect 11468 36812 11704 37048
rect 11789 36812 12025 37048
rect 12110 36812 12346 37048
rect 12431 36812 12667 37048
rect 12752 36812 12988 37048
rect 13073 36812 13309 37048
rect 13394 36812 13630 37048
rect 13715 36812 13951 37048
rect 14036 36812 14272 37048
rect 14357 36812 14593 37048
rect 14678 36812 14914 37048
rect 14999 36812 15235 37048
rect 15320 36812 15556 37048
rect 215 36488 451 36724
rect 537 36488 773 36724
rect 859 36488 1095 36724
rect 1181 36488 1417 36724
rect 1503 36488 1739 36724
rect 1825 36488 2061 36724
rect 2147 36488 2383 36724
rect 2469 36488 2705 36724
rect 2791 36488 3027 36724
rect 3113 36488 3349 36724
rect 3435 36488 3671 36724
rect 3757 36488 3993 36724
rect 4079 36488 4315 36724
rect 4401 36488 4637 36724
rect 4723 36488 4959 36724
rect 5045 36488 5281 36724
rect 5367 36488 5603 36724
rect 5689 36488 5925 36724
rect 6011 36488 6247 36724
rect 6332 36488 6568 36724
rect 6653 36488 6889 36724
rect 6974 36488 7210 36724
rect 7295 36488 7531 36724
rect 7616 36488 7852 36724
rect 7937 36488 8173 36724
rect 8258 36488 8494 36724
rect 8579 36488 8815 36724
rect 8900 36488 9136 36724
rect 9221 36488 9457 36724
rect 9542 36488 9778 36724
rect 9863 36488 10099 36724
rect 10184 36488 10420 36724
rect 10505 36488 10741 36724
rect 10826 36488 11062 36724
rect 11147 36488 11383 36724
rect 11468 36488 11704 36724
rect 11789 36488 12025 36724
rect 12110 36488 12346 36724
rect 12431 36488 12667 36724
rect 12752 36488 12988 36724
rect 13073 36488 13309 36724
rect 13394 36488 13630 36724
rect 13715 36488 13951 36724
rect 14036 36488 14272 36724
rect 14357 36488 14593 36724
rect 14678 36488 14914 36724
rect 14999 36488 15235 36724
rect 15320 36488 15556 36724
rect 215 36164 451 36400
rect 537 36164 773 36400
rect 859 36164 1095 36400
rect 1181 36164 1417 36400
rect 1503 36164 1739 36400
rect 1825 36164 2061 36400
rect 2147 36164 2383 36400
rect 2469 36164 2705 36400
rect 2791 36164 3027 36400
rect 3113 36164 3349 36400
rect 3435 36164 3671 36400
rect 3757 36164 3993 36400
rect 4079 36164 4315 36400
rect 4401 36164 4637 36400
rect 4723 36164 4959 36400
rect 5045 36164 5281 36400
rect 5367 36164 5603 36400
rect 5689 36164 5925 36400
rect 6011 36164 6247 36400
rect 6332 36164 6568 36400
rect 6653 36164 6889 36400
rect 6974 36164 7210 36400
rect 7295 36164 7531 36400
rect 7616 36164 7852 36400
rect 7937 36164 8173 36400
rect 8258 36164 8494 36400
rect 8579 36164 8815 36400
rect 8900 36164 9136 36400
rect 9221 36164 9457 36400
rect 9542 36164 9778 36400
rect 9863 36164 10099 36400
rect 10184 36164 10420 36400
rect 10505 36164 10741 36400
rect 10826 36164 11062 36400
rect 11147 36164 11383 36400
rect 11468 36164 11704 36400
rect 11789 36164 12025 36400
rect 12110 36164 12346 36400
rect 12431 36164 12667 36400
rect 12752 36164 12988 36400
rect 13073 36164 13309 36400
rect 13394 36164 13630 36400
rect 13715 36164 13951 36400
rect 14036 36164 14272 36400
rect 14357 36164 14593 36400
rect 14678 36164 14914 36400
rect 14999 36164 15235 36400
rect 15320 36164 15556 36400
rect 215 35840 451 36076
rect 537 35840 773 36076
rect 859 35840 1095 36076
rect 1181 35840 1417 36076
rect 1503 35840 1739 36076
rect 1825 35840 2061 36076
rect 2147 35840 2383 36076
rect 2469 35840 2705 36076
rect 2791 35840 3027 36076
rect 3113 35840 3349 36076
rect 3435 35840 3671 36076
rect 3757 35840 3993 36076
rect 4079 35840 4315 36076
rect 4401 35840 4637 36076
rect 4723 35840 4959 36076
rect 5045 35840 5281 36076
rect 5367 35840 5603 36076
rect 5689 35840 5925 36076
rect 6011 35840 6247 36076
rect 6332 35840 6568 36076
rect 6653 35840 6889 36076
rect 6974 35840 7210 36076
rect 7295 35840 7531 36076
rect 7616 35840 7852 36076
rect 7937 35840 8173 36076
rect 8258 35840 8494 36076
rect 8579 35840 8815 36076
rect 8900 35840 9136 36076
rect 9221 35840 9457 36076
rect 9542 35840 9778 36076
rect 9863 35840 10099 36076
rect 10184 35840 10420 36076
rect 10505 35840 10741 36076
rect 10826 35840 11062 36076
rect 11147 35840 11383 36076
rect 11468 35840 11704 36076
rect 11789 35840 12025 36076
rect 12110 35840 12346 36076
rect 12431 35840 12667 36076
rect 12752 35840 12988 36076
rect 13073 35840 13309 36076
rect 13394 35840 13630 36076
rect 13715 35840 13951 36076
rect 14036 35840 14272 36076
rect 14357 35840 14593 36076
rect 14678 35840 14914 36076
rect 14999 35840 15235 36076
rect 15320 35840 15556 36076
rect 215 35516 451 35752
rect 537 35516 773 35752
rect 859 35516 1095 35752
rect 1181 35516 1417 35752
rect 1503 35516 1739 35752
rect 1825 35516 2061 35752
rect 2147 35516 2383 35752
rect 2469 35516 2705 35752
rect 2791 35516 3027 35752
rect 3113 35516 3349 35752
rect 3435 35516 3671 35752
rect 3757 35516 3993 35752
rect 4079 35516 4315 35752
rect 4401 35516 4637 35752
rect 4723 35516 4959 35752
rect 5045 35516 5281 35752
rect 5367 35516 5603 35752
rect 5689 35516 5925 35752
rect 6011 35516 6247 35752
rect 6332 35516 6568 35752
rect 6653 35516 6889 35752
rect 6974 35516 7210 35752
rect 7295 35516 7531 35752
rect 7616 35516 7852 35752
rect 7937 35516 8173 35752
rect 8258 35516 8494 35752
rect 8579 35516 8815 35752
rect 8900 35516 9136 35752
rect 9221 35516 9457 35752
rect 9542 35516 9778 35752
rect 9863 35516 10099 35752
rect 10184 35516 10420 35752
rect 10505 35516 10741 35752
rect 10826 35516 11062 35752
rect 11147 35516 11383 35752
rect 11468 35516 11704 35752
rect 11789 35516 12025 35752
rect 12110 35516 12346 35752
rect 12431 35516 12667 35752
rect 12752 35516 12988 35752
rect 13073 35516 13309 35752
rect 13394 35516 13630 35752
rect 13715 35516 13951 35752
rect 14036 35516 14272 35752
rect 14357 35516 14593 35752
rect 14678 35516 14914 35752
rect 14999 35516 15235 35752
rect 15320 35516 15556 35752
rect 215 35192 451 35428
rect 537 35192 773 35428
rect 859 35192 1095 35428
rect 1181 35192 1417 35428
rect 1503 35192 1739 35428
rect 1825 35192 2061 35428
rect 2147 35192 2383 35428
rect 2469 35192 2705 35428
rect 2791 35192 3027 35428
rect 3113 35192 3349 35428
rect 3435 35192 3671 35428
rect 3757 35192 3993 35428
rect 4079 35192 4315 35428
rect 4401 35192 4637 35428
rect 4723 35192 4959 35428
rect 5045 35192 5281 35428
rect 5367 35192 5603 35428
rect 5689 35192 5925 35428
rect 6011 35192 6247 35428
rect 6332 35192 6568 35428
rect 6653 35192 6889 35428
rect 6974 35192 7210 35428
rect 7295 35192 7531 35428
rect 7616 35192 7852 35428
rect 7937 35192 8173 35428
rect 8258 35192 8494 35428
rect 8579 35192 8815 35428
rect 8900 35192 9136 35428
rect 9221 35192 9457 35428
rect 9542 35192 9778 35428
rect 9863 35192 10099 35428
rect 10184 35192 10420 35428
rect 10505 35192 10741 35428
rect 10826 35192 11062 35428
rect 11147 35192 11383 35428
rect 11468 35192 11704 35428
rect 11789 35192 12025 35428
rect 12110 35192 12346 35428
rect 12431 35192 12667 35428
rect 12752 35192 12988 35428
rect 13073 35192 13309 35428
rect 13394 35192 13630 35428
rect 13715 35192 13951 35428
rect 14036 35192 14272 35428
rect 14357 35192 14593 35428
rect 14678 35192 14914 35428
rect 14999 35192 15235 35428
rect 15320 35192 15556 35428
rect 215 18736 451 18972
rect 538 18736 774 18972
rect 861 18736 1097 18972
rect 1184 18736 1420 18972
rect 1507 18736 1743 18972
rect 1830 18736 2066 18972
rect 2153 18736 2389 18972
rect 2476 18736 2712 18972
rect 2799 18736 3035 18972
rect 3122 18736 3358 18972
rect 3445 18736 3681 18972
rect 3768 18736 4004 18972
rect 4091 18736 4327 18972
rect 4414 18736 4650 18972
rect 4737 18736 4973 18972
rect 5060 18736 5296 18972
rect 5383 18736 5619 18972
rect 5706 18736 5942 18972
rect 6029 18736 6265 18972
rect 6351 18736 6587 18972
rect 6673 18736 6909 18972
rect 6995 18736 7231 18972
rect 7317 18736 7553 18972
rect 7639 18736 7875 18972
rect 7961 18736 8197 18972
rect 8283 18736 8519 18972
rect 8605 18736 8841 18972
rect 8927 18736 9163 18972
rect 9249 18736 9485 18972
rect 9571 18736 9807 18972
rect 9893 18736 10129 18972
rect 10215 18736 10451 18972
rect 10537 18736 10773 18972
rect 10859 18736 11095 18972
rect 11181 18736 11417 18972
rect 11503 18736 11739 18972
rect 11825 18736 12061 18972
rect 12147 18736 12383 18972
rect 12469 18736 12705 18972
rect 12791 18736 13027 18972
rect 13113 18736 13349 18972
rect 13435 18736 13671 18972
rect 13757 18736 13993 18972
rect 14079 18736 14315 18972
rect 14401 18736 14637 18972
rect 14723 18736 14959 18972
rect 15045 18736 15281 18972
rect 15367 18736 15603 18972
rect 215 18400 451 18636
rect 538 18400 774 18636
rect 861 18400 1097 18636
rect 1184 18400 1420 18636
rect 1507 18400 1743 18636
rect 1830 18400 2066 18636
rect 2153 18400 2389 18636
rect 2476 18400 2712 18636
rect 2799 18400 3035 18636
rect 3122 18400 3358 18636
rect 3445 18400 3681 18636
rect 3768 18400 4004 18636
rect 4091 18400 4327 18636
rect 4414 18400 4650 18636
rect 4737 18400 4973 18636
rect 5060 18400 5296 18636
rect 5383 18400 5619 18636
rect 5706 18400 5942 18636
rect 6029 18400 6265 18636
rect 6351 18400 6587 18636
rect 6673 18400 6909 18636
rect 6995 18400 7231 18636
rect 7317 18400 7553 18636
rect 7639 18400 7875 18636
rect 7961 18400 8197 18636
rect 8283 18400 8519 18636
rect 8605 18400 8841 18636
rect 8927 18400 9163 18636
rect 9249 18400 9485 18636
rect 9571 18400 9807 18636
rect 9893 18400 10129 18636
rect 10215 18400 10451 18636
rect 10537 18400 10773 18636
rect 10859 18400 11095 18636
rect 11181 18400 11417 18636
rect 11503 18400 11739 18636
rect 11825 18400 12061 18636
rect 12147 18400 12383 18636
rect 12469 18400 12705 18636
rect 12791 18400 13027 18636
rect 13113 18400 13349 18636
rect 13435 18400 13671 18636
rect 13757 18400 13993 18636
rect 14079 18400 14315 18636
rect 14401 18400 14637 18636
rect 14723 18400 14959 18636
rect 15045 18400 15281 18636
rect 15367 18400 15603 18636
rect 215 18064 451 18300
rect 538 18064 774 18300
rect 861 18064 1097 18300
rect 1184 18064 1420 18300
rect 1507 18064 1743 18300
rect 1830 18064 2066 18300
rect 2153 18064 2389 18300
rect 2476 18064 2712 18300
rect 2799 18064 3035 18300
rect 3122 18064 3358 18300
rect 3445 18064 3681 18300
rect 3768 18064 4004 18300
rect 4091 18064 4327 18300
rect 4414 18064 4650 18300
rect 4737 18064 4973 18300
rect 5060 18064 5296 18300
rect 5383 18064 5619 18300
rect 5706 18064 5942 18300
rect 6029 18064 6265 18300
rect 6351 18064 6587 18300
rect 6673 18064 6909 18300
rect 6995 18064 7231 18300
rect 7317 18064 7553 18300
rect 7639 18064 7875 18300
rect 7961 18064 8197 18300
rect 8283 18064 8519 18300
rect 8605 18064 8841 18300
rect 8927 18064 9163 18300
rect 9249 18064 9485 18300
rect 9571 18064 9807 18300
rect 9893 18064 10129 18300
rect 10215 18064 10451 18300
rect 10537 18064 10773 18300
rect 10859 18064 11095 18300
rect 11181 18064 11417 18300
rect 11503 18064 11739 18300
rect 11825 18064 12061 18300
rect 12147 18064 12383 18300
rect 12469 18064 12705 18300
rect 12791 18064 13027 18300
rect 13113 18064 13349 18300
rect 13435 18064 13671 18300
rect 13757 18064 13993 18300
rect 14079 18064 14315 18300
rect 14401 18064 14637 18300
rect 14723 18064 14959 18300
rect 15045 18064 15281 18300
rect 15367 18064 15603 18300
rect 215 17728 451 17964
rect 538 17728 774 17964
rect 861 17728 1097 17964
rect 1184 17728 1420 17964
rect 1507 17728 1743 17964
rect 1830 17728 2066 17964
rect 2153 17728 2389 17964
rect 2476 17728 2712 17964
rect 2799 17728 3035 17964
rect 3122 17728 3358 17964
rect 3445 17728 3681 17964
rect 3768 17728 4004 17964
rect 4091 17728 4327 17964
rect 4414 17728 4650 17964
rect 4737 17728 4973 17964
rect 5060 17728 5296 17964
rect 5383 17728 5619 17964
rect 5706 17728 5942 17964
rect 6029 17728 6265 17964
rect 6351 17728 6587 17964
rect 6673 17728 6909 17964
rect 6995 17728 7231 17964
rect 7317 17728 7553 17964
rect 7639 17728 7875 17964
rect 7961 17728 8197 17964
rect 8283 17728 8519 17964
rect 8605 17728 8841 17964
rect 8927 17728 9163 17964
rect 9249 17728 9485 17964
rect 9571 17728 9807 17964
rect 9893 17728 10129 17964
rect 10215 17728 10451 17964
rect 10537 17728 10773 17964
rect 10859 17728 11095 17964
rect 11181 17728 11417 17964
rect 11503 17728 11739 17964
rect 11825 17728 12061 17964
rect 12147 17728 12383 17964
rect 12469 17728 12705 17964
rect 12791 17728 13027 17964
rect 13113 17728 13349 17964
rect 13435 17728 13671 17964
rect 13757 17728 13993 17964
rect 14079 17728 14315 17964
rect 14401 17728 14637 17964
rect 14723 17728 14959 17964
rect 15045 17728 15281 17964
rect 15367 17728 15603 17964
rect 215 17392 451 17628
rect 538 17392 774 17628
rect 861 17392 1097 17628
rect 1184 17392 1420 17628
rect 1507 17392 1743 17628
rect 1830 17392 2066 17628
rect 2153 17392 2389 17628
rect 2476 17392 2712 17628
rect 2799 17392 3035 17628
rect 3122 17392 3358 17628
rect 3445 17392 3681 17628
rect 3768 17392 4004 17628
rect 4091 17392 4327 17628
rect 4414 17392 4650 17628
rect 4737 17392 4973 17628
rect 5060 17392 5296 17628
rect 5383 17392 5619 17628
rect 5706 17392 5942 17628
rect 6029 17392 6265 17628
rect 6351 17392 6587 17628
rect 6673 17392 6909 17628
rect 6995 17392 7231 17628
rect 7317 17392 7553 17628
rect 7639 17392 7875 17628
rect 7961 17392 8197 17628
rect 8283 17392 8519 17628
rect 8605 17392 8841 17628
rect 8927 17392 9163 17628
rect 9249 17392 9485 17628
rect 9571 17392 9807 17628
rect 9893 17392 10129 17628
rect 10215 17392 10451 17628
rect 10537 17392 10773 17628
rect 10859 17392 11095 17628
rect 11181 17392 11417 17628
rect 11503 17392 11739 17628
rect 11825 17392 12061 17628
rect 12147 17392 12383 17628
rect 12469 17392 12705 17628
rect 12791 17392 13027 17628
rect 13113 17392 13349 17628
rect 13435 17392 13671 17628
rect 13757 17392 13993 17628
rect 14079 17392 14315 17628
rect 14401 17392 14637 17628
rect 14723 17392 14959 17628
rect 15045 17392 15281 17628
rect 15367 17392 15603 17628
rect 215 17056 451 17292
rect 538 17056 774 17292
rect 861 17056 1097 17292
rect 1184 17056 1420 17292
rect 1507 17056 1743 17292
rect 1830 17056 2066 17292
rect 2153 17056 2389 17292
rect 2476 17056 2712 17292
rect 2799 17056 3035 17292
rect 3122 17056 3358 17292
rect 3445 17056 3681 17292
rect 3768 17056 4004 17292
rect 4091 17056 4327 17292
rect 4414 17056 4650 17292
rect 4737 17056 4973 17292
rect 5060 17056 5296 17292
rect 5383 17056 5619 17292
rect 5706 17056 5942 17292
rect 6029 17056 6265 17292
rect 6351 17056 6587 17292
rect 6673 17056 6909 17292
rect 6995 17056 7231 17292
rect 7317 17056 7553 17292
rect 7639 17056 7875 17292
rect 7961 17056 8197 17292
rect 8283 17056 8519 17292
rect 8605 17056 8841 17292
rect 8927 17056 9163 17292
rect 9249 17056 9485 17292
rect 9571 17056 9807 17292
rect 9893 17056 10129 17292
rect 10215 17056 10451 17292
rect 10537 17056 10773 17292
rect 10859 17056 11095 17292
rect 11181 17056 11417 17292
rect 11503 17056 11739 17292
rect 11825 17056 12061 17292
rect 12147 17056 12383 17292
rect 12469 17056 12705 17292
rect 12791 17056 13027 17292
rect 13113 17056 13349 17292
rect 13435 17056 13671 17292
rect 13757 17056 13993 17292
rect 14079 17056 14315 17292
rect 14401 17056 14637 17292
rect 14723 17056 14959 17292
rect 15045 17056 15281 17292
rect 15367 17056 15603 17292
rect 215 16720 451 16956
rect 538 16720 774 16956
rect 861 16720 1097 16956
rect 1184 16720 1420 16956
rect 1507 16720 1743 16956
rect 1830 16720 2066 16956
rect 2153 16720 2389 16956
rect 2476 16720 2712 16956
rect 2799 16720 3035 16956
rect 3122 16720 3358 16956
rect 3445 16720 3681 16956
rect 3768 16720 4004 16956
rect 4091 16720 4327 16956
rect 4414 16720 4650 16956
rect 4737 16720 4973 16956
rect 5060 16720 5296 16956
rect 5383 16720 5619 16956
rect 5706 16720 5942 16956
rect 6029 16720 6265 16956
rect 6351 16720 6587 16956
rect 6673 16720 6909 16956
rect 6995 16720 7231 16956
rect 7317 16720 7553 16956
rect 7639 16720 7875 16956
rect 7961 16720 8197 16956
rect 8283 16720 8519 16956
rect 8605 16720 8841 16956
rect 8927 16720 9163 16956
rect 9249 16720 9485 16956
rect 9571 16720 9807 16956
rect 9893 16720 10129 16956
rect 10215 16720 10451 16956
rect 10537 16720 10773 16956
rect 10859 16720 11095 16956
rect 11181 16720 11417 16956
rect 11503 16720 11739 16956
rect 11825 16720 12061 16956
rect 12147 16720 12383 16956
rect 12469 16720 12705 16956
rect 12791 16720 13027 16956
rect 13113 16720 13349 16956
rect 13435 16720 13671 16956
rect 13757 16720 13993 16956
rect 14079 16720 14315 16956
rect 14401 16720 14637 16956
rect 14723 16720 14959 16956
rect 15045 16720 15281 16956
rect 15367 16720 15603 16956
rect 215 16384 451 16620
rect 538 16384 774 16620
rect 861 16384 1097 16620
rect 1184 16384 1420 16620
rect 1507 16384 1743 16620
rect 1830 16384 2066 16620
rect 2153 16384 2389 16620
rect 2476 16384 2712 16620
rect 2799 16384 3035 16620
rect 3122 16384 3358 16620
rect 3445 16384 3681 16620
rect 3768 16384 4004 16620
rect 4091 16384 4327 16620
rect 4414 16384 4650 16620
rect 4737 16384 4973 16620
rect 5060 16384 5296 16620
rect 5383 16384 5619 16620
rect 5706 16384 5942 16620
rect 6029 16384 6265 16620
rect 6351 16384 6587 16620
rect 6673 16384 6909 16620
rect 6995 16384 7231 16620
rect 7317 16384 7553 16620
rect 7639 16384 7875 16620
rect 7961 16384 8197 16620
rect 8283 16384 8519 16620
rect 8605 16384 8841 16620
rect 8927 16384 9163 16620
rect 9249 16384 9485 16620
rect 9571 16384 9807 16620
rect 9893 16384 10129 16620
rect 10215 16384 10451 16620
rect 10537 16384 10773 16620
rect 10859 16384 11095 16620
rect 11181 16384 11417 16620
rect 11503 16384 11739 16620
rect 11825 16384 12061 16620
rect 12147 16384 12383 16620
rect 12469 16384 12705 16620
rect 12791 16384 13027 16620
rect 13113 16384 13349 16620
rect 13435 16384 13671 16620
rect 13757 16384 13993 16620
rect 14079 16384 14315 16620
rect 14401 16384 14637 16620
rect 14723 16384 14959 16620
rect 15045 16384 15281 16620
rect 15367 16384 15603 16620
rect 215 16048 451 16284
rect 538 16048 774 16284
rect 861 16048 1097 16284
rect 1184 16048 1420 16284
rect 1507 16048 1743 16284
rect 1830 16048 2066 16284
rect 2153 16048 2389 16284
rect 2476 16048 2712 16284
rect 2799 16048 3035 16284
rect 3122 16048 3358 16284
rect 3445 16048 3681 16284
rect 3768 16048 4004 16284
rect 4091 16048 4327 16284
rect 4414 16048 4650 16284
rect 4737 16048 4973 16284
rect 5060 16048 5296 16284
rect 5383 16048 5619 16284
rect 5706 16048 5942 16284
rect 6029 16048 6265 16284
rect 6351 16048 6587 16284
rect 6673 16048 6909 16284
rect 6995 16048 7231 16284
rect 7317 16048 7553 16284
rect 7639 16048 7875 16284
rect 7961 16048 8197 16284
rect 8283 16048 8519 16284
rect 8605 16048 8841 16284
rect 8927 16048 9163 16284
rect 9249 16048 9485 16284
rect 9571 16048 9807 16284
rect 9893 16048 10129 16284
rect 10215 16048 10451 16284
rect 10537 16048 10773 16284
rect 10859 16048 11095 16284
rect 11181 16048 11417 16284
rect 11503 16048 11739 16284
rect 11825 16048 12061 16284
rect 12147 16048 12383 16284
rect 12469 16048 12705 16284
rect 12791 16048 13027 16284
rect 13113 16048 13349 16284
rect 13435 16048 13671 16284
rect 13757 16048 13993 16284
rect 14079 16048 14315 16284
rect 14401 16048 14637 16284
rect 14723 16048 14959 16284
rect 15045 16048 15281 16284
rect 15367 16048 15603 16284
rect 215 15712 451 15948
rect 538 15712 774 15948
rect 861 15712 1097 15948
rect 1184 15712 1420 15948
rect 1507 15712 1743 15948
rect 1830 15712 2066 15948
rect 2153 15712 2389 15948
rect 2476 15712 2712 15948
rect 2799 15712 3035 15948
rect 3122 15712 3358 15948
rect 3445 15712 3681 15948
rect 3768 15712 4004 15948
rect 4091 15712 4327 15948
rect 4414 15712 4650 15948
rect 4737 15712 4973 15948
rect 5060 15712 5296 15948
rect 5383 15712 5619 15948
rect 5706 15712 5942 15948
rect 6029 15712 6265 15948
rect 6351 15712 6587 15948
rect 6673 15712 6909 15948
rect 6995 15712 7231 15948
rect 7317 15712 7553 15948
rect 7639 15712 7875 15948
rect 7961 15712 8197 15948
rect 8283 15712 8519 15948
rect 8605 15712 8841 15948
rect 8927 15712 9163 15948
rect 9249 15712 9485 15948
rect 9571 15712 9807 15948
rect 9893 15712 10129 15948
rect 10215 15712 10451 15948
rect 10537 15712 10773 15948
rect 10859 15712 11095 15948
rect 11181 15712 11417 15948
rect 11503 15712 11739 15948
rect 11825 15712 12061 15948
rect 12147 15712 12383 15948
rect 12469 15712 12705 15948
rect 12791 15712 13027 15948
rect 13113 15712 13349 15948
rect 13435 15712 13671 15948
rect 13757 15712 13993 15948
rect 14079 15712 14315 15948
rect 14401 15712 14637 15948
rect 14723 15712 14959 15948
rect 15045 15712 15281 15948
rect 15367 15712 15603 15948
rect 215 15376 451 15612
rect 538 15376 774 15612
rect 861 15376 1097 15612
rect 1184 15376 1420 15612
rect 1507 15376 1743 15612
rect 1830 15376 2066 15612
rect 2153 15376 2389 15612
rect 2476 15376 2712 15612
rect 2799 15376 3035 15612
rect 3122 15376 3358 15612
rect 3445 15376 3681 15612
rect 3768 15376 4004 15612
rect 4091 15376 4327 15612
rect 4414 15376 4650 15612
rect 4737 15376 4973 15612
rect 5060 15376 5296 15612
rect 5383 15376 5619 15612
rect 5706 15376 5942 15612
rect 6029 15376 6265 15612
rect 6351 15376 6587 15612
rect 6673 15376 6909 15612
rect 6995 15376 7231 15612
rect 7317 15376 7553 15612
rect 7639 15376 7875 15612
rect 7961 15376 8197 15612
rect 8283 15376 8519 15612
rect 8605 15376 8841 15612
rect 8927 15376 9163 15612
rect 9249 15376 9485 15612
rect 9571 15376 9807 15612
rect 9893 15376 10129 15612
rect 10215 15376 10451 15612
rect 10537 15376 10773 15612
rect 10859 15376 11095 15612
rect 11181 15376 11417 15612
rect 11503 15376 11739 15612
rect 11825 15376 12061 15612
rect 12147 15376 12383 15612
rect 12469 15376 12705 15612
rect 12791 15376 13027 15612
rect 13113 15376 13349 15612
rect 13435 15376 13671 15612
rect 13757 15376 13993 15612
rect 14079 15376 14315 15612
rect 14401 15376 14637 15612
rect 14723 15376 14959 15612
rect 15045 15376 15281 15612
rect 15367 15376 15603 15612
rect 215 15040 451 15276
rect 538 15040 774 15276
rect 861 15040 1097 15276
rect 1184 15040 1420 15276
rect 1507 15040 1743 15276
rect 1830 15040 2066 15276
rect 2153 15040 2389 15276
rect 2476 15040 2712 15276
rect 2799 15040 3035 15276
rect 3122 15040 3358 15276
rect 3445 15040 3681 15276
rect 3768 15040 4004 15276
rect 4091 15040 4327 15276
rect 4414 15040 4650 15276
rect 4737 15040 4973 15276
rect 5060 15040 5296 15276
rect 5383 15040 5619 15276
rect 5706 15040 5942 15276
rect 6029 15040 6265 15276
rect 6351 15040 6587 15276
rect 6673 15040 6909 15276
rect 6995 15040 7231 15276
rect 7317 15040 7553 15276
rect 7639 15040 7875 15276
rect 7961 15040 8197 15276
rect 8283 15040 8519 15276
rect 8605 15040 8841 15276
rect 8927 15040 9163 15276
rect 9249 15040 9485 15276
rect 9571 15040 9807 15276
rect 9893 15040 10129 15276
rect 10215 15040 10451 15276
rect 10537 15040 10773 15276
rect 10859 15040 11095 15276
rect 11181 15040 11417 15276
rect 11503 15040 11739 15276
rect 11825 15040 12061 15276
rect 12147 15040 12383 15276
rect 12469 15040 12705 15276
rect 12791 15040 13027 15276
rect 13113 15040 13349 15276
rect 13435 15040 13671 15276
rect 13757 15040 13993 15276
rect 14079 15040 14315 15276
rect 14401 15040 14637 15276
rect 14723 15040 14959 15276
rect 15045 15040 15281 15276
rect 15367 15040 15603 15276
rect 215 14704 451 14940
rect 538 14704 774 14940
rect 861 14704 1097 14940
rect 1184 14704 1420 14940
rect 1507 14704 1743 14940
rect 1830 14704 2066 14940
rect 2153 14704 2389 14940
rect 2476 14704 2712 14940
rect 2799 14704 3035 14940
rect 3122 14704 3358 14940
rect 3445 14704 3681 14940
rect 3768 14704 4004 14940
rect 4091 14704 4327 14940
rect 4414 14704 4650 14940
rect 4737 14704 4973 14940
rect 5060 14704 5296 14940
rect 5383 14704 5619 14940
rect 5706 14704 5942 14940
rect 6029 14704 6265 14940
rect 6351 14704 6587 14940
rect 6673 14704 6909 14940
rect 6995 14704 7231 14940
rect 7317 14704 7553 14940
rect 7639 14704 7875 14940
rect 7961 14704 8197 14940
rect 8283 14704 8519 14940
rect 8605 14704 8841 14940
rect 8927 14704 9163 14940
rect 9249 14704 9485 14940
rect 9571 14704 9807 14940
rect 9893 14704 10129 14940
rect 10215 14704 10451 14940
rect 10537 14704 10773 14940
rect 10859 14704 11095 14940
rect 11181 14704 11417 14940
rect 11503 14704 11739 14940
rect 11825 14704 12061 14940
rect 12147 14704 12383 14940
rect 12469 14704 12705 14940
rect 12791 14704 13027 14940
rect 13113 14704 13349 14940
rect 13435 14704 13671 14940
rect 13757 14704 13993 14940
rect 14079 14704 14315 14940
rect 14401 14704 14637 14940
rect 14723 14704 14959 14940
rect 15045 14704 15281 14940
rect 15367 14704 15603 14940
rect 215 14368 451 14604
rect 538 14368 774 14604
rect 861 14368 1097 14604
rect 1184 14368 1420 14604
rect 1507 14368 1743 14604
rect 1830 14368 2066 14604
rect 2153 14368 2389 14604
rect 2476 14368 2712 14604
rect 2799 14368 3035 14604
rect 3122 14368 3358 14604
rect 3445 14368 3681 14604
rect 3768 14368 4004 14604
rect 4091 14368 4327 14604
rect 4414 14368 4650 14604
rect 4737 14368 4973 14604
rect 5060 14368 5296 14604
rect 5383 14368 5619 14604
rect 5706 14368 5942 14604
rect 6029 14368 6265 14604
rect 6351 14368 6587 14604
rect 6673 14368 6909 14604
rect 6995 14368 7231 14604
rect 7317 14368 7553 14604
rect 7639 14368 7875 14604
rect 7961 14368 8197 14604
rect 8283 14368 8519 14604
rect 8605 14368 8841 14604
rect 8927 14368 9163 14604
rect 9249 14368 9485 14604
rect 9571 14368 9807 14604
rect 9893 14368 10129 14604
rect 10215 14368 10451 14604
rect 10537 14368 10773 14604
rect 10859 14368 11095 14604
rect 11181 14368 11417 14604
rect 11503 14368 11739 14604
rect 11825 14368 12061 14604
rect 12147 14368 12383 14604
rect 12469 14368 12705 14604
rect 12791 14368 13027 14604
rect 13113 14368 13349 14604
rect 13435 14368 13671 14604
rect 13757 14368 13993 14604
rect 14079 14368 14315 14604
rect 14401 14368 14637 14604
rect 14723 14368 14959 14604
rect 15045 14368 15281 14604
rect 15367 14368 15603 14604
rect 215 14032 451 14268
rect 538 14032 774 14268
rect 861 14032 1097 14268
rect 1184 14032 1420 14268
rect 1507 14032 1743 14268
rect 1830 14032 2066 14268
rect 2153 14032 2389 14268
rect 2476 14032 2712 14268
rect 2799 14032 3035 14268
rect 3122 14032 3358 14268
rect 3445 14032 3681 14268
rect 3768 14032 4004 14268
rect 4091 14032 4327 14268
rect 4414 14032 4650 14268
rect 4737 14032 4973 14268
rect 5060 14032 5296 14268
rect 5383 14032 5619 14268
rect 5706 14032 5942 14268
rect 6029 14032 6265 14268
rect 6351 14032 6587 14268
rect 6673 14032 6909 14268
rect 6995 14032 7231 14268
rect 7317 14032 7553 14268
rect 7639 14032 7875 14268
rect 7961 14032 8197 14268
rect 8283 14032 8519 14268
rect 8605 14032 8841 14268
rect 8927 14032 9163 14268
rect 9249 14032 9485 14268
rect 9571 14032 9807 14268
rect 9893 14032 10129 14268
rect 10215 14032 10451 14268
rect 10537 14032 10773 14268
rect 10859 14032 11095 14268
rect 11181 14032 11417 14268
rect 11503 14032 11739 14268
rect 11825 14032 12061 14268
rect 12147 14032 12383 14268
rect 12469 14032 12705 14268
rect 12791 14032 13027 14268
rect 13113 14032 13349 14268
rect 13435 14032 13671 14268
rect 13757 14032 13993 14268
rect 14079 14032 14315 14268
rect 14401 14032 14637 14268
rect 14723 14032 14959 14268
rect 15045 14032 15281 14268
rect 15367 14032 15603 14268
rect 216 13427 452 13663
rect 538 13427 774 13663
rect 860 13427 1096 13663
rect 1182 13427 1418 13663
rect 1504 13427 1740 13663
rect 1826 13427 2062 13663
rect 2148 13427 2384 13663
rect 2470 13427 2706 13663
rect 2792 13427 3028 13663
rect 3114 13427 3350 13663
rect 3436 13427 3672 13663
rect 3758 13427 3994 13663
rect 4080 13427 4316 13663
rect 4402 13427 4638 13663
rect 4724 13427 4960 13663
rect 5046 13427 5282 13663
rect 5368 13427 5604 13663
rect 5690 13427 5926 13663
rect 6012 13427 6248 13663
rect 6333 13427 6569 13663
rect 6654 13427 6890 13663
rect 6975 13427 7211 13663
rect 7296 13427 7532 13663
rect 7617 13427 7853 13663
rect 7938 13427 8174 13663
rect 8259 13637 8333 13663
rect 8333 13637 8397 13663
rect 8397 13637 8417 13663
rect 8417 13637 8481 13663
rect 8481 13637 8495 13663
rect 8580 13637 8585 13663
rect 8585 13637 8649 13663
rect 8649 13637 8669 13663
rect 8669 13637 8733 13663
rect 8733 13637 8816 13663
rect 8259 13620 8495 13637
rect 8580 13620 8816 13637
rect 8259 13556 8333 13620
rect 8333 13556 8397 13620
rect 8397 13556 8417 13620
rect 8417 13556 8481 13620
rect 8481 13556 8495 13620
rect 8580 13556 8585 13620
rect 8585 13556 8649 13620
rect 8649 13556 8669 13620
rect 8669 13556 8733 13620
rect 8733 13556 8816 13620
rect 8259 13539 8495 13556
rect 8580 13539 8816 13556
rect 8259 13475 8333 13539
rect 8333 13475 8397 13539
rect 8397 13475 8417 13539
rect 8417 13475 8481 13539
rect 8481 13475 8495 13539
rect 8580 13475 8585 13539
rect 8585 13475 8649 13539
rect 8649 13475 8669 13539
rect 8669 13475 8733 13539
rect 8733 13475 8816 13539
rect 8259 13458 8495 13475
rect 8580 13458 8816 13475
rect 8259 13427 8333 13458
rect 8333 13427 8397 13458
rect 8397 13427 8417 13458
rect 8417 13427 8481 13458
rect 8481 13427 8495 13458
rect 8580 13427 8585 13458
rect 8585 13427 8649 13458
rect 8649 13427 8669 13458
rect 8669 13427 8733 13458
rect 8733 13427 8816 13458
rect 8901 13427 9137 13663
rect 9222 13427 9458 13663
rect 9543 13427 9779 13663
rect 9864 13427 10100 13663
rect 10185 13427 10421 13663
rect 10506 13427 10742 13663
rect 10827 13427 11063 13663
rect 11148 13427 11384 13663
rect 11469 13427 11705 13663
rect 11790 13427 12026 13663
rect 12111 13427 12347 13663
rect 12432 13427 12668 13663
rect 12753 13427 12989 13663
rect 13074 13427 13310 13663
rect 13395 13427 13631 13663
rect 13716 13427 13952 13663
rect 14037 13427 14273 13663
rect 14358 13427 14594 13663
rect 14679 13427 14915 13663
rect 15000 13427 15236 13663
rect 15321 13427 15557 13663
rect 216 12861 452 13097
rect 538 12861 774 13097
rect 860 12861 1096 13097
rect 1182 12861 1418 13097
rect 1504 12861 1740 13097
rect 1826 12861 2062 13097
rect 2148 12861 2384 13097
rect 2470 12861 2706 13097
rect 2792 12861 3028 13097
rect 3114 12861 3350 13097
rect 3436 12861 3672 13097
rect 3758 12861 3994 13097
rect 4080 12861 4316 13097
rect 4402 12861 4638 13097
rect 4724 12861 4960 13097
rect 5046 12861 5282 13097
rect 5368 12861 5604 13097
rect 5690 12861 5926 13097
rect 6012 12861 6248 13097
rect 6333 12861 6569 13097
rect 6654 12861 6890 13097
rect 6975 12861 7211 13097
rect 7296 12861 7532 13097
rect 7617 12861 7853 13097
rect 7938 12861 8174 13097
rect 8259 13069 8333 13097
rect 8333 13069 8397 13097
rect 8397 13069 8417 13097
rect 8417 13069 8481 13097
rect 8481 13069 8495 13097
rect 8580 13069 8585 13097
rect 8585 13069 8649 13097
rect 8649 13069 8669 13097
rect 8669 13069 8733 13097
rect 8733 13069 8816 13097
rect 8259 13051 8495 13069
rect 8580 13051 8816 13069
rect 8259 12987 8333 13051
rect 8333 12987 8397 13051
rect 8397 12987 8417 13051
rect 8417 12987 8481 13051
rect 8481 12987 8495 13051
rect 8580 12987 8585 13051
rect 8585 12987 8649 13051
rect 8649 12987 8669 13051
rect 8669 12987 8733 13051
rect 8733 12987 8816 13051
rect 8259 12969 8495 12987
rect 8580 12969 8816 12987
rect 8259 12905 8333 12969
rect 8333 12905 8397 12969
rect 8397 12905 8417 12969
rect 8417 12905 8481 12969
rect 8481 12905 8495 12969
rect 8580 12905 8585 12969
rect 8585 12905 8649 12969
rect 8649 12905 8669 12969
rect 8669 12905 8733 12969
rect 8733 12905 8816 12969
rect 8259 12887 8495 12905
rect 8580 12887 8816 12905
rect 8259 12861 8333 12887
rect 8333 12861 8397 12887
rect 8397 12861 8417 12887
rect 8417 12861 8481 12887
rect 8481 12861 8495 12887
rect 8580 12861 8585 12887
rect 8585 12861 8649 12887
rect 8649 12861 8669 12887
rect 8669 12861 8733 12887
rect 8733 12861 8816 12887
rect 8901 12861 9137 13097
rect 9222 12861 9458 13097
rect 9543 12861 9779 13097
rect 9864 12861 10100 13097
rect 10185 12861 10421 13097
rect 10506 12861 10742 13097
rect 10827 12861 11063 13097
rect 11148 12861 11384 13097
rect 11469 12861 11705 13097
rect 11790 12861 12026 13097
rect 12111 12861 12347 13097
rect 12432 12861 12668 13097
rect 12753 12861 12989 13097
rect 13074 12861 13310 13097
rect 13395 12861 13631 13097
rect 13716 12861 13952 13097
rect 14037 12861 14273 13097
rect 14358 12861 14594 13097
rect 14679 12861 14915 13097
rect 15000 12861 15236 13097
rect 15321 12861 15557 13097
rect 215 12257 451 12493
rect 537 12257 773 12493
rect 859 12257 1095 12493
rect 1181 12257 1417 12493
rect 1503 12257 1739 12493
rect 1825 12257 2061 12493
rect 2147 12257 2383 12493
rect 2469 12257 2705 12493
rect 2791 12257 3027 12493
rect 3113 12257 3349 12493
rect 3435 12257 3671 12493
rect 3757 12257 3993 12493
rect 4079 12257 4315 12493
rect 4401 12257 4637 12493
rect 4723 12257 4959 12493
rect 5045 12257 5281 12493
rect 5367 12257 5603 12493
rect 5689 12257 5925 12493
rect 6011 12257 6247 12493
rect 6332 12257 6568 12493
rect 6653 12257 6889 12493
rect 6974 12257 7210 12493
rect 7295 12257 7531 12493
rect 7616 12257 7852 12493
rect 7937 12257 8173 12493
rect 8258 12257 8494 12493
rect 8579 12257 8815 12493
rect 8900 12257 9136 12493
rect 9221 12257 9457 12493
rect 9542 12257 9778 12493
rect 9863 12257 10099 12493
rect 10184 12257 10420 12493
rect 10505 12257 10741 12493
rect 10826 12257 11062 12493
rect 11147 12257 11383 12493
rect 11468 12257 11704 12493
rect 11789 12257 12025 12493
rect 12110 12257 12346 12493
rect 12431 12257 12667 12493
rect 12752 12257 12988 12493
rect 13073 12257 13309 12493
rect 13394 12257 13630 12493
rect 13715 12257 13951 12493
rect 14036 12257 14272 12493
rect 14357 12257 14593 12493
rect 14678 12257 14914 12493
rect 14999 12257 15235 12493
rect 15320 12257 15556 12493
rect 215 11691 451 11927
rect 537 11691 773 11927
rect 859 11691 1095 11927
rect 1181 11691 1417 11927
rect 1503 11691 1739 11927
rect 1825 11691 2061 11927
rect 2147 11691 2383 11927
rect 2469 11691 2705 11927
rect 2791 11691 3027 11927
rect 3113 11691 3349 11927
rect 3435 11691 3671 11927
rect 3757 11691 3993 11927
rect 4079 11691 4315 11927
rect 4401 11691 4637 11927
rect 4723 11691 4959 11927
rect 5045 11691 5281 11927
rect 5367 11691 5603 11927
rect 5689 11691 5925 11927
rect 6011 11691 6247 11927
rect 6332 11691 6568 11927
rect 6653 11691 6889 11927
rect 6974 11691 7210 11927
rect 7295 11691 7531 11927
rect 7616 11691 7852 11927
rect 7937 11691 8173 11927
rect 8258 11691 8494 11927
rect 8579 11691 8815 11927
rect 8900 11691 9136 11927
rect 9221 11691 9457 11927
rect 9542 11691 9778 11927
rect 9863 11691 10099 11927
rect 10184 11691 10420 11927
rect 10505 11691 10741 11927
rect 10826 11691 11062 11927
rect 11147 11691 11383 11927
rect 11468 11691 11704 11927
rect 11789 11691 12025 11927
rect 12110 11691 12346 11927
rect 12431 11691 12667 11927
rect 12752 11691 12988 11927
rect 13073 11691 13309 11927
rect 13394 11691 13630 11927
rect 13715 11691 13951 11927
rect 14036 11691 14272 11927
rect 14357 11691 14593 11927
rect 14678 11691 14914 11927
rect 14999 11691 15235 11927
rect 15320 11691 15556 11927
rect 215 10329 451 10565
rect 537 10329 773 10565
rect 859 10329 1095 10565
rect 1181 10329 1417 10565
rect 1503 10329 1739 10565
rect 1825 10329 2061 10565
rect 2147 10329 2383 10565
rect 2469 10329 2705 10565
rect 2791 10329 3027 10565
rect 3113 10329 3349 10565
rect 3435 10329 3671 10565
rect 3757 10329 3993 10565
rect 4079 10329 4315 10565
rect 4401 10329 4637 10565
rect 4723 10329 4959 10565
rect 5045 10329 5281 10565
rect 5367 10329 5603 10565
rect 5689 10329 5925 10565
rect 6011 10329 6247 10565
rect 6332 10329 6568 10565
rect 6653 10329 6889 10565
rect 6974 10329 7210 10565
rect 7295 10329 7531 10565
rect 7616 10329 7852 10565
rect 7937 10329 8173 10565
rect 8258 10329 8494 10565
rect 8579 10329 8815 10565
rect 8900 10329 9136 10565
rect 9221 10329 9457 10565
rect 9542 10329 9778 10565
rect 9863 10329 10099 10565
rect 10184 10329 10420 10565
rect 10505 10329 10741 10565
rect 10826 10329 11062 10565
rect 11147 10329 11383 10565
rect 11468 10329 11704 10565
rect 11789 10329 12025 10565
rect 12110 10329 12346 10565
rect 12431 10329 12667 10565
rect 12752 10329 12988 10565
rect 13073 10329 13309 10565
rect 13394 10329 13630 10565
rect 13715 10329 13951 10565
rect 14036 10329 14272 10565
rect 14357 10329 14593 10565
rect 14678 10329 14914 10565
rect 14999 10329 15235 10565
rect 15320 10329 15556 10565
rect 216 9180 397 9203
rect 397 9180 452 9203
rect 538 9180 543 9203
rect 543 9180 561 9203
rect 561 9180 625 9203
rect 625 9180 643 9203
rect 643 9180 707 9203
rect 707 9180 725 9203
rect 725 9180 774 9203
rect 860 9180 871 9203
rect 871 9180 889 9203
rect 889 9180 953 9203
rect 953 9180 971 9203
rect 971 9180 1035 9203
rect 1035 9180 1053 9203
rect 1053 9180 1096 9203
rect 1182 9180 1199 9203
rect 1199 9180 1217 9203
rect 1217 9180 1281 9203
rect 1281 9180 1299 9203
rect 1299 9180 1363 9203
rect 1363 9180 1381 9203
rect 1381 9180 1418 9203
rect 1504 9180 1527 9203
rect 1527 9180 1545 9203
rect 1545 9180 1609 9203
rect 1609 9180 1627 9203
rect 1627 9180 1691 9203
rect 1691 9180 1709 9203
rect 1709 9180 1740 9203
rect 1826 9180 1855 9203
rect 1855 9180 1873 9203
rect 1873 9180 1937 9203
rect 1937 9180 1955 9203
rect 1955 9180 2019 9203
rect 2019 9180 2037 9203
rect 2037 9180 2062 9203
rect 2148 9180 2183 9203
rect 2183 9180 2201 9203
rect 2201 9180 2265 9203
rect 2265 9180 2282 9203
rect 2282 9180 2346 9203
rect 2346 9180 2363 9203
rect 2363 9180 2384 9203
rect 2470 9180 2553 9203
rect 2553 9180 2617 9203
rect 2617 9180 2635 9203
rect 2635 9180 2699 9203
rect 2699 9180 2706 9203
rect 2792 9180 2799 9203
rect 2799 9180 2863 9203
rect 2863 9180 2881 9203
rect 2881 9180 2945 9203
rect 2945 9180 2963 9203
rect 2963 9180 3027 9203
rect 3027 9180 3028 9203
rect 3114 9180 3127 9203
rect 3127 9180 3191 9203
rect 3191 9180 3209 9203
rect 3209 9180 3273 9203
rect 3273 9180 3290 9203
rect 3290 9180 3350 9203
rect 3436 9180 3452 9203
rect 3452 9180 3516 9203
rect 3516 9180 3533 9203
rect 3533 9180 3597 9203
rect 3597 9180 3614 9203
rect 3614 9180 3672 9203
rect 3758 9180 3759 9203
rect 3759 9180 3776 9203
rect 3776 9180 3840 9203
rect 3840 9180 3857 9203
rect 3857 9180 3921 9203
rect 3921 9180 3938 9203
rect 3938 9180 3994 9203
rect 4080 9180 4083 9203
rect 4083 9180 4100 9203
rect 4100 9180 4164 9203
rect 4164 9180 4181 9203
rect 4181 9180 4245 9203
rect 4245 9180 4262 9203
rect 4262 9180 4316 9203
rect 4402 9180 4407 9203
rect 4407 9180 4424 9203
rect 4424 9180 4488 9203
rect 4488 9180 4505 9203
rect 4505 9180 4569 9203
rect 4569 9180 4638 9203
rect 4724 9180 4759 9203
rect 4759 9180 4777 9203
rect 4777 9180 4841 9203
rect 4841 9180 4859 9203
rect 4859 9180 4923 9203
rect 4923 9180 4941 9203
rect 4941 9180 4960 9203
rect 5046 9180 5087 9203
rect 5087 9180 5105 9203
rect 5105 9180 5169 9203
rect 5169 9180 5187 9203
rect 5187 9180 5251 9203
rect 5251 9180 5269 9203
rect 5269 9180 5282 9203
rect 5368 9180 5415 9203
rect 5415 9180 5433 9203
rect 5433 9180 5497 9203
rect 5497 9180 5515 9203
rect 5515 9180 5579 9203
rect 5579 9180 5597 9203
rect 5597 9180 5604 9203
rect 5690 9180 5743 9203
rect 5743 9180 5760 9203
rect 5760 9180 5824 9203
rect 5824 9180 5841 9203
rect 5841 9180 5905 9203
rect 5905 9180 5922 9203
rect 5922 9180 5926 9203
rect 6012 9180 6067 9203
rect 6067 9180 6084 9203
rect 6084 9180 6148 9203
rect 6148 9180 6165 9203
rect 6165 9180 6229 9203
rect 6229 9180 6246 9203
rect 6246 9180 6248 9203
rect 6333 9180 6391 9203
rect 6391 9180 6408 9203
rect 6408 9180 6472 9203
rect 6472 9180 6489 9203
rect 6489 9180 6553 9203
rect 6553 9180 6569 9203
rect 6654 9180 6715 9203
rect 6715 9180 6732 9203
rect 6732 9180 6796 9203
rect 6796 9180 6813 9203
rect 6813 9180 6877 9203
rect 6877 9180 6890 9203
rect 6975 9180 7039 9203
rect 7039 9180 7056 9203
rect 7056 9180 7120 9203
rect 7120 9180 7137 9203
rect 7137 9180 7201 9203
rect 7201 9180 7211 9203
rect 7296 9180 7299 9203
rect 7299 9180 7363 9203
rect 7363 9180 7380 9203
rect 7380 9180 7444 9203
rect 7444 9180 7461 9203
rect 7461 9180 7525 9203
rect 7525 9180 7532 9203
rect 7617 9180 7623 9203
rect 7623 9180 7687 9203
rect 7687 9180 7813 9203
rect 216 9158 452 9180
rect 538 9158 774 9180
rect 860 9158 1096 9180
rect 1182 9158 1418 9180
rect 1504 9158 1740 9180
rect 1826 9158 2062 9180
rect 2148 9158 2384 9180
rect 2470 9158 2706 9180
rect 2792 9158 3028 9180
rect 3114 9158 3350 9180
rect 3436 9158 3672 9180
rect 3758 9158 3994 9180
rect 4080 9158 4316 9180
rect 4402 9158 4638 9180
rect 4724 9158 4960 9180
rect 5046 9158 5282 9180
rect 5368 9158 5604 9180
rect 5690 9158 5926 9180
rect 6012 9158 6248 9180
rect 6333 9158 6569 9180
rect 6654 9158 6890 9180
rect 6975 9158 7211 9180
rect 7296 9158 7532 9180
rect 7617 9177 7813 9180
rect 7813 9177 7853 9203
rect 7938 9177 7961 9203
rect 7961 9177 7981 9203
rect 7981 9177 8045 9203
rect 8045 9177 8065 9203
rect 8065 9177 8129 9203
rect 8129 9177 8149 9203
rect 8149 9177 8174 9203
rect 7617 9158 7853 9177
rect 216 9094 397 9158
rect 397 9094 452 9158
rect 538 9094 543 9158
rect 543 9094 561 9158
rect 561 9094 625 9158
rect 625 9094 643 9158
rect 643 9094 707 9158
rect 707 9094 725 9158
rect 725 9094 774 9158
rect 860 9094 871 9158
rect 871 9094 889 9158
rect 889 9094 953 9158
rect 953 9094 971 9158
rect 971 9094 1035 9158
rect 1035 9094 1053 9158
rect 1053 9094 1096 9158
rect 1182 9094 1199 9158
rect 1199 9094 1217 9158
rect 1217 9094 1281 9158
rect 1281 9094 1299 9158
rect 1299 9094 1363 9158
rect 1363 9094 1381 9158
rect 1381 9094 1418 9158
rect 1504 9094 1527 9158
rect 1527 9094 1545 9158
rect 1545 9094 1609 9158
rect 1609 9094 1627 9158
rect 1627 9094 1691 9158
rect 1691 9094 1709 9158
rect 1709 9094 1740 9158
rect 1826 9094 1855 9158
rect 1855 9094 1873 9158
rect 1873 9094 1937 9158
rect 1937 9094 1955 9158
rect 1955 9094 2019 9158
rect 2019 9094 2037 9158
rect 2037 9094 2062 9158
rect 2148 9094 2183 9158
rect 2183 9094 2201 9158
rect 2201 9094 2265 9158
rect 2265 9094 2282 9158
rect 2282 9094 2346 9158
rect 2346 9094 2363 9158
rect 2363 9094 2384 9158
rect 2470 9094 2553 9158
rect 2553 9094 2617 9158
rect 2617 9094 2635 9158
rect 2635 9094 2699 9158
rect 2699 9094 2706 9158
rect 2792 9094 2799 9158
rect 2799 9094 2863 9158
rect 2863 9094 2881 9158
rect 2881 9094 2945 9158
rect 2945 9094 2963 9158
rect 2963 9094 3027 9158
rect 3027 9094 3028 9158
rect 3114 9094 3127 9158
rect 3127 9094 3191 9158
rect 3191 9094 3209 9158
rect 3209 9094 3273 9158
rect 3273 9094 3290 9158
rect 3290 9094 3350 9158
rect 3436 9094 3452 9158
rect 3452 9094 3516 9158
rect 3516 9094 3533 9158
rect 3533 9094 3597 9158
rect 3597 9094 3614 9158
rect 3614 9094 3672 9158
rect 3758 9094 3759 9158
rect 3759 9094 3776 9158
rect 3776 9094 3840 9158
rect 3840 9094 3857 9158
rect 3857 9094 3921 9158
rect 3921 9094 3938 9158
rect 3938 9094 3994 9158
rect 4080 9094 4083 9158
rect 4083 9094 4100 9158
rect 4100 9094 4164 9158
rect 4164 9094 4181 9158
rect 4181 9094 4245 9158
rect 4245 9094 4262 9158
rect 4262 9094 4316 9158
rect 4402 9094 4407 9158
rect 4407 9094 4424 9158
rect 4424 9094 4488 9158
rect 4488 9094 4505 9158
rect 4505 9094 4569 9158
rect 4569 9094 4638 9158
rect 4724 9094 4759 9158
rect 4759 9094 4777 9158
rect 4777 9094 4841 9158
rect 4841 9094 4859 9158
rect 4859 9094 4923 9158
rect 4923 9094 4941 9158
rect 4941 9094 4960 9158
rect 5046 9094 5087 9158
rect 5087 9094 5105 9158
rect 5105 9094 5169 9158
rect 5169 9094 5187 9158
rect 5187 9094 5251 9158
rect 5251 9094 5269 9158
rect 5269 9094 5282 9158
rect 5368 9094 5415 9158
rect 5415 9094 5433 9158
rect 5433 9094 5497 9158
rect 5497 9094 5515 9158
rect 5515 9094 5579 9158
rect 5579 9094 5597 9158
rect 5597 9094 5604 9158
rect 5690 9094 5743 9158
rect 5743 9094 5760 9158
rect 5760 9094 5824 9158
rect 5824 9094 5841 9158
rect 5841 9094 5905 9158
rect 5905 9094 5922 9158
rect 5922 9094 5926 9158
rect 6012 9094 6067 9158
rect 6067 9094 6084 9158
rect 6084 9094 6148 9158
rect 6148 9094 6165 9158
rect 6165 9094 6229 9158
rect 6229 9094 6246 9158
rect 6246 9094 6248 9158
rect 6333 9094 6391 9158
rect 6391 9094 6408 9158
rect 6408 9094 6472 9158
rect 6472 9094 6489 9158
rect 6489 9094 6553 9158
rect 6553 9094 6569 9158
rect 6654 9094 6715 9158
rect 6715 9094 6732 9158
rect 6732 9094 6796 9158
rect 6796 9094 6813 9158
rect 6813 9094 6877 9158
rect 6877 9094 6890 9158
rect 6975 9094 7039 9158
rect 7039 9094 7056 9158
rect 7056 9094 7120 9158
rect 7120 9094 7137 9158
rect 7137 9094 7201 9158
rect 7201 9094 7211 9158
rect 7296 9094 7299 9158
rect 7299 9094 7363 9158
rect 7363 9094 7380 9158
rect 7380 9094 7444 9158
rect 7444 9094 7461 9158
rect 7461 9094 7525 9158
rect 7525 9094 7532 9158
rect 7617 9094 7623 9158
rect 7623 9094 7687 9158
rect 7687 9156 7853 9158
rect 7938 9156 8174 9177
rect 7687 9094 7813 9156
rect 216 9072 452 9094
rect 538 9072 774 9094
rect 860 9072 1096 9094
rect 1182 9072 1418 9094
rect 1504 9072 1740 9094
rect 1826 9072 2062 9094
rect 2148 9072 2384 9094
rect 2470 9072 2706 9094
rect 2792 9072 3028 9094
rect 3114 9072 3350 9094
rect 3436 9072 3672 9094
rect 3758 9072 3994 9094
rect 4080 9072 4316 9094
rect 4402 9072 4638 9094
rect 4724 9072 4960 9094
rect 5046 9072 5282 9094
rect 5368 9072 5604 9094
rect 5690 9072 5926 9094
rect 6012 9072 6248 9094
rect 6333 9072 6569 9094
rect 6654 9072 6890 9094
rect 6975 9072 7211 9094
rect 7296 9072 7532 9094
rect 7617 9092 7813 9094
rect 7813 9092 7853 9156
rect 7938 9092 7961 9156
rect 7961 9092 7981 9156
rect 7981 9092 8045 9156
rect 8045 9092 8065 9156
rect 8065 9092 8129 9156
rect 8129 9092 8149 9156
rect 8149 9092 8174 9156
rect 7617 9072 7853 9092
rect 216 9008 397 9072
rect 397 9008 452 9072
rect 538 9008 543 9072
rect 543 9008 561 9072
rect 561 9008 625 9072
rect 625 9008 643 9072
rect 643 9008 707 9072
rect 707 9008 725 9072
rect 725 9008 774 9072
rect 860 9008 871 9072
rect 871 9008 889 9072
rect 889 9008 953 9072
rect 953 9008 971 9072
rect 971 9008 1035 9072
rect 1035 9008 1053 9072
rect 1053 9008 1096 9072
rect 1182 9008 1199 9072
rect 1199 9008 1217 9072
rect 1217 9008 1281 9072
rect 1281 9008 1299 9072
rect 1299 9008 1363 9072
rect 1363 9008 1381 9072
rect 1381 9008 1418 9072
rect 1504 9008 1527 9072
rect 1527 9008 1545 9072
rect 1545 9008 1609 9072
rect 1609 9008 1627 9072
rect 1627 9008 1691 9072
rect 1691 9008 1709 9072
rect 1709 9008 1740 9072
rect 1826 9008 1855 9072
rect 1855 9008 1873 9072
rect 1873 9008 1937 9072
rect 1937 9008 1955 9072
rect 1955 9008 2019 9072
rect 2019 9008 2037 9072
rect 2037 9008 2062 9072
rect 2148 9008 2183 9072
rect 2183 9008 2201 9072
rect 2201 9008 2265 9072
rect 2265 9008 2282 9072
rect 2282 9008 2346 9072
rect 2346 9008 2363 9072
rect 2363 9008 2384 9072
rect 2470 9008 2553 9072
rect 2553 9008 2617 9072
rect 2617 9008 2635 9072
rect 2635 9008 2699 9072
rect 2699 9008 2706 9072
rect 2792 9008 2799 9072
rect 2799 9008 2863 9072
rect 2863 9008 2881 9072
rect 2881 9008 2945 9072
rect 2945 9008 2963 9072
rect 2963 9008 3027 9072
rect 3027 9008 3028 9072
rect 3114 9008 3127 9072
rect 3127 9008 3191 9072
rect 3191 9008 3209 9072
rect 3209 9008 3273 9072
rect 3273 9008 3290 9072
rect 3290 9008 3350 9072
rect 3436 9008 3452 9072
rect 3452 9008 3516 9072
rect 3516 9008 3533 9072
rect 3533 9008 3597 9072
rect 3597 9008 3614 9072
rect 3614 9008 3672 9072
rect 3758 9008 3759 9072
rect 3759 9008 3776 9072
rect 3776 9008 3840 9072
rect 3840 9008 3857 9072
rect 3857 9008 3921 9072
rect 3921 9008 3938 9072
rect 3938 9008 3994 9072
rect 4080 9008 4083 9072
rect 4083 9008 4100 9072
rect 4100 9008 4164 9072
rect 4164 9008 4181 9072
rect 4181 9008 4245 9072
rect 4245 9008 4262 9072
rect 4262 9008 4316 9072
rect 4402 9008 4407 9072
rect 4407 9008 4424 9072
rect 4424 9008 4488 9072
rect 4488 9008 4505 9072
rect 4505 9008 4569 9072
rect 4569 9008 4638 9072
rect 4724 9008 4759 9072
rect 4759 9008 4777 9072
rect 4777 9008 4841 9072
rect 4841 9008 4859 9072
rect 4859 9008 4923 9072
rect 4923 9008 4941 9072
rect 4941 9008 4960 9072
rect 5046 9008 5087 9072
rect 5087 9008 5105 9072
rect 5105 9008 5169 9072
rect 5169 9008 5187 9072
rect 5187 9008 5251 9072
rect 5251 9008 5269 9072
rect 5269 9008 5282 9072
rect 5368 9008 5415 9072
rect 5415 9008 5433 9072
rect 5433 9008 5497 9072
rect 5497 9008 5515 9072
rect 5515 9008 5579 9072
rect 5579 9008 5597 9072
rect 5597 9008 5604 9072
rect 5690 9008 5743 9072
rect 5743 9008 5760 9072
rect 5760 9008 5824 9072
rect 5824 9008 5841 9072
rect 5841 9008 5905 9072
rect 5905 9008 5922 9072
rect 5922 9008 5926 9072
rect 6012 9008 6067 9072
rect 6067 9008 6084 9072
rect 6084 9008 6148 9072
rect 6148 9008 6165 9072
rect 6165 9008 6229 9072
rect 6229 9008 6246 9072
rect 6246 9008 6248 9072
rect 6333 9008 6391 9072
rect 6391 9008 6408 9072
rect 6408 9008 6472 9072
rect 6472 9008 6489 9072
rect 6489 9008 6553 9072
rect 6553 9008 6569 9072
rect 6654 9008 6715 9072
rect 6715 9008 6732 9072
rect 6732 9008 6796 9072
rect 6796 9008 6813 9072
rect 6813 9008 6877 9072
rect 6877 9008 6890 9072
rect 6975 9008 7039 9072
rect 7039 9008 7056 9072
rect 7056 9008 7120 9072
rect 7120 9008 7137 9072
rect 7137 9008 7201 9072
rect 7201 9008 7211 9072
rect 7296 9008 7299 9072
rect 7299 9008 7363 9072
rect 7363 9008 7380 9072
rect 7380 9008 7444 9072
rect 7444 9008 7461 9072
rect 7461 9008 7525 9072
rect 7525 9008 7532 9072
rect 7617 9008 7623 9072
rect 7623 9008 7687 9072
rect 7687 9071 7853 9072
rect 7938 9071 8174 9092
rect 7687 9008 7813 9071
rect 216 8986 452 9008
rect 538 8986 774 9008
rect 860 8986 1096 9008
rect 1182 8986 1418 9008
rect 1504 8986 1740 9008
rect 1826 8986 2062 9008
rect 2148 8986 2384 9008
rect 2470 8986 2706 9008
rect 2792 8986 3028 9008
rect 3114 8986 3350 9008
rect 3436 8986 3672 9008
rect 3758 8986 3994 9008
rect 4080 8986 4316 9008
rect 4402 8986 4638 9008
rect 4724 8986 4960 9008
rect 5046 8986 5282 9008
rect 5368 8986 5604 9008
rect 5690 8986 5926 9008
rect 6012 8986 6248 9008
rect 6333 8986 6569 9008
rect 6654 8986 6890 9008
rect 6975 8986 7211 9008
rect 7296 8986 7532 9008
rect 7617 9007 7813 9008
rect 7813 9007 7853 9071
rect 7938 9007 7961 9071
rect 7961 9007 7981 9071
rect 7981 9007 8045 9071
rect 8045 9007 8065 9071
rect 8065 9007 8129 9071
rect 8129 9007 8149 9071
rect 8149 9007 8174 9071
rect 7617 8986 7853 9007
rect 7938 8986 8174 9007
rect 216 8967 397 8986
rect 397 8967 452 8986
rect 538 8967 543 8986
rect 543 8967 561 8986
rect 561 8967 625 8986
rect 625 8967 643 8986
rect 643 8967 707 8986
rect 707 8967 725 8986
rect 725 8967 774 8986
rect 860 8967 871 8986
rect 871 8967 889 8986
rect 889 8967 953 8986
rect 953 8967 971 8986
rect 971 8967 1035 8986
rect 1035 8967 1053 8986
rect 1053 8967 1096 8986
rect 1182 8967 1199 8986
rect 1199 8967 1217 8986
rect 1217 8967 1281 8986
rect 1281 8967 1299 8986
rect 1299 8967 1363 8986
rect 1363 8967 1381 8986
rect 1381 8967 1418 8986
rect 1504 8967 1527 8986
rect 1527 8967 1545 8986
rect 1545 8967 1609 8986
rect 1609 8967 1627 8986
rect 1627 8967 1691 8986
rect 1691 8967 1709 8986
rect 1709 8967 1740 8986
rect 1826 8967 1855 8986
rect 1855 8967 1873 8986
rect 1873 8967 1937 8986
rect 1937 8967 1955 8986
rect 1955 8967 2019 8986
rect 2019 8967 2037 8986
rect 2037 8967 2062 8986
rect 2148 8967 2183 8986
rect 2183 8967 2201 8986
rect 2201 8967 2265 8986
rect 2265 8967 2282 8986
rect 2282 8967 2346 8986
rect 2346 8967 2363 8986
rect 2363 8967 2384 8986
rect 2470 8967 2553 8986
rect 2553 8967 2617 8986
rect 2617 8967 2635 8986
rect 2635 8967 2699 8986
rect 2699 8967 2706 8986
rect 2792 8967 2799 8986
rect 2799 8967 2863 8986
rect 2863 8967 2881 8986
rect 2881 8967 2945 8986
rect 2945 8967 2963 8986
rect 2963 8967 3027 8986
rect 3027 8967 3028 8986
rect 3114 8967 3127 8986
rect 3127 8967 3191 8986
rect 3191 8967 3209 8986
rect 3209 8967 3273 8986
rect 3273 8967 3290 8986
rect 3290 8967 3350 8986
rect 3436 8967 3452 8986
rect 3452 8967 3516 8986
rect 3516 8967 3533 8986
rect 3533 8967 3597 8986
rect 3597 8967 3614 8986
rect 3614 8967 3672 8986
rect 3758 8967 3759 8986
rect 3759 8967 3776 8986
rect 3776 8967 3840 8986
rect 3840 8967 3857 8986
rect 3857 8967 3921 8986
rect 3921 8967 3938 8986
rect 3938 8967 3994 8986
rect 4080 8967 4083 8986
rect 4083 8967 4100 8986
rect 4100 8967 4164 8986
rect 4164 8967 4181 8986
rect 4181 8967 4245 8986
rect 4245 8967 4262 8986
rect 4262 8967 4316 8986
rect 4402 8967 4407 8986
rect 4407 8967 4424 8986
rect 4424 8967 4488 8986
rect 4488 8967 4505 8986
rect 4505 8967 4569 8986
rect 4569 8967 4638 8986
rect 4724 8967 4759 8986
rect 4759 8967 4777 8986
rect 4777 8967 4841 8986
rect 4841 8967 4859 8986
rect 4859 8967 4923 8986
rect 4923 8967 4941 8986
rect 4941 8967 4960 8986
rect 5046 8967 5087 8986
rect 5087 8967 5105 8986
rect 5105 8967 5169 8986
rect 5169 8967 5187 8986
rect 5187 8967 5251 8986
rect 5251 8967 5269 8986
rect 5269 8967 5282 8986
rect 5368 8967 5415 8986
rect 5415 8967 5433 8986
rect 5433 8967 5497 8986
rect 5497 8967 5515 8986
rect 5515 8967 5579 8986
rect 5579 8967 5597 8986
rect 5597 8967 5604 8986
rect 5690 8967 5743 8986
rect 5743 8967 5760 8986
rect 5760 8967 5824 8986
rect 5824 8967 5841 8986
rect 5841 8967 5905 8986
rect 5905 8967 5922 8986
rect 5922 8967 5926 8986
rect 6012 8967 6067 8986
rect 6067 8967 6084 8986
rect 6084 8967 6148 8986
rect 6148 8967 6165 8986
rect 6165 8967 6229 8986
rect 6229 8967 6246 8986
rect 6246 8967 6248 8986
rect 6333 8967 6391 8986
rect 6391 8967 6408 8986
rect 6408 8967 6472 8986
rect 6472 8967 6489 8986
rect 6489 8967 6553 8986
rect 6553 8967 6569 8986
rect 6654 8967 6715 8986
rect 6715 8967 6732 8986
rect 6732 8967 6796 8986
rect 6796 8967 6813 8986
rect 6813 8967 6877 8986
rect 6877 8967 6890 8986
rect 6975 8967 7039 8986
rect 7039 8967 7056 8986
rect 7056 8967 7120 8986
rect 7120 8967 7137 8986
rect 7137 8967 7201 8986
rect 7201 8967 7211 8986
rect 7296 8967 7299 8986
rect 7299 8967 7363 8986
rect 7363 8967 7380 8986
rect 7380 8967 7444 8986
rect 7444 8967 7461 8986
rect 7461 8967 7525 8986
rect 7525 8967 7532 8986
rect 7617 8967 7623 8986
rect 7623 8967 7687 8986
rect 7687 8967 7813 8986
rect 7813 8967 7853 8986
rect 7938 8967 7961 8986
rect 7961 8967 7981 8986
rect 7981 8967 8045 8986
rect 8045 8967 8065 8986
rect 8065 8967 8129 8986
rect 8129 8967 8149 8986
rect 8149 8967 8174 8986
rect 8259 8967 8495 9203
rect 8580 8967 8816 9203
rect 8901 9180 8923 9203
rect 8923 9180 8940 9203
rect 8940 9180 9004 9203
rect 9004 9180 9021 9203
rect 9021 9180 9085 9203
rect 9085 9180 9102 9203
rect 9102 9180 9137 9203
rect 9222 9180 9247 9203
rect 9247 9180 9264 9203
rect 9264 9180 9328 9203
rect 9328 9180 9345 9203
rect 9345 9180 9409 9203
rect 9409 9180 9426 9203
rect 9426 9180 9458 9203
rect 9543 9180 9571 9203
rect 9571 9180 9588 9203
rect 9588 9180 9652 9203
rect 9652 9180 9669 9203
rect 9669 9180 9733 9203
rect 9733 9180 9750 9203
rect 9750 9180 9779 9203
rect 9864 9180 9895 9203
rect 9895 9180 9912 9203
rect 9912 9180 9976 9203
rect 9976 9180 9993 9203
rect 9993 9180 10057 9203
rect 10057 9180 10073 9203
rect 10073 9180 10100 9203
rect 10185 9180 10217 9203
rect 10217 9180 10233 9203
rect 10233 9180 10297 9203
rect 10297 9180 10313 9203
rect 10313 9180 10377 9203
rect 10377 9180 10393 9203
rect 10393 9180 10421 9203
rect 10506 9180 10537 9203
rect 10537 9180 10553 9203
rect 10553 9180 10617 9203
rect 10617 9180 10633 9203
rect 10633 9180 10697 9203
rect 10697 9180 10713 9203
rect 10713 9180 10742 9203
rect 10827 9180 10857 9203
rect 10857 9180 10873 9203
rect 10873 9180 10937 9203
rect 10937 9180 10953 9203
rect 10953 9180 11017 9203
rect 11017 9180 11033 9203
rect 11033 9180 11063 9203
rect 11148 9180 11177 9203
rect 11177 9180 11193 9203
rect 11193 9180 11257 9203
rect 11257 9180 11273 9203
rect 11273 9180 11337 9203
rect 11337 9180 11353 9203
rect 11353 9180 11384 9203
rect 11469 9180 11497 9203
rect 11497 9180 11513 9203
rect 11513 9180 11577 9203
rect 11577 9180 11593 9203
rect 11593 9180 11657 9203
rect 11657 9180 11673 9203
rect 11673 9180 11705 9203
rect 11790 9180 11817 9203
rect 11817 9180 11833 9203
rect 11833 9180 11897 9203
rect 11897 9180 11913 9203
rect 11913 9180 11977 9203
rect 11977 9180 12026 9203
rect 8901 9158 9137 9180
rect 9222 9158 9458 9180
rect 9543 9158 9779 9180
rect 9864 9158 10100 9180
rect 10185 9158 10421 9180
rect 10506 9158 10742 9180
rect 10827 9158 11063 9180
rect 11148 9158 11384 9180
rect 11469 9158 11705 9180
rect 11790 9158 12026 9180
rect 8901 9094 8923 9158
rect 8923 9094 8940 9158
rect 8940 9094 9004 9158
rect 9004 9094 9021 9158
rect 9021 9094 9085 9158
rect 9085 9094 9102 9158
rect 9102 9094 9137 9158
rect 9222 9094 9247 9158
rect 9247 9094 9264 9158
rect 9264 9094 9328 9158
rect 9328 9094 9345 9158
rect 9345 9094 9409 9158
rect 9409 9094 9426 9158
rect 9426 9094 9458 9158
rect 9543 9094 9571 9158
rect 9571 9094 9588 9158
rect 9588 9094 9652 9158
rect 9652 9094 9669 9158
rect 9669 9094 9733 9158
rect 9733 9094 9750 9158
rect 9750 9094 9779 9158
rect 9864 9094 9895 9158
rect 9895 9094 9912 9158
rect 9912 9094 9976 9158
rect 9976 9094 9993 9158
rect 9993 9094 10057 9158
rect 10057 9094 10073 9158
rect 10073 9094 10100 9158
rect 10185 9094 10217 9158
rect 10217 9094 10233 9158
rect 10233 9094 10297 9158
rect 10297 9094 10313 9158
rect 10313 9094 10377 9158
rect 10377 9094 10393 9158
rect 10393 9094 10421 9158
rect 10506 9094 10537 9158
rect 10537 9094 10553 9158
rect 10553 9094 10617 9158
rect 10617 9094 10633 9158
rect 10633 9094 10697 9158
rect 10697 9094 10713 9158
rect 10713 9094 10742 9158
rect 10827 9094 10857 9158
rect 10857 9094 10873 9158
rect 10873 9094 10937 9158
rect 10937 9094 10953 9158
rect 10953 9094 11017 9158
rect 11017 9094 11033 9158
rect 11033 9094 11063 9158
rect 11148 9094 11177 9158
rect 11177 9094 11193 9158
rect 11193 9094 11257 9158
rect 11257 9094 11273 9158
rect 11273 9094 11337 9158
rect 11337 9094 11353 9158
rect 11353 9094 11384 9158
rect 11469 9094 11497 9158
rect 11497 9094 11513 9158
rect 11513 9094 11577 9158
rect 11577 9094 11593 9158
rect 11593 9094 11657 9158
rect 11657 9094 11673 9158
rect 11673 9094 11705 9158
rect 11790 9094 11817 9158
rect 11817 9094 11833 9158
rect 11833 9094 11897 9158
rect 11897 9094 11913 9158
rect 11913 9094 11977 9158
rect 11977 9094 12026 9158
rect 8901 9072 9137 9094
rect 9222 9072 9458 9094
rect 9543 9072 9779 9094
rect 9864 9072 10100 9094
rect 10185 9072 10421 9094
rect 10506 9072 10742 9094
rect 10827 9072 11063 9094
rect 11148 9072 11384 9094
rect 11469 9072 11705 9094
rect 11790 9072 12026 9094
rect 8901 9008 8923 9072
rect 8923 9008 8940 9072
rect 8940 9008 9004 9072
rect 9004 9008 9021 9072
rect 9021 9008 9085 9072
rect 9085 9008 9102 9072
rect 9102 9008 9137 9072
rect 9222 9008 9247 9072
rect 9247 9008 9264 9072
rect 9264 9008 9328 9072
rect 9328 9008 9345 9072
rect 9345 9008 9409 9072
rect 9409 9008 9426 9072
rect 9426 9008 9458 9072
rect 9543 9008 9571 9072
rect 9571 9008 9588 9072
rect 9588 9008 9652 9072
rect 9652 9008 9669 9072
rect 9669 9008 9733 9072
rect 9733 9008 9750 9072
rect 9750 9008 9779 9072
rect 9864 9008 9895 9072
rect 9895 9008 9912 9072
rect 9912 9008 9976 9072
rect 9976 9008 9993 9072
rect 9993 9008 10057 9072
rect 10057 9008 10073 9072
rect 10073 9008 10100 9072
rect 10185 9008 10217 9072
rect 10217 9008 10233 9072
rect 10233 9008 10297 9072
rect 10297 9008 10313 9072
rect 10313 9008 10377 9072
rect 10377 9008 10393 9072
rect 10393 9008 10421 9072
rect 10506 9008 10537 9072
rect 10537 9008 10553 9072
rect 10553 9008 10617 9072
rect 10617 9008 10633 9072
rect 10633 9008 10697 9072
rect 10697 9008 10713 9072
rect 10713 9008 10742 9072
rect 10827 9008 10857 9072
rect 10857 9008 10873 9072
rect 10873 9008 10937 9072
rect 10937 9008 10953 9072
rect 10953 9008 11017 9072
rect 11017 9008 11033 9072
rect 11033 9008 11063 9072
rect 11148 9008 11177 9072
rect 11177 9008 11193 9072
rect 11193 9008 11257 9072
rect 11257 9008 11273 9072
rect 11273 9008 11337 9072
rect 11337 9008 11353 9072
rect 11353 9008 11384 9072
rect 11469 9008 11497 9072
rect 11497 9008 11513 9072
rect 11513 9008 11577 9072
rect 11577 9008 11593 9072
rect 11593 9008 11657 9072
rect 11657 9008 11673 9072
rect 11673 9008 11705 9072
rect 11790 9008 11817 9072
rect 11817 9008 11833 9072
rect 11833 9008 11897 9072
rect 11897 9008 11913 9072
rect 11913 9008 11977 9072
rect 11977 9008 12026 9072
rect 8901 8986 9137 9008
rect 9222 8986 9458 9008
rect 9543 8986 9779 9008
rect 9864 8986 10100 9008
rect 10185 8986 10421 9008
rect 10506 8986 10742 9008
rect 10827 8986 11063 9008
rect 11148 8986 11384 9008
rect 11469 8986 11705 9008
rect 11790 8986 12026 9008
rect 8901 8967 8923 8986
rect 8923 8967 8940 8986
rect 8940 8967 9004 8986
rect 9004 8967 9021 8986
rect 9021 8967 9085 8986
rect 9085 8967 9102 8986
rect 9102 8967 9137 8986
rect 9222 8967 9247 8986
rect 9247 8967 9264 8986
rect 9264 8967 9328 8986
rect 9328 8967 9345 8986
rect 9345 8967 9409 8986
rect 9409 8967 9426 8986
rect 9426 8967 9458 8986
rect 9543 8967 9571 8986
rect 9571 8967 9588 8986
rect 9588 8967 9652 8986
rect 9652 8967 9669 8986
rect 9669 8967 9733 8986
rect 9733 8967 9750 8986
rect 9750 8967 9779 8986
rect 9864 8967 9895 8986
rect 9895 8967 9912 8986
rect 9912 8967 9976 8986
rect 9976 8967 9993 8986
rect 9993 8967 10057 8986
rect 10057 8967 10073 8986
rect 10073 8967 10100 8986
rect 10185 8967 10217 8986
rect 10217 8967 10233 8986
rect 10233 8967 10297 8986
rect 10297 8967 10313 8986
rect 10313 8967 10377 8986
rect 10377 8967 10393 8986
rect 10393 8967 10421 8986
rect 10506 8967 10537 8986
rect 10537 8967 10553 8986
rect 10553 8967 10617 8986
rect 10617 8967 10633 8986
rect 10633 8967 10697 8986
rect 10697 8967 10713 8986
rect 10713 8967 10742 8986
rect 10827 8967 10857 8986
rect 10857 8967 10873 8986
rect 10873 8967 10937 8986
rect 10937 8967 10953 8986
rect 10953 8967 11017 8986
rect 11017 8967 11033 8986
rect 11033 8967 11063 8986
rect 11148 8967 11177 8986
rect 11177 8967 11193 8986
rect 11193 8967 11257 8986
rect 11257 8967 11273 8986
rect 11273 8967 11337 8986
rect 11337 8967 11353 8986
rect 11353 8967 11384 8986
rect 11469 8967 11497 8986
rect 11497 8967 11513 8986
rect 11513 8967 11577 8986
rect 11577 8967 11593 8986
rect 11593 8967 11657 8986
rect 11657 8967 11673 8986
rect 11673 8967 11705 8986
rect 11790 8967 11817 8986
rect 11817 8967 11833 8986
rect 11833 8967 11897 8986
rect 11897 8967 11913 8986
rect 11913 8967 11977 8986
rect 11977 8967 12026 8986
rect 12111 9180 12165 9203
rect 12165 9180 12229 9203
rect 12229 9180 12246 9203
rect 12246 9180 12310 9203
rect 12310 9180 12327 9203
rect 12327 9180 12347 9203
rect 12432 9180 12472 9203
rect 12472 9180 12489 9203
rect 12489 9180 12553 9203
rect 12553 9180 12570 9203
rect 12570 9180 12634 9203
rect 12634 9180 12651 9203
rect 12651 9180 12668 9203
rect 12753 9180 12796 9203
rect 12796 9180 12813 9203
rect 12813 9180 12877 9203
rect 12877 9180 12894 9203
rect 12894 9180 12958 9203
rect 12958 9180 12975 9203
rect 12975 9180 12989 9203
rect 13074 9180 13120 9203
rect 13120 9180 13137 9203
rect 13137 9180 13201 9203
rect 13201 9180 13218 9203
rect 13218 9180 13282 9203
rect 13282 9180 13299 9203
rect 13299 9180 13310 9203
rect 13395 9180 13444 9203
rect 13444 9180 13461 9203
rect 13461 9180 13525 9203
rect 13525 9180 13542 9203
rect 13542 9180 13606 9203
rect 13606 9180 13623 9203
rect 13623 9180 13631 9203
rect 13716 9180 13768 9203
rect 13768 9180 13785 9203
rect 13785 9180 13849 9203
rect 13849 9180 13866 9203
rect 13866 9180 13930 9203
rect 13930 9180 13947 9203
rect 13947 9180 13952 9203
rect 14037 9180 14092 9203
rect 14092 9180 14109 9203
rect 14109 9180 14173 9203
rect 14173 9180 14190 9203
rect 14190 9180 14254 9203
rect 14254 9180 14271 9203
rect 14271 9180 14273 9203
rect 14358 9180 14416 9203
rect 14416 9180 14433 9203
rect 14433 9180 14497 9203
rect 14497 9180 14513 9203
rect 14513 9180 14577 9203
rect 14577 9180 14593 9203
rect 14593 9180 14594 9203
rect 14679 9180 14737 9203
rect 14737 9180 14753 9203
rect 14753 9180 14817 9203
rect 14817 9180 14833 9203
rect 14833 9180 14897 9203
rect 14897 9180 14913 9203
rect 14913 9180 14915 9203
rect 15000 9180 15057 9203
rect 15057 9180 15073 9203
rect 15073 9180 15137 9203
rect 15137 9180 15153 9203
rect 15153 9180 15217 9203
rect 15217 9180 15233 9203
rect 15233 9180 15236 9203
rect 15321 9180 15377 9203
rect 15377 9180 15393 9203
rect 15393 9180 15457 9203
rect 15457 9180 15473 9203
rect 15473 9180 15537 9203
rect 15537 9180 15553 9203
rect 15553 9180 15557 9203
rect 12111 9158 12347 9180
rect 12432 9158 12668 9180
rect 12753 9158 12989 9180
rect 13074 9158 13310 9180
rect 13395 9158 13631 9180
rect 13716 9158 13952 9180
rect 14037 9158 14273 9180
rect 14358 9158 14594 9180
rect 14679 9158 14915 9180
rect 15000 9158 15236 9180
rect 15321 9158 15557 9180
rect 12111 9094 12165 9158
rect 12165 9094 12229 9158
rect 12229 9094 12246 9158
rect 12246 9094 12310 9158
rect 12310 9094 12327 9158
rect 12327 9094 12347 9158
rect 12432 9094 12472 9158
rect 12472 9094 12489 9158
rect 12489 9094 12553 9158
rect 12553 9094 12570 9158
rect 12570 9094 12634 9158
rect 12634 9094 12651 9158
rect 12651 9094 12668 9158
rect 12753 9094 12796 9158
rect 12796 9094 12813 9158
rect 12813 9094 12877 9158
rect 12877 9094 12894 9158
rect 12894 9094 12958 9158
rect 12958 9094 12975 9158
rect 12975 9094 12989 9158
rect 13074 9094 13120 9158
rect 13120 9094 13137 9158
rect 13137 9094 13201 9158
rect 13201 9094 13218 9158
rect 13218 9094 13282 9158
rect 13282 9094 13299 9158
rect 13299 9094 13310 9158
rect 13395 9094 13444 9158
rect 13444 9094 13461 9158
rect 13461 9094 13525 9158
rect 13525 9094 13542 9158
rect 13542 9094 13606 9158
rect 13606 9094 13623 9158
rect 13623 9094 13631 9158
rect 13716 9094 13768 9158
rect 13768 9094 13785 9158
rect 13785 9094 13849 9158
rect 13849 9094 13866 9158
rect 13866 9094 13930 9158
rect 13930 9094 13947 9158
rect 13947 9094 13952 9158
rect 14037 9094 14092 9158
rect 14092 9094 14109 9158
rect 14109 9094 14173 9158
rect 14173 9094 14190 9158
rect 14190 9094 14254 9158
rect 14254 9094 14271 9158
rect 14271 9094 14273 9158
rect 14358 9094 14416 9158
rect 14416 9094 14433 9158
rect 14433 9094 14497 9158
rect 14497 9094 14513 9158
rect 14513 9094 14577 9158
rect 14577 9094 14593 9158
rect 14593 9094 14594 9158
rect 14679 9094 14737 9158
rect 14737 9094 14753 9158
rect 14753 9094 14817 9158
rect 14817 9094 14833 9158
rect 14833 9094 14897 9158
rect 14897 9094 14913 9158
rect 14913 9094 14915 9158
rect 15000 9094 15057 9158
rect 15057 9094 15073 9158
rect 15073 9094 15137 9158
rect 15137 9094 15153 9158
rect 15153 9094 15217 9158
rect 15217 9094 15233 9158
rect 15233 9094 15236 9158
rect 15321 9094 15377 9158
rect 15377 9094 15393 9158
rect 15393 9094 15457 9158
rect 15457 9094 15473 9158
rect 15473 9094 15537 9158
rect 15537 9094 15553 9158
rect 15553 9094 15557 9158
rect 12111 9072 12347 9094
rect 12432 9072 12668 9094
rect 12753 9072 12989 9094
rect 13074 9072 13310 9094
rect 13395 9072 13631 9094
rect 13716 9072 13952 9094
rect 14037 9072 14273 9094
rect 14358 9072 14594 9094
rect 14679 9072 14915 9094
rect 15000 9072 15236 9094
rect 15321 9072 15557 9094
rect 12111 9008 12165 9072
rect 12165 9008 12229 9072
rect 12229 9008 12246 9072
rect 12246 9008 12310 9072
rect 12310 9008 12327 9072
rect 12327 9008 12347 9072
rect 12432 9008 12472 9072
rect 12472 9008 12489 9072
rect 12489 9008 12553 9072
rect 12553 9008 12570 9072
rect 12570 9008 12634 9072
rect 12634 9008 12651 9072
rect 12651 9008 12668 9072
rect 12753 9008 12796 9072
rect 12796 9008 12813 9072
rect 12813 9008 12877 9072
rect 12877 9008 12894 9072
rect 12894 9008 12958 9072
rect 12958 9008 12975 9072
rect 12975 9008 12989 9072
rect 13074 9008 13120 9072
rect 13120 9008 13137 9072
rect 13137 9008 13201 9072
rect 13201 9008 13218 9072
rect 13218 9008 13282 9072
rect 13282 9008 13299 9072
rect 13299 9008 13310 9072
rect 13395 9008 13444 9072
rect 13444 9008 13461 9072
rect 13461 9008 13525 9072
rect 13525 9008 13542 9072
rect 13542 9008 13606 9072
rect 13606 9008 13623 9072
rect 13623 9008 13631 9072
rect 13716 9008 13768 9072
rect 13768 9008 13785 9072
rect 13785 9008 13849 9072
rect 13849 9008 13866 9072
rect 13866 9008 13930 9072
rect 13930 9008 13947 9072
rect 13947 9008 13952 9072
rect 14037 9008 14092 9072
rect 14092 9008 14109 9072
rect 14109 9008 14173 9072
rect 14173 9008 14190 9072
rect 14190 9008 14254 9072
rect 14254 9008 14271 9072
rect 14271 9008 14273 9072
rect 14358 9008 14416 9072
rect 14416 9008 14433 9072
rect 14433 9008 14497 9072
rect 14497 9008 14513 9072
rect 14513 9008 14577 9072
rect 14577 9008 14593 9072
rect 14593 9008 14594 9072
rect 14679 9008 14737 9072
rect 14737 9008 14753 9072
rect 14753 9008 14817 9072
rect 14817 9008 14833 9072
rect 14833 9008 14897 9072
rect 14897 9008 14913 9072
rect 14913 9008 14915 9072
rect 15000 9008 15057 9072
rect 15057 9008 15073 9072
rect 15073 9008 15137 9072
rect 15137 9008 15153 9072
rect 15153 9008 15217 9072
rect 15217 9008 15233 9072
rect 15233 9008 15236 9072
rect 15321 9008 15377 9072
rect 15377 9008 15393 9072
rect 15393 9008 15457 9072
rect 15457 9008 15473 9072
rect 15473 9008 15537 9072
rect 15537 9008 15553 9072
rect 15553 9008 15557 9072
rect 12111 8986 12347 9008
rect 12432 8986 12668 9008
rect 12753 8986 12989 9008
rect 13074 8986 13310 9008
rect 13395 8986 13631 9008
rect 13716 8986 13952 9008
rect 14037 8986 14273 9008
rect 14358 8986 14594 9008
rect 14679 8986 14915 9008
rect 15000 8986 15236 9008
rect 15321 8986 15557 9008
rect 12111 8967 12165 8986
rect 12165 8967 12229 8986
rect 12229 8967 12246 8986
rect 12246 8967 12310 8986
rect 12310 8967 12327 8986
rect 12327 8967 12347 8986
rect 12432 8967 12472 8986
rect 12472 8967 12489 8986
rect 12489 8967 12553 8986
rect 12553 8967 12570 8986
rect 12570 8967 12634 8986
rect 12634 8967 12651 8986
rect 12651 8967 12668 8986
rect 12753 8967 12796 8986
rect 12796 8967 12813 8986
rect 12813 8967 12877 8986
rect 12877 8967 12894 8986
rect 12894 8967 12958 8986
rect 12958 8967 12975 8986
rect 12975 8967 12989 8986
rect 13074 8967 13120 8986
rect 13120 8967 13137 8986
rect 13137 8967 13201 8986
rect 13201 8967 13218 8986
rect 13218 8967 13282 8986
rect 13282 8967 13299 8986
rect 13299 8967 13310 8986
rect 13395 8967 13444 8986
rect 13444 8967 13461 8986
rect 13461 8967 13525 8986
rect 13525 8967 13542 8986
rect 13542 8967 13606 8986
rect 13606 8967 13623 8986
rect 13623 8967 13631 8986
rect 13716 8967 13768 8986
rect 13768 8967 13785 8986
rect 13785 8967 13849 8986
rect 13849 8967 13866 8986
rect 13866 8967 13930 8986
rect 13930 8967 13947 8986
rect 13947 8967 13952 8986
rect 14037 8967 14092 8986
rect 14092 8967 14109 8986
rect 14109 8967 14173 8986
rect 14173 8967 14190 8986
rect 14190 8967 14254 8986
rect 14254 8967 14271 8986
rect 14271 8967 14273 8986
rect 14358 8967 14416 8986
rect 14416 8967 14433 8986
rect 14433 8967 14497 8986
rect 14497 8967 14513 8986
rect 14513 8967 14577 8986
rect 14577 8967 14593 8986
rect 14593 8967 14594 8986
rect 14679 8967 14737 8986
rect 14737 8967 14753 8986
rect 14753 8967 14817 8986
rect 14817 8967 14833 8986
rect 14833 8967 14897 8986
rect 14897 8967 14913 8986
rect 14913 8967 14915 8986
rect 15000 8967 15057 8986
rect 15057 8967 15073 8986
rect 15073 8967 15137 8986
rect 15137 8967 15153 8986
rect 15153 8967 15217 8986
rect 15217 8967 15233 8986
rect 15233 8967 15236 8986
rect 15321 8967 15377 8986
rect 15377 8967 15393 8986
rect 15393 8967 15457 8986
rect 15457 8967 15473 8986
rect 15473 8967 15537 8986
rect 15537 8967 15553 8986
rect 15553 8967 15557 8986
rect 216 8578 397 8597
rect 397 8578 452 8597
rect 538 8578 543 8597
rect 543 8578 561 8597
rect 561 8578 625 8597
rect 625 8578 643 8597
rect 643 8578 707 8597
rect 707 8578 725 8597
rect 725 8578 774 8597
rect 860 8578 871 8597
rect 871 8578 889 8597
rect 889 8578 953 8597
rect 953 8578 971 8597
rect 971 8578 1035 8597
rect 1035 8578 1053 8597
rect 1053 8578 1096 8597
rect 1182 8578 1199 8597
rect 1199 8578 1217 8597
rect 1217 8578 1281 8597
rect 1281 8578 1299 8597
rect 1299 8578 1363 8597
rect 1363 8578 1381 8597
rect 1381 8578 1418 8597
rect 1504 8578 1527 8597
rect 1527 8578 1545 8597
rect 1545 8578 1609 8597
rect 1609 8578 1627 8597
rect 1627 8578 1691 8597
rect 1691 8578 1709 8597
rect 1709 8578 1740 8597
rect 1826 8578 1855 8597
rect 1855 8578 1873 8597
rect 1873 8578 1937 8597
rect 1937 8578 1955 8597
rect 1955 8578 2019 8597
rect 2019 8578 2037 8597
rect 2037 8578 2062 8597
rect 2148 8578 2183 8597
rect 2183 8578 2201 8597
rect 2201 8578 2265 8597
rect 2265 8578 2282 8597
rect 2282 8578 2346 8597
rect 2346 8578 2363 8597
rect 2363 8578 2384 8597
rect 2470 8578 2553 8597
rect 2553 8578 2617 8597
rect 2617 8578 2635 8597
rect 2635 8578 2699 8597
rect 2699 8578 2706 8597
rect 2792 8578 2799 8597
rect 2799 8578 2863 8597
rect 2863 8578 2881 8597
rect 2881 8578 2945 8597
rect 2945 8578 2963 8597
rect 2963 8578 3027 8597
rect 3027 8578 3028 8597
rect 3114 8578 3127 8597
rect 3127 8578 3191 8597
rect 3191 8578 3209 8597
rect 3209 8578 3273 8597
rect 3273 8578 3290 8597
rect 3290 8578 3350 8597
rect 3436 8578 3452 8597
rect 3452 8578 3516 8597
rect 3516 8578 3533 8597
rect 3533 8578 3597 8597
rect 3597 8578 3614 8597
rect 3614 8578 3672 8597
rect 3758 8578 3759 8597
rect 3759 8578 3776 8597
rect 3776 8578 3840 8597
rect 3840 8578 3857 8597
rect 3857 8578 3921 8597
rect 3921 8578 3938 8597
rect 3938 8578 3994 8597
rect 4080 8578 4083 8597
rect 4083 8578 4100 8597
rect 4100 8578 4164 8597
rect 4164 8578 4181 8597
rect 4181 8578 4245 8597
rect 4245 8578 4262 8597
rect 4262 8578 4316 8597
rect 4402 8578 4407 8597
rect 4407 8578 4424 8597
rect 4424 8578 4488 8597
rect 4488 8578 4505 8597
rect 4505 8578 4569 8597
rect 4569 8578 4638 8597
rect 4724 8578 4759 8597
rect 4759 8578 4777 8597
rect 4777 8578 4841 8597
rect 4841 8578 4859 8597
rect 4859 8578 4923 8597
rect 4923 8578 4941 8597
rect 4941 8578 4960 8597
rect 5046 8578 5087 8597
rect 5087 8578 5105 8597
rect 5105 8578 5169 8597
rect 5169 8578 5187 8597
rect 5187 8578 5251 8597
rect 5251 8578 5269 8597
rect 5269 8578 5282 8597
rect 5368 8578 5415 8597
rect 5415 8578 5433 8597
rect 5433 8578 5497 8597
rect 5497 8578 5515 8597
rect 5515 8578 5579 8597
rect 5579 8578 5597 8597
rect 5597 8578 5604 8597
rect 5690 8578 5743 8597
rect 5743 8578 5760 8597
rect 5760 8578 5824 8597
rect 5824 8578 5841 8597
rect 5841 8578 5905 8597
rect 5905 8578 5922 8597
rect 5922 8578 5926 8597
rect 6012 8578 6067 8597
rect 6067 8578 6084 8597
rect 6084 8578 6148 8597
rect 6148 8578 6165 8597
rect 6165 8578 6229 8597
rect 6229 8578 6246 8597
rect 6246 8578 6248 8597
rect 6333 8578 6391 8597
rect 6391 8578 6408 8597
rect 6408 8578 6472 8597
rect 6472 8578 6489 8597
rect 6489 8578 6553 8597
rect 6553 8578 6569 8597
rect 6654 8578 6715 8597
rect 6715 8578 6732 8597
rect 6732 8578 6796 8597
rect 6796 8578 6813 8597
rect 6813 8578 6877 8597
rect 6877 8578 6890 8597
rect 6975 8578 7039 8597
rect 7039 8578 7056 8597
rect 7056 8578 7120 8597
rect 7120 8578 7137 8597
rect 7137 8578 7201 8597
rect 7201 8578 7211 8597
rect 7296 8578 7299 8597
rect 7299 8578 7363 8597
rect 7363 8578 7380 8597
rect 7380 8578 7444 8597
rect 7444 8578 7461 8597
rect 7461 8578 7525 8597
rect 7525 8578 7532 8597
rect 7617 8578 7623 8597
rect 7623 8578 7687 8597
rect 7687 8581 7813 8597
rect 7813 8581 7853 8597
rect 7938 8581 7961 8597
rect 7961 8581 7981 8597
rect 7981 8581 8045 8597
rect 8045 8581 8065 8597
rect 8065 8581 8129 8597
rect 8129 8581 8149 8597
rect 8149 8581 8174 8597
rect 7687 8578 7853 8581
rect 216 8556 452 8578
rect 538 8556 774 8578
rect 860 8556 1096 8578
rect 1182 8556 1418 8578
rect 1504 8556 1740 8578
rect 1826 8556 2062 8578
rect 2148 8556 2384 8578
rect 2470 8556 2706 8578
rect 2792 8556 3028 8578
rect 3114 8556 3350 8578
rect 3436 8556 3672 8578
rect 3758 8556 3994 8578
rect 4080 8556 4316 8578
rect 4402 8556 4638 8578
rect 4724 8556 4960 8578
rect 5046 8556 5282 8578
rect 5368 8556 5604 8578
rect 5690 8556 5926 8578
rect 6012 8556 6248 8578
rect 6333 8556 6569 8578
rect 6654 8556 6890 8578
rect 6975 8556 7211 8578
rect 7296 8556 7532 8578
rect 7617 8559 7853 8578
rect 7938 8559 8174 8581
rect 7617 8556 7813 8559
rect 216 8492 397 8556
rect 397 8492 452 8556
rect 538 8492 543 8556
rect 543 8492 561 8556
rect 561 8492 625 8556
rect 625 8492 643 8556
rect 643 8492 707 8556
rect 707 8492 725 8556
rect 725 8492 774 8556
rect 860 8492 871 8556
rect 871 8492 889 8556
rect 889 8492 953 8556
rect 953 8492 971 8556
rect 971 8492 1035 8556
rect 1035 8492 1053 8556
rect 1053 8492 1096 8556
rect 1182 8492 1199 8556
rect 1199 8492 1217 8556
rect 1217 8492 1281 8556
rect 1281 8492 1299 8556
rect 1299 8492 1363 8556
rect 1363 8492 1381 8556
rect 1381 8492 1418 8556
rect 1504 8492 1527 8556
rect 1527 8492 1545 8556
rect 1545 8492 1609 8556
rect 1609 8492 1627 8556
rect 1627 8492 1691 8556
rect 1691 8492 1709 8556
rect 1709 8492 1740 8556
rect 1826 8492 1855 8556
rect 1855 8492 1873 8556
rect 1873 8492 1937 8556
rect 1937 8492 1955 8556
rect 1955 8492 2019 8556
rect 2019 8492 2037 8556
rect 2037 8492 2062 8556
rect 2148 8492 2183 8556
rect 2183 8492 2201 8556
rect 2201 8492 2265 8556
rect 2265 8492 2282 8556
rect 2282 8492 2346 8556
rect 2346 8492 2363 8556
rect 2363 8492 2384 8556
rect 2470 8492 2553 8556
rect 2553 8492 2617 8556
rect 2617 8492 2635 8556
rect 2635 8492 2699 8556
rect 2699 8492 2706 8556
rect 2792 8492 2799 8556
rect 2799 8492 2863 8556
rect 2863 8492 2881 8556
rect 2881 8492 2945 8556
rect 2945 8492 2963 8556
rect 2963 8492 3027 8556
rect 3027 8492 3028 8556
rect 3114 8492 3127 8556
rect 3127 8492 3191 8556
rect 3191 8492 3209 8556
rect 3209 8492 3273 8556
rect 3273 8492 3290 8556
rect 3290 8492 3350 8556
rect 3436 8492 3452 8556
rect 3452 8492 3516 8556
rect 3516 8492 3533 8556
rect 3533 8492 3597 8556
rect 3597 8492 3614 8556
rect 3614 8492 3672 8556
rect 3758 8492 3759 8556
rect 3759 8492 3776 8556
rect 3776 8492 3840 8556
rect 3840 8492 3857 8556
rect 3857 8492 3921 8556
rect 3921 8492 3938 8556
rect 3938 8492 3994 8556
rect 4080 8492 4083 8556
rect 4083 8492 4100 8556
rect 4100 8492 4164 8556
rect 4164 8492 4181 8556
rect 4181 8492 4245 8556
rect 4245 8492 4262 8556
rect 4262 8492 4316 8556
rect 4402 8492 4407 8556
rect 4407 8492 4424 8556
rect 4424 8492 4488 8556
rect 4488 8492 4505 8556
rect 4505 8492 4569 8556
rect 4569 8492 4638 8556
rect 4724 8492 4759 8556
rect 4759 8492 4777 8556
rect 4777 8492 4841 8556
rect 4841 8492 4859 8556
rect 4859 8492 4923 8556
rect 4923 8492 4941 8556
rect 4941 8492 4960 8556
rect 5046 8492 5087 8556
rect 5087 8492 5105 8556
rect 5105 8492 5169 8556
rect 5169 8492 5187 8556
rect 5187 8492 5251 8556
rect 5251 8492 5269 8556
rect 5269 8492 5282 8556
rect 5368 8492 5415 8556
rect 5415 8492 5433 8556
rect 5433 8492 5497 8556
rect 5497 8492 5515 8556
rect 5515 8492 5579 8556
rect 5579 8492 5597 8556
rect 5597 8492 5604 8556
rect 5690 8492 5743 8556
rect 5743 8492 5760 8556
rect 5760 8492 5824 8556
rect 5824 8492 5841 8556
rect 5841 8492 5905 8556
rect 5905 8492 5922 8556
rect 5922 8492 5926 8556
rect 6012 8492 6067 8556
rect 6067 8492 6084 8556
rect 6084 8492 6148 8556
rect 6148 8492 6165 8556
rect 6165 8492 6229 8556
rect 6229 8492 6246 8556
rect 6246 8492 6248 8556
rect 6333 8492 6391 8556
rect 6391 8492 6408 8556
rect 6408 8492 6472 8556
rect 6472 8492 6489 8556
rect 6489 8492 6553 8556
rect 6553 8492 6569 8556
rect 6654 8492 6715 8556
rect 6715 8492 6732 8556
rect 6732 8492 6796 8556
rect 6796 8492 6813 8556
rect 6813 8492 6877 8556
rect 6877 8492 6890 8556
rect 6975 8492 7039 8556
rect 7039 8492 7056 8556
rect 7056 8492 7120 8556
rect 7120 8492 7137 8556
rect 7137 8492 7201 8556
rect 7201 8492 7211 8556
rect 7296 8492 7299 8556
rect 7299 8492 7363 8556
rect 7363 8492 7380 8556
rect 7380 8492 7444 8556
rect 7444 8492 7461 8556
rect 7461 8492 7525 8556
rect 7525 8492 7532 8556
rect 7617 8492 7623 8556
rect 7623 8492 7687 8556
rect 7687 8495 7813 8556
rect 7813 8495 7853 8559
rect 7938 8495 7961 8559
rect 7961 8495 7981 8559
rect 7981 8495 8045 8559
rect 8045 8495 8065 8559
rect 8065 8495 8129 8559
rect 8129 8495 8149 8559
rect 8149 8495 8174 8559
rect 7687 8492 7853 8495
rect 216 8470 452 8492
rect 538 8470 774 8492
rect 860 8470 1096 8492
rect 1182 8470 1418 8492
rect 1504 8470 1740 8492
rect 1826 8470 2062 8492
rect 2148 8470 2384 8492
rect 2470 8470 2706 8492
rect 2792 8470 3028 8492
rect 3114 8470 3350 8492
rect 3436 8470 3672 8492
rect 3758 8470 3994 8492
rect 4080 8470 4316 8492
rect 4402 8470 4638 8492
rect 4724 8470 4960 8492
rect 5046 8470 5282 8492
rect 5368 8470 5604 8492
rect 5690 8470 5926 8492
rect 6012 8470 6248 8492
rect 6333 8470 6569 8492
rect 6654 8470 6890 8492
rect 6975 8470 7211 8492
rect 7296 8470 7532 8492
rect 7617 8473 7853 8492
rect 7938 8473 8174 8495
rect 7617 8470 7813 8473
rect 216 8406 397 8470
rect 397 8406 452 8470
rect 538 8406 543 8470
rect 543 8406 561 8470
rect 561 8406 625 8470
rect 625 8406 643 8470
rect 643 8406 707 8470
rect 707 8406 725 8470
rect 725 8406 774 8470
rect 860 8406 871 8470
rect 871 8406 889 8470
rect 889 8406 953 8470
rect 953 8406 971 8470
rect 971 8406 1035 8470
rect 1035 8406 1053 8470
rect 1053 8406 1096 8470
rect 1182 8406 1199 8470
rect 1199 8406 1217 8470
rect 1217 8406 1281 8470
rect 1281 8406 1299 8470
rect 1299 8406 1363 8470
rect 1363 8406 1381 8470
rect 1381 8406 1418 8470
rect 1504 8406 1527 8470
rect 1527 8406 1545 8470
rect 1545 8406 1609 8470
rect 1609 8406 1627 8470
rect 1627 8406 1691 8470
rect 1691 8406 1709 8470
rect 1709 8406 1740 8470
rect 1826 8406 1855 8470
rect 1855 8406 1873 8470
rect 1873 8406 1937 8470
rect 1937 8406 1955 8470
rect 1955 8406 2019 8470
rect 2019 8406 2037 8470
rect 2037 8406 2062 8470
rect 2148 8406 2183 8470
rect 2183 8406 2201 8470
rect 2201 8406 2265 8470
rect 2265 8406 2282 8470
rect 2282 8406 2346 8470
rect 2346 8406 2363 8470
rect 2363 8406 2384 8470
rect 2470 8406 2553 8470
rect 2553 8406 2617 8470
rect 2617 8406 2635 8470
rect 2635 8406 2699 8470
rect 2699 8406 2706 8470
rect 2792 8406 2799 8470
rect 2799 8406 2863 8470
rect 2863 8406 2881 8470
rect 2881 8406 2945 8470
rect 2945 8406 2963 8470
rect 2963 8406 3027 8470
rect 3027 8406 3028 8470
rect 3114 8406 3127 8470
rect 3127 8406 3191 8470
rect 3191 8406 3209 8470
rect 3209 8406 3273 8470
rect 3273 8406 3290 8470
rect 3290 8406 3350 8470
rect 3436 8406 3452 8470
rect 3452 8406 3516 8470
rect 3516 8406 3533 8470
rect 3533 8406 3597 8470
rect 3597 8406 3614 8470
rect 3614 8406 3672 8470
rect 3758 8406 3759 8470
rect 3759 8406 3776 8470
rect 3776 8406 3840 8470
rect 3840 8406 3857 8470
rect 3857 8406 3921 8470
rect 3921 8406 3938 8470
rect 3938 8406 3994 8470
rect 4080 8406 4083 8470
rect 4083 8406 4100 8470
rect 4100 8406 4164 8470
rect 4164 8406 4181 8470
rect 4181 8406 4245 8470
rect 4245 8406 4262 8470
rect 4262 8406 4316 8470
rect 4402 8406 4407 8470
rect 4407 8406 4424 8470
rect 4424 8406 4488 8470
rect 4488 8406 4505 8470
rect 4505 8406 4569 8470
rect 4569 8406 4638 8470
rect 4724 8406 4759 8470
rect 4759 8406 4777 8470
rect 4777 8406 4841 8470
rect 4841 8406 4859 8470
rect 4859 8406 4923 8470
rect 4923 8406 4941 8470
rect 4941 8406 4960 8470
rect 5046 8406 5087 8470
rect 5087 8406 5105 8470
rect 5105 8406 5169 8470
rect 5169 8406 5187 8470
rect 5187 8406 5251 8470
rect 5251 8406 5269 8470
rect 5269 8406 5282 8470
rect 5368 8406 5415 8470
rect 5415 8406 5433 8470
rect 5433 8406 5497 8470
rect 5497 8406 5515 8470
rect 5515 8406 5579 8470
rect 5579 8406 5597 8470
rect 5597 8406 5604 8470
rect 5690 8406 5743 8470
rect 5743 8406 5760 8470
rect 5760 8406 5824 8470
rect 5824 8406 5841 8470
rect 5841 8406 5905 8470
rect 5905 8406 5922 8470
rect 5922 8406 5926 8470
rect 6012 8406 6067 8470
rect 6067 8406 6084 8470
rect 6084 8406 6148 8470
rect 6148 8406 6165 8470
rect 6165 8406 6229 8470
rect 6229 8406 6246 8470
rect 6246 8406 6248 8470
rect 6333 8406 6391 8470
rect 6391 8406 6408 8470
rect 6408 8406 6472 8470
rect 6472 8406 6489 8470
rect 6489 8406 6553 8470
rect 6553 8406 6569 8470
rect 6654 8406 6715 8470
rect 6715 8406 6732 8470
rect 6732 8406 6796 8470
rect 6796 8406 6813 8470
rect 6813 8406 6877 8470
rect 6877 8406 6890 8470
rect 6975 8406 7039 8470
rect 7039 8406 7056 8470
rect 7056 8406 7120 8470
rect 7120 8406 7137 8470
rect 7137 8406 7201 8470
rect 7201 8406 7211 8470
rect 7296 8406 7299 8470
rect 7299 8406 7363 8470
rect 7363 8406 7380 8470
rect 7380 8406 7444 8470
rect 7444 8406 7461 8470
rect 7461 8406 7525 8470
rect 7525 8406 7532 8470
rect 7617 8406 7623 8470
rect 7623 8406 7687 8470
rect 7687 8409 7813 8470
rect 7813 8409 7853 8473
rect 7938 8409 7961 8473
rect 7961 8409 7981 8473
rect 7981 8409 8045 8473
rect 8045 8409 8065 8473
rect 8065 8409 8129 8473
rect 8129 8409 8149 8473
rect 8149 8409 8174 8473
rect 7687 8406 7853 8409
rect 216 8384 452 8406
rect 538 8384 774 8406
rect 860 8384 1096 8406
rect 1182 8384 1418 8406
rect 1504 8384 1740 8406
rect 1826 8384 2062 8406
rect 2148 8384 2384 8406
rect 2470 8384 2706 8406
rect 2792 8384 3028 8406
rect 3114 8384 3350 8406
rect 3436 8384 3672 8406
rect 3758 8384 3994 8406
rect 4080 8384 4316 8406
rect 4402 8384 4638 8406
rect 4724 8384 4960 8406
rect 5046 8384 5282 8406
rect 5368 8384 5604 8406
rect 5690 8384 5926 8406
rect 6012 8384 6248 8406
rect 6333 8384 6569 8406
rect 6654 8384 6890 8406
rect 6975 8384 7211 8406
rect 7296 8384 7532 8406
rect 7617 8387 7853 8406
rect 7938 8387 8174 8409
rect 7617 8384 7813 8387
rect 216 8361 397 8384
rect 397 8361 452 8384
rect 538 8361 543 8384
rect 543 8361 561 8384
rect 561 8361 625 8384
rect 625 8361 643 8384
rect 643 8361 707 8384
rect 707 8361 725 8384
rect 725 8361 774 8384
rect 860 8361 871 8384
rect 871 8361 889 8384
rect 889 8361 953 8384
rect 953 8361 971 8384
rect 971 8361 1035 8384
rect 1035 8361 1053 8384
rect 1053 8361 1096 8384
rect 1182 8361 1199 8384
rect 1199 8361 1217 8384
rect 1217 8361 1281 8384
rect 1281 8361 1299 8384
rect 1299 8361 1363 8384
rect 1363 8361 1381 8384
rect 1381 8361 1418 8384
rect 1504 8361 1527 8384
rect 1527 8361 1545 8384
rect 1545 8361 1609 8384
rect 1609 8361 1627 8384
rect 1627 8361 1691 8384
rect 1691 8361 1709 8384
rect 1709 8361 1740 8384
rect 1826 8361 1855 8384
rect 1855 8361 1873 8384
rect 1873 8361 1937 8384
rect 1937 8361 1955 8384
rect 1955 8361 2019 8384
rect 2019 8361 2037 8384
rect 2037 8361 2062 8384
rect 2148 8361 2183 8384
rect 2183 8361 2201 8384
rect 2201 8361 2265 8384
rect 2265 8361 2282 8384
rect 2282 8361 2346 8384
rect 2346 8361 2363 8384
rect 2363 8361 2384 8384
rect 2470 8361 2553 8384
rect 2553 8361 2617 8384
rect 2617 8361 2635 8384
rect 2635 8361 2699 8384
rect 2699 8361 2706 8384
rect 2792 8361 2799 8384
rect 2799 8361 2863 8384
rect 2863 8361 2881 8384
rect 2881 8361 2945 8384
rect 2945 8361 2963 8384
rect 2963 8361 3027 8384
rect 3027 8361 3028 8384
rect 3114 8361 3127 8384
rect 3127 8361 3191 8384
rect 3191 8361 3209 8384
rect 3209 8361 3273 8384
rect 3273 8361 3290 8384
rect 3290 8361 3350 8384
rect 3436 8361 3452 8384
rect 3452 8361 3516 8384
rect 3516 8361 3533 8384
rect 3533 8361 3597 8384
rect 3597 8361 3614 8384
rect 3614 8361 3672 8384
rect 3758 8361 3759 8384
rect 3759 8361 3776 8384
rect 3776 8361 3840 8384
rect 3840 8361 3857 8384
rect 3857 8361 3921 8384
rect 3921 8361 3938 8384
rect 3938 8361 3994 8384
rect 4080 8361 4083 8384
rect 4083 8361 4100 8384
rect 4100 8361 4164 8384
rect 4164 8361 4181 8384
rect 4181 8361 4245 8384
rect 4245 8361 4262 8384
rect 4262 8361 4316 8384
rect 4402 8361 4407 8384
rect 4407 8361 4424 8384
rect 4424 8361 4488 8384
rect 4488 8361 4505 8384
rect 4505 8361 4569 8384
rect 4569 8361 4638 8384
rect 4724 8361 4759 8384
rect 4759 8361 4777 8384
rect 4777 8361 4841 8384
rect 4841 8361 4859 8384
rect 4859 8361 4923 8384
rect 4923 8361 4941 8384
rect 4941 8361 4960 8384
rect 5046 8361 5087 8384
rect 5087 8361 5105 8384
rect 5105 8361 5169 8384
rect 5169 8361 5187 8384
rect 5187 8361 5251 8384
rect 5251 8361 5269 8384
rect 5269 8361 5282 8384
rect 5368 8361 5415 8384
rect 5415 8361 5433 8384
rect 5433 8361 5497 8384
rect 5497 8361 5515 8384
rect 5515 8361 5579 8384
rect 5579 8361 5597 8384
rect 5597 8361 5604 8384
rect 5690 8361 5743 8384
rect 5743 8361 5760 8384
rect 5760 8361 5824 8384
rect 5824 8361 5841 8384
rect 5841 8361 5905 8384
rect 5905 8361 5922 8384
rect 5922 8361 5926 8384
rect 6012 8361 6067 8384
rect 6067 8361 6084 8384
rect 6084 8361 6148 8384
rect 6148 8361 6165 8384
rect 6165 8361 6229 8384
rect 6229 8361 6246 8384
rect 6246 8361 6248 8384
rect 6333 8361 6391 8384
rect 6391 8361 6408 8384
rect 6408 8361 6472 8384
rect 6472 8361 6489 8384
rect 6489 8361 6553 8384
rect 6553 8361 6569 8384
rect 6654 8361 6715 8384
rect 6715 8361 6732 8384
rect 6732 8361 6796 8384
rect 6796 8361 6813 8384
rect 6813 8361 6877 8384
rect 6877 8361 6890 8384
rect 6975 8361 7039 8384
rect 7039 8361 7056 8384
rect 7056 8361 7120 8384
rect 7120 8361 7137 8384
rect 7137 8361 7201 8384
rect 7201 8361 7211 8384
rect 7296 8361 7299 8384
rect 7299 8361 7363 8384
rect 7363 8361 7380 8384
rect 7380 8361 7444 8384
rect 7444 8361 7461 8384
rect 7461 8361 7525 8384
rect 7525 8361 7532 8384
rect 7617 8361 7623 8384
rect 7623 8361 7687 8384
rect 7687 8361 7813 8384
rect 7813 8361 7853 8387
rect 7938 8361 7961 8387
rect 7961 8361 7981 8387
rect 7981 8361 8045 8387
rect 8045 8361 8065 8387
rect 8065 8361 8129 8387
rect 8129 8361 8149 8387
rect 8149 8361 8174 8387
rect 8259 8361 8495 8597
rect 8580 8361 8816 8597
rect 8901 8578 8923 8597
rect 8923 8578 8940 8597
rect 8940 8578 9004 8597
rect 9004 8578 9021 8597
rect 9021 8578 9085 8597
rect 9085 8578 9102 8597
rect 9102 8578 9137 8597
rect 9222 8578 9247 8597
rect 9247 8578 9264 8597
rect 9264 8578 9328 8597
rect 9328 8578 9345 8597
rect 9345 8578 9409 8597
rect 9409 8578 9426 8597
rect 9426 8578 9458 8597
rect 9543 8578 9571 8597
rect 9571 8578 9588 8597
rect 9588 8578 9652 8597
rect 9652 8578 9669 8597
rect 9669 8578 9733 8597
rect 9733 8578 9750 8597
rect 9750 8578 9779 8597
rect 9864 8578 9895 8597
rect 9895 8578 9912 8597
rect 9912 8578 9976 8597
rect 9976 8578 9993 8597
rect 9993 8578 10057 8597
rect 10057 8578 10073 8597
rect 10073 8578 10100 8597
rect 10185 8578 10217 8597
rect 10217 8578 10233 8597
rect 10233 8578 10297 8597
rect 10297 8578 10313 8597
rect 10313 8578 10377 8597
rect 10377 8578 10393 8597
rect 10393 8578 10421 8597
rect 10506 8578 10537 8597
rect 10537 8578 10553 8597
rect 10553 8578 10617 8597
rect 10617 8578 10633 8597
rect 10633 8578 10697 8597
rect 10697 8578 10713 8597
rect 10713 8578 10742 8597
rect 10827 8578 10857 8597
rect 10857 8578 10873 8597
rect 10873 8578 10937 8597
rect 10937 8578 10953 8597
rect 10953 8578 11017 8597
rect 11017 8578 11033 8597
rect 11033 8578 11063 8597
rect 11148 8578 11177 8597
rect 11177 8578 11193 8597
rect 11193 8578 11257 8597
rect 11257 8578 11273 8597
rect 11273 8578 11337 8597
rect 11337 8578 11353 8597
rect 11353 8578 11384 8597
rect 11469 8578 11497 8597
rect 11497 8578 11513 8597
rect 11513 8578 11577 8597
rect 11577 8578 11593 8597
rect 11593 8578 11657 8597
rect 11657 8578 11673 8597
rect 11673 8578 11705 8597
rect 11790 8578 11817 8597
rect 11817 8578 11833 8597
rect 11833 8578 11897 8597
rect 11897 8578 11913 8597
rect 11913 8578 11977 8597
rect 11977 8578 12026 8597
rect 8901 8556 9137 8578
rect 9222 8556 9458 8578
rect 9543 8556 9779 8578
rect 9864 8556 10100 8578
rect 10185 8556 10421 8578
rect 10506 8556 10742 8578
rect 10827 8556 11063 8578
rect 11148 8556 11384 8578
rect 11469 8556 11705 8578
rect 11790 8556 12026 8578
rect 8901 8492 8923 8556
rect 8923 8492 8940 8556
rect 8940 8492 9004 8556
rect 9004 8492 9021 8556
rect 9021 8492 9085 8556
rect 9085 8492 9102 8556
rect 9102 8492 9137 8556
rect 9222 8492 9247 8556
rect 9247 8492 9264 8556
rect 9264 8492 9328 8556
rect 9328 8492 9345 8556
rect 9345 8492 9409 8556
rect 9409 8492 9426 8556
rect 9426 8492 9458 8556
rect 9543 8492 9571 8556
rect 9571 8492 9588 8556
rect 9588 8492 9652 8556
rect 9652 8492 9669 8556
rect 9669 8492 9733 8556
rect 9733 8492 9750 8556
rect 9750 8492 9779 8556
rect 9864 8492 9895 8556
rect 9895 8492 9912 8556
rect 9912 8492 9976 8556
rect 9976 8492 9993 8556
rect 9993 8492 10057 8556
rect 10057 8492 10073 8556
rect 10073 8492 10100 8556
rect 10185 8492 10217 8556
rect 10217 8492 10233 8556
rect 10233 8492 10297 8556
rect 10297 8492 10313 8556
rect 10313 8492 10377 8556
rect 10377 8492 10393 8556
rect 10393 8492 10421 8556
rect 10506 8492 10537 8556
rect 10537 8492 10553 8556
rect 10553 8492 10617 8556
rect 10617 8492 10633 8556
rect 10633 8492 10697 8556
rect 10697 8492 10713 8556
rect 10713 8492 10742 8556
rect 10827 8492 10857 8556
rect 10857 8492 10873 8556
rect 10873 8492 10937 8556
rect 10937 8492 10953 8556
rect 10953 8492 11017 8556
rect 11017 8492 11033 8556
rect 11033 8492 11063 8556
rect 11148 8492 11177 8556
rect 11177 8492 11193 8556
rect 11193 8492 11257 8556
rect 11257 8492 11273 8556
rect 11273 8492 11337 8556
rect 11337 8492 11353 8556
rect 11353 8492 11384 8556
rect 11469 8492 11497 8556
rect 11497 8492 11513 8556
rect 11513 8492 11577 8556
rect 11577 8492 11593 8556
rect 11593 8492 11657 8556
rect 11657 8492 11673 8556
rect 11673 8492 11705 8556
rect 11790 8492 11817 8556
rect 11817 8492 11833 8556
rect 11833 8492 11897 8556
rect 11897 8492 11913 8556
rect 11913 8492 11977 8556
rect 11977 8492 12026 8556
rect 8901 8470 9137 8492
rect 9222 8470 9458 8492
rect 9543 8470 9779 8492
rect 9864 8470 10100 8492
rect 10185 8470 10421 8492
rect 10506 8470 10742 8492
rect 10827 8470 11063 8492
rect 11148 8470 11384 8492
rect 11469 8470 11705 8492
rect 11790 8470 12026 8492
rect 8901 8406 8923 8470
rect 8923 8406 8940 8470
rect 8940 8406 9004 8470
rect 9004 8406 9021 8470
rect 9021 8406 9085 8470
rect 9085 8406 9102 8470
rect 9102 8406 9137 8470
rect 9222 8406 9247 8470
rect 9247 8406 9264 8470
rect 9264 8406 9328 8470
rect 9328 8406 9345 8470
rect 9345 8406 9409 8470
rect 9409 8406 9426 8470
rect 9426 8406 9458 8470
rect 9543 8406 9571 8470
rect 9571 8406 9588 8470
rect 9588 8406 9652 8470
rect 9652 8406 9669 8470
rect 9669 8406 9733 8470
rect 9733 8406 9750 8470
rect 9750 8406 9779 8470
rect 9864 8406 9895 8470
rect 9895 8406 9912 8470
rect 9912 8406 9976 8470
rect 9976 8406 9993 8470
rect 9993 8406 10057 8470
rect 10057 8406 10073 8470
rect 10073 8406 10100 8470
rect 10185 8406 10217 8470
rect 10217 8406 10233 8470
rect 10233 8406 10297 8470
rect 10297 8406 10313 8470
rect 10313 8406 10377 8470
rect 10377 8406 10393 8470
rect 10393 8406 10421 8470
rect 10506 8406 10537 8470
rect 10537 8406 10553 8470
rect 10553 8406 10617 8470
rect 10617 8406 10633 8470
rect 10633 8406 10697 8470
rect 10697 8406 10713 8470
rect 10713 8406 10742 8470
rect 10827 8406 10857 8470
rect 10857 8406 10873 8470
rect 10873 8406 10937 8470
rect 10937 8406 10953 8470
rect 10953 8406 11017 8470
rect 11017 8406 11033 8470
rect 11033 8406 11063 8470
rect 11148 8406 11177 8470
rect 11177 8406 11193 8470
rect 11193 8406 11257 8470
rect 11257 8406 11273 8470
rect 11273 8406 11337 8470
rect 11337 8406 11353 8470
rect 11353 8406 11384 8470
rect 11469 8406 11497 8470
rect 11497 8406 11513 8470
rect 11513 8406 11577 8470
rect 11577 8406 11593 8470
rect 11593 8406 11657 8470
rect 11657 8406 11673 8470
rect 11673 8406 11705 8470
rect 11790 8406 11817 8470
rect 11817 8406 11833 8470
rect 11833 8406 11897 8470
rect 11897 8406 11913 8470
rect 11913 8406 11977 8470
rect 11977 8406 12026 8470
rect 8901 8384 9137 8406
rect 9222 8384 9458 8406
rect 9543 8384 9779 8406
rect 9864 8384 10100 8406
rect 10185 8384 10421 8406
rect 10506 8384 10742 8406
rect 10827 8384 11063 8406
rect 11148 8384 11384 8406
rect 11469 8384 11705 8406
rect 11790 8384 12026 8406
rect 8901 8361 8923 8384
rect 8923 8361 8940 8384
rect 8940 8361 9004 8384
rect 9004 8361 9021 8384
rect 9021 8361 9085 8384
rect 9085 8361 9102 8384
rect 9102 8361 9137 8384
rect 9222 8361 9247 8384
rect 9247 8361 9264 8384
rect 9264 8361 9328 8384
rect 9328 8361 9345 8384
rect 9345 8361 9409 8384
rect 9409 8361 9426 8384
rect 9426 8361 9458 8384
rect 9543 8361 9571 8384
rect 9571 8361 9588 8384
rect 9588 8361 9652 8384
rect 9652 8361 9669 8384
rect 9669 8361 9733 8384
rect 9733 8361 9750 8384
rect 9750 8361 9779 8384
rect 9864 8361 9895 8384
rect 9895 8361 9912 8384
rect 9912 8361 9976 8384
rect 9976 8361 9993 8384
rect 9993 8361 10057 8384
rect 10057 8361 10073 8384
rect 10073 8361 10100 8384
rect 10185 8361 10217 8384
rect 10217 8361 10233 8384
rect 10233 8361 10297 8384
rect 10297 8361 10313 8384
rect 10313 8361 10377 8384
rect 10377 8361 10393 8384
rect 10393 8361 10421 8384
rect 10506 8361 10537 8384
rect 10537 8361 10553 8384
rect 10553 8361 10617 8384
rect 10617 8361 10633 8384
rect 10633 8361 10697 8384
rect 10697 8361 10713 8384
rect 10713 8361 10742 8384
rect 10827 8361 10857 8384
rect 10857 8361 10873 8384
rect 10873 8361 10937 8384
rect 10937 8361 10953 8384
rect 10953 8361 11017 8384
rect 11017 8361 11033 8384
rect 11033 8361 11063 8384
rect 11148 8361 11177 8384
rect 11177 8361 11193 8384
rect 11193 8361 11257 8384
rect 11257 8361 11273 8384
rect 11273 8361 11337 8384
rect 11337 8361 11353 8384
rect 11353 8361 11384 8384
rect 11469 8361 11497 8384
rect 11497 8361 11513 8384
rect 11513 8361 11577 8384
rect 11577 8361 11593 8384
rect 11593 8361 11657 8384
rect 11657 8361 11673 8384
rect 11673 8361 11705 8384
rect 11790 8361 11817 8384
rect 11817 8361 11833 8384
rect 11833 8361 11897 8384
rect 11897 8361 11913 8384
rect 11913 8361 11977 8384
rect 11977 8361 12026 8384
rect 12111 8578 12165 8597
rect 12165 8578 12229 8597
rect 12229 8578 12246 8597
rect 12246 8578 12310 8597
rect 12310 8578 12327 8597
rect 12327 8578 12347 8597
rect 12432 8578 12472 8597
rect 12472 8578 12489 8597
rect 12489 8578 12553 8597
rect 12553 8578 12570 8597
rect 12570 8578 12634 8597
rect 12634 8578 12651 8597
rect 12651 8578 12668 8597
rect 12753 8578 12796 8597
rect 12796 8578 12813 8597
rect 12813 8578 12877 8597
rect 12877 8578 12894 8597
rect 12894 8578 12958 8597
rect 12958 8578 12975 8597
rect 12975 8578 12989 8597
rect 13074 8578 13120 8597
rect 13120 8578 13137 8597
rect 13137 8578 13201 8597
rect 13201 8578 13218 8597
rect 13218 8578 13282 8597
rect 13282 8578 13299 8597
rect 13299 8578 13310 8597
rect 13395 8578 13444 8597
rect 13444 8578 13461 8597
rect 13461 8578 13525 8597
rect 13525 8578 13542 8597
rect 13542 8578 13606 8597
rect 13606 8578 13623 8597
rect 13623 8578 13631 8597
rect 13716 8578 13768 8597
rect 13768 8578 13785 8597
rect 13785 8578 13849 8597
rect 13849 8578 13866 8597
rect 13866 8578 13930 8597
rect 13930 8578 13947 8597
rect 13947 8578 13952 8597
rect 14037 8578 14092 8597
rect 14092 8578 14109 8597
rect 14109 8578 14173 8597
rect 14173 8578 14190 8597
rect 14190 8578 14254 8597
rect 14254 8578 14271 8597
rect 14271 8578 14273 8597
rect 14358 8578 14416 8597
rect 14416 8578 14433 8597
rect 14433 8578 14497 8597
rect 14497 8578 14513 8597
rect 14513 8578 14577 8597
rect 14577 8578 14593 8597
rect 14593 8578 14594 8597
rect 14679 8578 14737 8597
rect 14737 8578 14753 8597
rect 14753 8578 14817 8597
rect 14817 8578 14833 8597
rect 14833 8578 14897 8597
rect 14897 8578 14913 8597
rect 14913 8578 14915 8597
rect 15000 8578 15057 8597
rect 15057 8578 15073 8597
rect 15073 8578 15137 8597
rect 15137 8578 15153 8597
rect 15153 8578 15217 8597
rect 15217 8578 15233 8597
rect 15233 8578 15236 8597
rect 15321 8578 15377 8597
rect 15377 8578 15393 8597
rect 15393 8578 15457 8597
rect 15457 8578 15473 8597
rect 15473 8578 15537 8597
rect 15537 8578 15553 8597
rect 15553 8578 15557 8597
rect 12111 8556 12347 8578
rect 12432 8556 12668 8578
rect 12753 8556 12989 8578
rect 13074 8556 13310 8578
rect 13395 8556 13631 8578
rect 13716 8556 13952 8578
rect 14037 8556 14273 8578
rect 14358 8556 14594 8578
rect 14679 8556 14915 8578
rect 15000 8556 15236 8578
rect 15321 8556 15557 8578
rect 12111 8492 12165 8556
rect 12165 8492 12229 8556
rect 12229 8492 12246 8556
rect 12246 8492 12310 8556
rect 12310 8492 12327 8556
rect 12327 8492 12347 8556
rect 12432 8492 12472 8556
rect 12472 8492 12489 8556
rect 12489 8492 12553 8556
rect 12553 8492 12570 8556
rect 12570 8492 12634 8556
rect 12634 8492 12651 8556
rect 12651 8492 12668 8556
rect 12753 8492 12796 8556
rect 12796 8492 12813 8556
rect 12813 8492 12877 8556
rect 12877 8492 12894 8556
rect 12894 8492 12958 8556
rect 12958 8492 12975 8556
rect 12975 8492 12989 8556
rect 13074 8492 13120 8556
rect 13120 8492 13137 8556
rect 13137 8492 13201 8556
rect 13201 8492 13218 8556
rect 13218 8492 13282 8556
rect 13282 8492 13299 8556
rect 13299 8492 13310 8556
rect 13395 8492 13444 8556
rect 13444 8492 13461 8556
rect 13461 8492 13525 8556
rect 13525 8492 13542 8556
rect 13542 8492 13606 8556
rect 13606 8492 13623 8556
rect 13623 8492 13631 8556
rect 13716 8492 13768 8556
rect 13768 8492 13785 8556
rect 13785 8492 13849 8556
rect 13849 8492 13866 8556
rect 13866 8492 13930 8556
rect 13930 8492 13947 8556
rect 13947 8492 13952 8556
rect 14037 8492 14092 8556
rect 14092 8492 14109 8556
rect 14109 8492 14173 8556
rect 14173 8492 14190 8556
rect 14190 8492 14254 8556
rect 14254 8492 14271 8556
rect 14271 8492 14273 8556
rect 14358 8492 14416 8556
rect 14416 8492 14433 8556
rect 14433 8492 14497 8556
rect 14497 8492 14513 8556
rect 14513 8492 14577 8556
rect 14577 8492 14593 8556
rect 14593 8492 14594 8556
rect 14679 8492 14737 8556
rect 14737 8492 14753 8556
rect 14753 8492 14817 8556
rect 14817 8492 14833 8556
rect 14833 8492 14897 8556
rect 14897 8492 14913 8556
rect 14913 8492 14915 8556
rect 15000 8492 15057 8556
rect 15057 8492 15073 8556
rect 15073 8492 15137 8556
rect 15137 8492 15153 8556
rect 15153 8492 15217 8556
rect 15217 8492 15233 8556
rect 15233 8492 15236 8556
rect 15321 8492 15377 8556
rect 15377 8492 15393 8556
rect 15393 8492 15457 8556
rect 15457 8492 15473 8556
rect 15473 8492 15537 8556
rect 15537 8492 15553 8556
rect 15553 8492 15557 8556
rect 12111 8470 12347 8492
rect 12432 8470 12668 8492
rect 12753 8470 12989 8492
rect 13074 8470 13310 8492
rect 13395 8470 13631 8492
rect 13716 8470 13952 8492
rect 14037 8470 14273 8492
rect 14358 8470 14594 8492
rect 14679 8470 14915 8492
rect 15000 8470 15236 8492
rect 15321 8470 15557 8492
rect 12111 8406 12165 8470
rect 12165 8406 12229 8470
rect 12229 8406 12246 8470
rect 12246 8406 12310 8470
rect 12310 8406 12327 8470
rect 12327 8406 12347 8470
rect 12432 8406 12472 8470
rect 12472 8406 12489 8470
rect 12489 8406 12553 8470
rect 12553 8406 12570 8470
rect 12570 8406 12634 8470
rect 12634 8406 12651 8470
rect 12651 8406 12668 8470
rect 12753 8406 12796 8470
rect 12796 8406 12813 8470
rect 12813 8406 12877 8470
rect 12877 8406 12894 8470
rect 12894 8406 12958 8470
rect 12958 8406 12975 8470
rect 12975 8406 12989 8470
rect 13074 8406 13120 8470
rect 13120 8406 13137 8470
rect 13137 8406 13201 8470
rect 13201 8406 13218 8470
rect 13218 8406 13282 8470
rect 13282 8406 13299 8470
rect 13299 8406 13310 8470
rect 13395 8406 13444 8470
rect 13444 8406 13461 8470
rect 13461 8406 13525 8470
rect 13525 8406 13542 8470
rect 13542 8406 13606 8470
rect 13606 8406 13623 8470
rect 13623 8406 13631 8470
rect 13716 8406 13768 8470
rect 13768 8406 13785 8470
rect 13785 8406 13849 8470
rect 13849 8406 13866 8470
rect 13866 8406 13930 8470
rect 13930 8406 13947 8470
rect 13947 8406 13952 8470
rect 14037 8406 14092 8470
rect 14092 8406 14109 8470
rect 14109 8406 14173 8470
rect 14173 8406 14190 8470
rect 14190 8406 14254 8470
rect 14254 8406 14271 8470
rect 14271 8406 14273 8470
rect 14358 8406 14416 8470
rect 14416 8406 14433 8470
rect 14433 8406 14497 8470
rect 14497 8406 14513 8470
rect 14513 8406 14577 8470
rect 14577 8406 14593 8470
rect 14593 8406 14594 8470
rect 14679 8406 14737 8470
rect 14737 8406 14753 8470
rect 14753 8406 14817 8470
rect 14817 8406 14833 8470
rect 14833 8406 14897 8470
rect 14897 8406 14913 8470
rect 14913 8406 14915 8470
rect 15000 8406 15057 8470
rect 15057 8406 15073 8470
rect 15073 8406 15137 8470
rect 15137 8406 15153 8470
rect 15153 8406 15217 8470
rect 15217 8406 15233 8470
rect 15233 8406 15236 8470
rect 15321 8406 15377 8470
rect 15377 8406 15393 8470
rect 15393 8406 15457 8470
rect 15457 8406 15473 8470
rect 15473 8406 15537 8470
rect 15537 8406 15553 8470
rect 15553 8406 15557 8470
rect 12111 8384 12347 8406
rect 12432 8384 12668 8406
rect 12753 8384 12989 8406
rect 13074 8384 13310 8406
rect 13395 8384 13631 8406
rect 13716 8384 13952 8406
rect 14037 8384 14273 8406
rect 14358 8384 14594 8406
rect 14679 8384 14915 8406
rect 15000 8384 15236 8406
rect 15321 8384 15557 8406
rect 12111 8361 12165 8384
rect 12165 8361 12229 8384
rect 12229 8361 12246 8384
rect 12246 8361 12310 8384
rect 12310 8361 12327 8384
rect 12327 8361 12347 8384
rect 12432 8361 12472 8384
rect 12472 8361 12489 8384
rect 12489 8361 12553 8384
rect 12553 8361 12570 8384
rect 12570 8361 12634 8384
rect 12634 8361 12651 8384
rect 12651 8361 12668 8384
rect 12753 8361 12796 8384
rect 12796 8361 12813 8384
rect 12813 8361 12877 8384
rect 12877 8361 12894 8384
rect 12894 8361 12958 8384
rect 12958 8361 12975 8384
rect 12975 8361 12989 8384
rect 13074 8361 13120 8384
rect 13120 8361 13137 8384
rect 13137 8361 13201 8384
rect 13201 8361 13218 8384
rect 13218 8361 13282 8384
rect 13282 8361 13299 8384
rect 13299 8361 13310 8384
rect 13395 8361 13444 8384
rect 13444 8361 13461 8384
rect 13461 8361 13525 8384
rect 13525 8361 13542 8384
rect 13542 8361 13606 8384
rect 13606 8361 13623 8384
rect 13623 8361 13631 8384
rect 13716 8361 13768 8384
rect 13768 8361 13785 8384
rect 13785 8361 13849 8384
rect 13849 8361 13866 8384
rect 13866 8361 13930 8384
rect 13930 8361 13947 8384
rect 13947 8361 13952 8384
rect 14037 8361 14092 8384
rect 14092 8361 14109 8384
rect 14109 8361 14173 8384
rect 14173 8361 14190 8384
rect 14190 8361 14254 8384
rect 14254 8361 14271 8384
rect 14271 8361 14273 8384
rect 14358 8361 14416 8384
rect 14416 8361 14433 8384
rect 14433 8361 14497 8384
rect 14497 8361 14513 8384
rect 14513 8361 14577 8384
rect 14577 8361 14593 8384
rect 14593 8361 14594 8384
rect 14679 8361 14737 8384
rect 14737 8361 14753 8384
rect 14753 8361 14817 8384
rect 14817 8361 14833 8384
rect 14833 8361 14897 8384
rect 14897 8361 14913 8384
rect 14913 8361 14915 8384
rect 15000 8361 15057 8384
rect 15057 8361 15073 8384
rect 15073 8361 15137 8384
rect 15137 8361 15153 8384
rect 15153 8361 15217 8384
rect 15217 8361 15233 8384
rect 15233 8361 15236 8384
rect 15321 8361 15377 8384
rect 15377 8361 15393 8384
rect 15393 8361 15457 8384
rect 15457 8361 15473 8384
rect 15473 8361 15537 8384
rect 15537 8361 15553 8384
rect 15553 8361 15557 8384
rect 215 7757 451 7993
rect 537 7757 773 7993
rect 859 7757 1095 7993
rect 1181 7757 1417 7993
rect 1503 7757 1739 7993
rect 1825 7757 2061 7993
rect 2147 7757 2383 7993
rect 2469 7757 2705 7993
rect 2791 7757 3027 7993
rect 3113 7757 3349 7993
rect 3435 7757 3671 7993
rect 3757 7757 3993 7993
rect 4079 7757 4315 7993
rect 4401 7757 4637 7993
rect 4723 7757 4959 7993
rect 5045 7757 5281 7993
rect 5367 7757 5603 7993
rect 5689 7757 5925 7993
rect 6011 7757 6247 7993
rect 6332 7757 6568 7993
rect 6653 7757 6889 7993
rect 6974 7757 7210 7993
rect 7295 7757 7531 7993
rect 7616 7757 7852 7993
rect 7937 7757 8173 7993
rect 8258 7757 8494 7993
rect 8579 7757 8815 7993
rect 8900 7757 9136 7993
rect 9221 7757 9457 7993
rect 9542 7757 9778 7993
rect 9863 7757 10099 7993
rect 10184 7757 10420 7993
rect 10505 7757 10741 7993
rect 10826 7757 11062 7993
rect 11147 7757 11383 7993
rect 11468 7757 11704 7993
rect 11789 7757 12025 7993
rect 12110 7757 12346 7993
rect 12431 7757 12667 7993
rect 12752 7757 12988 7993
rect 13073 7757 13309 7993
rect 13394 7757 13630 7993
rect 13715 7757 13951 7993
rect 14036 7757 14272 7993
rect 14357 7757 14593 7993
rect 14678 7757 14914 7993
rect 14999 7757 15235 7993
rect 15320 7757 15556 7993
rect 215 7391 451 7627
rect 537 7391 773 7627
rect 859 7391 1095 7627
rect 1181 7391 1417 7627
rect 1503 7391 1739 7627
rect 1825 7391 2061 7627
rect 2147 7391 2383 7627
rect 2469 7391 2705 7627
rect 2791 7391 3027 7627
rect 3113 7391 3349 7627
rect 3435 7391 3671 7627
rect 3757 7391 3993 7627
rect 4079 7391 4315 7627
rect 4401 7391 4637 7627
rect 4723 7391 4959 7627
rect 5045 7391 5281 7627
rect 5367 7391 5603 7627
rect 5689 7391 5925 7627
rect 6011 7391 6247 7627
rect 6332 7391 6568 7627
rect 6653 7391 6889 7627
rect 6974 7391 7210 7627
rect 7295 7391 7531 7627
rect 7616 7391 7852 7627
rect 7937 7391 8173 7627
rect 8258 7391 8494 7627
rect 8579 7391 8815 7627
rect 8900 7391 9136 7627
rect 9221 7391 9457 7627
rect 9542 7391 9778 7627
rect 9863 7391 10099 7627
rect 10184 7391 10420 7627
rect 10505 7391 10741 7627
rect 10826 7391 11062 7627
rect 11147 7391 11383 7627
rect 11468 7391 11704 7627
rect 11789 7391 12025 7627
rect 12110 7391 12346 7627
rect 12431 7391 12667 7627
rect 12752 7391 12988 7627
rect 13073 7391 13309 7627
rect 13394 7391 13630 7627
rect 13715 7391 13951 7627
rect 14036 7391 14272 7627
rect 14357 7391 14593 7627
rect 14678 7391 14914 7627
rect 14999 7391 15235 7627
rect 15320 7391 15556 7627
rect 215 6787 451 7023
rect 537 6787 773 7023
rect 859 6787 1095 7023
rect 1181 6787 1417 7023
rect 1503 6787 1739 7023
rect 1825 6787 2061 7023
rect 2147 6787 2383 7023
rect 2469 6787 2705 7023
rect 2791 6787 3027 7023
rect 3113 6787 3349 7023
rect 3435 6787 3671 7023
rect 3757 6787 3993 7023
rect 4079 6787 4315 7023
rect 4401 6787 4637 7023
rect 4723 6787 4959 7023
rect 5045 6787 5281 7023
rect 5367 6787 5603 7023
rect 5689 6787 5925 7023
rect 6011 6787 6247 7023
rect 6332 6787 6568 7023
rect 6653 6787 6889 7023
rect 6974 6787 7210 7023
rect 7295 6787 7531 7023
rect 7616 6787 7852 7023
rect 7937 6787 8173 7023
rect 8258 6787 8494 7023
rect 8579 6787 8815 7023
rect 8900 6787 9136 7023
rect 9221 6787 9457 7023
rect 9542 6787 9778 7023
rect 9863 6787 10099 7023
rect 10184 6787 10420 7023
rect 10505 6787 10741 7023
rect 10826 6787 11062 7023
rect 11147 6787 11383 7023
rect 11468 6787 11704 7023
rect 11789 6787 12025 7023
rect 12110 6787 12346 7023
rect 12431 6787 12667 7023
rect 12752 6787 12988 7023
rect 13073 6787 13309 7023
rect 13394 6787 13630 7023
rect 13715 6787 13951 7023
rect 14036 6787 14272 7023
rect 14357 6787 14593 7023
rect 14678 6787 14914 7023
rect 14999 6787 15235 7023
rect 15320 6787 15556 7023
rect 215 6421 451 6657
rect 537 6421 773 6657
rect 859 6421 1095 6657
rect 1181 6421 1417 6657
rect 1503 6421 1739 6657
rect 1825 6421 2061 6657
rect 2147 6421 2383 6657
rect 2469 6421 2705 6657
rect 2791 6421 3027 6657
rect 3113 6421 3349 6657
rect 3435 6421 3671 6657
rect 3757 6421 3993 6657
rect 4079 6421 4315 6657
rect 4401 6421 4637 6657
rect 4723 6421 4959 6657
rect 5045 6421 5281 6657
rect 5367 6421 5603 6657
rect 5689 6421 5925 6657
rect 6011 6421 6247 6657
rect 6332 6421 6568 6657
rect 6653 6421 6889 6657
rect 6974 6421 7210 6657
rect 7295 6421 7531 6657
rect 7616 6421 7852 6657
rect 7937 6421 8173 6657
rect 8258 6421 8494 6657
rect 8579 6421 8815 6657
rect 8900 6421 9136 6657
rect 9221 6421 9457 6657
rect 9542 6421 9778 6657
rect 9863 6421 10099 6657
rect 10184 6421 10420 6657
rect 10505 6421 10741 6657
rect 10826 6421 11062 6657
rect 11147 6421 11383 6657
rect 11468 6421 11704 6657
rect 11789 6421 12025 6657
rect 12110 6421 12346 6657
rect 12431 6421 12667 6657
rect 12752 6421 12988 6657
rect 13073 6421 13309 6657
rect 13394 6421 13630 6657
rect 13715 6421 13951 6657
rect 14036 6421 14272 6657
rect 14357 6421 14593 6657
rect 14678 6421 14914 6657
rect 14999 6421 15235 6657
rect 15320 6421 15556 6657
rect 215 5817 451 6053
rect 537 5817 773 6053
rect 859 5817 1095 6053
rect 1181 5817 1417 6053
rect 1503 5817 1739 6053
rect 1825 5817 2061 6053
rect 2147 5817 2383 6053
rect 2469 5817 2705 6053
rect 2791 5817 3027 6053
rect 3113 5817 3349 6053
rect 3435 5817 3671 6053
rect 3757 5817 3993 6053
rect 4079 5817 4315 6053
rect 4401 5817 4637 6053
rect 4723 5817 4959 6053
rect 5045 5817 5281 6053
rect 5367 5817 5603 6053
rect 5689 5817 5925 6053
rect 6011 5817 6247 6053
rect 6332 5817 6568 6053
rect 6653 5817 6889 6053
rect 6974 5817 7210 6053
rect 7295 5817 7531 6053
rect 7616 5817 7852 6053
rect 7937 5817 8173 6053
rect 8258 5817 8494 6053
rect 8579 5817 8815 6053
rect 8900 5817 9136 6053
rect 9221 5817 9457 6053
rect 9542 5817 9778 6053
rect 9863 5817 10099 6053
rect 10184 5817 10420 6053
rect 10505 5817 10741 6053
rect 10826 5817 11062 6053
rect 11147 5817 11383 6053
rect 11468 5817 11704 6053
rect 11789 5817 12025 6053
rect 12110 5817 12346 6053
rect 12431 5817 12667 6053
rect 12752 5817 12988 6053
rect 13073 5817 13309 6053
rect 13394 5817 13630 6053
rect 13715 5817 13951 6053
rect 14036 5817 14272 6053
rect 14357 5817 14593 6053
rect 14678 5817 14914 6053
rect 14999 5817 15235 6053
rect 15320 5817 15556 6053
rect 215 5211 451 5447
rect 537 5211 773 5447
rect 859 5211 1095 5447
rect 1181 5211 1417 5447
rect 1503 5211 1739 5447
rect 1825 5211 2061 5447
rect 2147 5211 2383 5447
rect 2469 5211 2705 5447
rect 2791 5211 3027 5447
rect 3113 5211 3349 5447
rect 3435 5211 3671 5447
rect 3757 5211 3993 5447
rect 4079 5211 4315 5447
rect 4401 5211 4637 5447
rect 4723 5211 4959 5447
rect 5045 5211 5281 5447
rect 5367 5211 5603 5447
rect 5689 5211 5925 5447
rect 6011 5211 6247 5447
rect 6332 5211 6568 5447
rect 6653 5211 6889 5447
rect 6974 5211 7210 5447
rect 7295 5211 7531 5447
rect 7616 5211 7852 5447
rect 7937 5211 8173 5447
rect 8258 5211 8494 5447
rect 8579 5211 8815 5447
rect 8900 5211 9136 5447
rect 9221 5211 9457 5447
rect 9542 5211 9778 5447
rect 9863 5211 10099 5447
rect 10184 5211 10420 5447
rect 10505 5211 10741 5447
rect 10826 5211 11062 5447
rect 11147 5211 11383 5447
rect 11468 5211 11704 5447
rect 11789 5211 12025 5447
rect 12110 5211 12346 5447
rect 12431 5211 12667 5447
rect 12752 5211 12988 5447
rect 13073 5211 13309 5447
rect 13394 5211 13630 5447
rect 13715 5211 13951 5447
rect 14036 5211 14272 5447
rect 14357 5211 14593 5447
rect 14678 5211 14914 5447
rect 14999 5211 15235 5447
rect 15320 5211 15556 5447
rect 215 4607 451 4843
rect 537 4607 773 4843
rect 859 4607 1095 4843
rect 1181 4607 1417 4843
rect 1503 4607 1739 4843
rect 1825 4607 2061 4843
rect 2147 4607 2383 4843
rect 2469 4607 2705 4843
rect 2791 4607 3027 4843
rect 3113 4607 3349 4843
rect 3435 4607 3671 4843
rect 3757 4607 3993 4843
rect 4079 4607 4315 4843
rect 4401 4607 4637 4843
rect 4723 4607 4959 4843
rect 5045 4607 5281 4843
rect 5367 4607 5603 4843
rect 5689 4607 5925 4843
rect 6011 4607 6247 4843
rect 6332 4607 6568 4843
rect 6653 4607 6889 4843
rect 6974 4607 7210 4843
rect 7295 4607 7531 4843
rect 7616 4607 7852 4843
rect 7937 4607 8173 4843
rect 8258 4607 8494 4843
rect 8579 4607 8815 4843
rect 8900 4607 9136 4843
rect 9221 4607 9457 4843
rect 9542 4607 9778 4843
rect 9863 4607 10099 4843
rect 10184 4607 10420 4843
rect 10505 4607 10741 4843
rect 10826 4607 11062 4843
rect 11147 4607 11383 4843
rect 11468 4607 11704 4843
rect 11789 4607 12025 4843
rect 12110 4607 12346 4843
rect 12431 4607 12667 4843
rect 12752 4607 12988 4843
rect 13073 4607 13309 4843
rect 13394 4607 13630 4843
rect 13715 4607 13951 4843
rect 14036 4607 14272 4843
rect 14357 4607 14593 4843
rect 14678 4607 14914 4843
rect 14999 4607 15235 4843
rect 15320 4607 15556 4843
rect 215 4001 451 4237
rect 537 4001 773 4237
rect 859 4001 1095 4237
rect 1181 4001 1417 4237
rect 1503 4001 1739 4237
rect 1825 4001 2061 4237
rect 2147 4001 2383 4237
rect 2469 4001 2705 4237
rect 2791 4001 3027 4237
rect 3113 4001 3349 4237
rect 3435 4001 3671 4237
rect 3757 4001 3993 4237
rect 4079 4001 4315 4237
rect 4401 4001 4637 4237
rect 4723 4001 4959 4237
rect 5045 4001 5281 4237
rect 5367 4001 5603 4237
rect 5689 4001 5925 4237
rect 6011 4001 6247 4237
rect 6332 4001 6568 4237
rect 6653 4001 6889 4237
rect 6974 4001 7210 4237
rect 7295 4001 7531 4237
rect 7616 4001 7852 4237
rect 7937 4001 8173 4237
rect 8258 4001 8494 4237
rect 8579 4001 8815 4237
rect 8900 4001 9136 4237
rect 9221 4001 9457 4237
rect 9542 4001 9778 4237
rect 9863 4001 10099 4237
rect 10184 4001 10420 4237
rect 10505 4001 10741 4237
rect 10826 4001 11062 4237
rect 11147 4001 11383 4237
rect 11468 4001 11704 4237
rect 11789 4001 12025 4237
rect 12110 4001 12346 4237
rect 12431 4001 12667 4237
rect 12752 4001 12988 4237
rect 13073 4001 13309 4237
rect 13394 4001 13630 4237
rect 13715 4001 13951 4237
rect 14036 4001 14272 4237
rect 14357 4001 14593 4237
rect 14678 4001 14914 4237
rect 14999 4001 15235 4237
rect 15320 4001 15556 4237
rect 215 3397 451 3633
rect 537 3397 773 3633
rect 859 3397 1095 3633
rect 1181 3397 1417 3633
rect 1503 3397 1739 3633
rect 1825 3397 2061 3633
rect 2147 3397 2383 3633
rect 2469 3397 2705 3633
rect 2791 3397 3027 3633
rect 3113 3397 3349 3633
rect 3435 3397 3671 3633
rect 3757 3397 3993 3633
rect 4079 3397 4315 3633
rect 4401 3397 4637 3633
rect 4723 3397 4959 3633
rect 5045 3397 5281 3633
rect 5367 3397 5603 3633
rect 5689 3397 5925 3633
rect 6011 3397 6247 3633
rect 6332 3397 6568 3633
rect 6653 3397 6889 3633
rect 6974 3397 7210 3633
rect 7295 3397 7531 3633
rect 7616 3397 7852 3633
rect 7937 3397 8173 3633
rect 8258 3397 8494 3633
rect 8579 3397 8815 3633
rect 8900 3397 9136 3633
rect 9221 3397 9457 3633
rect 9542 3397 9778 3633
rect 9863 3397 10099 3633
rect 10184 3397 10420 3633
rect 10505 3397 10741 3633
rect 10826 3397 11062 3633
rect 11147 3397 11383 3633
rect 11468 3397 11704 3633
rect 11789 3397 12025 3633
rect 12110 3397 12346 3633
rect 12431 3397 12667 3633
rect 12752 3397 12988 3633
rect 13073 3397 13309 3633
rect 13394 3397 13630 3633
rect 13715 3397 13951 3633
rect 14036 3397 14272 3633
rect 14357 3397 14593 3633
rect 14678 3397 14914 3633
rect 14999 3397 15235 3633
rect 15320 3397 15556 3633
rect 215 3031 451 3267
rect 537 3031 773 3267
rect 859 3031 1095 3267
rect 1181 3031 1417 3267
rect 1503 3031 1739 3267
rect 1825 3031 2061 3267
rect 2147 3031 2383 3267
rect 2469 3031 2705 3267
rect 2791 3031 3027 3267
rect 3113 3031 3349 3267
rect 3435 3031 3671 3267
rect 3757 3031 3993 3267
rect 4079 3031 4315 3267
rect 4401 3031 4637 3267
rect 4723 3031 4959 3267
rect 5045 3031 5281 3267
rect 5367 3031 5603 3267
rect 5689 3031 5925 3267
rect 6011 3031 6247 3267
rect 6332 3031 6568 3267
rect 6653 3031 6889 3267
rect 6974 3031 7210 3267
rect 7295 3031 7531 3267
rect 7616 3031 7852 3267
rect 7937 3031 8173 3267
rect 8258 3031 8494 3267
rect 8579 3031 8815 3267
rect 8900 3031 9136 3267
rect 9221 3031 9457 3267
rect 9542 3031 9778 3267
rect 9863 3031 10099 3267
rect 10184 3031 10420 3267
rect 10505 3031 10741 3267
rect 10826 3031 11062 3267
rect 11147 3031 11383 3267
rect 11468 3031 11704 3267
rect 11789 3031 12025 3267
rect 12110 3031 12346 3267
rect 12431 3031 12667 3267
rect 12752 3031 12988 3267
rect 13073 3031 13309 3267
rect 13394 3031 13630 3267
rect 13715 3031 13951 3267
rect 14036 3031 14272 3267
rect 14357 3031 14593 3267
rect 14678 3031 14914 3267
rect 14999 3031 15235 3267
rect 15320 3031 15556 3267
rect 215 2427 451 2663
rect 537 2637 547 2663
rect 547 2637 611 2663
rect 611 2637 659 2663
rect 659 2637 723 2663
rect 723 2637 771 2663
rect 771 2637 773 2663
rect 859 2637 883 2663
rect 883 2637 947 2663
rect 947 2637 1095 2663
rect 537 2579 773 2637
rect 859 2579 1095 2637
rect 537 2515 547 2579
rect 547 2515 611 2579
rect 611 2515 659 2579
rect 659 2515 723 2579
rect 723 2515 771 2579
rect 771 2515 773 2579
rect 859 2515 883 2579
rect 883 2515 947 2579
rect 947 2515 1095 2579
rect 537 2457 773 2515
rect 859 2457 1095 2515
rect 537 2427 547 2457
rect 547 2427 611 2457
rect 611 2427 659 2457
rect 659 2427 723 2457
rect 723 2427 771 2457
rect 771 2427 773 2457
rect 859 2427 883 2457
rect 883 2427 947 2457
rect 947 2427 1095 2457
rect 1181 2427 1417 2663
rect 1503 2427 1739 2663
rect 1825 2427 2061 2663
rect 2147 2427 2383 2663
rect 2469 2427 2705 2663
rect 2791 2427 3027 2663
rect 3113 2427 3349 2663
rect 3435 2427 3671 2663
rect 3757 2427 3993 2663
rect 4079 2427 4315 2663
rect 4401 2427 4637 2663
rect 4723 2427 4959 2663
rect 5045 2427 5281 2663
rect 5367 2427 5603 2663
rect 5689 2427 5925 2663
rect 6011 2427 6247 2663
rect 6332 2427 6568 2663
rect 6653 2427 6889 2663
rect 6974 2427 7210 2663
rect 7295 2427 7531 2663
rect 7616 2427 7852 2663
rect 7937 2427 8173 2663
rect 8258 2427 8494 2663
rect 8579 2427 8815 2663
rect 8900 2427 9136 2663
rect 9221 2427 9457 2663
rect 9542 2427 9778 2663
rect 9863 2427 10099 2663
rect 10184 2427 10420 2663
rect 10505 2427 10741 2663
rect 10826 2427 11062 2663
rect 11147 2427 11383 2663
rect 11468 2637 11674 2663
rect 11674 2637 11704 2663
rect 11468 2579 11704 2637
rect 11468 2515 11674 2579
rect 11674 2515 11704 2579
rect 11468 2457 11704 2515
rect 11468 2427 11674 2457
rect 11674 2427 11704 2457
rect 11789 2427 12025 2663
rect 12110 2427 12346 2663
rect 12431 2427 12667 2663
rect 12752 2427 12988 2663
rect 13073 2427 13309 2663
rect 13394 2427 13630 2663
rect 13715 2427 13951 2663
rect 14036 2427 14272 2663
rect 14357 2427 14593 2663
rect 14678 2427 14914 2663
rect 14999 2427 15235 2663
rect 15320 2427 15556 2663
rect 215 1821 451 2057
rect 537 2027 547 2057
rect 547 2027 611 2057
rect 611 2027 659 2057
rect 659 2027 723 2057
rect 723 2027 771 2057
rect 771 2027 773 2057
rect 859 2027 883 2057
rect 883 2027 947 2057
rect 947 2027 1095 2057
rect 537 1969 773 2027
rect 859 1969 1095 2027
rect 537 1905 547 1969
rect 547 1905 611 1969
rect 611 1905 659 1969
rect 659 1905 723 1969
rect 723 1905 771 1969
rect 771 1905 773 1969
rect 859 1905 883 1969
rect 883 1905 947 1969
rect 947 1905 1095 1969
rect 537 1847 773 1905
rect 859 1847 1095 1905
rect 537 1821 547 1847
rect 547 1821 611 1847
rect 611 1821 659 1847
rect 659 1821 723 1847
rect 723 1821 771 1847
rect 771 1821 773 1847
rect 859 1821 883 1847
rect 883 1821 947 1847
rect 947 1821 1095 1847
rect 1181 1821 1417 2057
rect 1503 1821 1739 2057
rect 1825 1821 2061 2057
rect 2147 1821 2383 2057
rect 2469 1821 2705 2057
rect 2791 1821 3027 2057
rect 3113 1821 3349 2057
rect 3435 1821 3671 2057
rect 3757 1821 3993 2057
rect 4079 1821 4315 2057
rect 4401 1821 4637 2057
rect 4723 1821 4959 2057
rect 5045 1821 5281 2057
rect 5367 1821 5603 2057
rect 5689 1821 5925 2057
rect 6011 1821 6247 2057
rect 6332 1821 6568 2057
rect 6653 1821 6889 2057
rect 6974 1821 7210 2057
rect 7295 1821 7531 2057
rect 7616 1821 7852 2057
rect 7937 1821 8173 2057
rect 8258 1821 8494 2057
rect 8579 1821 8815 2057
rect 8900 1821 9136 2057
rect 9221 1821 9457 2057
rect 9542 1821 9778 2057
rect 9863 1821 10099 2057
rect 10184 1821 10420 2057
rect 10505 1821 10741 2057
rect 10826 1821 11062 2057
rect 11147 1821 11383 2057
rect 11468 2027 11674 2057
rect 11674 2027 11704 2057
rect 11468 1969 11704 2027
rect 11468 1905 11674 1969
rect 11674 1905 11704 1969
rect 11468 1847 11704 1905
rect 11468 1821 11674 1847
rect 11674 1821 11704 1847
rect 11789 1821 12025 2057
rect 12110 1821 12346 2057
rect 12431 1821 12667 2057
rect 12752 1821 12988 2057
rect 13073 1821 13309 2057
rect 13394 1821 13630 2057
rect 13715 1821 13951 2057
rect 14036 1821 14272 2057
rect 14357 1821 14593 2057
rect 14678 1821 14914 2057
rect 14999 1821 15235 2057
rect 15320 1821 15556 2057
rect 215 1216 451 1452
rect 537 1216 773 1452
rect 859 1216 1095 1452
rect 1181 1216 1417 1452
rect 1503 1216 1739 1452
rect 1825 1216 2061 1452
rect 2147 1216 2383 1452
rect 2469 1216 2705 1452
rect 2791 1216 3027 1452
rect 3113 1216 3349 1452
rect 3435 1216 3671 1452
rect 3757 1216 3993 1452
rect 4079 1216 4315 1452
rect 4401 1216 4637 1452
rect 4723 1216 4959 1452
rect 5045 1216 5281 1452
rect 5367 1216 5603 1452
rect 5689 1216 5925 1452
rect 6011 1216 6247 1452
rect 6332 1216 6568 1452
rect 6653 1216 6889 1452
rect 6974 1216 7210 1452
rect 7295 1216 7531 1452
rect 7616 1216 7852 1452
rect 7937 1216 8173 1452
rect 8258 1216 8494 1452
rect 8579 1216 8815 1452
rect 8900 1216 9136 1452
rect 9221 1216 9457 1452
rect 9542 1216 9778 1452
rect 9863 1216 10099 1452
rect 10184 1216 10420 1452
rect 10505 1216 10741 1452
rect 10826 1216 11062 1452
rect 11147 1216 11383 1452
rect 11468 1216 11704 1452
rect 11789 1216 12025 1452
rect 12110 1216 12346 1452
rect 12431 1216 12667 1452
rect 12752 1216 12988 1452
rect 13073 1216 13309 1452
rect 13394 1216 13630 1452
rect 13715 1216 13951 1452
rect 14036 1216 14272 1452
rect 14357 1216 14593 1452
rect 14678 1216 14914 1452
rect 14999 1216 15235 1452
rect 15320 1216 15556 1452
rect 215 834 451 1070
rect 537 834 773 1070
rect 859 834 1095 1070
rect 1181 834 1417 1070
rect 1503 834 1739 1070
rect 1825 834 2061 1070
rect 2147 834 2383 1070
rect 2469 834 2705 1070
rect 2791 834 3027 1070
rect 3113 834 3349 1070
rect 3435 834 3671 1070
rect 3757 834 3993 1070
rect 4079 834 4315 1070
rect 4401 834 4637 1070
rect 4723 834 4959 1070
rect 5045 834 5281 1070
rect 5367 834 5603 1070
rect 5689 834 5925 1070
rect 6011 834 6247 1070
rect 6332 834 6568 1070
rect 6653 834 6889 1070
rect 6974 834 7210 1070
rect 7295 834 7531 1070
rect 7616 834 7852 1070
rect 7937 834 8173 1070
rect 8258 834 8494 1070
rect 8579 834 8815 1070
rect 8900 834 9136 1070
rect 9221 834 9457 1070
rect 9542 834 9778 1070
rect 9863 834 10099 1070
rect 10184 834 10420 1070
rect 10505 834 10741 1070
rect 10826 834 11062 1070
rect 11147 834 11383 1070
rect 11468 834 11704 1070
rect 11789 834 12025 1070
rect 12110 834 12346 1070
rect 12431 834 12667 1070
rect 12752 834 12988 1070
rect 13073 834 13309 1070
rect 13394 834 13630 1070
rect 13715 834 13951 1070
rect 14036 834 14272 1070
rect 14357 834 14593 1070
rect 14678 834 14914 1070
rect 14999 834 15235 1070
rect 15320 834 15556 1070
rect 215 452 451 688
rect 537 452 773 688
rect 859 452 1095 688
rect 1181 452 1417 688
rect 1503 452 1739 688
rect 1825 452 2061 688
rect 2147 452 2383 688
rect 2469 452 2705 688
rect 2791 452 3027 688
rect 3113 452 3349 688
rect 3435 452 3671 688
rect 3757 452 3993 688
rect 4079 452 4315 688
rect 4401 452 4637 688
rect 4723 452 4959 688
rect 5045 452 5281 688
rect 5367 452 5603 688
rect 5689 452 5925 688
rect 6011 452 6247 688
rect 6332 452 6568 688
rect 6653 452 6889 688
rect 6974 452 7210 688
rect 7295 452 7531 688
rect 7616 452 7852 688
rect 7937 452 8173 688
rect 8258 452 8494 688
rect 8579 452 8815 688
rect 8900 452 9136 688
rect 9221 452 9457 688
rect 9542 452 9778 688
rect 9863 452 10099 688
rect 10184 452 10420 688
rect 10505 452 10741 688
rect 10826 452 11062 688
rect 11147 452 11383 688
rect 11468 452 11704 688
rect 11789 452 12025 688
rect 12110 452 12346 688
rect 12431 452 12667 688
rect 12752 452 12988 688
rect 13073 452 13309 688
rect 13394 452 13630 688
rect 13715 452 13951 688
rect 14036 452 14272 688
rect 14357 452 14593 688
rect 14678 452 14914 688
rect 14999 452 15235 688
rect 15320 452 15556 688
<< metal5 >>
rect 0 39964 16000 40000
rect 0 39728 215 39964
rect 451 39728 537 39964
rect 773 39728 859 39964
rect 1095 39728 1181 39964
rect 1417 39728 1503 39964
rect 1739 39728 1825 39964
rect 2061 39728 2147 39964
rect 2383 39728 2469 39964
rect 2705 39728 2791 39964
rect 3027 39728 3113 39964
rect 3349 39728 3435 39964
rect 3671 39728 3757 39964
rect 3993 39728 4079 39964
rect 4315 39728 4401 39964
rect 4637 39728 4723 39964
rect 4959 39728 5045 39964
rect 5281 39728 5367 39964
rect 5603 39728 5689 39964
rect 5925 39728 6011 39964
rect 6247 39728 6332 39964
rect 6568 39728 6653 39964
rect 6889 39728 6974 39964
rect 7210 39728 7295 39964
rect 7531 39728 7616 39964
rect 7852 39728 7937 39964
rect 8173 39728 8258 39964
rect 8494 39728 8579 39964
rect 8815 39728 8900 39964
rect 9136 39728 9221 39964
rect 9457 39728 9542 39964
rect 9778 39728 9863 39964
rect 10099 39728 10184 39964
rect 10420 39728 10505 39964
rect 10741 39728 10826 39964
rect 11062 39728 11147 39964
rect 11383 39728 11468 39964
rect 11704 39728 11789 39964
rect 12025 39728 12110 39964
rect 12346 39728 12431 39964
rect 12667 39728 12752 39964
rect 12988 39728 13073 39964
rect 13309 39728 13394 39964
rect 13630 39728 13715 39964
rect 13951 39728 14036 39964
rect 14272 39728 14357 39964
rect 14593 39728 14678 39964
rect 14914 39728 14999 39964
rect 15235 39728 15320 39964
rect 15556 39728 16000 39964
rect 0 39640 16000 39728
rect 0 39404 215 39640
rect 451 39404 537 39640
rect 773 39404 859 39640
rect 1095 39404 1181 39640
rect 1417 39404 1503 39640
rect 1739 39404 1825 39640
rect 2061 39404 2147 39640
rect 2383 39404 2469 39640
rect 2705 39404 2791 39640
rect 3027 39404 3113 39640
rect 3349 39404 3435 39640
rect 3671 39404 3757 39640
rect 3993 39404 4079 39640
rect 4315 39404 4401 39640
rect 4637 39404 4723 39640
rect 4959 39404 5045 39640
rect 5281 39404 5367 39640
rect 5603 39404 5689 39640
rect 5925 39404 6011 39640
rect 6247 39404 6332 39640
rect 6568 39404 6653 39640
rect 6889 39404 6974 39640
rect 7210 39404 7295 39640
rect 7531 39404 7616 39640
rect 7852 39404 7937 39640
rect 8173 39404 8258 39640
rect 8494 39404 8579 39640
rect 8815 39404 8900 39640
rect 9136 39404 9221 39640
rect 9457 39404 9542 39640
rect 9778 39404 9863 39640
rect 10099 39404 10184 39640
rect 10420 39404 10505 39640
rect 10741 39404 10826 39640
rect 11062 39404 11147 39640
rect 11383 39404 11468 39640
rect 11704 39404 11789 39640
rect 12025 39404 12110 39640
rect 12346 39404 12431 39640
rect 12667 39404 12752 39640
rect 12988 39404 13073 39640
rect 13309 39404 13394 39640
rect 13630 39404 13715 39640
rect 13951 39404 14036 39640
rect 14272 39404 14357 39640
rect 14593 39404 14678 39640
rect 14914 39404 14999 39640
rect 15235 39404 15320 39640
rect 15556 39404 16000 39640
rect 0 39316 16000 39404
rect 0 39080 215 39316
rect 451 39080 537 39316
rect 773 39080 859 39316
rect 1095 39080 1181 39316
rect 1417 39080 1503 39316
rect 1739 39080 1825 39316
rect 2061 39080 2147 39316
rect 2383 39080 2469 39316
rect 2705 39080 2791 39316
rect 3027 39080 3113 39316
rect 3349 39080 3435 39316
rect 3671 39080 3757 39316
rect 3993 39080 4079 39316
rect 4315 39080 4401 39316
rect 4637 39080 4723 39316
rect 4959 39080 5045 39316
rect 5281 39080 5367 39316
rect 5603 39080 5689 39316
rect 5925 39080 6011 39316
rect 6247 39080 6332 39316
rect 6568 39080 6653 39316
rect 6889 39080 6974 39316
rect 7210 39080 7295 39316
rect 7531 39080 7616 39316
rect 7852 39080 7937 39316
rect 8173 39080 8258 39316
rect 8494 39080 8579 39316
rect 8815 39080 8900 39316
rect 9136 39080 9221 39316
rect 9457 39080 9542 39316
rect 9778 39080 9863 39316
rect 10099 39080 10184 39316
rect 10420 39080 10505 39316
rect 10741 39080 10826 39316
rect 11062 39080 11147 39316
rect 11383 39080 11468 39316
rect 11704 39080 11789 39316
rect 12025 39080 12110 39316
rect 12346 39080 12431 39316
rect 12667 39080 12752 39316
rect 12988 39080 13073 39316
rect 13309 39080 13394 39316
rect 13630 39080 13715 39316
rect 13951 39080 14036 39316
rect 14272 39080 14357 39316
rect 14593 39080 14678 39316
rect 14914 39080 14999 39316
rect 15235 39080 15320 39316
rect 15556 39080 16000 39316
rect 0 38992 16000 39080
rect 0 38756 215 38992
rect 451 38756 537 38992
rect 773 38756 859 38992
rect 1095 38756 1181 38992
rect 1417 38756 1503 38992
rect 1739 38756 1825 38992
rect 2061 38756 2147 38992
rect 2383 38756 2469 38992
rect 2705 38756 2791 38992
rect 3027 38756 3113 38992
rect 3349 38756 3435 38992
rect 3671 38756 3757 38992
rect 3993 38756 4079 38992
rect 4315 38756 4401 38992
rect 4637 38756 4723 38992
rect 4959 38756 5045 38992
rect 5281 38756 5367 38992
rect 5603 38756 5689 38992
rect 5925 38756 6011 38992
rect 6247 38756 6332 38992
rect 6568 38756 6653 38992
rect 6889 38756 6974 38992
rect 7210 38756 7295 38992
rect 7531 38756 7616 38992
rect 7852 38756 7937 38992
rect 8173 38756 8258 38992
rect 8494 38756 8579 38992
rect 8815 38756 8900 38992
rect 9136 38756 9221 38992
rect 9457 38756 9542 38992
rect 9778 38756 9863 38992
rect 10099 38756 10184 38992
rect 10420 38756 10505 38992
rect 10741 38756 10826 38992
rect 11062 38756 11147 38992
rect 11383 38756 11468 38992
rect 11704 38756 11789 38992
rect 12025 38756 12110 38992
rect 12346 38756 12431 38992
rect 12667 38756 12752 38992
rect 12988 38756 13073 38992
rect 13309 38756 13394 38992
rect 13630 38756 13715 38992
rect 13951 38756 14036 38992
rect 14272 38756 14357 38992
rect 14593 38756 14678 38992
rect 14914 38756 14999 38992
rect 15235 38756 15320 38992
rect 15556 38756 16000 38992
rect 0 38668 16000 38756
rect 0 38432 215 38668
rect 451 38432 537 38668
rect 773 38432 859 38668
rect 1095 38432 1181 38668
rect 1417 38432 1503 38668
rect 1739 38432 1825 38668
rect 2061 38432 2147 38668
rect 2383 38432 2469 38668
rect 2705 38432 2791 38668
rect 3027 38432 3113 38668
rect 3349 38432 3435 38668
rect 3671 38432 3757 38668
rect 3993 38432 4079 38668
rect 4315 38432 4401 38668
rect 4637 38432 4723 38668
rect 4959 38432 5045 38668
rect 5281 38432 5367 38668
rect 5603 38432 5689 38668
rect 5925 38432 6011 38668
rect 6247 38432 6332 38668
rect 6568 38432 6653 38668
rect 6889 38432 6974 38668
rect 7210 38432 7295 38668
rect 7531 38432 7616 38668
rect 7852 38432 7937 38668
rect 8173 38432 8258 38668
rect 8494 38432 8579 38668
rect 8815 38432 8900 38668
rect 9136 38432 9221 38668
rect 9457 38432 9542 38668
rect 9778 38432 9863 38668
rect 10099 38432 10184 38668
rect 10420 38432 10505 38668
rect 10741 38432 10826 38668
rect 11062 38432 11147 38668
rect 11383 38432 11468 38668
rect 11704 38432 11789 38668
rect 12025 38432 12110 38668
rect 12346 38432 12431 38668
rect 12667 38432 12752 38668
rect 12988 38432 13073 38668
rect 13309 38432 13394 38668
rect 13630 38432 13715 38668
rect 13951 38432 14036 38668
rect 14272 38432 14357 38668
rect 14593 38432 14678 38668
rect 14914 38432 14999 38668
rect 15235 38432 15320 38668
rect 15556 38432 16000 38668
rect 0 38344 16000 38432
rect 0 38108 215 38344
rect 451 38108 537 38344
rect 773 38108 859 38344
rect 1095 38108 1181 38344
rect 1417 38108 1503 38344
rect 1739 38108 1825 38344
rect 2061 38108 2147 38344
rect 2383 38108 2469 38344
rect 2705 38108 2791 38344
rect 3027 38108 3113 38344
rect 3349 38108 3435 38344
rect 3671 38108 3757 38344
rect 3993 38108 4079 38344
rect 4315 38108 4401 38344
rect 4637 38108 4723 38344
rect 4959 38108 5045 38344
rect 5281 38108 5367 38344
rect 5603 38108 5689 38344
rect 5925 38108 6011 38344
rect 6247 38108 6332 38344
rect 6568 38108 6653 38344
rect 6889 38108 6974 38344
rect 7210 38108 7295 38344
rect 7531 38108 7616 38344
rect 7852 38108 7937 38344
rect 8173 38108 8258 38344
rect 8494 38108 8579 38344
rect 8815 38108 8900 38344
rect 9136 38108 9221 38344
rect 9457 38108 9542 38344
rect 9778 38108 9863 38344
rect 10099 38108 10184 38344
rect 10420 38108 10505 38344
rect 10741 38108 10826 38344
rect 11062 38108 11147 38344
rect 11383 38108 11468 38344
rect 11704 38108 11789 38344
rect 12025 38108 12110 38344
rect 12346 38108 12431 38344
rect 12667 38108 12752 38344
rect 12988 38108 13073 38344
rect 13309 38108 13394 38344
rect 13630 38108 13715 38344
rect 13951 38108 14036 38344
rect 14272 38108 14357 38344
rect 14593 38108 14678 38344
rect 14914 38108 14999 38344
rect 15235 38108 15320 38344
rect 15556 38108 16000 38344
rect 0 38020 16000 38108
rect 0 37784 215 38020
rect 451 37784 537 38020
rect 773 37784 859 38020
rect 1095 37784 1181 38020
rect 1417 37784 1503 38020
rect 1739 37784 1825 38020
rect 2061 37784 2147 38020
rect 2383 37784 2469 38020
rect 2705 37784 2791 38020
rect 3027 37784 3113 38020
rect 3349 37784 3435 38020
rect 3671 37784 3757 38020
rect 3993 37784 4079 38020
rect 4315 37784 4401 38020
rect 4637 37784 4723 38020
rect 4959 37784 5045 38020
rect 5281 37784 5367 38020
rect 5603 37784 5689 38020
rect 5925 37784 6011 38020
rect 6247 37784 6332 38020
rect 6568 37784 6653 38020
rect 6889 37784 6974 38020
rect 7210 37784 7295 38020
rect 7531 37784 7616 38020
rect 7852 37784 7937 38020
rect 8173 37784 8258 38020
rect 8494 37784 8579 38020
rect 8815 37784 8900 38020
rect 9136 37784 9221 38020
rect 9457 37784 9542 38020
rect 9778 37784 9863 38020
rect 10099 37784 10184 38020
rect 10420 37784 10505 38020
rect 10741 37784 10826 38020
rect 11062 37784 11147 38020
rect 11383 37784 11468 38020
rect 11704 37784 11789 38020
rect 12025 37784 12110 38020
rect 12346 37784 12431 38020
rect 12667 37784 12752 38020
rect 12988 37784 13073 38020
rect 13309 37784 13394 38020
rect 13630 37784 13715 38020
rect 13951 37784 14036 38020
rect 14272 37784 14357 38020
rect 14593 37784 14678 38020
rect 14914 37784 14999 38020
rect 15235 37784 15320 38020
rect 15556 37784 16000 38020
rect 0 37696 16000 37784
rect 0 37460 215 37696
rect 451 37460 537 37696
rect 773 37460 859 37696
rect 1095 37460 1181 37696
rect 1417 37460 1503 37696
rect 1739 37460 1825 37696
rect 2061 37460 2147 37696
rect 2383 37460 2469 37696
rect 2705 37460 2791 37696
rect 3027 37460 3113 37696
rect 3349 37460 3435 37696
rect 3671 37460 3757 37696
rect 3993 37460 4079 37696
rect 4315 37460 4401 37696
rect 4637 37460 4723 37696
rect 4959 37460 5045 37696
rect 5281 37460 5367 37696
rect 5603 37460 5689 37696
rect 5925 37460 6011 37696
rect 6247 37460 6332 37696
rect 6568 37460 6653 37696
rect 6889 37460 6974 37696
rect 7210 37460 7295 37696
rect 7531 37460 7616 37696
rect 7852 37460 7937 37696
rect 8173 37460 8258 37696
rect 8494 37460 8579 37696
rect 8815 37460 8900 37696
rect 9136 37460 9221 37696
rect 9457 37460 9542 37696
rect 9778 37460 9863 37696
rect 10099 37460 10184 37696
rect 10420 37460 10505 37696
rect 10741 37460 10826 37696
rect 11062 37460 11147 37696
rect 11383 37460 11468 37696
rect 11704 37460 11789 37696
rect 12025 37460 12110 37696
rect 12346 37460 12431 37696
rect 12667 37460 12752 37696
rect 12988 37460 13073 37696
rect 13309 37460 13394 37696
rect 13630 37460 13715 37696
rect 13951 37460 14036 37696
rect 14272 37460 14357 37696
rect 14593 37460 14678 37696
rect 14914 37460 14999 37696
rect 15235 37460 15320 37696
rect 15556 37460 16000 37696
rect 0 37372 16000 37460
rect 0 37136 215 37372
rect 451 37136 537 37372
rect 773 37136 859 37372
rect 1095 37136 1181 37372
rect 1417 37136 1503 37372
rect 1739 37136 1825 37372
rect 2061 37136 2147 37372
rect 2383 37136 2469 37372
rect 2705 37136 2791 37372
rect 3027 37136 3113 37372
rect 3349 37136 3435 37372
rect 3671 37136 3757 37372
rect 3993 37136 4079 37372
rect 4315 37136 4401 37372
rect 4637 37136 4723 37372
rect 4959 37136 5045 37372
rect 5281 37136 5367 37372
rect 5603 37136 5689 37372
rect 5925 37136 6011 37372
rect 6247 37136 6332 37372
rect 6568 37136 6653 37372
rect 6889 37136 6974 37372
rect 7210 37136 7295 37372
rect 7531 37136 7616 37372
rect 7852 37136 7937 37372
rect 8173 37136 8258 37372
rect 8494 37136 8579 37372
rect 8815 37136 8900 37372
rect 9136 37136 9221 37372
rect 9457 37136 9542 37372
rect 9778 37136 9863 37372
rect 10099 37136 10184 37372
rect 10420 37136 10505 37372
rect 10741 37136 10826 37372
rect 11062 37136 11147 37372
rect 11383 37136 11468 37372
rect 11704 37136 11789 37372
rect 12025 37136 12110 37372
rect 12346 37136 12431 37372
rect 12667 37136 12752 37372
rect 12988 37136 13073 37372
rect 13309 37136 13394 37372
rect 13630 37136 13715 37372
rect 13951 37136 14036 37372
rect 14272 37136 14357 37372
rect 14593 37136 14678 37372
rect 14914 37136 14999 37372
rect 15235 37136 15320 37372
rect 15556 37136 16000 37372
rect 0 37048 16000 37136
rect 0 36812 215 37048
rect 451 36812 537 37048
rect 773 36812 859 37048
rect 1095 36812 1181 37048
rect 1417 36812 1503 37048
rect 1739 36812 1825 37048
rect 2061 36812 2147 37048
rect 2383 36812 2469 37048
rect 2705 36812 2791 37048
rect 3027 36812 3113 37048
rect 3349 36812 3435 37048
rect 3671 36812 3757 37048
rect 3993 36812 4079 37048
rect 4315 36812 4401 37048
rect 4637 36812 4723 37048
rect 4959 36812 5045 37048
rect 5281 36812 5367 37048
rect 5603 36812 5689 37048
rect 5925 36812 6011 37048
rect 6247 36812 6332 37048
rect 6568 36812 6653 37048
rect 6889 36812 6974 37048
rect 7210 36812 7295 37048
rect 7531 36812 7616 37048
rect 7852 36812 7937 37048
rect 8173 36812 8258 37048
rect 8494 36812 8579 37048
rect 8815 36812 8900 37048
rect 9136 36812 9221 37048
rect 9457 36812 9542 37048
rect 9778 36812 9863 37048
rect 10099 36812 10184 37048
rect 10420 36812 10505 37048
rect 10741 36812 10826 37048
rect 11062 36812 11147 37048
rect 11383 36812 11468 37048
rect 11704 36812 11789 37048
rect 12025 36812 12110 37048
rect 12346 36812 12431 37048
rect 12667 36812 12752 37048
rect 12988 36812 13073 37048
rect 13309 36812 13394 37048
rect 13630 36812 13715 37048
rect 13951 36812 14036 37048
rect 14272 36812 14357 37048
rect 14593 36812 14678 37048
rect 14914 36812 14999 37048
rect 15235 36812 15320 37048
rect 15556 36812 16000 37048
rect 0 36724 16000 36812
rect 0 36488 215 36724
rect 451 36488 537 36724
rect 773 36488 859 36724
rect 1095 36488 1181 36724
rect 1417 36488 1503 36724
rect 1739 36488 1825 36724
rect 2061 36488 2147 36724
rect 2383 36488 2469 36724
rect 2705 36488 2791 36724
rect 3027 36488 3113 36724
rect 3349 36488 3435 36724
rect 3671 36488 3757 36724
rect 3993 36488 4079 36724
rect 4315 36488 4401 36724
rect 4637 36488 4723 36724
rect 4959 36488 5045 36724
rect 5281 36488 5367 36724
rect 5603 36488 5689 36724
rect 5925 36488 6011 36724
rect 6247 36488 6332 36724
rect 6568 36488 6653 36724
rect 6889 36488 6974 36724
rect 7210 36488 7295 36724
rect 7531 36488 7616 36724
rect 7852 36488 7937 36724
rect 8173 36488 8258 36724
rect 8494 36488 8579 36724
rect 8815 36488 8900 36724
rect 9136 36488 9221 36724
rect 9457 36488 9542 36724
rect 9778 36488 9863 36724
rect 10099 36488 10184 36724
rect 10420 36488 10505 36724
rect 10741 36488 10826 36724
rect 11062 36488 11147 36724
rect 11383 36488 11468 36724
rect 11704 36488 11789 36724
rect 12025 36488 12110 36724
rect 12346 36488 12431 36724
rect 12667 36488 12752 36724
rect 12988 36488 13073 36724
rect 13309 36488 13394 36724
rect 13630 36488 13715 36724
rect 13951 36488 14036 36724
rect 14272 36488 14357 36724
rect 14593 36488 14678 36724
rect 14914 36488 14999 36724
rect 15235 36488 15320 36724
rect 15556 36488 16000 36724
rect 0 36400 16000 36488
rect 0 36164 215 36400
rect 451 36164 537 36400
rect 773 36164 859 36400
rect 1095 36164 1181 36400
rect 1417 36164 1503 36400
rect 1739 36164 1825 36400
rect 2061 36164 2147 36400
rect 2383 36164 2469 36400
rect 2705 36164 2791 36400
rect 3027 36164 3113 36400
rect 3349 36164 3435 36400
rect 3671 36164 3757 36400
rect 3993 36164 4079 36400
rect 4315 36164 4401 36400
rect 4637 36164 4723 36400
rect 4959 36164 5045 36400
rect 5281 36164 5367 36400
rect 5603 36164 5689 36400
rect 5925 36164 6011 36400
rect 6247 36164 6332 36400
rect 6568 36164 6653 36400
rect 6889 36164 6974 36400
rect 7210 36164 7295 36400
rect 7531 36164 7616 36400
rect 7852 36164 7937 36400
rect 8173 36164 8258 36400
rect 8494 36164 8579 36400
rect 8815 36164 8900 36400
rect 9136 36164 9221 36400
rect 9457 36164 9542 36400
rect 9778 36164 9863 36400
rect 10099 36164 10184 36400
rect 10420 36164 10505 36400
rect 10741 36164 10826 36400
rect 11062 36164 11147 36400
rect 11383 36164 11468 36400
rect 11704 36164 11789 36400
rect 12025 36164 12110 36400
rect 12346 36164 12431 36400
rect 12667 36164 12752 36400
rect 12988 36164 13073 36400
rect 13309 36164 13394 36400
rect 13630 36164 13715 36400
rect 13951 36164 14036 36400
rect 14272 36164 14357 36400
rect 14593 36164 14678 36400
rect 14914 36164 14999 36400
rect 15235 36164 15320 36400
rect 15556 36164 16000 36400
rect 0 36076 16000 36164
rect 0 35840 215 36076
rect 451 35840 537 36076
rect 773 35840 859 36076
rect 1095 35840 1181 36076
rect 1417 35840 1503 36076
rect 1739 35840 1825 36076
rect 2061 35840 2147 36076
rect 2383 35840 2469 36076
rect 2705 35840 2791 36076
rect 3027 35840 3113 36076
rect 3349 35840 3435 36076
rect 3671 35840 3757 36076
rect 3993 35840 4079 36076
rect 4315 35840 4401 36076
rect 4637 35840 4723 36076
rect 4959 35840 5045 36076
rect 5281 35840 5367 36076
rect 5603 35840 5689 36076
rect 5925 35840 6011 36076
rect 6247 35840 6332 36076
rect 6568 35840 6653 36076
rect 6889 35840 6974 36076
rect 7210 35840 7295 36076
rect 7531 35840 7616 36076
rect 7852 35840 7937 36076
rect 8173 35840 8258 36076
rect 8494 35840 8579 36076
rect 8815 35840 8900 36076
rect 9136 35840 9221 36076
rect 9457 35840 9542 36076
rect 9778 35840 9863 36076
rect 10099 35840 10184 36076
rect 10420 35840 10505 36076
rect 10741 35840 10826 36076
rect 11062 35840 11147 36076
rect 11383 35840 11468 36076
rect 11704 35840 11789 36076
rect 12025 35840 12110 36076
rect 12346 35840 12431 36076
rect 12667 35840 12752 36076
rect 12988 35840 13073 36076
rect 13309 35840 13394 36076
rect 13630 35840 13715 36076
rect 13951 35840 14036 36076
rect 14272 35840 14357 36076
rect 14593 35840 14678 36076
rect 14914 35840 14999 36076
rect 15235 35840 15320 36076
rect 15556 35840 16000 36076
rect 0 35752 16000 35840
rect 0 35516 215 35752
rect 451 35516 537 35752
rect 773 35516 859 35752
rect 1095 35516 1181 35752
rect 1417 35516 1503 35752
rect 1739 35516 1825 35752
rect 2061 35516 2147 35752
rect 2383 35516 2469 35752
rect 2705 35516 2791 35752
rect 3027 35516 3113 35752
rect 3349 35516 3435 35752
rect 3671 35516 3757 35752
rect 3993 35516 4079 35752
rect 4315 35516 4401 35752
rect 4637 35516 4723 35752
rect 4959 35516 5045 35752
rect 5281 35516 5367 35752
rect 5603 35516 5689 35752
rect 5925 35516 6011 35752
rect 6247 35516 6332 35752
rect 6568 35516 6653 35752
rect 6889 35516 6974 35752
rect 7210 35516 7295 35752
rect 7531 35516 7616 35752
rect 7852 35516 7937 35752
rect 8173 35516 8258 35752
rect 8494 35516 8579 35752
rect 8815 35516 8900 35752
rect 9136 35516 9221 35752
rect 9457 35516 9542 35752
rect 9778 35516 9863 35752
rect 10099 35516 10184 35752
rect 10420 35516 10505 35752
rect 10741 35516 10826 35752
rect 11062 35516 11147 35752
rect 11383 35516 11468 35752
rect 11704 35516 11789 35752
rect 12025 35516 12110 35752
rect 12346 35516 12431 35752
rect 12667 35516 12752 35752
rect 12988 35516 13073 35752
rect 13309 35516 13394 35752
rect 13630 35516 13715 35752
rect 13951 35516 14036 35752
rect 14272 35516 14357 35752
rect 14593 35516 14678 35752
rect 14914 35516 14999 35752
rect 15235 35516 15320 35752
rect 15556 35516 16000 35752
rect 0 35428 16000 35516
rect 0 35192 215 35428
rect 451 35192 537 35428
rect 773 35192 859 35428
rect 1095 35192 1181 35428
rect 1417 35192 1503 35428
rect 1739 35192 1825 35428
rect 2061 35192 2147 35428
rect 2383 35192 2469 35428
rect 2705 35192 2791 35428
rect 3027 35192 3113 35428
rect 3349 35192 3435 35428
rect 3671 35192 3757 35428
rect 3993 35192 4079 35428
rect 4315 35192 4401 35428
rect 4637 35192 4723 35428
rect 4959 35192 5045 35428
rect 5281 35192 5367 35428
rect 5603 35192 5689 35428
rect 5925 35192 6011 35428
rect 6247 35192 6332 35428
rect 6568 35192 6653 35428
rect 6889 35192 6974 35428
rect 7210 35192 7295 35428
rect 7531 35192 7616 35428
rect 7852 35192 7937 35428
rect 8173 35192 8258 35428
rect 8494 35192 8579 35428
rect 8815 35192 8900 35428
rect 9136 35192 9221 35428
rect 9457 35192 9542 35428
rect 9778 35192 9863 35428
rect 10099 35192 10184 35428
rect 10420 35192 10505 35428
rect 10741 35192 10826 35428
rect 11062 35192 11147 35428
rect 11383 35192 11468 35428
rect 11704 35192 11789 35428
rect 12025 35192 12110 35428
rect 12346 35192 12431 35428
rect 12667 35192 12752 35428
rect 12988 35192 13073 35428
rect 13309 35192 13394 35428
rect 13630 35192 13715 35428
rect 13951 35192 14036 35428
rect 14272 35192 14357 35428
rect 14593 35192 14678 35428
rect 14914 35192 14999 35428
rect 15235 35192 15320 35428
rect 15556 35192 16000 35428
rect 0 35157 16000 35192
rect 0 18972 16000 18997
rect 0 18736 215 18972
rect 451 18736 538 18972
rect 774 18736 861 18972
rect 1097 18736 1184 18972
rect 1420 18736 1507 18972
rect 1743 18736 1830 18972
rect 2066 18736 2153 18972
rect 2389 18736 2476 18972
rect 2712 18736 2799 18972
rect 3035 18736 3122 18972
rect 3358 18736 3445 18972
rect 3681 18736 3768 18972
rect 4004 18736 4091 18972
rect 4327 18736 4414 18972
rect 4650 18736 4737 18972
rect 4973 18736 5060 18972
rect 5296 18736 5383 18972
rect 5619 18736 5706 18972
rect 5942 18736 6029 18972
rect 6265 18736 6351 18972
rect 6587 18736 6673 18972
rect 6909 18736 6995 18972
rect 7231 18736 7317 18972
rect 7553 18736 7639 18972
rect 7875 18736 7961 18972
rect 8197 18736 8283 18972
rect 8519 18736 8605 18972
rect 8841 18736 8927 18972
rect 9163 18736 9249 18972
rect 9485 18736 9571 18972
rect 9807 18736 9893 18972
rect 10129 18736 10215 18972
rect 10451 18736 10537 18972
rect 10773 18736 10859 18972
rect 11095 18736 11181 18972
rect 11417 18736 11503 18972
rect 11739 18736 11825 18972
rect 12061 18736 12147 18972
rect 12383 18736 12469 18972
rect 12705 18736 12791 18972
rect 13027 18736 13113 18972
rect 13349 18736 13435 18972
rect 13671 18736 13757 18972
rect 13993 18736 14079 18972
rect 14315 18736 14401 18972
rect 14637 18736 14723 18972
rect 14959 18736 15045 18972
rect 15281 18736 15367 18972
rect 15603 18736 16000 18972
rect 0 18636 16000 18736
rect 0 18400 215 18636
rect 451 18400 538 18636
rect 774 18400 861 18636
rect 1097 18400 1184 18636
rect 1420 18400 1507 18636
rect 1743 18400 1830 18636
rect 2066 18400 2153 18636
rect 2389 18400 2476 18636
rect 2712 18400 2799 18636
rect 3035 18400 3122 18636
rect 3358 18400 3445 18636
rect 3681 18400 3768 18636
rect 4004 18400 4091 18636
rect 4327 18400 4414 18636
rect 4650 18400 4737 18636
rect 4973 18400 5060 18636
rect 5296 18400 5383 18636
rect 5619 18400 5706 18636
rect 5942 18400 6029 18636
rect 6265 18400 6351 18636
rect 6587 18400 6673 18636
rect 6909 18400 6995 18636
rect 7231 18400 7317 18636
rect 7553 18400 7639 18636
rect 7875 18400 7961 18636
rect 8197 18400 8283 18636
rect 8519 18400 8605 18636
rect 8841 18400 8927 18636
rect 9163 18400 9249 18636
rect 9485 18400 9571 18636
rect 9807 18400 9893 18636
rect 10129 18400 10215 18636
rect 10451 18400 10537 18636
rect 10773 18400 10859 18636
rect 11095 18400 11181 18636
rect 11417 18400 11503 18636
rect 11739 18400 11825 18636
rect 12061 18400 12147 18636
rect 12383 18400 12469 18636
rect 12705 18400 12791 18636
rect 13027 18400 13113 18636
rect 13349 18400 13435 18636
rect 13671 18400 13757 18636
rect 13993 18400 14079 18636
rect 14315 18400 14401 18636
rect 14637 18400 14723 18636
rect 14959 18400 15045 18636
rect 15281 18400 15367 18636
rect 15603 18400 16000 18636
rect 0 18300 16000 18400
rect 0 18064 215 18300
rect 451 18064 538 18300
rect 774 18064 861 18300
rect 1097 18064 1184 18300
rect 1420 18064 1507 18300
rect 1743 18064 1830 18300
rect 2066 18064 2153 18300
rect 2389 18064 2476 18300
rect 2712 18064 2799 18300
rect 3035 18064 3122 18300
rect 3358 18064 3445 18300
rect 3681 18064 3768 18300
rect 4004 18064 4091 18300
rect 4327 18064 4414 18300
rect 4650 18064 4737 18300
rect 4973 18064 5060 18300
rect 5296 18064 5383 18300
rect 5619 18064 5706 18300
rect 5942 18064 6029 18300
rect 6265 18064 6351 18300
rect 6587 18064 6673 18300
rect 6909 18064 6995 18300
rect 7231 18064 7317 18300
rect 7553 18064 7639 18300
rect 7875 18064 7961 18300
rect 8197 18064 8283 18300
rect 8519 18064 8605 18300
rect 8841 18064 8927 18300
rect 9163 18064 9249 18300
rect 9485 18064 9571 18300
rect 9807 18064 9893 18300
rect 10129 18064 10215 18300
rect 10451 18064 10537 18300
rect 10773 18064 10859 18300
rect 11095 18064 11181 18300
rect 11417 18064 11503 18300
rect 11739 18064 11825 18300
rect 12061 18064 12147 18300
rect 12383 18064 12469 18300
rect 12705 18064 12791 18300
rect 13027 18064 13113 18300
rect 13349 18064 13435 18300
rect 13671 18064 13757 18300
rect 13993 18064 14079 18300
rect 14315 18064 14401 18300
rect 14637 18064 14723 18300
rect 14959 18064 15045 18300
rect 15281 18064 15367 18300
rect 15603 18064 16000 18300
rect 0 17964 16000 18064
rect 0 17728 215 17964
rect 451 17728 538 17964
rect 774 17728 861 17964
rect 1097 17728 1184 17964
rect 1420 17728 1507 17964
rect 1743 17728 1830 17964
rect 2066 17728 2153 17964
rect 2389 17728 2476 17964
rect 2712 17728 2799 17964
rect 3035 17728 3122 17964
rect 3358 17728 3445 17964
rect 3681 17728 3768 17964
rect 4004 17728 4091 17964
rect 4327 17728 4414 17964
rect 4650 17728 4737 17964
rect 4973 17728 5060 17964
rect 5296 17728 5383 17964
rect 5619 17728 5706 17964
rect 5942 17728 6029 17964
rect 6265 17728 6351 17964
rect 6587 17728 6673 17964
rect 6909 17728 6995 17964
rect 7231 17728 7317 17964
rect 7553 17728 7639 17964
rect 7875 17728 7961 17964
rect 8197 17728 8283 17964
rect 8519 17728 8605 17964
rect 8841 17728 8927 17964
rect 9163 17728 9249 17964
rect 9485 17728 9571 17964
rect 9807 17728 9893 17964
rect 10129 17728 10215 17964
rect 10451 17728 10537 17964
rect 10773 17728 10859 17964
rect 11095 17728 11181 17964
rect 11417 17728 11503 17964
rect 11739 17728 11825 17964
rect 12061 17728 12147 17964
rect 12383 17728 12469 17964
rect 12705 17728 12791 17964
rect 13027 17728 13113 17964
rect 13349 17728 13435 17964
rect 13671 17728 13757 17964
rect 13993 17728 14079 17964
rect 14315 17728 14401 17964
rect 14637 17728 14723 17964
rect 14959 17728 15045 17964
rect 15281 17728 15367 17964
rect 15603 17728 16000 17964
rect 0 17628 16000 17728
rect 0 17392 215 17628
rect 451 17392 538 17628
rect 774 17392 861 17628
rect 1097 17392 1184 17628
rect 1420 17392 1507 17628
rect 1743 17392 1830 17628
rect 2066 17392 2153 17628
rect 2389 17392 2476 17628
rect 2712 17392 2799 17628
rect 3035 17392 3122 17628
rect 3358 17392 3445 17628
rect 3681 17392 3768 17628
rect 4004 17392 4091 17628
rect 4327 17392 4414 17628
rect 4650 17392 4737 17628
rect 4973 17392 5060 17628
rect 5296 17392 5383 17628
rect 5619 17392 5706 17628
rect 5942 17392 6029 17628
rect 6265 17392 6351 17628
rect 6587 17392 6673 17628
rect 6909 17392 6995 17628
rect 7231 17392 7317 17628
rect 7553 17392 7639 17628
rect 7875 17392 7961 17628
rect 8197 17392 8283 17628
rect 8519 17392 8605 17628
rect 8841 17392 8927 17628
rect 9163 17392 9249 17628
rect 9485 17392 9571 17628
rect 9807 17392 9893 17628
rect 10129 17392 10215 17628
rect 10451 17392 10537 17628
rect 10773 17392 10859 17628
rect 11095 17392 11181 17628
rect 11417 17392 11503 17628
rect 11739 17392 11825 17628
rect 12061 17392 12147 17628
rect 12383 17392 12469 17628
rect 12705 17392 12791 17628
rect 13027 17392 13113 17628
rect 13349 17392 13435 17628
rect 13671 17392 13757 17628
rect 13993 17392 14079 17628
rect 14315 17392 14401 17628
rect 14637 17392 14723 17628
rect 14959 17392 15045 17628
rect 15281 17392 15367 17628
rect 15603 17392 16000 17628
rect 0 17292 16000 17392
rect 0 17056 215 17292
rect 451 17056 538 17292
rect 774 17056 861 17292
rect 1097 17056 1184 17292
rect 1420 17056 1507 17292
rect 1743 17056 1830 17292
rect 2066 17056 2153 17292
rect 2389 17056 2476 17292
rect 2712 17056 2799 17292
rect 3035 17056 3122 17292
rect 3358 17056 3445 17292
rect 3681 17056 3768 17292
rect 4004 17056 4091 17292
rect 4327 17056 4414 17292
rect 4650 17056 4737 17292
rect 4973 17056 5060 17292
rect 5296 17056 5383 17292
rect 5619 17056 5706 17292
rect 5942 17056 6029 17292
rect 6265 17056 6351 17292
rect 6587 17056 6673 17292
rect 6909 17056 6995 17292
rect 7231 17056 7317 17292
rect 7553 17056 7639 17292
rect 7875 17056 7961 17292
rect 8197 17056 8283 17292
rect 8519 17056 8605 17292
rect 8841 17056 8927 17292
rect 9163 17056 9249 17292
rect 9485 17056 9571 17292
rect 9807 17056 9893 17292
rect 10129 17056 10215 17292
rect 10451 17056 10537 17292
rect 10773 17056 10859 17292
rect 11095 17056 11181 17292
rect 11417 17056 11503 17292
rect 11739 17056 11825 17292
rect 12061 17056 12147 17292
rect 12383 17056 12469 17292
rect 12705 17056 12791 17292
rect 13027 17056 13113 17292
rect 13349 17056 13435 17292
rect 13671 17056 13757 17292
rect 13993 17056 14079 17292
rect 14315 17056 14401 17292
rect 14637 17056 14723 17292
rect 14959 17056 15045 17292
rect 15281 17056 15367 17292
rect 15603 17056 16000 17292
rect 0 16956 16000 17056
rect 0 16720 215 16956
rect 451 16720 538 16956
rect 774 16720 861 16956
rect 1097 16720 1184 16956
rect 1420 16720 1507 16956
rect 1743 16720 1830 16956
rect 2066 16720 2153 16956
rect 2389 16720 2476 16956
rect 2712 16720 2799 16956
rect 3035 16720 3122 16956
rect 3358 16720 3445 16956
rect 3681 16720 3768 16956
rect 4004 16720 4091 16956
rect 4327 16720 4414 16956
rect 4650 16720 4737 16956
rect 4973 16720 5060 16956
rect 5296 16720 5383 16956
rect 5619 16720 5706 16956
rect 5942 16720 6029 16956
rect 6265 16720 6351 16956
rect 6587 16720 6673 16956
rect 6909 16720 6995 16956
rect 7231 16720 7317 16956
rect 7553 16720 7639 16956
rect 7875 16720 7961 16956
rect 8197 16720 8283 16956
rect 8519 16720 8605 16956
rect 8841 16720 8927 16956
rect 9163 16720 9249 16956
rect 9485 16720 9571 16956
rect 9807 16720 9893 16956
rect 10129 16720 10215 16956
rect 10451 16720 10537 16956
rect 10773 16720 10859 16956
rect 11095 16720 11181 16956
rect 11417 16720 11503 16956
rect 11739 16720 11825 16956
rect 12061 16720 12147 16956
rect 12383 16720 12469 16956
rect 12705 16720 12791 16956
rect 13027 16720 13113 16956
rect 13349 16720 13435 16956
rect 13671 16720 13757 16956
rect 13993 16720 14079 16956
rect 14315 16720 14401 16956
rect 14637 16720 14723 16956
rect 14959 16720 15045 16956
rect 15281 16720 15367 16956
rect 15603 16720 16000 16956
rect 0 16620 16000 16720
rect 0 16384 215 16620
rect 451 16384 538 16620
rect 774 16384 861 16620
rect 1097 16384 1184 16620
rect 1420 16384 1507 16620
rect 1743 16384 1830 16620
rect 2066 16384 2153 16620
rect 2389 16384 2476 16620
rect 2712 16384 2799 16620
rect 3035 16384 3122 16620
rect 3358 16384 3445 16620
rect 3681 16384 3768 16620
rect 4004 16384 4091 16620
rect 4327 16384 4414 16620
rect 4650 16384 4737 16620
rect 4973 16384 5060 16620
rect 5296 16384 5383 16620
rect 5619 16384 5706 16620
rect 5942 16384 6029 16620
rect 6265 16384 6351 16620
rect 6587 16384 6673 16620
rect 6909 16384 6995 16620
rect 7231 16384 7317 16620
rect 7553 16384 7639 16620
rect 7875 16384 7961 16620
rect 8197 16384 8283 16620
rect 8519 16384 8605 16620
rect 8841 16384 8927 16620
rect 9163 16384 9249 16620
rect 9485 16384 9571 16620
rect 9807 16384 9893 16620
rect 10129 16384 10215 16620
rect 10451 16384 10537 16620
rect 10773 16384 10859 16620
rect 11095 16384 11181 16620
rect 11417 16384 11503 16620
rect 11739 16384 11825 16620
rect 12061 16384 12147 16620
rect 12383 16384 12469 16620
rect 12705 16384 12791 16620
rect 13027 16384 13113 16620
rect 13349 16384 13435 16620
rect 13671 16384 13757 16620
rect 13993 16384 14079 16620
rect 14315 16384 14401 16620
rect 14637 16384 14723 16620
rect 14959 16384 15045 16620
rect 15281 16384 15367 16620
rect 15603 16384 16000 16620
rect 0 16284 16000 16384
rect 0 16048 215 16284
rect 451 16048 538 16284
rect 774 16048 861 16284
rect 1097 16048 1184 16284
rect 1420 16048 1507 16284
rect 1743 16048 1830 16284
rect 2066 16048 2153 16284
rect 2389 16048 2476 16284
rect 2712 16048 2799 16284
rect 3035 16048 3122 16284
rect 3358 16048 3445 16284
rect 3681 16048 3768 16284
rect 4004 16048 4091 16284
rect 4327 16048 4414 16284
rect 4650 16048 4737 16284
rect 4973 16048 5060 16284
rect 5296 16048 5383 16284
rect 5619 16048 5706 16284
rect 5942 16048 6029 16284
rect 6265 16048 6351 16284
rect 6587 16048 6673 16284
rect 6909 16048 6995 16284
rect 7231 16048 7317 16284
rect 7553 16048 7639 16284
rect 7875 16048 7961 16284
rect 8197 16048 8283 16284
rect 8519 16048 8605 16284
rect 8841 16048 8927 16284
rect 9163 16048 9249 16284
rect 9485 16048 9571 16284
rect 9807 16048 9893 16284
rect 10129 16048 10215 16284
rect 10451 16048 10537 16284
rect 10773 16048 10859 16284
rect 11095 16048 11181 16284
rect 11417 16048 11503 16284
rect 11739 16048 11825 16284
rect 12061 16048 12147 16284
rect 12383 16048 12469 16284
rect 12705 16048 12791 16284
rect 13027 16048 13113 16284
rect 13349 16048 13435 16284
rect 13671 16048 13757 16284
rect 13993 16048 14079 16284
rect 14315 16048 14401 16284
rect 14637 16048 14723 16284
rect 14959 16048 15045 16284
rect 15281 16048 15367 16284
rect 15603 16048 16000 16284
rect 0 15948 16000 16048
rect 0 15712 215 15948
rect 451 15712 538 15948
rect 774 15712 861 15948
rect 1097 15712 1184 15948
rect 1420 15712 1507 15948
rect 1743 15712 1830 15948
rect 2066 15712 2153 15948
rect 2389 15712 2476 15948
rect 2712 15712 2799 15948
rect 3035 15712 3122 15948
rect 3358 15712 3445 15948
rect 3681 15712 3768 15948
rect 4004 15712 4091 15948
rect 4327 15712 4414 15948
rect 4650 15712 4737 15948
rect 4973 15712 5060 15948
rect 5296 15712 5383 15948
rect 5619 15712 5706 15948
rect 5942 15712 6029 15948
rect 6265 15712 6351 15948
rect 6587 15712 6673 15948
rect 6909 15712 6995 15948
rect 7231 15712 7317 15948
rect 7553 15712 7639 15948
rect 7875 15712 7961 15948
rect 8197 15712 8283 15948
rect 8519 15712 8605 15948
rect 8841 15712 8927 15948
rect 9163 15712 9249 15948
rect 9485 15712 9571 15948
rect 9807 15712 9893 15948
rect 10129 15712 10215 15948
rect 10451 15712 10537 15948
rect 10773 15712 10859 15948
rect 11095 15712 11181 15948
rect 11417 15712 11503 15948
rect 11739 15712 11825 15948
rect 12061 15712 12147 15948
rect 12383 15712 12469 15948
rect 12705 15712 12791 15948
rect 13027 15712 13113 15948
rect 13349 15712 13435 15948
rect 13671 15712 13757 15948
rect 13993 15712 14079 15948
rect 14315 15712 14401 15948
rect 14637 15712 14723 15948
rect 14959 15712 15045 15948
rect 15281 15712 15367 15948
rect 15603 15712 16000 15948
rect 0 15612 16000 15712
rect 0 15376 215 15612
rect 451 15376 538 15612
rect 774 15376 861 15612
rect 1097 15376 1184 15612
rect 1420 15376 1507 15612
rect 1743 15376 1830 15612
rect 2066 15376 2153 15612
rect 2389 15376 2476 15612
rect 2712 15376 2799 15612
rect 3035 15376 3122 15612
rect 3358 15376 3445 15612
rect 3681 15376 3768 15612
rect 4004 15376 4091 15612
rect 4327 15376 4414 15612
rect 4650 15376 4737 15612
rect 4973 15376 5060 15612
rect 5296 15376 5383 15612
rect 5619 15376 5706 15612
rect 5942 15376 6029 15612
rect 6265 15376 6351 15612
rect 6587 15376 6673 15612
rect 6909 15376 6995 15612
rect 7231 15376 7317 15612
rect 7553 15376 7639 15612
rect 7875 15376 7961 15612
rect 8197 15376 8283 15612
rect 8519 15376 8605 15612
rect 8841 15376 8927 15612
rect 9163 15376 9249 15612
rect 9485 15376 9571 15612
rect 9807 15376 9893 15612
rect 10129 15376 10215 15612
rect 10451 15376 10537 15612
rect 10773 15376 10859 15612
rect 11095 15376 11181 15612
rect 11417 15376 11503 15612
rect 11739 15376 11825 15612
rect 12061 15376 12147 15612
rect 12383 15376 12469 15612
rect 12705 15376 12791 15612
rect 13027 15376 13113 15612
rect 13349 15376 13435 15612
rect 13671 15376 13757 15612
rect 13993 15376 14079 15612
rect 14315 15376 14401 15612
rect 14637 15376 14723 15612
rect 14959 15376 15045 15612
rect 15281 15376 15367 15612
rect 15603 15376 16000 15612
rect 0 15276 16000 15376
rect 0 15040 215 15276
rect 451 15040 538 15276
rect 774 15040 861 15276
rect 1097 15040 1184 15276
rect 1420 15040 1507 15276
rect 1743 15040 1830 15276
rect 2066 15040 2153 15276
rect 2389 15040 2476 15276
rect 2712 15040 2799 15276
rect 3035 15040 3122 15276
rect 3358 15040 3445 15276
rect 3681 15040 3768 15276
rect 4004 15040 4091 15276
rect 4327 15040 4414 15276
rect 4650 15040 4737 15276
rect 4973 15040 5060 15276
rect 5296 15040 5383 15276
rect 5619 15040 5706 15276
rect 5942 15040 6029 15276
rect 6265 15040 6351 15276
rect 6587 15040 6673 15276
rect 6909 15040 6995 15276
rect 7231 15040 7317 15276
rect 7553 15040 7639 15276
rect 7875 15040 7961 15276
rect 8197 15040 8283 15276
rect 8519 15040 8605 15276
rect 8841 15040 8927 15276
rect 9163 15040 9249 15276
rect 9485 15040 9571 15276
rect 9807 15040 9893 15276
rect 10129 15040 10215 15276
rect 10451 15040 10537 15276
rect 10773 15040 10859 15276
rect 11095 15040 11181 15276
rect 11417 15040 11503 15276
rect 11739 15040 11825 15276
rect 12061 15040 12147 15276
rect 12383 15040 12469 15276
rect 12705 15040 12791 15276
rect 13027 15040 13113 15276
rect 13349 15040 13435 15276
rect 13671 15040 13757 15276
rect 13993 15040 14079 15276
rect 14315 15040 14401 15276
rect 14637 15040 14723 15276
rect 14959 15040 15045 15276
rect 15281 15040 15367 15276
rect 15603 15040 16000 15276
rect 0 14940 16000 15040
rect 0 14704 215 14940
rect 451 14704 538 14940
rect 774 14704 861 14940
rect 1097 14704 1184 14940
rect 1420 14704 1507 14940
rect 1743 14704 1830 14940
rect 2066 14704 2153 14940
rect 2389 14704 2476 14940
rect 2712 14704 2799 14940
rect 3035 14704 3122 14940
rect 3358 14704 3445 14940
rect 3681 14704 3768 14940
rect 4004 14704 4091 14940
rect 4327 14704 4414 14940
rect 4650 14704 4737 14940
rect 4973 14704 5060 14940
rect 5296 14704 5383 14940
rect 5619 14704 5706 14940
rect 5942 14704 6029 14940
rect 6265 14704 6351 14940
rect 6587 14704 6673 14940
rect 6909 14704 6995 14940
rect 7231 14704 7317 14940
rect 7553 14704 7639 14940
rect 7875 14704 7961 14940
rect 8197 14704 8283 14940
rect 8519 14704 8605 14940
rect 8841 14704 8927 14940
rect 9163 14704 9249 14940
rect 9485 14704 9571 14940
rect 9807 14704 9893 14940
rect 10129 14704 10215 14940
rect 10451 14704 10537 14940
rect 10773 14704 10859 14940
rect 11095 14704 11181 14940
rect 11417 14704 11503 14940
rect 11739 14704 11825 14940
rect 12061 14704 12147 14940
rect 12383 14704 12469 14940
rect 12705 14704 12791 14940
rect 13027 14704 13113 14940
rect 13349 14704 13435 14940
rect 13671 14704 13757 14940
rect 13993 14704 14079 14940
rect 14315 14704 14401 14940
rect 14637 14704 14723 14940
rect 14959 14704 15045 14940
rect 15281 14704 15367 14940
rect 15603 14704 16000 14940
rect 0 14604 16000 14704
rect 0 14368 215 14604
rect 451 14368 538 14604
rect 774 14368 861 14604
rect 1097 14368 1184 14604
rect 1420 14368 1507 14604
rect 1743 14368 1830 14604
rect 2066 14368 2153 14604
rect 2389 14368 2476 14604
rect 2712 14368 2799 14604
rect 3035 14368 3122 14604
rect 3358 14368 3445 14604
rect 3681 14368 3768 14604
rect 4004 14368 4091 14604
rect 4327 14368 4414 14604
rect 4650 14368 4737 14604
rect 4973 14368 5060 14604
rect 5296 14368 5383 14604
rect 5619 14368 5706 14604
rect 5942 14368 6029 14604
rect 6265 14368 6351 14604
rect 6587 14368 6673 14604
rect 6909 14368 6995 14604
rect 7231 14368 7317 14604
rect 7553 14368 7639 14604
rect 7875 14368 7961 14604
rect 8197 14368 8283 14604
rect 8519 14368 8605 14604
rect 8841 14368 8927 14604
rect 9163 14368 9249 14604
rect 9485 14368 9571 14604
rect 9807 14368 9893 14604
rect 10129 14368 10215 14604
rect 10451 14368 10537 14604
rect 10773 14368 10859 14604
rect 11095 14368 11181 14604
rect 11417 14368 11503 14604
rect 11739 14368 11825 14604
rect 12061 14368 12147 14604
rect 12383 14368 12469 14604
rect 12705 14368 12791 14604
rect 13027 14368 13113 14604
rect 13349 14368 13435 14604
rect 13671 14368 13757 14604
rect 13993 14368 14079 14604
rect 14315 14368 14401 14604
rect 14637 14368 14723 14604
rect 14959 14368 15045 14604
rect 15281 14368 15367 14604
rect 15603 14368 16000 14604
rect 0 14268 16000 14368
rect 0 14032 215 14268
rect 451 14032 538 14268
rect 774 14032 861 14268
rect 1097 14032 1184 14268
rect 1420 14032 1507 14268
rect 1743 14032 1830 14268
rect 2066 14032 2153 14268
rect 2389 14032 2476 14268
rect 2712 14032 2799 14268
rect 3035 14032 3122 14268
rect 3358 14032 3445 14268
rect 3681 14032 3768 14268
rect 4004 14032 4091 14268
rect 4327 14032 4414 14268
rect 4650 14032 4737 14268
rect 4973 14032 5060 14268
rect 5296 14032 5383 14268
rect 5619 14032 5706 14268
rect 5942 14032 6029 14268
rect 6265 14032 6351 14268
rect 6587 14032 6673 14268
rect 6909 14032 6995 14268
rect 7231 14032 7317 14268
rect 7553 14032 7639 14268
rect 7875 14032 7961 14268
rect 8197 14032 8283 14268
rect 8519 14032 8605 14268
rect 8841 14032 8927 14268
rect 9163 14032 9249 14268
rect 9485 14032 9571 14268
rect 9807 14032 9893 14268
rect 10129 14032 10215 14268
rect 10451 14032 10537 14268
rect 10773 14032 10859 14268
rect 11095 14032 11181 14268
rect 11417 14032 11503 14268
rect 11739 14032 11825 14268
rect 12061 14032 12147 14268
rect 12383 14032 12469 14268
rect 12705 14032 12791 14268
rect 13027 14032 13113 14268
rect 13349 14032 13435 14268
rect 13671 14032 13757 14268
rect 13993 14032 14079 14268
rect 14315 14032 14401 14268
rect 14637 14032 14723 14268
rect 14959 14032 15045 14268
rect 15281 14032 15367 14268
rect 15603 14032 16000 14268
rect 0 14007 16000 14032
rect 0 13663 16000 13687
rect 0 13427 216 13663
rect 452 13427 538 13663
rect 774 13427 860 13663
rect 1096 13427 1182 13663
rect 1418 13427 1504 13663
rect 1740 13427 1826 13663
rect 2062 13427 2148 13663
rect 2384 13427 2470 13663
rect 2706 13427 2792 13663
rect 3028 13427 3114 13663
rect 3350 13427 3436 13663
rect 3672 13427 3758 13663
rect 3994 13427 4080 13663
rect 4316 13427 4402 13663
rect 4638 13427 4724 13663
rect 4960 13427 5046 13663
rect 5282 13427 5368 13663
rect 5604 13427 5690 13663
rect 5926 13427 6012 13663
rect 6248 13427 6333 13663
rect 6569 13427 6654 13663
rect 6890 13427 6975 13663
rect 7211 13427 7296 13663
rect 7532 13427 7617 13663
rect 7853 13427 7938 13663
rect 8174 13427 8259 13663
rect 8495 13427 8580 13663
rect 8816 13427 8901 13663
rect 9137 13427 9222 13663
rect 9458 13427 9543 13663
rect 9779 13427 9864 13663
rect 10100 13427 10185 13663
rect 10421 13427 10506 13663
rect 10742 13427 10827 13663
rect 11063 13427 11148 13663
rect 11384 13427 11469 13663
rect 11705 13427 11790 13663
rect 12026 13427 12111 13663
rect 12347 13427 12432 13663
rect 12668 13427 12753 13663
rect 12989 13427 13074 13663
rect 13310 13427 13395 13663
rect 13631 13427 13716 13663
rect 13952 13427 14037 13663
rect 14273 13427 14358 13663
rect 14594 13427 14679 13663
rect 14915 13427 15000 13663
rect 15236 13427 15321 13663
rect 15557 13427 16000 13663
rect 0 13097 16000 13427
rect 0 12861 216 13097
rect 452 12861 538 13097
rect 774 12861 860 13097
rect 1096 12861 1182 13097
rect 1418 12861 1504 13097
rect 1740 12861 1826 13097
rect 2062 12861 2148 13097
rect 2384 12861 2470 13097
rect 2706 12861 2792 13097
rect 3028 12861 3114 13097
rect 3350 12861 3436 13097
rect 3672 12861 3758 13097
rect 3994 12861 4080 13097
rect 4316 12861 4402 13097
rect 4638 12861 4724 13097
rect 4960 12861 5046 13097
rect 5282 12861 5368 13097
rect 5604 12861 5690 13097
rect 5926 12861 6012 13097
rect 6248 12861 6333 13097
rect 6569 12861 6654 13097
rect 6890 12861 6975 13097
rect 7211 12861 7296 13097
rect 7532 12861 7617 13097
rect 7853 12861 7938 13097
rect 8174 12861 8259 13097
rect 8495 12861 8580 13097
rect 8816 12861 8901 13097
rect 9137 12861 9222 13097
rect 9458 12861 9543 13097
rect 9779 12861 9864 13097
rect 10100 12861 10185 13097
rect 10421 12861 10506 13097
rect 10742 12861 10827 13097
rect 11063 12861 11148 13097
rect 11384 12861 11469 13097
rect 11705 12861 11790 13097
rect 12026 12861 12111 13097
rect 12347 12861 12432 13097
rect 12668 12861 12753 13097
rect 12989 12861 13074 13097
rect 13310 12861 13395 13097
rect 13631 12861 13716 13097
rect 13952 12861 14037 13097
rect 14273 12861 14358 13097
rect 14594 12861 14679 13097
rect 14915 12861 15000 13097
rect 15236 12861 15321 13097
rect 15557 12861 16000 13097
rect 0 12837 16000 12861
rect 0 12493 16000 12517
rect 0 12257 215 12493
rect 451 12257 537 12493
rect 773 12257 859 12493
rect 1095 12257 1181 12493
rect 1417 12257 1503 12493
rect 1739 12257 1825 12493
rect 2061 12257 2147 12493
rect 2383 12257 2469 12493
rect 2705 12257 2791 12493
rect 3027 12257 3113 12493
rect 3349 12257 3435 12493
rect 3671 12257 3757 12493
rect 3993 12257 4079 12493
rect 4315 12257 4401 12493
rect 4637 12257 4723 12493
rect 4959 12257 5045 12493
rect 5281 12257 5367 12493
rect 5603 12257 5689 12493
rect 5925 12257 6011 12493
rect 6247 12257 6332 12493
rect 6568 12257 6653 12493
rect 6889 12257 6974 12493
rect 7210 12257 7295 12493
rect 7531 12257 7616 12493
rect 7852 12257 7937 12493
rect 8173 12257 8258 12493
rect 8494 12257 8579 12493
rect 8815 12257 8900 12493
rect 9136 12257 9221 12493
rect 9457 12257 9542 12493
rect 9778 12257 9863 12493
rect 10099 12257 10184 12493
rect 10420 12257 10505 12493
rect 10741 12257 10826 12493
rect 11062 12257 11147 12493
rect 11383 12257 11468 12493
rect 11704 12257 11789 12493
rect 12025 12257 12110 12493
rect 12346 12257 12431 12493
rect 12667 12257 12752 12493
rect 12988 12257 13073 12493
rect 13309 12257 13394 12493
rect 13630 12257 13715 12493
rect 13951 12257 14036 12493
rect 14272 12257 14357 12493
rect 14593 12257 14678 12493
rect 14914 12257 14999 12493
rect 15235 12257 15320 12493
rect 15556 12257 16000 12493
rect 0 11927 16000 12257
rect 0 11691 215 11927
rect 451 11691 537 11927
rect 773 11691 859 11927
rect 1095 11691 1181 11927
rect 1417 11691 1503 11927
rect 1739 11691 1825 11927
rect 2061 11691 2147 11927
rect 2383 11691 2469 11927
rect 2705 11691 2791 11927
rect 3027 11691 3113 11927
rect 3349 11691 3435 11927
rect 3671 11691 3757 11927
rect 3993 11691 4079 11927
rect 4315 11691 4401 11927
rect 4637 11691 4723 11927
rect 4959 11691 5045 11927
rect 5281 11691 5367 11927
rect 5603 11691 5689 11927
rect 5925 11691 6011 11927
rect 6247 11691 6332 11927
rect 6568 11691 6653 11927
rect 6889 11691 6974 11927
rect 7210 11691 7295 11927
rect 7531 11691 7616 11927
rect 7852 11691 7937 11927
rect 8173 11691 8258 11927
rect 8494 11691 8579 11927
rect 8815 11691 8900 11927
rect 9136 11691 9221 11927
rect 9457 11691 9542 11927
rect 9778 11691 9863 11927
rect 10099 11691 10184 11927
rect 10420 11691 10505 11927
rect 10741 11691 10826 11927
rect 11062 11691 11147 11927
rect 11383 11691 11468 11927
rect 11704 11691 11789 11927
rect 12025 11691 12110 11927
rect 12346 11691 12431 11927
rect 12667 11691 12752 11927
rect 12988 11691 13073 11927
rect 13309 11691 13394 11927
rect 13630 11691 13715 11927
rect 13951 11691 14036 11927
rect 14272 11691 14357 11927
rect 14593 11691 14678 11927
rect 14914 11691 14999 11927
rect 15235 11691 15320 11927
rect 15556 11691 16000 11927
rect 0 11667 16000 11691
rect 0 10565 16000 11347
rect 0 10329 215 10565
rect 451 10329 537 10565
rect 773 10329 859 10565
rect 1095 10329 1181 10565
rect 1417 10329 1503 10565
rect 1739 10329 1825 10565
rect 2061 10329 2147 10565
rect 2383 10329 2469 10565
rect 2705 10329 2791 10565
rect 3027 10329 3113 10565
rect 3349 10329 3435 10565
rect 3671 10329 3757 10565
rect 3993 10329 4079 10565
rect 4315 10329 4401 10565
rect 4637 10329 4723 10565
rect 4959 10329 5045 10565
rect 5281 10329 5367 10565
rect 5603 10329 5689 10565
rect 5925 10329 6011 10565
rect 6247 10329 6332 10565
rect 6568 10329 6653 10565
rect 6889 10329 6974 10565
rect 7210 10329 7295 10565
rect 7531 10329 7616 10565
rect 7852 10329 7937 10565
rect 8173 10329 8258 10565
rect 8494 10329 8579 10565
rect 8815 10329 8900 10565
rect 9136 10329 9221 10565
rect 9457 10329 9542 10565
rect 9778 10329 9863 10565
rect 10099 10329 10184 10565
rect 10420 10329 10505 10565
rect 10741 10329 10826 10565
rect 11062 10329 11147 10565
rect 11383 10329 11468 10565
rect 11704 10329 11789 10565
rect 12025 10329 12110 10565
rect 12346 10329 12431 10565
rect 12667 10329 12752 10565
rect 12988 10329 13073 10565
rect 13309 10329 13394 10565
rect 13630 10329 13715 10565
rect 13951 10329 14036 10565
rect 14272 10329 14357 10565
rect 14593 10329 14678 10565
rect 14914 10329 14999 10565
rect 15235 10329 15320 10565
rect 15556 10329 16000 10565
rect 0 9547 16000 10329
rect 0 9203 16000 9227
rect 0 8967 216 9203
rect 452 8967 538 9203
rect 774 8967 860 9203
rect 1096 8967 1182 9203
rect 1418 8967 1504 9203
rect 1740 8967 1826 9203
rect 2062 8967 2148 9203
rect 2384 8967 2470 9203
rect 2706 8967 2792 9203
rect 3028 8967 3114 9203
rect 3350 8967 3436 9203
rect 3672 8967 3758 9203
rect 3994 8967 4080 9203
rect 4316 8967 4402 9203
rect 4638 8967 4724 9203
rect 4960 8967 5046 9203
rect 5282 8967 5368 9203
rect 5604 8967 5690 9203
rect 5926 8967 6012 9203
rect 6248 8967 6333 9203
rect 6569 8967 6654 9203
rect 6890 8967 6975 9203
rect 7211 8967 7296 9203
rect 7532 8967 7617 9203
rect 7853 8967 7938 9203
rect 8174 8967 8259 9203
rect 8495 8967 8580 9203
rect 8816 8967 8901 9203
rect 9137 8967 9222 9203
rect 9458 8967 9543 9203
rect 9779 8967 9864 9203
rect 10100 8967 10185 9203
rect 10421 8967 10506 9203
rect 10742 8967 10827 9203
rect 11063 8967 11148 9203
rect 11384 8967 11469 9203
rect 11705 8967 11790 9203
rect 12026 8967 12111 9203
rect 12347 8967 12432 9203
rect 12668 8967 12753 9203
rect 12989 8967 13074 9203
rect 13310 8967 13395 9203
rect 13631 8967 13716 9203
rect 13952 8967 14037 9203
rect 14273 8967 14358 9203
rect 14594 8967 14679 9203
rect 14915 8967 15000 9203
rect 15236 8967 15321 9203
rect 15557 8967 16000 9203
rect 0 8597 16000 8967
rect 0 8361 216 8597
rect 452 8361 538 8597
rect 774 8361 860 8597
rect 1096 8361 1182 8597
rect 1418 8361 1504 8597
rect 1740 8361 1826 8597
rect 2062 8361 2148 8597
rect 2384 8361 2470 8597
rect 2706 8361 2792 8597
rect 3028 8361 3114 8597
rect 3350 8361 3436 8597
rect 3672 8361 3758 8597
rect 3994 8361 4080 8597
rect 4316 8361 4402 8597
rect 4638 8361 4724 8597
rect 4960 8361 5046 8597
rect 5282 8361 5368 8597
rect 5604 8361 5690 8597
rect 5926 8361 6012 8597
rect 6248 8361 6333 8597
rect 6569 8361 6654 8597
rect 6890 8361 6975 8597
rect 7211 8361 7296 8597
rect 7532 8361 7617 8597
rect 7853 8361 7938 8597
rect 8174 8361 8259 8597
rect 8495 8361 8580 8597
rect 8816 8361 8901 8597
rect 9137 8361 9222 8597
rect 9458 8361 9543 8597
rect 9779 8361 9864 8597
rect 10100 8361 10185 8597
rect 10421 8361 10506 8597
rect 10742 8361 10827 8597
rect 11063 8361 11148 8597
rect 11384 8361 11469 8597
rect 11705 8361 11790 8597
rect 12026 8361 12111 8597
rect 12347 8361 12432 8597
rect 12668 8361 12753 8597
rect 12989 8361 13074 8597
rect 13310 8361 13395 8597
rect 13631 8361 13716 8597
rect 13952 8361 14037 8597
rect 14273 8361 14358 8597
rect 14594 8361 14679 8597
rect 14915 8361 15000 8597
rect 15236 8361 15321 8597
rect 15557 8361 16000 8597
rect 0 8337 16000 8361
rect 0 7993 16000 8017
rect 0 7757 215 7993
rect 451 7757 537 7993
rect 773 7757 859 7993
rect 1095 7757 1181 7993
rect 1417 7757 1503 7993
rect 1739 7757 1825 7993
rect 2061 7757 2147 7993
rect 2383 7757 2469 7993
rect 2705 7757 2791 7993
rect 3027 7757 3113 7993
rect 3349 7757 3435 7993
rect 3671 7757 3757 7993
rect 3993 7757 4079 7993
rect 4315 7757 4401 7993
rect 4637 7757 4723 7993
rect 4959 7757 5045 7993
rect 5281 7757 5367 7993
rect 5603 7757 5689 7993
rect 5925 7757 6011 7993
rect 6247 7757 6332 7993
rect 6568 7757 6653 7993
rect 6889 7757 6974 7993
rect 7210 7757 7295 7993
rect 7531 7757 7616 7993
rect 7852 7757 7937 7993
rect 8173 7757 8258 7993
rect 8494 7757 8579 7993
rect 8815 7757 8900 7993
rect 9136 7757 9221 7993
rect 9457 7757 9542 7993
rect 9778 7757 9863 7993
rect 10099 7757 10184 7993
rect 10420 7757 10505 7993
rect 10741 7757 10826 7993
rect 11062 7757 11147 7993
rect 11383 7757 11468 7993
rect 11704 7757 11789 7993
rect 12025 7757 12110 7993
rect 12346 7757 12431 7993
rect 12667 7757 12752 7993
rect 12988 7757 13073 7993
rect 13309 7757 13394 7993
rect 13630 7757 13715 7993
rect 13951 7757 14036 7993
rect 14272 7757 14357 7993
rect 14593 7757 14678 7993
rect 14914 7757 14999 7993
rect 15235 7757 15320 7993
rect 15556 7757 16000 7993
rect 0 7627 16000 7757
rect 0 7391 215 7627
rect 451 7391 537 7627
rect 773 7391 859 7627
rect 1095 7391 1181 7627
rect 1417 7391 1503 7627
rect 1739 7391 1825 7627
rect 2061 7391 2147 7627
rect 2383 7391 2469 7627
rect 2705 7391 2791 7627
rect 3027 7391 3113 7627
rect 3349 7391 3435 7627
rect 3671 7391 3757 7627
rect 3993 7391 4079 7627
rect 4315 7391 4401 7627
rect 4637 7391 4723 7627
rect 4959 7391 5045 7627
rect 5281 7391 5367 7627
rect 5603 7391 5689 7627
rect 5925 7391 6011 7627
rect 6247 7391 6332 7627
rect 6568 7391 6653 7627
rect 6889 7391 6974 7627
rect 7210 7391 7295 7627
rect 7531 7391 7616 7627
rect 7852 7391 7937 7627
rect 8173 7391 8258 7627
rect 8494 7391 8579 7627
rect 8815 7391 8900 7627
rect 9136 7391 9221 7627
rect 9457 7391 9542 7627
rect 9778 7391 9863 7627
rect 10099 7391 10184 7627
rect 10420 7391 10505 7627
rect 10741 7391 10826 7627
rect 11062 7391 11147 7627
rect 11383 7391 11468 7627
rect 11704 7391 11789 7627
rect 12025 7391 12110 7627
rect 12346 7391 12431 7627
rect 12667 7391 12752 7627
rect 12988 7391 13073 7627
rect 13309 7391 13394 7627
rect 13630 7391 13715 7627
rect 13951 7391 14036 7627
rect 14272 7391 14357 7627
rect 14593 7391 14678 7627
rect 14914 7391 14999 7627
rect 15235 7391 15320 7627
rect 15556 7391 16000 7627
rect 0 7367 16000 7391
rect 0 7023 16000 7047
rect 0 6787 215 7023
rect 451 6787 537 7023
rect 773 6787 859 7023
rect 1095 6787 1181 7023
rect 1417 6787 1503 7023
rect 1739 6787 1825 7023
rect 2061 6787 2147 7023
rect 2383 6787 2469 7023
rect 2705 6787 2791 7023
rect 3027 6787 3113 7023
rect 3349 6787 3435 7023
rect 3671 6787 3757 7023
rect 3993 6787 4079 7023
rect 4315 6787 4401 7023
rect 4637 6787 4723 7023
rect 4959 6787 5045 7023
rect 5281 6787 5367 7023
rect 5603 6787 5689 7023
rect 5925 6787 6011 7023
rect 6247 6787 6332 7023
rect 6568 6787 6653 7023
rect 6889 6787 6974 7023
rect 7210 6787 7295 7023
rect 7531 6787 7616 7023
rect 7852 6787 7937 7023
rect 8173 6787 8258 7023
rect 8494 6787 8579 7023
rect 8815 6787 8900 7023
rect 9136 6787 9221 7023
rect 9457 6787 9542 7023
rect 9778 6787 9863 7023
rect 10099 6787 10184 7023
rect 10420 6787 10505 7023
rect 10741 6787 10826 7023
rect 11062 6787 11147 7023
rect 11383 6787 11468 7023
rect 11704 6787 11789 7023
rect 12025 6787 12110 7023
rect 12346 6787 12431 7023
rect 12667 6787 12752 7023
rect 12988 6787 13073 7023
rect 13309 6787 13394 7023
rect 13630 6787 13715 7023
rect 13951 6787 14036 7023
rect 14272 6787 14357 7023
rect 14593 6787 14678 7023
rect 14914 6787 14999 7023
rect 15235 6787 15320 7023
rect 15556 6787 16000 7023
rect 0 6657 16000 6787
rect 0 6421 215 6657
rect 451 6421 537 6657
rect 773 6421 859 6657
rect 1095 6421 1181 6657
rect 1417 6421 1503 6657
rect 1739 6421 1825 6657
rect 2061 6421 2147 6657
rect 2383 6421 2469 6657
rect 2705 6421 2791 6657
rect 3027 6421 3113 6657
rect 3349 6421 3435 6657
rect 3671 6421 3757 6657
rect 3993 6421 4079 6657
rect 4315 6421 4401 6657
rect 4637 6421 4723 6657
rect 4959 6421 5045 6657
rect 5281 6421 5367 6657
rect 5603 6421 5689 6657
rect 5925 6421 6011 6657
rect 6247 6421 6332 6657
rect 6568 6421 6653 6657
rect 6889 6421 6974 6657
rect 7210 6421 7295 6657
rect 7531 6421 7616 6657
rect 7852 6421 7937 6657
rect 8173 6421 8258 6657
rect 8494 6421 8579 6657
rect 8815 6421 8900 6657
rect 9136 6421 9221 6657
rect 9457 6421 9542 6657
rect 9778 6421 9863 6657
rect 10099 6421 10184 6657
rect 10420 6421 10505 6657
rect 10741 6421 10826 6657
rect 11062 6421 11147 6657
rect 11383 6421 11468 6657
rect 11704 6421 11789 6657
rect 12025 6421 12110 6657
rect 12346 6421 12431 6657
rect 12667 6421 12752 6657
rect 12988 6421 13073 6657
rect 13309 6421 13394 6657
rect 13630 6421 13715 6657
rect 13951 6421 14036 6657
rect 14272 6421 14357 6657
rect 14593 6421 14678 6657
rect 14914 6421 14999 6657
rect 15235 6421 15320 6657
rect 15556 6421 16000 6657
rect 0 6397 16000 6421
rect 0 6053 16000 6077
rect 0 5817 215 6053
rect 451 5817 537 6053
rect 773 5817 859 6053
rect 1095 5817 1181 6053
rect 1417 5817 1503 6053
rect 1739 5817 1825 6053
rect 2061 5817 2147 6053
rect 2383 5817 2469 6053
rect 2705 5817 2791 6053
rect 3027 5817 3113 6053
rect 3349 5817 3435 6053
rect 3671 5817 3757 6053
rect 3993 5817 4079 6053
rect 4315 5817 4401 6053
rect 4637 5817 4723 6053
rect 4959 5817 5045 6053
rect 5281 5817 5367 6053
rect 5603 5817 5689 6053
rect 5925 5817 6011 6053
rect 6247 5817 6332 6053
rect 6568 5817 6653 6053
rect 6889 5817 6974 6053
rect 7210 5817 7295 6053
rect 7531 5817 7616 6053
rect 7852 5817 7937 6053
rect 8173 5817 8258 6053
rect 8494 5817 8579 6053
rect 8815 5817 8900 6053
rect 9136 5817 9221 6053
rect 9457 5817 9542 6053
rect 9778 5817 9863 6053
rect 10099 5817 10184 6053
rect 10420 5817 10505 6053
rect 10741 5817 10826 6053
rect 11062 5817 11147 6053
rect 11383 5817 11468 6053
rect 11704 5817 11789 6053
rect 12025 5817 12110 6053
rect 12346 5817 12431 6053
rect 12667 5817 12752 6053
rect 12988 5817 13073 6053
rect 13309 5817 13394 6053
rect 13630 5817 13715 6053
rect 13951 5817 14036 6053
rect 14272 5817 14357 6053
rect 14593 5817 14678 6053
rect 14914 5817 14999 6053
rect 15235 5817 15320 6053
rect 15556 5817 16000 6053
rect 0 5447 16000 5817
rect 0 5211 215 5447
rect 451 5211 537 5447
rect 773 5211 859 5447
rect 1095 5211 1181 5447
rect 1417 5211 1503 5447
rect 1739 5211 1825 5447
rect 2061 5211 2147 5447
rect 2383 5211 2469 5447
rect 2705 5211 2791 5447
rect 3027 5211 3113 5447
rect 3349 5211 3435 5447
rect 3671 5211 3757 5447
rect 3993 5211 4079 5447
rect 4315 5211 4401 5447
rect 4637 5211 4723 5447
rect 4959 5211 5045 5447
rect 5281 5211 5367 5447
rect 5603 5211 5689 5447
rect 5925 5211 6011 5447
rect 6247 5211 6332 5447
rect 6568 5211 6653 5447
rect 6889 5211 6974 5447
rect 7210 5211 7295 5447
rect 7531 5211 7616 5447
rect 7852 5211 7937 5447
rect 8173 5211 8258 5447
rect 8494 5211 8579 5447
rect 8815 5211 8900 5447
rect 9136 5211 9221 5447
rect 9457 5211 9542 5447
rect 9778 5211 9863 5447
rect 10099 5211 10184 5447
rect 10420 5211 10505 5447
rect 10741 5211 10826 5447
rect 11062 5211 11147 5447
rect 11383 5211 11468 5447
rect 11704 5211 11789 5447
rect 12025 5211 12110 5447
rect 12346 5211 12431 5447
rect 12667 5211 12752 5447
rect 12988 5211 13073 5447
rect 13309 5211 13394 5447
rect 13630 5211 13715 5447
rect 13951 5211 14036 5447
rect 14272 5211 14357 5447
rect 14593 5211 14678 5447
rect 14914 5211 14999 5447
rect 15235 5211 15320 5447
rect 15556 5211 16000 5447
rect 0 5187 16000 5211
rect 0 4843 16000 4867
rect 0 4607 215 4843
rect 451 4607 537 4843
rect 773 4607 859 4843
rect 1095 4607 1181 4843
rect 1417 4607 1503 4843
rect 1739 4607 1825 4843
rect 2061 4607 2147 4843
rect 2383 4607 2469 4843
rect 2705 4607 2791 4843
rect 3027 4607 3113 4843
rect 3349 4607 3435 4843
rect 3671 4607 3757 4843
rect 3993 4607 4079 4843
rect 4315 4607 4401 4843
rect 4637 4607 4723 4843
rect 4959 4607 5045 4843
rect 5281 4607 5367 4843
rect 5603 4607 5689 4843
rect 5925 4607 6011 4843
rect 6247 4607 6332 4843
rect 6568 4607 6653 4843
rect 6889 4607 6974 4843
rect 7210 4607 7295 4843
rect 7531 4607 7616 4843
rect 7852 4607 7937 4843
rect 8173 4607 8258 4843
rect 8494 4607 8579 4843
rect 8815 4607 8900 4843
rect 9136 4607 9221 4843
rect 9457 4607 9542 4843
rect 9778 4607 9863 4843
rect 10099 4607 10184 4843
rect 10420 4607 10505 4843
rect 10741 4607 10826 4843
rect 11062 4607 11147 4843
rect 11383 4607 11468 4843
rect 11704 4607 11789 4843
rect 12025 4607 12110 4843
rect 12346 4607 12431 4843
rect 12667 4607 12752 4843
rect 12988 4607 13073 4843
rect 13309 4607 13394 4843
rect 13630 4607 13715 4843
rect 13951 4607 14036 4843
rect 14272 4607 14357 4843
rect 14593 4607 14678 4843
rect 14914 4607 14999 4843
rect 15235 4607 15320 4843
rect 15556 4607 16000 4843
rect 0 4237 16000 4607
rect 0 4001 215 4237
rect 451 4001 537 4237
rect 773 4001 859 4237
rect 1095 4001 1181 4237
rect 1417 4001 1503 4237
rect 1739 4001 1825 4237
rect 2061 4001 2147 4237
rect 2383 4001 2469 4237
rect 2705 4001 2791 4237
rect 3027 4001 3113 4237
rect 3349 4001 3435 4237
rect 3671 4001 3757 4237
rect 3993 4001 4079 4237
rect 4315 4001 4401 4237
rect 4637 4001 4723 4237
rect 4959 4001 5045 4237
rect 5281 4001 5367 4237
rect 5603 4001 5689 4237
rect 5925 4001 6011 4237
rect 6247 4001 6332 4237
rect 6568 4001 6653 4237
rect 6889 4001 6974 4237
rect 7210 4001 7295 4237
rect 7531 4001 7616 4237
rect 7852 4001 7937 4237
rect 8173 4001 8258 4237
rect 8494 4001 8579 4237
rect 8815 4001 8900 4237
rect 9136 4001 9221 4237
rect 9457 4001 9542 4237
rect 9778 4001 9863 4237
rect 10099 4001 10184 4237
rect 10420 4001 10505 4237
rect 10741 4001 10826 4237
rect 11062 4001 11147 4237
rect 11383 4001 11468 4237
rect 11704 4001 11789 4237
rect 12025 4001 12110 4237
rect 12346 4001 12431 4237
rect 12667 4001 12752 4237
rect 12988 4001 13073 4237
rect 13309 4001 13394 4237
rect 13630 4001 13715 4237
rect 13951 4001 14036 4237
rect 14272 4001 14357 4237
rect 14593 4001 14678 4237
rect 14914 4001 14999 4237
rect 15235 4001 15320 4237
rect 15556 4001 16000 4237
rect 0 3977 16000 4001
rect 0 3633 16000 3657
rect 0 3397 215 3633
rect 451 3397 537 3633
rect 773 3397 859 3633
rect 1095 3397 1181 3633
rect 1417 3397 1503 3633
rect 1739 3397 1825 3633
rect 2061 3397 2147 3633
rect 2383 3397 2469 3633
rect 2705 3397 2791 3633
rect 3027 3397 3113 3633
rect 3349 3397 3435 3633
rect 3671 3397 3757 3633
rect 3993 3397 4079 3633
rect 4315 3397 4401 3633
rect 4637 3397 4723 3633
rect 4959 3397 5045 3633
rect 5281 3397 5367 3633
rect 5603 3397 5689 3633
rect 5925 3397 6011 3633
rect 6247 3397 6332 3633
rect 6568 3397 6653 3633
rect 6889 3397 6974 3633
rect 7210 3397 7295 3633
rect 7531 3397 7616 3633
rect 7852 3397 7937 3633
rect 8173 3397 8258 3633
rect 8494 3397 8579 3633
rect 8815 3397 8900 3633
rect 9136 3397 9221 3633
rect 9457 3397 9542 3633
rect 9778 3397 9863 3633
rect 10099 3397 10184 3633
rect 10420 3397 10505 3633
rect 10741 3397 10826 3633
rect 11062 3397 11147 3633
rect 11383 3397 11468 3633
rect 11704 3397 11789 3633
rect 12025 3397 12110 3633
rect 12346 3397 12431 3633
rect 12667 3397 12752 3633
rect 12988 3397 13073 3633
rect 13309 3397 13394 3633
rect 13630 3397 13715 3633
rect 13951 3397 14036 3633
rect 14272 3397 14357 3633
rect 14593 3397 14678 3633
rect 14914 3397 14999 3633
rect 15235 3397 15320 3633
rect 15556 3397 16000 3633
rect 0 3267 16000 3397
rect 0 3031 215 3267
rect 451 3031 537 3267
rect 773 3031 859 3267
rect 1095 3031 1181 3267
rect 1417 3031 1503 3267
rect 1739 3031 1825 3267
rect 2061 3031 2147 3267
rect 2383 3031 2469 3267
rect 2705 3031 2791 3267
rect 3027 3031 3113 3267
rect 3349 3031 3435 3267
rect 3671 3031 3757 3267
rect 3993 3031 4079 3267
rect 4315 3031 4401 3267
rect 4637 3031 4723 3267
rect 4959 3031 5045 3267
rect 5281 3031 5367 3267
rect 5603 3031 5689 3267
rect 5925 3031 6011 3267
rect 6247 3031 6332 3267
rect 6568 3031 6653 3267
rect 6889 3031 6974 3267
rect 7210 3031 7295 3267
rect 7531 3031 7616 3267
rect 7852 3031 7937 3267
rect 8173 3031 8258 3267
rect 8494 3031 8579 3267
rect 8815 3031 8900 3267
rect 9136 3031 9221 3267
rect 9457 3031 9542 3267
rect 9778 3031 9863 3267
rect 10099 3031 10184 3267
rect 10420 3031 10505 3267
rect 10741 3031 10826 3267
rect 11062 3031 11147 3267
rect 11383 3031 11468 3267
rect 11704 3031 11789 3267
rect 12025 3031 12110 3267
rect 12346 3031 12431 3267
rect 12667 3031 12752 3267
rect 12988 3031 13073 3267
rect 13309 3031 13394 3267
rect 13630 3031 13715 3267
rect 13951 3031 14036 3267
rect 14272 3031 14357 3267
rect 14593 3031 14678 3267
rect 14914 3031 14999 3267
rect 15235 3031 15320 3267
rect 15556 3031 16000 3267
rect 0 3007 16000 3031
rect 0 2663 16000 2687
rect 0 2427 215 2663
rect 451 2427 537 2663
rect 773 2427 859 2663
rect 1095 2427 1181 2663
rect 1417 2427 1503 2663
rect 1739 2427 1825 2663
rect 2061 2427 2147 2663
rect 2383 2427 2469 2663
rect 2705 2427 2791 2663
rect 3027 2427 3113 2663
rect 3349 2427 3435 2663
rect 3671 2427 3757 2663
rect 3993 2427 4079 2663
rect 4315 2427 4401 2663
rect 4637 2427 4723 2663
rect 4959 2427 5045 2663
rect 5281 2427 5367 2663
rect 5603 2427 5689 2663
rect 5925 2427 6011 2663
rect 6247 2427 6332 2663
rect 6568 2427 6653 2663
rect 6889 2427 6974 2663
rect 7210 2427 7295 2663
rect 7531 2427 7616 2663
rect 7852 2427 7937 2663
rect 8173 2427 8258 2663
rect 8494 2427 8579 2663
rect 8815 2427 8900 2663
rect 9136 2427 9221 2663
rect 9457 2427 9542 2663
rect 9778 2427 9863 2663
rect 10099 2427 10184 2663
rect 10420 2427 10505 2663
rect 10741 2427 10826 2663
rect 11062 2427 11147 2663
rect 11383 2427 11468 2663
rect 11704 2427 11789 2663
rect 12025 2427 12110 2663
rect 12346 2427 12431 2663
rect 12667 2427 12752 2663
rect 12988 2427 13073 2663
rect 13309 2427 13394 2663
rect 13630 2427 13715 2663
rect 13951 2427 14036 2663
rect 14272 2427 14357 2663
rect 14593 2427 14678 2663
rect 14914 2427 14999 2663
rect 15235 2427 15320 2663
rect 15556 2427 16000 2663
rect 0 2057 16000 2427
rect 0 1821 215 2057
rect 451 1821 537 2057
rect 773 1821 859 2057
rect 1095 1821 1181 2057
rect 1417 1821 1503 2057
rect 1739 1821 1825 2057
rect 2061 1821 2147 2057
rect 2383 1821 2469 2057
rect 2705 1821 2791 2057
rect 3027 1821 3113 2057
rect 3349 1821 3435 2057
rect 3671 1821 3757 2057
rect 3993 1821 4079 2057
rect 4315 1821 4401 2057
rect 4637 1821 4723 2057
rect 4959 1821 5045 2057
rect 5281 1821 5367 2057
rect 5603 1821 5689 2057
rect 5925 1821 6011 2057
rect 6247 1821 6332 2057
rect 6568 1821 6653 2057
rect 6889 1821 6974 2057
rect 7210 1821 7295 2057
rect 7531 1821 7616 2057
rect 7852 1821 7937 2057
rect 8173 1821 8258 2057
rect 8494 1821 8579 2057
rect 8815 1821 8900 2057
rect 9136 1821 9221 2057
rect 9457 1821 9542 2057
rect 9778 1821 9863 2057
rect 10099 1821 10184 2057
rect 10420 1821 10505 2057
rect 10741 1821 10826 2057
rect 11062 1821 11147 2057
rect 11383 1821 11468 2057
rect 11704 1821 11789 2057
rect 12025 1821 12110 2057
rect 12346 1821 12431 2057
rect 12667 1821 12752 2057
rect 12988 1821 13073 2057
rect 13309 1821 13394 2057
rect 13630 1821 13715 2057
rect 13951 1821 14036 2057
rect 14272 1821 14357 2057
rect 14593 1821 14678 2057
rect 14914 1821 14999 2057
rect 15235 1821 15320 2057
rect 15556 1821 16000 2057
rect 0 1797 16000 1821
rect 0 1452 16000 1477
rect 0 1216 215 1452
rect 451 1216 537 1452
rect 773 1216 859 1452
rect 1095 1216 1181 1452
rect 1417 1216 1503 1452
rect 1739 1216 1825 1452
rect 2061 1216 2147 1452
rect 2383 1216 2469 1452
rect 2705 1216 2791 1452
rect 3027 1216 3113 1452
rect 3349 1216 3435 1452
rect 3671 1216 3757 1452
rect 3993 1216 4079 1452
rect 4315 1216 4401 1452
rect 4637 1216 4723 1452
rect 4959 1216 5045 1452
rect 5281 1216 5367 1452
rect 5603 1216 5689 1452
rect 5925 1216 6011 1452
rect 6247 1216 6332 1452
rect 6568 1216 6653 1452
rect 6889 1216 6974 1452
rect 7210 1216 7295 1452
rect 7531 1216 7616 1452
rect 7852 1216 7937 1452
rect 8173 1216 8258 1452
rect 8494 1216 8579 1452
rect 8815 1216 8900 1452
rect 9136 1216 9221 1452
rect 9457 1216 9542 1452
rect 9778 1216 9863 1452
rect 10099 1216 10184 1452
rect 10420 1216 10505 1452
rect 10741 1216 10826 1452
rect 11062 1216 11147 1452
rect 11383 1216 11468 1452
rect 11704 1216 11789 1452
rect 12025 1216 12110 1452
rect 12346 1216 12431 1452
rect 12667 1216 12752 1452
rect 12988 1216 13073 1452
rect 13309 1216 13394 1452
rect 13630 1216 13715 1452
rect 13951 1216 14036 1452
rect 14272 1216 14357 1452
rect 14593 1216 14678 1452
rect 14914 1216 14999 1452
rect 15235 1216 15320 1452
rect 15556 1216 16000 1452
rect 0 1070 16000 1216
rect 0 834 215 1070
rect 451 834 537 1070
rect 773 834 859 1070
rect 1095 834 1181 1070
rect 1417 834 1503 1070
rect 1739 834 1825 1070
rect 2061 834 2147 1070
rect 2383 834 2469 1070
rect 2705 834 2791 1070
rect 3027 834 3113 1070
rect 3349 834 3435 1070
rect 3671 834 3757 1070
rect 3993 834 4079 1070
rect 4315 834 4401 1070
rect 4637 834 4723 1070
rect 4959 834 5045 1070
rect 5281 834 5367 1070
rect 5603 834 5689 1070
rect 5925 834 6011 1070
rect 6247 834 6332 1070
rect 6568 834 6653 1070
rect 6889 834 6974 1070
rect 7210 834 7295 1070
rect 7531 834 7616 1070
rect 7852 834 7937 1070
rect 8173 834 8258 1070
rect 8494 834 8579 1070
rect 8815 834 8900 1070
rect 9136 834 9221 1070
rect 9457 834 9542 1070
rect 9778 834 9863 1070
rect 10099 834 10184 1070
rect 10420 834 10505 1070
rect 10741 834 10826 1070
rect 11062 834 11147 1070
rect 11383 834 11468 1070
rect 11704 834 11789 1070
rect 12025 834 12110 1070
rect 12346 834 12431 1070
rect 12667 834 12752 1070
rect 12988 834 13073 1070
rect 13309 834 13394 1070
rect 13630 834 13715 1070
rect 13951 834 14036 1070
rect 14272 834 14357 1070
rect 14593 834 14678 1070
rect 14914 834 14999 1070
rect 15235 834 15320 1070
rect 15556 834 16000 1070
rect 0 688 16000 834
rect 0 452 215 688
rect 451 452 537 688
rect 773 452 859 688
rect 1095 452 1181 688
rect 1417 452 1503 688
rect 1739 452 1825 688
rect 2061 452 2147 688
rect 2383 452 2469 688
rect 2705 452 2791 688
rect 3027 452 3113 688
rect 3349 452 3435 688
rect 3671 452 3757 688
rect 3993 452 4079 688
rect 4315 452 4401 688
rect 4637 452 4723 688
rect 4959 452 5045 688
rect 5281 452 5367 688
rect 5603 452 5689 688
rect 5925 452 6011 688
rect 6247 452 6332 688
rect 6568 452 6653 688
rect 6889 452 6974 688
rect 7210 452 7295 688
rect 7531 452 7616 688
rect 7852 452 7937 688
rect 8173 452 8258 688
rect 8494 452 8579 688
rect 8815 452 8900 688
rect 9136 452 9221 688
rect 9457 452 9542 688
rect 9778 452 9863 688
rect 10099 452 10184 688
rect 10420 452 10505 688
rect 10741 452 10826 688
rect 11062 452 11147 688
rect 11383 452 11468 688
rect 11704 452 11789 688
rect 12025 452 12110 688
rect 12346 452 12431 688
rect 12667 452 12752 688
rect 12988 452 13073 688
rect 13309 452 13394 688
rect 13630 452 13715 688
rect 13951 452 14036 688
rect 14272 452 14357 688
rect 14593 452 14678 688
rect 14914 452 14999 688
rect 15235 452 15320 688
rect 15556 452 16000 688
rect 0 427 16000 452
use nfet_CDNS_52468879185592  nfet_CDNS_52468879185592_0
timestamp 1707688321
transform 0 1 7315 1 0 487
box -79 -32 335 632
use sky130_fd_io__gpiovrefv2_ctl  sky130_fd_io__gpiovrefv2_ctl_0
timestamp 1707688321
transform 1 0 1420 0 1 5
box -92 0 10574 4277
use sky130_fd_io__gpiovrefv2_decoder_5_32  sky130_fd_io__gpiovrefv2_decoder_5_32_0
timestamp 1707688321
transform 0 -1 9525 1 0 1278
box 0 -160 38722 2696
use sky130_fd_io__gpiovrefv2_res_ladder  sky130_fd_io__gpiovrefv2_res_ladder_0
timestamp 1707688321
transform 1 0 643 0 1 1203
box -278 -967 15000 38783
<< labels >>
flabel comment s 13403 25375 13403 25375 0 FreeSans 10000 90 0 0 M3 shield
flabel comment s 10595 25375 10595 25375 0 FreeSans 10000 90 0 0 M3 shield
flabel comment s 5764 25375 5764 25375 0 FreeSans 10000 90 0 0 M3 shield
flabel comment s 3457 25375 3457 25375 0 FreeSans 10000 90 0 0 M3 shield
flabel comment s 1428 25375 1428 25375 0 FreeSans 10000 90 0 0 M3 shield
flabel metal1 s 7497 0 7625 128 3 FreeSans 200 0 0 0 vinref
port 10 nsew signal bidirectional
flabel metal1 s 1231 0 1283 128 3 FreeSans 200 0 0 0 ref_sel<4>
port 2 nsew signal input
flabel metal1 s 979 0 1031 128 3 FreeSans 200 0 0 0 ref_sel<3>
port 3 nsew signal input
flabel metal1 s 13080 0 13132 128 3 FreeSans 200 0 0 0 ref_sel<1>
port 4 nsew signal input
flabel metal1 s 6059 0 6111 128 3 FreeSans 200 0 0 0 vrefgen_en
port 5 nsew signal input
flabel metal1 s 6347 0 6399 128 3 FreeSans 200 0 0 0 hld_h_n
port 6 nsew signal input
flabel metal1 s 6547 0 6599 128 3 FreeSans 200 0 0 0 enable_h
port 7 nsew signal input
flabel metal1 s 6745 0 6797 128 3 FreeSans 200 0 0 0 ref_sel<2>
port 8 nsew signal input
flabel metal1 s 12099 0 12151 128 3 FreeSans 200 0 0 0 ref_sel<0>
port 9 nsew signal input
flabel metal5 s 0 12837 254 13687 3 FreeSans 520 0 0 0 vddio_q
port 11 nsew power bidirectional
flabel metal5 s 0 14007 254 18997 3 FreeSans 520 0 0 0 vddio
port 12 nsew power bidirectional
flabel metal5 s 0 35157 254 40000 3 FreeSans 520 0 0 0 vssio
port 13 nsew ground bidirectional
flabel metal5 s 0 9547 254 11347 3 FreeSans 520 0 0 0 vssa
port 14 nsew ground bidirectional
flabel metal5 s 0 1797 254 2687 3 FreeSans 520 0 0 0 vccd
port 15 nsew power bidirectional
flabel metal5 s 0 7367 254 8017 3 FreeSans 520 0 0 0 vssa
port 14 nsew ground bidirectional
flabel metal5 s 0 3977 254 4867 3 FreeSans 520 0 0 0 vddio
port 12 nsew power bidirectional
flabel metal5 s 0 427 254 1477 3 FreeSans 520 0 0 0 vcchib
port 16 nsew power bidirectional
flabel metal5 s 0 6397 254 7047 3 FreeSans 520 0 0 0 vswitch
port 17 nsew power bidirectional
flabel metal5 s 0 5187 254 6077 3 FreeSans 520 0 0 0 vssio
port 13 nsew ground bidirectional
flabel metal5 s 0 11667 254 12517 3 FreeSans 520 0 0 0 vssio_q
port 18 nsew ground bidirectional
flabel metal5 s 0 3007 193 3657 3 FreeSans 520 0 0 0 vdda
port 19 nsew power bidirectional
flabel metal5 s 0 8337 254 9227 3 FreeSans 520 0 0 0 vssd
port 20 nsew ground bidirectional
flabel metal5 s 15746 9547 16000 11347 3 FreeSans 520 180 0 0 vssa
port 14 nsew ground bidirectional
flabel metal5 s 15746 8337 16000 9227 3 FreeSans 520 180 0 0 vssd
port 20 nsew ground bidirectional
flabel metal5 s 15807 3007 16000 3657 3 FreeSans 520 180 0 0 vdda
port 19 nsew power bidirectional
flabel metal5 s 15746 5187 16000 6077 3 FreeSans 520 180 0 0 vssio
port 13 nsew ground bidirectional
flabel metal5 s 15746 6397 16000 7047 3 FreeSans 520 180 0 0 vswitch
port 17 nsew power bidirectional
flabel metal5 s 15746 427 16000 1477 3 FreeSans 520 180 0 0 vcchib
port 16 nsew power bidirectional
flabel metal5 s 15746 3977 16000 4867 3 FreeSans 520 180 0 0 vddio
port 12 nsew power bidirectional
flabel metal5 s 15746 7367 16000 8017 3 FreeSans 520 180 0 0 vssa
port 14 nsew ground bidirectional
flabel metal5 s 15746 1797 16000 2687 3 FreeSans 520 180 0 0 vccd
port 15 nsew power bidirectional
flabel metal5 s 15746 11667 16000 12517 3 FreeSans 520 180 0 0 vssio_q
port 18 nsew ground bidirectional
flabel metal5 s 15746 14007 16000 18997 3 FreeSans 520 180 0 0 vddio
port 12 nsew power bidirectional
flabel metal5 s 15746 12837 16000 13687 3 FreeSans 520 180 0 0 vddio_q
port 11 nsew power bidirectional
flabel metal5 s 15746 35157 16000 40000 3 FreeSans 520 180 0 0 vssio
port 13 nsew ground bidirectional
flabel metal4 s 0 12817 254 13707 3 FreeSans 520 0 0 0 vddio_q
port 11 nsew power bidirectional
flabel metal4 s 0 14007 254 19000 3 FreeSans 520 0 0 0 vddio
port 12 nsew power bidirectional
flabel metal4 s 0 35157 254 39999 3 FreeSans 520 0 0 0 vssio
port 13 nsew ground bidirectional
flabel metal4 s 0 9673 254 10269 3 FreeSans 520 0 0 0 amuxbus_b
port 21 nsew signal bidirectional
flabel metal4 s 0 1777 254 2707 3 FreeSans 520 0 0 0 vccd
port 15 nsew power bidirectional
flabel metal4 s 0 7347 254 8037 3 FreeSans 520 0 0 0 vssa
port 14 nsew ground bidirectional
flabel metal4 s 0 3957 254 4887 3 FreeSans 520 0 0 0 vddio
port 12 nsew power bidirectional
flabel metal4 s 0 407 254 1497 3 FreeSans 520 0 0 0 vcchib
port 16 nsew power bidirectional
flabel metal4 s 0 6377 254 7067 3 FreeSans 520 0 0 0 vswitch
port 17 nsew power bidirectional
flabel metal4 s 0 5167 254 6097 3 FreeSans 520 0 0 0 vssio
port 13 nsew ground bidirectional
flabel metal4 s 0 11647 254 12537 3 FreeSans 520 0 0 0 vssio_q
port 18 nsew ground bidirectional
flabel metal4 s 0 2987 193 3677 3 FreeSans 520 0 0 0 vdda
port 19 nsew power bidirectional
flabel metal4 s 0 8317 254 9247 3 FreeSans 520 0 0 0 vssd
port 20 nsew ground bidirectional
flabel metal4 s 0 10625 254 11221 3 FreeSans 520 0 0 0 amuxbus_a
port 22 nsew signal bidirectional
flabel metal4 s 0 11281 254 11347 3 FreeSans 520 0 0 0 vssa
port 14 nsew ground bidirectional
flabel metal4 s 0 10329 254 10565 3 FreeSans 520 0 0 0 vssa
port 14 nsew ground bidirectional
flabel metal4 s 0 9547 254 9613 3 FreeSans 520 0 0 0 vssa
port 14 nsew ground bidirectional
flabel metal4 s 15746 11281 16000 11347 3 FreeSans 520 180 0 0 vssa
port 14 nsew ground bidirectional
flabel metal4 s 15746 10329 16000 10565 3 FreeSans 520 180 0 0 vssa
port 14 nsew ground bidirectional
flabel metal4 s 15746 9547 16000 9613 3 FreeSans 520 180 0 0 vssa
port 14 nsew ground bidirectional
flabel metal4 s 15746 10625 16000 11221 3 FreeSans 520 180 0 0 amuxbus_a
port 22 nsew signal bidirectional
flabel metal4 s 15746 8317 16000 9247 3 FreeSans 520 180 0 0 vssd
port 20 nsew ground bidirectional
flabel metal4 s 15807 2987 16000 3677 3 FreeSans 520 180 0 0 vdda
port 19 nsew power bidirectional
flabel metal4 s 15746 11647 16000 12537 3 FreeSans 520 180 0 0 vssio_q
port 18 nsew ground bidirectional
flabel metal4 s 15746 5167 16000 6097 3 FreeSans 520 180 0 0 vssio
port 13 nsew ground bidirectional
flabel metal4 s 15746 6377 16000 7067 3 FreeSans 520 180 0 0 vswitch
port 17 nsew power bidirectional
flabel metal4 s 15746 407 16000 1497 3 FreeSans 520 180 0 0 vcchib
port 16 nsew power bidirectional
flabel metal4 s 15746 3957 16000 4887 3 FreeSans 520 180 0 0 vddio
port 12 nsew power bidirectional
flabel metal4 s 15746 7347 16000 8037 3 FreeSans 520 180 0 0 vssa
port 14 nsew ground bidirectional
flabel metal4 s 15746 12817 16000 13707 3 FreeSans 520 180 0 0 vddio_q
port 11 nsew power bidirectional
flabel metal4 s 15746 1777 16000 2707 3 FreeSans 520 180 0 0 vccd
port 15 nsew power bidirectional
flabel metal4 s 15746 9673 16000 10269 3 FreeSans 520 180 0 0 amuxbus_b
port 21 nsew signal bidirectional
flabel metal4 s 15746 35157 16000 39999 3 FreeSans 520 180 0 0 vssio
port 13 nsew ground bidirectional
flabel metal4 s 15746 14007 16000 19000 3 FreeSans 520 180 0 0 vddio
port 12 nsew power bidirectional
flabel metal2 s 6745 0 6797 128 3 FreeSans 200 0 0 0 ref_sel<2>
port 8 nsew signal input
flabel metal2 s 6547 0 6599 128 3 FreeSans 200 0 0 0 enable_h
port 7 nsew signal input
flabel metal2 s 6059 0 6111 128 3 FreeSans 200 0 0 0 vrefgen_en
port 5 nsew signal input
flabel metal2 s 6347 0 6399 128 3 FreeSans 200 0 0 0 hld_h_n
port 6 nsew signal input
flabel metal2 s 12099 0 12151 128 3 FreeSans 200 0 0 0 ref_sel<0>
port 9 nsew signal input
flabel metal2 s 7497 0 7625 128 3 FreeSans 200 0 0 0 vinref
port 10 nsew signal bidirectional
flabel metal2 s 1231 0 1283 128 3 FreeSans 200 0 0 0 ref_sel<4>
port 2 nsew signal input
flabel metal2 s 979 0 1031 128 3 FreeSans 200 0 0 0 ref_sel<3>
port 3 nsew signal input
flabel metal2 s 13080 0 13132 128 3 FreeSans 200 0 0 0 ref_sel<1>
port 4 nsew signal input
rlabel metal1 s 6745 0 6797 3007 1 ref_sel<2>
port 8 nsew signal input
rlabel metal1 s 6547 0 6599 465 1 enable_h
port 7 nsew signal input
rlabel metal1 s 5983 547 6111 599 1 vrefgen_en
port 5 nsew signal input
rlabel metal1 s 6031 541 6111 547 1 vrefgen_en
port 5 nsew signal input
rlabel metal1 s 6045 527 6111 541 1 vrefgen_en
port 5 nsew signal input
rlabel metal1 s 6059 513 6111 527 1 vrefgen_en
port 5 nsew signal input
rlabel metal1 s 6059 0 6111 513 1 vrefgen_en
port 5 nsew signal input
rlabel metal1 s 6347 0 6399 465 1 hld_h_n
port 6 nsew signal input
rlabel metal1 s 11899 710 12080 720 1 ref_sel<0>
port 9 nsew signal input
rlabel metal1 s 11899 696 12090 710 1 ref_sel<0>
port 9 nsew signal input
rlabel metal1 s 11899 682 12104 696 1 ref_sel<0>
port 9 nsew signal input
rlabel metal1 s 11899 668 12118 682 1 ref_sel<0>
port 9 nsew signal input
rlabel metal1 s 12059 667 12132 668 1 ref_sel<0>
port 9 nsew signal input
rlabel metal1 s 12068 658 12133 667 1 ref_sel<0>
port 9 nsew signal input
rlabel metal1 s 12077 649 12142 658 1 ref_sel<0>
port 9 nsew signal input
rlabel metal1 s 12088 638 12151 649 1 ref_sel<0>
port 9 nsew signal input
rlabel metal1 s 12099 627 12151 638 1 ref_sel<0>
port 9 nsew signal input
rlabel metal1 s 12099 0 12151 627 1 ref_sel<0>
port 9 nsew signal input
rlabel metal1 s 7497 0 7625 128 1 vinref
port 10 nsew signal bidirectional
rlabel metal1 s 1231 0 1283 128 1 ref_sel<4>
port 2 nsew signal input
rlabel metal1 s 979 0 1031 128 1 ref_sel<3>
port 3 nsew signal input
rlabel metal1 s 13080 0 13132 128 1 ref_sel<1>
port 4 nsew signal input
rlabel metal4 s 0 8317 16000 9247 1 vssd
port 20 nsew ground bidirectional
rlabel metal4 s 0 2987 16000 3677 1 vdda
port 19 nsew power bidirectional
rlabel metal4 s 0 6377 16000 7067 1 vswitch
port 17 nsew power bidirectional
rlabel metal4 s 0 407 16000 1497 1 vcchib
port 16 nsew power bidirectional
rlabel metal5 s 0 9547 16000 11347 1 vssa
port 14 nsew ground bidirectional
rlabel metal4 s 0 7347 16000 8037 1 vssa
port 14 nsew ground bidirectional
rlabel metal4 s 0 9547 16000 9613 1 vssa
port 14 nsew ground bidirectional
rlabel metal4 s 0 10329 16000 10565 1 vssa
port 14 nsew ground bidirectional
rlabel metal4 s 0 11281 16000 11347 1 vssa
port 14 nsew ground bidirectional
rlabel metal4 s 0 1777 16000 2707 1 vccd
port 15 nsew power bidirectional
rlabel metal4 s 0 11647 16000 12537 1 vssio_q
port 18 nsew ground bidirectional
rlabel metal5 s 0 14007 16000 18997 1 vddio
port 12 nsew power bidirectional
rlabel metal4 s 0 3957 16000 4887 1 vddio
port 12 nsew power bidirectional
rlabel metal4 s 0 14007 16000 19000 1 vddio
port 12 nsew power bidirectional
rlabel metal4 s 0 12817 16000 13707 1 vddio_q
port 11 nsew power bidirectional
rlabel metal5 s 0 35157 16000 40000 1 vssio
port 13 nsew ground bidirectional
rlabel metal4 s 0 5167 16000 6097 1 vssio
port 13 nsew ground bidirectional
rlabel metal4 s 0 35157 16000 40000 1 vssio
port 13 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 16000 40000
string GDS_END 26381912
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 25924122
string LEFclass BLOCK
string LEFsymmetry R90
string path 200.325 207.925 200.325 231.175 
<< end >>
