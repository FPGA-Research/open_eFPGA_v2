magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< poly >>
rect 973 819 1091 836
rect 3131 819 3249 836
rect 973 803 1107 819
rect 973 769 989 803
rect 1023 769 1057 803
rect 1091 769 1107 803
rect 973 753 1107 769
rect 3115 803 3249 819
rect 3115 769 3131 803
rect 3165 769 3199 803
rect 3233 769 3249 803
rect 3115 753 3249 769
rect 973 736 1091 753
rect 3131 736 3249 753
<< polycont >>
rect 989 769 1023 803
rect 1057 769 1091 803
rect 3131 769 3165 803
rect 3199 769 3233 803
<< locali >>
rect 989 804 1091 819
rect 3131 804 3233 819
rect 1021 803 1059 804
rect 1023 769 1057 803
rect 3163 803 3201 804
rect 989 753 1091 769
rect 3165 769 3199 803
rect 3131 753 3233 769
<< viali >>
rect 987 803 1021 804
rect 1059 803 1093 804
rect 987 770 989 803
rect 989 770 1021 803
rect 1059 770 1091 803
rect 1091 770 1093 803
rect 3129 803 3163 804
rect 3201 803 3235 804
rect 3129 770 3131 803
rect 3131 770 3163 803
rect 3201 770 3233 803
rect 3233 770 3235 803
<< metal1 >>
tri -3732 12180 -3731 12181 se
tri -1939 12180 -1938 12181 sw
rect -4565 11680 -3518 11705
rect -4565 1127 -3700 11680
tri -3700 11498 -3518 11680 nw
rect -4565 1088 -3739 1127
tri -3739 1088 -3700 1127 nw
rect -4471 1054 -4345 1088
tri -4345 1054 -4311 1088 nw
rect -4471 1033 -4366 1054
tri -4366 1033 -4345 1054 nw
tri -2570 1033 -2549 1054 se
tri -2419 1033 -2398 1054 sw
tri -2058 1033 -2037 1054 se
tri -1907 1033 -1886 1054 sw
tri -766 1033 -745 1054 se
tri -615 1033 -594 1054 sw
tri -254 1033 -233 1054 se
tri -103 1033 -82 1054 sw
tri 1038 1033 1059 1054 se
tri 1189 1033 1210 1054 sw
tri 1550 1033 1571 1054 se
tri 1701 1033 1722 1054 sw
tri 2842 1033 2863 1054 se
tri 2993 1033 3014 1054 sw
tri 3354 1033 3375 1054 se
tri 3505 1033 3526 1054 sw
tri 4646 1033 4667 1054 se
tri 4797 1033 4818 1054 sw
tri 5158 1033 5179 1054 se
rect 5179 1033 5309 1054
tri 5309 1033 5330 1054 sw
tri 6450 1033 6471 1054 se
tri 6601 1033 6622 1054 sw
tri 6962 1033 6983 1054 se
tri 7113 1033 7134 1054 sw
tri 8254 1033 8275 1054 se
tri 8405 1033 8426 1054 sw
tri 8766 1033 8787 1054 se
tri 8917 1033 8938 1054 sw
tri 10209 1033 10230 1054 sw
tri 10570 1033 10591 1054 se
tri 10721 1033 10742 1054 sw
tri 11862 1033 11883 1054 se
tri 12013 1033 12034 1054 sw
tri 12374 1033 12395 1054 se
tri 12525 1033 12546 1054 sw
rect -4471 1032 -4367 1033
tri -4367 1032 -4366 1033 nw
tri -3629 1032 -3628 1033 se
rect -4471 974 -4425 1032
tri -4425 974 -4367 1032 nw
rect -3628 981 8526 1033
rect 8527 982 8528 1032
rect 8564 982 8565 1032
rect 8566 981 8970 1033
rect 9022 981 9038 1033
rect 9090 981 9096 1033
rect 10079 981 10395 1033
rect 10397 1032 10433 1033
rect 10396 982 10434 1032
rect 10397 981 10433 982
rect 10435 981 10746 1033
rect 10798 981 10814 1033
rect 10866 981 11229 1033
rect 11231 1032 11267 1033
rect 11230 982 11268 1032
rect 11231 981 11267 982
rect 11269 981 11715 1033
rect 11767 981 11783 1033
rect 11835 981 12199 1033
rect 12200 982 12201 1032
rect 12237 982 12238 1032
rect 12239 981 13116 1033
rect 13118 1032 13154 1033
rect 13117 982 13155 1032
rect 13118 981 13154 982
rect 13156 981 13687 1033
tri 13687 1032 13688 1033 sw
tri -3628 974 -3621 981 nw
tri 8268 974 8275 981 ne
rect 8275 974 8402 981
tri -4471 928 -4425 974 nw
tri 8275 951 8298 974 ne
rect 981 804 1099 816
rect 981 770 987 804
rect 1021 770 1059 804
rect 1093 770 1099 804
tri 953 620 981 648 se
rect 981 620 1099 770
rect 3119 804 3249 835
tri 8297 818 8298 819 se
rect 8298 818 8402 974
tri 8402 953 8430 981 nw
tri 10051 876 10079 904 se
rect 10079 877 10209 981
tri 10209 948 10242 981 nw
tri 13680 974 13687 981 ne
rect 13768 1000 13867 1032
tri 13867 1000 13899 1032 sw
rect 13768 999 13954 1000
tri 13954 999 13955 1000 sw
rect 13768 974 14018 999
tri 13834 948 13860 974 ne
rect 13860 948 14018 974
tri 13860 947 13861 948 ne
rect 13861 947 14018 948
tri 13435 904 13476 945 se
rect 13476 904 13699 945
tri 10209 877 10236 904 sw
tri 13408 877 13435 904 se
rect 13435 901 13699 904
tri 13699 901 13743 945 sw
rect 13435 889 13743 901
tri 13743 889 13755 901 sw
rect 13435 877 13501 889
tri 13501 877 13513 889 nw
tri 13672 877 13684 889 ne
rect 13684 877 13755 889
rect 10079 876 10236 877
tri 10236 876 10237 877 sw
tri 13390 876 13391 877 se
rect 13391 876 13500 877
tri 13500 876 13501 877 nw
tri 13684 876 13685 877 ne
rect 13685 876 13755 877
tri 13755 876 13768 889 sw
rect 10051 824 13448 876
tri 13448 824 13500 876 nw
tri 13685 824 13737 876 ne
rect 13737 824 13774 876
rect 10051 818 13442 824
tri 13442 818 13448 824 nw
tri 13588 818 13594 824 se
tri 13737 818 13743 824 ne
rect 13743 818 13774 824
tri 8295 816 8297 818 se
rect 8297 816 8402 818
tri 13586 816 13588 818 se
rect 13588 816 13594 818
rect 3119 770 3129 804
rect 3163 770 3201 804
rect 3235 770 3249 804
tri 8269 790 8295 816 se
rect 8295 790 8402 816
tri 13585 815 13586 816 se
rect 13586 815 13594 816
tri 8402 790 8427 815 sw
tri 13560 790 13585 815 se
rect 13585 790 13594 815
rect 3119 705 3249 770
rect 8267 733 13532 790
tri 14279 733 14291 745 se
tri 3249 705 3277 733 sw
tri 14251 705 14279 733 se
rect 14279 705 14291 733
rect 3119 703 13532 705
rect 3119 686 8970 703
tri 3119 648 3157 686 ne
rect 3157 651 8970 686
rect 9022 651 9038 703
rect 9090 651 10746 703
rect 10798 651 10814 703
rect 10866 651 11715 703
rect 11767 651 11783 703
rect 11835 651 13532 703
rect 3157 648 13532 651
tri 1099 620 1127 648 sw
tri 4573 287 4574 288 sw
tri 6378 287 6379 288 sw
tri 1772 283 1776 287 se
tri -40 250 -7 283 se
tri 953 250 986 283 sw
tri 1739 250 1772 283 se
rect 1772 250 1776 283
tri 2768 283 2772 287 sw
rect 4573 283 4574 287
tri 4574 283 4578 287 sw
tri 5376 283 5380 287 se
rect 2768 250 2772 283
tri 2772 250 2805 283 sw
rect 4573 250 4578 283
tri 4578 250 4611 283 sw
tri 5343 250 5376 283 se
rect 5376 250 5380 283
rect 6378 283 6379 287
tri 6379 283 6383 287 sw
tri 7188 283 7192 287 se
rect 6378 250 6383 283
tri 6383 250 6416 283 sw
tri 7155 250 7188 283 se
rect 7188 250 7192 283
tri 8184 283 8188 287 sw
tri 8990 283 8994 287 se
rect 8184 250 8188 283
tri 8188 250 8221 283 sw
tri 8957 250 8990 283 se
rect 8990 250 8994 283
tri 9986 283 9990 287 sw
tri 10794 283 10798 287 se
rect 9986 250 9990 283
tri 9990 250 10023 283 sw
tri 10761 250 10794 283 se
rect 10794 250 10798 283
tri 11790 283 11794 287 sw
tri 12592 283 12596 287 se
rect 11790 250 11794 283
tri 11794 250 11827 283 sw
tri 12559 250 12592 283 se
rect 12592 250 12596 283
tri 13444 250 13481 287 sw
tri 6051 -335 6057 -329 se
tri 6185 -335 6191 -329 sw
tri 2875 -461 2881 -455 ne
tri 3009 -461 3015 -455 nw
tri 5584 -461 5590 -455 ne
tri 5718 -461 5724 -455 nw
<< rmetal1 >>
rect 8526 1032 8528 1033
rect 8526 982 8527 1032
rect 8526 981 8528 982
rect 8564 1032 8566 1033
rect 8565 982 8566 1032
rect 8564 981 8566 982
rect 10395 1032 10397 1033
rect 10433 1032 10435 1033
rect 10395 982 10396 1032
rect 10434 982 10435 1032
rect 10395 981 10397 982
rect 10433 981 10435 982
rect 11229 1032 11231 1033
rect 11267 1032 11269 1033
rect 11229 982 11230 1032
rect 11268 982 11269 1032
rect 11229 981 11231 982
rect 11267 981 11269 982
rect 12199 1032 12201 1033
rect 12199 982 12200 1032
rect 12199 981 12201 982
rect 12237 1032 12239 1033
rect 12238 982 12239 1032
rect 12237 981 12239 982
rect 13116 1032 13118 1033
rect 13154 1032 13156 1033
rect 13116 982 13117 1032
rect 13155 982 13156 1032
rect 13116 981 13118 982
rect 13154 981 13156 982
<< via1 >>
rect 8970 981 9022 1033
rect 9038 981 9090 1033
rect 10746 981 10798 1033
rect 10814 981 10866 1033
rect 11715 981 11767 1033
rect 11783 981 11835 1033
rect 8970 651 9022 703
rect 9038 651 9090 703
rect 10746 651 10798 703
rect 10814 651 10866 703
rect 11715 651 11767 703
rect 11783 651 11835 703
<< metal2 >>
rect -714 20547 -136 20556
rect -714 20491 -711 20547
rect -655 20491 -625 20547
rect -569 20491 -539 20547
rect -483 20491 -453 20547
rect -397 20491 -367 20547
rect -311 20491 -281 20547
rect -225 20491 -195 20547
rect -139 20491 -136 20547
rect -714 20455 -136 20491
rect -714 20399 -711 20455
rect -655 20399 -625 20455
rect -569 20399 -539 20455
rect -483 20399 -453 20455
rect -397 20399 -367 20455
rect -311 20399 -281 20455
rect -225 20399 -195 20455
rect -139 20399 -136 20455
rect -714 20363 -136 20399
rect -714 20307 -711 20363
rect -655 20307 -625 20363
rect -569 20307 -539 20363
rect -483 20307 -453 20363
rect -397 20307 -367 20363
rect -311 20307 -281 20363
rect -225 20307 -195 20363
rect -139 20307 -136 20363
rect -714 20271 -136 20307
rect -714 20215 -711 20271
rect -655 20215 -625 20271
rect -569 20215 -539 20271
rect -483 20215 -453 20271
rect -397 20215 -367 20271
rect -311 20215 -281 20271
rect -225 20215 -195 20271
rect -139 20215 -136 20271
rect -714 20179 -136 20215
rect -714 20123 -711 20179
rect -655 20123 -625 20179
rect -569 20123 -539 20179
rect -483 20123 -453 20179
rect -397 20123 -367 20179
rect -311 20123 -281 20179
rect -225 20123 -195 20179
rect -139 20123 -136 20179
rect -714 20086 -136 20123
rect -714 20030 -711 20086
rect -655 20030 -625 20086
rect -569 20030 -539 20086
rect -483 20030 -453 20086
rect -397 20030 -367 20086
rect -311 20030 -281 20086
rect -225 20030 -195 20086
rect -139 20030 -136 20086
rect -714 19993 -136 20030
rect -714 19937 -711 19993
rect -655 19937 -625 19993
rect -569 19937 -539 19993
rect -483 19937 -453 19993
rect -397 19937 -367 19993
rect -311 19937 -281 19993
rect -225 19937 -195 19993
rect -139 19937 -136 19993
rect -714 19928 -136 19937
rect 1103 20550 1657 20559
rect 1103 20494 1106 20550
rect 1162 20494 1188 20550
rect 1244 20494 1270 20550
rect 1326 20494 1352 20550
rect 1408 20494 1434 20550
rect 1490 20494 1516 20550
rect 1572 20494 1598 20550
rect 1654 20494 1657 20550
rect 1103 20470 1657 20494
rect 1103 20414 1106 20470
rect 1162 20414 1188 20470
rect 1244 20414 1270 20470
rect 1326 20414 1352 20470
rect 1408 20414 1434 20470
rect 1490 20414 1516 20470
rect 1572 20414 1598 20470
rect 1654 20414 1657 20470
rect 1103 20390 1657 20414
rect 1103 20334 1106 20390
rect 1162 20334 1188 20390
rect 1244 20334 1270 20390
rect 1326 20334 1352 20390
rect 1408 20334 1434 20390
rect 1490 20334 1516 20390
rect 1572 20334 1598 20390
rect 1654 20334 1657 20390
rect 1103 20310 1657 20334
rect 1103 20254 1106 20310
rect 1162 20254 1188 20310
rect 1244 20254 1270 20310
rect 1326 20254 1352 20310
rect 1408 20254 1434 20310
rect 1490 20254 1516 20310
rect 1572 20254 1598 20310
rect 1654 20254 1657 20310
rect 1103 20230 1657 20254
rect 1103 20174 1106 20230
rect 1162 20174 1188 20230
rect 1244 20174 1270 20230
rect 1326 20174 1352 20230
rect 1408 20174 1434 20230
rect 1490 20174 1516 20230
rect 1572 20174 1598 20230
rect 1654 20174 1657 20230
rect 1103 20149 1657 20174
rect 1103 20093 1106 20149
rect 1162 20093 1188 20149
rect 1244 20093 1270 20149
rect 1326 20093 1352 20149
rect 1408 20093 1434 20149
rect 1490 20093 1516 20149
rect 1572 20093 1598 20149
rect 1654 20093 1657 20149
rect 1103 20068 1657 20093
rect 1103 20012 1106 20068
rect 1162 20012 1188 20068
rect 1244 20012 1270 20068
rect 1326 20012 1352 20068
rect 1408 20012 1434 20068
rect 1490 20012 1516 20068
rect 1572 20012 1598 20068
rect 1654 20012 1657 20068
rect 1103 19987 1657 20012
rect 1103 19931 1106 19987
rect 1162 19931 1188 19987
rect 1244 19931 1270 19987
rect 1326 19931 1352 19987
rect 1408 19931 1434 19987
rect 1490 19931 1516 19987
rect 1572 19931 1598 19987
rect 1654 19931 1657 19987
rect 1103 19906 1657 19931
rect 1103 19850 1106 19906
rect 1162 19850 1188 19906
rect 1244 19850 1270 19906
rect 1326 19850 1352 19906
rect 1408 19850 1434 19906
rect 1490 19850 1516 19906
rect 1572 19850 1598 19906
rect 1654 19850 1657 19906
rect 1103 19825 1657 19850
rect 1103 19769 1106 19825
rect 1162 19769 1188 19825
rect 1244 19769 1270 19825
rect 1326 19769 1352 19825
rect 1408 19769 1434 19825
rect 1490 19769 1516 19825
rect 1572 19769 1598 19825
rect 1654 19769 1657 19825
rect 1103 19744 1657 19769
rect 1103 19688 1106 19744
rect 1162 19688 1188 19744
rect 1244 19688 1270 19744
rect 1326 19688 1352 19744
rect 1408 19688 1434 19744
rect 1490 19688 1516 19744
rect 1572 19688 1598 19744
rect 1654 19688 1657 19744
rect 1103 19663 1657 19688
rect 1103 19607 1106 19663
rect 1162 19607 1188 19663
rect 1244 19607 1270 19663
rect 1326 19607 1352 19663
rect 1408 19607 1434 19663
rect 1490 19607 1516 19663
rect 1572 19607 1598 19663
rect 1654 19607 1657 19663
rect 1103 19582 1657 19607
rect 1103 19526 1106 19582
rect 1162 19526 1188 19582
rect 1244 19526 1270 19582
rect 1326 19526 1352 19582
rect 1408 19526 1434 19582
rect 1490 19526 1516 19582
rect 1572 19526 1598 19582
rect 1654 19526 1657 19582
rect 1103 19501 1657 19526
rect 1103 19445 1106 19501
rect 1162 19445 1188 19501
rect 1244 19445 1270 19501
rect 1326 19445 1352 19501
rect 1408 19445 1434 19501
rect 1490 19445 1516 19501
rect 1572 19445 1598 19501
rect 1654 19445 1657 19501
rect 1103 19420 1657 19445
rect 1103 19364 1106 19420
rect 1162 19364 1188 19420
rect 1244 19364 1270 19420
rect 1326 19364 1352 19420
rect 1408 19364 1434 19420
rect 1490 19364 1516 19420
rect 1572 19364 1598 19420
rect 1654 19364 1657 19420
rect 1103 19339 1657 19364
rect 1103 19283 1106 19339
rect 1162 19283 1188 19339
rect 1244 19283 1270 19339
rect 1326 19283 1352 19339
rect 1408 19283 1434 19339
rect 1490 19283 1516 19339
rect 1572 19283 1598 19339
rect 1654 19283 1657 19339
rect 1103 19258 1657 19283
rect 1103 19202 1106 19258
rect 1162 19202 1188 19258
rect 1244 19202 1270 19258
rect 1326 19202 1352 19258
rect 1408 19202 1434 19258
rect 1490 19202 1516 19258
rect 1572 19202 1598 19258
rect 1654 19202 1657 19258
rect 1103 19177 1657 19202
rect 1103 19121 1106 19177
rect 1162 19121 1188 19177
rect 1244 19121 1270 19177
rect 1326 19121 1352 19177
rect 1408 19121 1434 19177
rect 1490 19121 1516 19177
rect 1572 19121 1598 19177
rect 1654 19121 1657 19177
rect 1103 19096 1657 19121
rect 1103 19040 1106 19096
rect 1162 19040 1188 19096
rect 1244 19040 1270 19096
rect 1326 19040 1352 19096
rect 1408 19040 1434 19096
rect 1490 19040 1516 19096
rect 1572 19040 1598 19096
rect 1654 19040 1657 19096
rect 1103 19031 1657 19040
rect 2907 20550 3461 20559
rect 2907 20494 2910 20550
rect 2966 20494 2992 20550
rect 3048 20494 3074 20550
rect 3130 20494 3156 20550
rect 3212 20494 3238 20550
rect 3294 20494 3320 20550
rect 3376 20494 3402 20550
rect 3458 20494 3461 20550
rect 2907 20470 3461 20494
rect 2907 20414 2910 20470
rect 2966 20414 2992 20470
rect 3048 20414 3074 20470
rect 3130 20414 3156 20470
rect 3212 20414 3238 20470
rect 3294 20414 3320 20470
rect 3376 20414 3402 20470
rect 3458 20414 3461 20470
rect 2907 20390 3461 20414
rect 2907 20334 2910 20390
rect 2966 20334 2992 20390
rect 3048 20334 3074 20390
rect 3130 20334 3156 20390
rect 3212 20334 3238 20390
rect 3294 20334 3320 20390
rect 3376 20334 3402 20390
rect 3458 20334 3461 20390
rect 2907 20310 3461 20334
rect 2907 20254 2910 20310
rect 2966 20254 2992 20310
rect 3048 20254 3074 20310
rect 3130 20254 3156 20310
rect 3212 20254 3238 20310
rect 3294 20254 3320 20310
rect 3376 20254 3402 20310
rect 3458 20254 3461 20310
rect 2907 20230 3461 20254
rect 2907 20174 2910 20230
rect 2966 20174 2992 20230
rect 3048 20174 3074 20230
rect 3130 20174 3156 20230
rect 3212 20174 3238 20230
rect 3294 20174 3320 20230
rect 3376 20174 3402 20230
rect 3458 20174 3461 20230
rect 2907 20149 3461 20174
rect 2907 20093 2910 20149
rect 2966 20093 2992 20149
rect 3048 20093 3074 20149
rect 3130 20093 3156 20149
rect 3212 20093 3238 20149
rect 3294 20093 3320 20149
rect 3376 20093 3402 20149
rect 3458 20093 3461 20149
rect 2907 20068 3461 20093
rect 2907 20012 2910 20068
rect 2966 20012 2992 20068
rect 3048 20012 3074 20068
rect 3130 20012 3156 20068
rect 3212 20012 3238 20068
rect 3294 20012 3320 20068
rect 3376 20012 3402 20068
rect 3458 20012 3461 20068
rect 2907 19987 3461 20012
rect 2907 19931 2910 19987
rect 2966 19931 2992 19987
rect 3048 19931 3074 19987
rect 3130 19931 3156 19987
rect 3212 19931 3238 19987
rect 3294 19931 3320 19987
rect 3376 19931 3402 19987
rect 3458 19931 3461 19987
rect 2907 19906 3461 19931
rect 2907 19850 2910 19906
rect 2966 19850 2992 19906
rect 3048 19850 3074 19906
rect 3130 19850 3156 19906
rect 3212 19850 3238 19906
rect 3294 19850 3320 19906
rect 3376 19850 3402 19906
rect 3458 19850 3461 19906
rect 2907 19825 3461 19850
rect 2907 19769 2910 19825
rect 2966 19769 2992 19825
rect 3048 19769 3074 19825
rect 3130 19769 3156 19825
rect 3212 19769 3238 19825
rect 3294 19769 3320 19825
rect 3376 19769 3402 19825
rect 3458 19769 3461 19825
rect 2907 19744 3461 19769
rect 2907 19688 2910 19744
rect 2966 19688 2992 19744
rect 3048 19688 3074 19744
rect 3130 19688 3156 19744
rect 3212 19688 3238 19744
rect 3294 19688 3320 19744
rect 3376 19688 3402 19744
rect 3458 19688 3461 19744
rect 2907 19663 3461 19688
rect 2907 19607 2910 19663
rect 2966 19607 2992 19663
rect 3048 19607 3074 19663
rect 3130 19607 3156 19663
rect 3212 19607 3238 19663
rect 3294 19607 3320 19663
rect 3376 19607 3402 19663
rect 3458 19607 3461 19663
rect 2907 19582 3461 19607
rect 2907 19526 2910 19582
rect 2966 19526 2992 19582
rect 3048 19526 3074 19582
rect 3130 19526 3156 19582
rect 3212 19526 3238 19582
rect 3294 19526 3320 19582
rect 3376 19526 3402 19582
rect 3458 19526 3461 19582
rect 2907 19501 3461 19526
rect 2907 19445 2910 19501
rect 2966 19445 2992 19501
rect 3048 19445 3074 19501
rect 3130 19445 3156 19501
rect 3212 19445 3238 19501
rect 3294 19445 3320 19501
rect 3376 19445 3402 19501
rect 3458 19445 3461 19501
rect 2907 19420 3461 19445
rect 2907 19364 2910 19420
rect 2966 19364 2992 19420
rect 3048 19364 3074 19420
rect 3130 19364 3156 19420
rect 3212 19364 3238 19420
rect 3294 19364 3320 19420
rect 3376 19364 3402 19420
rect 3458 19364 3461 19420
rect 2907 19339 3461 19364
rect 2907 19283 2910 19339
rect 2966 19283 2992 19339
rect 3048 19283 3074 19339
rect 3130 19283 3156 19339
rect 3212 19283 3238 19339
rect 3294 19283 3320 19339
rect 3376 19283 3402 19339
rect 3458 19283 3461 19339
rect 2907 19258 3461 19283
rect 2907 19202 2910 19258
rect 2966 19202 2992 19258
rect 3048 19202 3074 19258
rect 3130 19202 3156 19258
rect 3212 19202 3238 19258
rect 3294 19202 3320 19258
rect 3376 19202 3402 19258
rect 3458 19202 3461 19258
rect 2907 19177 3461 19202
rect 2907 19121 2910 19177
rect 2966 19121 2992 19177
rect 3048 19121 3074 19177
rect 3130 19121 3156 19177
rect 3212 19121 3238 19177
rect 3294 19121 3320 19177
rect 3376 19121 3402 19177
rect 3458 19121 3461 19177
rect 2907 19096 3461 19121
rect 2907 19040 2910 19096
rect 2966 19040 2992 19096
rect 3048 19040 3074 19096
rect 3130 19040 3156 19096
rect 3212 19040 3238 19096
rect 3294 19040 3320 19096
rect 3376 19040 3402 19096
rect 3458 19040 3461 19096
rect 2907 19031 3461 19040
rect 4705 20550 5259 20559
rect 4705 20494 4708 20550
rect 4764 20494 4790 20550
rect 4846 20494 4872 20550
rect 4928 20494 4954 20550
rect 5010 20494 5036 20550
rect 5092 20494 5118 20550
rect 5174 20494 5200 20550
rect 5256 20494 5259 20550
rect 4705 20470 5259 20494
rect 4705 20414 4708 20470
rect 4764 20414 4790 20470
rect 4846 20414 4872 20470
rect 4928 20414 4954 20470
rect 5010 20414 5036 20470
rect 5092 20414 5118 20470
rect 5174 20414 5200 20470
rect 5256 20414 5259 20470
rect 4705 20390 5259 20414
rect 4705 20334 4708 20390
rect 4764 20334 4790 20390
rect 4846 20334 4872 20390
rect 4928 20334 4954 20390
rect 5010 20334 5036 20390
rect 5092 20334 5118 20390
rect 5174 20334 5200 20390
rect 5256 20334 5259 20390
rect 4705 20310 5259 20334
rect 4705 20254 4708 20310
rect 4764 20254 4790 20310
rect 4846 20254 4872 20310
rect 4928 20254 4954 20310
rect 5010 20254 5036 20310
rect 5092 20254 5118 20310
rect 5174 20254 5200 20310
rect 5256 20254 5259 20310
rect 4705 20230 5259 20254
rect 4705 20174 4708 20230
rect 4764 20174 4790 20230
rect 4846 20174 4872 20230
rect 4928 20174 4954 20230
rect 5010 20174 5036 20230
rect 5092 20174 5118 20230
rect 5174 20174 5200 20230
rect 5256 20174 5259 20230
rect 4705 20149 5259 20174
rect 4705 20093 4708 20149
rect 4764 20093 4790 20149
rect 4846 20093 4872 20149
rect 4928 20093 4954 20149
rect 5010 20093 5036 20149
rect 5092 20093 5118 20149
rect 5174 20093 5200 20149
rect 5256 20093 5259 20149
rect 4705 20068 5259 20093
rect 4705 20012 4708 20068
rect 4764 20012 4790 20068
rect 4846 20012 4872 20068
rect 4928 20012 4954 20068
rect 5010 20012 5036 20068
rect 5092 20012 5118 20068
rect 5174 20012 5200 20068
rect 5256 20012 5259 20068
rect 4705 19987 5259 20012
rect 4705 19931 4708 19987
rect 4764 19931 4790 19987
rect 4846 19931 4872 19987
rect 4928 19931 4954 19987
rect 5010 19931 5036 19987
rect 5092 19931 5118 19987
rect 5174 19931 5200 19987
rect 5256 19931 5259 19987
rect 4705 19906 5259 19931
rect 4705 19850 4708 19906
rect 4764 19850 4790 19906
rect 4846 19850 4872 19906
rect 4928 19850 4954 19906
rect 5010 19850 5036 19906
rect 5092 19850 5118 19906
rect 5174 19850 5200 19906
rect 5256 19850 5259 19906
rect 4705 19825 5259 19850
rect 4705 19769 4708 19825
rect 4764 19769 4790 19825
rect 4846 19769 4872 19825
rect 4928 19769 4954 19825
rect 5010 19769 5036 19825
rect 5092 19769 5118 19825
rect 5174 19769 5200 19825
rect 5256 19769 5259 19825
rect 4705 19744 5259 19769
rect 4705 19688 4708 19744
rect 4764 19688 4790 19744
rect 4846 19688 4872 19744
rect 4928 19688 4954 19744
rect 5010 19688 5036 19744
rect 5092 19688 5118 19744
rect 5174 19688 5200 19744
rect 5256 19688 5259 19744
rect 4705 19663 5259 19688
rect 4705 19607 4708 19663
rect 4764 19607 4790 19663
rect 4846 19607 4872 19663
rect 4928 19607 4954 19663
rect 5010 19607 5036 19663
rect 5092 19607 5118 19663
rect 5174 19607 5200 19663
rect 5256 19607 5259 19663
rect 4705 19582 5259 19607
rect 4705 19526 4708 19582
rect 4764 19526 4790 19582
rect 4846 19526 4872 19582
rect 4928 19526 4954 19582
rect 5010 19526 5036 19582
rect 5092 19526 5118 19582
rect 5174 19526 5200 19582
rect 5256 19526 5259 19582
rect 4705 19501 5259 19526
rect 4705 19445 4708 19501
rect 4764 19445 4790 19501
rect 4846 19445 4872 19501
rect 4928 19445 4954 19501
rect 5010 19445 5036 19501
rect 5092 19445 5118 19501
rect 5174 19445 5200 19501
rect 5256 19445 5259 19501
rect 4705 19420 5259 19445
rect 4705 19364 4708 19420
rect 4764 19364 4790 19420
rect 4846 19364 4872 19420
rect 4928 19364 4954 19420
rect 5010 19364 5036 19420
rect 5092 19364 5118 19420
rect 5174 19364 5200 19420
rect 5256 19364 5259 19420
rect 4705 19339 5259 19364
rect 4705 19283 4708 19339
rect 4764 19283 4790 19339
rect 4846 19283 4872 19339
rect 4928 19283 4954 19339
rect 5010 19283 5036 19339
rect 5092 19283 5118 19339
rect 5174 19283 5200 19339
rect 5256 19283 5259 19339
rect 4705 19258 5259 19283
rect 4705 19202 4708 19258
rect 4764 19202 4790 19258
rect 4846 19202 4872 19258
rect 4928 19202 4954 19258
rect 5010 19202 5036 19258
rect 5092 19202 5118 19258
rect 5174 19202 5200 19258
rect 5256 19202 5259 19258
rect 4705 19177 5259 19202
rect 4705 19121 4708 19177
rect 4764 19121 4790 19177
rect 4846 19121 4872 19177
rect 4928 19121 4954 19177
rect 5010 19121 5036 19177
rect 5092 19121 5118 19177
rect 5174 19121 5200 19177
rect 5256 19121 5259 19177
rect 4705 19096 5259 19121
rect 4705 19040 4708 19096
rect 4764 19040 4790 19096
rect 4846 19040 4872 19096
rect 4928 19040 4954 19096
rect 5010 19040 5036 19096
rect 5092 19040 5118 19096
rect 5174 19040 5200 19096
rect 5256 19040 5259 19096
rect 4705 19031 5259 19040
rect 6378 20550 6754 20559
rect 6378 20149 6754 20174
rect 6434 20093 6458 20149
rect 6514 20093 6538 20149
rect 6594 20093 6618 20149
rect 6674 20093 6698 20149
rect 6378 20068 6754 20093
rect 6434 20012 6458 20068
rect 6514 20012 6538 20068
rect 6594 20012 6618 20068
rect 6674 20012 6698 20068
rect 6378 19987 6754 20012
rect 6434 19931 6458 19987
rect 6514 19931 6538 19987
rect 6594 19931 6618 19987
rect 6674 19931 6698 19987
rect 6378 19906 6754 19931
rect 6434 19850 6458 19906
rect 6514 19850 6538 19906
rect 6594 19850 6618 19906
rect 6674 19850 6698 19906
rect 6378 19825 6754 19850
rect 6434 19769 6458 19825
rect 6514 19769 6538 19825
rect 6594 19769 6618 19825
rect 6674 19769 6698 19825
rect 6378 19744 6754 19769
rect 6434 19688 6458 19744
rect 6514 19688 6538 19744
rect 6594 19688 6618 19744
rect 6674 19688 6698 19744
rect 6378 19663 6754 19688
rect 6434 19607 6458 19663
rect 6514 19607 6538 19663
rect 6594 19607 6618 19663
rect 6674 19607 6698 19663
rect 6378 19582 6754 19607
rect 6434 19526 6458 19582
rect 6514 19526 6538 19582
rect 6594 19526 6618 19582
rect 6674 19526 6698 19582
rect 6378 19501 6754 19526
rect 6434 19445 6458 19501
rect 6514 19445 6538 19501
rect 6594 19445 6618 19501
rect 6674 19445 6698 19501
rect 6378 19420 6754 19445
rect 6434 19364 6458 19420
rect 6514 19364 6538 19420
rect 6594 19364 6618 19420
rect 6674 19364 6698 19420
rect 6378 19339 6754 19364
rect 6434 19283 6458 19339
rect 6514 19283 6538 19339
rect 6594 19283 6618 19339
rect 6674 19283 6698 19339
rect 6378 19258 6754 19283
rect 6434 19202 6458 19258
rect 6514 19202 6538 19258
rect 6594 19202 6618 19258
rect 6674 19202 6698 19258
rect 6378 19177 6754 19202
rect 6434 19121 6458 19177
rect 6514 19121 6538 19177
rect 6594 19121 6618 19177
rect 6674 19121 6698 19177
rect 6378 19096 6754 19121
rect 6434 19040 6458 19096
rect 6514 19040 6538 19096
rect 6594 19040 6618 19096
rect 6674 19040 6698 19096
rect 6378 19031 6754 19040
rect 8067 20556 8327 20565
rect 8123 20500 8169 20556
rect 8225 20500 8271 20556
rect 8067 20475 8327 20500
rect 8123 20419 8169 20475
rect 8225 20419 8271 20475
rect 8067 20394 8327 20419
rect 8123 20338 8169 20394
rect 8225 20338 8271 20394
rect 8067 20313 8327 20338
rect 8123 20257 8169 20313
rect 8225 20257 8271 20313
rect 8067 20232 8327 20257
rect 8123 20176 8169 20232
rect 8225 20176 8271 20232
rect 8067 20151 8327 20176
rect 8123 20095 8169 20151
rect 8225 20095 8271 20151
rect 8067 20070 8327 20095
rect 8123 20014 8169 20070
rect 8225 20014 8271 20070
rect 8067 19989 8327 20014
rect 8123 19933 8169 19989
rect 8225 19933 8271 19989
rect 8067 19908 8327 19933
rect 8123 19852 8169 19908
rect 8225 19852 8271 19908
rect 8067 19827 8327 19852
rect 8123 19771 8169 19827
rect 8225 19771 8271 19827
rect 8067 19745 8327 19771
rect 8123 19689 8169 19745
rect 8225 19689 8271 19745
rect 8067 19663 8327 19689
rect 8123 19607 8169 19663
rect 8225 19607 8271 19663
rect 8067 19581 8327 19607
rect 8123 19525 8169 19581
rect 8225 19525 8271 19581
rect 8067 19499 8327 19525
rect 8123 19443 8169 19499
rect 8225 19443 8271 19499
rect 8067 19417 8327 19443
rect 8123 19361 8169 19417
rect 8225 19361 8271 19417
rect 8067 19335 8327 19361
rect 8123 19279 8169 19335
rect 8225 19279 8271 19335
rect 8067 19253 8327 19279
rect 8123 19197 8169 19253
rect 8225 19197 8271 19253
rect 8067 19171 8327 19197
rect 8123 19115 8169 19171
rect 8225 19115 8271 19171
rect 8067 19089 8327 19115
rect 8123 19033 8169 19089
rect 8225 19033 8271 19089
rect 8067 19024 8327 19033
rect 8894 20556 9142 20565
rect 8950 20500 8990 20556
rect 9046 20500 9086 20556
rect 8894 20475 9142 20500
rect 8950 20419 8990 20475
rect 9046 20419 9086 20475
rect 8894 20394 9142 20419
rect 8950 20338 8990 20394
rect 9046 20338 9086 20394
rect 8894 20313 9142 20338
rect 8950 20257 8990 20313
rect 9046 20257 9086 20313
rect 8894 20232 9142 20257
rect 8950 20176 8990 20232
rect 9046 20176 9086 20232
rect 8894 20151 9142 20176
rect 8950 20095 8990 20151
rect 9046 20095 9086 20151
rect 8894 20070 9142 20095
rect 8950 20014 8990 20070
rect 9046 20014 9086 20070
rect 8894 19989 9142 20014
rect 8950 19933 8990 19989
rect 9046 19933 9086 19989
rect 8894 19908 9142 19933
rect 8950 19852 8990 19908
rect 9046 19852 9086 19908
rect 8894 19827 9142 19852
rect 8950 19771 8990 19827
rect 9046 19771 9086 19827
rect 8894 19745 9142 19771
rect 8950 19689 8990 19745
rect 9046 19689 9086 19745
rect 8894 19663 9142 19689
rect 8950 19607 8990 19663
rect 9046 19607 9086 19663
rect 8894 19581 9142 19607
rect 8950 19525 8990 19581
rect 9046 19525 9086 19581
rect 8894 19499 9142 19525
rect 8950 19443 8990 19499
rect 9046 19443 9086 19499
rect 8894 19417 9142 19443
rect 8950 19361 8990 19417
rect 9046 19361 9086 19417
rect 8894 19335 9142 19361
rect 8950 19279 8990 19335
rect 9046 19279 9086 19335
rect 8894 19253 9142 19279
rect 8950 19197 8990 19253
rect 9046 19197 9086 19253
rect 8894 19171 9142 19197
rect 8950 19115 8990 19171
rect 9046 19115 9086 19171
rect 8894 19089 9142 19115
rect 8950 19033 8990 19089
rect 9046 19033 9086 19089
rect 10123 20550 10677 20559
rect 10123 20494 10126 20550
rect 10182 20494 10208 20550
rect 10264 20494 10290 20550
rect 10346 20494 10372 20550
rect 10428 20494 10454 20550
rect 10510 20494 10536 20550
rect 10592 20494 10618 20550
rect 10674 20494 10677 20550
rect 10123 20467 10677 20494
rect 10123 20411 10126 20467
rect 10182 20411 10208 20467
rect 10264 20411 10290 20467
rect 10346 20411 10372 20467
rect 10428 20411 10454 20467
rect 10510 20411 10536 20467
rect 10592 20411 10618 20467
rect 10674 20411 10677 20467
rect 10123 20384 10677 20411
rect 10123 20328 10126 20384
rect 10182 20328 10208 20384
rect 10264 20328 10290 20384
rect 10346 20328 10372 20384
rect 10428 20328 10454 20384
rect 10510 20328 10536 20384
rect 10592 20328 10618 20384
rect 10674 20328 10677 20384
rect 10123 20301 10677 20328
rect 10123 20245 10126 20301
rect 10182 20245 10208 20301
rect 10264 20245 10290 20301
rect 10346 20245 10372 20301
rect 10428 20245 10454 20301
rect 10510 20245 10536 20301
rect 10592 20245 10618 20301
rect 10674 20245 10677 20301
rect 10123 20217 10677 20245
rect 10123 20161 10126 20217
rect 10182 20161 10208 20217
rect 10264 20161 10290 20217
rect 10346 20161 10372 20217
rect 10428 20161 10454 20217
rect 10510 20161 10536 20217
rect 10592 20161 10618 20217
rect 10674 20161 10677 20217
rect 10123 20133 10677 20161
rect 10123 20077 10126 20133
rect 10182 20077 10208 20133
rect 10264 20077 10290 20133
rect 10346 20077 10372 20133
rect 10428 20077 10454 20133
rect 10510 20077 10536 20133
rect 10592 20077 10618 20133
rect 10674 20077 10677 20133
rect 10123 20049 10677 20077
rect 10123 19993 10126 20049
rect 10182 19993 10208 20049
rect 10264 19993 10290 20049
rect 10346 19993 10372 20049
rect 10428 19993 10454 20049
rect 10510 19993 10536 20049
rect 10592 19993 10618 20049
rect 10674 19993 10677 20049
rect 10123 19965 10677 19993
rect 10123 19909 10126 19965
rect 10182 19909 10208 19965
rect 10264 19909 10290 19965
rect 10346 19909 10372 19965
rect 10428 19909 10454 19965
rect 10510 19909 10536 19965
rect 10592 19909 10618 19965
rect 10674 19909 10677 19965
rect 10123 19881 10677 19909
rect 10123 19825 10126 19881
rect 10182 19825 10208 19881
rect 10264 19825 10290 19881
rect 10346 19825 10372 19881
rect 10428 19825 10454 19881
rect 10510 19825 10536 19881
rect 10592 19825 10618 19881
rect 10674 19825 10677 19881
rect 10123 19797 10677 19825
rect 10123 19741 10126 19797
rect 10182 19741 10208 19797
rect 10264 19741 10290 19797
rect 10346 19741 10372 19797
rect 10428 19741 10454 19797
rect 10510 19741 10536 19797
rect 10592 19741 10618 19797
rect 10674 19741 10677 19797
rect 10123 19713 10677 19741
rect 10123 19657 10126 19713
rect 10182 19657 10208 19713
rect 10264 19657 10290 19713
rect 10346 19657 10372 19713
rect 10428 19657 10454 19713
rect 10510 19657 10536 19713
rect 10592 19657 10618 19713
rect 10674 19657 10677 19713
rect 10123 19629 10677 19657
rect 10123 19573 10126 19629
rect 10182 19573 10208 19629
rect 10264 19573 10290 19629
rect 10346 19573 10372 19629
rect 10428 19573 10454 19629
rect 10510 19573 10536 19629
rect 10592 19573 10618 19629
rect 10674 19573 10677 19629
rect 10123 19545 10677 19573
rect 10123 19489 10126 19545
rect 10182 19489 10208 19545
rect 10264 19489 10290 19545
rect 10346 19489 10372 19545
rect 10428 19489 10454 19545
rect 10510 19489 10536 19545
rect 10592 19489 10618 19545
rect 10674 19489 10677 19545
rect 10123 19461 10677 19489
rect 10123 19405 10126 19461
rect 10182 19405 10208 19461
rect 10264 19405 10290 19461
rect 10346 19405 10372 19461
rect 10428 19405 10454 19461
rect 10510 19405 10536 19461
rect 10592 19405 10618 19461
rect 10674 19405 10677 19461
rect 10123 19377 10677 19405
rect 10123 19321 10126 19377
rect 10182 19321 10208 19377
rect 10264 19321 10290 19377
rect 10346 19321 10372 19377
rect 10428 19321 10454 19377
rect 10510 19321 10536 19377
rect 10592 19321 10618 19377
rect 10674 19321 10677 19377
rect 10123 19293 10677 19321
rect 10123 19237 10126 19293
rect 10182 19237 10208 19293
rect 10264 19237 10290 19293
rect 10346 19237 10372 19293
rect 10428 19237 10454 19293
rect 10510 19237 10536 19293
rect 10592 19237 10618 19293
rect 10674 19237 10677 19293
rect 10123 19209 10677 19237
rect 10123 19153 10126 19209
rect 10182 19153 10208 19209
rect 10264 19153 10290 19209
rect 10346 19153 10372 19209
rect 10428 19153 10454 19209
rect 10510 19153 10536 19209
rect 10592 19153 10618 19209
rect 10674 19153 10677 19209
rect 10123 19125 10677 19153
rect 10123 19069 10126 19125
rect 10182 19069 10208 19125
rect 10264 19069 10290 19125
rect 10346 19069 10372 19125
rect 10428 19069 10454 19125
rect 10510 19069 10536 19125
rect 10592 19069 10618 19125
rect 10674 19069 10677 19125
rect 10123 19060 10677 19069
rect 11924 20550 12478 20559
rect 11924 20494 11927 20550
rect 11983 20494 12009 20550
rect 12065 20494 12091 20550
rect 12147 20494 12173 20550
rect 12229 20494 12255 20550
rect 12311 20494 12337 20550
rect 12393 20494 12419 20550
rect 12475 20494 12478 20550
rect 11924 20467 12478 20494
rect 11924 20411 11927 20467
rect 11983 20411 12009 20467
rect 12065 20411 12091 20467
rect 12147 20411 12173 20467
rect 12229 20411 12255 20467
rect 12311 20411 12337 20467
rect 12393 20411 12419 20467
rect 12475 20411 12478 20467
rect 11924 20384 12478 20411
rect 11924 20328 11927 20384
rect 11983 20328 12009 20384
rect 12065 20328 12091 20384
rect 12147 20328 12173 20384
rect 12229 20328 12255 20384
rect 12311 20328 12337 20384
rect 12393 20328 12419 20384
rect 12475 20328 12478 20384
rect 11924 20301 12478 20328
rect 11924 20245 11927 20301
rect 11983 20245 12009 20301
rect 12065 20245 12091 20301
rect 12147 20245 12173 20301
rect 12229 20245 12255 20301
rect 12311 20245 12337 20301
rect 12393 20245 12419 20301
rect 12475 20245 12478 20301
rect 11924 20217 12478 20245
rect 11924 20161 11927 20217
rect 11983 20161 12009 20217
rect 12065 20161 12091 20217
rect 12147 20161 12173 20217
rect 12229 20161 12255 20217
rect 12311 20161 12337 20217
rect 12393 20161 12419 20217
rect 12475 20161 12478 20217
rect 11924 20133 12478 20161
rect 11924 20077 11927 20133
rect 11983 20077 12009 20133
rect 12065 20077 12091 20133
rect 12147 20077 12173 20133
rect 12229 20077 12255 20133
rect 12311 20077 12337 20133
rect 12393 20077 12419 20133
rect 12475 20077 12478 20133
rect 11924 20049 12478 20077
rect 11924 19993 11927 20049
rect 11983 19993 12009 20049
rect 12065 19993 12091 20049
rect 12147 19993 12173 20049
rect 12229 19993 12255 20049
rect 12311 19993 12337 20049
rect 12393 19993 12419 20049
rect 12475 19993 12478 20049
rect 11924 19965 12478 19993
rect 11924 19909 11927 19965
rect 11983 19909 12009 19965
rect 12065 19909 12091 19965
rect 12147 19909 12173 19965
rect 12229 19909 12255 19965
rect 12311 19909 12337 19965
rect 12393 19909 12419 19965
rect 12475 19909 12478 19965
rect 11924 19881 12478 19909
rect 11924 19825 11927 19881
rect 11983 19825 12009 19881
rect 12065 19825 12091 19881
rect 12147 19825 12173 19881
rect 12229 19825 12255 19881
rect 12311 19825 12337 19881
rect 12393 19825 12419 19881
rect 12475 19825 12478 19881
rect 11924 19797 12478 19825
rect 11924 19741 11927 19797
rect 11983 19741 12009 19797
rect 12065 19741 12091 19797
rect 12147 19741 12173 19797
rect 12229 19741 12255 19797
rect 12311 19741 12337 19797
rect 12393 19741 12419 19797
rect 12475 19741 12478 19797
rect 11924 19713 12478 19741
rect 11924 19657 11927 19713
rect 11983 19657 12009 19713
rect 12065 19657 12091 19713
rect 12147 19657 12173 19713
rect 12229 19657 12255 19713
rect 12311 19657 12337 19713
rect 12393 19657 12419 19713
rect 12475 19657 12478 19713
rect 11924 19629 12478 19657
rect 11924 19573 11927 19629
rect 11983 19573 12009 19629
rect 12065 19573 12091 19629
rect 12147 19573 12173 19629
rect 12229 19573 12255 19629
rect 12311 19573 12337 19629
rect 12393 19573 12419 19629
rect 12475 19573 12478 19629
rect 11924 19545 12478 19573
rect 11924 19489 11927 19545
rect 11983 19489 12009 19545
rect 12065 19489 12091 19545
rect 12147 19489 12173 19545
rect 12229 19489 12255 19545
rect 12311 19489 12337 19545
rect 12393 19489 12419 19545
rect 12475 19489 12478 19545
rect 11924 19461 12478 19489
rect 11924 19405 11927 19461
rect 11983 19405 12009 19461
rect 12065 19405 12091 19461
rect 12147 19405 12173 19461
rect 12229 19405 12255 19461
rect 12311 19405 12337 19461
rect 12393 19405 12419 19461
rect 12475 19405 12478 19461
rect 11924 19377 12478 19405
rect 11924 19321 11927 19377
rect 11983 19321 12009 19377
rect 12065 19321 12091 19377
rect 12147 19321 12173 19377
rect 12229 19321 12255 19377
rect 12311 19321 12337 19377
rect 12393 19321 12419 19377
rect 12475 19321 12478 19377
rect 11924 19293 12478 19321
rect 11924 19237 11927 19293
rect 11983 19237 12009 19293
rect 12065 19237 12091 19293
rect 12147 19237 12173 19293
rect 12229 19237 12255 19293
rect 12311 19237 12337 19293
rect 12393 19237 12419 19293
rect 12475 19237 12478 19293
rect 11924 19209 12478 19237
rect 11924 19153 11927 19209
rect 11983 19153 12009 19209
rect 12065 19153 12091 19209
rect 12147 19153 12173 19209
rect 12229 19153 12255 19209
rect 12311 19153 12337 19209
rect 12393 19153 12419 19209
rect 12475 19153 12478 19209
rect 11924 19125 12478 19153
rect 11924 19069 11927 19125
rect 11983 19069 12009 19125
rect 12065 19069 12091 19125
rect 12147 19069 12173 19125
rect 12229 19069 12255 19125
rect 12311 19069 12337 19125
rect 12393 19069 12419 19125
rect 12475 19069 12478 19125
rect 11924 19060 12478 19069
rect 8894 19024 9142 19033
tri -639 12842 -421 13060 se
rect -421 12842 -122 13060
rect 2903 13046 3469 13055
rect 2903 12990 2906 13046
rect 2962 12990 2990 13046
rect 3046 12990 3074 13046
rect 3130 12990 3158 13046
rect 3214 12990 3242 13046
rect 3298 12990 3326 13046
rect 3382 12990 3410 13046
rect 3466 12990 3469 13046
rect 2903 12957 3469 12990
rect -724 12833 -122 12842
rect -724 12777 -714 12833
rect -658 12777 -626 12833
rect -570 12777 -538 12833
rect -482 12777 -450 12833
rect -394 12777 -362 12833
rect -306 12777 -274 12833
rect -218 12777 -186 12833
rect -130 12777 -122 12833
rect -724 12753 -122 12777
rect -724 12697 -714 12753
rect -658 12697 -626 12753
rect -570 12697 -538 12753
rect -482 12697 -450 12753
rect -394 12697 -362 12753
rect -306 12697 -274 12753
rect -218 12697 -186 12753
rect -130 12697 -122 12753
rect -724 12673 -122 12697
rect -724 12617 -714 12673
rect -658 12617 -626 12673
rect -570 12617 -538 12673
rect -482 12617 -450 12673
rect -394 12617 -362 12673
rect -306 12617 -274 12673
rect -218 12617 -186 12673
rect -130 12617 -122 12673
rect -724 12593 -122 12617
rect -724 12537 -714 12593
rect -658 12537 -626 12593
rect -570 12537 -538 12593
rect -482 12537 -450 12593
rect -394 12537 -362 12593
rect -306 12537 -274 12593
rect -218 12537 -186 12593
rect -130 12537 -122 12593
rect -724 12513 -122 12537
rect -724 12457 -714 12513
rect -658 12457 -626 12513
rect -570 12457 -538 12513
rect -482 12457 -450 12513
rect -394 12457 -362 12513
rect -306 12457 -274 12513
rect -218 12457 -186 12513
rect -130 12457 -122 12513
rect 1106 12927 1657 12929
rect 1106 12871 1115 12927
rect 1171 12871 1211 12927
rect 1267 12871 1307 12927
rect 1363 12871 1402 12927
rect 1458 12871 1497 12927
rect 1553 12871 1592 12927
rect 1648 12871 1657 12927
rect 1106 12843 1657 12871
rect 1106 12787 1115 12843
rect 1171 12787 1211 12843
rect 1267 12787 1307 12843
rect 1363 12787 1402 12843
rect 1458 12787 1497 12843
rect 1553 12787 1592 12843
rect 1648 12787 1657 12843
rect 1106 12759 1657 12787
rect 1106 12703 1115 12759
rect 1171 12703 1211 12759
rect 1267 12703 1307 12759
rect 1363 12703 1402 12759
rect 1458 12703 1497 12759
rect 1553 12703 1592 12759
rect 1648 12703 1657 12759
rect 1106 12675 1657 12703
rect 1106 12619 1115 12675
rect 1171 12619 1211 12675
rect 1267 12619 1307 12675
rect 1363 12619 1402 12675
rect 1458 12619 1497 12675
rect 1553 12619 1592 12675
rect 1648 12619 1657 12675
rect 1106 12591 1657 12619
rect 1106 12535 1115 12591
rect 1171 12535 1211 12591
rect 1267 12535 1307 12591
rect 1363 12535 1402 12591
rect 1458 12535 1497 12591
rect 1553 12535 1592 12591
rect 1648 12535 1657 12591
rect 1106 12507 1657 12535
rect -724 12433 -122 12457
tri 1075 12449 1106 12480 ne
rect 1106 12451 1115 12507
rect 1171 12451 1211 12507
rect 1267 12451 1307 12507
rect 1363 12451 1402 12507
rect 1458 12451 1497 12507
rect 1553 12451 1592 12507
rect 1648 12451 1657 12507
rect 2903 12901 2906 12957
rect 2962 12901 2990 12957
rect 3046 12901 3074 12957
rect 3130 12901 3158 12957
rect 3214 12901 3242 12957
rect 3298 12901 3326 12957
rect 3382 12901 3410 12957
rect 3466 12901 3469 12957
rect 2903 12868 3469 12901
rect 2903 12812 2906 12868
rect 2962 12812 2990 12868
rect 3046 12812 3074 12868
rect 3130 12812 3158 12868
rect 3214 12812 3242 12868
rect 3298 12812 3326 12868
rect 3382 12812 3410 12868
rect 3466 12812 3469 12868
rect 2903 12779 3469 12812
rect 2903 12723 2906 12779
rect 2962 12723 2990 12779
rect 3046 12723 3074 12779
rect 3130 12723 3158 12779
rect 3214 12723 3242 12779
rect 3298 12723 3326 12779
rect 3382 12723 3410 12779
rect 3466 12723 3469 12779
rect 2903 12690 3469 12723
rect 2903 12634 2906 12690
rect 2962 12634 2990 12690
rect 3046 12634 3074 12690
rect 3130 12634 3158 12690
rect 3214 12634 3242 12690
rect 3298 12634 3326 12690
rect 3382 12634 3410 12690
rect 3466 12634 3469 12690
rect 2903 12601 3469 12634
rect 2903 12545 2906 12601
rect 2962 12545 2990 12601
rect 3046 12545 3074 12601
rect 3130 12545 3158 12601
rect 3214 12545 3242 12601
rect 3298 12545 3326 12601
rect 3382 12545 3410 12601
rect 3466 12545 3469 12601
rect 2903 12511 3469 12545
rect 1106 12449 1657 12451
tri 1657 12449 1688 12480 nw
rect 2903 12455 2906 12511
rect 2962 12455 2990 12511
rect 3046 12455 3074 12511
rect 3130 12455 3158 12511
rect 3214 12455 3242 12511
rect 3298 12455 3326 12511
rect 3382 12455 3410 12511
rect 3466 12455 3469 12511
rect 4701 13046 5267 13055
rect 4701 12990 4704 13046
rect 4760 12990 4788 13046
rect 4844 12990 4872 13046
rect 4928 12990 4956 13046
rect 5012 12990 5040 13046
rect 5096 12990 5124 13046
rect 5180 12990 5208 13046
rect 5264 12990 5267 13046
rect 4701 12957 5267 12990
rect 4701 12901 4704 12957
rect 4760 12901 4788 12957
rect 4844 12901 4872 12957
rect 4928 12901 4956 12957
rect 5012 12901 5040 12957
rect 5096 12901 5124 12957
rect 5180 12901 5208 12957
rect 5264 12901 5267 12957
rect 4701 12868 5267 12901
rect 4701 12812 4704 12868
rect 4760 12812 4788 12868
rect 4844 12812 4872 12868
rect 4928 12812 4956 12868
rect 5012 12812 5040 12868
rect 5096 12812 5124 12868
rect 5180 12812 5208 12868
rect 5264 12812 5267 12868
rect 4701 12779 5267 12812
rect 4701 12723 4704 12779
rect 4760 12723 4788 12779
rect 4844 12723 4872 12779
rect 4928 12723 4956 12779
rect 5012 12723 5040 12779
rect 5096 12723 5124 12779
rect 5180 12723 5208 12779
rect 5264 12723 5267 12779
rect 4701 12690 5267 12723
rect 4701 12634 4704 12690
rect 4760 12634 4788 12690
rect 4844 12634 4872 12690
rect 4928 12634 4956 12690
rect 5012 12634 5040 12690
rect 5096 12634 5124 12690
rect 5180 12634 5208 12690
rect 5264 12634 5267 12690
rect 4701 12601 5267 12634
rect 4701 12545 4704 12601
rect 4760 12545 4788 12601
rect 4844 12545 4872 12601
rect 4928 12545 4956 12601
rect 5012 12545 5040 12601
rect 5096 12545 5124 12601
rect 5180 12545 5208 12601
rect 5264 12545 5267 12601
rect 4701 12511 5267 12545
rect 2903 12446 3469 12455
tri 4667 12446 4701 12480 ne
rect 4701 12455 4704 12511
rect 4760 12455 4788 12511
rect 4844 12455 4872 12511
rect 4928 12455 4956 12511
rect 5012 12455 5040 12511
rect 5096 12455 5124 12511
rect 5180 12455 5208 12511
rect 5264 12455 5267 12511
rect 6508 13046 7074 13055
rect 6508 12990 6511 13046
rect 6567 12990 6595 13046
rect 6651 12990 6679 13046
rect 6735 12990 6763 13046
rect 6819 12990 6847 13046
rect 6903 12990 6931 13046
rect 6987 12990 7015 13046
rect 7071 12990 7074 13046
rect 6508 12957 7074 12990
rect 6508 12901 6511 12957
rect 6567 12901 6595 12957
rect 6651 12901 6679 12957
rect 6735 12901 6763 12957
rect 6819 12901 6847 12957
rect 6903 12901 6931 12957
rect 6987 12901 7015 12957
rect 7071 12901 7074 12957
rect 6508 12868 7074 12901
rect 6508 12812 6511 12868
rect 6567 12812 6595 12868
rect 6651 12812 6679 12868
rect 6735 12812 6763 12868
rect 6819 12812 6847 12868
rect 6903 12812 6931 12868
rect 6987 12812 7015 12868
rect 7071 12812 7074 12868
rect 6508 12779 7074 12812
rect 6508 12723 6511 12779
rect 6567 12723 6595 12779
rect 6651 12723 6679 12779
rect 6735 12723 6763 12779
rect 6819 12723 6847 12779
rect 6903 12723 6931 12779
rect 6987 12723 7015 12779
rect 7071 12723 7074 12779
rect 6508 12690 7074 12723
rect 6508 12634 6511 12690
rect 6567 12634 6595 12690
rect 6651 12634 6679 12690
rect 6735 12634 6763 12690
rect 6819 12634 6847 12690
rect 6903 12634 6931 12690
rect 6987 12634 7015 12690
rect 7071 12634 7074 12690
rect 6508 12601 7074 12634
rect 6508 12545 6511 12601
rect 6567 12545 6595 12601
rect 6651 12545 6679 12601
rect 6735 12545 6763 12601
rect 6819 12545 6847 12601
rect 6903 12545 6931 12601
rect 6987 12545 7015 12601
rect 7071 12545 7074 12601
rect 6508 12511 7074 12545
rect 4701 12446 5267 12455
tri 5267 12446 5301 12480 nw
tri 6474 12446 6508 12480 ne
rect 6508 12455 6511 12511
rect 6567 12455 6595 12511
rect 6651 12455 6679 12511
rect 6735 12455 6763 12511
rect 6819 12455 6847 12511
rect 6903 12455 6931 12511
rect 6987 12455 7015 12511
rect 7071 12455 7074 12511
rect 8323 13045 8885 13054
rect 8323 12989 8324 13045
rect 8380 12989 8408 13045
rect 8464 12989 8492 13045
rect 8548 12989 8576 13045
rect 8632 12989 8660 13045
rect 8716 12989 8744 13045
rect 8800 12989 8828 13045
rect 8884 12989 8885 13045
rect 8323 12965 8885 12989
rect 8323 12909 8324 12965
rect 8380 12909 8408 12965
rect 8464 12909 8492 12965
rect 8548 12909 8576 12965
rect 8632 12909 8660 12965
rect 8716 12909 8744 12965
rect 8800 12909 8828 12965
rect 8884 12909 8885 12965
rect 8323 12885 8885 12909
rect 8323 12829 8324 12885
rect 8380 12829 8408 12885
rect 8464 12829 8492 12885
rect 8548 12829 8576 12885
rect 8632 12829 8660 12885
rect 8716 12829 8744 12885
rect 8800 12829 8828 12885
rect 8884 12829 8885 12885
rect 8323 12805 8885 12829
rect 8323 12749 8324 12805
rect 8380 12749 8408 12805
rect 8464 12749 8492 12805
rect 8548 12749 8576 12805
rect 8632 12749 8660 12805
rect 8716 12749 8744 12805
rect 8800 12749 8828 12805
rect 8884 12749 8885 12805
rect 8323 12725 8885 12749
rect 8323 12669 8324 12725
rect 8380 12669 8408 12725
rect 8464 12669 8492 12725
rect 8548 12669 8576 12725
rect 8632 12669 8660 12725
rect 8716 12669 8744 12725
rect 8800 12669 8828 12725
rect 8884 12669 8885 12725
rect 8323 12645 8885 12669
rect 8323 12589 8324 12645
rect 8380 12589 8408 12645
rect 8464 12589 8492 12645
rect 8548 12589 8576 12645
rect 8632 12589 8660 12645
rect 8716 12589 8744 12645
rect 8800 12589 8828 12645
rect 8884 12589 8885 12645
rect 8323 12565 8885 12589
rect 8323 12509 8324 12565
rect 8380 12509 8408 12565
rect 8464 12509 8492 12565
rect 8548 12509 8576 12565
rect 8632 12509 8660 12565
rect 8716 12509 8744 12565
rect 8800 12509 8828 12565
rect 8884 12509 8885 12565
rect 8323 12485 8885 12509
rect 6508 12446 7074 12455
tri 7074 12446 7108 12480 nw
rect -724 12377 -714 12433
rect -658 12377 -626 12433
rect -570 12377 -538 12433
rect -482 12377 -450 12433
rect -394 12377 -362 12433
rect -306 12377 -274 12433
rect -218 12377 -186 12433
rect -130 12377 -122 12433
rect -724 12353 -122 12377
rect -724 12297 -714 12353
rect -658 12297 -626 12353
rect -570 12297 -538 12353
rect -482 12297 -450 12353
rect -394 12297 -362 12353
rect -306 12297 -274 12353
rect -218 12297 -186 12353
rect -130 12297 -122 12353
rect -724 12273 -122 12297
rect -724 12217 -714 12273
rect -658 12217 -626 12273
rect -570 12217 -538 12273
rect -482 12217 -450 12273
rect -394 12217 -362 12273
rect -306 12217 -274 12273
rect -218 12217 -186 12273
rect -130 12217 -122 12273
rect -724 12193 -122 12217
tri -4109 12177 -4105 12181 se
rect -4105 12177 -1939 12181
tri -4311 11975 -4109 12177 se
rect -4109 12168 -1939 12177
rect -4109 12112 -2511 12168
rect -2455 12112 -2405 12168
rect -2349 12112 -2299 12168
rect -2243 12112 -2193 12168
rect -2137 12112 -1939 12168
rect -4109 12085 -1939 12112
rect -4109 12029 -2511 12085
rect -2455 12029 -2405 12085
rect -2349 12029 -2299 12085
rect -2243 12029 -2193 12085
rect -2137 12029 -1939 12085
rect -4109 12001 -1939 12029
rect -4109 11975 -2511 12001
rect -4311 11945 -2511 11975
rect -2455 11945 -2405 12001
rect -2349 11945 -2299 12001
rect -2243 11945 -2193 12001
rect -2137 11945 -1939 12001
rect -4311 11917 -1939 11945
rect -4311 11861 -2511 11917
rect -2455 11861 -2405 11917
rect -2349 11861 -2299 11917
rect -2243 11861 -2193 11917
rect -2137 11861 -1939 11917
rect -4311 11833 -1939 11861
rect -4311 11777 -2511 11833
rect -2455 11777 -2405 11833
rect -2349 11777 -2299 11833
rect -2243 11777 -2193 11833
rect -2137 11777 -1939 11833
rect -4311 11749 -1939 11777
rect -4311 11693 -2511 11749
rect -2455 11693 -2405 11749
rect -2349 11693 -2299 11749
rect -2243 11693 -2193 11749
rect -2137 11693 -1939 11749
rect -4311 5139 -1939 11693
rect -3750 5027 -3657 5139
tri -3657 5027 -3545 5139 nw
tri -2726 5027 -2614 5139 ne
rect -2614 5027 -2051 5139
tri -2051 5027 -1939 5139 nw
rect -724 12137 -714 12193
rect -658 12137 -626 12193
rect -570 12137 -538 12193
rect -482 12137 -450 12193
rect -394 12137 -362 12193
rect -306 12137 -274 12193
rect -218 12137 -186 12193
rect -130 12137 -122 12193
rect -724 12113 -122 12137
rect 8323 12429 8324 12485
rect 8380 12429 8408 12485
rect 8464 12429 8492 12485
rect 8548 12429 8576 12485
rect 8632 12429 8660 12485
rect 8716 12429 8744 12485
rect 8800 12429 8828 12485
rect 8884 12429 8885 12485
rect 10119 13046 10685 13055
rect 10119 12990 10122 13046
rect 10178 12990 10206 13046
rect 10262 12990 10290 13046
rect 10346 12990 10374 13046
rect 10430 12990 10458 13046
rect 10514 12990 10542 13046
rect 10598 12990 10626 13046
rect 10682 12990 10685 13046
rect 10119 12957 10685 12990
rect 10119 12901 10122 12957
rect 10178 12901 10206 12957
rect 10262 12901 10290 12957
rect 10346 12901 10374 12957
rect 10430 12901 10458 12957
rect 10514 12901 10542 12957
rect 10598 12901 10626 12957
rect 10682 12901 10685 12957
rect 10119 12868 10685 12901
rect 10119 12812 10122 12868
rect 10178 12812 10206 12868
rect 10262 12812 10290 12868
rect 10346 12812 10374 12868
rect 10430 12812 10458 12868
rect 10514 12812 10542 12868
rect 10598 12812 10626 12868
rect 10682 12812 10685 12868
rect 10119 12779 10685 12812
rect 10119 12723 10122 12779
rect 10178 12723 10206 12779
rect 10262 12723 10290 12779
rect 10346 12723 10374 12779
rect 10430 12723 10458 12779
rect 10514 12723 10542 12779
rect 10598 12723 10626 12779
rect 10682 12723 10685 12779
rect 10119 12690 10685 12723
rect 10119 12634 10122 12690
rect 10178 12634 10206 12690
rect 10262 12634 10290 12690
rect 10346 12634 10374 12690
rect 10430 12634 10458 12690
rect 10514 12634 10542 12690
rect 10598 12634 10626 12690
rect 10682 12634 10685 12690
rect 10119 12601 10685 12634
rect 10119 12545 10122 12601
rect 10178 12545 10206 12601
rect 10262 12545 10290 12601
rect 10346 12545 10374 12601
rect 10430 12545 10458 12601
rect 10514 12545 10542 12601
rect 10598 12545 10626 12601
rect 10682 12545 10685 12601
rect 10119 12511 10685 12545
tri 10085 12446 10119 12480 ne
rect 10119 12455 10122 12511
rect 10178 12455 10206 12511
rect 10262 12455 10290 12511
rect 10346 12455 10374 12511
rect 10430 12455 10458 12511
rect 10514 12455 10542 12511
rect 10598 12455 10626 12511
rect 10682 12455 10685 12511
rect 11920 13046 12486 13055
rect 11920 12990 11923 13046
rect 11979 12990 12007 13046
rect 12063 12990 12091 13046
rect 12147 12990 12175 13046
rect 12231 12990 12259 13046
rect 12315 12990 12343 13046
rect 12399 12990 12427 13046
rect 12483 12990 12486 13046
rect 11920 12963 12486 12990
rect 11920 12907 11923 12963
rect 11979 12907 12007 12963
rect 12063 12907 12091 12963
rect 12147 12907 12175 12963
rect 12231 12907 12259 12963
rect 12315 12907 12343 12963
rect 12399 12907 12427 12963
rect 12483 12907 12486 12963
rect 11920 12880 12486 12907
rect 11920 12824 11923 12880
rect 11979 12824 12007 12880
rect 12063 12824 12091 12880
rect 12147 12824 12175 12880
rect 12231 12824 12259 12880
rect 12315 12824 12343 12880
rect 12399 12824 12427 12880
rect 12483 12824 12486 12880
rect 11920 12797 12486 12824
rect 11920 12741 11923 12797
rect 11979 12741 12007 12797
rect 12063 12741 12091 12797
rect 12147 12741 12175 12797
rect 12231 12741 12259 12797
rect 12315 12741 12343 12797
rect 12399 12741 12427 12797
rect 12483 12741 12486 12797
rect 11920 12713 12486 12741
rect 11920 12657 11923 12713
rect 11979 12657 12007 12713
rect 12063 12657 12091 12713
rect 12147 12657 12175 12713
rect 12231 12657 12259 12713
rect 12315 12657 12343 12713
rect 12399 12657 12427 12713
rect 12483 12657 12486 12713
rect 11920 12629 12486 12657
rect 11920 12573 11923 12629
rect 11979 12573 12007 12629
rect 12063 12573 12091 12629
rect 12147 12573 12175 12629
rect 12231 12573 12259 12629
rect 12315 12573 12343 12629
rect 12399 12573 12427 12629
rect 12483 12573 12486 12629
rect 11920 12545 12486 12573
rect 11920 12489 11923 12545
rect 11979 12489 12007 12545
rect 12063 12489 12091 12545
rect 12147 12489 12175 12545
rect 12231 12489 12259 12545
rect 12315 12489 12343 12545
rect 12399 12489 12427 12545
rect 12483 12489 12486 12545
rect 11920 12480 12486 12489
rect 10119 12446 10685 12455
tri 10685 12446 10719 12480 nw
rect 8323 12405 8885 12429
rect 8323 12349 8324 12405
rect 8380 12349 8408 12405
rect 8464 12349 8492 12405
rect 8548 12349 8576 12405
rect 8632 12349 8660 12405
rect 8716 12349 8744 12405
rect 8800 12349 8828 12405
rect 8884 12349 8885 12405
rect 8323 12325 8885 12349
rect 8323 12269 8324 12325
rect 8380 12269 8408 12325
rect 8464 12269 8492 12325
rect 8548 12269 8576 12325
rect 8632 12269 8660 12325
rect 8716 12269 8744 12325
rect 8800 12269 8828 12325
rect 8884 12269 8885 12325
rect 8323 12245 8885 12269
rect 8323 12189 8324 12245
rect 8380 12189 8408 12245
rect 8464 12189 8492 12245
rect 8548 12189 8576 12245
rect 8632 12189 8660 12245
rect 8716 12189 8744 12245
rect 8800 12189 8828 12245
rect 8884 12189 8885 12245
rect 8323 12165 8885 12189
rect -724 12057 -714 12113
rect -658 12057 -626 12113
rect -570 12057 -538 12113
rect -482 12057 -450 12113
rect -394 12057 -362 12113
rect -306 12057 -274 12113
rect -218 12057 -186 12113
rect -130 12057 -122 12113
rect -724 12033 -122 12057
rect -724 11977 -714 12033
rect -658 11977 -626 12033
rect -570 11977 -538 12033
rect -482 11977 -450 12033
rect -394 11977 -362 12033
rect -306 11977 -274 12033
rect -218 11977 -186 12033
rect -130 11977 -122 12033
rect -724 11953 -122 11977
rect -724 11897 -714 11953
rect -658 11897 -626 11953
rect -570 11897 -538 11953
rect -482 11897 -450 11953
rect -394 11897 -362 11953
rect -306 11897 -274 11953
rect -218 11897 -186 11953
rect -130 11897 -122 11953
rect -724 11873 -122 11897
rect -724 11817 -714 11873
rect -658 11817 -626 11873
rect -570 11817 -538 11873
rect -482 11817 -450 11873
rect -394 11817 -362 11873
rect -306 11817 -274 11873
rect -218 11817 -186 11873
rect -130 11817 -122 11873
rect -724 11793 -122 11817
rect -724 11737 -714 11793
rect -658 11737 -626 11793
rect -570 11737 -538 11793
rect -482 11737 -450 11793
rect -394 11737 -362 11793
rect -306 11737 -274 11793
rect -218 11737 -186 11793
rect -130 11737 -122 11793
rect -724 11713 -122 11737
rect -724 11657 -714 11713
rect -658 11657 -626 11713
rect -570 11657 -538 11713
rect -482 11657 -450 11713
rect -394 11657 -362 11713
rect -306 11657 -274 11713
rect -218 11657 -186 11713
rect -130 11657 -122 11713
rect -724 11633 -122 11657
rect -724 11577 -714 11633
rect -658 11577 -626 11633
rect -570 11577 -538 11633
rect -482 11577 -450 11633
rect -394 11577 -362 11633
rect -306 11577 -274 11633
rect -218 11577 -186 11633
rect -130 11577 -122 11633
rect -724 11553 -122 11577
rect -724 11497 -714 11553
rect -658 11497 -626 11553
rect -570 11497 -538 11553
rect -482 11497 -450 11553
rect -394 11497 -362 11553
rect -306 11497 -274 11553
rect -218 11497 -186 11553
rect -130 11497 -122 11553
rect -724 11473 -122 11497
rect -724 11417 -714 11473
rect -658 11417 -626 11473
rect -570 11417 -538 11473
rect -482 11417 -450 11473
rect -394 11417 -362 11473
rect -306 11417 -274 11473
rect -218 11417 -186 11473
rect -130 11417 -122 11473
rect -724 11393 -122 11417
rect -724 11337 -714 11393
rect -658 11337 -626 11393
rect -570 11337 -538 11393
rect -482 11337 -450 11393
rect -394 11337 -362 11393
rect -306 11337 -274 11393
rect -218 11337 -186 11393
rect -130 11337 -122 11393
rect -724 11313 -122 11337
rect -724 11257 -714 11313
rect -658 11257 -626 11313
rect -570 11257 -538 11313
rect -482 11257 -450 11313
rect -394 11257 -362 11313
rect -306 11257 -274 11313
rect -218 11257 -186 11313
rect -130 11257 -122 11313
rect -724 11233 -122 11257
rect -724 11177 -714 11233
rect -658 11177 -626 11233
rect -570 11177 -538 11233
rect -482 11177 -450 11233
rect -394 11177 -362 11233
rect -306 11177 -274 11233
rect -218 11177 -186 11233
rect -130 11177 -122 11233
rect -724 11153 -122 11177
rect -724 11097 -714 11153
rect -658 11097 -626 11153
rect -570 11097 -538 11153
rect -482 11097 -450 11153
rect -394 11097 -362 11153
rect -306 11097 -274 11153
rect -218 11097 -186 11153
rect -130 11097 -122 11153
rect -724 11073 -122 11097
rect -724 11017 -714 11073
rect -658 11017 -626 11073
rect -570 11017 -538 11073
rect -482 11017 -450 11073
rect -394 11017 -362 11073
rect -306 11017 -274 11073
rect -218 11017 -186 11073
rect -130 11017 -122 11073
rect -724 10993 -122 11017
rect -724 10937 -714 10993
rect -658 10937 -626 10993
rect -570 10937 -538 10993
rect -482 10937 -450 10993
rect -394 10937 -362 10993
rect -306 10937 -274 10993
rect -218 10937 -186 10993
rect -130 10937 -122 10993
rect -724 10913 -122 10937
rect -724 10857 -714 10913
rect -658 10857 -626 10913
rect -570 10857 -538 10913
rect -482 10857 -450 10913
rect -394 10857 -362 10913
rect -306 10857 -274 10913
rect -218 10857 -186 10913
rect -130 10857 -122 10913
rect -724 10833 -122 10857
rect -724 10777 -714 10833
rect -658 10777 -626 10833
rect -570 10777 -538 10833
rect -482 10777 -450 10833
rect -394 10777 -362 10833
rect -306 10777 -274 10833
rect -218 10777 -186 10833
rect -130 10777 -122 10833
rect -724 10753 -122 10777
rect -724 10697 -714 10753
rect -658 10697 -626 10753
rect -570 10697 -538 10753
rect -482 10697 -450 10753
rect -394 10697 -362 10753
rect -306 10697 -274 10753
rect -218 10697 -186 10753
rect -130 10697 -122 10753
rect -724 10673 -122 10697
rect -724 10617 -714 10673
rect -658 10617 -626 10673
rect -570 10617 -538 10673
rect -482 10617 -450 10673
rect -394 10617 -362 10673
rect -306 10617 -274 10673
rect -218 10617 -186 10673
rect -130 10617 -122 10673
rect -724 10593 -122 10617
rect -724 10537 -714 10593
rect -658 10537 -626 10593
rect -570 10537 -538 10593
rect -482 10537 -450 10593
rect -394 10537 -362 10593
rect -306 10537 -274 10593
rect -218 10537 -186 10593
rect -130 10537 -122 10593
rect -724 10513 -122 10537
rect -724 10457 -714 10513
rect -658 10457 -626 10513
rect -570 10457 -538 10513
rect -482 10457 -450 10513
rect -394 10457 -362 10513
rect -306 10457 -274 10513
rect -218 10457 -186 10513
rect -130 10457 -122 10513
rect -724 10433 -122 10457
rect -724 10377 -714 10433
rect -658 10377 -626 10433
rect -570 10377 -538 10433
rect -482 10377 -450 10433
rect -394 10377 -362 10433
rect -306 10377 -274 10433
rect -218 10377 -186 10433
rect -130 10377 -122 10433
rect -724 10353 -122 10377
rect -724 10297 -714 10353
rect -658 10297 -626 10353
rect -570 10297 -538 10353
rect -482 10297 -450 10353
rect -394 10297 -362 10353
rect -306 10297 -274 10353
rect -218 10297 -186 10353
rect -130 10297 -122 10353
rect -724 10273 -122 10297
rect -724 10217 -714 10273
rect -658 10217 -626 10273
rect -570 10217 -538 10273
rect -482 10217 -450 10273
rect -394 10217 -362 10273
rect -306 10217 -274 10273
rect -218 10217 -186 10273
rect -130 10217 -122 10273
rect -724 10193 -122 10217
rect -724 10137 -714 10193
rect -658 10137 -626 10193
rect -570 10137 -538 10193
rect -482 10137 -450 10193
rect -394 10137 -362 10193
rect -306 10137 -274 10193
rect -218 10137 -186 10193
rect -130 10137 -122 10193
rect -724 10113 -122 10137
rect -724 10057 -714 10113
rect -658 10057 -626 10113
rect -570 10057 -538 10113
rect -482 10057 -450 10113
rect -394 10057 -362 10113
rect -306 10057 -274 10113
rect -218 10057 -186 10113
rect -130 10057 -122 10113
rect -724 10033 -122 10057
rect -724 9977 -714 10033
rect -658 9977 -626 10033
rect -570 9977 -538 10033
rect -482 9977 -450 10033
rect -394 9977 -362 10033
rect -306 9977 -274 10033
rect -218 9977 -186 10033
rect -130 9977 -122 10033
rect -724 9953 -122 9977
rect -724 9897 -714 9953
rect -658 9897 -626 9953
rect -570 9897 -538 9953
rect -482 9897 -450 9953
rect -394 9897 -362 9953
rect -306 9897 -274 9953
rect -218 9897 -186 9953
rect -130 9897 -122 9953
rect -724 9873 -122 9897
rect -724 9817 -714 9873
rect -658 9817 -626 9873
rect -570 9817 -538 9873
rect -482 9817 -450 9873
rect -394 9817 -362 9873
rect -306 9817 -274 9873
rect -218 9817 -186 9873
rect -130 9817 -122 9873
rect -724 9793 -122 9817
rect -724 9737 -714 9793
rect -658 9737 -626 9793
rect -570 9737 -538 9793
rect -482 9737 -450 9793
rect -394 9737 -362 9793
rect -306 9737 -274 9793
rect -218 9737 -186 9793
rect -130 9737 -122 9793
rect -724 9713 -122 9737
rect -724 9657 -714 9713
rect -658 9657 -626 9713
rect -570 9657 -538 9713
rect -482 9657 -450 9713
rect -394 9657 -362 9713
rect -306 9657 -274 9713
rect -218 9657 -186 9713
rect -130 9657 -122 9713
rect -724 9633 -122 9657
rect -724 9577 -714 9633
rect -658 9577 -626 9633
rect -570 9577 -538 9633
rect -482 9577 -450 9633
rect -394 9577 -362 9633
rect -306 9577 -274 9633
rect -218 9577 -186 9633
rect -130 9577 -122 9633
rect -724 9553 -122 9577
rect -724 9497 -714 9553
rect -658 9497 -626 9553
rect -570 9497 -538 9553
rect -482 9497 -450 9553
rect -394 9497 -362 9553
rect -306 9497 -274 9553
rect -218 9497 -186 9553
rect -130 9497 -122 9553
rect -724 9473 -122 9497
rect -724 9417 -714 9473
rect -658 9417 -626 9473
rect -570 9417 -538 9473
rect -482 9417 -450 9473
rect -394 9417 -362 9473
rect -306 9417 -274 9473
rect -218 9417 -186 9473
rect -130 9417 -122 9473
rect -724 9393 -122 9417
rect -724 9337 -714 9393
rect -658 9337 -626 9393
rect -570 9337 -538 9393
rect -482 9337 -450 9393
rect -394 9337 -362 9393
rect -306 9337 -274 9393
rect -218 9337 -186 9393
rect -130 9337 -122 9393
rect -724 9313 -122 9337
rect -724 9257 -714 9313
rect -658 9257 -626 9313
rect -570 9257 -538 9313
rect -482 9257 -450 9313
rect -394 9257 -362 9313
rect -306 9257 -274 9313
rect -218 9257 -186 9313
rect -130 9257 -122 9313
rect -724 9233 -122 9257
rect -724 9177 -714 9233
rect -658 9177 -626 9233
rect -570 9177 -538 9233
rect -482 9177 -450 9233
rect -394 9177 -362 9233
rect -306 9177 -274 9233
rect -218 9177 -186 9233
rect -130 9177 -122 9233
rect -724 9153 -122 9177
rect -724 9097 -714 9153
rect -658 9097 -626 9153
rect -570 9097 -538 9153
rect -482 9097 -450 9153
rect -394 9097 -362 9153
rect -306 9097 -274 9153
rect -218 9097 -186 9153
rect -130 9097 -122 9153
rect -724 9073 -122 9097
rect -724 9017 -714 9073
rect -658 9017 -626 9073
rect -570 9017 -538 9073
rect -482 9017 -450 9073
rect -394 9017 -362 9073
rect -306 9017 -274 9073
rect -218 9017 -186 9073
rect -130 9017 -122 9073
rect -724 8993 -122 9017
rect -724 8937 -714 8993
rect -658 8937 -626 8993
rect -570 8937 -538 8993
rect -482 8937 -450 8993
rect -394 8937 -362 8993
rect -306 8937 -274 8993
rect -218 8937 -186 8993
rect -130 8937 -122 8993
rect -724 8913 -122 8937
rect -724 8857 -714 8913
rect -658 8857 -626 8913
rect -570 8857 -538 8913
rect -482 8857 -450 8913
rect -394 8857 -362 8913
rect -306 8857 -274 8913
rect -218 8857 -186 8913
rect -130 8857 -122 8913
rect -724 8833 -122 8857
rect -724 8777 -714 8833
rect -658 8777 -626 8833
rect -570 8777 -538 8833
rect -482 8777 -450 8833
rect -394 8777 -362 8833
rect -306 8777 -274 8833
rect -218 8777 -186 8833
rect -130 8777 -122 8833
rect -724 8753 -122 8777
rect -724 8697 -714 8753
rect -658 8697 -626 8753
rect -570 8697 -538 8753
rect -482 8697 -450 8753
rect -394 8697 -362 8753
rect -306 8697 -274 8753
rect -218 8697 -186 8753
rect -130 8697 -122 8753
rect -724 8673 -122 8697
rect -724 8617 -714 8673
rect -658 8617 -626 8673
rect -570 8617 -538 8673
rect -482 8617 -450 8673
rect -394 8617 -362 8673
rect -306 8617 -274 8673
rect -218 8617 -186 8673
rect -130 8617 -122 8673
rect -724 8593 -122 8617
rect -724 8537 -714 8593
rect -658 8537 -626 8593
rect -570 8537 -538 8593
rect -482 8537 -450 8593
rect -394 8537 -362 8593
rect -306 8537 -274 8593
rect -218 8537 -186 8593
rect -130 8537 -122 8593
rect -724 8513 -122 8537
rect -724 8457 -714 8513
rect -658 8457 -626 8513
rect -570 8457 -538 8513
rect -482 8457 -450 8513
rect -394 8457 -362 8513
rect -306 8457 -274 8513
rect -218 8457 -186 8513
rect -130 8457 -122 8513
rect -724 8433 -122 8457
rect -724 8377 -714 8433
rect -658 8377 -626 8433
rect -570 8377 -538 8433
rect -482 8377 -450 8433
rect -394 8377 -362 8433
rect -306 8377 -274 8433
rect -218 8377 -186 8433
rect -130 8377 -122 8433
rect -724 8353 -122 8377
rect -724 8297 -714 8353
rect -658 8297 -626 8353
rect -570 8297 -538 8353
rect -482 8297 -450 8353
rect -394 8297 -362 8353
rect -306 8297 -274 8353
rect -218 8297 -186 8353
rect -130 8297 -122 8353
rect -724 8273 -122 8297
rect -724 8217 -714 8273
rect -658 8217 -626 8273
rect -570 8217 -538 8273
rect -482 8217 -450 8273
rect -394 8217 -362 8273
rect -306 8217 -274 8273
rect -218 8217 -186 8273
rect -130 8217 -122 8273
rect -724 8193 -122 8217
rect -724 8137 -714 8193
rect -658 8137 -626 8193
rect -570 8137 -538 8193
rect -482 8137 -450 8193
rect -394 8137 -362 8193
rect -306 8137 -274 8193
rect -218 8137 -186 8193
rect -130 8137 -122 8193
rect -724 8113 -122 8137
rect -724 8057 -714 8113
rect -658 8057 -626 8113
rect -570 8057 -538 8113
rect -482 8057 -450 8113
rect -394 8057 -362 8113
rect -306 8057 -274 8113
rect -218 8057 -186 8113
rect -130 8057 -122 8113
rect -724 8033 -122 8057
rect -724 7977 -714 8033
rect -658 7977 -626 8033
rect -570 7977 -538 8033
rect -482 7977 -450 8033
rect -394 7977 -362 8033
rect -306 7977 -274 8033
rect -218 7977 -186 8033
rect -130 7977 -122 8033
rect -724 7953 -122 7977
rect -724 7897 -714 7953
rect -658 7897 -626 7953
rect -570 7897 -538 7953
rect -482 7897 -450 7953
rect -394 7897 -362 7953
rect -306 7897 -274 7953
rect -218 7897 -186 7953
rect -130 7897 -122 7953
rect -724 7873 -122 7897
rect -724 7817 -714 7873
rect -658 7817 -626 7873
rect -570 7817 -538 7873
rect -482 7817 -450 7873
rect -394 7817 -362 7873
rect -306 7817 -274 7873
rect -218 7817 -186 7873
rect -130 7817 -122 7873
rect -724 7793 -122 7817
rect -724 7737 -714 7793
rect -658 7737 -626 7793
rect -570 7737 -538 7793
rect -482 7737 -450 7793
rect -394 7737 -362 7793
rect -306 7737 -274 7793
rect -218 7737 -186 7793
rect -130 7737 -122 7793
rect -724 7713 -122 7737
rect -724 7657 -714 7713
rect -658 7657 -626 7713
rect -570 7657 -538 7713
rect -482 7657 -450 7713
rect -394 7657 -362 7713
rect -306 7657 -274 7713
rect -218 7657 -186 7713
rect -130 7657 -122 7713
rect -724 7633 -122 7657
rect -724 7577 -714 7633
rect -658 7577 -626 7633
rect -570 7577 -538 7633
rect -482 7577 -450 7633
rect -394 7577 -362 7633
rect -306 7577 -274 7633
rect -218 7577 -186 7633
rect -130 7577 -122 7633
rect -724 7553 -122 7577
rect -724 7497 -714 7553
rect -658 7497 -626 7553
rect -570 7497 -538 7553
rect -482 7497 -450 7553
rect -394 7497 -362 7553
rect -306 7497 -274 7553
rect -218 7497 -186 7553
rect -130 7497 -122 7553
rect -724 7473 -122 7497
rect -724 7417 -714 7473
rect -658 7417 -626 7473
rect -570 7417 -538 7473
rect -482 7417 -450 7473
rect -394 7417 -362 7473
rect -306 7417 -274 7473
rect -218 7417 -186 7473
rect -130 7417 -122 7473
rect -724 7393 -122 7417
rect -724 7337 -714 7393
rect -658 7337 -626 7393
rect -570 7337 -538 7393
rect -482 7337 -450 7393
rect -394 7337 -362 7393
rect -306 7337 -274 7393
rect -218 7337 -186 7393
rect -130 7337 -122 7393
rect -724 7313 -122 7337
rect -724 7257 -714 7313
rect -658 7257 -626 7313
rect -570 7257 -538 7313
rect -482 7257 -450 7313
rect -394 7257 -362 7313
rect -306 7257 -274 7313
rect -218 7257 -186 7313
rect -130 7257 -122 7313
rect -724 7233 -122 7257
rect -724 7177 -714 7233
rect -658 7177 -626 7233
rect -570 7177 -538 7233
rect -482 7177 -450 7233
rect -394 7177 -362 7233
rect -306 7177 -274 7233
rect -218 7177 -186 7233
rect -130 7177 -122 7233
rect -724 7153 -122 7177
rect -724 7097 -714 7153
rect -658 7097 -626 7153
rect -570 7097 -538 7153
rect -482 7097 -450 7153
rect -394 7097 -362 7153
rect -306 7097 -274 7153
rect -218 7097 -186 7153
rect -130 7097 -122 7153
rect -724 7073 -122 7097
rect -724 7017 -714 7073
rect -658 7017 -626 7073
rect -570 7017 -538 7073
rect -482 7017 -450 7073
rect -394 7017 -362 7073
rect -306 7017 -274 7073
rect -218 7017 -186 7073
rect -130 7017 -122 7073
rect -724 6993 -122 7017
rect -724 6937 -714 6993
rect -658 6937 -626 6993
rect -570 6937 -538 6993
rect -482 6937 -450 6993
rect -394 6937 -362 6993
rect -306 6937 -274 6993
rect -218 6937 -186 6993
rect -130 6937 -122 6993
rect -724 6912 -122 6937
rect -724 6856 -714 6912
rect -658 6856 -626 6912
rect -570 6856 -538 6912
rect -482 6856 -450 6912
rect -394 6856 -362 6912
rect -306 6856 -274 6912
rect -218 6856 -186 6912
rect -130 6856 -122 6912
rect -724 6831 -122 6856
rect -724 6775 -714 6831
rect -658 6775 -626 6831
rect -570 6775 -538 6831
rect -482 6775 -450 6831
rect -394 6775 -362 6831
rect -306 6775 -274 6831
rect -218 6775 -186 6831
rect -130 6775 -122 6831
rect -724 6750 -122 6775
rect -724 6694 -714 6750
rect -658 6694 -626 6750
rect -570 6694 -538 6750
rect -482 6694 -450 6750
rect -394 6694 -362 6750
rect -306 6694 -274 6750
rect -218 6694 -186 6750
rect -130 6694 -122 6750
rect -724 6669 -122 6694
rect -724 6613 -714 6669
rect -658 6613 -626 6669
rect -570 6613 -538 6669
rect -482 6613 -450 6669
rect -394 6613 -362 6669
rect -306 6613 -274 6669
rect -218 6613 -186 6669
rect -130 6613 -122 6669
rect -724 6588 -122 6613
rect -724 6532 -714 6588
rect -658 6532 -626 6588
rect -570 6532 -538 6588
rect -482 6532 -450 6588
rect -394 6532 -362 6588
rect -306 6532 -274 6588
rect -218 6532 -186 6588
rect -130 6532 -122 6588
rect -724 6507 -122 6532
rect -724 6451 -714 6507
rect -658 6451 -626 6507
rect -570 6451 -538 6507
rect -482 6451 -450 6507
rect -394 6451 -362 6507
rect -306 6451 -274 6507
rect -218 6451 -186 6507
rect -130 6451 -122 6507
rect -724 6426 -122 6451
rect -724 6370 -714 6426
rect -658 6370 -626 6426
rect -570 6370 -538 6426
rect -482 6370 -450 6426
rect -394 6370 -362 6426
rect -306 6370 -274 6426
rect -218 6370 -186 6426
rect -130 6370 -122 6426
rect -724 6345 -122 6370
rect -724 6289 -714 6345
rect -658 6289 -626 6345
rect -570 6289 -538 6345
rect -482 6289 -450 6345
rect -394 6289 -362 6345
rect -306 6289 -274 6345
rect -218 6289 -186 6345
rect -130 6289 -122 6345
rect -724 6264 -122 6289
rect -724 6208 -714 6264
rect -658 6208 -626 6264
rect -570 6208 -538 6264
rect -482 6208 -450 6264
rect -394 6208 -362 6264
rect -306 6208 -274 6264
rect -218 6208 -186 6264
rect -130 6208 -122 6264
rect -724 6183 -122 6208
rect -724 6127 -714 6183
rect -658 6127 -626 6183
rect -570 6127 -538 6183
rect -482 6127 -450 6183
rect -394 6127 -362 6183
rect -306 6127 -274 6183
rect -218 6127 -186 6183
rect -130 6127 -122 6183
rect -724 6102 -122 6127
rect -724 6046 -714 6102
rect -658 6046 -626 6102
rect -570 6046 -538 6102
rect -482 6046 -450 6102
rect -394 6046 -362 6102
rect -306 6046 -274 6102
rect -218 6046 -186 6102
rect -130 6046 -122 6102
rect -724 6021 -122 6046
rect -724 5965 -714 6021
rect -658 5965 -626 6021
rect -570 5965 -538 6021
rect -482 5965 -450 6021
rect -394 5965 -362 6021
rect -306 5965 -274 6021
rect -218 5965 -186 6021
rect -130 5965 -122 6021
rect -724 5940 -122 5965
rect -724 5884 -714 5940
rect -658 5884 -626 5940
rect -570 5884 -538 5940
rect -482 5884 -450 5940
rect -394 5884 -362 5940
rect -306 5884 -274 5940
rect -218 5884 -186 5940
rect -130 5884 -122 5940
rect -724 5859 -122 5884
rect -724 5803 -714 5859
rect -658 5803 -626 5859
rect -570 5803 -538 5859
rect -482 5803 -450 5859
rect -394 5803 -362 5859
rect -306 5803 -274 5859
rect -218 5803 -186 5859
rect -130 5803 -122 5859
rect -724 5778 -122 5803
rect -724 5722 -714 5778
rect -658 5722 -626 5778
rect -570 5722 -538 5778
rect -482 5722 -450 5778
rect -394 5722 -362 5778
rect -306 5722 -274 5778
rect -218 5722 -186 5778
rect -130 5722 -122 5778
rect -724 5697 -122 5722
rect -724 5641 -714 5697
rect -658 5641 -626 5697
rect -570 5641 -538 5697
rect -482 5641 -450 5697
rect -394 5641 -362 5697
rect -306 5641 -274 5697
rect -218 5641 -186 5697
rect -130 5641 -122 5697
rect -724 5616 -122 5641
rect -724 5560 -714 5616
rect -658 5560 -626 5616
rect -570 5560 -538 5616
rect -482 5560 -450 5616
rect -394 5560 -362 5616
rect -306 5560 -274 5616
rect -218 5560 -186 5616
rect -130 5560 -122 5616
rect -724 5535 -122 5560
rect -724 5479 -714 5535
rect -658 5479 -626 5535
rect -570 5479 -538 5535
rect -482 5479 -450 5535
rect -394 5479 -362 5535
rect -306 5479 -274 5535
rect -218 5479 -186 5535
rect -130 5479 -122 5535
rect -724 5454 -122 5479
rect -724 5398 -714 5454
rect -658 5398 -626 5454
rect -570 5398 -538 5454
rect -482 5398 -450 5454
rect -394 5398 -362 5454
rect -306 5398 -274 5454
rect -218 5398 -186 5454
rect -130 5398 -122 5454
rect -724 5373 -122 5398
rect -724 5317 -714 5373
rect -658 5317 -626 5373
rect -570 5317 -538 5373
rect -482 5317 -450 5373
rect -394 5317 -362 5373
rect -306 5317 -274 5373
rect -218 5317 -186 5373
rect -130 5317 -122 5373
rect -724 5292 -122 5317
rect -724 5236 -714 5292
rect -658 5236 -626 5292
rect -570 5236 -538 5292
rect -482 5236 -450 5292
rect -394 5236 -362 5292
rect -306 5236 -274 5292
rect -218 5236 -186 5292
rect -130 5236 -122 5292
rect -724 5211 -122 5236
rect -724 5155 -714 5211
rect -658 5155 -626 5211
rect -570 5155 -538 5211
rect -482 5155 -450 5211
rect -394 5155 -362 5211
rect -306 5155 -274 5211
rect -218 5155 -186 5211
rect -130 5155 -122 5211
rect 1094 5210 1670 12116
rect 2898 11335 3474 11680
rect 4699 5210 5275 12116
rect 6506 5210 7082 12116
rect 8323 12109 8324 12165
rect 8380 12109 8408 12165
rect 8464 12109 8492 12165
rect 8548 12109 8576 12165
rect 8632 12109 8660 12165
rect 8716 12109 8744 12165
rect 8800 12109 8828 12165
rect 8884 12109 8885 12165
rect 8323 12085 8885 12109
rect 8323 12029 8324 12085
rect 8380 12029 8408 12085
rect 8464 12029 8492 12085
rect 8548 12029 8576 12085
rect 8632 12029 8660 12085
rect 8716 12029 8744 12085
rect 8800 12029 8828 12085
rect 8884 12029 8885 12085
rect 8323 12005 8885 12029
rect 8323 11949 8324 12005
rect 8380 11949 8408 12005
rect 8464 11949 8492 12005
rect 8548 11949 8576 12005
rect 8632 11949 8660 12005
rect 8716 11949 8744 12005
rect 8800 11949 8828 12005
rect 8884 11949 8885 12005
rect 8323 11925 8885 11949
rect 8323 11869 8324 11925
rect 8380 11869 8408 11925
rect 8464 11869 8492 11925
rect 8548 11869 8576 11925
rect 8632 11869 8660 11925
rect 8716 11869 8744 11925
rect 8800 11869 8828 11925
rect 8884 11869 8885 11925
rect 8323 11845 8885 11869
rect 8323 11789 8324 11845
rect 8380 11789 8408 11845
rect 8464 11789 8492 11845
rect 8548 11789 8576 11845
rect 8632 11789 8660 11845
rect 8716 11789 8744 11845
rect 8800 11789 8828 11845
rect 8884 11789 8885 11845
rect 8323 11765 8885 11789
rect 8323 11709 8324 11765
rect 8380 11709 8408 11765
rect 8464 11709 8492 11765
rect 8548 11709 8576 11765
rect 8632 11709 8660 11765
rect 8716 11709 8744 11765
rect 8800 11709 8828 11765
rect 8884 11709 8885 11765
rect 8323 11685 8885 11709
rect 8323 11629 8324 11685
rect 8380 11629 8408 11685
rect 8464 11629 8492 11685
rect 8548 11629 8576 11685
rect 8632 11629 8660 11685
rect 8716 11629 8744 11685
rect 8800 11629 8828 11685
rect 8884 11629 8885 11685
rect 8323 11605 8885 11629
rect 8323 11549 8324 11605
rect 8380 11549 8408 11605
rect 8464 11549 8492 11605
rect 8548 11549 8576 11605
rect 8632 11549 8660 11605
rect 8716 11549 8744 11605
rect 8800 11549 8828 11605
rect 8884 11549 8885 11605
rect 8323 11525 8885 11549
rect 8323 11469 8324 11525
rect 8380 11469 8408 11525
rect 8464 11469 8492 11525
rect 8548 11469 8576 11525
rect 8632 11469 8660 11525
rect 8716 11469 8744 11525
rect 8800 11469 8828 11525
rect 8884 11469 8885 11525
rect 8323 11445 8885 11469
rect 8323 11389 8324 11445
rect 8380 11389 8408 11445
rect 8464 11389 8492 11445
rect 8548 11389 8576 11445
rect 8632 11389 8660 11445
rect 8716 11389 8744 11445
rect 8800 11389 8828 11445
rect 8884 11389 8885 11445
rect 8323 11365 8885 11389
rect 8323 11309 8324 11365
rect 8380 11309 8408 11365
rect 8464 11309 8492 11365
rect 8548 11309 8576 11365
rect 8632 11309 8660 11365
rect 8716 11309 8744 11365
rect 8800 11309 8828 11365
rect 8884 11309 8885 11365
rect 8323 11285 8885 11309
rect 8323 11229 8324 11285
rect 8380 11229 8408 11285
rect 8464 11229 8492 11285
rect 8548 11229 8576 11285
rect 8632 11229 8660 11285
rect 8716 11229 8744 11285
rect 8800 11229 8828 11285
rect 8884 11229 8885 11285
rect 8323 11205 8885 11229
rect 8323 11149 8324 11205
rect 8380 11149 8408 11205
rect 8464 11149 8492 11205
rect 8548 11149 8576 11205
rect 8632 11149 8660 11205
rect 8716 11149 8744 11205
rect 8800 11149 8828 11205
rect 8884 11149 8885 11205
rect 8323 11125 8885 11149
rect 8323 11069 8324 11125
rect 8380 11069 8408 11125
rect 8464 11069 8492 11125
rect 8548 11069 8576 11125
rect 8632 11069 8660 11125
rect 8716 11069 8744 11125
rect 8800 11069 8828 11125
rect 8884 11069 8885 11125
rect 8323 11045 8885 11069
rect 8323 10989 8324 11045
rect 8380 10989 8408 11045
rect 8464 10989 8492 11045
rect 8548 10989 8576 11045
rect 8632 10989 8660 11045
rect 8716 10989 8744 11045
rect 8800 10989 8828 11045
rect 8884 10989 8885 11045
rect 8323 10965 8885 10989
rect 8323 10909 8324 10965
rect 8380 10909 8408 10965
rect 8464 10909 8492 10965
rect 8548 10909 8576 10965
rect 8632 10909 8660 10965
rect 8716 10909 8744 10965
rect 8800 10909 8828 10965
rect 8884 10909 8885 10965
rect 8323 10885 8885 10909
rect 8323 10829 8324 10885
rect 8380 10829 8408 10885
rect 8464 10829 8492 10885
rect 8548 10829 8576 10885
rect 8632 10829 8660 10885
rect 8716 10829 8744 10885
rect 8800 10829 8828 10885
rect 8884 10829 8885 10885
rect 8323 10805 8885 10829
rect 8323 10749 8324 10805
rect 8380 10749 8408 10805
rect 8464 10749 8492 10805
rect 8548 10749 8576 10805
rect 8632 10749 8660 10805
rect 8716 10749 8744 10805
rect 8800 10749 8828 10805
rect 8884 10749 8885 10805
rect 8323 10725 8885 10749
rect 8323 10669 8324 10725
rect 8380 10669 8408 10725
rect 8464 10669 8492 10725
rect 8548 10669 8576 10725
rect 8632 10669 8660 10725
rect 8716 10669 8744 10725
rect 8800 10669 8828 10725
rect 8884 10669 8885 10725
rect 8323 10645 8885 10669
rect 8323 10589 8324 10645
rect 8380 10589 8408 10645
rect 8464 10589 8492 10645
rect 8548 10589 8576 10645
rect 8632 10589 8660 10645
rect 8716 10589 8744 10645
rect 8800 10589 8828 10645
rect 8884 10589 8885 10645
rect 8323 10565 8885 10589
rect 8323 10509 8324 10565
rect 8380 10509 8408 10565
rect 8464 10509 8492 10565
rect 8548 10509 8576 10565
rect 8632 10509 8660 10565
rect 8716 10509 8744 10565
rect 8800 10509 8828 10565
rect 8884 10509 8885 10565
rect 8323 10485 8885 10509
rect 8323 10429 8324 10485
rect 8380 10429 8408 10485
rect 8464 10429 8492 10485
rect 8548 10429 8576 10485
rect 8632 10429 8660 10485
rect 8716 10429 8744 10485
rect 8800 10429 8828 10485
rect 8884 10429 8885 10485
rect 8323 10405 8885 10429
rect 8323 10349 8324 10405
rect 8380 10349 8408 10405
rect 8464 10349 8492 10405
rect 8548 10349 8576 10405
rect 8632 10349 8660 10405
rect 8716 10349 8744 10405
rect 8800 10349 8828 10405
rect 8884 10349 8885 10405
rect 8323 10325 8885 10349
rect 8323 10269 8324 10325
rect 8380 10269 8408 10325
rect 8464 10269 8492 10325
rect 8548 10269 8576 10325
rect 8632 10269 8660 10325
rect 8716 10269 8744 10325
rect 8800 10269 8828 10325
rect 8884 10269 8885 10325
rect 8323 10245 8885 10269
rect 8323 10189 8324 10245
rect 8380 10189 8408 10245
rect 8464 10189 8492 10245
rect 8548 10189 8576 10245
rect 8632 10189 8660 10245
rect 8716 10189 8744 10245
rect 8800 10189 8828 10245
rect 8884 10189 8885 10245
rect 8323 10165 8885 10189
rect 8323 10109 8324 10165
rect 8380 10109 8408 10165
rect 8464 10109 8492 10165
rect 8548 10109 8576 10165
rect 8632 10109 8660 10165
rect 8716 10109 8744 10165
rect 8800 10109 8828 10165
rect 8884 10109 8885 10165
rect 8323 10085 8885 10109
rect 8323 10029 8324 10085
rect 8380 10029 8408 10085
rect 8464 10029 8492 10085
rect 8548 10029 8576 10085
rect 8632 10029 8660 10085
rect 8716 10029 8744 10085
rect 8800 10029 8828 10085
rect 8884 10029 8885 10085
rect 8323 10005 8885 10029
rect 8323 9949 8324 10005
rect 8380 9949 8408 10005
rect 8464 9949 8492 10005
rect 8548 9949 8576 10005
rect 8632 9949 8660 10005
rect 8716 9949 8744 10005
rect 8800 9949 8828 10005
rect 8884 9949 8885 10005
rect 8323 9925 8885 9949
rect 8323 9869 8324 9925
rect 8380 9869 8408 9925
rect 8464 9869 8492 9925
rect 8548 9869 8576 9925
rect 8632 9869 8660 9925
rect 8716 9869 8744 9925
rect 8800 9869 8828 9925
rect 8884 9869 8885 9925
rect 8323 9845 8885 9869
rect 8323 9789 8324 9845
rect 8380 9789 8408 9845
rect 8464 9789 8492 9845
rect 8548 9789 8576 9845
rect 8632 9789 8660 9845
rect 8716 9789 8744 9845
rect 8800 9789 8828 9845
rect 8884 9789 8885 9845
rect 8323 9765 8885 9789
rect 8323 9709 8324 9765
rect 8380 9709 8408 9765
rect 8464 9709 8492 9765
rect 8548 9709 8576 9765
rect 8632 9709 8660 9765
rect 8716 9709 8744 9765
rect 8800 9709 8828 9765
rect 8884 9709 8885 9765
rect 8323 9685 8885 9709
rect 8323 9629 8324 9685
rect 8380 9629 8408 9685
rect 8464 9629 8492 9685
rect 8548 9629 8576 9685
rect 8632 9629 8660 9685
rect 8716 9629 8744 9685
rect 8800 9629 8828 9685
rect 8884 9629 8885 9685
rect 8323 9605 8885 9629
rect 8323 9549 8324 9605
rect 8380 9549 8408 9605
rect 8464 9549 8492 9605
rect 8548 9549 8576 9605
rect 8632 9549 8660 9605
rect 8716 9549 8744 9605
rect 8800 9549 8828 9605
rect 8884 9549 8885 9605
rect 8323 9524 8885 9549
rect 8323 9468 8324 9524
rect 8380 9468 8408 9524
rect 8464 9468 8492 9524
rect 8548 9468 8576 9524
rect 8632 9468 8660 9524
rect 8716 9468 8744 9524
rect 8800 9468 8828 9524
rect 8884 9468 8885 9524
rect 8323 9443 8885 9468
rect 8323 9387 8324 9443
rect 8380 9387 8408 9443
rect 8464 9387 8492 9443
rect 8548 9387 8576 9443
rect 8632 9387 8660 9443
rect 8716 9387 8744 9443
rect 8800 9387 8828 9443
rect 8884 9387 8885 9443
rect 8323 9362 8885 9387
rect 8323 9306 8324 9362
rect 8380 9306 8408 9362
rect 8464 9306 8492 9362
rect 8548 9306 8576 9362
rect 8632 9306 8660 9362
rect 8716 9306 8744 9362
rect 8800 9306 8828 9362
rect 8884 9306 8885 9362
rect 8323 9281 8885 9306
rect 8323 9225 8324 9281
rect 8380 9225 8408 9281
rect 8464 9225 8492 9281
rect 8548 9225 8576 9281
rect 8632 9225 8660 9281
rect 8716 9225 8744 9281
rect 8800 9225 8828 9281
rect 8884 9225 8885 9281
rect 8323 9200 8885 9225
rect 8323 9144 8324 9200
rect 8380 9144 8408 9200
rect 8464 9144 8492 9200
rect 8548 9144 8576 9200
rect 8632 9144 8660 9200
rect 8716 9144 8744 9200
rect 8800 9144 8828 9200
rect 8884 9144 8885 9200
rect 8323 9119 8885 9144
rect 8323 9063 8324 9119
rect 8380 9063 8408 9119
rect 8464 9063 8492 9119
rect 8548 9063 8576 9119
rect 8632 9063 8660 9119
rect 8716 9063 8744 9119
rect 8800 9063 8828 9119
rect 8884 9063 8885 9119
rect 8323 9038 8885 9063
rect 8323 8982 8324 9038
rect 8380 8982 8408 9038
rect 8464 8982 8492 9038
rect 8548 8982 8576 9038
rect 8632 8982 8660 9038
rect 8716 8982 8744 9038
rect 8800 8982 8828 9038
rect 8884 8982 8885 9038
rect 8323 8957 8885 8982
rect 8323 8901 8324 8957
rect 8380 8901 8408 8957
rect 8464 8901 8492 8957
rect 8548 8901 8576 8957
rect 8632 8901 8660 8957
rect 8716 8901 8744 8957
rect 8800 8901 8828 8957
rect 8884 8901 8885 8957
rect 8323 8876 8885 8901
rect 8323 8820 8324 8876
rect 8380 8820 8408 8876
rect 8464 8820 8492 8876
rect 8548 8820 8576 8876
rect 8632 8820 8660 8876
rect 8716 8820 8744 8876
rect 8800 8820 8828 8876
rect 8884 8820 8885 8876
rect 8323 8795 8885 8820
rect 8323 8739 8324 8795
rect 8380 8739 8408 8795
rect 8464 8739 8492 8795
rect 8548 8739 8576 8795
rect 8632 8739 8660 8795
rect 8716 8739 8744 8795
rect 8800 8739 8828 8795
rect 8884 8739 8885 8795
rect 8323 8714 8885 8739
rect 8323 8658 8324 8714
rect 8380 8658 8408 8714
rect 8464 8658 8492 8714
rect 8548 8658 8576 8714
rect 8632 8658 8660 8714
rect 8716 8658 8744 8714
rect 8800 8658 8828 8714
rect 8884 8658 8885 8714
rect 8323 8633 8885 8658
rect 8323 8577 8324 8633
rect 8380 8577 8408 8633
rect 8464 8577 8492 8633
rect 8548 8577 8576 8633
rect 8632 8577 8660 8633
rect 8716 8577 8744 8633
rect 8800 8577 8828 8633
rect 8884 8577 8885 8633
rect 8323 8552 8885 8577
rect 8323 8496 8324 8552
rect 8380 8496 8408 8552
rect 8464 8496 8492 8552
rect 8548 8496 8576 8552
rect 8632 8496 8660 8552
rect 8716 8496 8744 8552
rect 8800 8496 8828 8552
rect 8884 8496 8885 8552
rect 8323 8471 8885 8496
rect 8323 8415 8324 8471
rect 8380 8415 8408 8471
rect 8464 8415 8492 8471
rect 8548 8415 8576 8471
rect 8632 8415 8660 8471
rect 8716 8415 8744 8471
rect 8800 8415 8828 8471
rect 8884 8415 8885 8471
rect 8323 8390 8885 8415
rect 8323 8334 8324 8390
rect 8380 8334 8408 8390
rect 8464 8334 8492 8390
rect 8548 8334 8576 8390
rect 8632 8334 8660 8390
rect 8716 8334 8744 8390
rect 8800 8334 8828 8390
rect 8884 8334 8885 8390
rect 8323 8309 8885 8334
rect 8323 8253 8324 8309
rect 8380 8253 8408 8309
rect 8464 8253 8492 8309
rect 8548 8253 8576 8309
rect 8632 8253 8660 8309
rect 8716 8253 8744 8309
rect 8800 8253 8828 8309
rect 8884 8253 8885 8309
rect 8323 8228 8885 8253
rect 8323 8172 8324 8228
rect 8380 8172 8408 8228
rect 8464 8172 8492 8228
rect 8548 8172 8576 8228
rect 8632 8172 8660 8228
rect 8716 8172 8744 8228
rect 8800 8172 8828 8228
rect 8884 8172 8885 8228
rect 8323 8147 8885 8172
rect 8323 8091 8324 8147
rect 8380 8091 8408 8147
rect 8464 8091 8492 8147
rect 8548 8091 8576 8147
rect 8632 8091 8660 8147
rect 8716 8091 8744 8147
rect 8800 8091 8828 8147
rect 8884 8091 8885 8147
rect 8323 8066 8885 8091
rect 8323 8010 8324 8066
rect 8380 8010 8408 8066
rect 8464 8010 8492 8066
rect 8548 8010 8576 8066
rect 8632 8010 8660 8066
rect 8716 8010 8744 8066
rect 8800 8010 8828 8066
rect 8884 8010 8885 8066
rect 8323 7985 8885 8010
rect 8323 7929 8324 7985
rect 8380 7929 8408 7985
rect 8464 7929 8492 7985
rect 8548 7929 8576 7985
rect 8632 7929 8660 7985
rect 8716 7929 8744 7985
rect 8800 7929 8828 7985
rect 8884 7929 8885 7985
rect 8323 7904 8885 7929
rect 8323 7848 8324 7904
rect 8380 7848 8408 7904
rect 8464 7848 8492 7904
rect 8548 7848 8576 7904
rect 8632 7848 8660 7904
rect 8716 7848 8744 7904
rect 8800 7848 8828 7904
rect 8884 7848 8885 7904
rect 8323 7823 8885 7848
rect 8323 7767 8324 7823
rect 8380 7767 8408 7823
rect 8464 7767 8492 7823
rect 8548 7767 8576 7823
rect 8632 7767 8660 7823
rect 8716 7767 8744 7823
rect 8800 7767 8828 7823
rect 8884 7767 8885 7823
rect 8323 7742 8885 7767
rect 8323 7686 8324 7742
rect 8380 7686 8408 7742
rect 8464 7686 8492 7742
rect 8548 7686 8576 7742
rect 8632 7686 8660 7742
rect 8716 7686 8744 7742
rect 8800 7686 8828 7742
rect 8884 7686 8885 7742
rect 8323 7661 8885 7686
rect 8323 7605 8324 7661
rect 8380 7605 8408 7661
rect 8464 7605 8492 7661
rect 8548 7605 8576 7661
rect 8632 7605 8660 7661
rect 8716 7605 8744 7661
rect 8800 7605 8828 7661
rect 8884 7605 8885 7661
rect 8323 7580 8885 7605
rect 8323 7524 8324 7580
rect 8380 7524 8408 7580
rect 8464 7524 8492 7580
rect 8548 7524 8576 7580
rect 8632 7524 8660 7580
rect 8716 7524 8744 7580
rect 8800 7524 8828 7580
rect 8884 7524 8885 7580
rect 8323 7499 8885 7524
rect 8323 7443 8324 7499
rect 8380 7443 8408 7499
rect 8464 7443 8492 7499
rect 8548 7443 8576 7499
rect 8632 7443 8660 7499
rect 8716 7443 8744 7499
rect 8800 7443 8828 7499
rect 8884 7443 8885 7499
rect 8323 7418 8885 7443
rect 8323 7362 8324 7418
rect 8380 7362 8408 7418
rect 8464 7362 8492 7418
rect 8548 7362 8576 7418
rect 8632 7362 8660 7418
rect 8716 7362 8744 7418
rect 8800 7362 8828 7418
rect 8884 7362 8885 7418
rect 8323 7337 8885 7362
rect 8323 7281 8324 7337
rect 8380 7281 8408 7337
rect 8464 7281 8492 7337
rect 8548 7281 8576 7337
rect 8632 7281 8660 7337
rect 8716 7281 8744 7337
rect 8800 7281 8828 7337
rect 8884 7281 8885 7337
rect 8323 7256 8885 7281
rect 8323 7200 8324 7256
rect 8380 7200 8408 7256
rect 8464 7200 8492 7256
rect 8548 7200 8576 7256
rect 8632 7200 8660 7256
rect 8716 7200 8744 7256
rect 8800 7200 8828 7256
rect 8884 7200 8885 7256
rect 8323 7175 8885 7200
rect 8323 7119 8324 7175
rect 8380 7119 8408 7175
rect 8464 7119 8492 7175
rect 8548 7119 8576 7175
rect 8632 7119 8660 7175
rect 8716 7119 8744 7175
rect 8800 7119 8828 7175
rect 8884 7119 8885 7175
rect 8323 7094 8885 7119
rect 8323 7038 8324 7094
rect 8380 7038 8408 7094
rect 8464 7038 8492 7094
rect 8548 7038 8576 7094
rect 8632 7038 8660 7094
rect 8716 7038 8744 7094
rect 8800 7038 8828 7094
rect 8884 7038 8885 7094
rect 8323 7013 8885 7038
rect 8323 6957 8324 7013
rect 8380 6957 8408 7013
rect 8464 6957 8492 7013
rect 8548 6957 8576 7013
rect 8632 6957 8660 7013
rect 8716 6957 8744 7013
rect 8800 6957 8828 7013
rect 8884 6957 8885 7013
rect 8323 6932 8885 6957
rect 8323 6876 8324 6932
rect 8380 6876 8408 6932
rect 8464 6876 8492 6932
rect 8548 6876 8576 6932
rect 8632 6876 8660 6932
rect 8716 6876 8744 6932
rect 8800 6876 8828 6932
rect 8884 6876 8885 6932
rect 8323 6851 8885 6876
rect 8323 6795 8324 6851
rect 8380 6795 8408 6851
rect 8464 6795 8492 6851
rect 8548 6795 8576 6851
rect 8632 6795 8660 6851
rect 8716 6795 8744 6851
rect 8800 6795 8828 6851
rect 8884 6795 8885 6851
rect 8323 6770 8885 6795
rect 8323 6714 8324 6770
rect 8380 6714 8408 6770
rect 8464 6714 8492 6770
rect 8548 6714 8576 6770
rect 8632 6714 8660 6770
rect 8716 6714 8744 6770
rect 8800 6714 8828 6770
rect 8884 6714 8885 6770
rect 8323 6689 8885 6714
rect 8323 6633 8324 6689
rect 8380 6633 8408 6689
rect 8464 6633 8492 6689
rect 8548 6633 8576 6689
rect 8632 6633 8660 6689
rect 8716 6633 8744 6689
rect 8800 6633 8828 6689
rect 8884 6633 8885 6689
rect 8323 6608 8885 6633
rect 8323 6552 8324 6608
rect 8380 6552 8408 6608
rect 8464 6552 8492 6608
rect 8548 6552 8576 6608
rect 8632 6552 8660 6608
rect 8716 6552 8744 6608
rect 8800 6552 8828 6608
rect 8884 6552 8885 6608
rect 8323 6527 8885 6552
rect 8323 6471 8324 6527
rect 8380 6471 8408 6527
rect 8464 6471 8492 6527
rect 8548 6471 8576 6527
rect 8632 6471 8660 6527
rect 8716 6471 8744 6527
rect 8800 6471 8828 6527
rect 8884 6471 8885 6527
rect 8323 6446 8885 6471
rect 8323 6390 8324 6446
rect 8380 6390 8408 6446
rect 8464 6390 8492 6446
rect 8548 6390 8576 6446
rect 8632 6390 8660 6446
rect 8716 6390 8744 6446
rect 8800 6390 8828 6446
rect 8884 6390 8885 6446
rect 8323 6365 8885 6390
rect 8323 6309 8324 6365
rect 8380 6309 8408 6365
rect 8464 6309 8492 6365
rect 8548 6309 8576 6365
rect 8632 6309 8660 6365
rect 8716 6309 8744 6365
rect 8800 6309 8828 6365
rect 8884 6309 8885 6365
rect 8323 6284 8885 6309
rect 8323 6228 8324 6284
rect 8380 6228 8408 6284
rect 8464 6228 8492 6284
rect 8548 6228 8576 6284
rect 8632 6228 8660 6284
rect 8716 6228 8744 6284
rect 8800 6228 8828 6284
rect 8884 6228 8885 6284
rect 8323 6203 8885 6228
rect 8323 6147 8324 6203
rect 8380 6147 8408 6203
rect 8464 6147 8492 6203
rect 8548 6147 8576 6203
rect 8632 6147 8660 6203
rect 8716 6147 8744 6203
rect 8800 6147 8828 6203
rect 8884 6147 8885 6203
rect 8323 6122 8885 6147
rect 8323 6066 8324 6122
rect 8380 6066 8408 6122
rect 8464 6066 8492 6122
rect 8548 6066 8576 6122
rect 8632 6066 8660 6122
rect 8716 6066 8744 6122
rect 8800 6066 8828 6122
rect 8884 6066 8885 6122
rect 8323 6041 8885 6066
rect 8323 5985 8324 6041
rect 8380 5985 8408 6041
rect 8464 5985 8492 6041
rect 8548 5985 8576 6041
rect 8632 5985 8660 6041
rect 8716 5985 8744 6041
rect 8800 5985 8828 6041
rect 8884 5985 8885 6041
rect 8323 5960 8885 5985
rect 8323 5904 8324 5960
rect 8380 5904 8408 5960
rect 8464 5904 8492 5960
rect 8548 5904 8576 5960
rect 8632 5904 8660 5960
rect 8716 5904 8744 5960
rect 8800 5904 8828 5960
rect 8884 5904 8885 5960
rect 8323 5879 8885 5904
rect 8323 5823 8324 5879
rect 8380 5823 8408 5879
rect 8464 5823 8492 5879
rect 8548 5823 8576 5879
rect 8632 5823 8660 5879
rect 8716 5823 8744 5879
rect 8800 5823 8828 5879
rect 8884 5823 8885 5879
rect 8323 5798 8885 5823
rect 8323 5742 8324 5798
rect 8380 5742 8408 5798
rect 8464 5742 8492 5798
rect 8548 5742 8576 5798
rect 8632 5742 8660 5798
rect 8716 5742 8744 5798
rect 8800 5742 8828 5798
rect 8884 5742 8885 5798
rect 8323 5717 8885 5742
rect 8323 5661 8324 5717
rect 8380 5661 8408 5717
rect 8464 5661 8492 5717
rect 8548 5661 8576 5717
rect 8632 5661 8660 5717
rect 8716 5661 8744 5717
rect 8800 5661 8828 5717
rect 8884 5661 8885 5717
rect 8323 5636 8885 5661
rect 8323 5580 8324 5636
rect 8380 5580 8408 5636
rect 8464 5580 8492 5636
rect 8548 5580 8576 5636
rect 8632 5580 8660 5636
rect 8716 5580 8744 5636
rect 8800 5580 8828 5636
rect 8884 5580 8885 5636
rect 8323 5555 8885 5580
rect 8323 5499 8324 5555
rect 8380 5499 8408 5555
rect 8464 5499 8492 5555
rect 8548 5499 8576 5555
rect 8632 5499 8660 5555
rect 8716 5499 8744 5555
rect 8800 5499 8828 5555
rect 8884 5499 8885 5555
rect 8323 5474 8885 5499
rect 8323 5418 8324 5474
rect 8380 5418 8408 5474
rect 8464 5418 8492 5474
rect 8548 5418 8576 5474
rect 8632 5418 8660 5474
rect 8716 5418 8744 5474
rect 8800 5418 8828 5474
rect 8884 5418 8885 5474
rect 8323 5393 8885 5418
rect 8323 5337 8324 5393
rect 8380 5337 8408 5393
rect 8464 5337 8492 5393
rect 8548 5337 8576 5393
rect 8632 5337 8660 5393
rect 8716 5337 8744 5393
rect 8800 5337 8828 5393
rect 8884 5337 8885 5393
rect 8323 5312 8885 5337
rect 8323 5256 8324 5312
rect 8380 5256 8408 5312
rect 8464 5256 8492 5312
rect 8548 5256 8576 5312
rect 8632 5256 8660 5312
rect 8716 5256 8744 5312
rect 8800 5256 8828 5312
rect 8884 5256 8885 5312
rect 8323 5231 8885 5256
tri 195 5191 214 5210 ne
rect 214 5191 216 5210
tri 752 5191 771 5210 nw
tri 1999 5191 2018 5210 ne
rect 2018 5191 2020 5210
tri 2556 5191 2575 5210 nw
tri 3803 5191 3822 5210 ne
rect 3822 5191 3824 5210
tri 4360 5191 4379 5210 nw
tri 5607 5191 5626 5210 ne
rect 5626 5191 5628 5210
tri 6164 5191 6183 5210 nw
tri 7411 5191 7430 5210 ne
rect 7430 5191 7433 5210
tri 7969 5193 7986 5210 nw
tri 214 5189 216 5191 ne
tri 2018 5189 2020 5191 ne
tri 3822 5189 3824 5191 ne
tri 5626 5189 5628 5191 ne
tri 7430 5189 7432 5191 ne
rect 7432 5189 7433 5191
tri 7432 5188 7433 5189 ne
rect -724 5130 -122 5155
rect -724 5074 -714 5130
rect -658 5074 -626 5130
rect -570 5074 -538 5130
rect -482 5074 -450 5130
rect -394 5074 -362 5130
rect -306 5074 -274 5130
rect -218 5074 -186 5130
rect -130 5074 -122 5130
rect 8323 5175 8324 5231
rect 8380 5175 8408 5231
rect 8464 5175 8492 5231
rect 8548 5175 8576 5231
rect 8632 5175 8660 5231
rect 8716 5175 8744 5231
rect 8800 5175 8828 5231
rect 8884 5175 8885 5231
rect 10116 5210 10692 12116
tri 9212 5188 9234 5210 ne
tri 9770 5193 9787 5210 nw
tri 11025 5193 11042 5210 ne
rect 11042 5193 11047 5210
tri 11583 5196 11597 5210 nw
tri 11042 5188 11047 5193 ne
rect 8323 5150 8885 5175
rect 8323 5094 8324 5150
rect 8380 5094 8408 5150
rect 8464 5094 8492 5150
rect 8548 5094 8576 5150
rect 8632 5094 8660 5150
rect 8716 5094 8744 5150
rect 8800 5094 8828 5150
rect 8884 5094 8885 5150
rect -724 5049 -122 5074
tri -3750 4934 -3657 5027 nw
tri -2614 4942 -2529 5027 ne
rect -2529 4942 -2136 5027
tri -2136 4942 -2051 5027 nw
rect -724 4993 -714 5049
rect -658 4993 -626 5049
rect -570 4993 -538 5049
rect -482 4993 -450 5049
rect -394 4993 -362 5049
rect -306 4993 -274 5049
rect -218 4993 -186 5049
rect -130 5027 -122 5049
tri -122 5027 -59 5090 sw
rect 8323 5069 8885 5094
rect -130 4993 -59 5027
rect -724 4968 -59 4993
tri -2529 4939 -2526 4942 ne
rect -2526 3016 -2136 4942
rect -724 4912 -714 4968
rect -658 4912 -626 4968
rect -570 4912 -538 4968
rect -482 4912 -450 4968
rect -394 4912 -362 4968
rect -306 4912 -274 4968
rect -218 4912 -186 4968
rect -130 4934 -59 4968
tri -59 4934 34 5027 sw
rect 8323 5013 8324 5069
rect 8380 5013 8408 5069
rect 8464 5013 8492 5069
rect 8548 5013 8576 5069
rect 8632 5013 8660 5069
rect 8716 5013 8744 5069
rect 8800 5013 8828 5069
rect 8884 5013 8885 5069
rect 8323 4988 8885 5013
rect -130 4912 34 4934
rect -724 4887 34 4912
rect -724 4831 -714 4887
rect -658 4831 -626 4887
rect -570 4831 -538 4887
rect -482 4831 -450 4887
rect -394 4831 -362 4887
rect -306 4831 -274 4887
rect -218 4831 -186 4887
rect -130 4879 34 4887
tri 34 4879 89 4934 sw
rect 8323 4932 8324 4988
rect 8380 4932 8408 4988
rect 8464 4932 8492 4988
rect 8548 4932 8576 4988
rect 8632 4932 8660 4988
rect 8716 4932 8744 4988
rect 8800 4932 8828 4988
rect 8884 4932 8885 4988
tri 11564 4934 11657 5027 se
rect 11657 4934 11859 12440
rect 11919 5139 12495 12180
rect 8323 4907 8885 4932
rect -130 4839 89 4879
tri 89 4839 129 4879 sw
rect 8323 4851 8324 4907
rect 8380 4851 8408 4907
rect 8464 4851 8492 4907
rect 8548 4851 8576 4907
rect 8632 4851 8660 4907
rect 8716 4851 8744 4907
rect 8800 4851 8828 4907
rect 8884 4851 8885 4907
tri 11509 4879 11564 4934 se
rect 11564 4879 11859 4934
tri 11859 4879 12007 5027 sw
tri 12411 4879 12559 5027 se
rect -130 4831 -122 4839
rect -724 4806 -122 4831
rect -724 4750 -714 4806
rect -658 4750 -626 4806
rect -570 4750 -538 4806
rect -482 4750 -450 4806
rect -394 4750 -362 4806
rect -306 4750 -274 4806
rect -218 4750 -186 4806
rect -130 4750 -122 4806
tri -1577 4729 -1567 4739 se
tri -1055 4729 -1046 4738 sw
rect -724 4725 -122 4750
rect -724 4669 -714 4725
rect -658 4669 -626 4725
rect -570 4669 -538 4725
rect -482 4669 -450 4725
rect -394 4669 -362 4725
rect -306 4669 -274 4725
rect -218 4669 -186 4725
rect -130 4669 -122 4725
rect -724 4644 -122 4669
rect -724 4588 -714 4644
rect -658 4588 -626 4644
rect -570 4588 -538 4644
rect -482 4588 -450 4644
rect -394 4588 -362 4644
rect -306 4588 -274 4644
rect -218 4588 -186 4644
rect -130 4588 -122 4644
rect -724 4563 -122 4588
rect -724 4507 -714 4563
rect -658 4507 -626 4563
rect -570 4507 -538 4563
rect -482 4507 -450 4563
rect -394 4507 -362 4563
rect -306 4507 -274 4563
rect -218 4507 -186 4563
rect -130 4507 -122 4563
rect -724 4482 -122 4507
rect -724 4426 -714 4482
rect -658 4426 -626 4482
rect -570 4426 -538 4482
rect -482 4426 -450 4482
rect -394 4426 -362 4482
rect -306 4426 -274 4482
rect -218 4426 -186 4482
rect -130 4426 -122 4482
rect -724 4401 -122 4426
rect -724 4345 -714 4401
rect -658 4345 -626 4401
rect -570 4345 -538 4401
rect -482 4345 -450 4401
rect -394 4345 -362 4401
rect -306 4345 -274 4401
rect -218 4345 -186 4401
rect -130 4345 -122 4401
rect -724 4320 -122 4345
rect -724 4264 -714 4320
rect -658 4264 -626 4320
rect -570 4264 -538 4320
rect -482 4264 -450 4320
rect -394 4264 -362 4320
rect -306 4264 -274 4320
rect -218 4264 -186 4320
rect -130 4264 -122 4320
rect -724 4239 -122 4264
rect -724 4183 -714 4239
rect -658 4183 -626 4239
rect -570 4183 -538 4239
rect -482 4183 -450 4239
rect -394 4183 -362 4239
rect -306 4183 -274 4239
rect -218 4183 -186 4239
rect -130 4183 -122 4239
rect -724 4158 -122 4183
rect -724 4102 -714 4158
rect -658 4102 -626 4158
rect -570 4102 -538 4158
rect -482 4102 -450 4158
rect -394 4102 -362 4158
rect -306 4102 -274 4158
rect -218 4102 -186 4158
rect -130 4102 -122 4158
rect -724 4077 -122 4102
rect -724 4021 -714 4077
rect -658 4021 -626 4077
rect -570 4021 -538 4077
rect -482 4021 -450 4077
rect -394 4021 -362 4077
rect -306 4021 -274 4077
rect -218 4021 -186 4077
rect -130 4021 -122 4077
rect -724 3996 -122 4021
rect -724 3940 -714 3996
rect -658 3940 -626 3996
rect -570 3940 -538 3996
rect -482 3940 -450 3996
rect -394 3940 -362 3996
rect -306 3940 -274 3996
rect -218 3940 -186 3996
rect -130 3940 -122 3996
rect -724 3915 -122 3940
rect -724 3859 -714 3915
rect -658 3859 -626 3915
rect -570 3859 -538 3915
rect -482 3859 -450 3915
rect -394 3859 -362 3915
rect -306 3859 -274 3915
rect -218 3859 -186 3915
rect -130 3859 -122 3915
rect -724 3834 -122 3859
rect -724 3778 -714 3834
rect -658 3778 -626 3834
rect -570 3778 -538 3834
rect -482 3778 -450 3834
rect -394 3778 -362 3834
rect -306 3778 -274 3834
rect -218 3778 -186 3834
rect -130 3778 -122 3834
rect -724 3753 -122 3778
rect -724 3697 -714 3753
rect -658 3697 -626 3753
rect -570 3697 -538 3753
rect -482 3697 -450 3753
rect -394 3697 -362 3753
rect -306 3697 -274 3753
rect -218 3697 -186 3753
rect -130 3697 -122 3753
rect -724 3672 -122 3697
rect -724 3616 -714 3672
rect -658 3616 -626 3672
rect -570 3616 -538 3672
rect -482 3616 -450 3672
rect -394 3616 -362 3672
rect -306 3616 -274 3672
rect -218 3616 -186 3672
rect -130 3616 -122 3672
rect -724 3591 -122 3616
rect -724 3535 -714 3591
rect -658 3535 -626 3591
rect -570 3535 -538 3591
rect -482 3535 -450 3591
rect -394 3535 -362 3591
rect -306 3535 -274 3591
rect -218 3535 -186 3591
rect -130 3535 -122 3591
rect 8323 4826 8885 4851
rect 11657 4839 11859 4879
rect 12559 4839 12761 12440
tri 12761 4879 12909 5027 sw
tri 13313 4879 13461 5027 se
rect 13461 4839 13663 12440
tri 13663 4879 13811 5027 sw
tri 14251 4879 14399 5027 se
rect 8323 4770 8324 4826
rect 8380 4770 8408 4826
rect 8464 4770 8492 4826
rect 8548 4770 8576 4826
rect 8632 4770 8660 4826
rect 8716 4770 8744 4826
rect 8800 4770 8828 4826
rect 8884 4770 8885 4826
rect 8323 4745 8885 4770
rect 8323 4689 8324 4745
rect 8380 4689 8408 4745
rect 8464 4689 8492 4745
rect 8548 4689 8576 4745
rect 8632 4689 8660 4745
rect 8716 4689 8744 4745
rect 8800 4689 8828 4745
rect 8884 4689 8885 4745
rect 8323 4664 8885 4689
rect 8323 4608 8324 4664
rect 8380 4608 8408 4664
rect 8464 4608 8492 4664
rect 8548 4608 8576 4664
rect 8632 4608 8660 4664
rect 8716 4608 8744 4664
rect 8800 4608 8828 4664
rect 8884 4608 8885 4664
rect 8323 4583 8885 4608
rect 8323 4527 8324 4583
rect 8380 4527 8408 4583
rect 8464 4527 8492 4583
rect 8548 4527 8576 4583
rect 8632 4527 8660 4583
rect 8716 4527 8744 4583
rect 8800 4527 8828 4583
rect 8884 4527 8885 4583
rect 8323 4502 8885 4527
rect 8323 4446 8324 4502
rect 8380 4446 8408 4502
rect 8464 4446 8492 4502
rect 8548 4446 8576 4502
rect 8632 4446 8660 4502
rect 8716 4446 8744 4502
rect 8800 4446 8828 4502
rect 8884 4446 8885 4502
rect 8323 4421 8885 4446
rect 8323 4365 8324 4421
rect 8380 4365 8408 4421
rect 8464 4365 8492 4421
rect 8548 4365 8576 4421
rect 8632 4365 8660 4421
rect 8716 4365 8744 4421
rect 8800 4365 8828 4421
rect 8884 4365 8885 4421
rect 8323 4340 8885 4365
rect 8323 4284 8324 4340
rect 8380 4284 8408 4340
rect 8464 4284 8492 4340
rect 8548 4284 8576 4340
rect 8632 4284 8660 4340
rect 8716 4284 8744 4340
rect 8800 4284 8828 4340
rect 8884 4284 8885 4340
rect 8323 4259 8885 4284
rect 8323 4203 8324 4259
rect 8380 4203 8408 4259
rect 8464 4203 8492 4259
rect 8548 4203 8576 4259
rect 8632 4203 8660 4259
rect 8716 4203 8744 4259
rect 8800 4203 8828 4259
rect 8884 4203 8885 4259
rect 8323 4178 8885 4203
rect 8323 4122 8324 4178
rect 8380 4122 8408 4178
rect 8464 4122 8492 4178
rect 8548 4122 8576 4178
rect 8632 4122 8660 4178
rect 8716 4122 8744 4178
rect 8800 4122 8828 4178
rect 8884 4122 8885 4178
rect 8323 4097 8885 4122
rect 8323 4041 8324 4097
rect 8380 4041 8408 4097
rect 8464 4041 8492 4097
rect 8548 4041 8576 4097
rect 8632 4041 8660 4097
rect 8716 4041 8744 4097
rect 8800 4041 8828 4097
rect 8884 4041 8885 4097
rect 14399 4086 15130 13060
rect 8323 4016 8885 4041
rect 8323 3960 8324 4016
rect 8380 3960 8408 4016
rect 8464 3960 8492 4016
rect 8548 3960 8576 4016
rect 8632 3960 8660 4016
rect 8716 3960 8744 4016
rect 8800 3960 8828 4016
rect 8884 3960 8885 4016
rect 8323 3935 8885 3960
rect 8323 3879 8324 3935
rect 8380 3879 8408 3935
rect 8464 3879 8492 3935
rect 8548 3879 8576 3935
rect 8632 3879 8660 3935
rect 8716 3879 8744 3935
rect 8800 3879 8828 3935
rect 8884 3879 8885 3935
rect 8323 3854 8885 3879
rect 8323 3798 8324 3854
rect 8380 3798 8408 3854
rect 8464 3798 8492 3854
rect 8548 3798 8576 3854
rect 8632 3798 8660 3854
rect 8716 3798 8744 3854
rect 8800 3798 8828 3854
rect 8884 3798 8885 3854
tri 14431 3831 14686 4086 nw
rect 8323 3773 8885 3798
rect 8323 3717 8324 3773
rect 8380 3717 8408 3773
rect 8464 3717 8492 3773
rect 8548 3717 8576 3773
rect 8632 3717 8660 3773
rect 8716 3717 8744 3773
rect 8800 3717 8828 3773
rect 8884 3717 8885 3773
rect 8323 3692 8885 3717
rect 8323 3636 8324 3692
rect 8380 3636 8408 3692
rect 8464 3636 8492 3692
rect 8548 3636 8576 3692
rect 8632 3636 8660 3692
rect 8716 3636 8744 3692
rect 8800 3636 8828 3692
rect 8884 3636 8885 3692
rect 8323 3611 8885 3636
rect 8323 3555 8324 3611
rect 8380 3555 8408 3611
rect 8464 3555 8492 3611
rect 8548 3555 8576 3611
rect 8632 3555 8660 3611
rect 8716 3555 8744 3611
rect 8800 3555 8828 3611
rect 8884 3555 8885 3611
rect 8323 3546 8885 3555
rect -724 3510 -122 3535
rect -724 3454 -714 3510
rect -658 3454 -626 3510
rect -570 3454 -538 3510
rect -482 3454 -450 3510
rect -394 3454 -362 3510
rect -306 3454 -274 3510
rect -218 3454 -186 3510
rect -130 3454 -122 3510
rect -724 3429 -122 3454
rect -724 3373 -714 3429
rect -658 3373 -626 3429
rect -570 3373 -538 3429
rect -482 3373 -450 3429
rect -394 3373 -362 3429
rect -306 3373 -274 3429
rect -218 3373 -186 3429
rect -130 3373 -122 3429
rect -724 3348 -122 3373
rect -724 3292 -714 3348
rect -658 3292 -626 3348
rect -570 3292 -538 3348
rect -482 3292 -450 3348
rect -394 3292 -362 3348
rect -306 3292 -274 3348
rect -218 3292 -186 3348
rect -130 3292 -122 3348
rect -724 3267 -122 3292
rect -724 3211 -714 3267
rect -658 3211 -626 3267
rect -570 3211 -538 3267
rect -482 3211 -450 3267
rect -394 3211 -362 3267
rect -306 3211 -274 3267
rect -218 3211 -186 3267
rect -130 3211 -122 3267
rect -724 3192 -122 3211
tri -2136 3016 -1970 3182 sw
tri -4330 2972 -4286 3016 se
rect -2526 2992 -1970 3016
tri -1970 2992 -1946 3016 sw
tri -3750 2972 -3730 2992 sw
rect -4330 0 -3730 2972
rect -2526 2972 -1946 2992
tri -1946 2972 -1926 2992 sw
rect -2526 0 -1926 2972
rect -722 0 -122 2972
tri -31 0 -26 5 se
rect 1082 0 1682 2972
rect 2886 0 3486 2972
rect 4690 229 5272 2972
rect 6494 0 7094 2972
rect 8298 0 8898 2972
rect 8964 981 8970 1033
rect 9022 981 9038 1033
rect 9090 981 9096 1033
rect 9005 929 9057 981
rect 9006 927 9056 928
rect 9005 891 9057 927
rect 9006 890 9056 891
rect 9005 703 9057 889
rect 8964 651 8970 703
rect 9022 651 9038 703
rect 9090 651 9096 703
rect 10102 34 10702 2972
rect 10740 981 10746 1033
rect 10798 981 10814 1033
rect 10866 981 10872 1033
rect 11709 981 11715 1033
rect 11767 981 11783 1033
rect 11835 981 11841 1033
rect 10781 929 10833 981
rect 10782 927 10832 928
rect 11750 929 11802 981
rect 11751 927 11801 928
rect 10782 890 10832 891
rect 10781 703 10833 889
rect 11751 890 11801 891
rect 11750 703 11802 889
rect 10740 651 10746 703
rect 10798 651 10814 703
rect 10866 651 10872 703
rect 11709 651 11715 703
rect 11767 651 11783 703
rect 11835 651 11841 703
rect 11906 0 12506 2972
rect 13710 1100 14310 2972
rect 13710 981 14191 1100
tri 14191 981 14310 1100 nw
rect 13710 0 14175 981
tri 14175 965 14191 981 nw
tri -4326 -18 -4308 0 ne
rect -4308 -18 -4299 0
tri -4308 -27 -4299 -18 ne
rect -3763 -18 -3754 0
tri -3754 -18 -3736 0 nw
tri -2526 -18 -2508 0 ne
rect -1972 -18 -1963 0
tri -1963 -18 -1945 0 nw
tri -715 -18 -697 0 ne
rect -697 -18 -688 0
tri -3763 -27 -3754 -18 nw
tri -1972 -27 -1963 -18 nw
tri -697 -27 -688 -18 ne
tri -152 -27 -125 0 nw
<< rmetal2 >>
rect 9005 928 9057 929
rect 9005 927 9006 928
rect 9056 927 9057 928
rect 9005 890 9006 891
rect 9056 890 9057 891
rect 9005 889 9057 890
rect 10781 928 10833 929
rect 10781 927 10782 928
rect 10832 927 10833 928
rect 11750 928 11802 929
rect 11750 927 11751 928
rect 11801 927 11802 928
rect 10781 890 10782 891
rect 10832 890 10833 891
rect 10781 889 10833 890
rect 11750 890 11751 891
rect 11801 890 11802 891
rect 11750 889 11802 890
<< via2 >>
rect -711 20491 -655 20547
rect -625 20491 -569 20547
rect -539 20491 -483 20547
rect -453 20491 -397 20547
rect -367 20491 -311 20547
rect -281 20491 -225 20547
rect -195 20491 -139 20547
rect -711 20399 -655 20455
rect -625 20399 -569 20455
rect -539 20399 -483 20455
rect -453 20399 -397 20455
rect -367 20399 -311 20455
rect -281 20399 -225 20455
rect -195 20399 -139 20455
rect -711 20307 -655 20363
rect -625 20307 -569 20363
rect -539 20307 -483 20363
rect -453 20307 -397 20363
rect -367 20307 -311 20363
rect -281 20307 -225 20363
rect -195 20307 -139 20363
rect -711 20215 -655 20271
rect -625 20215 -569 20271
rect -539 20215 -483 20271
rect -453 20215 -397 20271
rect -367 20215 -311 20271
rect -281 20215 -225 20271
rect -195 20215 -139 20271
rect -711 20123 -655 20179
rect -625 20123 -569 20179
rect -539 20123 -483 20179
rect -453 20123 -397 20179
rect -367 20123 -311 20179
rect -281 20123 -225 20179
rect -195 20123 -139 20179
rect -711 20030 -655 20086
rect -625 20030 -569 20086
rect -539 20030 -483 20086
rect -453 20030 -397 20086
rect -367 20030 -311 20086
rect -281 20030 -225 20086
rect -195 20030 -139 20086
rect -711 19937 -655 19993
rect -625 19937 -569 19993
rect -539 19937 -483 19993
rect -453 19937 -397 19993
rect -367 19937 -311 19993
rect -281 19937 -225 19993
rect -195 19937 -139 19993
rect 1106 20494 1162 20550
rect 1188 20494 1244 20550
rect 1270 20494 1326 20550
rect 1352 20494 1408 20550
rect 1434 20494 1490 20550
rect 1516 20494 1572 20550
rect 1598 20494 1654 20550
rect 1106 20414 1162 20470
rect 1188 20414 1244 20470
rect 1270 20414 1326 20470
rect 1352 20414 1408 20470
rect 1434 20414 1490 20470
rect 1516 20414 1572 20470
rect 1598 20414 1654 20470
rect 1106 20334 1162 20390
rect 1188 20334 1244 20390
rect 1270 20334 1326 20390
rect 1352 20334 1408 20390
rect 1434 20334 1490 20390
rect 1516 20334 1572 20390
rect 1598 20334 1654 20390
rect 1106 20254 1162 20310
rect 1188 20254 1244 20310
rect 1270 20254 1326 20310
rect 1352 20254 1408 20310
rect 1434 20254 1490 20310
rect 1516 20254 1572 20310
rect 1598 20254 1654 20310
rect 1106 20174 1162 20230
rect 1188 20174 1244 20230
rect 1270 20174 1326 20230
rect 1352 20174 1408 20230
rect 1434 20174 1490 20230
rect 1516 20174 1572 20230
rect 1598 20174 1654 20230
rect 1106 20093 1162 20149
rect 1188 20093 1244 20149
rect 1270 20093 1326 20149
rect 1352 20093 1408 20149
rect 1434 20093 1490 20149
rect 1516 20093 1572 20149
rect 1598 20093 1654 20149
rect 1106 20012 1162 20068
rect 1188 20012 1244 20068
rect 1270 20012 1326 20068
rect 1352 20012 1408 20068
rect 1434 20012 1490 20068
rect 1516 20012 1572 20068
rect 1598 20012 1654 20068
rect 1106 19931 1162 19987
rect 1188 19931 1244 19987
rect 1270 19931 1326 19987
rect 1352 19931 1408 19987
rect 1434 19931 1490 19987
rect 1516 19931 1572 19987
rect 1598 19931 1654 19987
rect 1106 19850 1162 19906
rect 1188 19850 1244 19906
rect 1270 19850 1326 19906
rect 1352 19850 1408 19906
rect 1434 19850 1490 19906
rect 1516 19850 1572 19906
rect 1598 19850 1654 19906
rect 1106 19769 1162 19825
rect 1188 19769 1244 19825
rect 1270 19769 1326 19825
rect 1352 19769 1408 19825
rect 1434 19769 1490 19825
rect 1516 19769 1572 19825
rect 1598 19769 1654 19825
rect 1106 19688 1162 19744
rect 1188 19688 1244 19744
rect 1270 19688 1326 19744
rect 1352 19688 1408 19744
rect 1434 19688 1490 19744
rect 1516 19688 1572 19744
rect 1598 19688 1654 19744
rect 1106 19607 1162 19663
rect 1188 19607 1244 19663
rect 1270 19607 1326 19663
rect 1352 19607 1408 19663
rect 1434 19607 1490 19663
rect 1516 19607 1572 19663
rect 1598 19607 1654 19663
rect 1106 19526 1162 19582
rect 1188 19526 1244 19582
rect 1270 19526 1326 19582
rect 1352 19526 1408 19582
rect 1434 19526 1490 19582
rect 1516 19526 1572 19582
rect 1598 19526 1654 19582
rect 1106 19445 1162 19501
rect 1188 19445 1244 19501
rect 1270 19445 1326 19501
rect 1352 19445 1408 19501
rect 1434 19445 1490 19501
rect 1516 19445 1572 19501
rect 1598 19445 1654 19501
rect 1106 19364 1162 19420
rect 1188 19364 1244 19420
rect 1270 19364 1326 19420
rect 1352 19364 1408 19420
rect 1434 19364 1490 19420
rect 1516 19364 1572 19420
rect 1598 19364 1654 19420
rect 1106 19283 1162 19339
rect 1188 19283 1244 19339
rect 1270 19283 1326 19339
rect 1352 19283 1408 19339
rect 1434 19283 1490 19339
rect 1516 19283 1572 19339
rect 1598 19283 1654 19339
rect 1106 19202 1162 19258
rect 1188 19202 1244 19258
rect 1270 19202 1326 19258
rect 1352 19202 1408 19258
rect 1434 19202 1490 19258
rect 1516 19202 1572 19258
rect 1598 19202 1654 19258
rect 1106 19121 1162 19177
rect 1188 19121 1244 19177
rect 1270 19121 1326 19177
rect 1352 19121 1408 19177
rect 1434 19121 1490 19177
rect 1516 19121 1572 19177
rect 1598 19121 1654 19177
rect 1106 19040 1162 19096
rect 1188 19040 1244 19096
rect 1270 19040 1326 19096
rect 1352 19040 1408 19096
rect 1434 19040 1490 19096
rect 1516 19040 1572 19096
rect 1598 19040 1654 19096
rect 2910 20494 2966 20550
rect 2992 20494 3048 20550
rect 3074 20494 3130 20550
rect 3156 20494 3212 20550
rect 3238 20494 3294 20550
rect 3320 20494 3376 20550
rect 3402 20494 3458 20550
rect 2910 20414 2966 20470
rect 2992 20414 3048 20470
rect 3074 20414 3130 20470
rect 3156 20414 3212 20470
rect 3238 20414 3294 20470
rect 3320 20414 3376 20470
rect 3402 20414 3458 20470
rect 2910 20334 2966 20390
rect 2992 20334 3048 20390
rect 3074 20334 3130 20390
rect 3156 20334 3212 20390
rect 3238 20334 3294 20390
rect 3320 20334 3376 20390
rect 3402 20334 3458 20390
rect 2910 20254 2966 20310
rect 2992 20254 3048 20310
rect 3074 20254 3130 20310
rect 3156 20254 3212 20310
rect 3238 20254 3294 20310
rect 3320 20254 3376 20310
rect 3402 20254 3458 20310
rect 2910 20174 2966 20230
rect 2992 20174 3048 20230
rect 3074 20174 3130 20230
rect 3156 20174 3212 20230
rect 3238 20174 3294 20230
rect 3320 20174 3376 20230
rect 3402 20174 3458 20230
rect 2910 20093 2966 20149
rect 2992 20093 3048 20149
rect 3074 20093 3130 20149
rect 3156 20093 3212 20149
rect 3238 20093 3294 20149
rect 3320 20093 3376 20149
rect 3402 20093 3458 20149
rect 2910 20012 2966 20068
rect 2992 20012 3048 20068
rect 3074 20012 3130 20068
rect 3156 20012 3212 20068
rect 3238 20012 3294 20068
rect 3320 20012 3376 20068
rect 3402 20012 3458 20068
rect 2910 19931 2966 19987
rect 2992 19931 3048 19987
rect 3074 19931 3130 19987
rect 3156 19931 3212 19987
rect 3238 19931 3294 19987
rect 3320 19931 3376 19987
rect 3402 19931 3458 19987
rect 2910 19850 2966 19906
rect 2992 19850 3048 19906
rect 3074 19850 3130 19906
rect 3156 19850 3212 19906
rect 3238 19850 3294 19906
rect 3320 19850 3376 19906
rect 3402 19850 3458 19906
rect 2910 19769 2966 19825
rect 2992 19769 3048 19825
rect 3074 19769 3130 19825
rect 3156 19769 3212 19825
rect 3238 19769 3294 19825
rect 3320 19769 3376 19825
rect 3402 19769 3458 19825
rect 2910 19688 2966 19744
rect 2992 19688 3048 19744
rect 3074 19688 3130 19744
rect 3156 19688 3212 19744
rect 3238 19688 3294 19744
rect 3320 19688 3376 19744
rect 3402 19688 3458 19744
rect 2910 19607 2966 19663
rect 2992 19607 3048 19663
rect 3074 19607 3130 19663
rect 3156 19607 3212 19663
rect 3238 19607 3294 19663
rect 3320 19607 3376 19663
rect 3402 19607 3458 19663
rect 2910 19526 2966 19582
rect 2992 19526 3048 19582
rect 3074 19526 3130 19582
rect 3156 19526 3212 19582
rect 3238 19526 3294 19582
rect 3320 19526 3376 19582
rect 3402 19526 3458 19582
rect 2910 19445 2966 19501
rect 2992 19445 3048 19501
rect 3074 19445 3130 19501
rect 3156 19445 3212 19501
rect 3238 19445 3294 19501
rect 3320 19445 3376 19501
rect 3402 19445 3458 19501
rect 2910 19364 2966 19420
rect 2992 19364 3048 19420
rect 3074 19364 3130 19420
rect 3156 19364 3212 19420
rect 3238 19364 3294 19420
rect 3320 19364 3376 19420
rect 3402 19364 3458 19420
rect 2910 19283 2966 19339
rect 2992 19283 3048 19339
rect 3074 19283 3130 19339
rect 3156 19283 3212 19339
rect 3238 19283 3294 19339
rect 3320 19283 3376 19339
rect 3402 19283 3458 19339
rect 2910 19202 2966 19258
rect 2992 19202 3048 19258
rect 3074 19202 3130 19258
rect 3156 19202 3212 19258
rect 3238 19202 3294 19258
rect 3320 19202 3376 19258
rect 3402 19202 3458 19258
rect 2910 19121 2966 19177
rect 2992 19121 3048 19177
rect 3074 19121 3130 19177
rect 3156 19121 3212 19177
rect 3238 19121 3294 19177
rect 3320 19121 3376 19177
rect 3402 19121 3458 19177
rect 2910 19040 2966 19096
rect 2992 19040 3048 19096
rect 3074 19040 3130 19096
rect 3156 19040 3212 19096
rect 3238 19040 3294 19096
rect 3320 19040 3376 19096
rect 3402 19040 3458 19096
rect 4708 20494 4764 20550
rect 4790 20494 4846 20550
rect 4872 20494 4928 20550
rect 4954 20494 5010 20550
rect 5036 20494 5092 20550
rect 5118 20494 5174 20550
rect 5200 20494 5256 20550
rect 4708 20414 4764 20470
rect 4790 20414 4846 20470
rect 4872 20414 4928 20470
rect 4954 20414 5010 20470
rect 5036 20414 5092 20470
rect 5118 20414 5174 20470
rect 5200 20414 5256 20470
rect 4708 20334 4764 20390
rect 4790 20334 4846 20390
rect 4872 20334 4928 20390
rect 4954 20334 5010 20390
rect 5036 20334 5092 20390
rect 5118 20334 5174 20390
rect 5200 20334 5256 20390
rect 4708 20254 4764 20310
rect 4790 20254 4846 20310
rect 4872 20254 4928 20310
rect 4954 20254 5010 20310
rect 5036 20254 5092 20310
rect 5118 20254 5174 20310
rect 5200 20254 5256 20310
rect 4708 20174 4764 20230
rect 4790 20174 4846 20230
rect 4872 20174 4928 20230
rect 4954 20174 5010 20230
rect 5036 20174 5092 20230
rect 5118 20174 5174 20230
rect 5200 20174 5256 20230
rect 4708 20093 4764 20149
rect 4790 20093 4846 20149
rect 4872 20093 4928 20149
rect 4954 20093 5010 20149
rect 5036 20093 5092 20149
rect 5118 20093 5174 20149
rect 5200 20093 5256 20149
rect 4708 20012 4764 20068
rect 4790 20012 4846 20068
rect 4872 20012 4928 20068
rect 4954 20012 5010 20068
rect 5036 20012 5092 20068
rect 5118 20012 5174 20068
rect 5200 20012 5256 20068
rect 4708 19931 4764 19987
rect 4790 19931 4846 19987
rect 4872 19931 4928 19987
rect 4954 19931 5010 19987
rect 5036 19931 5092 19987
rect 5118 19931 5174 19987
rect 5200 19931 5256 19987
rect 4708 19850 4764 19906
rect 4790 19850 4846 19906
rect 4872 19850 4928 19906
rect 4954 19850 5010 19906
rect 5036 19850 5092 19906
rect 5118 19850 5174 19906
rect 5200 19850 5256 19906
rect 4708 19769 4764 19825
rect 4790 19769 4846 19825
rect 4872 19769 4928 19825
rect 4954 19769 5010 19825
rect 5036 19769 5092 19825
rect 5118 19769 5174 19825
rect 5200 19769 5256 19825
rect 4708 19688 4764 19744
rect 4790 19688 4846 19744
rect 4872 19688 4928 19744
rect 4954 19688 5010 19744
rect 5036 19688 5092 19744
rect 5118 19688 5174 19744
rect 5200 19688 5256 19744
rect 4708 19607 4764 19663
rect 4790 19607 4846 19663
rect 4872 19607 4928 19663
rect 4954 19607 5010 19663
rect 5036 19607 5092 19663
rect 5118 19607 5174 19663
rect 5200 19607 5256 19663
rect 4708 19526 4764 19582
rect 4790 19526 4846 19582
rect 4872 19526 4928 19582
rect 4954 19526 5010 19582
rect 5036 19526 5092 19582
rect 5118 19526 5174 19582
rect 5200 19526 5256 19582
rect 4708 19445 4764 19501
rect 4790 19445 4846 19501
rect 4872 19445 4928 19501
rect 4954 19445 5010 19501
rect 5036 19445 5092 19501
rect 5118 19445 5174 19501
rect 5200 19445 5256 19501
rect 4708 19364 4764 19420
rect 4790 19364 4846 19420
rect 4872 19364 4928 19420
rect 4954 19364 5010 19420
rect 5036 19364 5092 19420
rect 5118 19364 5174 19420
rect 5200 19364 5256 19420
rect 4708 19283 4764 19339
rect 4790 19283 4846 19339
rect 4872 19283 4928 19339
rect 4954 19283 5010 19339
rect 5036 19283 5092 19339
rect 5118 19283 5174 19339
rect 5200 19283 5256 19339
rect 4708 19202 4764 19258
rect 4790 19202 4846 19258
rect 4872 19202 4928 19258
rect 4954 19202 5010 19258
rect 5036 19202 5092 19258
rect 5118 19202 5174 19258
rect 5200 19202 5256 19258
rect 4708 19121 4764 19177
rect 4790 19121 4846 19177
rect 4872 19121 4928 19177
rect 4954 19121 5010 19177
rect 5036 19121 5092 19177
rect 5118 19121 5174 19177
rect 5200 19121 5256 19177
rect 4708 19040 4764 19096
rect 4790 19040 4846 19096
rect 4872 19040 4928 19096
rect 4954 19040 5010 19096
rect 5036 19040 5092 19096
rect 5118 19040 5174 19096
rect 5200 19040 5256 19096
rect 6378 20174 6754 20550
rect 6378 20093 6434 20149
rect 6458 20093 6514 20149
rect 6538 20093 6594 20149
rect 6618 20093 6674 20149
rect 6698 20093 6754 20149
rect 6378 20012 6434 20068
rect 6458 20012 6514 20068
rect 6538 20012 6594 20068
rect 6618 20012 6674 20068
rect 6698 20012 6754 20068
rect 6378 19931 6434 19987
rect 6458 19931 6514 19987
rect 6538 19931 6594 19987
rect 6618 19931 6674 19987
rect 6698 19931 6754 19987
rect 6378 19850 6434 19906
rect 6458 19850 6514 19906
rect 6538 19850 6594 19906
rect 6618 19850 6674 19906
rect 6698 19850 6754 19906
rect 6378 19769 6434 19825
rect 6458 19769 6514 19825
rect 6538 19769 6594 19825
rect 6618 19769 6674 19825
rect 6698 19769 6754 19825
rect 6378 19688 6434 19744
rect 6458 19688 6514 19744
rect 6538 19688 6594 19744
rect 6618 19688 6674 19744
rect 6698 19688 6754 19744
rect 6378 19607 6434 19663
rect 6458 19607 6514 19663
rect 6538 19607 6594 19663
rect 6618 19607 6674 19663
rect 6698 19607 6754 19663
rect 6378 19526 6434 19582
rect 6458 19526 6514 19582
rect 6538 19526 6594 19582
rect 6618 19526 6674 19582
rect 6698 19526 6754 19582
rect 6378 19445 6434 19501
rect 6458 19445 6514 19501
rect 6538 19445 6594 19501
rect 6618 19445 6674 19501
rect 6698 19445 6754 19501
rect 6378 19364 6434 19420
rect 6458 19364 6514 19420
rect 6538 19364 6594 19420
rect 6618 19364 6674 19420
rect 6698 19364 6754 19420
rect 6378 19283 6434 19339
rect 6458 19283 6514 19339
rect 6538 19283 6594 19339
rect 6618 19283 6674 19339
rect 6698 19283 6754 19339
rect 6378 19202 6434 19258
rect 6458 19202 6514 19258
rect 6538 19202 6594 19258
rect 6618 19202 6674 19258
rect 6698 19202 6754 19258
rect 6378 19121 6434 19177
rect 6458 19121 6514 19177
rect 6538 19121 6594 19177
rect 6618 19121 6674 19177
rect 6698 19121 6754 19177
rect 6378 19040 6434 19096
rect 6458 19040 6514 19096
rect 6538 19040 6594 19096
rect 6618 19040 6674 19096
rect 6698 19040 6754 19096
rect 8067 20500 8123 20556
rect 8169 20500 8225 20556
rect 8271 20500 8327 20556
rect 8067 20419 8123 20475
rect 8169 20419 8225 20475
rect 8271 20419 8327 20475
rect 8067 20338 8123 20394
rect 8169 20338 8225 20394
rect 8271 20338 8327 20394
rect 8067 20257 8123 20313
rect 8169 20257 8225 20313
rect 8271 20257 8327 20313
rect 8067 20176 8123 20232
rect 8169 20176 8225 20232
rect 8271 20176 8327 20232
rect 8067 20095 8123 20151
rect 8169 20095 8225 20151
rect 8271 20095 8327 20151
rect 8067 20014 8123 20070
rect 8169 20014 8225 20070
rect 8271 20014 8327 20070
rect 8067 19933 8123 19989
rect 8169 19933 8225 19989
rect 8271 19933 8327 19989
rect 8067 19852 8123 19908
rect 8169 19852 8225 19908
rect 8271 19852 8327 19908
rect 8067 19771 8123 19827
rect 8169 19771 8225 19827
rect 8271 19771 8327 19827
rect 8067 19689 8123 19745
rect 8169 19689 8225 19745
rect 8271 19689 8327 19745
rect 8067 19607 8123 19663
rect 8169 19607 8225 19663
rect 8271 19607 8327 19663
rect 8067 19525 8123 19581
rect 8169 19525 8225 19581
rect 8271 19525 8327 19581
rect 8067 19443 8123 19499
rect 8169 19443 8225 19499
rect 8271 19443 8327 19499
rect 8067 19361 8123 19417
rect 8169 19361 8225 19417
rect 8271 19361 8327 19417
rect 8067 19279 8123 19335
rect 8169 19279 8225 19335
rect 8271 19279 8327 19335
rect 8067 19197 8123 19253
rect 8169 19197 8225 19253
rect 8271 19197 8327 19253
rect 8067 19115 8123 19171
rect 8169 19115 8225 19171
rect 8271 19115 8327 19171
rect 8067 19033 8123 19089
rect 8169 19033 8225 19089
rect 8271 19033 8327 19089
rect 8894 20500 8950 20556
rect 8990 20500 9046 20556
rect 9086 20500 9142 20556
rect 8894 20419 8950 20475
rect 8990 20419 9046 20475
rect 9086 20419 9142 20475
rect 8894 20338 8950 20394
rect 8990 20338 9046 20394
rect 9086 20338 9142 20394
rect 8894 20257 8950 20313
rect 8990 20257 9046 20313
rect 9086 20257 9142 20313
rect 8894 20176 8950 20232
rect 8990 20176 9046 20232
rect 9086 20176 9142 20232
rect 8894 20095 8950 20151
rect 8990 20095 9046 20151
rect 9086 20095 9142 20151
rect 8894 20014 8950 20070
rect 8990 20014 9046 20070
rect 9086 20014 9142 20070
rect 8894 19933 8950 19989
rect 8990 19933 9046 19989
rect 9086 19933 9142 19989
rect 8894 19852 8950 19908
rect 8990 19852 9046 19908
rect 9086 19852 9142 19908
rect 8894 19771 8950 19827
rect 8990 19771 9046 19827
rect 9086 19771 9142 19827
rect 8894 19689 8950 19745
rect 8990 19689 9046 19745
rect 9086 19689 9142 19745
rect 8894 19607 8950 19663
rect 8990 19607 9046 19663
rect 9086 19607 9142 19663
rect 8894 19525 8950 19581
rect 8990 19525 9046 19581
rect 9086 19525 9142 19581
rect 8894 19443 8950 19499
rect 8990 19443 9046 19499
rect 9086 19443 9142 19499
rect 8894 19361 8950 19417
rect 8990 19361 9046 19417
rect 9086 19361 9142 19417
rect 8894 19279 8950 19335
rect 8990 19279 9046 19335
rect 9086 19279 9142 19335
rect 8894 19197 8950 19253
rect 8990 19197 9046 19253
rect 9086 19197 9142 19253
rect 8894 19115 8950 19171
rect 8990 19115 9046 19171
rect 9086 19115 9142 19171
rect 8894 19033 8950 19089
rect 8990 19033 9046 19089
rect 9086 19033 9142 19089
rect 10126 20494 10182 20550
rect 10208 20494 10264 20550
rect 10290 20494 10346 20550
rect 10372 20494 10428 20550
rect 10454 20494 10510 20550
rect 10536 20494 10592 20550
rect 10618 20494 10674 20550
rect 10126 20411 10182 20467
rect 10208 20411 10264 20467
rect 10290 20411 10346 20467
rect 10372 20411 10428 20467
rect 10454 20411 10510 20467
rect 10536 20411 10592 20467
rect 10618 20411 10674 20467
rect 10126 20328 10182 20384
rect 10208 20328 10264 20384
rect 10290 20328 10346 20384
rect 10372 20328 10428 20384
rect 10454 20328 10510 20384
rect 10536 20328 10592 20384
rect 10618 20328 10674 20384
rect 10126 20245 10182 20301
rect 10208 20245 10264 20301
rect 10290 20245 10346 20301
rect 10372 20245 10428 20301
rect 10454 20245 10510 20301
rect 10536 20245 10592 20301
rect 10618 20245 10674 20301
rect 10126 20161 10182 20217
rect 10208 20161 10264 20217
rect 10290 20161 10346 20217
rect 10372 20161 10428 20217
rect 10454 20161 10510 20217
rect 10536 20161 10592 20217
rect 10618 20161 10674 20217
rect 10126 20077 10182 20133
rect 10208 20077 10264 20133
rect 10290 20077 10346 20133
rect 10372 20077 10428 20133
rect 10454 20077 10510 20133
rect 10536 20077 10592 20133
rect 10618 20077 10674 20133
rect 10126 19993 10182 20049
rect 10208 19993 10264 20049
rect 10290 19993 10346 20049
rect 10372 19993 10428 20049
rect 10454 19993 10510 20049
rect 10536 19993 10592 20049
rect 10618 19993 10674 20049
rect 10126 19909 10182 19965
rect 10208 19909 10264 19965
rect 10290 19909 10346 19965
rect 10372 19909 10428 19965
rect 10454 19909 10510 19965
rect 10536 19909 10592 19965
rect 10618 19909 10674 19965
rect 10126 19825 10182 19881
rect 10208 19825 10264 19881
rect 10290 19825 10346 19881
rect 10372 19825 10428 19881
rect 10454 19825 10510 19881
rect 10536 19825 10592 19881
rect 10618 19825 10674 19881
rect 10126 19741 10182 19797
rect 10208 19741 10264 19797
rect 10290 19741 10346 19797
rect 10372 19741 10428 19797
rect 10454 19741 10510 19797
rect 10536 19741 10592 19797
rect 10618 19741 10674 19797
rect 10126 19657 10182 19713
rect 10208 19657 10264 19713
rect 10290 19657 10346 19713
rect 10372 19657 10428 19713
rect 10454 19657 10510 19713
rect 10536 19657 10592 19713
rect 10618 19657 10674 19713
rect 10126 19573 10182 19629
rect 10208 19573 10264 19629
rect 10290 19573 10346 19629
rect 10372 19573 10428 19629
rect 10454 19573 10510 19629
rect 10536 19573 10592 19629
rect 10618 19573 10674 19629
rect 10126 19489 10182 19545
rect 10208 19489 10264 19545
rect 10290 19489 10346 19545
rect 10372 19489 10428 19545
rect 10454 19489 10510 19545
rect 10536 19489 10592 19545
rect 10618 19489 10674 19545
rect 10126 19405 10182 19461
rect 10208 19405 10264 19461
rect 10290 19405 10346 19461
rect 10372 19405 10428 19461
rect 10454 19405 10510 19461
rect 10536 19405 10592 19461
rect 10618 19405 10674 19461
rect 10126 19321 10182 19377
rect 10208 19321 10264 19377
rect 10290 19321 10346 19377
rect 10372 19321 10428 19377
rect 10454 19321 10510 19377
rect 10536 19321 10592 19377
rect 10618 19321 10674 19377
rect 10126 19237 10182 19293
rect 10208 19237 10264 19293
rect 10290 19237 10346 19293
rect 10372 19237 10428 19293
rect 10454 19237 10510 19293
rect 10536 19237 10592 19293
rect 10618 19237 10674 19293
rect 10126 19153 10182 19209
rect 10208 19153 10264 19209
rect 10290 19153 10346 19209
rect 10372 19153 10428 19209
rect 10454 19153 10510 19209
rect 10536 19153 10592 19209
rect 10618 19153 10674 19209
rect 10126 19069 10182 19125
rect 10208 19069 10264 19125
rect 10290 19069 10346 19125
rect 10372 19069 10428 19125
rect 10454 19069 10510 19125
rect 10536 19069 10592 19125
rect 10618 19069 10674 19125
rect 11927 20494 11983 20550
rect 12009 20494 12065 20550
rect 12091 20494 12147 20550
rect 12173 20494 12229 20550
rect 12255 20494 12311 20550
rect 12337 20494 12393 20550
rect 12419 20494 12475 20550
rect 11927 20411 11983 20467
rect 12009 20411 12065 20467
rect 12091 20411 12147 20467
rect 12173 20411 12229 20467
rect 12255 20411 12311 20467
rect 12337 20411 12393 20467
rect 12419 20411 12475 20467
rect 11927 20328 11983 20384
rect 12009 20328 12065 20384
rect 12091 20328 12147 20384
rect 12173 20328 12229 20384
rect 12255 20328 12311 20384
rect 12337 20328 12393 20384
rect 12419 20328 12475 20384
rect 11927 20245 11983 20301
rect 12009 20245 12065 20301
rect 12091 20245 12147 20301
rect 12173 20245 12229 20301
rect 12255 20245 12311 20301
rect 12337 20245 12393 20301
rect 12419 20245 12475 20301
rect 11927 20161 11983 20217
rect 12009 20161 12065 20217
rect 12091 20161 12147 20217
rect 12173 20161 12229 20217
rect 12255 20161 12311 20217
rect 12337 20161 12393 20217
rect 12419 20161 12475 20217
rect 11927 20077 11983 20133
rect 12009 20077 12065 20133
rect 12091 20077 12147 20133
rect 12173 20077 12229 20133
rect 12255 20077 12311 20133
rect 12337 20077 12393 20133
rect 12419 20077 12475 20133
rect 11927 19993 11983 20049
rect 12009 19993 12065 20049
rect 12091 19993 12147 20049
rect 12173 19993 12229 20049
rect 12255 19993 12311 20049
rect 12337 19993 12393 20049
rect 12419 19993 12475 20049
rect 11927 19909 11983 19965
rect 12009 19909 12065 19965
rect 12091 19909 12147 19965
rect 12173 19909 12229 19965
rect 12255 19909 12311 19965
rect 12337 19909 12393 19965
rect 12419 19909 12475 19965
rect 11927 19825 11983 19881
rect 12009 19825 12065 19881
rect 12091 19825 12147 19881
rect 12173 19825 12229 19881
rect 12255 19825 12311 19881
rect 12337 19825 12393 19881
rect 12419 19825 12475 19881
rect 11927 19741 11983 19797
rect 12009 19741 12065 19797
rect 12091 19741 12147 19797
rect 12173 19741 12229 19797
rect 12255 19741 12311 19797
rect 12337 19741 12393 19797
rect 12419 19741 12475 19797
rect 11927 19657 11983 19713
rect 12009 19657 12065 19713
rect 12091 19657 12147 19713
rect 12173 19657 12229 19713
rect 12255 19657 12311 19713
rect 12337 19657 12393 19713
rect 12419 19657 12475 19713
rect 11927 19573 11983 19629
rect 12009 19573 12065 19629
rect 12091 19573 12147 19629
rect 12173 19573 12229 19629
rect 12255 19573 12311 19629
rect 12337 19573 12393 19629
rect 12419 19573 12475 19629
rect 11927 19489 11983 19545
rect 12009 19489 12065 19545
rect 12091 19489 12147 19545
rect 12173 19489 12229 19545
rect 12255 19489 12311 19545
rect 12337 19489 12393 19545
rect 12419 19489 12475 19545
rect 11927 19405 11983 19461
rect 12009 19405 12065 19461
rect 12091 19405 12147 19461
rect 12173 19405 12229 19461
rect 12255 19405 12311 19461
rect 12337 19405 12393 19461
rect 12419 19405 12475 19461
rect 11927 19321 11983 19377
rect 12009 19321 12065 19377
rect 12091 19321 12147 19377
rect 12173 19321 12229 19377
rect 12255 19321 12311 19377
rect 12337 19321 12393 19377
rect 12419 19321 12475 19377
rect 11927 19237 11983 19293
rect 12009 19237 12065 19293
rect 12091 19237 12147 19293
rect 12173 19237 12229 19293
rect 12255 19237 12311 19293
rect 12337 19237 12393 19293
rect 12419 19237 12475 19293
rect 11927 19153 11983 19209
rect 12009 19153 12065 19209
rect 12091 19153 12147 19209
rect 12173 19153 12229 19209
rect 12255 19153 12311 19209
rect 12337 19153 12393 19209
rect 12419 19153 12475 19209
rect 11927 19069 11983 19125
rect 12009 19069 12065 19125
rect 12091 19069 12147 19125
rect 12173 19069 12229 19125
rect 12255 19069 12311 19125
rect 12337 19069 12393 19125
rect 12419 19069 12475 19125
rect 2906 12990 2962 13046
rect 2990 12990 3046 13046
rect 3074 12990 3130 13046
rect 3158 12990 3214 13046
rect 3242 12990 3298 13046
rect 3326 12990 3382 13046
rect 3410 12990 3466 13046
rect -714 12777 -658 12833
rect -626 12777 -570 12833
rect -538 12777 -482 12833
rect -450 12777 -394 12833
rect -362 12777 -306 12833
rect -274 12777 -218 12833
rect -186 12777 -130 12833
rect -714 12697 -658 12753
rect -626 12697 -570 12753
rect -538 12697 -482 12753
rect -450 12697 -394 12753
rect -362 12697 -306 12753
rect -274 12697 -218 12753
rect -186 12697 -130 12753
rect -714 12617 -658 12673
rect -626 12617 -570 12673
rect -538 12617 -482 12673
rect -450 12617 -394 12673
rect -362 12617 -306 12673
rect -274 12617 -218 12673
rect -186 12617 -130 12673
rect -714 12537 -658 12593
rect -626 12537 -570 12593
rect -538 12537 -482 12593
rect -450 12537 -394 12593
rect -362 12537 -306 12593
rect -274 12537 -218 12593
rect -186 12537 -130 12593
rect -714 12457 -658 12513
rect -626 12457 -570 12513
rect -538 12457 -482 12513
rect -450 12457 -394 12513
rect -362 12457 -306 12513
rect -274 12457 -218 12513
rect -186 12457 -130 12513
rect 1115 12871 1171 12927
rect 1211 12871 1267 12927
rect 1307 12871 1363 12927
rect 1402 12871 1458 12927
rect 1497 12871 1553 12927
rect 1592 12871 1648 12927
rect 1115 12787 1171 12843
rect 1211 12787 1267 12843
rect 1307 12787 1363 12843
rect 1402 12787 1458 12843
rect 1497 12787 1553 12843
rect 1592 12787 1648 12843
rect 1115 12703 1171 12759
rect 1211 12703 1267 12759
rect 1307 12703 1363 12759
rect 1402 12703 1458 12759
rect 1497 12703 1553 12759
rect 1592 12703 1648 12759
rect 1115 12619 1171 12675
rect 1211 12619 1267 12675
rect 1307 12619 1363 12675
rect 1402 12619 1458 12675
rect 1497 12619 1553 12675
rect 1592 12619 1648 12675
rect 1115 12535 1171 12591
rect 1211 12535 1267 12591
rect 1307 12535 1363 12591
rect 1402 12535 1458 12591
rect 1497 12535 1553 12591
rect 1592 12535 1648 12591
rect 1115 12451 1171 12507
rect 1211 12451 1267 12507
rect 1307 12451 1363 12507
rect 1402 12451 1458 12507
rect 1497 12451 1553 12507
rect 1592 12451 1648 12507
rect 2906 12901 2962 12957
rect 2990 12901 3046 12957
rect 3074 12901 3130 12957
rect 3158 12901 3214 12957
rect 3242 12901 3298 12957
rect 3326 12901 3382 12957
rect 3410 12901 3466 12957
rect 2906 12812 2962 12868
rect 2990 12812 3046 12868
rect 3074 12812 3130 12868
rect 3158 12812 3214 12868
rect 3242 12812 3298 12868
rect 3326 12812 3382 12868
rect 3410 12812 3466 12868
rect 2906 12723 2962 12779
rect 2990 12723 3046 12779
rect 3074 12723 3130 12779
rect 3158 12723 3214 12779
rect 3242 12723 3298 12779
rect 3326 12723 3382 12779
rect 3410 12723 3466 12779
rect 2906 12634 2962 12690
rect 2990 12634 3046 12690
rect 3074 12634 3130 12690
rect 3158 12634 3214 12690
rect 3242 12634 3298 12690
rect 3326 12634 3382 12690
rect 3410 12634 3466 12690
rect 2906 12545 2962 12601
rect 2990 12545 3046 12601
rect 3074 12545 3130 12601
rect 3158 12545 3214 12601
rect 3242 12545 3298 12601
rect 3326 12545 3382 12601
rect 3410 12545 3466 12601
rect 2906 12455 2962 12511
rect 2990 12455 3046 12511
rect 3074 12455 3130 12511
rect 3158 12455 3214 12511
rect 3242 12455 3298 12511
rect 3326 12455 3382 12511
rect 3410 12455 3466 12511
rect 4704 12990 4760 13046
rect 4788 12990 4844 13046
rect 4872 12990 4928 13046
rect 4956 12990 5012 13046
rect 5040 12990 5096 13046
rect 5124 12990 5180 13046
rect 5208 12990 5264 13046
rect 4704 12901 4760 12957
rect 4788 12901 4844 12957
rect 4872 12901 4928 12957
rect 4956 12901 5012 12957
rect 5040 12901 5096 12957
rect 5124 12901 5180 12957
rect 5208 12901 5264 12957
rect 4704 12812 4760 12868
rect 4788 12812 4844 12868
rect 4872 12812 4928 12868
rect 4956 12812 5012 12868
rect 5040 12812 5096 12868
rect 5124 12812 5180 12868
rect 5208 12812 5264 12868
rect 4704 12723 4760 12779
rect 4788 12723 4844 12779
rect 4872 12723 4928 12779
rect 4956 12723 5012 12779
rect 5040 12723 5096 12779
rect 5124 12723 5180 12779
rect 5208 12723 5264 12779
rect 4704 12634 4760 12690
rect 4788 12634 4844 12690
rect 4872 12634 4928 12690
rect 4956 12634 5012 12690
rect 5040 12634 5096 12690
rect 5124 12634 5180 12690
rect 5208 12634 5264 12690
rect 4704 12545 4760 12601
rect 4788 12545 4844 12601
rect 4872 12545 4928 12601
rect 4956 12545 5012 12601
rect 5040 12545 5096 12601
rect 5124 12545 5180 12601
rect 5208 12545 5264 12601
rect 4704 12455 4760 12511
rect 4788 12455 4844 12511
rect 4872 12455 4928 12511
rect 4956 12455 5012 12511
rect 5040 12455 5096 12511
rect 5124 12455 5180 12511
rect 5208 12455 5264 12511
rect 6511 12990 6567 13046
rect 6595 12990 6651 13046
rect 6679 12990 6735 13046
rect 6763 12990 6819 13046
rect 6847 12990 6903 13046
rect 6931 12990 6987 13046
rect 7015 12990 7071 13046
rect 6511 12901 6567 12957
rect 6595 12901 6651 12957
rect 6679 12901 6735 12957
rect 6763 12901 6819 12957
rect 6847 12901 6903 12957
rect 6931 12901 6987 12957
rect 7015 12901 7071 12957
rect 6511 12812 6567 12868
rect 6595 12812 6651 12868
rect 6679 12812 6735 12868
rect 6763 12812 6819 12868
rect 6847 12812 6903 12868
rect 6931 12812 6987 12868
rect 7015 12812 7071 12868
rect 6511 12723 6567 12779
rect 6595 12723 6651 12779
rect 6679 12723 6735 12779
rect 6763 12723 6819 12779
rect 6847 12723 6903 12779
rect 6931 12723 6987 12779
rect 7015 12723 7071 12779
rect 6511 12634 6567 12690
rect 6595 12634 6651 12690
rect 6679 12634 6735 12690
rect 6763 12634 6819 12690
rect 6847 12634 6903 12690
rect 6931 12634 6987 12690
rect 7015 12634 7071 12690
rect 6511 12545 6567 12601
rect 6595 12545 6651 12601
rect 6679 12545 6735 12601
rect 6763 12545 6819 12601
rect 6847 12545 6903 12601
rect 6931 12545 6987 12601
rect 7015 12545 7071 12601
rect 6511 12455 6567 12511
rect 6595 12455 6651 12511
rect 6679 12455 6735 12511
rect 6763 12455 6819 12511
rect 6847 12455 6903 12511
rect 6931 12455 6987 12511
rect 7015 12455 7071 12511
rect 8324 12989 8380 13045
rect 8408 12989 8464 13045
rect 8492 12989 8548 13045
rect 8576 12989 8632 13045
rect 8660 12989 8716 13045
rect 8744 12989 8800 13045
rect 8828 12989 8884 13045
rect 8324 12909 8380 12965
rect 8408 12909 8464 12965
rect 8492 12909 8548 12965
rect 8576 12909 8632 12965
rect 8660 12909 8716 12965
rect 8744 12909 8800 12965
rect 8828 12909 8884 12965
rect 8324 12829 8380 12885
rect 8408 12829 8464 12885
rect 8492 12829 8548 12885
rect 8576 12829 8632 12885
rect 8660 12829 8716 12885
rect 8744 12829 8800 12885
rect 8828 12829 8884 12885
rect 8324 12749 8380 12805
rect 8408 12749 8464 12805
rect 8492 12749 8548 12805
rect 8576 12749 8632 12805
rect 8660 12749 8716 12805
rect 8744 12749 8800 12805
rect 8828 12749 8884 12805
rect 8324 12669 8380 12725
rect 8408 12669 8464 12725
rect 8492 12669 8548 12725
rect 8576 12669 8632 12725
rect 8660 12669 8716 12725
rect 8744 12669 8800 12725
rect 8828 12669 8884 12725
rect 8324 12589 8380 12645
rect 8408 12589 8464 12645
rect 8492 12589 8548 12645
rect 8576 12589 8632 12645
rect 8660 12589 8716 12645
rect 8744 12589 8800 12645
rect 8828 12589 8884 12645
rect 8324 12509 8380 12565
rect 8408 12509 8464 12565
rect 8492 12509 8548 12565
rect 8576 12509 8632 12565
rect 8660 12509 8716 12565
rect 8744 12509 8800 12565
rect 8828 12509 8884 12565
rect -714 12377 -658 12433
rect -626 12377 -570 12433
rect -538 12377 -482 12433
rect -450 12377 -394 12433
rect -362 12377 -306 12433
rect -274 12377 -218 12433
rect -186 12377 -130 12433
rect -714 12297 -658 12353
rect -626 12297 -570 12353
rect -538 12297 -482 12353
rect -450 12297 -394 12353
rect -362 12297 -306 12353
rect -274 12297 -218 12353
rect -186 12297 -130 12353
rect -714 12217 -658 12273
rect -626 12217 -570 12273
rect -538 12217 -482 12273
rect -450 12217 -394 12273
rect -362 12217 -306 12273
rect -274 12217 -218 12273
rect -186 12217 -130 12273
rect -2511 12112 -2455 12168
rect -2405 12112 -2349 12168
rect -2299 12112 -2243 12168
rect -2193 12112 -2137 12168
rect -2511 12029 -2455 12085
rect -2405 12029 -2349 12085
rect -2299 12029 -2243 12085
rect -2193 12029 -2137 12085
rect -2511 11945 -2455 12001
rect -2405 11945 -2349 12001
rect -2299 11945 -2243 12001
rect -2193 11945 -2137 12001
rect -2511 11861 -2455 11917
rect -2405 11861 -2349 11917
rect -2299 11861 -2243 11917
rect -2193 11861 -2137 11917
rect -2511 11777 -2455 11833
rect -2405 11777 -2349 11833
rect -2299 11777 -2243 11833
rect -2193 11777 -2137 11833
rect -2511 11693 -2455 11749
rect -2405 11693 -2349 11749
rect -2299 11693 -2243 11749
rect -2193 11693 -2137 11749
rect -714 12137 -658 12193
rect -626 12137 -570 12193
rect -538 12137 -482 12193
rect -450 12137 -394 12193
rect -362 12137 -306 12193
rect -274 12137 -218 12193
rect -186 12137 -130 12193
rect 8324 12429 8380 12485
rect 8408 12429 8464 12485
rect 8492 12429 8548 12485
rect 8576 12429 8632 12485
rect 8660 12429 8716 12485
rect 8744 12429 8800 12485
rect 8828 12429 8884 12485
rect 10122 12990 10178 13046
rect 10206 12990 10262 13046
rect 10290 12990 10346 13046
rect 10374 12990 10430 13046
rect 10458 12990 10514 13046
rect 10542 12990 10598 13046
rect 10626 12990 10682 13046
rect 10122 12901 10178 12957
rect 10206 12901 10262 12957
rect 10290 12901 10346 12957
rect 10374 12901 10430 12957
rect 10458 12901 10514 12957
rect 10542 12901 10598 12957
rect 10626 12901 10682 12957
rect 10122 12812 10178 12868
rect 10206 12812 10262 12868
rect 10290 12812 10346 12868
rect 10374 12812 10430 12868
rect 10458 12812 10514 12868
rect 10542 12812 10598 12868
rect 10626 12812 10682 12868
rect 10122 12723 10178 12779
rect 10206 12723 10262 12779
rect 10290 12723 10346 12779
rect 10374 12723 10430 12779
rect 10458 12723 10514 12779
rect 10542 12723 10598 12779
rect 10626 12723 10682 12779
rect 10122 12634 10178 12690
rect 10206 12634 10262 12690
rect 10290 12634 10346 12690
rect 10374 12634 10430 12690
rect 10458 12634 10514 12690
rect 10542 12634 10598 12690
rect 10626 12634 10682 12690
rect 10122 12545 10178 12601
rect 10206 12545 10262 12601
rect 10290 12545 10346 12601
rect 10374 12545 10430 12601
rect 10458 12545 10514 12601
rect 10542 12545 10598 12601
rect 10626 12545 10682 12601
rect 10122 12455 10178 12511
rect 10206 12455 10262 12511
rect 10290 12455 10346 12511
rect 10374 12455 10430 12511
rect 10458 12455 10514 12511
rect 10542 12455 10598 12511
rect 10626 12455 10682 12511
rect 11923 12990 11979 13046
rect 12007 12990 12063 13046
rect 12091 12990 12147 13046
rect 12175 12990 12231 13046
rect 12259 12990 12315 13046
rect 12343 12990 12399 13046
rect 12427 12990 12483 13046
rect 11923 12907 11979 12963
rect 12007 12907 12063 12963
rect 12091 12907 12147 12963
rect 12175 12907 12231 12963
rect 12259 12907 12315 12963
rect 12343 12907 12399 12963
rect 12427 12907 12483 12963
rect 11923 12824 11979 12880
rect 12007 12824 12063 12880
rect 12091 12824 12147 12880
rect 12175 12824 12231 12880
rect 12259 12824 12315 12880
rect 12343 12824 12399 12880
rect 12427 12824 12483 12880
rect 11923 12741 11979 12797
rect 12007 12741 12063 12797
rect 12091 12741 12147 12797
rect 12175 12741 12231 12797
rect 12259 12741 12315 12797
rect 12343 12741 12399 12797
rect 12427 12741 12483 12797
rect 11923 12657 11979 12713
rect 12007 12657 12063 12713
rect 12091 12657 12147 12713
rect 12175 12657 12231 12713
rect 12259 12657 12315 12713
rect 12343 12657 12399 12713
rect 12427 12657 12483 12713
rect 11923 12573 11979 12629
rect 12007 12573 12063 12629
rect 12091 12573 12147 12629
rect 12175 12573 12231 12629
rect 12259 12573 12315 12629
rect 12343 12573 12399 12629
rect 12427 12573 12483 12629
rect 11923 12489 11979 12545
rect 12007 12489 12063 12545
rect 12091 12489 12147 12545
rect 12175 12489 12231 12545
rect 12259 12489 12315 12545
rect 12343 12489 12399 12545
rect 12427 12489 12483 12545
rect 8324 12349 8380 12405
rect 8408 12349 8464 12405
rect 8492 12349 8548 12405
rect 8576 12349 8632 12405
rect 8660 12349 8716 12405
rect 8744 12349 8800 12405
rect 8828 12349 8884 12405
rect 8324 12269 8380 12325
rect 8408 12269 8464 12325
rect 8492 12269 8548 12325
rect 8576 12269 8632 12325
rect 8660 12269 8716 12325
rect 8744 12269 8800 12325
rect 8828 12269 8884 12325
rect 8324 12189 8380 12245
rect 8408 12189 8464 12245
rect 8492 12189 8548 12245
rect 8576 12189 8632 12245
rect 8660 12189 8716 12245
rect 8744 12189 8800 12245
rect 8828 12189 8884 12245
rect -714 12057 -658 12113
rect -626 12057 -570 12113
rect -538 12057 -482 12113
rect -450 12057 -394 12113
rect -362 12057 -306 12113
rect -274 12057 -218 12113
rect -186 12057 -130 12113
rect -714 11977 -658 12033
rect -626 11977 -570 12033
rect -538 11977 -482 12033
rect -450 11977 -394 12033
rect -362 11977 -306 12033
rect -274 11977 -218 12033
rect -186 11977 -130 12033
rect -714 11897 -658 11953
rect -626 11897 -570 11953
rect -538 11897 -482 11953
rect -450 11897 -394 11953
rect -362 11897 -306 11953
rect -274 11897 -218 11953
rect -186 11897 -130 11953
rect -714 11817 -658 11873
rect -626 11817 -570 11873
rect -538 11817 -482 11873
rect -450 11817 -394 11873
rect -362 11817 -306 11873
rect -274 11817 -218 11873
rect -186 11817 -130 11873
rect -714 11737 -658 11793
rect -626 11737 -570 11793
rect -538 11737 -482 11793
rect -450 11737 -394 11793
rect -362 11737 -306 11793
rect -274 11737 -218 11793
rect -186 11737 -130 11793
rect -714 11657 -658 11713
rect -626 11657 -570 11713
rect -538 11657 -482 11713
rect -450 11657 -394 11713
rect -362 11657 -306 11713
rect -274 11657 -218 11713
rect -186 11657 -130 11713
rect -714 11577 -658 11633
rect -626 11577 -570 11633
rect -538 11577 -482 11633
rect -450 11577 -394 11633
rect -362 11577 -306 11633
rect -274 11577 -218 11633
rect -186 11577 -130 11633
rect -714 11497 -658 11553
rect -626 11497 -570 11553
rect -538 11497 -482 11553
rect -450 11497 -394 11553
rect -362 11497 -306 11553
rect -274 11497 -218 11553
rect -186 11497 -130 11553
rect -714 11417 -658 11473
rect -626 11417 -570 11473
rect -538 11417 -482 11473
rect -450 11417 -394 11473
rect -362 11417 -306 11473
rect -274 11417 -218 11473
rect -186 11417 -130 11473
rect -714 11337 -658 11393
rect -626 11337 -570 11393
rect -538 11337 -482 11393
rect -450 11337 -394 11393
rect -362 11337 -306 11393
rect -274 11337 -218 11393
rect -186 11337 -130 11393
rect -714 11257 -658 11313
rect -626 11257 -570 11313
rect -538 11257 -482 11313
rect -450 11257 -394 11313
rect -362 11257 -306 11313
rect -274 11257 -218 11313
rect -186 11257 -130 11313
rect -714 11177 -658 11233
rect -626 11177 -570 11233
rect -538 11177 -482 11233
rect -450 11177 -394 11233
rect -362 11177 -306 11233
rect -274 11177 -218 11233
rect -186 11177 -130 11233
rect -714 11097 -658 11153
rect -626 11097 -570 11153
rect -538 11097 -482 11153
rect -450 11097 -394 11153
rect -362 11097 -306 11153
rect -274 11097 -218 11153
rect -186 11097 -130 11153
rect -714 11017 -658 11073
rect -626 11017 -570 11073
rect -538 11017 -482 11073
rect -450 11017 -394 11073
rect -362 11017 -306 11073
rect -274 11017 -218 11073
rect -186 11017 -130 11073
rect -714 10937 -658 10993
rect -626 10937 -570 10993
rect -538 10937 -482 10993
rect -450 10937 -394 10993
rect -362 10937 -306 10993
rect -274 10937 -218 10993
rect -186 10937 -130 10993
rect -714 10857 -658 10913
rect -626 10857 -570 10913
rect -538 10857 -482 10913
rect -450 10857 -394 10913
rect -362 10857 -306 10913
rect -274 10857 -218 10913
rect -186 10857 -130 10913
rect -714 10777 -658 10833
rect -626 10777 -570 10833
rect -538 10777 -482 10833
rect -450 10777 -394 10833
rect -362 10777 -306 10833
rect -274 10777 -218 10833
rect -186 10777 -130 10833
rect -714 10697 -658 10753
rect -626 10697 -570 10753
rect -538 10697 -482 10753
rect -450 10697 -394 10753
rect -362 10697 -306 10753
rect -274 10697 -218 10753
rect -186 10697 -130 10753
rect -714 10617 -658 10673
rect -626 10617 -570 10673
rect -538 10617 -482 10673
rect -450 10617 -394 10673
rect -362 10617 -306 10673
rect -274 10617 -218 10673
rect -186 10617 -130 10673
rect -714 10537 -658 10593
rect -626 10537 -570 10593
rect -538 10537 -482 10593
rect -450 10537 -394 10593
rect -362 10537 -306 10593
rect -274 10537 -218 10593
rect -186 10537 -130 10593
rect -714 10457 -658 10513
rect -626 10457 -570 10513
rect -538 10457 -482 10513
rect -450 10457 -394 10513
rect -362 10457 -306 10513
rect -274 10457 -218 10513
rect -186 10457 -130 10513
rect -714 10377 -658 10433
rect -626 10377 -570 10433
rect -538 10377 -482 10433
rect -450 10377 -394 10433
rect -362 10377 -306 10433
rect -274 10377 -218 10433
rect -186 10377 -130 10433
rect -714 10297 -658 10353
rect -626 10297 -570 10353
rect -538 10297 -482 10353
rect -450 10297 -394 10353
rect -362 10297 -306 10353
rect -274 10297 -218 10353
rect -186 10297 -130 10353
rect -714 10217 -658 10273
rect -626 10217 -570 10273
rect -538 10217 -482 10273
rect -450 10217 -394 10273
rect -362 10217 -306 10273
rect -274 10217 -218 10273
rect -186 10217 -130 10273
rect -714 10137 -658 10193
rect -626 10137 -570 10193
rect -538 10137 -482 10193
rect -450 10137 -394 10193
rect -362 10137 -306 10193
rect -274 10137 -218 10193
rect -186 10137 -130 10193
rect -714 10057 -658 10113
rect -626 10057 -570 10113
rect -538 10057 -482 10113
rect -450 10057 -394 10113
rect -362 10057 -306 10113
rect -274 10057 -218 10113
rect -186 10057 -130 10113
rect -714 9977 -658 10033
rect -626 9977 -570 10033
rect -538 9977 -482 10033
rect -450 9977 -394 10033
rect -362 9977 -306 10033
rect -274 9977 -218 10033
rect -186 9977 -130 10033
rect -714 9897 -658 9953
rect -626 9897 -570 9953
rect -538 9897 -482 9953
rect -450 9897 -394 9953
rect -362 9897 -306 9953
rect -274 9897 -218 9953
rect -186 9897 -130 9953
rect -714 9817 -658 9873
rect -626 9817 -570 9873
rect -538 9817 -482 9873
rect -450 9817 -394 9873
rect -362 9817 -306 9873
rect -274 9817 -218 9873
rect -186 9817 -130 9873
rect -714 9737 -658 9793
rect -626 9737 -570 9793
rect -538 9737 -482 9793
rect -450 9737 -394 9793
rect -362 9737 -306 9793
rect -274 9737 -218 9793
rect -186 9737 -130 9793
rect -714 9657 -658 9713
rect -626 9657 -570 9713
rect -538 9657 -482 9713
rect -450 9657 -394 9713
rect -362 9657 -306 9713
rect -274 9657 -218 9713
rect -186 9657 -130 9713
rect -714 9577 -658 9633
rect -626 9577 -570 9633
rect -538 9577 -482 9633
rect -450 9577 -394 9633
rect -362 9577 -306 9633
rect -274 9577 -218 9633
rect -186 9577 -130 9633
rect -714 9497 -658 9553
rect -626 9497 -570 9553
rect -538 9497 -482 9553
rect -450 9497 -394 9553
rect -362 9497 -306 9553
rect -274 9497 -218 9553
rect -186 9497 -130 9553
rect -714 9417 -658 9473
rect -626 9417 -570 9473
rect -538 9417 -482 9473
rect -450 9417 -394 9473
rect -362 9417 -306 9473
rect -274 9417 -218 9473
rect -186 9417 -130 9473
rect -714 9337 -658 9393
rect -626 9337 -570 9393
rect -538 9337 -482 9393
rect -450 9337 -394 9393
rect -362 9337 -306 9393
rect -274 9337 -218 9393
rect -186 9337 -130 9393
rect -714 9257 -658 9313
rect -626 9257 -570 9313
rect -538 9257 -482 9313
rect -450 9257 -394 9313
rect -362 9257 -306 9313
rect -274 9257 -218 9313
rect -186 9257 -130 9313
rect -714 9177 -658 9233
rect -626 9177 -570 9233
rect -538 9177 -482 9233
rect -450 9177 -394 9233
rect -362 9177 -306 9233
rect -274 9177 -218 9233
rect -186 9177 -130 9233
rect -714 9097 -658 9153
rect -626 9097 -570 9153
rect -538 9097 -482 9153
rect -450 9097 -394 9153
rect -362 9097 -306 9153
rect -274 9097 -218 9153
rect -186 9097 -130 9153
rect -714 9017 -658 9073
rect -626 9017 -570 9073
rect -538 9017 -482 9073
rect -450 9017 -394 9073
rect -362 9017 -306 9073
rect -274 9017 -218 9073
rect -186 9017 -130 9073
rect -714 8937 -658 8993
rect -626 8937 -570 8993
rect -538 8937 -482 8993
rect -450 8937 -394 8993
rect -362 8937 -306 8993
rect -274 8937 -218 8993
rect -186 8937 -130 8993
rect -714 8857 -658 8913
rect -626 8857 -570 8913
rect -538 8857 -482 8913
rect -450 8857 -394 8913
rect -362 8857 -306 8913
rect -274 8857 -218 8913
rect -186 8857 -130 8913
rect -714 8777 -658 8833
rect -626 8777 -570 8833
rect -538 8777 -482 8833
rect -450 8777 -394 8833
rect -362 8777 -306 8833
rect -274 8777 -218 8833
rect -186 8777 -130 8833
rect -714 8697 -658 8753
rect -626 8697 -570 8753
rect -538 8697 -482 8753
rect -450 8697 -394 8753
rect -362 8697 -306 8753
rect -274 8697 -218 8753
rect -186 8697 -130 8753
rect -714 8617 -658 8673
rect -626 8617 -570 8673
rect -538 8617 -482 8673
rect -450 8617 -394 8673
rect -362 8617 -306 8673
rect -274 8617 -218 8673
rect -186 8617 -130 8673
rect -714 8537 -658 8593
rect -626 8537 -570 8593
rect -538 8537 -482 8593
rect -450 8537 -394 8593
rect -362 8537 -306 8593
rect -274 8537 -218 8593
rect -186 8537 -130 8593
rect -714 8457 -658 8513
rect -626 8457 -570 8513
rect -538 8457 -482 8513
rect -450 8457 -394 8513
rect -362 8457 -306 8513
rect -274 8457 -218 8513
rect -186 8457 -130 8513
rect -714 8377 -658 8433
rect -626 8377 -570 8433
rect -538 8377 -482 8433
rect -450 8377 -394 8433
rect -362 8377 -306 8433
rect -274 8377 -218 8433
rect -186 8377 -130 8433
rect -714 8297 -658 8353
rect -626 8297 -570 8353
rect -538 8297 -482 8353
rect -450 8297 -394 8353
rect -362 8297 -306 8353
rect -274 8297 -218 8353
rect -186 8297 -130 8353
rect -714 8217 -658 8273
rect -626 8217 -570 8273
rect -538 8217 -482 8273
rect -450 8217 -394 8273
rect -362 8217 -306 8273
rect -274 8217 -218 8273
rect -186 8217 -130 8273
rect -714 8137 -658 8193
rect -626 8137 -570 8193
rect -538 8137 -482 8193
rect -450 8137 -394 8193
rect -362 8137 -306 8193
rect -274 8137 -218 8193
rect -186 8137 -130 8193
rect -714 8057 -658 8113
rect -626 8057 -570 8113
rect -538 8057 -482 8113
rect -450 8057 -394 8113
rect -362 8057 -306 8113
rect -274 8057 -218 8113
rect -186 8057 -130 8113
rect -714 7977 -658 8033
rect -626 7977 -570 8033
rect -538 7977 -482 8033
rect -450 7977 -394 8033
rect -362 7977 -306 8033
rect -274 7977 -218 8033
rect -186 7977 -130 8033
rect -714 7897 -658 7953
rect -626 7897 -570 7953
rect -538 7897 -482 7953
rect -450 7897 -394 7953
rect -362 7897 -306 7953
rect -274 7897 -218 7953
rect -186 7897 -130 7953
rect -714 7817 -658 7873
rect -626 7817 -570 7873
rect -538 7817 -482 7873
rect -450 7817 -394 7873
rect -362 7817 -306 7873
rect -274 7817 -218 7873
rect -186 7817 -130 7873
rect -714 7737 -658 7793
rect -626 7737 -570 7793
rect -538 7737 -482 7793
rect -450 7737 -394 7793
rect -362 7737 -306 7793
rect -274 7737 -218 7793
rect -186 7737 -130 7793
rect -714 7657 -658 7713
rect -626 7657 -570 7713
rect -538 7657 -482 7713
rect -450 7657 -394 7713
rect -362 7657 -306 7713
rect -274 7657 -218 7713
rect -186 7657 -130 7713
rect -714 7577 -658 7633
rect -626 7577 -570 7633
rect -538 7577 -482 7633
rect -450 7577 -394 7633
rect -362 7577 -306 7633
rect -274 7577 -218 7633
rect -186 7577 -130 7633
rect -714 7497 -658 7553
rect -626 7497 -570 7553
rect -538 7497 -482 7553
rect -450 7497 -394 7553
rect -362 7497 -306 7553
rect -274 7497 -218 7553
rect -186 7497 -130 7553
rect -714 7417 -658 7473
rect -626 7417 -570 7473
rect -538 7417 -482 7473
rect -450 7417 -394 7473
rect -362 7417 -306 7473
rect -274 7417 -218 7473
rect -186 7417 -130 7473
rect -714 7337 -658 7393
rect -626 7337 -570 7393
rect -538 7337 -482 7393
rect -450 7337 -394 7393
rect -362 7337 -306 7393
rect -274 7337 -218 7393
rect -186 7337 -130 7393
rect -714 7257 -658 7313
rect -626 7257 -570 7313
rect -538 7257 -482 7313
rect -450 7257 -394 7313
rect -362 7257 -306 7313
rect -274 7257 -218 7313
rect -186 7257 -130 7313
rect -714 7177 -658 7233
rect -626 7177 -570 7233
rect -538 7177 -482 7233
rect -450 7177 -394 7233
rect -362 7177 -306 7233
rect -274 7177 -218 7233
rect -186 7177 -130 7233
rect -714 7097 -658 7153
rect -626 7097 -570 7153
rect -538 7097 -482 7153
rect -450 7097 -394 7153
rect -362 7097 -306 7153
rect -274 7097 -218 7153
rect -186 7097 -130 7153
rect -714 7017 -658 7073
rect -626 7017 -570 7073
rect -538 7017 -482 7073
rect -450 7017 -394 7073
rect -362 7017 -306 7073
rect -274 7017 -218 7073
rect -186 7017 -130 7073
rect -714 6937 -658 6993
rect -626 6937 -570 6993
rect -538 6937 -482 6993
rect -450 6937 -394 6993
rect -362 6937 -306 6993
rect -274 6937 -218 6993
rect -186 6937 -130 6993
rect -714 6856 -658 6912
rect -626 6856 -570 6912
rect -538 6856 -482 6912
rect -450 6856 -394 6912
rect -362 6856 -306 6912
rect -274 6856 -218 6912
rect -186 6856 -130 6912
rect -714 6775 -658 6831
rect -626 6775 -570 6831
rect -538 6775 -482 6831
rect -450 6775 -394 6831
rect -362 6775 -306 6831
rect -274 6775 -218 6831
rect -186 6775 -130 6831
rect -714 6694 -658 6750
rect -626 6694 -570 6750
rect -538 6694 -482 6750
rect -450 6694 -394 6750
rect -362 6694 -306 6750
rect -274 6694 -218 6750
rect -186 6694 -130 6750
rect -714 6613 -658 6669
rect -626 6613 -570 6669
rect -538 6613 -482 6669
rect -450 6613 -394 6669
rect -362 6613 -306 6669
rect -274 6613 -218 6669
rect -186 6613 -130 6669
rect -714 6532 -658 6588
rect -626 6532 -570 6588
rect -538 6532 -482 6588
rect -450 6532 -394 6588
rect -362 6532 -306 6588
rect -274 6532 -218 6588
rect -186 6532 -130 6588
rect -714 6451 -658 6507
rect -626 6451 -570 6507
rect -538 6451 -482 6507
rect -450 6451 -394 6507
rect -362 6451 -306 6507
rect -274 6451 -218 6507
rect -186 6451 -130 6507
rect -714 6370 -658 6426
rect -626 6370 -570 6426
rect -538 6370 -482 6426
rect -450 6370 -394 6426
rect -362 6370 -306 6426
rect -274 6370 -218 6426
rect -186 6370 -130 6426
rect -714 6289 -658 6345
rect -626 6289 -570 6345
rect -538 6289 -482 6345
rect -450 6289 -394 6345
rect -362 6289 -306 6345
rect -274 6289 -218 6345
rect -186 6289 -130 6345
rect -714 6208 -658 6264
rect -626 6208 -570 6264
rect -538 6208 -482 6264
rect -450 6208 -394 6264
rect -362 6208 -306 6264
rect -274 6208 -218 6264
rect -186 6208 -130 6264
rect -714 6127 -658 6183
rect -626 6127 -570 6183
rect -538 6127 -482 6183
rect -450 6127 -394 6183
rect -362 6127 -306 6183
rect -274 6127 -218 6183
rect -186 6127 -130 6183
rect -714 6046 -658 6102
rect -626 6046 -570 6102
rect -538 6046 -482 6102
rect -450 6046 -394 6102
rect -362 6046 -306 6102
rect -274 6046 -218 6102
rect -186 6046 -130 6102
rect -714 5965 -658 6021
rect -626 5965 -570 6021
rect -538 5965 -482 6021
rect -450 5965 -394 6021
rect -362 5965 -306 6021
rect -274 5965 -218 6021
rect -186 5965 -130 6021
rect -714 5884 -658 5940
rect -626 5884 -570 5940
rect -538 5884 -482 5940
rect -450 5884 -394 5940
rect -362 5884 -306 5940
rect -274 5884 -218 5940
rect -186 5884 -130 5940
rect -714 5803 -658 5859
rect -626 5803 -570 5859
rect -538 5803 -482 5859
rect -450 5803 -394 5859
rect -362 5803 -306 5859
rect -274 5803 -218 5859
rect -186 5803 -130 5859
rect -714 5722 -658 5778
rect -626 5722 -570 5778
rect -538 5722 -482 5778
rect -450 5722 -394 5778
rect -362 5722 -306 5778
rect -274 5722 -218 5778
rect -186 5722 -130 5778
rect -714 5641 -658 5697
rect -626 5641 -570 5697
rect -538 5641 -482 5697
rect -450 5641 -394 5697
rect -362 5641 -306 5697
rect -274 5641 -218 5697
rect -186 5641 -130 5697
rect -714 5560 -658 5616
rect -626 5560 -570 5616
rect -538 5560 -482 5616
rect -450 5560 -394 5616
rect -362 5560 -306 5616
rect -274 5560 -218 5616
rect -186 5560 -130 5616
rect -714 5479 -658 5535
rect -626 5479 -570 5535
rect -538 5479 -482 5535
rect -450 5479 -394 5535
rect -362 5479 -306 5535
rect -274 5479 -218 5535
rect -186 5479 -130 5535
rect -714 5398 -658 5454
rect -626 5398 -570 5454
rect -538 5398 -482 5454
rect -450 5398 -394 5454
rect -362 5398 -306 5454
rect -274 5398 -218 5454
rect -186 5398 -130 5454
rect -714 5317 -658 5373
rect -626 5317 -570 5373
rect -538 5317 -482 5373
rect -450 5317 -394 5373
rect -362 5317 -306 5373
rect -274 5317 -218 5373
rect -186 5317 -130 5373
rect -714 5236 -658 5292
rect -626 5236 -570 5292
rect -538 5236 -482 5292
rect -450 5236 -394 5292
rect -362 5236 -306 5292
rect -274 5236 -218 5292
rect -186 5236 -130 5292
rect -714 5155 -658 5211
rect -626 5155 -570 5211
rect -538 5155 -482 5211
rect -450 5155 -394 5211
rect -362 5155 -306 5211
rect -274 5155 -218 5211
rect -186 5155 -130 5211
rect 8324 12109 8380 12165
rect 8408 12109 8464 12165
rect 8492 12109 8548 12165
rect 8576 12109 8632 12165
rect 8660 12109 8716 12165
rect 8744 12109 8800 12165
rect 8828 12109 8884 12165
rect 8324 12029 8380 12085
rect 8408 12029 8464 12085
rect 8492 12029 8548 12085
rect 8576 12029 8632 12085
rect 8660 12029 8716 12085
rect 8744 12029 8800 12085
rect 8828 12029 8884 12085
rect 8324 11949 8380 12005
rect 8408 11949 8464 12005
rect 8492 11949 8548 12005
rect 8576 11949 8632 12005
rect 8660 11949 8716 12005
rect 8744 11949 8800 12005
rect 8828 11949 8884 12005
rect 8324 11869 8380 11925
rect 8408 11869 8464 11925
rect 8492 11869 8548 11925
rect 8576 11869 8632 11925
rect 8660 11869 8716 11925
rect 8744 11869 8800 11925
rect 8828 11869 8884 11925
rect 8324 11789 8380 11845
rect 8408 11789 8464 11845
rect 8492 11789 8548 11845
rect 8576 11789 8632 11845
rect 8660 11789 8716 11845
rect 8744 11789 8800 11845
rect 8828 11789 8884 11845
rect 8324 11709 8380 11765
rect 8408 11709 8464 11765
rect 8492 11709 8548 11765
rect 8576 11709 8632 11765
rect 8660 11709 8716 11765
rect 8744 11709 8800 11765
rect 8828 11709 8884 11765
rect 8324 11629 8380 11685
rect 8408 11629 8464 11685
rect 8492 11629 8548 11685
rect 8576 11629 8632 11685
rect 8660 11629 8716 11685
rect 8744 11629 8800 11685
rect 8828 11629 8884 11685
rect 8324 11549 8380 11605
rect 8408 11549 8464 11605
rect 8492 11549 8548 11605
rect 8576 11549 8632 11605
rect 8660 11549 8716 11605
rect 8744 11549 8800 11605
rect 8828 11549 8884 11605
rect 8324 11469 8380 11525
rect 8408 11469 8464 11525
rect 8492 11469 8548 11525
rect 8576 11469 8632 11525
rect 8660 11469 8716 11525
rect 8744 11469 8800 11525
rect 8828 11469 8884 11525
rect 8324 11389 8380 11445
rect 8408 11389 8464 11445
rect 8492 11389 8548 11445
rect 8576 11389 8632 11445
rect 8660 11389 8716 11445
rect 8744 11389 8800 11445
rect 8828 11389 8884 11445
rect 8324 11309 8380 11365
rect 8408 11309 8464 11365
rect 8492 11309 8548 11365
rect 8576 11309 8632 11365
rect 8660 11309 8716 11365
rect 8744 11309 8800 11365
rect 8828 11309 8884 11365
rect 8324 11229 8380 11285
rect 8408 11229 8464 11285
rect 8492 11229 8548 11285
rect 8576 11229 8632 11285
rect 8660 11229 8716 11285
rect 8744 11229 8800 11285
rect 8828 11229 8884 11285
rect 8324 11149 8380 11205
rect 8408 11149 8464 11205
rect 8492 11149 8548 11205
rect 8576 11149 8632 11205
rect 8660 11149 8716 11205
rect 8744 11149 8800 11205
rect 8828 11149 8884 11205
rect 8324 11069 8380 11125
rect 8408 11069 8464 11125
rect 8492 11069 8548 11125
rect 8576 11069 8632 11125
rect 8660 11069 8716 11125
rect 8744 11069 8800 11125
rect 8828 11069 8884 11125
rect 8324 10989 8380 11045
rect 8408 10989 8464 11045
rect 8492 10989 8548 11045
rect 8576 10989 8632 11045
rect 8660 10989 8716 11045
rect 8744 10989 8800 11045
rect 8828 10989 8884 11045
rect 8324 10909 8380 10965
rect 8408 10909 8464 10965
rect 8492 10909 8548 10965
rect 8576 10909 8632 10965
rect 8660 10909 8716 10965
rect 8744 10909 8800 10965
rect 8828 10909 8884 10965
rect 8324 10829 8380 10885
rect 8408 10829 8464 10885
rect 8492 10829 8548 10885
rect 8576 10829 8632 10885
rect 8660 10829 8716 10885
rect 8744 10829 8800 10885
rect 8828 10829 8884 10885
rect 8324 10749 8380 10805
rect 8408 10749 8464 10805
rect 8492 10749 8548 10805
rect 8576 10749 8632 10805
rect 8660 10749 8716 10805
rect 8744 10749 8800 10805
rect 8828 10749 8884 10805
rect 8324 10669 8380 10725
rect 8408 10669 8464 10725
rect 8492 10669 8548 10725
rect 8576 10669 8632 10725
rect 8660 10669 8716 10725
rect 8744 10669 8800 10725
rect 8828 10669 8884 10725
rect 8324 10589 8380 10645
rect 8408 10589 8464 10645
rect 8492 10589 8548 10645
rect 8576 10589 8632 10645
rect 8660 10589 8716 10645
rect 8744 10589 8800 10645
rect 8828 10589 8884 10645
rect 8324 10509 8380 10565
rect 8408 10509 8464 10565
rect 8492 10509 8548 10565
rect 8576 10509 8632 10565
rect 8660 10509 8716 10565
rect 8744 10509 8800 10565
rect 8828 10509 8884 10565
rect 8324 10429 8380 10485
rect 8408 10429 8464 10485
rect 8492 10429 8548 10485
rect 8576 10429 8632 10485
rect 8660 10429 8716 10485
rect 8744 10429 8800 10485
rect 8828 10429 8884 10485
rect 8324 10349 8380 10405
rect 8408 10349 8464 10405
rect 8492 10349 8548 10405
rect 8576 10349 8632 10405
rect 8660 10349 8716 10405
rect 8744 10349 8800 10405
rect 8828 10349 8884 10405
rect 8324 10269 8380 10325
rect 8408 10269 8464 10325
rect 8492 10269 8548 10325
rect 8576 10269 8632 10325
rect 8660 10269 8716 10325
rect 8744 10269 8800 10325
rect 8828 10269 8884 10325
rect 8324 10189 8380 10245
rect 8408 10189 8464 10245
rect 8492 10189 8548 10245
rect 8576 10189 8632 10245
rect 8660 10189 8716 10245
rect 8744 10189 8800 10245
rect 8828 10189 8884 10245
rect 8324 10109 8380 10165
rect 8408 10109 8464 10165
rect 8492 10109 8548 10165
rect 8576 10109 8632 10165
rect 8660 10109 8716 10165
rect 8744 10109 8800 10165
rect 8828 10109 8884 10165
rect 8324 10029 8380 10085
rect 8408 10029 8464 10085
rect 8492 10029 8548 10085
rect 8576 10029 8632 10085
rect 8660 10029 8716 10085
rect 8744 10029 8800 10085
rect 8828 10029 8884 10085
rect 8324 9949 8380 10005
rect 8408 9949 8464 10005
rect 8492 9949 8548 10005
rect 8576 9949 8632 10005
rect 8660 9949 8716 10005
rect 8744 9949 8800 10005
rect 8828 9949 8884 10005
rect 8324 9869 8380 9925
rect 8408 9869 8464 9925
rect 8492 9869 8548 9925
rect 8576 9869 8632 9925
rect 8660 9869 8716 9925
rect 8744 9869 8800 9925
rect 8828 9869 8884 9925
rect 8324 9789 8380 9845
rect 8408 9789 8464 9845
rect 8492 9789 8548 9845
rect 8576 9789 8632 9845
rect 8660 9789 8716 9845
rect 8744 9789 8800 9845
rect 8828 9789 8884 9845
rect 8324 9709 8380 9765
rect 8408 9709 8464 9765
rect 8492 9709 8548 9765
rect 8576 9709 8632 9765
rect 8660 9709 8716 9765
rect 8744 9709 8800 9765
rect 8828 9709 8884 9765
rect 8324 9629 8380 9685
rect 8408 9629 8464 9685
rect 8492 9629 8548 9685
rect 8576 9629 8632 9685
rect 8660 9629 8716 9685
rect 8744 9629 8800 9685
rect 8828 9629 8884 9685
rect 8324 9549 8380 9605
rect 8408 9549 8464 9605
rect 8492 9549 8548 9605
rect 8576 9549 8632 9605
rect 8660 9549 8716 9605
rect 8744 9549 8800 9605
rect 8828 9549 8884 9605
rect 8324 9468 8380 9524
rect 8408 9468 8464 9524
rect 8492 9468 8548 9524
rect 8576 9468 8632 9524
rect 8660 9468 8716 9524
rect 8744 9468 8800 9524
rect 8828 9468 8884 9524
rect 8324 9387 8380 9443
rect 8408 9387 8464 9443
rect 8492 9387 8548 9443
rect 8576 9387 8632 9443
rect 8660 9387 8716 9443
rect 8744 9387 8800 9443
rect 8828 9387 8884 9443
rect 8324 9306 8380 9362
rect 8408 9306 8464 9362
rect 8492 9306 8548 9362
rect 8576 9306 8632 9362
rect 8660 9306 8716 9362
rect 8744 9306 8800 9362
rect 8828 9306 8884 9362
rect 8324 9225 8380 9281
rect 8408 9225 8464 9281
rect 8492 9225 8548 9281
rect 8576 9225 8632 9281
rect 8660 9225 8716 9281
rect 8744 9225 8800 9281
rect 8828 9225 8884 9281
rect 8324 9144 8380 9200
rect 8408 9144 8464 9200
rect 8492 9144 8548 9200
rect 8576 9144 8632 9200
rect 8660 9144 8716 9200
rect 8744 9144 8800 9200
rect 8828 9144 8884 9200
rect 8324 9063 8380 9119
rect 8408 9063 8464 9119
rect 8492 9063 8548 9119
rect 8576 9063 8632 9119
rect 8660 9063 8716 9119
rect 8744 9063 8800 9119
rect 8828 9063 8884 9119
rect 8324 8982 8380 9038
rect 8408 8982 8464 9038
rect 8492 8982 8548 9038
rect 8576 8982 8632 9038
rect 8660 8982 8716 9038
rect 8744 8982 8800 9038
rect 8828 8982 8884 9038
rect 8324 8901 8380 8957
rect 8408 8901 8464 8957
rect 8492 8901 8548 8957
rect 8576 8901 8632 8957
rect 8660 8901 8716 8957
rect 8744 8901 8800 8957
rect 8828 8901 8884 8957
rect 8324 8820 8380 8876
rect 8408 8820 8464 8876
rect 8492 8820 8548 8876
rect 8576 8820 8632 8876
rect 8660 8820 8716 8876
rect 8744 8820 8800 8876
rect 8828 8820 8884 8876
rect 8324 8739 8380 8795
rect 8408 8739 8464 8795
rect 8492 8739 8548 8795
rect 8576 8739 8632 8795
rect 8660 8739 8716 8795
rect 8744 8739 8800 8795
rect 8828 8739 8884 8795
rect 8324 8658 8380 8714
rect 8408 8658 8464 8714
rect 8492 8658 8548 8714
rect 8576 8658 8632 8714
rect 8660 8658 8716 8714
rect 8744 8658 8800 8714
rect 8828 8658 8884 8714
rect 8324 8577 8380 8633
rect 8408 8577 8464 8633
rect 8492 8577 8548 8633
rect 8576 8577 8632 8633
rect 8660 8577 8716 8633
rect 8744 8577 8800 8633
rect 8828 8577 8884 8633
rect 8324 8496 8380 8552
rect 8408 8496 8464 8552
rect 8492 8496 8548 8552
rect 8576 8496 8632 8552
rect 8660 8496 8716 8552
rect 8744 8496 8800 8552
rect 8828 8496 8884 8552
rect 8324 8415 8380 8471
rect 8408 8415 8464 8471
rect 8492 8415 8548 8471
rect 8576 8415 8632 8471
rect 8660 8415 8716 8471
rect 8744 8415 8800 8471
rect 8828 8415 8884 8471
rect 8324 8334 8380 8390
rect 8408 8334 8464 8390
rect 8492 8334 8548 8390
rect 8576 8334 8632 8390
rect 8660 8334 8716 8390
rect 8744 8334 8800 8390
rect 8828 8334 8884 8390
rect 8324 8253 8380 8309
rect 8408 8253 8464 8309
rect 8492 8253 8548 8309
rect 8576 8253 8632 8309
rect 8660 8253 8716 8309
rect 8744 8253 8800 8309
rect 8828 8253 8884 8309
rect 8324 8172 8380 8228
rect 8408 8172 8464 8228
rect 8492 8172 8548 8228
rect 8576 8172 8632 8228
rect 8660 8172 8716 8228
rect 8744 8172 8800 8228
rect 8828 8172 8884 8228
rect 8324 8091 8380 8147
rect 8408 8091 8464 8147
rect 8492 8091 8548 8147
rect 8576 8091 8632 8147
rect 8660 8091 8716 8147
rect 8744 8091 8800 8147
rect 8828 8091 8884 8147
rect 8324 8010 8380 8066
rect 8408 8010 8464 8066
rect 8492 8010 8548 8066
rect 8576 8010 8632 8066
rect 8660 8010 8716 8066
rect 8744 8010 8800 8066
rect 8828 8010 8884 8066
rect 8324 7929 8380 7985
rect 8408 7929 8464 7985
rect 8492 7929 8548 7985
rect 8576 7929 8632 7985
rect 8660 7929 8716 7985
rect 8744 7929 8800 7985
rect 8828 7929 8884 7985
rect 8324 7848 8380 7904
rect 8408 7848 8464 7904
rect 8492 7848 8548 7904
rect 8576 7848 8632 7904
rect 8660 7848 8716 7904
rect 8744 7848 8800 7904
rect 8828 7848 8884 7904
rect 8324 7767 8380 7823
rect 8408 7767 8464 7823
rect 8492 7767 8548 7823
rect 8576 7767 8632 7823
rect 8660 7767 8716 7823
rect 8744 7767 8800 7823
rect 8828 7767 8884 7823
rect 8324 7686 8380 7742
rect 8408 7686 8464 7742
rect 8492 7686 8548 7742
rect 8576 7686 8632 7742
rect 8660 7686 8716 7742
rect 8744 7686 8800 7742
rect 8828 7686 8884 7742
rect 8324 7605 8380 7661
rect 8408 7605 8464 7661
rect 8492 7605 8548 7661
rect 8576 7605 8632 7661
rect 8660 7605 8716 7661
rect 8744 7605 8800 7661
rect 8828 7605 8884 7661
rect 8324 7524 8380 7580
rect 8408 7524 8464 7580
rect 8492 7524 8548 7580
rect 8576 7524 8632 7580
rect 8660 7524 8716 7580
rect 8744 7524 8800 7580
rect 8828 7524 8884 7580
rect 8324 7443 8380 7499
rect 8408 7443 8464 7499
rect 8492 7443 8548 7499
rect 8576 7443 8632 7499
rect 8660 7443 8716 7499
rect 8744 7443 8800 7499
rect 8828 7443 8884 7499
rect 8324 7362 8380 7418
rect 8408 7362 8464 7418
rect 8492 7362 8548 7418
rect 8576 7362 8632 7418
rect 8660 7362 8716 7418
rect 8744 7362 8800 7418
rect 8828 7362 8884 7418
rect 8324 7281 8380 7337
rect 8408 7281 8464 7337
rect 8492 7281 8548 7337
rect 8576 7281 8632 7337
rect 8660 7281 8716 7337
rect 8744 7281 8800 7337
rect 8828 7281 8884 7337
rect 8324 7200 8380 7256
rect 8408 7200 8464 7256
rect 8492 7200 8548 7256
rect 8576 7200 8632 7256
rect 8660 7200 8716 7256
rect 8744 7200 8800 7256
rect 8828 7200 8884 7256
rect 8324 7119 8380 7175
rect 8408 7119 8464 7175
rect 8492 7119 8548 7175
rect 8576 7119 8632 7175
rect 8660 7119 8716 7175
rect 8744 7119 8800 7175
rect 8828 7119 8884 7175
rect 8324 7038 8380 7094
rect 8408 7038 8464 7094
rect 8492 7038 8548 7094
rect 8576 7038 8632 7094
rect 8660 7038 8716 7094
rect 8744 7038 8800 7094
rect 8828 7038 8884 7094
rect 8324 6957 8380 7013
rect 8408 6957 8464 7013
rect 8492 6957 8548 7013
rect 8576 6957 8632 7013
rect 8660 6957 8716 7013
rect 8744 6957 8800 7013
rect 8828 6957 8884 7013
rect 8324 6876 8380 6932
rect 8408 6876 8464 6932
rect 8492 6876 8548 6932
rect 8576 6876 8632 6932
rect 8660 6876 8716 6932
rect 8744 6876 8800 6932
rect 8828 6876 8884 6932
rect 8324 6795 8380 6851
rect 8408 6795 8464 6851
rect 8492 6795 8548 6851
rect 8576 6795 8632 6851
rect 8660 6795 8716 6851
rect 8744 6795 8800 6851
rect 8828 6795 8884 6851
rect 8324 6714 8380 6770
rect 8408 6714 8464 6770
rect 8492 6714 8548 6770
rect 8576 6714 8632 6770
rect 8660 6714 8716 6770
rect 8744 6714 8800 6770
rect 8828 6714 8884 6770
rect 8324 6633 8380 6689
rect 8408 6633 8464 6689
rect 8492 6633 8548 6689
rect 8576 6633 8632 6689
rect 8660 6633 8716 6689
rect 8744 6633 8800 6689
rect 8828 6633 8884 6689
rect 8324 6552 8380 6608
rect 8408 6552 8464 6608
rect 8492 6552 8548 6608
rect 8576 6552 8632 6608
rect 8660 6552 8716 6608
rect 8744 6552 8800 6608
rect 8828 6552 8884 6608
rect 8324 6471 8380 6527
rect 8408 6471 8464 6527
rect 8492 6471 8548 6527
rect 8576 6471 8632 6527
rect 8660 6471 8716 6527
rect 8744 6471 8800 6527
rect 8828 6471 8884 6527
rect 8324 6390 8380 6446
rect 8408 6390 8464 6446
rect 8492 6390 8548 6446
rect 8576 6390 8632 6446
rect 8660 6390 8716 6446
rect 8744 6390 8800 6446
rect 8828 6390 8884 6446
rect 8324 6309 8380 6365
rect 8408 6309 8464 6365
rect 8492 6309 8548 6365
rect 8576 6309 8632 6365
rect 8660 6309 8716 6365
rect 8744 6309 8800 6365
rect 8828 6309 8884 6365
rect 8324 6228 8380 6284
rect 8408 6228 8464 6284
rect 8492 6228 8548 6284
rect 8576 6228 8632 6284
rect 8660 6228 8716 6284
rect 8744 6228 8800 6284
rect 8828 6228 8884 6284
rect 8324 6147 8380 6203
rect 8408 6147 8464 6203
rect 8492 6147 8548 6203
rect 8576 6147 8632 6203
rect 8660 6147 8716 6203
rect 8744 6147 8800 6203
rect 8828 6147 8884 6203
rect 8324 6066 8380 6122
rect 8408 6066 8464 6122
rect 8492 6066 8548 6122
rect 8576 6066 8632 6122
rect 8660 6066 8716 6122
rect 8744 6066 8800 6122
rect 8828 6066 8884 6122
rect 8324 5985 8380 6041
rect 8408 5985 8464 6041
rect 8492 5985 8548 6041
rect 8576 5985 8632 6041
rect 8660 5985 8716 6041
rect 8744 5985 8800 6041
rect 8828 5985 8884 6041
rect 8324 5904 8380 5960
rect 8408 5904 8464 5960
rect 8492 5904 8548 5960
rect 8576 5904 8632 5960
rect 8660 5904 8716 5960
rect 8744 5904 8800 5960
rect 8828 5904 8884 5960
rect 8324 5823 8380 5879
rect 8408 5823 8464 5879
rect 8492 5823 8548 5879
rect 8576 5823 8632 5879
rect 8660 5823 8716 5879
rect 8744 5823 8800 5879
rect 8828 5823 8884 5879
rect 8324 5742 8380 5798
rect 8408 5742 8464 5798
rect 8492 5742 8548 5798
rect 8576 5742 8632 5798
rect 8660 5742 8716 5798
rect 8744 5742 8800 5798
rect 8828 5742 8884 5798
rect 8324 5661 8380 5717
rect 8408 5661 8464 5717
rect 8492 5661 8548 5717
rect 8576 5661 8632 5717
rect 8660 5661 8716 5717
rect 8744 5661 8800 5717
rect 8828 5661 8884 5717
rect 8324 5580 8380 5636
rect 8408 5580 8464 5636
rect 8492 5580 8548 5636
rect 8576 5580 8632 5636
rect 8660 5580 8716 5636
rect 8744 5580 8800 5636
rect 8828 5580 8884 5636
rect 8324 5499 8380 5555
rect 8408 5499 8464 5555
rect 8492 5499 8548 5555
rect 8576 5499 8632 5555
rect 8660 5499 8716 5555
rect 8744 5499 8800 5555
rect 8828 5499 8884 5555
rect 8324 5418 8380 5474
rect 8408 5418 8464 5474
rect 8492 5418 8548 5474
rect 8576 5418 8632 5474
rect 8660 5418 8716 5474
rect 8744 5418 8800 5474
rect 8828 5418 8884 5474
rect 8324 5337 8380 5393
rect 8408 5337 8464 5393
rect 8492 5337 8548 5393
rect 8576 5337 8632 5393
rect 8660 5337 8716 5393
rect 8744 5337 8800 5393
rect 8828 5337 8884 5393
rect 8324 5256 8380 5312
rect 8408 5256 8464 5312
rect 8492 5256 8548 5312
rect 8576 5256 8632 5312
rect 8660 5256 8716 5312
rect 8744 5256 8800 5312
rect 8828 5256 8884 5312
rect -714 5074 -658 5130
rect -626 5074 -570 5130
rect -538 5074 -482 5130
rect -450 5074 -394 5130
rect -362 5074 -306 5130
rect -274 5074 -218 5130
rect -186 5074 -130 5130
rect 8324 5175 8380 5231
rect 8408 5175 8464 5231
rect 8492 5175 8548 5231
rect 8576 5175 8632 5231
rect 8660 5175 8716 5231
rect 8744 5175 8800 5231
rect 8828 5175 8884 5231
rect 8324 5094 8380 5150
rect 8408 5094 8464 5150
rect 8492 5094 8548 5150
rect 8576 5094 8632 5150
rect 8660 5094 8716 5150
rect 8744 5094 8800 5150
rect 8828 5094 8884 5150
rect -714 4993 -658 5049
rect -626 4993 -570 5049
rect -538 4993 -482 5049
rect -450 4993 -394 5049
rect -362 4993 -306 5049
rect -274 4993 -218 5049
rect -186 4993 -130 5049
rect -714 4912 -658 4968
rect -626 4912 -570 4968
rect -538 4912 -482 4968
rect -450 4912 -394 4968
rect -362 4912 -306 4968
rect -274 4912 -218 4968
rect -186 4912 -130 4968
rect 8324 5013 8380 5069
rect 8408 5013 8464 5069
rect 8492 5013 8548 5069
rect 8576 5013 8632 5069
rect 8660 5013 8716 5069
rect 8744 5013 8800 5069
rect 8828 5013 8884 5069
rect -714 4831 -658 4887
rect -626 4831 -570 4887
rect -538 4831 -482 4887
rect -450 4831 -394 4887
rect -362 4831 -306 4887
rect -274 4831 -218 4887
rect -186 4831 -130 4887
rect 8324 4932 8380 4988
rect 8408 4932 8464 4988
rect 8492 4932 8548 4988
rect 8576 4932 8632 4988
rect 8660 4932 8716 4988
rect 8744 4932 8800 4988
rect 8828 4932 8884 4988
rect 8324 4851 8380 4907
rect 8408 4851 8464 4907
rect 8492 4851 8548 4907
rect 8576 4851 8632 4907
rect 8660 4851 8716 4907
rect 8744 4851 8800 4907
rect 8828 4851 8884 4907
rect -714 4750 -658 4806
rect -626 4750 -570 4806
rect -538 4750 -482 4806
rect -450 4750 -394 4806
rect -362 4750 -306 4806
rect -274 4750 -218 4806
rect -186 4750 -130 4806
rect -714 4669 -658 4725
rect -626 4669 -570 4725
rect -538 4669 -482 4725
rect -450 4669 -394 4725
rect -362 4669 -306 4725
rect -274 4669 -218 4725
rect -186 4669 -130 4725
rect -714 4588 -658 4644
rect -626 4588 -570 4644
rect -538 4588 -482 4644
rect -450 4588 -394 4644
rect -362 4588 -306 4644
rect -274 4588 -218 4644
rect -186 4588 -130 4644
rect -714 4507 -658 4563
rect -626 4507 -570 4563
rect -538 4507 -482 4563
rect -450 4507 -394 4563
rect -362 4507 -306 4563
rect -274 4507 -218 4563
rect -186 4507 -130 4563
rect -714 4426 -658 4482
rect -626 4426 -570 4482
rect -538 4426 -482 4482
rect -450 4426 -394 4482
rect -362 4426 -306 4482
rect -274 4426 -218 4482
rect -186 4426 -130 4482
rect -714 4345 -658 4401
rect -626 4345 -570 4401
rect -538 4345 -482 4401
rect -450 4345 -394 4401
rect -362 4345 -306 4401
rect -274 4345 -218 4401
rect -186 4345 -130 4401
rect -714 4264 -658 4320
rect -626 4264 -570 4320
rect -538 4264 -482 4320
rect -450 4264 -394 4320
rect -362 4264 -306 4320
rect -274 4264 -218 4320
rect -186 4264 -130 4320
rect -714 4183 -658 4239
rect -626 4183 -570 4239
rect -538 4183 -482 4239
rect -450 4183 -394 4239
rect -362 4183 -306 4239
rect -274 4183 -218 4239
rect -186 4183 -130 4239
rect -714 4102 -658 4158
rect -626 4102 -570 4158
rect -538 4102 -482 4158
rect -450 4102 -394 4158
rect -362 4102 -306 4158
rect -274 4102 -218 4158
rect -186 4102 -130 4158
rect -714 4021 -658 4077
rect -626 4021 -570 4077
rect -538 4021 -482 4077
rect -450 4021 -394 4077
rect -362 4021 -306 4077
rect -274 4021 -218 4077
rect -186 4021 -130 4077
rect -714 3940 -658 3996
rect -626 3940 -570 3996
rect -538 3940 -482 3996
rect -450 3940 -394 3996
rect -362 3940 -306 3996
rect -274 3940 -218 3996
rect -186 3940 -130 3996
rect -714 3859 -658 3915
rect -626 3859 -570 3915
rect -538 3859 -482 3915
rect -450 3859 -394 3915
rect -362 3859 -306 3915
rect -274 3859 -218 3915
rect -186 3859 -130 3915
rect -714 3778 -658 3834
rect -626 3778 -570 3834
rect -538 3778 -482 3834
rect -450 3778 -394 3834
rect -362 3778 -306 3834
rect -274 3778 -218 3834
rect -186 3778 -130 3834
rect -714 3697 -658 3753
rect -626 3697 -570 3753
rect -538 3697 -482 3753
rect -450 3697 -394 3753
rect -362 3697 -306 3753
rect -274 3697 -218 3753
rect -186 3697 -130 3753
rect -714 3616 -658 3672
rect -626 3616 -570 3672
rect -538 3616 -482 3672
rect -450 3616 -394 3672
rect -362 3616 -306 3672
rect -274 3616 -218 3672
rect -186 3616 -130 3672
rect -714 3535 -658 3591
rect -626 3535 -570 3591
rect -538 3535 -482 3591
rect -450 3535 -394 3591
rect -362 3535 -306 3591
rect -274 3535 -218 3591
rect -186 3535 -130 3591
rect 8324 4770 8380 4826
rect 8408 4770 8464 4826
rect 8492 4770 8548 4826
rect 8576 4770 8632 4826
rect 8660 4770 8716 4826
rect 8744 4770 8800 4826
rect 8828 4770 8884 4826
rect 8324 4689 8380 4745
rect 8408 4689 8464 4745
rect 8492 4689 8548 4745
rect 8576 4689 8632 4745
rect 8660 4689 8716 4745
rect 8744 4689 8800 4745
rect 8828 4689 8884 4745
rect 8324 4608 8380 4664
rect 8408 4608 8464 4664
rect 8492 4608 8548 4664
rect 8576 4608 8632 4664
rect 8660 4608 8716 4664
rect 8744 4608 8800 4664
rect 8828 4608 8884 4664
rect 8324 4527 8380 4583
rect 8408 4527 8464 4583
rect 8492 4527 8548 4583
rect 8576 4527 8632 4583
rect 8660 4527 8716 4583
rect 8744 4527 8800 4583
rect 8828 4527 8884 4583
rect 8324 4446 8380 4502
rect 8408 4446 8464 4502
rect 8492 4446 8548 4502
rect 8576 4446 8632 4502
rect 8660 4446 8716 4502
rect 8744 4446 8800 4502
rect 8828 4446 8884 4502
rect 8324 4365 8380 4421
rect 8408 4365 8464 4421
rect 8492 4365 8548 4421
rect 8576 4365 8632 4421
rect 8660 4365 8716 4421
rect 8744 4365 8800 4421
rect 8828 4365 8884 4421
rect 8324 4284 8380 4340
rect 8408 4284 8464 4340
rect 8492 4284 8548 4340
rect 8576 4284 8632 4340
rect 8660 4284 8716 4340
rect 8744 4284 8800 4340
rect 8828 4284 8884 4340
rect 8324 4203 8380 4259
rect 8408 4203 8464 4259
rect 8492 4203 8548 4259
rect 8576 4203 8632 4259
rect 8660 4203 8716 4259
rect 8744 4203 8800 4259
rect 8828 4203 8884 4259
rect 8324 4122 8380 4178
rect 8408 4122 8464 4178
rect 8492 4122 8548 4178
rect 8576 4122 8632 4178
rect 8660 4122 8716 4178
rect 8744 4122 8800 4178
rect 8828 4122 8884 4178
rect 8324 4041 8380 4097
rect 8408 4041 8464 4097
rect 8492 4041 8548 4097
rect 8576 4041 8632 4097
rect 8660 4041 8716 4097
rect 8744 4041 8800 4097
rect 8828 4041 8884 4097
rect 8324 3960 8380 4016
rect 8408 3960 8464 4016
rect 8492 3960 8548 4016
rect 8576 3960 8632 4016
rect 8660 3960 8716 4016
rect 8744 3960 8800 4016
rect 8828 3960 8884 4016
rect 8324 3879 8380 3935
rect 8408 3879 8464 3935
rect 8492 3879 8548 3935
rect 8576 3879 8632 3935
rect 8660 3879 8716 3935
rect 8744 3879 8800 3935
rect 8828 3879 8884 3935
rect 8324 3798 8380 3854
rect 8408 3798 8464 3854
rect 8492 3798 8548 3854
rect 8576 3798 8632 3854
rect 8660 3798 8716 3854
rect 8744 3798 8800 3854
rect 8828 3798 8884 3854
rect 8324 3717 8380 3773
rect 8408 3717 8464 3773
rect 8492 3717 8548 3773
rect 8576 3717 8632 3773
rect 8660 3717 8716 3773
rect 8744 3717 8800 3773
rect 8828 3717 8884 3773
rect 8324 3636 8380 3692
rect 8408 3636 8464 3692
rect 8492 3636 8548 3692
rect 8576 3636 8632 3692
rect 8660 3636 8716 3692
rect 8744 3636 8800 3692
rect 8828 3636 8884 3692
rect 8324 3555 8380 3611
rect 8408 3555 8464 3611
rect 8492 3555 8548 3611
rect 8576 3555 8632 3611
rect 8660 3555 8716 3611
rect 8744 3555 8800 3611
rect 8828 3555 8884 3611
rect -714 3454 -658 3510
rect -626 3454 -570 3510
rect -538 3454 -482 3510
rect -450 3454 -394 3510
rect -362 3454 -306 3510
rect -274 3454 -218 3510
rect -186 3454 -130 3510
rect -714 3373 -658 3429
rect -626 3373 -570 3429
rect -538 3373 -482 3429
rect -450 3373 -394 3429
rect -362 3373 -306 3429
rect -274 3373 -218 3429
rect -186 3373 -130 3429
rect -714 3292 -658 3348
rect -626 3292 -570 3348
rect -538 3292 -482 3348
rect -450 3292 -394 3348
rect -362 3292 -306 3348
rect -274 3292 -218 3348
rect -186 3292 -130 3348
rect -714 3211 -658 3267
rect -626 3211 -570 3267
rect -538 3211 -482 3267
rect -450 3211 -394 3267
rect -362 3211 -306 3267
rect -274 3211 -218 3267
rect -186 3211 -130 3267
<< metal3 >>
rect -722 20547 -122 20566
rect -722 20491 -711 20547
rect -655 20491 -625 20547
rect -569 20491 -539 20547
rect -483 20491 -453 20547
rect -397 20491 -367 20547
rect -311 20491 -281 20547
rect -225 20491 -195 20547
rect -139 20491 -122 20547
rect -722 20455 -122 20491
rect -722 20399 -711 20455
rect -655 20399 -625 20455
rect -569 20399 -539 20455
rect -483 20399 -453 20455
rect -397 20399 -367 20455
rect -311 20399 -281 20455
rect -225 20399 -195 20455
rect -139 20399 -122 20455
rect -722 20363 -122 20399
rect -722 20307 -711 20363
rect -655 20307 -625 20363
rect -569 20307 -539 20363
rect -483 20307 -453 20363
rect -397 20307 -367 20363
rect -311 20307 -281 20363
rect -225 20307 -195 20363
rect -139 20307 -122 20363
rect -722 20271 -122 20307
rect -722 20215 -711 20271
rect -655 20215 -625 20271
rect -569 20215 -539 20271
rect -483 20215 -453 20271
rect -397 20215 -367 20271
rect -311 20215 -281 20271
rect -225 20215 -195 20271
rect -139 20215 -122 20271
rect -722 20179 -122 20215
rect -722 20123 -711 20179
rect -655 20123 -625 20179
rect -569 20123 -539 20179
rect -483 20123 -453 20179
rect -397 20123 -367 20179
rect -311 20123 -281 20179
rect -225 20123 -195 20179
rect -139 20123 -122 20179
rect -722 20086 -122 20123
rect -722 20030 -711 20086
rect -655 20030 -625 20086
rect -569 20030 -539 20086
rect -483 20030 -453 20086
rect -397 20030 -367 20086
rect -311 20030 -281 20086
rect -225 20030 -195 20086
rect -139 20030 -122 20086
rect -722 19993 -122 20030
rect -722 19937 -711 19993
rect -655 19937 -625 19993
rect -569 19937 -539 19993
rect -483 19937 -453 19993
rect -397 19937 -367 19993
rect -311 19937 -281 19993
rect -225 19937 -195 19993
rect -139 19937 -122 19993
rect -722 12833 -122 19937
rect 1094 20550 1670 20567
rect 1094 20494 1106 20550
rect 1162 20494 1188 20550
rect 1244 20494 1270 20550
rect 1326 20494 1352 20550
rect 1408 20494 1434 20550
rect 1490 20494 1516 20550
rect 1572 20494 1598 20550
rect 1654 20494 1670 20550
rect 1094 20470 1670 20494
rect 1094 20414 1106 20470
rect 1162 20414 1188 20470
rect 1244 20414 1270 20470
rect 1326 20414 1352 20470
rect 1408 20414 1434 20470
rect 1490 20414 1516 20470
rect 1572 20414 1598 20470
rect 1654 20414 1670 20470
rect 1094 20390 1670 20414
rect 1094 20334 1106 20390
rect 1162 20334 1188 20390
rect 1244 20334 1270 20390
rect 1326 20334 1352 20390
rect 1408 20334 1434 20390
rect 1490 20334 1516 20390
rect 1572 20334 1598 20390
rect 1654 20334 1670 20390
rect 1094 20310 1670 20334
rect 1094 20254 1106 20310
rect 1162 20254 1188 20310
rect 1244 20254 1270 20310
rect 1326 20254 1352 20310
rect 1408 20254 1434 20310
rect 1490 20254 1516 20310
rect 1572 20254 1598 20310
rect 1654 20254 1670 20310
rect 1094 20230 1670 20254
rect 1094 20174 1106 20230
rect 1162 20174 1188 20230
rect 1244 20174 1270 20230
rect 1326 20174 1352 20230
rect 1408 20174 1434 20230
rect 1490 20174 1516 20230
rect 1572 20174 1598 20230
rect 1654 20174 1670 20230
rect 1094 20149 1670 20174
rect 1094 20093 1106 20149
rect 1162 20093 1188 20149
rect 1244 20093 1270 20149
rect 1326 20093 1352 20149
rect 1408 20093 1434 20149
rect 1490 20093 1516 20149
rect 1572 20093 1598 20149
rect 1654 20093 1670 20149
rect 1094 20068 1670 20093
rect 1094 20012 1106 20068
rect 1162 20012 1188 20068
rect 1244 20012 1270 20068
rect 1326 20012 1352 20068
rect 1408 20012 1434 20068
rect 1490 20012 1516 20068
rect 1572 20012 1598 20068
rect 1654 20012 1670 20068
rect 1094 19987 1670 20012
rect 1094 19931 1106 19987
rect 1162 19931 1188 19987
rect 1244 19931 1270 19987
rect 1326 19931 1352 19987
rect 1408 19931 1434 19987
rect 1490 19931 1516 19987
rect 1572 19931 1598 19987
rect 1654 19931 1670 19987
rect 1094 19906 1670 19931
rect 1094 19850 1106 19906
rect 1162 19850 1188 19906
rect 1244 19850 1270 19906
rect 1326 19850 1352 19906
rect 1408 19850 1434 19906
rect 1490 19850 1516 19906
rect 1572 19850 1598 19906
rect 1654 19850 1670 19906
rect 1094 19825 1670 19850
rect 1094 19769 1106 19825
rect 1162 19769 1188 19825
rect 1244 19769 1270 19825
rect 1326 19769 1352 19825
rect 1408 19769 1434 19825
rect 1490 19769 1516 19825
rect 1572 19769 1598 19825
rect 1654 19769 1670 19825
rect 1094 19744 1670 19769
rect 1094 19688 1106 19744
rect 1162 19688 1188 19744
rect 1244 19688 1270 19744
rect 1326 19688 1352 19744
rect 1408 19688 1434 19744
rect 1490 19688 1516 19744
rect 1572 19688 1598 19744
rect 1654 19688 1670 19744
rect 1094 19663 1670 19688
rect 1094 19607 1106 19663
rect 1162 19607 1188 19663
rect 1244 19607 1270 19663
rect 1326 19607 1352 19663
rect 1408 19607 1434 19663
rect 1490 19607 1516 19663
rect 1572 19607 1598 19663
rect 1654 19607 1670 19663
rect 1094 19582 1670 19607
rect 1094 19526 1106 19582
rect 1162 19526 1188 19582
rect 1244 19526 1270 19582
rect 1326 19526 1352 19582
rect 1408 19526 1434 19582
rect 1490 19526 1516 19582
rect 1572 19526 1598 19582
rect 1654 19526 1670 19582
rect 1094 19501 1670 19526
rect 1094 19445 1106 19501
rect 1162 19445 1188 19501
rect 1244 19445 1270 19501
rect 1326 19445 1352 19501
rect 1408 19445 1434 19501
rect 1490 19445 1516 19501
rect 1572 19445 1598 19501
rect 1654 19445 1670 19501
rect 1094 19420 1670 19445
rect 1094 19364 1106 19420
rect 1162 19364 1188 19420
rect 1244 19364 1270 19420
rect 1326 19364 1352 19420
rect 1408 19364 1434 19420
rect 1490 19364 1516 19420
rect 1572 19364 1598 19420
rect 1654 19364 1670 19420
rect 1094 19339 1670 19364
rect 1094 19283 1106 19339
rect 1162 19283 1188 19339
rect 1244 19283 1270 19339
rect 1326 19283 1352 19339
rect 1408 19283 1434 19339
rect 1490 19283 1516 19339
rect 1572 19283 1598 19339
rect 1654 19283 1670 19339
rect 1094 19258 1670 19283
rect 1094 19202 1106 19258
rect 1162 19202 1188 19258
rect 1244 19202 1270 19258
rect 1326 19202 1352 19258
rect 1408 19202 1434 19258
rect 1490 19202 1516 19258
rect 1572 19202 1598 19258
rect 1654 19202 1670 19258
rect 1094 19177 1670 19202
rect 1094 19121 1106 19177
rect 1162 19121 1188 19177
rect 1244 19121 1270 19177
rect 1326 19121 1352 19177
rect 1408 19121 1434 19177
rect 1490 19121 1516 19177
rect 1572 19121 1598 19177
rect 1654 19121 1670 19177
rect 1094 19096 1670 19121
rect 1094 19040 1106 19096
rect 1162 19040 1188 19096
rect 1244 19040 1270 19096
rect 1326 19040 1352 19096
rect 1408 19040 1434 19096
rect 1490 19040 1516 19096
rect 1572 19040 1598 19096
rect 1654 19040 1670 19096
rect 211 18409 217 18445
rect -722 12777 -714 12833
rect -658 12777 -626 12833
rect -570 12777 -538 12833
rect -482 12777 -450 12833
rect -394 12777 -362 12833
rect -306 12777 -274 12833
rect -218 12777 -186 12833
rect -130 12777 -122 12833
rect -722 12753 -122 12777
rect -722 12697 -714 12753
rect -658 12697 -626 12753
rect -570 12697 -538 12753
rect -482 12697 -450 12753
rect -394 12697 -362 12753
rect -306 12697 -274 12753
rect -218 12697 -186 12753
rect -130 12697 -122 12753
rect -722 12673 -122 12697
rect -722 12617 -714 12673
rect -658 12617 -626 12673
rect -570 12617 -538 12673
rect -482 12617 -450 12673
rect -394 12617 -362 12673
rect -306 12617 -274 12673
rect -218 12617 -186 12673
rect -130 12617 -122 12673
rect -722 12593 -122 12617
rect -722 12537 -714 12593
rect -658 12537 -626 12593
rect -570 12537 -538 12593
rect -482 12537 -450 12593
rect -394 12537 -362 12593
rect -306 12537 -274 12593
rect -218 12537 -186 12593
rect -130 12537 -122 12593
rect -722 12513 -122 12537
rect -722 12457 -714 12513
rect -658 12457 -626 12513
rect -570 12457 -538 12513
rect -482 12457 -450 12513
rect -394 12457 -362 12513
rect -306 12457 -274 12513
rect -218 12457 -186 12513
rect -130 12457 -122 12513
rect -722 12433 -122 12457
rect -722 12377 -714 12433
rect -658 12377 -626 12433
rect -570 12377 -538 12433
rect -482 12377 -450 12433
rect -394 12377 -362 12433
rect -306 12377 -274 12433
rect -218 12377 -186 12433
rect -130 12377 -122 12433
rect -722 12353 -122 12377
rect -722 12297 -714 12353
rect -658 12297 -626 12353
rect -570 12297 -538 12353
rect -482 12297 -450 12353
rect -394 12297 -362 12353
rect -306 12297 -274 12353
rect -218 12297 -186 12353
rect -130 12297 -122 12353
rect -722 12273 -122 12297
rect -722 12217 -714 12273
rect -658 12217 -626 12273
rect -570 12217 -538 12273
rect -482 12217 -450 12273
rect -394 12217 -362 12273
rect -306 12217 -274 12273
rect -218 12217 -186 12273
rect -130 12217 -122 12273
rect -722 12193 -122 12217
rect -2517 12168 -2131 12181
rect -2517 12112 -2511 12168
rect -2455 12112 -2405 12168
rect -2349 12112 -2299 12168
rect -2243 12112 -2193 12168
rect -2137 12112 -2131 12168
rect -2517 12085 -2131 12112
rect -2517 12029 -2511 12085
rect -2455 12029 -2405 12085
rect -2349 12029 -2299 12085
rect -2243 12029 -2193 12085
rect -2137 12029 -2131 12085
rect -2517 12001 -2131 12029
rect -2517 11945 -2511 12001
rect -2455 11945 -2405 12001
rect -2349 11945 -2299 12001
rect -2243 11945 -2193 12001
rect -2137 11945 -2131 12001
rect -4308 2988 -3745 11945
rect -2517 11917 -2131 11945
rect -2517 11861 -2511 11917
rect -2455 11861 -2405 11917
rect -2349 11861 -2299 11917
rect -2243 11861 -2193 11917
rect -2137 11861 -2131 11917
rect -2517 11833 -2131 11861
rect -2517 11777 -2511 11833
rect -2455 11777 -2405 11833
rect -2349 11777 -2299 11833
rect -2243 11777 -2193 11833
rect -2137 11777 -2131 11833
rect -2517 11749 -2131 11777
rect -2517 11693 -2511 11749
rect -2455 11693 -2405 11749
rect -2349 11693 -2299 11749
rect -2243 11693 -2193 11749
rect -2137 11693 -2131 11749
rect -2517 11242 -2131 11693
rect -722 12137 -714 12193
rect -658 12137 -626 12193
rect -570 12137 -538 12193
rect -482 12137 -450 12193
rect -394 12137 -362 12193
rect -306 12137 -274 12193
rect -218 12137 -186 12193
rect -130 12137 -122 12193
rect -722 12113 -122 12137
rect -722 12057 -714 12113
rect -658 12057 -626 12113
rect -570 12057 -538 12113
rect -482 12057 -450 12113
rect -394 12057 -362 12113
rect -306 12057 -274 12113
rect -218 12057 -186 12113
rect -130 12057 -122 12113
rect -722 12033 -122 12057
rect -722 11977 -714 12033
rect -658 11977 -626 12033
rect -570 11977 -538 12033
rect -482 11977 -450 12033
rect -394 11977 -362 12033
rect -306 11977 -274 12033
rect -218 11977 -186 12033
rect -130 11977 -122 12033
rect -722 11953 -122 11977
rect -722 11897 -714 11953
rect -658 11897 -626 11953
rect -570 11897 -538 11953
rect -482 11897 -450 11953
rect -394 11897 -362 11953
rect -306 11897 -274 11953
rect -218 11897 -186 11953
rect -130 11897 -122 11953
rect -722 11873 -122 11897
rect -722 11817 -714 11873
rect -658 11817 -626 11873
rect -570 11817 -538 11873
rect -482 11817 -450 11873
rect -394 11817 -362 11873
rect -306 11817 -274 11873
rect -218 11817 -186 11873
rect -130 11817 -122 11873
rect -722 11793 -122 11817
rect -722 11737 -714 11793
rect -658 11737 -626 11793
rect -570 11737 -538 11793
rect -482 11737 -450 11793
rect -394 11737 -362 11793
rect -306 11737 -274 11793
rect -218 11737 -186 11793
rect -130 11737 -122 11793
rect -722 11713 -122 11737
rect -722 11657 -714 11713
rect -658 11657 -626 11713
rect -570 11657 -538 11713
rect -482 11657 -450 11713
rect -394 11657 -362 11713
rect -306 11657 -274 11713
rect -218 11657 -186 11713
rect -130 11657 -122 11713
rect -722 11633 -122 11657
rect -722 11577 -714 11633
rect -658 11577 -626 11633
rect -570 11577 -538 11633
rect -482 11577 -450 11633
rect -394 11577 -362 11633
rect -306 11577 -274 11633
rect -218 11577 -186 11633
rect -130 11577 -122 11633
rect -722 11553 -122 11577
rect -722 11497 -714 11553
rect -658 11497 -626 11553
rect -570 11497 -538 11553
rect -482 11497 -450 11553
rect -394 11497 -362 11553
rect -306 11497 -274 11553
rect -218 11497 -186 11553
rect -130 11497 -122 11553
rect -722 11473 -122 11497
rect -722 11417 -714 11473
rect -658 11417 -626 11473
rect -570 11417 -538 11473
rect -482 11417 -450 11473
rect -394 11417 -362 11473
rect -306 11417 -274 11473
rect -218 11417 -186 11473
rect -130 11417 -122 11473
rect -722 11393 -122 11417
tri -3405 4725 -3404 4726 se
tri -2860 4725 -2859 4726 sw
rect -1598 3526 -1038 11355
rect -722 11337 -714 11393
rect -658 11337 -626 11393
rect -570 11337 -538 11393
rect -482 11337 -450 11393
rect -394 11337 -362 11393
rect -306 11337 -274 11393
rect -218 11337 -186 11393
rect -130 11337 -122 11393
rect -722 11313 -122 11337
rect -722 11257 -714 11313
rect -658 11257 -626 11313
rect -570 11257 -538 11313
rect -482 11257 -450 11313
rect -394 11257 -362 11313
rect -306 11257 -274 11313
rect -218 11257 -186 11313
rect -130 11257 -122 11313
rect -722 11233 -122 11257
rect -722 11177 -714 11233
rect -658 11177 -626 11233
rect -570 11177 -538 11233
rect -482 11177 -450 11233
rect -394 11177 -362 11233
rect -306 11177 -274 11233
rect -218 11177 -186 11233
rect -130 11177 -122 11233
rect -722 11153 -122 11177
rect -722 11097 -714 11153
rect -658 11097 -626 11153
rect -570 11097 -538 11153
rect -482 11097 -450 11153
rect -394 11097 -362 11153
rect -306 11097 -274 11153
rect -218 11097 -186 11153
rect -130 11097 -122 11153
rect -722 11073 -122 11097
rect -722 11017 -714 11073
rect -658 11017 -626 11073
rect -570 11017 -538 11073
rect -482 11017 -450 11073
rect -394 11017 -362 11073
rect -306 11017 -274 11073
rect -218 11017 -186 11073
rect -130 11017 -122 11073
rect -722 10993 -122 11017
rect -722 10937 -714 10993
rect -658 10937 -626 10993
rect -570 10937 -538 10993
rect -482 10937 -450 10993
rect -394 10937 -362 10993
rect -306 10937 -274 10993
rect -218 10937 -186 10993
rect -130 10937 -122 10993
rect -722 10913 -122 10937
rect -722 10857 -714 10913
rect -658 10857 -626 10913
rect -570 10857 -538 10913
rect -482 10857 -450 10913
rect -394 10857 -362 10913
rect -306 10857 -274 10913
rect -218 10857 -186 10913
rect -130 10857 -122 10913
rect -722 10833 -122 10857
rect -722 10777 -714 10833
rect -658 10777 -626 10833
rect -570 10777 -538 10833
rect -482 10777 -450 10833
rect -394 10777 -362 10833
rect -306 10777 -274 10833
rect -218 10777 -186 10833
rect -130 10777 -122 10833
rect -722 10753 -122 10777
rect -722 10697 -714 10753
rect -658 10697 -626 10753
rect -570 10697 -538 10753
rect -482 10697 -450 10753
rect -394 10697 -362 10753
rect -306 10697 -274 10753
rect -218 10697 -186 10753
rect -130 10697 -122 10753
rect -722 10673 -122 10697
rect -722 10617 -714 10673
rect -658 10617 -626 10673
rect -570 10617 -538 10673
rect -482 10617 -450 10673
rect -394 10617 -362 10673
rect -306 10617 -274 10673
rect -218 10617 -186 10673
rect -130 10617 -122 10673
rect -722 10593 -122 10617
rect -722 10537 -714 10593
rect -658 10537 -626 10593
rect -570 10537 -538 10593
rect -482 10537 -450 10593
rect -394 10537 -362 10593
rect -306 10537 -274 10593
rect -218 10537 -186 10593
rect -130 10537 -122 10593
rect -722 10513 -122 10537
rect -722 10457 -714 10513
rect -658 10457 -626 10513
rect -570 10457 -538 10513
rect -482 10457 -450 10513
rect -394 10457 -362 10513
rect -306 10457 -274 10513
rect -218 10457 -186 10513
rect -130 10457 -122 10513
rect -722 10433 -122 10457
rect -722 10377 -714 10433
rect -658 10377 -626 10433
rect -570 10377 -538 10433
rect -482 10377 -450 10433
rect -394 10377 -362 10433
rect -306 10377 -274 10433
rect -218 10377 -186 10433
rect -130 10377 -122 10433
rect -722 10353 -122 10377
rect -722 10297 -714 10353
rect -658 10297 -626 10353
rect -570 10297 -538 10353
rect -482 10297 -450 10353
rect -394 10297 -362 10353
rect -306 10297 -274 10353
rect -218 10297 -186 10353
rect -130 10297 -122 10353
rect -722 10273 -122 10297
rect -722 10217 -714 10273
rect -658 10217 -626 10273
rect -570 10217 -538 10273
rect -482 10217 -450 10273
rect -394 10217 -362 10273
rect -306 10217 -274 10273
rect -218 10217 -186 10273
rect -130 10217 -122 10273
rect -722 10193 -122 10217
rect -722 10137 -714 10193
rect -658 10137 -626 10193
rect -570 10137 -538 10193
rect -482 10137 -450 10193
rect -394 10137 -362 10193
rect -306 10137 -274 10193
rect -218 10137 -186 10193
rect -130 10137 -122 10193
rect -722 10113 -122 10137
rect -722 10057 -714 10113
rect -658 10057 -626 10113
rect -570 10057 -538 10113
rect -482 10057 -450 10113
rect -394 10057 -362 10113
rect -306 10057 -274 10113
rect -218 10057 -186 10113
rect -130 10057 -122 10113
rect -722 10033 -122 10057
rect -722 9977 -714 10033
rect -658 9977 -626 10033
rect -570 9977 -538 10033
rect -482 9977 -450 10033
rect -394 9977 -362 10033
rect -306 9977 -274 10033
rect -218 9977 -186 10033
rect -130 9977 -122 10033
rect -722 9953 -122 9977
rect -722 9897 -714 9953
rect -658 9897 -626 9953
rect -570 9897 -538 9953
rect -482 9897 -450 9953
rect -394 9897 -362 9953
rect -306 9897 -274 9953
rect -218 9897 -186 9953
rect -130 9897 -122 9953
rect -722 9873 -122 9897
rect -722 9817 -714 9873
rect -658 9817 -626 9873
rect -570 9817 -538 9873
rect -482 9817 -450 9873
rect -394 9817 -362 9873
rect -306 9817 -274 9873
rect -218 9817 -186 9873
rect -130 9817 -122 9873
rect -722 9793 -122 9817
rect -722 9737 -714 9793
rect -658 9737 -626 9793
rect -570 9737 -538 9793
rect -482 9737 -450 9793
rect -394 9737 -362 9793
rect -306 9737 -274 9793
rect -218 9737 -186 9793
rect -130 9737 -122 9793
rect -722 9713 -122 9737
rect -722 9657 -714 9713
rect -658 9657 -626 9713
rect -570 9657 -538 9713
rect -482 9657 -450 9713
rect -394 9657 -362 9713
rect -306 9657 -274 9713
rect -218 9657 -186 9713
rect -130 9657 -122 9713
rect -722 9633 -122 9657
rect -722 9577 -714 9633
rect -658 9577 -626 9633
rect -570 9577 -538 9633
rect -482 9577 -450 9633
rect -394 9577 -362 9633
rect -306 9577 -274 9633
rect -218 9577 -186 9633
rect -130 9577 -122 9633
rect -722 9553 -122 9577
rect -722 9497 -714 9553
rect -658 9497 -626 9553
rect -570 9497 -538 9553
rect -482 9497 -450 9553
rect -394 9497 -362 9553
rect -306 9497 -274 9553
rect -218 9497 -186 9553
rect -130 9497 -122 9553
rect -722 9473 -122 9497
rect -722 9417 -714 9473
rect -658 9417 -626 9473
rect -570 9417 -538 9473
rect -482 9417 -450 9473
rect -394 9417 -362 9473
rect -306 9417 -274 9473
rect -218 9417 -186 9473
rect -130 9417 -122 9473
rect -722 9393 -122 9417
rect -722 9337 -714 9393
rect -658 9337 -626 9393
rect -570 9337 -538 9393
rect -482 9337 -450 9393
rect -394 9337 -362 9393
rect -306 9337 -274 9393
rect -218 9337 -186 9393
rect -130 9337 -122 9393
rect -722 9313 -122 9337
rect -722 9257 -714 9313
rect -658 9257 -626 9313
rect -570 9257 -538 9313
rect -482 9257 -450 9313
rect -394 9257 -362 9313
rect -306 9257 -274 9313
rect -218 9257 -186 9313
rect -130 9257 -122 9313
rect -722 9233 -122 9257
rect -722 9177 -714 9233
rect -658 9177 -626 9233
rect -570 9177 -538 9233
rect -482 9177 -450 9233
rect -394 9177 -362 9233
rect -306 9177 -274 9233
rect -218 9177 -186 9233
rect -130 9177 -122 9233
rect -722 9153 -122 9177
rect -722 9097 -714 9153
rect -658 9097 -626 9153
rect -570 9097 -538 9153
rect -482 9097 -450 9153
rect -394 9097 -362 9153
rect -306 9097 -274 9153
rect -218 9097 -186 9153
rect -130 9097 -122 9153
rect -722 9073 -122 9097
rect -722 9017 -714 9073
rect -658 9017 -626 9073
rect -570 9017 -538 9073
rect -482 9017 -450 9073
rect -394 9017 -362 9073
rect -306 9017 -274 9073
rect -218 9017 -186 9073
rect -130 9017 -122 9073
rect -722 8993 -122 9017
rect -722 8937 -714 8993
rect -658 8937 -626 8993
rect -570 8937 -538 8993
rect -482 8937 -450 8993
rect -394 8937 -362 8993
rect -306 8937 -274 8993
rect -218 8937 -186 8993
rect -130 8937 -122 8993
rect -722 8913 -122 8937
rect -722 8857 -714 8913
rect -658 8857 -626 8913
rect -570 8857 -538 8913
rect -482 8857 -450 8913
rect -394 8857 -362 8913
rect -306 8857 -274 8913
rect -218 8857 -186 8913
rect -130 8857 -122 8913
rect -722 8833 -122 8857
rect -722 8777 -714 8833
rect -658 8777 -626 8833
rect -570 8777 -538 8833
rect -482 8777 -450 8833
rect -394 8777 -362 8833
rect -306 8777 -274 8833
rect -218 8777 -186 8833
rect -130 8777 -122 8833
rect -722 8753 -122 8777
rect -722 8697 -714 8753
rect -658 8697 -626 8753
rect -570 8697 -538 8753
rect -482 8697 -450 8753
rect -394 8697 -362 8753
rect -306 8697 -274 8753
rect -218 8697 -186 8753
rect -130 8697 -122 8753
rect -722 8673 -122 8697
rect -722 8617 -714 8673
rect -658 8617 -626 8673
rect -570 8617 -538 8673
rect -482 8617 -450 8673
rect -394 8617 -362 8673
rect -306 8617 -274 8673
rect -218 8617 -186 8673
rect -130 8617 -122 8673
rect -722 8593 -122 8617
rect -722 8537 -714 8593
rect -658 8537 -626 8593
rect -570 8537 -538 8593
rect -482 8537 -450 8593
rect -394 8537 -362 8593
rect -306 8537 -274 8593
rect -218 8537 -186 8593
rect -130 8537 -122 8593
rect -722 8513 -122 8537
rect -722 8457 -714 8513
rect -658 8457 -626 8513
rect -570 8457 -538 8513
rect -482 8457 -450 8513
rect -394 8457 -362 8513
rect -306 8457 -274 8513
rect -218 8457 -186 8513
rect -130 8457 -122 8513
rect -722 8433 -122 8457
rect -722 8377 -714 8433
rect -658 8377 -626 8433
rect -570 8377 -538 8433
rect -482 8377 -450 8433
rect -394 8377 -362 8433
rect -306 8377 -274 8433
rect -218 8377 -186 8433
rect -130 8377 -122 8433
rect -722 8353 -122 8377
rect -722 8297 -714 8353
rect -658 8297 -626 8353
rect -570 8297 -538 8353
rect -482 8297 -450 8353
rect -394 8297 -362 8353
rect -306 8297 -274 8353
rect -218 8297 -186 8353
rect -130 8297 -122 8353
rect -722 8273 -122 8297
rect -722 8217 -714 8273
rect -658 8217 -626 8273
rect -570 8217 -538 8273
rect -482 8217 -450 8273
rect -394 8217 -362 8273
rect -306 8217 -274 8273
rect -218 8217 -186 8273
rect -130 8217 -122 8273
rect -722 8193 -122 8217
rect -722 8137 -714 8193
rect -658 8137 -626 8193
rect -570 8137 -538 8193
rect -482 8137 -450 8193
rect -394 8137 -362 8193
rect -306 8137 -274 8193
rect -218 8137 -186 8193
rect -130 8137 -122 8193
rect -722 8113 -122 8137
rect -722 8057 -714 8113
rect -658 8057 -626 8113
rect -570 8057 -538 8113
rect -482 8057 -450 8113
rect -394 8057 -362 8113
rect -306 8057 -274 8113
rect -218 8057 -186 8113
rect -130 8057 -122 8113
rect -722 8033 -122 8057
rect -722 7977 -714 8033
rect -658 7977 -626 8033
rect -570 7977 -538 8033
rect -482 7977 -450 8033
rect -394 7977 -362 8033
rect -306 7977 -274 8033
rect -218 7977 -186 8033
rect -130 7977 -122 8033
rect -722 7953 -122 7977
rect -722 7897 -714 7953
rect -658 7897 -626 7953
rect -570 7897 -538 7953
rect -482 7897 -450 7953
rect -394 7897 -362 7953
rect -306 7897 -274 7953
rect -218 7897 -186 7953
rect -130 7897 -122 7953
rect -722 7873 -122 7897
rect -722 7817 -714 7873
rect -658 7817 -626 7873
rect -570 7817 -538 7873
rect -482 7817 -450 7873
rect -394 7817 -362 7873
rect -306 7817 -274 7873
rect -218 7817 -186 7873
rect -130 7817 -122 7873
rect -722 7793 -122 7817
rect -722 7737 -714 7793
rect -658 7737 -626 7793
rect -570 7737 -538 7793
rect -482 7737 -450 7793
rect -394 7737 -362 7793
rect -306 7737 -274 7793
rect -218 7737 -186 7793
rect -130 7737 -122 7793
rect -722 7713 -122 7737
rect -722 7657 -714 7713
rect -658 7657 -626 7713
rect -570 7657 -538 7713
rect -482 7657 -450 7713
rect -394 7657 -362 7713
rect -306 7657 -274 7713
rect -218 7657 -186 7713
rect -130 7657 -122 7713
rect -722 7633 -122 7657
rect -722 7577 -714 7633
rect -658 7577 -626 7633
rect -570 7577 -538 7633
rect -482 7577 -450 7633
rect -394 7577 -362 7633
rect -306 7577 -274 7633
rect -218 7577 -186 7633
rect -130 7577 -122 7633
rect -722 7553 -122 7577
rect -722 7497 -714 7553
rect -658 7497 -626 7553
rect -570 7497 -538 7553
rect -482 7497 -450 7553
rect -394 7497 -362 7553
rect -306 7497 -274 7553
rect -218 7497 -186 7553
rect -130 7497 -122 7553
rect -722 7473 -122 7497
rect -722 7417 -714 7473
rect -658 7417 -626 7473
rect -570 7417 -538 7473
rect -482 7417 -450 7473
rect -394 7417 -362 7473
rect -306 7417 -274 7473
rect -218 7417 -186 7473
rect -130 7417 -122 7473
rect -722 7393 -122 7417
rect -722 7337 -714 7393
rect -658 7337 -626 7393
rect -570 7337 -538 7393
rect -482 7337 -450 7393
rect -394 7337 -362 7393
rect -306 7337 -274 7393
rect -218 7337 -186 7393
rect -130 7337 -122 7393
rect -722 7313 -122 7337
rect -722 7257 -714 7313
rect -658 7257 -626 7313
rect -570 7257 -538 7313
rect -482 7257 -450 7313
rect -394 7257 -362 7313
rect -306 7257 -274 7313
rect -218 7257 -186 7313
rect -130 7257 -122 7313
rect -722 7233 -122 7257
rect -722 7177 -714 7233
rect -658 7177 -626 7233
rect -570 7177 -538 7233
rect -482 7177 -450 7233
rect -394 7177 -362 7233
rect -306 7177 -274 7233
rect -218 7177 -186 7233
rect -130 7177 -122 7233
rect -722 7153 -122 7177
rect -722 7097 -714 7153
rect -658 7097 -626 7153
rect -570 7097 -538 7153
rect -482 7097 -450 7153
rect -394 7097 -362 7153
rect -306 7097 -274 7153
rect -218 7097 -186 7153
rect -130 7097 -122 7153
rect -722 7073 -122 7097
rect -722 7017 -714 7073
rect -658 7017 -626 7073
rect -570 7017 -538 7073
rect -482 7017 -450 7073
rect -394 7017 -362 7073
rect -306 7017 -274 7073
rect -218 7017 -186 7073
rect -130 7017 -122 7073
rect -722 6993 -122 7017
rect -722 6937 -714 6993
rect -658 6937 -626 6993
rect -570 6937 -538 6993
rect -482 6937 -450 6993
rect -394 6937 -362 6993
rect -306 6937 -274 6993
rect -218 6937 -186 6993
rect -130 6937 -122 6993
rect -722 6912 -122 6937
rect -722 6856 -714 6912
rect -658 6856 -626 6912
rect -570 6856 -538 6912
rect -482 6856 -450 6912
rect -394 6856 -362 6912
rect -306 6856 -274 6912
rect -218 6856 -186 6912
rect -130 6856 -122 6912
rect -722 6831 -122 6856
rect -722 6775 -714 6831
rect -658 6775 -626 6831
rect -570 6775 -538 6831
rect -482 6775 -450 6831
rect -394 6775 -362 6831
rect -306 6775 -274 6831
rect -218 6775 -186 6831
rect -130 6775 -122 6831
rect -722 6750 -122 6775
rect -722 6694 -714 6750
rect -658 6694 -626 6750
rect -570 6694 -538 6750
rect -482 6694 -450 6750
rect -394 6694 -362 6750
rect -306 6694 -274 6750
rect -218 6694 -186 6750
rect -130 6694 -122 6750
rect -722 6669 -122 6694
rect -722 6613 -714 6669
rect -658 6613 -626 6669
rect -570 6613 -538 6669
rect -482 6613 -450 6669
rect -394 6613 -362 6669
rect -306 6613 -274 6669
rect -218 6613 -186 6669
rect -130 6613 -122 6669
rect -722 6588 -122 6613
rect -722 6532 -714 6588
rect -658 6532 -626 6588
rect -570 6532 -538 6588
rect -482 6532 -450 6588
rect -394 6532 -362 6588
rect -306 6532 -274 6588
rect -218 6532 -186 6588
rect -130 6532 -122 6588
rect -722 6507 -122 6532
rect -722 6451 -714 6507
rect -658 6451 -626 6507
rect -570 6451 -538 6507
rect -482 6451 -450 6507
rect -394 6451 -362 6507
rect -306 6451 -274 6507
rect -218 6451 -186 6507
rect -130 6451 -122 6507
rect -722 6426 -122 6451
rect -722 6370 -714 6426
rect -658 6370 -626 6426
rect -570 6370 -538 6426
rect -482 6370 -450 6426
rect -394 6370 -362 6426
rect -306 6370 -274 6426
rect -218 6370 -186 6426
rect -130 6370 -122 6426
rect -722 6345 -122 6370
rect -722 6289 -714 6345
rect -658 6289 -626 6345
rect -570 6289 -538 6345
rect -482 6289 -450 6345
rect -394 6289 -362 6345
rect -306 6289 -274 6345
rect -218 6289 -186 6345
rect -130 6289 -122 6345
rect -722 6264 -122 6289
rect -722 6208 -714 6264
rect -658 6208 -626 6264
rect -570 6208 -538 6264
rect -482 6208 -450 6264
rect -394 6208 -362 6264
rect -306 6208 -274 6264
rect -218 6208 -186 6264
rect -130 6208 -122 6264
rect -722 6183 -122 6208
rect -722 6127 -714 6183
rect -658 6127 -626 6183
rect -570 6127 -538 6183
rect -482 6127 -450 6183
rect -394 6127 -362 6183
rect -306 6127 -274 6183
rect -218 6127 -186 6183
rect -130 6127 -122 6183
rect -722 6102 -122 6127
rect -722 6046 -714 6102
rect -658 6046 -626 6102
rect -570 6046 -538 6102
rect -482 6046 -450 6102
rect -394 6046 -362 6102
rect -306 6046 -274 6102
rect -218 6046 -186 6102
rect -130 6046 -122 6102
rect -722 6021 -122 6046
rect -722 5965 -714 6021
rect -658 5965 -626 6021
rect -570 5965 -538 6021
rect -482 5965 -450 6021
rect -394 5965 -362 6021
rect -306 5965 -274 6021
rect -218 5965 -186 6021
rect -130 5965 -122 6021
rect -722 5940 -122 5965
rect -722 5884 -714 5940
rect -658 5884 -626 5940
rect -570 5884 -538 5940
rect -482 5884 -450 5940
rect -394 5884 -362 5940
rect -306 5884 -274 5940
rect -218 5884 -186 5940
rect -130 5884 -122 5940
rect -722 5859 -122 5884
rect -722 5803 -714 5859
rect -658 5803 -626 5859
rect -570 5803 -538 5859
rect -482 5803 -450 5859
rect -394 5803 -362 5859
rect -306 5803 -274 5859
rect -218 5803 -186 5859
rect -130 5803 -122 5859
rect -722 5778 -122 5803
rect -722 5722 -714 5778
rect -658 5722 -626 5778
rect -570 5722 -538 5778
rect -482 5722 -450 5778
rect -394 5722 -362 5778
rect -306 5722 -274 5778
rect -218 5722 -186 5778
rect -130 5722 -122 5778
rect -722 5697 -122 5722
rect -722 5641 -714 5697
rect -658 5641 -626 5697
rect -570 5641 -538 5697
rect -482 5641 -450 5697
rect -394 5641 -362 5697
rect -306 5641 -274 5697
rect -218 5641 -186 5697
rect -130 5641 -122 5697
rect -722 5616 -122 5641
rect -722 5560 -714 5616
rect -658 5560 -626 5616
rect -570 5560 -538 5616
rect -482 5560 -450 5616
rect -394 5560 -362 5616
rect -306 5560 -274 5616
rect -218 5560 -186 5616
rect -130 5560 -122 5616
rect -722 5535 -122 5560
rect -722 5479 -714 5535
rect -658 5479 -626 5535
rect -570 5479 -538 5535
rect -482 5479 -450 5535
rect -394 5479 -362 5535
rect -306 5479 -274 5535
rect -218 5479 -186 5535
rect -130 5479 -122 5535
rect -722 5454 -122 5479
rect -722 5398 -714 5454
rect -658 5398 -626 5454
rect -570 5398 -538 5454
rect -482 5398 -450 5454
rect -394 5398 -362 5454
rect -306 5398 -274 5454
rect -218 5398 -186 5454
rect -130 5398 -122 5454
rect -722 5373 -122 5398
rect -722 5317 -714 5373
rect -658 5317 -626 5373
rect -570 5317 -538 5373
rect -482 5317 -450 5373
rect -394 5317 -362 5373
rect -306 5317 -274 5373
rect -218 5317 -186 5373
rect -130 5317 -122 5373
rect -722 5292 -122 5317
rect -722 5236 -714 5292
rect -658 5236 -626 5292
rect -570 5236 -538 5292
rect -482 5236 -450 5292
rect -394 5236 -362 5292
rect -306 5236 -274 5292
rect -218 5236 -186 5292
rect -130 5236 -122 5292
rect -722 5211 -122 5236
rect -722 5155 -714 5211
rect -658 5155 -626 5211
rect -570 5155 -538 5211
rect -482 5155 -450 5211
rect -394 5155 -362 5211
rect -306 5155 -274 5211
rect -218 5155 -186 5211
rect -130 5155 -122 5211
rect -722 5130 -122 5155
rect -722 5074 -714 5130
rect -658 5074 -626 5130
rect -570 5074 -538 5130
rect -482 5074 -450 5130
rect -394 5074 -362 5130
rect -306 5074 -274 5130
rect -218 5074 -186 5130
rect -130 5074 -122 5130
rect -722 5049 -122 5074
rect -722 4993 -714 5049
rect -658 4993 -626 5049
rect -570 4993 -538 5049
rect -482 4993 -450 5049
rect -394 4993 -362 5049
rect -306 4993 -274 5049
rect -218 4993 -186 5049
rect -130 4993 -122 5049
rect -722 4968 -122 4993
rect -722 4912 -714 4968
rect -658 4912 -626 4968
rect -570 4912 -538 4968
rect -482 4912 -450 4968
rect -394 4912 -362 4968
rect -306 4912 -274 4968
rect -218 4912 -186 4968
rect -130 4912 -122 4968
rect -722 4887 -122 4912
rect -722 4831 -714 4887
rect -658 4831 -626 4887
rect -570 4831 -538 4887
rect -482 4831 -450 4887
rect -394 4831 -362 4887
rect -306 4831 -274 4887
rect -218 4831 -186 4887
rect -130 4831 -122 4887
rect -722 4806 -122 4831
rect -722 4750 -714 4806
rect -658 4750 -626 4806
rect -570 4750 -538 4806
rect -482 4750 -450 4806
rect -394 4750 -362 4806
rect -306 4750 -274 4806
rect -218 4750 -186 4806
rect -130 4750 -122 4806
rect -722 4725 -122 4750
rect -722 4669 -714 4725
rect -658 4669 -626 4725
rect -570 4669 -538 4725
rect -482 4669 -450 4725
rect -394 4669 -362 4725
rect -306 4669 -274 4725
rect -218 4669 -186 4725
rect -130 4669 -122 4725
rect -722 4644 -122 4669
rect -722 4588 -714 4644
rect -658 4588 -626 4644
rect -570 4588 -538 4644
rect -482 4588 -450 4644
rect -394 4588 -362 4644
rect -306 4588 -274 4644
rect -218 4588 -186 4644
rect -130 4588 -122 4644
rect -722 4563 -122 4588
rect -722 4507 -714 4563
rect -658 4507 -626 4563
rect -570 4507 -538 4563
rect -482 4507 -450 4563
rect -394 4507 -362 4563
rect -306 4507 -274 4563
rect -218 4507 -186 4563
rect -130 4507 -122 4563
rect -722 4482 -122 4507
rect -722 4426 -714 4482
rect -658 4426 -626 4482
rect -570 4426 -538 4482
rect -482 4426 -450 4482
rect -394 4426 -362 4482
rect -306 4426 -274 4482
rect -218 4426 -186 4482
rect -130 4426 -122 4482
rect -722 4401 -122 4426
rect -722 4345 -714 4401
rect -658 4345 -626 4401
rect -570 4345 -538 4401
rect -482 4345 -450 4401
rect -394 4345 -362 4401
rect -306 4345 -274 4401
rect -218 4345 -186 4401
rect -130 4345 -122 4401
rect -722 4320 -122 4345
rect -722 4264 -714 4320
rect -658 4264 -626 4320
rect -570 4264 -538 4320
rect -482 4264 -450 4320
rect -394 4264 -362 4320
rect -306 4264 -274 4320
rect -218 4264 -186 4320
rect -130 4264 -122 4320
rect -722 4239 -122 4264
rect -722 4183 -714 4239
rect -658 4183 -626 4239
rect -570 4183 -538 4239
rect -482 4183 -450 4239
rect -394 4183 -362 4239
rect -306 4183 -274 4239
rect -218 4183 -186 4239
rect -130 4183 -122 4239
rect -722 4158 -122 4183
rect -722 4102 -714 4158
rect -658 4102 -626 4158
rect -570 4102 -538 4158
rect -482 4102 -450 4158
rect -394 4102 -362 4158
rect -306 4102 -274 4158
rect -218 4102 -186 4158
rect -130 4102 -122 4158
rect -722 4077 -122 4102
rect -722 4021 -714 4077
rect -658 4021 -626 4077
rect -570 4021 -538 4077
rect -482 4021 -450 4077
rect -394 4021 -362 4077
rect -306 4021 -274 4077
rect -218 4021 -186 4077
rect -130 4021 -122 4077
rect -722 3996 -122 4021
rect -722 3940 -714 3996
rect -658 3940 -626 3996
rect -570 3940 -538 3996
rect -482 3940 -450 3996
rect -394 3940 -362 3996
rect -306 3940 -274 3996
rect -218 3940 -186 3996
rect -130 3940 -122 3996
rect -722 3915 -122 3940
rect -722 3859 -714 3915
rect -658 3859 -626 3915
rect -570 3859 -538 3915
rect -482 3859 -450 3915
rect -394 3859 -362 3915
rect -306 3859 -274 3915
rect -218 3859 -186 3915
rect -130 3859 -122 3915
rect -722 3834 -122 3859
rect -722 3778 -714 3834
rect -658 3778 -626 3834
rect -570 3778 -538 3834
rect -482 3778 -450 3834
rect -394 3778 -362 3834
rect -306 3778 -274 3834
rect -218 3778 -186 3834
rect -130 3778 -122 3834
rect -722 3753 -122 3778
rect -722 3697 -714 3753
rect -658 3697 -626 3753
rect -570 3697 -538 3753
rect -482 3697 -450 3753
rect -394 3697 -362 3753
rect -306 3697 -274 3753
rect -218 3697 -186 3753
rect -130 3697 -122 3753
rect -722 3672 -122 3697
rect -722 3616 -714 3672
rect -658 3616 -626 3672
rect -570 3616 -538 3672
rect -482 3616 -450 3672
rect -394 3616 -362 3672
rect -306 3616 -274 3672
rect -218 3616 -186 3672
rect -130 3616 -122 3672
rect -722 3591 -122 3616
rect -722 3535 -714 3591
rect -658 3535 -626 3591
rect -570 3535 -538 3591
rect -482 3535 -450 3591
rect -394 3535 -362 3591
rect -306 3535 -274 3591
rect -218 3535 -186 3591
rect -130 3535 -122 3591
rect -722 3510 -122 3535
rect 209 18381 217 18409
rect 281 18381 313 18445
rect 377 18381 409 18445
rect 473 18381 505 18445
rect 569 18381 601 18445
rect 665 18381 696 18445
rect 760 18409 766 18445
rect 760 18381 769 18409
rect 209 18357 769 18381
rect 209 18293 217 18357
rect 281 18293 313 18357
rect 377 18293 409 18357
rect 473 18293 505 18357
rect 569 18293 601 18357
rect 665 18293 696 18357
rect 760 18293 769 18357
rect 209 18269 769 18293
rect 209 18205 217 18269
rect 281 18205 313 18269
rect 377 18205 409 18269
rect 473 18205 505 18269
rect 569 18205 601 18269
rect 665 18205 696 18269
rect 760 18205 769 18269
rect 209 18181 769 18205
rect 209 18117 217 18181
rect 281 18117 313 18181
rect 377 18117 409 18181
rect 473 18117 505 18181
rect 569 18117 601 18181
rect 665 18117 696 18181
rect 760 18117 769 18181
rect 209 18093 769 18117
rect 209 18029 217 18093
rect 281 18029 313 18093
rect 377 18029 409 18093
rect 473 18029 505 18093
rect 569 18029 601 18093
rect 665 18029 696 18093
rect 760 18029 769 18093
rect 209 3526 769 18029
rect 1094 12927 1670 19040
rect 2898 20550 3474 20567
rect 2898 20494 2910 20550
rect 2966 20494 2992 20550
rect 3048 20494 3074 20550
rect 3130 20494 3156 20550
rect 3212 20494 3238 20550
rect 3294 20494 3320 20550
rect 3376 20494 3402 20550
rect 3458 20494 3474 20550
rect 2898 20470 3474 20494
rect 2898 20414 2910 20470
rect 2966 20414 2992 20470
rect 3048 20414 3074 20470
rect 3130 20414 3156 20470
rect 3212 20414 3238 20470
rect 3294 20414 3320 20470
rect 3376 20414 3402 20470
rect 3458 20414 3474 20470
rect 2898 20390 3474 20414
rect 2898 20334 2910 20390
rect 2966 20334 2992 20390
rect 3048 20334 3074 20390
rect 3130 20334 3156 20390
rect 3212 20334 3238 20390
rect 3294 20334 3320 20390
rect 3376 20334 3402 20390
rect 3458 20334 3474 20390
rect 2898 20310 3474 20334
rect 2898 20254 2910 20310
rect 2966 20254 2992 20310
rect 3048 20254 3074 20310
rect 3130 20254 3156 20310
rect 3212 20254 3238 20310
rect 3294 20254 3320 20310
rect 3376 20254 3402 20310
rect 3458 20254 3474 20310
rect 2898 20230 3474 20254
rect 2898 20174 2910 20230
rect 2966 20174 2992 20230
rect 3048 20174 3074 20230
rect 3130 20174 3156 20230
rect 3212 20174 3238 20230
rect 3294 20174 3320 20230
rect 3376 20174 3402 20230
rect 3458 20174 3474 20230
rect 2898 20149 3474 20174
rect 2898 20093 2910 20149
rect 2966 20093 2992 20149
rect 3048 20093 3074 20149
rect 3130 20093 3156 20149
rect 3212 20093 3238 20149
rect 3294 20093 3320 20149
rect 3376 20093 3402 20149
rect 3458 20093 3474 20149
rect 2898 20068 3474 20093
rect 2898 20012 2910 20068
rect 2966 20012 2992 20068
rect 3048 20012 3074 20068
rect 3130 20012 3156 20068
rect 3212 20012 3238 20068
rect 3294 20012 3320 20068
rect 3376 20012 3402 20068
rect 3458 20012 3474 20068
rect 2898 19987 3474 20012
rect 2898 19931 2910 19987
rect 2966 19931 2992 19987
rect 3048 19931 3074 19987
rect 3130 19931 3156 19987
rect 3212 19931 3238 19987
rect 3294 19931 3320 19987
rect 3376 19931 3402 19987
rect 3458 19931 3474 19987
rect 2898 19906 3474 19931
rect 2898 19850 2910 19906
rect 2966 19850 2992 19906
rect 3048 19850 3074 19906
rect 3130 19850 3156 19906
rect 3212 19850 3238 19906
rect 3294 19850 3320 19906
rect 3376 19850 3402 19906
rect 3458 19850 3474 19906
rect 2898 19825 3474 19850
rect 2898 19769 2910 19825
rect 2966 19769 2992 19825
rect 3048 19769 3074 19825
rect 3130 19769 3156 19825
rect 3212 19769 3238 19825
rect 3294 19769 3320 19825
rect 3376 19769 3402 19825
rect 3458 19769 3474 19825
rect 2898 19744 3474 19769
rect 2898 19688 2910 19744
rect 2966 19688 2992 19744
rect 3048 19688 3074 19744
rect 3130 19688 3156 19744
rect 3212 19688 3238 19744
rect 3294 19688 3320 19744
rect 3376 19688 3402 19744
rect 3458 19688 3474 19744
rect 2898 19663 3474 19688
rect 2898 19607 2910 19663
rect 2966 19607 2992 19663
rect 3048 19607 3074 19663
rect 3130 19607 3156 19663
rect 3212 19607 3238 19663
rect 3294 19607 3320 19663
rect 3376 19607 3402 19663
rect 3458 19607 3474 19663
rect 2898 19582 3474 19607
rect 2898 19526 2910 19582
rect 2966 19526 2992 19582
rect 3048 19526 3074 19582
rect 3130 19526 3156 19582
rect 3212 19526 3238 19582
rect 3294 19526 3320 19582
rect 3376 19526 3402 19582
rect 3458 19526 3474 19582
rect 2898 19501 3474 19526
rect 2898 19445 2910 19501
rect 2966 19445 2992 19501
rect 3048 19445 3074 19501
rect 3130 19445 3156 19501
rect 3212 19445 3238 19501
rect 3294 19445 3320 19501
rect 3376 19445 3402 19501
rect 3458 19445 3474 19501
rect 2898 19420 3474 19445
rect 2898 19364 2910 19420
rect 2966 19364 2992 19420
rect 3048 19364 3074 19420
rect 3130 19364 3156 19420
rect 3212 19364 3238 19420
rect 3294 19364 3320 19420
rect 3376 19364 3402 19420
rect 3458 19364 3474 19420
rect 2898 19339 3474 19364
rect 2898 19283 2910 19339
rect 2966 19283 2992 19339
rect 3048 19283 3074 19339
rect 3130 19283 3156 19339
rect 3212 19283 3238 19339
rect 3294 19283 3320 19339
rect 3376 19283 3402 19339
rect 3458 19283 3474 19339
rect 2898 19258 3474 19283
rect 2898 19202 2910 19258
rect 2966 19202 2992 19258
rect 3048 19202 3074 19258
rect 3130 19202 3156 19258
rect 3212 19202 3238 19258
rect 3294 19202 3320 19258
rect 3376 19202 3402 19258
rect 3458 19202 3474 19258
rect 2898 19177 3474 19202
rect 2898 19121 2910 19177
rect 2966 19121 2992 19177
rect 3048 19121 3074 19177
rect 3130 19121 3156 19177
rect 3212 19121 3238 19177
rect 3294 19121 3320 19177
rect 3376 19121 3402 19177
rect 3458 19121 3474 19177
rect 2898 19096 3474 19121
rect 2898 19040 2910 19096
rect 2966 19040 2992 19096
rect 3048 19040 3074 19096
rect 3130 19040 3156 19096
rect 3212 19040 3238 19096
rect 3294 19040 3320 19096
rect 3376 19040 3402 19096
rect 3458 19040 3474 19096
rect 2898 18904 3474 19040
tri 2898 18860 2942 18904 ne
rect 2942 18860 3474 18904
tri 2942 18790 3012 18860 ne
rect 3012 18824 3438 18860
tri 3438 18824 3474 18860 nw
rect 4696 20550 5272 20567
rect 4696 20494 4708 20550
rect 4764 20494 4790 20550
rect 4846 20494 4872 20550
rect 4928 20494 4954 20550
rect 5010 20494 5036 20550
rect 5092 20494 5118 20550
rect 5174 20494 5200 20550
rect 5256 20494 5272 20550
rect 4696 20470 5272 20494
rect 4696 20414 4708 20470
rect 4764 20414 4790 20470
rect 4846 20414 4872 20470
rect 4928 20414 4954 20470
rect 5010 20414 5036 20470
rect 5092 20414 5118 20470
rect 5174 20414 5200 20470
rect 5256 20414 5272 20470
rect 4696 20390 5272 20414
rect 4696 20334 4708 20390
rect 4764 20334 4790 20390
rect 4846 20334 4872 20390
rect 4928 20334 4954 20390
rect 5010 20334 5036 20390
rect 5092 20334 5118 20390
rect 5174 20334 5200 20390
rect 5256 20334 5272 20390
rect 4696 20310 5272 20334
rect 4696 20254 4708 20310
rect 4764 20254 4790 20310
rect 4846 20254 4872 20310
rect 4928 20254 4954 20310
rect 5010 20254 5036 20310
rect 5092 20254 5118 20310
rect 5174 20254 5200 20310
rect 5256 20254 5272 20310
rect 4696 20230 5272 20254
rect 4696 20174 4708 20230
rect 4764 20174 4790 20230
rect 4846 20174 4872 20230
rect 4928 20174 4954 20230
rect 5010 20174 5036 20230
rect 5092 20174 5118 20230
rect 5174 20174 5200 20230
rect 5256 20174 5272 20230
rect 4696 20149 5272 20174
rect 4696 20093 4708 20149
rect 4764 20093 4790 20149
rect 4846 20093 4872 20149
rect 4928 20093 4954 20149
rect 5010 20093 5036 20149
rect 5092 20093 5118 20149
rect 5174 20093 5200 20149
rect 5256 20093 5272 20149
rect 4696 20068 5272 20093
rect 4696 20012 4708 20068
rect 4764 20012 4790 20068
rect 4846 20012 4872 20068
rect 4928 20012 4954 20068
rect 5010 20012 5036 20068
rect 5092 20012 5118 20068
rect 5174 20012 5200 20068
rect 5256 20012 5272 20068
rect 4696 19987 5272 20012
rect 4696 19931 4708 19987
rect 4764 19931 4790 19987
rect 4846 19931 4872 19987
rect 4928 19931 4954 19987
rect 5010 19931 5036 19987
rect 5092 19931 5118 19987
rect 5174 19931 5200 19987
rect 5256 19931 5272 19987
rect 4696 19906 5272 19931
rect 4696 19850 4708 19906
rect 4764 19850 4790 19906
rect 4846 19850 4872 19906
rect 4928 19850 4954 19906
rect 5010 19850 5036 19906
rect 5092 19850 5118 19906
rect 5174 19850 5200 19906
rect 5256 19850 5272 19906
rect 4696 19825 5272 19850
rect 4696 19769 4708 19825
rect 4764 19769 4790 19825
rect 4846 19769 4872 19825
rect 4928 19769 4954 19825
rect 5010 19769 5036 19825
rect 5092 19769 5118 19825
rect 5174 19769 5200 19825
rect 5256 19769 5272 19825
rect 4696 19744 5272 19769
rect 4696 19688 4708 19744
rect 4764 19688 4790 19744
rect 4846 19688 4872 19744
rect 4928 19688 4954 19744
rect 5010 19688 5036 19744
rect 5092 19688 5118 19744
rect 5174 19688 5200 19744
rect 5256 19688 5272 19744
rect 4696 19663 5272 19688
rect 4696 19607 4708 19663
rect 4764 19607 4790 19663
rect 4846 19607 4872 19663
rect 4928 19607 4954 19663
rect 5010 19607 5036 19663
rect 5092 19607 5118 19663
rect 5174 19607 5200 19663
rect 5256 19607 5272 19663
rect 4696 19582 5272 19607
rect 4696 19526 4708 19582
rect 4764 19526 4790 19582
rect 4846 19526 4872 19582
rect 4928 19526 4954 19582
rect 5010 19526 5036 19582
rect 5092 19526 5118 19582
rect 5174 19526 5200 19582
rect 5256 19526 5272 19582
rect 4696 19501 5272 19526
rect 4696 19445 4708 19501
rect 4764 19445 4790 19501
rect 4846 19445 4872 19501
rect 4928 19445 4954 19501
rect 5010 19445 5036 19501
rect 5092 19445 5118 19501
rect 5174 19445 5200 19501
rect 5256 19445 5272 19501
rect 4696 19420 5272 19445
rect 4696 19364 4708 19420
rect 4764 19364 4790 19420
rect 4846 19364 4872 19420
rect 4928 19364 4954 19420
rect 5010 19364 5036 19420
rect 5092 19364 5118 19420
rect 5174 19364 5200 19420
rect 5256 19364 5272 19420
rect 4696 19339 5272 19364
rect 4696 19283 4708 19339
rect 4764 19283 4790 19339
rect 4846 19283 4872 19339
rect 4928 19283 4954 19339
rect 5010 19283 5036 19339
rect 5092 19283 5118 19339
rect 5174 19283 5200 19339
rect 5256 19283 5272 19339
rect 4696 19258 5272 19283
rect 4696 19202 4708 19258
rect 4764 19202 4790 19258
rect 4846 19202 4872 19258
rect 4928 19202 4954 19258
rect 5010 19202 5036 19258
rect 5092 19202 5118 19258
rect 5174 19202 5200 19258
rect 5256 19202 5272 19258
rect 4696 19177 5272 19202
rect 4696 19121 4708 19177
rect 4764 19121 4790 19177
rect 4846 19121 4872 19177
rect 4928 19121 4954 19177
rect 5010 19121 5036 19177
rect 5092 19121 5118 19177
rect 5174 19121 5200 19177
rect 5256 19121 5272 19177
rect 4696 19096 5272 19121
rect 4696 19040 4708 19096
rect 4764 19040 4790 19096
rect 4846 19040 4872 19096
rect 4928 19040 4954 19096
rect 5010 19040 5036 19096
rect 5092 19040 5118 19096
rect 5174 19040 5200 19096
rect 5256 19040 5272 19096
rect 4696 18942 5272 19040
rect 6370 20550 6759 20567
rect 6370 20174 6378 20550
rect 6754 20174 6759 20550
rect 6370 20149 6759 20174
rect 6370 20093 6378 20149
rect 6434 20093 6458 20149
rect 6514 20093 6538 20149
rect 6594 20093 6618 20149
rect 6674 20093 6698 20149
rect 6754 20093 6759 20149
rect 6370 20068 6759 20093
rect 6370 20012 6378 20068
rect 6434 20012 6458 20068
rect 6514 20012 6538 20068
rect 6594 20012 6618 20068
rect 6674 20012 6698 20068
rect 6754 20012 6759 20068
rect 6370 19987 6759 20012
rect 6370 19931 6378 19987
rect 6434 19931 6458 19987
rect 6514 19931 6538 19987
rect 6594 19931 6618 19987
rect 6674 19931 6698 19987
rect 6754 19931 6759 19987
rect 6370 19906 6759 19931
rect 6370 19850 6378 19906
rect 6434 19850 6458 19906
rect 6514 19850 6538 19906
rect 6594 19850 6618 19906
rect 6674 19850 6698 19906
rect 6754 19850 6759 19906
rect 6370 19825 6759 19850
rect 6370 19769 6378 19825
rect 6434 19769 6458 19825
rect 6514 19769 6538 19825
rect 6594 19769 6618 19825
rect 6674 19769 6698 19825
rect 6754 19769 6759 19825
rect 6370 19744 6759 19769
rect 6370 19688 6378 19744
rect 6434 19688 6458 19744
rect 6514 19688 6538 19744
rect 6594 19688 6618 19744
rect 6674 19688 6698 19744
rect 6754 19688 6759 19744
rect 6370 19663 6759 19688
rect 6370 19607 6378 19663
rect 6434 19607 6458 19663
rect 6514 19607 6538 19663
rect 6594 19607 6618 19663
rect 6674 19607 6698 19663
rect 6754 19607 6759 19663
rect 6370 19582 6759 19607
rect 6370 19526 6378 19582
rect 6434 19526 6458 19582
rect 6514 19526 6538 19582
rect 6594 19526 6618 19582
rect 6674 19526 6698 19582
rect 6754 19526 6759 19582
rect 6370 19501 6759 19526
rect 6370 19445 6378 19501
rect 6434 19445 6458 19501
rect 6514 19445 6538 19501
rect 6594 19445 6618 19501
rect 6674 19445 6698 19501
rect 6754 19445 6759 19501
rect 6370 19420 6759 19445
rect 6370 19364 6378 19420
rect 6434 19364 6458 19420
rect 6514 19364 6538 19420
rect 6594 19364 6618 19420
rect 6674 19364 6698 19420
rect 6754 19364 6759 19420
rect 6370 19339 6759 19364
rect 6370 19283 6378 19339
rect 6434 19283 6458 19339
rect 6514 19283 6538 19339
rect 6594 19283 6618 19339
rect 6674 19283 6698 19339
rect 6754 19283 6759 19339
rect 6370 19258 6759 19283
rect 6370 19202 6378 19258
rect 6434 19202 6458 19258
rect 6514 19202 6538 19258
rect 6594 19202 6618 19258
rect 6674 19202 6698 19258
rect 6754 19202 6759 19258
rect 6370 19177 6759 19202
rect 6370 19121 6378 19177
rect 6434 19121 6458 19177
rect 6514 19121 6538 19177
rect 6594 19121 6618 19177
rect 6674 19121 6698 19177
rect 6754 19121 6759 19177
rect 6370 19096 6759 19121
rect 6370 19040 6378 19096
rect 6434 19040 6458 19096
rect 6514 19040 6538 19096
rect 6594 19040 6618 19096
rect 6674 19040 6698 19096
rect 6754 19040 6759 19096
rect 6370 19019 6759 19040
rect 4696 18887 5051 18942
tri 4696 18824 4759 18887 ne
rect 3012 18790 3404 18824
tri 3404 18790 3438 18824 nw
tri 3012 18785 3017 18790 ne
rect 2018 18409 2024 18445
rect 1094 12871 1115 12927
rect 1171 12871 1211 12927
rect 1267 12871 1307 12927
rect 1363 12871 1402 12927
rect 1458 12871 1497 12927
rect 1553 12871 1592 12927
rect 1648 12871 1670 12927
rect 1094 12843 1670 12871
rect 1094 12787 1115 12843
rect 1171 12787 1211 12843
rect 1267 12787 1307 12843
rect 1363 12787 1402 12843
rect 1458 12787 1497 12843
rect 1553 12787 1592 12843
rect 1648 12787 1670 12843
rect 1094 12759 1670 12787
rect 1094 12703 1115 12759
rect 1171 12703 1211 12759
rect 1267 12703 1307 12759
rect 1363 12703 1402 12759
rect 1458 12703 1497 12759
rect 1553 12703 1592 12759
rect 1648 12703 1670 12759
rect 1094 12675 1670 12703
rect 1094 12619 1115 12675
rect 1171 12619 1211 12675
rect 1267 12619 1307 12675
rect 1363 12619 1402 12675
rect 1458 12619 1497 12675
rect 1553 12619 1592 12675
rect 1648 12619 1670 12675
rect 1094 12591 1670 12619
rect 1094 12535 1115 12591
rect 1171 12535 1211 12591
rect 1267 12535 1307 12591
rect 1363 12535 1402 12591
rect 1458 12535 1497 12591
rect 1553 12535 1592 12591
rect 1648 12535 1670 12591
rect 1094 12507 1670 12535
rect 1094 12451 1115 12507
rect 1171 12451 1211 12507
rect 1267 12451 1307 12507
rect 1363 12451 1402 12507
rect 1458 12451 1497 12507
rect 1553 12451 1592 12507
rect 1648 12451 1670 12507
rect 1094 12440 1670 12451
rect 2013 18381 2024 18409
rect 2088 18381 2120 18445
rect 2184 18381 2216 18445
rect 2280 18381 2312 18445
rect 2376 18381 2408 18445
rect 2472 18381 2503 18445
rect 2567 18381 2573 18445
rect 2013 18357 2573 18381
rect 2013 18293 2024 18357
rect 2088 18293 2120 18357
rect 2184 18293 2216 18357
rect 2280 18293 2312 18357
rect 2376 18293 2408 18357
rect 2472 18293 2503 18357
rect 2567 18293 2573 18357
tri 2950 18347 3017 18414 se
rect 3017 18409 3404 18790
tri 4727 18445 4759 18477 se
rect 4759 18445 5051 18887
tri 5051 18793 5200 18942 nw
rect 6370 18885 6706 19019
tri 6706 18966 6759 19019 nw
rect 8061 20556 8334 20566
rect 8061 20500 8067 20556
rect 8123 20500 8169 20556
rect 8225 20500 8271 20556
rect 8327 20500 8334 20556
rect 8061 20475 8334 20500
rect 8061 20419 8067 20475
rect 8123 20419 8169 20475
rect 8225 20419 8271 20475
rect 8327 20419 8334 20475
rect 8061 20394 8334 20419
rect 8061 20338 8067 20394
rect 8123 20338 8169 20394
rect 8225 20338 8271 20394
rect 8327 20338 8334 20394
rect 8061 20313 8334 20338
rect 8061 20257 8067 20313
rect 8123 20257 8169 20313
rect 8225 20257 8271 20313
rect 8327 20257 8334 20313
rect 8061 20232 8334 20257
rect 8061 20176 8067 20232
rect 8123 20176 8169 20232
rect 8225 20176 8271 20232
rect 8327 20176 8334 20232
rect 8061 20151 8334 20176
rect 8061 20095 8067 20151
rect 8123 20095 8169 20151
rect 8225 20095 8271 20151
rect 8327 20095 8334 20151
rect 8061 20070 8334 20095
rect 8061 20014 8067 20070
rect 8123 20014 8169 20070
rect 8225 20014 8271 20070
rect 8327 20014 8334 20070
rect 8061 19989 8334 20014
rect 8061 19933 8067 19989
rect 8123 19933 8169 19989
rect 8225 19933 8271 19989
rect 8327 19933 8334 19989
rect 8061 19908 8334 19933
rect 8061 19852 8067 19908
rect 8123 19852 8169 19908
rect 8225 19852 8271 19908
rect 8327 19852 8334 19908
rect 8061 19827 8334 19852
rect 8061 19771 8067 19827
rect 8123 19771 8169 19827
rect 8225 19771 8271 19827
rect 8327 19771 8334 19827
rect 8061 19745 8334 19771
rect 8061 19689 8067 19745
rect 8123 19689 8169 19745
rect 8225 19689 8271 19745
rect 8327 19689 8334 19745
rect 8061 19663 8334 19689
rect 8061 19607 8067 19663
rect 8123 19607 8169 19663
rect 8225 19607 8271 19663
rect 8327 19607 8334 19663
rect 8061 19581 8334 19607
rect 8061 19525 8067 19581
rect 8123 19525 8169 19581
rect 8225 19525 8271 19581
rect 8327 19525 8334 19581
rect 8061 19499 8334 19525
rect 8061 19443 8067 19499
rect 8123 19443 8169 19499
rect 8225 19443 8271 19499
rect 8327 19443 8334 19499
rect 8061 19417 8334 19443
rect 8061 19361 8067 19417
rect 8123 19361 8169 19417
rect 8225 19361 8271 19417
rect 8327 19361 8334 19417
rect 8061 19335 8334 19361
rect 8061 19279 8067 19335
rect 8123 19279 8169 19335
rect 8225 19279 8271 19335
rect 8327 19279 8334 19335
rect 8061 19253 8334 19279
rect 8061 19197 8067 19253
rect 8123 19197 8169 19253
rect 8225 19197 8271 19253
rect 8327 19197 8334 19253
rect 8061 19171 8334 19197
rect 8061 19115 8067 19171
rect 8123 19115 8169 19171
rect 8225 19115 8271 19171
rect 8327 19115 8334 19171
rect 8061 19089 8334 19115
rect 8061 19033 8067 19089
rect 8123 19033 8169 19089
rect 8225 19033 8271 19089
rect 8327 19033 8334 19089
tri 6370 18847 6408 18885 ne
tri 3404 18409 3412 18417 sw
rect 3813 18409 3819 18445
rect 3017 18347 3412 18409
tri 3412 18347 3474 18409 sw
rect 2013 18269 2573 18293
rect 2013 18205 2024 18269
rect 2088 18205 2120 18269
rect 2184 18205 2216 18269
rect 2280 18205 2312 18269
rect 2376 18205 2408 18269
rect 2472 18205 2503 18269
rect 2567 18205 2573 18269
rect 2013 18181 2573 18205
rect 2013 18117 2024 18181
rect 2088 18117 2120 18181
rect 2184 18117 2216 18181
rect 2280 18117 2312 18181
rect 2376 18117 2408 18181
rect 2472 18117 2503 18181
rect 2567 18117 2573 18181
rect 2013 18093 2573 18117
rect 2013 18029 2024 18093
rect 2088 18029 2120 18093
rect 2184 18029 2216 18093
rect 2280 18029 2312 18093
rect 2376 18029 2408 18093
rect 2472 18029 2503 18093
rect 2567 18029 2573 18093
rect -722 3454 -714 3510
rect -658 3454 -626 3510
rect -570 3454 -538 3510
rect -482 3454 -450 3510
rect -394 3454 -362 3510
rect -306 3454 -274 3510
rect -218 3454 -186 3510
rect -130 3454 -122 3510
rect -722 3429 -122 3454
rect -722 3373 -714 3429
rect -658 3373 -626 3429
rect -570 3373 -538 3429
rect -482 3373 -450 3429
rect -394 3373 -362 3429
rect -306 3373 -274 3429
rect -218 3373 -186 3429
rect -130 3373 -122 3429
rect -722 3348 -122 3373
rect -722 3292 -714 3348
rect -658 3292 -626 3348
rect -570 3292 -538 3348
rect -482 3292 -450 3348
rect -394 3292 -362 3348
rect -306 3292 -274 3348
rect -218 3292 -186 3348
rect -130 3292 -122 3348
rect -722 3267 -122 3292
rect -722 3211 -714 3267
rect -658 3211 -626 3267
rect -570 3211 -538 3267
rect -482 3211 -450 3267
rect -394 3211 -362 3267
rect -306 3211 -274 3267
rect -218 3211 -186 3267
rect -130 3211 -122 3267
rect -722 3194 -122 3211
rect 1094 3173 1670 12080
rect 2013 3526 2573 18029
tri 2898 18295 2950 18347 se
rect 2950 18295 3474 18347
rect 2898 13046 3474 18295
rect 2898 12990 2906 13046
rect 2962 12990 2990 13046
rect 3046 12990 3074 13046
rect 3130 12990 3158 13046
rect 3214 12990 3242 13046
rect 3298 12990 3326 13046
rect 3382 12990 3410 13046
rect 3466 12990 3474 13046
rect 2898 12957 3474 12990
rect 2898 12901 2906 12957
rect 2962 12901 2990 12957
rect 3046 12901 3074 12957
rect 3130 12901 3158 12957
rect 3214 12901 3242 12957
rect 3298 12901 3326 12957
rect 3382 12901 3410 12957
rect 3466 12901 3474 12957
rect 2898 12868 3474 12901
rect 2898 12812 2906 12868
rect 2962 12812 2990 12868
rect 3046 12812 3074 12868
rect 3130 12812 3158 12868
rect 3214 12812 3242 12868
rect 3298 12812 3326 12868
rect 3382 12812 3410 12868
rect 3466 12812 3474 12868
rect 2898 12779 3474 12812
rect 2898 12723 2906 12779
rect 2962 12723 2990 12779
rect 3046 12723 3074 12779
rect 3130 12723 3158 12779
rect 3214 12723 3242 12779
rect 3298 12723 3326 12779
rect 3382 12723 3410 12779
rect 3466 12723 3474 12779
rect 2898 12690 3474 12723
rect 2898 12634 2906 12690
rect 2962 12634 2990 12690
rect 3046 12634 3074 12690
rect 3130 12634 3158 12690
rect 3214 12634 3242 12690
rect 3298 12634 3326 12690
rect 3382 12634 3410 12690
rect 3466 12634 3474 12690
rect 2898 12601 3474 12634
rect 2898 12545 2906 12601
rect 2962 12545 2990 12601
rect 3046 12545 3074 12601
rect 3130 12545 3158 12601
rect 3214 12545 3242 12601
rect 3298 12545 3326 12601
rect 3382 12545 3410 12601
rect 3466 12545 3474 12601
rect 2898 12511 3474 12545
rect 2898 12455 2906 12511
rect 2962 12455 2990 12511
rect 3046 12455 3074 12511
rect 3130 12455 3158 12511
rect 3214 12455 3242 12511
rect 3298 12455 3326 12511
rect 3382 12455 3410 12511
rect 3466 12455 3474 12511
rect 2898 12444 3474 12455
rect 3811 18381 3819 18409
rect 3883 18381 3915 18445
rect 3979 18381 4011 18445
rect 4075 18381 4107 18445
rect 4171 18381 4203 18445
rect 4267 18381 4298 18445
rect 4362 18409 4368 18445
tri 4699 18417 4727 18445 se
rect 4727 18417 5051 18445
tri 4696 18414 4699 18417 se
rect 4699 18414 5051 18417
rect 4696 18409 5051 18414
tri 5051 18409 5059 18417 sw
rect 5623 18409 5629 18445
rect 4362 18381 4371 18409
rect 3811 18357 4371 18381
rect 3811 18293 3819 18357
rect 3883 18293 3915 18357
rect 3979 18293 4011 18357
rect 4075 18293 4107 18357
rect 4171 18293 4203 18357
rect 4267 18293 4298 18357
rect 4362 18293 4371 18357
rect 3811 18269 4371 18293
rect 3811 18205 3819 18269
rect 3883 18205 3915 18269
rect 3979 18205 4011 18269
rect 4075 18205 4107 18269
rect 4171 18205 4203 18269
rect 4267 18205 4298 18269
rect 4362 18205 4371 18269
rect 3811 18181 4371 18205
rect 3811 18117 3819 18181
rect 3883 18117 3915 18181
rect 3979 18117 4011 18181
rect 4075 18117 4107 18181
rect 4171 18117 4203 18181
rect 4267 18117 4298 18181
rect 4362 18117 4371 18181
rect 3811 18093 4371 18117
rect 3811 18029 3819 18093
rect 3883 18029 3915 18093
rect 3979 18029 4011 18093
rect 4075 18029 4107 18093
rect 4171 18029 4203 18093
rect 4267 18029 4298 18093
rect 4362 18029 4371 18093
tri 1670 3173 1673 3176 sw
rect 2898 3173 3474 12080
rect 3811 3526 4371 18029
rect 4696 18255 5059 18409
tri 5059 18255 5213 18409 sw
rect 5618 18381 5629 18409
rect 5693 18381 5725 18445
rect 5789 18381 5821 18445
rect 5885 18381 5917 18445
rect 5981 18381 6013 18445
rect 6077 18381 6108 18445
rect 6172 18381 6178 18445
rect 5618 18357 6178 18381
rect 5618 18293 5629 18357
rect 5693 18293 5725 18357
rect 5789 18293 5821 18357
rect 5885 18293 5917 18357
rect 5981 18293 6013 18357
rect 6077 18293 6108 18357
rect 6172 18293 6178 18357
rect 5618 18269 6178 18293
rect 4696 13046 5272 18255
rect 4696 12990 4704 13046
rect 4760 12990 4788 13046
rect 4844 12990 4872 13046
rect 4928 12990 4956 13046
rect 5012 12990 5040 13046
rect 5096 12990 5124 13046
rect 5180 12990 5208 13046
rect 5264 12990 5272 13046
rect 4696 12957 5272 12990
rect 4696 12901 4704 12957
rect 4760 12901 4788 12957
rect 4844 12901 4872 12957
rect 4928 12901 4956 12957
rect 5012 12901 5040 12957
rect 5096 12901 5124 12957
rect 5180 12901 5208 12957
rect 5264 12901 5272 12957
rect 4696 12868 5272 12901
rect 4696 12812 4704 12868
rect 4760 12812 4788 12868
rect 4844 12812 4872 12868
rect 4928 12812 4956 12868
rect 5012 12812 5040 12868
rect 5096 12812 5124 12868
rect 5180 12812 5208 12868
rect 5264 12812 5272 12868
rect 4696 12779 5272 12812
rect 4696 12723 4704 12779
rect 4760 12723 4788 12779
rect 4844 12723 4872 12779
rect 4928 12723 4956 12779
rect 5012 12723 5040 12779
rect 5096 12723 5124 12779
rect 5180 12723 5208 12779
rect 5264 12723 5272 12779
rect 4696 12690 5272 12723
rect 4696 12634 4704 12690
rect 4760 12634 4788 12690
rect 4844 12634 4872 12690
rect 4928 12634 4956 12690
rect 5012 12634 5040 12690
rect 5096 12634 5124 12690
rect 5180 12634 5208 12690
rect 5264 12634 5272 12690
rect 4696 12601 5272 12634
rect 4696 12545 4704 12601
rect 4760 12545 4788 12601
rect 4844 12545 4872 12601
rect 4928 12545 4956 12601
rect 5012 12545 5040 12601
rect 5096 12545 5124 12601
rect 5180 12545 5208 12601
rect 5264 12545 5272 12601
rect 4696 12511 5272 12545
rect 4696 12455 4704 12511
rect 4760 12455 4788 12511
rect 4844 12455 4872 12511
rect 4928 12455 4956 12511
rect 5012 12455 5040 12511
rect 5096 12455 5124 12511
rect 5180 12455 5208 12511
rect 5264 12455 5272 12511
rect 4696 12444 5272 12455
rect 5618 18205 5629 18269
rect 5693 18205 5725 18269
rect 5789 18205 5821 18269
rect 5885 18205 5917 18269
rect 5981 18205 6013 18269
rect 6077 18205 6108 18269
rect 6172 18205 6178 18269
rect 5618 18181 6178 18205
rect 5618 18117 5629 18181
rect 5693 18117 5725 18181
rect 5789 18117 5821 18181
rect 5885 18117 5917 18181
rect 5981 18117 6013 18181
rect 6077 18117 6108 18181
rect 6172 18117 6178 18181
rect 5618 18093 6178 18117
rect 5618 18029 5629 18093
rect 5693 18029 5725 18093
rect 5789 18029 5821 18093
rect 5885 18029 5917 18093
rect 5981 18029 6013 18093
rect 6077 18029 6108 18093
rect 6172 18029 6178 18093
rect 6408 18126 6706 18885
rect 7421 18409 7427 18445
rect 7419 18381 7427 18409
rect 7491 18381 7523 18445
rect 7587 18381 7619 18445
rect 7683 18381 7715 18445
rect 7779 18381 7811 18445
rect 7875 18381 7906 18445
rect 7970 18409 7976 18445
rect 7970 18381 7979 18409
rect 7419 18357 7979 18381
tri 6408 18031 6503 18126 ne
tri 3474 3173 3477 3176 sw
rect 4699 3173 5275 12080
rect 5618 3526 6178 18029
rect 6503 17947 6706 18126
tri 6706 17947 7079 18320 sw
rect 6503 13046 7079 17947
rect 6503 12990 6511 13046
rect 6567 12990 6595 13046
rect 6651 12990 6679 13046
rect 6735 12990 6763 13046
rect 6819 12990 6847 13046
rect 6903 12990 6931 13046
rect 6987 12990 7015 13046
rect 7071 12990 7079 13046
rect 6503 12957 7079 12990
rect 6503 12901 6511 12957
rect 6567 12901 6595 12957
rect 6651 12901 6679 12957
rect 6735 12901 6763 12957
rect 6819 12901 6847 12957
rect 6903 12901 6931 12957
rect 6987 12901 7015 12957
rect 7071 12901 7079 12957
rect 6503 12868 7079 12901
rect 6503 12812 6511 12868
rect 6567 12812 6595 12868
rect 6651 12812 6679 12868
rect 6735 12812 6763 12868
rect 6819 12812 6847 12868
rect 6903 12812 6931 12868
rect 6987 12812 7015 12868
rect 7071 12812 7079 12868
rect 6503 12779 7079 12812
rect 6503 12723 6511 12779
rect 6567 12723 6595 12779
rect 6651 12723 6679 12779
rect 6735 12723 6763 12779
rect 6819 12723 6847 12779
rect 6903 12723 6931 12779
rect 6987 12723 7015 12779
rect 7071 12723 7079 12779
rect 6503 12690 7079 12723
rect 6503 12634 6511 12690
rect 6567 12634 6595 12690
rect 6651 12634 6679 12690
rect 6735 12634 6763 12690
rect 6819 12634 6847 12690
rect 6903 12634 6931 12690
rect 6987 12634 7015 12690
rect 7071 12634 7079 12690
rect 6503 12601 7079 12634
rect 6503 12545 6511 12601
rect 6567 12545 6595 12601
rect 6651 12545 6679 12601
rect 6735 12545 6763 12601
rect 6819 12545 6847 12601
rect 6903 12545 6931 12601
rect 6987 12545 7015 12601
rect 7071 12545 7079 12601
rect 6503 12511 7079 12545
rect 6503 12455 6511 12511
rect 6567 12455 6595 12511
rect 6651 12455 6679 12511
rect 6735 12455 6763 12511
rect 6819 12455 6847 12511
rect 6903 12455 6931 12511
rect 6987 12455 7015 12511
rect 7071 12455 7079 12511
rect 6503 12444 7079 12455
rect 7419 18293 7427 18357
rect 7491 18293 7523 18357
rect 7587 18293 7619 18357
rect 7683 18293 7715 18357
rect 7779 18293 7811 18357
rect 7875 18293 7906 18357
rect 7970 18293 7979 18357
rect 7419 18269 7979 18293
rect 7419 18205 7427 18269
rect 7491 18205 7523 18269
rect 7587 18205 7619 18269
rect 7683 18205 7715 18269
rect 7779 18205 7811 18269
rect 7875 18205 7906 18269
rect 7970 18205 7979 18269
rect 8061 18391 8334 19033
rect 8885 20556 9151 20566
rect 8885 20500 8894 20556
rect 8950 20500 8990 20556
rect 9046 20500 9086 20556
rect 9142 20500 9151 20556
rect 8885 20475 9151 20500
rect 8885 20419 8894 20475
rect 8950 20419 8990 20475
rect 9046 20419 9086 20475
rect 9142 20419 9151 20475
rect 8885 20394 9151 20419
rect 8885 20338 8894 20394
rect 8950 20338 8990 20394
rect 9046 20338 9086 20394
rect 9142 20338 9151 20394
rect 8885 20313 9151 20338
rect 8885 20257 8894 20313
rect 8950 20257 8990 20313
rect 9046 20257 9086 20313
rect 9142 20257 9151 20313
rect 8885 20232 9151 20257
rect 8885 20176 8894 20232
rect 8950 20176 8990 20232
rect 9046 20176 9086 20232
rect 9142 20176 9151 20232
rect 8885 20151 9151 20176
rect 8885 20095 8894 20151
rect 8950 20095 8990 20151
rect 9046 20095 9086 20151
rect 9142 20095 9151 20151
rect 8885 20070 9151 20095
rect 8885 20014 8894 20070
rect 8950 20014 8990 20070
rect 9046 20014 9086 20070
rect 9142 20014 9151 20070
rect 8885 19989 9151 20014
rect 8885 19933 8894 19989
rect 8950 19933 8990 19989
rect 9046 19933 9086 19989
rect 9142 19933 9151 19989
rect 8885 19908 9151 19933
rect 8885 19852 8894 19908
rect 8950 19852 8990 19908
rect 9046 19852 9086 19908
rect 9142 19852 9151 19908
rect 8885 19827 9151 19852
rect 8885 19771 8894 19827
rect 8950 19771 8990 19827
rect 9046 19771 9086 19827
rect 9142 19771 9151 19827
rect 8885 19745 9151 19771
rect 8885 19689 8894 19745
rect 8950 19689 8990 19745
rect 9046 19689 9086 19745
rect 9142 19689 9151 19745
rect 8885 19663 9151 19689
rect 8885 19607 8894 19663
rect 8950 19607 8990 19663
rect 9046 19607 9086 19663
rect 9142 19607 9151 19663
rect 8885 19581 9151 19607
rect 8885 19525 8894 19581
rect 8950 19525 8990 19581
rect 9046 19525 9086 19581
rect 9142 19525 9151 19581
rect 8885 19499 9151 19525
rect 8885 19443 8894 19499
rect 8950 19443 8990 19499
rect 9046 19443 9086 19499
rect 9142 19443 9151 19499
rect 8885 19417 9151 19443
rect 8885 19361 8894 19417
rect 8950 19361 8990 19417
rect 9046 19361 9086 19417
rect 9142 19361 9151 19417
rect 8885 19335 9151 19361
rect 8885 19279 8894 19335
rect 8950 19279 8990 19335
rect 9046 19279 9086 19335
rect 9142 19279 9151 19335
rect 8885 19253 9151 19279
rect 8885 19197 8894 19253
rect 8950 19197 8990 19253
rect 9046 19197 9086 19253
rect 9142 19197 9151 19253
rect 8885 19171 9151 19197
rect 8885 19115 8894 19171
rect 8950 19115 8990 19171
rect 9046 19115 9086 19171
rect 9142 19115 9151 19171
rect 8885 19089 9151 19115
rect 8885 19033 8894 19089
rect 8950 19033 8990 19089
rect 9046 19033 9086 19089
rect 9142 19033 9151 19089
tri 8334 18391 8350 18407 sw
rect 8061 18344 8350 18391
tri 8061 18243 8162 18344 ne
rect 8162 18243 8350 18344
tri 8350 18243 8498 18391 sw
tri 8737 18243 8885 18391 se
rect 8885 18271 9151 19033
rect 10114 20550 10690 20567
rect 10114 20494 10126 20550
rect 10182 20494 10208 20550
rect 10264 20494 10290 20550
rect 10346 20494 10372 20550
rect 10428 20494 10454 20550
rect 10510 20494 10536 20550
rect 10592 20494 10618 20550
rect 10674 20494 10690 20550
rect 10114 20467 10690 20494
rect 10114 20411 10126 20467
rect 10182 20411 10208 20467
rect 10264 20411 10290 20467
rect 10346 20411 10372 20467
rect 10428 20411 10454 20467
rect 10510 20411 10536 20467
rect 10592 20411 10618 20467
rect 10674 20411 10690 20467
rect 10114 20384 10690 20411
rect 10114 20328 10126 20384
rect 10182 20328 10208 20384
rect 10264 20328 10290 20384
rect 10346 20328 10372 20384
rect 10428 20328 10454 20384
rect 10510 20328 10536 20384
rect 10592 20328 10618 20384
rect 10674 20328 10690 20384
rect 10114 20301 10690 20328
rect 10114 20245 10126 20301
rect 10182 20245 10208 20301
rect 10264 20245 10290 20301
rect 10346 20245 10372 20301
rect 10428 20245 10454 20301
rect 10510 20245 10536 20301
rect 10592 20245 10618 20301
rect 10674 20245 10690 20301
rect 10114 20217 10690 20245
rect 10114 20161 10126 20217
rect 10182 20161 10208 20217
rect 10264 20161 10290 20217
rect 10346 20161 10372 20217
rect 10428 20161 10454 20217
rect 10510 20161 10536 20217
rect 10592 20161 10618 20217
rect 10674 20161 10690 20217
rect 10114 20133 10690 20161
rect 10114 20077 10126 20133
rect 10182 20077 10208 20133
rect 10264 20077 10290 20133
rect 10346 20077 10372 20133
rect 10428 20077 10454 20133
rect 10510 20077 10536 20133
rect 10592 20077 10618 20133
rect 10674 20077 10690 20133
rect 10114 20049 10690 20077
rect 10114 19993 10126 20049
rect 10182 19993 10208 20049
rect 10264 19993 10290 20049
rect 10346 19993 10372 20049
rect 10428 19993 10454 20049
rect 10510 19993 10536 20049
rect 10592 19993 10618 20049
rect 10674 19993 10690 20049
rect 10114 19965 10690 19993
rect 10114 19909 10126 19965
rect 10182 19909 10208 19965
rect 10264 19909 10290 19965
rect 10346 19909 10372 19965
rect 10428 19909 10454 19965
rect 10510 19909 10536 19965
rect 10592 19909 10618 19965
rect 10674 19909 10690 19965
rect 10114 19881 10690 19909
rect 10114 19825 10126 19881
rect 10182 19825 10208 19881
rect 10264 19825 10290 19881
rect 10346 19825 10372 19881
rect 10428 19825 10454 19881
rect 10510 19825 10536 19881
rect 10592 19825 10618 19881
rect 10674 19825 10690 19881
rect 10114 19797 10690 19825
rect 10114 19741 10126 19797
rect 10182 19741 10208 19797
rect 10264 19741 10290 19797
rect 10346 19741 10372 19797
rect 10428 19741 10454 19797
rect 10510 19741 10536 19797
rect 10592 19741 10618 19797
rect 10674 19741 10690 19797
rect 10114 19713 10690 19741
rect 10114 19657 10126 19713
rect 10182 19657 10208 19713
rect 10264 19657 10290 19713
rect 10346 19657 10372 19713
rect 10428 19657 10454 19713
rect 10510 19657 10536 19713
rect 10592 19657 10618 19713
rect 10674 19657 10690 19713
rect 10114 19629 10690 19657
rect 10114 19573 10126 19629
rect 10182 19573 10208 19629
rect 10264 19573 10290 19629
rect 10346 19573 10372 19629
rect 10428 19573 10454 19629
rect 10510 19573 10536 19629
rect 10592 19573 10618 19629
rect 10674 19573 10690 19629
rect 10114 19545 10690 19573
rect 10114 19489 10126 19545
rect 10182 19489 10208 19545
rect 10264 19489 10290 19545
rect 10346 19489 10372 19545
rect 10428 19489 10454 19545
rect 10510 19489 10536 19545
rect 10592 19489 10618 19545
rect 10674 19489 10690 19545
rect 10114 19461 10690 19489
rect 10114 19405 10126 19461
rect 10182 19405 10208 19461
rect 10264 19405 10290 19461
rect 10346 19405 10372 19461
rect 10428 19405 10454 19461
rect 10510 19405 10536 19461
rect 10592 19405 10618 19461
rect 10674 19405 10690 19461
rect 10114 19377 10690 19405
rect 10114 19321 10126 19377
rect 10182 19321 10208 19377
rect 10264 19321 10290 19377
rect 10346 19321 10372 19377
rect 10428 19321 10454 19377
rect 10510 19321 10536 19377
rect 10592 19321 10618 19377
rect 10674 19321 10690 19377
rect 10114 19293 10690 19321
rect 10114 19237 10126 19293
rect 10182 19237 10208 19293
rect 10264 19237 10290 19293
rect 10346 19237 10372 19293
rect 10428 19237 10454 19293
rect 10510 19237 10536 19293
rect 10592 19237 10618 19293
rect 10674 19237 10690 19293
rect 10114 19209 10690 19237
rect 10114 19153 10126 19209
rect 10182 19153 10208 19209
rect 10264 19153 10290 19209
rect 10346 19153 10372 19209
rect 10428 19153 10454 19209
rect 10510 19153 10536 19209
rect 10592 19153 10618 19209
rect 10674 19153 10690 19209
rect 11915 20550 12491 20567
rect 11915 20494 11927 20550
rect 11983 20494 12009 20550
rect 12065 20494 12091 20550
rect 12147 20494 12173 20550
rect 12229 20494 12255 20550
rect 12311 20494 12337 20550
rect 12393 20494 12419 20550
rect 12475 20494 12491 20550
rect 11915 20467 12491 20494
rect 11915 20411 11927 20467
rect 11983 20411 12009 20467
rect 12065 20411 12091 20467
rect 12147 20411 12173 20467
rect 12229 20411 12255 20467
rect 12311 20411 12337 20467
rect 12393 20411 12419 20467
rect 12475 20411 12491 20467
rect 11915 20384 12491 20411
rect 11915 20328 11927 20384
rect 11983 20328 12009 20384
rect 12065 20328 12091 20384
rect 12147 20328 12173 20384
rect 12229 20328 12255 20384
rect 12311 20328 12337 20384
rect 12393 20328 12419 20384
rect 12475 20328 12491 20384
rect 11915 20301 12491 20328
rect 11915 20245 11927 20301
rect 11983 20245 12009 20301
rect 12065 20245 12091 20301
rect 12147 20245 12173 20301
rect 12229 20245 12255 20301
rect 12311 20245 12337 20301
rect 12393 20245 12419 20301
rect 12475 20245 12491 20301
rect 11915 20217 12491 20245
rect 11915 20161 11927 20217
rect 11983 20161 12009 20217
rect 12065 20161 12091 20217
rect 12147 20161 12173 20217
rect 12229 20161 12255 20217
rect 12311 20161 12337 20217
rect 12393 20161 12419 20217
rect 12475 20161 12491 20217
rect 11915 20133 12491 20161
rect 11915 20077 11927 20133
rect 11983 20077 12009 20133
rect 12065 20077 12091 20133
rect 12147 20077 12173 20133
rect 12229 20077 12255 20133
rect 12311 20077 12337 20133
rect 12393 20077 12419 20133
rect 12475 20077 12491 20133
rect 11915 20049 12491 20077
rect 11915 19993 11927 20049
rect 11983 19993 12009 20049
rect 12065 19993 12091 20049
rect 12147 19993 12173 20049
rect 12229 19993 12255 20049
rect 12311 19993 12337 20049
rect 12393 19993 12419 20049
rect 12475 19993 12491 20049
rect 11915 19965 12491 19993
rect 11915 19909 11927 19965
rect 11983 19909 12009 19965
rect 12065 19909 12091 19965
rect 12147 19909 12173 19965
rect 12229 19909 12255 19965
rect 12311 19909 12337 19965
rect 12393 19909 12419 19965
rect 12475 19909 12491 19965
rect 11915 19881 12491 19909
rect 11915 19825 11927 19881
rect 11983 19825 12009 19881
rect 12065 19825 12091 19881
rect 12147 19825 12173 19881
rect 12229 19825 12255 19881
rect 12311 19825 12337 19881
rect 12393 19825 12419 19881
rect 12475 19825 12491 19881
rect 11915 19797 12491 19825
rect 11915 19741 11927 19797
rect 11983 19741 12009 19797
rect 12065 19741 12091 19797
rect 12147 19741 12173 19797
rect 12229 19741 12255 19797
rect 12311 19741 12337 19797
rect 12393 19741 12419 19797
rect 12475 19741 12491 19797
rect 11915 19713 12491 19741
rect 11915 19657 11927 19713
rect 11983 19657 12009 19713
rect 12065 19657 12091 19713
rect 12147 19657 12173 19713
rect 12229 19657 12255 19713
rect 12311 19657 12337 19713
rect 12393 19657 12419 19713
rect 12475 19657 12491 19713
rect 11915 19629 12491 19657
rect 11915 19573 11927 19629
rect 11983 19573 12009 19629
rect 12065 19573 12091 19629
rect 12147 19573 12173 19629
rect 12229 19573 12255 19629
rect 12311 19573 12337 19629
rect 12393 19573 12419 19629
rect 12475 19573 12491 19629
rect 11915 19545 12491 19573
rect 11915 19489 11927 19545
rect 11983 19489 12009 19545
rect 12065 19489 12091 19545
rect 12147 19489 12173 19545
rect 12229 19489 12255 19545
rect 12311 19489 12337 19545
rect 12393 19489 12419 19545
rect 12475 19489 12491 19545
rect 11915 19461 12491 19489
rect 11915 19405 11927 19461
rect 11983 19405 12009 19461
rect 12065 19405 12091 19461
rect 12147 19405 12173 19461
rect 12229 19405 12255 19461
rect 12311 19405 12337 19461
rect 12393 19405 12419 19461
rect 12475 19405 12491 19461
rect 11915 19377 12491 19405
rect 11915 19321 11927 19377
rect 11983 19321 12009 19377
rect 12065 19321 12091 19377
rect 12147 19321 12173 19377
rect 12229 19321 12255 19377
rect 12311 19321 12337 19377
rect 12393 19321 12419 19377
rect 12475 19321 12491 19377
rect 11915 19293 12491 19321
rect 11915 19237 11927 19293
rect 11983 19237 12009 19293
rect 12065 19237 12091 19293
rect 12147 19237 12173 19293
rect 12229 19237 12255 19293
rect 12311 19237 12337 19293
rect 12393 19237 12419 19293
rect 12475 19237 12491 19293
rect 11915 19209 12491 19237
tri 10690 19153 10714 19177 sw
rect 11915 19153 11927 19209
rect 11983 19153 12009 19209
rect 12065 19153 12091 19209
rect 12147 19153 12173 19209
rect 12229 19153 12255 19209
rect 12311 19153 12337 19209
rect 12393 19153 12419 19209
rect 12475 19153 12491 19209
rect 10114 19125 10714 19153
tri 10714 19125 10742 19153 sw
rect 11915 19125 12491 19153
rect 10114 19069 10126 19125
rect 10182 19069 10208 19125
rect 10264 19069 10290 19125
rect 10346 19069 10372 19125
rect 10428 19069 10454 19125
rect 10510 19069 10536 19125
rect 10592 19069 10618 19125
rect 10674 19069 10742 19125
tri 10742 19069 10798 19125 sw
rect 11915 19069 11927 19125
rect 11983 19069 12009 19125
rect 12065 19069 12091 19125
rect 12147 19069 12173 19125
rect 12229 19069 12255 19125
rect 12311 19069 12337 19125
rect 12393 19069 12419 19125
rect 12475 19069 12491 19125
rect 10114 19064 10798 19069
tri 10798 19064 10803 19069 sw
rect 10114 19061 10803 19064
tri 10803 19061 10806 19064 sw
rect 10114 18943 10806 19061
tri 10358 18939 10362 18943 ne
rect 10362 18939 10806 18943
rect 11915 18939 12491 19069
tri 10362 18839 10462 18939 ne
rect 10462 18839 10806 18939
tri 12011 18839 12111 18939 ne
rect 12111 18839 12491 18939
tri 10462 18822 10479 18839 ne
rect 10479 18822 10806 18839
tri 12111 18822 12128 18839 ne
rect 12128 18822 12474 18839
tri 12474 18822 12491 18839 nw
tri 10479 18790 10511 18822 ne
tri 10501 18445 10511 18455 se
rect 10511 18445 10806 18822
tri 12128 18789 12161 18822 ne
rect 9231 18409 9237 18445
rect 8885 18243 9123 18271
tri 9123 18243 9151 18271 nw
rect 9229 18381 9237 18409
rect 9301 18381 9333 18445
rect 9397 18381 9429 18445
rect 9493 18381 9525 18445
rect 9589 18381 9621 18445
rect 9685 18381 9716 18445
rect 9780 18409 9786 18445
tri 10487 18431 10501 18445 se
rect 10501 18431 10806 18445
tri 10465 18409 10487 18431 se
rect 10487 18409 10806 18431
tri 12139 18409 12161 18431 se
rect 12161 18409 12474 18822
rect 9780 18381 9789 18409
tri 10449 18393 10465 18409 se
rect 10465 18393 10806 18409
tri 12123 18393 12139 18409 se
rect 12139 18393 12474 18409
rect 9229 18357 9789 18381
tri 10433 18377 10449 18393 se
rect 10449 18377 10806 18393
tri 12107 18377 12123 18393 se
rect 12123 18377 12474 18393
tri 12474 18377 12490 18393 sw
rect 9229 18293 9237 18357
rect 9301 18293 9333 18357
rect 9397 18293 9429 18357
rect 9493 18293 9525 18357
rect 9589 18293 9621 18357
rect 9685 18293 9716 18357
rect 9780 18293 9789 18357
rect 9229 18269 9789 18293
tri 10337 18281 10433 18377 se
rect 10433 18281 10806 18377
rect 7419 18181 7979 18205
rect 7419 18117 7427 18181
rect 7491 18117 7523 18181
rect 7587 18117 7619 18181
rect 7683 18117 7715 18181
rect 7779 18117 7811 18181
rect 7875 18117 7906 18181
rect 7970 18117 7979 18181
rect 7419 18093 7979 18117
tri 8162 18105 8300 18243 ne
rect 8300 18105 8985 18243
tri 8985 18105 9123 18243 nw
rect 9229 18205 9237 18269
rect 9301 18205 9333 18269
rect 9397 18205 9429 18269
rect 9493 18205 9525 18269
rect 9589 18205 9621 18269
rect 9685 18205 9716 18269
rect 9780 18205 9789 18269
rect 9229 18181 9789 18205
rect 9229 18117 9237 18181
rect 9301 18117 9333 18181
rect 9397 18117 9429 18181
rect 9493 18117 9525 18181
rect 9589 18117 9621 18181
rect 9685 18117 9716 18181
rect 9780 18117 9789 18181
rect 7419 18029 7427 18093
rect 7491 18029 7523 18093
rect 7587 18029 7619 18093
rect 7683 18029 7715 18093
rect 7779 18029 7811 18093
rect 7875 18029 7906 18093
rect 7970 18029 7979 18093
tri 5275 3173 5278 3176 sw
tri 1058 3137 1094 3173 se
rect 1094 3137 1673 3173
tri -3745 2988 -3596 3137 sw
tri -2666 2988 -2517 3137 se
tri -2131 2988 -1982 3137 sw
tri 909 2988 1058 3137 se
rect 1058 2988 1673 3137
tri 1673 2988 1858 3173 sw
tri 2713 2988 2898 3173 se
rect 2898 2988 3477 3173
tri 3477 2988 3662 3173 sw
tri 4514 2988 4699 3173 se
rect 4699 2988 5278 3173
tri 5278 2988 5463 3173 sw
tri 6321 2988 6506 3173 se
rect 6506 2988 7082 12080
rect 7419 3526 7979 18029
rect 8300 13045 8900 18105
tri 8900 18020 8985 18105 nw
rect 9229 18093 9789 18117
rect 9229 18029 9237 18093
rect 9301 18029 9333 18093
rect 9397 18029 9429 18093
rect 9493 18029 9525 18093
rect 9589 18029 9621 18093
rect 9685 18029 9716 18093
rect 9780 18029 9789 18093
rect 8300 12989 8324 13045
rect 8380 12989 8408 13045
rect 8464 12989 8492 13045
rect 8548 12989 8576 13045
rect 8632 12989 8660 13045
rect 8716 12989 8744 13045
rect 8800 12989 8828 13045
rect 8884 12989 8900 13045
rect 8300 12965 8900 12989
rect 8300 12909 8324 12965
rect 8380 12909 8408 12965
rect 8464 12909 8492 12965
rect 8548 12909 8576 12965
rect 8632 12909 8660 12965
rect 8716 12909 8744 12965
rect 8800 12909 8828 12965
rect 8884 12909 8900 12965
rect 8300 12885 8900 12909
rect 8300 12829 8324 12885
rect 8380 12829 8408 12885
rect 8464 12829 8492 12885
rect 8548 12829 8576 12885
rect 8632 12829 8660 12885
rect 8716 12829 8744 12885
rect 8800 12829 8828 12885
rect 8884 12829 8900 12885
rect 8300 12805 8900 12829
rect 8300 12749 8324 12805
rect 8380 12749 8408 12805
rect 8464 12749 8492 12805
rect 8548 12749 8576 12805
rect 8632 12749 8660 12805
rect 8716 12749 8744 12805
rect 8800 12749 8828 12805
rect 8884 12749 8900 12805
rect 8300 12725 8900 12749
rect 8300 12669 8324 12725
rect 8380 12669 8408 12725
rect 8464 12669 8492 12725
rect 8548 12669 8576 12725
rect 8632 12669 8660 12725
rect 8716 12669 8744 12725
rect 8800 12669 8828 12725
rect 8884 12669 8900 12725
rect 8300 12645 8900 12669
rect 8300 12589 8324 12645
rect 8380 12589 8408 12645
rect 8464 12589 8492 12645
rect 8548 12589 8576 12645
rect 8632 12589 8660 12645
rect 8716 12589 8744 12645
rect 8800 12589 8828 12645
rect 8884 12589 8900 12645
rect 8300 12565 8900 12589
rect 8300 12509 8324 12565
rect 8380 12509 8408 12565
rect 8464 12509 8492 12565
rect 8548 12509 8576 12565
rect 8632 12509 8660 12565
rect 8716 12509 8744 12565
rect 8800 12509 8828 12565
rect 8884 12509 8900 12565
rect 8300 12485 8900 12509
rect 8300 12429 8324 12485
rect 8380 12429 8408 12485
rect 8464 12429 8492 12485
rect 8548 12429 8576 12485
rect 8632 12429 8660 12485
rect 8716 12429 8744 12485
rect 8800 12429 8828 12485
rect 8884 12429 8900 12485
rect 8300 12405 8900 12429
rect 8300 12349 8324 12405
rect 8380 12349 8408 12405
rect 8464 12349 8492 12405
rect 8548 12349 8576 12405
rect 8632 12349 8660 12405
rect 8716 12349 8744 12405
rect 8800 12349 8828 12405
rect 8884 12349 8900 12405
rect 8300 12325 8900 12349
rect 8300 12269 8324 12325
rect 8380 12269 8408 12325
rect 8464 12269 8492 12325
rect 8548 12269 8576 12325
rect 8632 12269 8660 12325
rect 8716 12269 8744 12325
rect 8800 12269 8828 12325
rect 8884 12269 8900 12325
rect 8300 12245 8900 12269
rect 8300 12189 8324 12245
rect 8380 12189 8408 12245
rect 8464 12189 8492 12245
rect 8548 12189 8576 12245
rect 8632 12189 8660 12245
rect 8716 12189 8744 12245
rect 8800 12189 8828 12245
rect 8884 12189 8900 12245
rect 8300 12165 8900 12189
rect 8300 12109 8324 12165
rect 8380 12109 8408 12165
rect 8464 12109 8492 12165
rect 8548 12109 8576 12165
rect 8632 12109 8660 12165
rect 8716 12109 8744 12165
rect 8800 12109 8828 12165
rect 8884 12109 8900 12165
rect 8300 12085 8900 12109
rect 8300 12029 8324 12085
rect 8380 12029 8408 12085
rect 8464 12029 8492 12085
rect 8548 12029 8576 12085
rect 8632 12029 8660 12085
rect 8716 12029 8744 12085
rect 8800 12029 8828 12085
rect 8884 12029 8900 12085
rect 8300 12005 8900 12029
rect 8300 11949 8324 12005
rect 8380 11949 8408 12005
rect 8464 11949 8492 12005
rect 8548 11949 8576 12005
rect 8632 11949 8660 12005
rect 8716 11949 8744 12005
rect 8800 11949 8828 12005
rect 8884 11949 8900 12005
rect 8300 11925 8900 11949
rect 8300 11869 8324 11925
rect 8380 11869 8408 11925
rect 8464 11869 8492 11925
rect 8548 11869 8576 11925
rect 8632 11869 8660 11925
rect 8716 11869 8744 11925
rect 8800 11869 8828 11925
rect 8884 11869 8900 11925
rect 8300 11845 8900 11869
rect 8300 11789 8324 11845
rect 8380 11789 8408 11845
rect 8464 11789 8492 11845
rect 8548 11789 8576 11845
rect 8632 11789 8660 11845
rect 8716 11789 8744 11845
rect 8800 11789 8828 11845
rect 8884 11789 8900 11845
rect 8300 11765 8900 11789
rect 8300 11709 8324 11765
rect 8380 11709 8408 11765
rect 8464 11709 8492 11765
rect 8548 11709 8576 11765
rect 8632 11709 8660 11765
rect 8716 11709 8744 11765
rect 8800 11709 8828 11765
rect 8884 11709 8900 11765
rect 8300 11685 8900 11709
rect 8300 11629 8324 11685
rect 8380 11629 8408 11685
rect 8464 11629 8492 11685
rect 8548 11629 8576 11685
rect 8632 11629 8660 11685
rect 8716 11629 8744 11685
rect 8800 11629 8828 11685
rect 8884 11629 8900 11685
rect 8300 11605 8900 11629
rect 8300 11549 8324 11605
rect 8380 11549 8408 11605
rect 8464 11549 8492 11605
rect 8548 11549 8576 11605
rect 8632 11549 8660 11605
rect 8716 11549 8744 11605
rect 8800 11549 8828 11605
rect 8884 11549 8900 11605
rect 8300 11525 8900 11549
rect 8300 11469 8324 11525
rect 8380 11469 8408 11525
rect 8464 11469 8492 11525
rect 8548 11469 8576 11525
rect 8632 11469 8660 11525
rect 8716 11469 8744 11525
rect 8800 11469 8828 11525
rect 8884 11469 8900 11525
rect 8300 11445 8900 11469
rect 8300 11389 8324 11445
rect 8380 11389 8408 11445
rect 8464 11389 8492 11445
rect 8548 11389 8576 11445
rect 8632 11389 8660 11445
rect 8716 11389 8744 11445
rect 8800 11389 8828 11445
rect 8884 11389 8900 11445
rect 8300 11365 8900 11389
rect 8300 11309 8324 11365
rect 8380 11309 8408 11365
rect 8464 11309 8492 11365
rect 8548 11309 8576 11365
rect 8632 11309 8660 11365
rect 8716 11309 8744 11365
rect 8800 11309 8828 11365
rect 8884 11309 8900 11365
rect 8300 11285 8900 11309
rect 8300 11229 8324 11285
rect 8380 11229 8408 11285
rect 8464 11229 8492 11285
rect 8548 11229 8576 11285
rect 8632 11229 8660 11285
rect 8716 11229 8744 11285
rect 8800 11229 8828 11285
rect 8884 11229 8900 11285
rect 8300 11205 8900 11229
rect 8300 11149 8324 11205
rect 8380 11149 8408 11205
rect 8464 11149 8492 11205
rect 8548 11149 8576 11205
rect 8632 11149 8660 11205
rect 8716 11149 8744 11205
rect 8800 11149 8828 11205
rect 8884 11149 8900 11205
rect 8300 11125 8900 11149
rect 8300 11069 8324 11125
rect 8380 11069 8408 11125
rect 8464 11069 8492 11125
rect 8548 11069 8576 11125
rect 8632 11069 8660 11125
rect 8716 11069 8744 11125
rect 8800 11069 8828 11125
rect 8884 11069 8900 11125
rect 8300 11045 8900 11069
rect 8300 10989 8324 11045
rect 8380 10989 8408 11045
rect 8464 10989 8492 11045
rect 8548 10989 8576 11045
rect 8632 10989 8660 11045
rect 8716 10989 8744 11045
rect 8800 10989 8828 11045
rect 8884 10989 8900 11045
rect 8300 10965 8900 10989
rect 8300 10909 8324 10965
rect 8380 10909 8408 10965
rect 8464 10909 8492 10965
rect 8548 10909 8576 10965
rect 8632 10909 8660 10965
rect 8716 10909 8744 10965
rect 8800 10909 8828 10965
rect 8884 10909 8900 10965
rect 8300 10885 8900 10909
rect 8300 10829 8324 10885
rect 8380 10829 8408 10885
rect 8464 10829 8492 10885
rect 8548 10829 8576 10885
rect 8632 10829 8660 10885
rect 8716 10829 8744 10885
rect 8800 10829 8828 10885
rect 8884 10829 8900 10885
rect 8300 10805 8900 10829
rect 8300 10749 8324 10805
rect 8380 10749 8408 10805
rect 8464 10749 8492 10805
rect 8548 10749 8576 10805
rect 8632 10749 8660 10805
rect 8716 10749 8744 10805
rect 8800 10749 8828 10805
rect 8884 10749 8900 10805
rect 8300 10725 8900 10749
rect 8300 10669 8324 10725
rect 8380 10669 8408 10725
rect 8464 10669 8492 10725
rect 8548 10669 8576 10725
rect 8632 10669 8660 10725
rect 8716 10669 8744 10725
rect 8800 10669 8828 10725
rect 8884 10669 8900 10725
rect 8300 10645 8900 10669
rect 8300 10589 8324 10645
rect 8380 10589 8408 10645
rect 8464 10589 8492 10645
rect 8548 10589 8576 10645
rect 8632 10589 8660 10645
rect 8716 10589 8744 10645
rect 8800 10589 8828 10645
rect 8884 10589 8900 10645
rect 8300 10565 8900 10589
rect 8300 10509 8324 10565
rect 8380 10509 8408 10565
rect 8464 10509 8492 10565
rect 8548 10509 8576 10565
rect 8632 10509 8660 10565
rect 8716 10509 8744 10565
rect 8800 10509 8828 10565
rect 8884 10509 8900 10565
rect 8300 10485 8900 10509
rect 8300 10429 8324 10485
rect 8380 10429 8408 10485
rect 8464 10429 8492 10485
rect 8548 10429 8576 10485
rect 8632 10429 8660 10485
rect 8716 10429 8744 10485
rect 8800 10429 8828 10485
rect 8884 10429 8900 10485
rect 8300 10405 8900 10429
rect 8300 10349 8324 10405
rect 8380 10349 8408 10405
rect 8464 10349 8492 10405
rect 8548 10349 8576 10405
rect 8632 10349 8660 10405
rect 8716 10349 8744 10405
rect 8800 10349 8828 10405
rect 8884 10349 8900 10405
rect 8300 10325 8900 10349
rect 8300 10269 8324 10325
rect 8380 10269 8408 10325
rect 8464 10269 8492 10325
rect 8548 10269 8576 10325
rect 8632 10269 8660 10325
rect 8716 10269 8744 10325
rect 8800 10269 8828 10325
rect 8884 10269 8900 10325
rect 8300 10245 8900 10269
rect 8300 10189 8324 10245
rect 8380 10189 8408 10245
rect 8464 10189 8492 10245
rect 8548 10189 8576 10245
rect 8632 10189 8660 10245
rect 8716 10189 8744 10245
rect 8800 10189 8828 10245
rect 8884 10189 8900 10245
rect 8300 10165 8900 10189
rect 8300 10109 8324 10165
rect 8380 10109 8408 10165
rect 8464 10109 8492 10165
rect 8548 10109 8576 10165
rect 8632 10109 8660 10165
rect 8716 10109 8744 10165
rect 8800 10109 8828 10165
rect 8884 10109 8900 10165
rect 8300 10085 8900 10109
rect 8300 10029 8324 10085
rect 8380 10029 8408 10085
rect 8464 10029 8492 10085
rect 8548 10029 8576 10085
rect 8632 10029 8660 10085
rect 8716 10029 8744 10085
rect 8800 10029 8828 10085
rect 8884 10029 8900 10085
rect 8300 10005 8900 10029
rect 8300 9949 8324 10005
rect 8380 9949 8408 10005
rect 8464 9949 8492 10005
rect 8548 9949 8576 10005
rect 8632 9949 8660 10005
rect 8716 9949 8744 10005
rect 8800 9949 8828 10005
rect 8884 9949 8900 10005
rect 8300 9925 8900 9949
rect 8300 9869 8324 9925
rect 8380 9869 8408 9925
rect 8464 9869 8492 9925
rect 8548 9869 8576 9925
rect 8632 9869 8660 9925
rect 8716 9869 8744 9925
rect 8800 9869 8828 9925
rect 8884 9869 8900 9925
rect 8300 9845 8900 9869
rect 8300 9789 8324 9845
rect 8380 9789 8408 9845
rect 8464 9789 8492 9845
rect 8548 9789 8576 9845
rect 8632 9789 8660 9845
rect 8716 9789 8744 9845
rect 8800 9789 8828 9845
rect 8884 9789 8900 9845
rect 8300 9765 8900 9789
rect 8300 9709 8324 9765
rect 8380 9709 8408 9765
rect 8464 9709 8492 9765
rect 8548 9709 8576 9765
rect 8632 9709 8660 9765
rect 8716 9709 8744 9765
rect 8800 9709 8828 9765
rect 8884 9709 8900 9765
rect 8300 9685 8900 9709
rect 8300 9629 8324 9685
rect 8380 9629 8408 9685
rect 8464 9629 8492 9685
rect 8548 9629 8576 9685
rect 8632 9629 8660 9685
rect 8716 9629 8744 9685
rect 8800 9629 8828 9685
rect 8884 9629 8900 9685
rect 8300 9605 8900 9629
rect 8300 9549 8324 9605
rect 8380 9549 8408 9605
rect 8464 9549 8492 9605
rect 8548 9549 8576 9605
rect 8632 9549 8660 9605
rect 8716 9549 8744 9605
rect 8800 9549 8828 9605
rect 8884 9549 8900 9605
rect 8300 9524 8900 9549
rect 8300 9468 8324 9524
rect 8380 9468 8408 9524
rect 8464 9468 8492 9524
rect 8548 9468 8576 9524
rect 8632 9468 8660 9524
rect 8716 9468 8744 9524
rect 8800 9468 8828 9524
rect 8884 9468 8900 9524
rect 8300 9443 8900 9468
rect 8300 9387 8324 9443
rect 8380 9387 8408 9443
rect 8464 9387 8492 9443
rect 8548 9387 8576 9443
rect 8632 9387 8660 9443
rect 8716 9387 8744 9443
rect 8800 9387 8828 9443
rect 8884 9387 8900 9443
rect 8300 9362 8900 9387
rect 8300 9306 8324 9362
rect 8380 9306 8408 9362
rect 8464 9306 8492 9362
rect 8548 9306 8576 9362
rect 8632 9306 8660 9362
rect 8716 9306 8744 9362
rect 8800 9306 8828 9362
rect 8884 9306 8900 9362
rect 8300 9281 8900 9306
rect 8300 9225 8324 9281
rect 8380 9225 8408 9281
rect 8464 9225 8492 9281
rect 8548 9225 8576 9281
rect 8632 9225 8660 9281
rect 8716 9225 8744 9281
rect 8800 9225 8828 9281
rect 8884 9225 8900 9281
rect 8300 9200 8900 9225
rect 8300 9144 8324 9200
rect 8380 9144 8408 9200
rect 8464 9144 8492 9200
rect 8548 9144 8576 9200
rect 8632 9144 8660 9200
rect 8716 9144 8744 9200
rect 8800 9144 8828 9200
rect 8884 9144 8900 9200
rect 8300 9119 8900 9144
rect 8300 9063 8324 9119
rect 8380 9063 8408 9119
rect 8464 9063 8492 9119
rect 8548 9063 8576 9119
rect 8632 9063 8660 9119
rect 8716 9063 8744 9119
rect 8800 9063 8828 9119
rect 8884 9063 8900 9119
rect 8300 9038 8900 9063
rect 8300 8982 8324 9038
rect 8380 8982 8408 9038
rect 8464 8982 8492 9038
rect 8548 8982 8576 9038
rect 8632 8982 8660 9038
rect 8716 8982 8744 9038
rect 8800 8982 8828 9038
rect 8884 8982 8900 9038
rect 8300 8957 8900 8982
rect 8300 8901 8324 8957
rect 8380 8901 8408 8957
rect 8464 8901 8492 8957
rect 8548 8901 8576 8957
rect 8632 8901 8660 8957
rect 8716 8901 8744 8957
rect 8800 8901 8828 8957
rect 8884 8901 8900 8957
rect 8300 8876 8900 8901
rect 8300 8820 8324 8876
rect 8380 8820 8408 8876
rect 8464 8820 8492 8876
rect 8548 8820 8576 8876
rect 8632 8820 8660 8876
rect 8716 8820 8744 8876
rect 8800 8820 8828 8876
rect 8884 8820 8900 8876
rect 8300 8795 8900 8820
rect 8300 8739 8324 8795
rect 8380 8739 8408 8795
rect 8464 8739 8492 8795
rect 8548 8739 8576 8795
rect 8632 8739 8660 8795
rect 8716 8739 8744 8795
rect 8800 8739 8828 8795
rect 8884 8739 8900 8795
rect 8300 8714 8900 8739
rect 8300 8658 8324 8714
rect 8380 8658 8408 8714
rect 8464 8658 8492 8714
rect 8548 8658 8576 8714
rect 8632 8658 8660 8714
rect 8716 8658 8744 8714
rect 8800 8658 8828 8714
rect 8884 8658 8900 8714
rect 8300 8633 8900 8658
rect 8300 8577 8324 8633
rect 8380 8577 8408 8633
rect 8464 8577 8492 8633
rect 8548 8577 8576 8633
rect 8632 8577 8660 8633
rect 8716 8577 8744 8633
rect 8800 8577 8828 8633
rect 8884 8577 8900 8633
rect 8300 8552 8900 8577
rect 8300 8496 8324 8552
rect 8380 8496 8408 8552
rect 8464 8496 8492 8552
rect 8548 8496 8576 8552
rect 8632 8496 8660 8552
rect 8716 8496 8744 8552
rect 8800 8496 8828 8552
rect 8884 8496 8900 8552
rect 8300 8471 8900 8496
rect 8300 8415 8324 8471
rect 8380 8415 8408 8471
rect 8464 8415 8492 8471
rect 8548 8415 8576 8471
rect 8632 8415 8660 8471
rect 8716 8415 8744 8471
rect 8800 8415 8828 8471
rect 8884 8415 8900 8471
rect 8300 8390 8900 8415
rect 8300 8334 8324 8390
rect 8380 8334 8408 8390
rect 8464 8334 8492 8390
rect 8548 8334 8576 8390
rect 8632 8334 8660 8390
rect 8716 8334 8744 8390
rect 8800 8334 8828 8390
rect 8884 8334 8900 8390
rect 8300 8309 8900 8334
rect 8300 8253 8324 8309
rect 8380 8253 8408 8309
rect 8464 8253 8492 8309
rect 8548 8253 8576 8309
rect 8632 8253 8660 8309
rect 8716 8253 8744 8309
rect 8800 8253 8828 8309
rect 8884 8253 8900 8309
rect 8300 8228 8900 8253
rect 8300 8172 8324 8228
rect 8380 8172 8408 8228
rect 8464 8172 8492 8228
rect 8548 8172 8576 8228
rect 8632 8172 8660 8228
rect 8716 8172 8744 8228
rect 8800 8172 8828 8228
rect 8884 8172 8900 8228
rect 8300 8147 8900 8172
rect 8300 8091 8324 8147
rect 8380 8091 8408 8147
rect 8464 8091 8492 8147
rect 8548 8091 8576 8147
rect 8632 8091 8660 8147
rect 8716 8091 8744 8147
rect 8800 8091 8828 8147
rect 8884 8091 8900 8147
rect 8300 8066 8900 8091
rect 8300 8010 8324 8066
rect 8380 8010 8408 8066
rect 8464 8010 8492 8066
rect 8548 8010 8576 8066
rect 8632 8010 8660 8066
rect 8716 8010 8744 8066
rect 8800 8010 8828 8066
rect 8884 8010 8900 8066
rect 8300 7985 8900 8010
rect 8300 7929 8324 7985
rect 8380 7929 8408 7985
rect 8464 7929 8492 7985
rect 8548 7929 8576 7985
rect 8632 7929 8660 7985
rect 8716 7929 8744 7985
rect 8800 7929 8828 7985
rect 8884 7929 8900 7985
rect 8300 7904 8900 7929
rect 8300 7848 8324 7904
rect 8380 7848 8408 7904
rect 8464 7848 8492 7904
rect 8548 7848 8576 7904
rect 8632 7848 8660 7904
rect 8716 7848 8744 7904
rect 8800 7848 8828 7904
rect 8884 7848 8900 7904
rect 8300 7823 8900 7848
rect 8300 7767 8324 7823
rect 8380 7767 8408 7823
rect 8464 7767 8492 7823
rect 8548 7767 8576 7823
rect 8632 7767 8660 7823
rect 8716 7767 8744 7823
rect 8800 7767 8828 7823
rect 8884 7767 8900 7823
rect 8300 7742 8900 7767
rect 8300 7686 8324 7742
rect 8380 7686 8408 7742
rect 8464 7686 8492 7742
rect 8548 7686 8576 7742
rect 8632 7686 8660 7742
rect 8716 7686 8744 7742
rect 8800 7686 8828 7742
rect 8884 7686 8900 7742
rect 8300 7661 8900 7686
rect 8300 7605 8324 7661
rect 8380 7605 8408 7661
rect 8464 7605 8492 7661
rect 8548 7605 8576 7661
rect 8632 7605 8660 7661
rect 8716 7605 8744 7661
rect 8800 7605 8828 7661
rect 8884 7605 8900 7661
rect 8300 7580 8900 7605
rect 8300 7524 8324 7580
rect 8380 7524 8408 7580
rect 8464 7524 8492 7580
rect 8548 7524 8576 7580
rect 8632 7524 8660 7580
rect 8716 7524 8744 7580
rect 8800 7524 8828 7580
rect 8884 7524 8900 7580
rect 8300 7499 8900 7524
rect 8300 7443 8324 7499
rect 8380 7443 8408 7499
rect 8464 7443 8492 7499
rect 8548 7443 8576 7499
rect 8632 7443 8660 7499
rect 8716 7443 8744 7499
rect 8800 7443 8828 7499
rect 8884 7443 8900 7499
rect 8300 7418 8900 7443
rect 8300 7362 8324 7418
rect 8380 7362 8408 7418
rect 8464 7362 8492 7418
rect 8548 7362 8576 7418
rect 8632 7362 8660 7418
rect 8716 7362 8744 7418
rect 8800 7362 8828 7418
rect 8884 7362 8900 7418
rect 8300 7337 8900 7362
rect 8300 7281 8324 7337
rect 8380 7281 8408 7337
rect 8464 7281 8492 7337
rect 8548 7281 8576 7337
rect 8632 7281 8660 7337
rect 8716 7281 8744 7337
rect 8800 7281 8828 7337
rect 8884 7281 8900 7337
rect 8300 7256 8900 7281
rect 8300 7200 8324 7256
rect 8380 7200 8408 7256
rect 8464 7200 8492 7256
rect 8548 7200 8576 7256
rect 8632 7200 8660 7256
rect 8716 7200 8744 7256
rect 8800 7200 8828 7256
rect 8884 7200 8900 7256
rect 8300 7175 8900 7200
rect 8300 7119 8324 7175
rect 8380 7119 8408 7175
rect 8464 7119 8492 7175
rect 8548 7119 8576 7175
rect 8632 7119 8660 7175
rect 8716 7119 8744 7175
rect 8800 7119 8828 7175
rect 8884 7119 8900 7175
rect 8300 7094 8900 7119
rect 8300 7038 8324 7094
rect 8380 7038 8408 7094
rect 8464 7038 8492 7094
rect 8548 7038 8576 7094
rect 8632 7038 8660 7094
rect 8716 7038 8744 7094
rect 8800 7038 8828 7094
rect 8884 7038 8900 7094
rect 8300 7013 8900 7038
rect 8300 6957 8324 7013
rect 8380 6957 8408 7013
rect 8464 6957 8492 7013
rect 8548 6957 8576 7013
rect 8632 6957 8660 7013
rect 8716 6957 8744 7013
rect 8800 6957 8828 7013
rect 8884 6957 8900 7013
rect 8300 6932 8900 6957
rect 8300 6876 8324 6932
rect 8380 6876 8408 6932
rect 8464 6876 8492 6932
rect 8548 6876 8576 6932
rect 8632 6876 8660 6932
rect 8716 6876 8744 6932
rect 8800 6876 8828 6932
rect 8884 6876 8900 6932
rect 8300 6851 8900 6876
rect 8300 6795 8324 6851
rect 8380 6795 8408 6851
rect 8464 6795 8492 6851
rect 8548 6795 8576 6851
rect 8632 6795 8660 6851
rect 8716 6795 8744 6851
rect 8800 6795 8828 6851
rect 8884 6795 8900 6851
rect 8300 6770 8900 6795
rect 8300 6714 8324 6770
rect 8380 6714 8408 6770
rect 8464 6714 8492 6770
rect 8548 6714 8576 6770
rect 8632 6714 8660 6770
rect 8716 6714 8744 6770
rect 8800 6714 8828 6770
rect 8884 6714 8900 6770
rect 8300 6689 8900 6714
rect 8300 6633 8324 6689
rect 8380 6633 8408 6689
rect 8464 6633 8492 6689
rect 8548 6633 8576 6689
rect 8632 6633 8660 6689
rect 8716 6633 8744 6689
rect 8800 6633 8828 6689
rect 8884 6633 8900 6689
rect 8300 6608 8900 6633
rect 8300 6552 8324 6608
rect 8380 6552 8408 6608
rect 8464 6552 8492 6608
rect 8548 6552 8576 6608
rect 8632 6552 8660 6608
rect 8716 6552 8744 6608
rect 8800 6552 8828 6608
rect 8884 6552 8900 6608
rect 8300 6527 8900 6552
rect 8300 6471 8324 6527
rect 8380 6471 8408 6527
rect 8464 6471 8492 6527
rect 8548 6471 8576 6527
rect 8632 6471 8660 6527
rect 8716 6471 8744 6527
rect 8800 6471 8828 6527
rect 8884 6471 8900 6527
rect 8300 6446 8900 6471
rect 8300 6390 8324 6446
rect 8380 6390 8408 6446
rect 8464 6390 8492 6446
rect 8548 6390 8576 6446
rect 8632 6390 8660 6446
rect 8716 6390 8744 6446
rect 8800 6390 8828 6446
rect 8884 6390 8900 6446
rect 8300 6365 8900 6390
rect 8300 6309 8324 6365
rect 8380 6309 8408 6365
rect 8464 6309 8492 6365
rect 8548 6309 8576 6365
rect 8632 6309 8660 6365
rect 8716 6309 8744 6365
rect 8800 6309 8828 6365
rect 8884 6309 8900 6365
rect 8300 6284 8900 6309
rect 8300 6228 8324 6284
rect 8380 6228 8408 6284
rect 8464 6228 8492 6284
rect 8548 6228 8576 6284
rect 8632 6228 8660 6284
rect 8716 6228 8744 6284
rect 8800 6228 8828 6284
rect 8884 6228 8900 6284
rect 8300 6203 8900 6228
rect 8300 6147 8324 6203
rect 8380 6147 8408 6203
rect 8464 6147 8492 6203
rect 8548 6147 8576 6203
rect 8632 6147 8660 6203
rect 8716 6147 8744 6203
rect 8800 6147 8828 6203
rect 8884 6147 8900 6203
rect 8300 6122 8900 6147
rect 8300 6066 8324 6122
rect 8380 6066 8408 6122
rect 8464 6066 8492 6122
rect 8548 6066 8576 6122
rect 8632 6066 8660 6122
rect 8716 6066 8744 6122
rect 8800 6066 8828 6122
rect 8884 6066 8900 6122
rect 8300 6041 8900 6066
rect 8300 5985 8324 6041
rect 8380 5985 8408 6041
rect 8464 5985 8492 6041
rect 8548 5985 8576 6041
rect 8632 5985 8660 6041
rect 8716 5985 8744 6041
rect 8800 5985 8828 6041
rect 8884 5985 8900 6041
rect 8300 5960 8900 5985
rect 8300 5904 8324 5960
rect 8380 5904 8408 5960
rect 8464 5904 8492 5960
rect 8548 5904 8576 5960
rect 8632 5904 8660 5960
rect 8716 5904 8744 5960
rect 8800 5904 8828 5960
rect 8884 5904 8900 5960
rect 8300 5879 8900 5904
rect 8300 5823 8324 5879
rect 8380 5823 8408 5879
rect 8464 5823 8492 5879
rect 8548 5823 8576 5879
rect 8632 5823 8660 5879
rect 8716 5823 8744 5879
rect 8800 5823 8828 5879
rect 8884 5823 8900 5879
rect 8300 5798 8900 5823
rect 8300 5742 8324 5798
rect 8380 5742 8408 5798
rect 8464 5742 8492 5798
rect 8548 5742 8576 5798
rect 8632 5742 8660 5798
rect 8716 5742 8744 5798
rect 8800 5742 8828 5798
rect 8884 5742 8900 5798
rect 8300 5717 8900 5742
rect 8300 5661 8324 5717
rect 8380 5661 8408 5717
rect 8464 5661 8492 5717
rect 8548 5661 8576 5717
rect 8632 5661 8660 5717
rect 8716 5661 8744 5717
rect 8800 5661 8828 5717
rect 8884 5661 8900 5717
rect 8300 5636 8900 5661
rect 8300 5580 8324 5636
rect 8380 5580 8408 5636
rect 8464 5580 8492 5636
rect 8548 5580 8576 5636
rect 8632 5580 8660 5636
rect 8716 5580 8744 5636
rect 8800 5580 8828 5636
rect 8884 5580 8900 5636
rect 8300 5555 8900 5580
rect 8300 5499 8324 5555
rect 8380 5499 8408 5555
rect 8464 5499 8492 5555
rect 8548 5499 8576 5555
rect 8632 5499 8660 5555
rect 8716 5499 8744 5555
rect 8800 5499 8828 5555
rect 8884 5499 8900 5555
rect 8300 5474 8900 5499
rect 8300 5418 8324 5474
rect 8380 5418 8408 5474
rect 8464 5418 8492 5474
rect 8548 5418 8576 5474
rect 8632 5418 8660 5474
rect 8716 5418 8744 5474
rect 8800 5418 8828 5474
rect 8884 5418 8900 5474
rect 8300 5393 8900 5418
rect 8300 5337 8324 5393
rect 8380 5337 8408 5393
rect 8464 5337 8492 5393
rect 8548 5337 8576 5393
rect 8632 5337 8660 5393
rect 8716 5337 8744 5393
rect 8800 5337 8828 5393
rect 8884 5337 8900 5393
rect 8300 5312 8900 5337
rect 8300 5256 8324 5312
rect 8380 5256 8408 5312
rect 8464 5256 8492 5312
rect 8548 5256 8576 5312
rect 8632 5256 8660 5312
rect 8716 5256 8744 5312
rect 8800 5256 8828 5312
rect 8884 5256 8900 5312
rect 8300 5231 8900 5256
rect 8300 5175 8324 5231
rect 8380 5175 8408 5231
rect 8464 5175 8492 5231
rect 8548 5175 8576 5231
rect 8632 5175 8660 5231
rect 8716 5175 8744 5231
rect 8800 5175 8828 5231
rect 8884 5175 8900 5231
rect 8300 5150 8900 5175
rect 8300 5094 8324 5150
rect 8380 5094 8408 5150
rect 8464 5094 8492 5150
rect 8548 5094 8576 5150
rect 8632 5094 8660 5150
rect 8716 5094 8744 5150
rect 8800 5094 8828 5150
rect 8884 5094 8900 5150
rect 8300 5069 8900 5094
rect 8300 5013 8324 5069
rect 8380 5013 8408 5069
rect 8464 5013 8492 5069
rect 8548 5013 8576 5069
rect 8632 5013 8660 5069
rect 8716 5013 8744 5069
rect 8800 5013 8828 5069
rect 8884 5013 8900 5069
rect 8300 4988 8900 5013
rect 8300 4932 8324 4988
rect 8380 4932 8408 4988
rect 8464 4932 8492 4988
rect 8548 4932 8576 4988
rect 8632 4932 8660 4988
rect 8716 4932 8744 4988
rect 8800 4932 8828 4988
rect 8884 4932 8900 4988
rect 8300 4907 8900 4932
rect 8300 4851 8324 4907
rect 8380 4851 8408 4907
rect 8464 4851 8492 4907
rect 8548 4851 8576 4907
rect 8632 4851 8660 4907
rect 8716 4851 8744 4907
rect 8800 4851 8828 4907
rect 8884 4851 8900 4907
rect 8300 4826 8900 4851
rect 8300 4770 8324 4826
rect 8380 4770 8408 4826
rect 8464 4770 8492 4826
rect 8548 4770 8576 4826
rect 8632 4770 8660 4826
rect 8716 4770 8744 4826
rect 8800 4770 8828 4826
rect 8884 4770 8900 4826
rect 8300 4745 8900 4770
rect 8300 4689 8324 4745
rect 8380 4689 8408 4745
rect 8464 4689 8492 4745
rect 8548 4689 8576 4745
rect 8632 4689 8660 4745
rect 8716 4689 8744 4745
rect 8800 4689 8828 4745
rect 8884 4689 8900 4745
rect 8300 4664 8900 4689
rect 8300 4608 8324 4664
rect 8380 4608 8408 4664
rect 8464 4608 8492 4664
rect 8548 4608 8576 4664
rect 8632 4608 8660 4664
rect 8716 4608 8744 4664
rect 8800 4608 8828 4664
rect 8884 4608 8900 4664
rect 8300 4583 8900 4608
rect 8300 4527 8324 4583
rect 8380 4527 8408 4583
rect 8464 4527 8492 4583
rect 8548 4527 8576 4583
rect 8632 4527 8660 4583
rect 8716 4527 8744 4583
rect 8800 4527 8828 4583
rect 8884 4527 8900 4583
rect 8300 4502 8900 4527
rect 8300 4446 8324 4502
rect 8380 4446 8408 4502
rect 8464 4446 8492 4502
rect 8548 4446 8576 4502
rect 8632 4446 8660 4502
rect 8716 4446 8744 4502
rect 8800 4446 8828 4502
rect 8884 4446 8900 4502
rect 8300 4421 8900 4446
rect 8300 4365 8324 4421
rect 8380 4365 8408 4421
rect 8464 4365 8492 4421
rect 8548 4365 8576 4421
rect 8632 4365 8660 4421
rect 8716 4365 8744 4421
rect 8800 4365 8828 4421
rect 8884 4365 8900 4421
rect 8300 4340 8900 4365
rect 8300 4284 8324 4340
rect 8380 4284 8408 4340
rect 8464 4284 8492 4340
rect 8548 4284 8576 4340
rect 8632 4284 8660 4340
rect 8716 4284 8744 4340
rect 8800 4284 8828 4340
rect 8884 4284 8900 4340
rect 8300 4259 8900 4284
rect 8300 4203 8324 4259
rect 8380 4203 8408 4259
rect 8464 4203 8492 4259
rect 8548 4203 8576 4259
rect 8632 4203 8660 4259
rect 8716 4203 8744 4259
rect 8800 4203 8828 4259
rect 8884 4203 8900 4259
rect 8300 4178 8900 4203
rect 8300 4122 8324 4178
rect 8380 4122 8408 4178
rect 8464 4122 8492 4178
rect 8548 4122 8576 4178
rect 8632 4122 8660 4178
rect 8716 4122 8744 4178
rect 8800 4122 8828 4178
rect 8884 4122 8900 4178
rect 8300 4097 8900 4122
rect 8300 4041 8324 4097
rect 8380 4041 8408 4097
rect 8464 4041 8492 4097
rect 8548 4041 8576 4097
rect 8632 4041 8660 4097
rect 8716 4041 8744 4097
rect 8800 4041 8828 4097
rect 8884 4041 8900 4097
rect 8300 4016 8900 4041
rect 8300 3960 8324 4016
rect 8380 3960 8408 4016
rect 8464 3960 8492 4016
rect 8548 3960 8576 4016
rect 8632 3960 8660 4016
rect 8716 3960 8744 4016
rect 8800 3960 8828 4016
rect 8884 3960 8900 4016
rect 8300 3935 8900 3960
rect 8300 3879 8324 3935
rect 8380 3879 8408 3935
rect 8464 3879 8492 3935
rect 8548 3879 8576 3935
rect 8632 3879 8660 3935
rect 8716 3879 8744 3935
rect 8800 3879 8828 3935
rect 8884 3879 8900 3935
rect 8300 3854 8900 3879
rect 8300 3798 8324 3854
rect 8380 3798 8408 3854
rect 8464 3798 8492 3854
rect 8548 3798 8576 3854
rect 8632 3798 8660 3854
rect 8716 3798 8744 3854
rect 8800 3798 8828 3854
rect 8884 3798 8900 3854
rect 8300 3773 8900 3798
rect 8300 3717 8324 3773
rect 8380 3717 8408 3773
rect 8464 3717 8492 3773
rect 8548 3717 8576 3773
rect 8632 3717 8660 3773
rect 8716 3717 8744 3773
rect 8800 3717 8828 3773
rect 8884 3717 8900 3773
rect 8300 3692 8900 3717
rect 8300 3636 8324 3692
rect 8380 3636 8408 3692
rect 8464 3636 8492 3692
rect 8548 3636 8576 3692
rect 8632 3636 8660 3692
rect 8716 3636 8744 3692
rect 8800 3636 8828 3692
rect 8884 3636 8900 3692
rect 8300 3611 8900 3636
rect 8300 3555 8324 3611
rect 8380 3555 8408 3611
rect 8464 3555 8492 3611
rect 8548 3555 8576 3611
rect 8632 3555 8660 3611
rect 8716 3555 8744 3611
rect 8800 3555 8828 3611
rect 8884 3555 8900 3611
rect 8300 3526 8900 3555
rect 9229 3526 9789 18029
rect 10114 17429 10806 18281
rect 10114 13046 10690 17429
tri 10690 17313 10806 17429 nw
rect 11030 18371 11590 18377
tri 12106 18376 12107 18377 se
rect 12107 18376 12490 18377
tri 12490 18376 12491 18377 sw
rect 11030 17347 11036 18371
rect 11580 17347 11590 18371
tri 12009 18279 12106 18376 se
rect 12106 18279 12491 18376
rect 11030 17330 11590 17347
rect 10114 12990 10122 13046
rect 10178 12990 10206 13046
rect 10262 12990 10290 13046
rect 10346 12990 10374 13046
rect 10430 12990 10458 13046
rect 10514 12990 10542 13046
rect 10598 12990 10626 13046
rect 10682 12990 10690 13046
rect 10114 12957 10690 12990
rect 10114 12901 10122 12957
rect 10178 12901 10206 12957
rect 10262 12901 10290 12957
rect 10346 12901 10374 12957
rect 10430 12901 10458 12957
rect 10514 12901 10542 12957
rect 10598 12901 10626 12957
rect 10682 12901 10690 12957
rect 10114 12868 10690 12901
rect 10114 12812 10122 12868
rect 10178 12812 10206 12868
rect 10262 12812 10290 12868
rect 10346 12812 10374 12868
rect 10430 12812 10458 12868
rect 10514 12812 10542 12868
rect 10598 12812 10626 12868
rect 10682 12812 10690 12868
rect 10114 12779 10690 12812
rect 10114 12723 10122 12779
rect 10178 12723 10206 12779
rect 10262 12723 10290 12779
rect 10346 12723 10374 12779
rect 10430 12723 10458 12779
rect 10514 12723 10542 12779
rect 10598 12723 10626 12779
rect 10682 12723 10690 12779
rect 10114 12690 10690 12723
rect 10114 12634 10122 12690
rect 10178 12634 10206 12690
rect 10262 12634 10290 12690
rect 10346 12634 10374 12690
rect 10430 12634 10458 12690
rect 10514 12634 10542 12690
rect 10598 12634 10626 12690
rect 10682 12634 10690 12690
rect 10114 12601 10690 12634
rect 10114 12545 10122 12601
rect 10178 12545 10206 12601
rect 10262 12545 10290 12601
rect 10346 12545 10374 12601
rect 10430 12545 10458 12601
rect 10514 12545 10542 12601
rect 10598 12545 10626 12601
rect 10682 12545 10690 12601
rect 10114 12511 10690 12545
rect 10114 12455 10122 12511
rect 10178 12455 10206 12511
rect 10262 12455 10290 12511
rect 10346 12455 10374 12511
rect 10430 12455 10458 12511
rect 10514 12455 10542 12511
rect 10598 12455 10626 12511
rect 10682 12455 10690 12511
rect 10114 12444 10690 12455
rect 11030 17266 11036 17330
rect 11100 17266 11116 17330
rect 11180 17266 11196 17330
rect 11260 17266 11276 17330
rect 11340 17266 11356 17330
rect 11420 17266 11436 17330
rect 11500 17266 11516 17330
rect 11580 17266 11590 17330
rect 11915 17286 12491 18279
tri 7082 2988 7270 3176 sw
tri 9931 2988 10116 3173 se
rect 10116 2988 10692 12080
rect 11030 3526 11590 17266
tri 12024 17143 12167 17286 ne
tri 12025 16436 12167 16578 se
rect 12167 16436 12491 17286
rect 11915 13046 12491 16436
rect 11915 12990 11923 13046
rect 11979 12990 12007 13046
rect 12063 12990 12091 13046
rect 12147 12990 12175 13046
rect 12231 12990 12259 13046
rect 12315 12990 12343 13046
rect 12399 12990 12427 13046
rect 12483 12990 12491 13046
rect 11915 12963 12491 12990
rect 11915 12907 11923 12963
rect 11979 12907 12007 12963
rect 12063 12907 12091 12963
rect 12147 12907 12175 12963
rect 12231 12907 12259 12963
rect 12315 12907 12343 12963
rect 12399 12907 12427 12963
rect 12483 12907 12491 12963
rect 11915 12880 12491 12907
rect 11915 12824 11923 12880
rect 11979 12824 12007 12880
rect 12063 12824 12091 12880
rect 12147 12824 12175 12880
rect 12231 12824 12259 12880
rect 12315 12824 12343 12880
rect 12399 12824 12427 12880
rect 12483 12824 12491 12880
rect 11915 12797 12491 12824
rect 11915 12741 11923 12797
rect 11979 12741 12007 12797
rect 12063 12741 12091 12797
rect 12147 12741 12175 12797
rect 12231 12741 12259 12797
rect 12315 12741 12343 12797
rect 12399 12741 12427 12797
rect 12483 12741 12491 12797
rect 11915 12713 12491 12741
rect 11915 12657 11923 12713
rect 11979 12657 12007 12713
rect 12063 12657 12091 12713
rect 12147 12657 12175 12713
rect 12231 12657 12259 12713
rect 12315 12657 12343 12713
rect 12399 12657 12427 12713
rect 12483 12657 12491 12713
rect 11915 12629 12491 12657
rect 11915 12573 11923 12629
rect 11979 12573 12007 12629
rect 12063 12573 12091 12629
rect 12147 12573 12175 12629
rect 12231 12573 12259 12629
rect 12315 12573 12343 12629
rect 12399 12573 12427 12629
rect 12483 12573 12491 12629
rect 11915 12545 12491 12573
rect 11915 12489 11923 12545
rect 11979 12489 12007 12545
rect 12063 12489 12091 12545
rect 12147 12489 12175 12545
rect 12231 12489 12259 12545
rect 12315 12489 12343 12545
rect 12399 12489 12427 12545
rect 12483 12489 12491 12545
rect 11915 12444 12491 12489
rect 12829 18371 13389 18377
rect 12829 17987 12837 18371
rect 13381 17987 13389 18371
rect 12829 17970 13389 17987
rect 12829 17906 12837 17970
rect 12901 17906 12917 17970
rect 12981 17906 12997 17970
rect 13061 17906 13077 17970
rect 13141 17906 13157 17970
rect 13221 17906 13237 17970
rect 13301 17906 13317 17970
rect 13381 17906 13389 17970
rect 12829 17889 13389 17906
rect 12829 17825 12837 17889
rect 12901 17825 12917 17889
rect 12981 17825 12997 17889
rect 13061 17825 13077 17889
rect 13141 17825 13157 17889
rect 13221 17825 13237 17889
rect 13301 17825 13317 17889
rect 13381 17825 13389 17889
rect 12829 17808 13389 17825
rect 12829 17744 12837 17808
rect 12901 17744 12917 17808
rect 12981 17744 12997 17808
rect 13061 17744 13077 17808
rect 13141 17744 13157 17808
rect 13221 17744 13237 17808
rect 13301 17744 13317 17808
rect 13381 17744 13389 17808
rect 12829 17727 13389 17744
rect 12829 17663 12837 17727
rect 12901 17663 12917 17727
rect 12981 17663 12997 17727
rect 13061 17663 13077 17727
rect 13141 17663 13157 17727
rect 13221 17663 13237 17727
rect 13301 17663 13317 17727
rect 13381 17663 13389 17727
rect 12829 17646 13389 17663
rect 12829 17582 12837 17646
rect 12901 17582 12917 17646
rect 12981 17582 12997 17646
rect 13061 17582 13077 17646
rect 13141 17582 13157 17646
rect 13221 17582 13237 17646
rect 13301 17582 13317 17646
rect 13381 17582 13389 17646
rect 12829 17565 13389 17582
rect 12829 17501 12837 17565
rect 12901 17501 12917 17565
rect 12981 17501 12997 17565
rect 13061 17501 13077 17565
rect 13141 17501 13157 17565
rect 13221 17501 13237 17565
rect 13301 17501 13317 17565
rect 13381 17501 13389 17565
rect 12829 17484 13389 17501
rect 12829 17420 12837 17484
rect 12901 17420 12917 17484
rect 12981 17420 12997 17484
rect 13061 17420 13077 17484
rect 13141 17420 13157 17484
rect 13221 17420 13237 17484
rect 13301 17420 13317 17484
rect 13381 17420 13389 17484
rect 12829 17403 13389 17420
rect 12829 17339 12837 17403
rect 12901 17339 12917 17403
rect 12981 17339 12997 17403
rect 13061 17339 13077 17403
rect 13141 17339 13157 17403
rect 13221 17339 13237 17403
rect 13301 17339 13317 17403
rect 13381 17339 13389 17403
rect 12829 17322 13389 17339
rect 12829 17258 12837 17322
rect 12901 17258 12917 17322
rect 12981 17258 12997 17322
rect 13061 17258 13077 17322
rect 13141 17258 13157 17322
rect 13221 17258 13237 17322
rect 13301 17258 13317 17322
rect 13381 17258 13389 17322
rect 12829 17241 13389 17258
rect 12829 17177 12837 17241
rect 12901 17177 12917 17241
rect 12981 17177 12997 17241
rect 13061 17177 13077 17241
rect 13141 17177 13157 17241
rect 13221 17177 13237 17241
rect 13301 17177 13317 17241
rect 13381 17177 13389 17241
rect 12829 17160 13389 17177
rect 12829 17096 12837 17160
rect 12901 17096 12917 17160
rect 12981 17096 12997 17160
rect 13061 17096 13077 17160
rect 13141 17096 13157 17160
rect 13221 17096 13237 17160
rect 13301 17096 13317 17160
rect 13381 17096 13389 17160
rect 12829 17079 13389 17096
rect 12829 17015 12837 17079
rect 12901 17015 12917 17079
rect 12981 17015 12997 17079
rect 13061 17015 13077 17079
rect 13141 17015 13157 17079
rect 13221 17015 13237 17079
rect 13301 17015 13317 17079
rect 13381 17015 13389 17079
rect 12829 16998 13389 17015
rect 12829 16934 12837 16998
rect 12901 16934 12917 16998
rect 12981 16934 12997 16998
rect 13061 16934 13077 16998
rect 13141 16934 13157 16998
rect 13221 16934 13237 16998
rect 13301 16934 13317 16998
rect 13381 16934 13389 16998
tri 10692 2988 10880 3176 sw
tri 11734 2988 11919 3173 se
rect 11919 2988 12495 12153
rect 12829 3526 13389 16934
tri 12495 2988 12683 3176 sw
tri 13522 2988 13671 3137 se
rect 13671 2988 14287 11850
tri 14287 2988 14436 3137 sw
rect -4308 2948 14287 2988
rect -4308 -800 13671 2948
rect 13721 1151 14287 2897
<< via3 >>
rect 217 18381 281 18445
rect 313 18381 377 18445
rect 409 18381 473 18445
rect 505 18381 569 18445
rect 601 18381 665 18445
rect 696 18381 760 18445
rect 217 18293 281 18357
rect 313 18293 377 18357
rect 409 18293 473 18357
rect 505 18293 569 18357
rect 601 18293 665 18357
rect 696 18293 760 18357
rect 217 18205 281 18269
rect 313 18205 377 18269
rect 409 18205 473 18269
rect 505 18205 569 18269
rect 601 18205 665 18269
rect 696 18205 760 18269
rect 217 18117 281 18181
rect 313 18117 377 18181
rect 409 18117 473 18181
rect 505 18117 569 18181
rect 601 18117 665 18181
rect 696 18117 760 18181
rect 217 18029 281 18093
rect 313 18029 377 18093
rect 409 18029 473 18093
rect 505 18029 569 18093
rect 601 18029 665 18093
rect 696 18029 760 18093
rect 2024 18381 2088 18445
rect 2120 18381 2184 18445
rect 2216 18381 2280 18445
rect 2312 18381 2376 18445
rect 2408 18381 2472 18445
rect 2503 18381 2567 18445
rect 2024 18293 2088 18357
rect 2120 18293 2184 18357
rect 2216 18293 2280 18357
rect 2312 18293 2376 18357
rect 2408 18293 2472 18357
rect 2503 18293 2567 18357
rect 2024 18205 2088 18269
rect 2120 18205 2184 18269
rect 2216 18205 2280 18269
rect 2312 18205 2376 18269
rect 2408 18205 2472 18269
rect 2503 18205 2567 18269
rect 2024 18117 2088 18181
rect 2120 18117 2184 18181
rect 2216 18117 2280 18181
rect 2312 18117 2376 18181
rect 2408 18117 2472 18181
rect 2503 18117 2567 18181
rect 2024 18029 2088 18093
rect 2120 18029 2184 18093
rect 2216 18029 2280 18093
rect 2312 18029 2376 18093
rect 2408 18029 2472 18093
rect 2503 18029 2567 18093
rect 3819 18381 3883 18445
rect 3915 18381 3979 18445
rect 4011 18381 4075 18445
rect 4107 18381 4171 18445
rect 4203 18381 4267 18445
rect 4298 18381 4362 18445
rect 3819 18293 3883 18357
rect 3915 18293 3979 18357
rect 4011 18293 4075 18357
rect 4107 18293 4171 18357
rect 4203 18293 4267 18357
rect 4298 18293 4362 18357
rect 3819 18205 3883 18269
rect 3915 18205 3979 18269
rect 4011 18205 4075 18269
rect 4107 18205 4171 18269
rect 4203 18205 4267 18269
rect 4298 18205 4362 18269
rect 3819 18117 3883 18181
rect 3915 18117 3979 18181
rect 4011 18117 4075 18181
rect 4107 18117 4171 18181
rect 4203 18117 4267 18181
rect 4298 18117 4362 18181
rect 3819 18029 3883 18093
rect 3915 18029 3979 18093
rect 4011 18029 4075 18093
rect 4107 18029 4171 18093
rect 4203 18029 4267 18093
rect 4298 18029 4362 18093
rect 5629 18381 5693 18445
rect 5725 18381 5789 18445
rect 5821 18381 5885 18445
rect 5917 18381 5981 18445
rect 6013 18381 6077 18445
rect 6108 18381 6172 18445
rect 5629 18293 5693 18357
rect 5725 18293 5789 18357
rect 5821 18293 5885 18357
rect 5917 18293 5981 18357
rect 6013 18293 6077 18357
rect 6108 18293 6172 18357
rect 5629 18205 5693 18269
rect 5725 18205 5789 18269
rect 5821 18205 5885 18269
rect 5917 18205 5981 18269
rect 6013 18205 6077 18269
rect 6108 18205 6172 18269
rect 5629 18117 5693 18181
rect 5725 18117 5789 18181
rect 5821 18117 5885 18181
rect 5917 18117 5981 18181
rect 6013 18117 6077 18181
rect 6108 18117 6172 18181
rect 5629 18029 5693 18093
rect 5725 18029 5789 18093
rect 5821 18029 5885 18093
rect 5917 18029 5981 18093
rect 6013 18029 6077 18093
rect 6108 18029 6172 18093
rect 7427 18381 7491 18445
rect 7523 18381 7587 18445
rect 7619 18381 7683 18445
rect 7715 18381 7779 18445
rect 7811 18381 7875 18445
rect 7906 18381 7970 18445
rect 7427 18293 7491 18357
rect 7523 18293 7587 18357
rect 7619 18293 7683 18357
rect 7715 18293 7779 18357
rect 7811 18293 7875 18357
rect 7906 18293 7970 18357
rect 7427 18205 7491 18269
rect 7523 18205 7587 18269
rect 7619 18205 7683 18269
rect 7715 18205 7779 18269
rect 7811 18205 7875 18269
rect 7906 18205 7970 18269
rect 9237 18381 9301 18445
rect 9333 18381 9397 18445
rect 9429 18381 9493 18445
rect 9525 18381 9589 18445
rect 9621 18381 9685 18445
rect 9716 18381 9780 18445
rect 9237 18293 9301 18357
rect 9333 18293 9397 18357
rect 9429 18293 9493 18357
rect 9525 18293 9589 18357
rect 9621 18293 9685 18357
rect 9716 18293 9780 18357
rect 7427 18117 7491 18181
rect 7523 18117 7587 18181
rect 7619 18117 7683 18181
rect 7715 18117 7779 18181
rect 7811 18117 7875 18181
rect 7906 18117 7970 18181
rect 9237 18205 9301 18269
rect 9333 18205 9397 18269
rect 9429 18205 9493 18269
rect 9525 18205 9589 18269
rect 9621 18205 9685 18269
rect 9716 18205 9780 18269
rect 9237 18117 9301 18181
rect 9333 18117 9397 18181
rect 9429 18117 9493 18181
rect 9525 18117 9589 18181
rect 9621 18117 9685 18181
rect 9716 18117 9780 18181
rect 7427 18029 7491 18093
rect 7523 18029 7587 18093
rect 7619 18029 7683 18093
rect 7715 18029 7779 18093
rect 7811 18029 7875 18093
rect 7906 18029 7970 18093
rect 9237 18029 9301 18093
rect 9333 18029 9397 18093
rect 9429 18029 9493 18093
rect 9525 18029 9589 18093
rect 9621 18029 9685 18093
rect 9716 18029 9780 18093
rect 11036 17347 11580 18371
rect 11036 17266 11100 17330
rect 11116 17266 11180 17330
rect 11196 17266 11260 17330
rect 11276 17266 11340 17330
rect 11356 17266 11420 17330
rect 11436 17266 11500 17330
rect 11516 17266 11580 17330
rect 12837 17987 13381 18371
rect 12837 17906 12901 17970
rect 12917 17906 12981 17970
rect 12997 17906 13061 17970
rect 13077 17906 13141 17970
rect 13157 17906 13221 17970
rect 13237 17906 13301 17970
rect 13317 17906 13381 17970
rect 12837 17825 12901 17889
rect 12917 17825 12981 17889
rect 12997 17825 13061 17889
rect 13077 17825 13141 17889
rect 13157 17825 13221 17889
rect 13237 17825 13301 17889
rect 13317 17825 13381 17889
rect 12837 17744 12901 17808
rect 12917 17744 12981 17808
rect 12997 17744 13061 17808
rect 13077 17744 13141 17808
rect 13157 17744 13221 17808
rect 13237 17744 13301 17808
rect 13317 17744 13381 17808
rect 12837 17663 12901 17727
rect 12917 17663 12981 17727
rect 12997 17663 13061 17727
rect 13077 17663 13141 17727
rect 13157 17663 13221 17727
rect 13237 17663 13301 17727
rect 13317 17663 13381 17727
rect 12837 17582 12901 17646
rect 12917 17582 12981 17646
rect 12997 17582 13061 17646
rect 13077 17582 13141 17646
rect 13157 17582 13221 17646
rect 13237 17582 13301 17646
rect 13317 17582 13381 17646
rect 12837 17501 12901 17565
rect 12917 17501 12981 17565
rect 12997 17501 13061 17565
rect 13077 17501 13141 17565
rect 13157 17501 13221 17565
rect 13237 17501 13301 17565
rect 13317 17501 13381 17565
rect 12837 17420 12901 17484
rect 12917 17420 12981 17484
rect 12997 17420 13061 17484
rect 13077 17420 13141 17484
rect 13157 17420 13221 17484
rect 13237 17420 13301 17484
rect 13317 17420 13381 17484
rect 12837 17339 12901 17403
rect 12917 17339 12981 17403
rect 12997 17339 13061 17403
rect 13077 17339 13141 17403
rect 13157 17339 13221 17403
rect 13237 17339 13301 17403
rect 13317 17339 13381 17403
rect 12837 17258 12901 17322
rect 12917 17258 12981 17322
rect 12997 17258 13061 17322
rect 13077 17258 13141 17322
rect 13157 17258 13221 17322
rect 13237 17258 13301 17322
rect 13317 17258 13381 17322
rect 12837 17177 12901 17241
rect 12917 17177 12981 17241
rect 12997 17177 13061 17241
rect 13077 17177 13141 17241
rect 13157 17177 13221 17241
rect 13237 17177 13301 17241
rect 13317 17177 13381 17241
rect 12837 17096 12901 17160
rect 12917 17096 12981 17160
rect 12997 17096 13061 17160
rect 13077 17096 13141 17160
rect 13157 17096 13221 17160
rect 13237 17096 13301 17160
rect 13317 17096 13381 17160
rect 12837 17015 12901 17079
rect 12917 17015 12981 17079
rect 12997 17015 13061 17079
rect 13077 17015 13141 17079
rect 13157 17015 13221 17079
rect 13237 17015 13301 17079
rect 13317 17015 13381 17079
rect 12837 16934 12901 16998
rect 12917 16934 12981 16998
rect 12997 16934 13061 16998
rect 13077 16934 13141 16998
rect 13157 16934 13221 16998
rect 13237 16934 13301 16998
rect 13317 16934 13381 16998
<< metal4 >>
rect 216 18445 761 18446
rect 216 18381 217 18445
rect 281 18381 313 18445
rect 377 18381 409 18445
rect 473 18381 505 18445
rect 569 18381 601 18445
rect 665 18381 696 18445
rect 760 18381 761 18445
rect 216 18357 761 18381
rect 216 18293 217 18357
rect 281 18293 313 18357
rect 377 18293 409 18357
rect 473 18293 505 18357
rect 569 18293 601 18357
rect 665 18293 696 18357
rect 760 18293 761 18357
rect 216 18269 761 18293
rect 216 18205 217 18269
rect 281 18205 313 18269
rect 377 18205 409 18269
rect 473 18205 505 18269
rect 569 18205 601 18269
rect 665 18205 696 18269
rect 760 18205 761 18269
rect 216 18181 761 18205
rect 216 18117 217 18181
rect 281 18117 313 18181
rect 377 18117 409 18181
rect 473 18117 505 18181
rect 569 18117 601 18181
rect 665 18117 696 18181
rect 760 18117 761 18181
rect 216 18093 761 18117
rect 216 18029 217 18093
rect 281 18029 313 18093
rect 377 18029 409 18093
rect 473 18029 505 18093
rect 569 18029 601 18093
rect 665 18029 696 18093
rect 760 18029 761 18093
rect 216 18028 761 18029
rect 2023 18445 2568 18446
rect 2023 18381 2024 18445
rect 2088 18381 2120 18445
rect 2184 18381 2216 18445
rect 2280 18381 2312 18445
rect 2376 18381 2408 18445
rect 2472 18381 2503 18445
rect 2567 18381 2568 18445
rect 2023 18357 2568 18381
rect 2023 18293 2024 18357
rect 2088 18293 2120 18357
rect 2184 18293 2216 18357
rect 2280 18293 2312 18357
rect 2376 18293 2408 18357
rect 2472 18293 2503 18357
rect 2567 18293 2568 18357
rect 2023 18269 2568 18293
rect 2023 18205 2024 18269
rect 2088 18205 2120 18269
rect 2184 18205 2216 18269
rect 2280 18205 2312 18269
rect 2376 18205 2408 18269
rect 2472 18205 2503 18269
rect 2567 18205 2568 18269
rect 2023 18181 2568 18205
rect 2023 18117 2024 18181
rect 2088 18117 2120 18181
rect 2184 18117 2216 18181
rect 2280 18117 2312 18181
rect 2376 18117 2408 18181
rect 2472 18117 2503 18181
rect 2567 18117 2568 18181
rect 2023 18093 2568 18117
rect 2023 18029 2024 18093
rect 2088 18029 2120 18093
rect 2184 18029 2216 18093
rect 2280 18029 2312 18093
rect 2376 18029 2408 18093
rect 2472 18029 2503 18093
rect 2567 18029 2568 18093
rect 2023 18028 2568 18029
rect 3818 18445 4363 18446
rect 3818 18381 3819 18445
rect 3883 18381 3915 18445
rect 3979 18381 4011 18445
rect 4075 18381 4107 18445
rect 4171 18381 4203 18445
rect 4267 18381 4298 18445
rect 4362 18381 4363 18445
rect 3818 18357 4363 18381
rect 3818 18293 3819 18357
rect 3883 18293 3915 18357
rect 3979 18293 4011 18357
rect 4075 18293 4107 18357
rect 4171 18293 4203 18357
rect 4267 18293 4298 18357
rect 4362 18293 4363 18357
rect 3818 18269 4363 18293
rect 3818 18205 3819 18269
rect 3883 18205 3915 18269
rect 3979 18205 4011 18269
rect 4075 18205 4107 18269
rect 4171 18205 4203 18269
rect 4267 18205 4298 18269
rect 4362 18205 4363 18269
rect 3818 18181 4363 18205
rect 3818 18117 3819 18181
rect 3883 18117 3915 18181
rect 3979 18117 4011 18181
rect 4075 18117 4107 18181
rect 4171 18117 4203 18181
rect 4267 18117 4298 18181
rect 4362 18117 4363 18181
rect 3818 18093 4363 18117
rect 3818 18029 3819 18093
rect 3883 18029 3915 18093
rect 3979 18029 4011 18093
rect 4075 18029 4107 18093
rect 4171 18029 4203 18093
rect 4267 18029 4298 18093
rect 4362 18029 4363 18093
rect 3818 18028 4363 18029
rect 5628 18445 6173 18446
rect 5628 18381 5629 18445
rect 5693 18381 5725 18445
rect 5789 18381 5821 18445
rect 5885 18381 5917 18445
rect 5981 18381 6013 18445
rect 6077 18381 6108 18445
rect 6172 18381 6173 18445
rect 5628 18357 6173 18381
rect 5628 18293 5629 18357
rect 5693 18293 5725 18357
rect 5789 18293 5821 18357
rect 5885 18293 5917 18357
rect 5981 18293 6013 18357
rect 6077 18293 6108 18357
rect 6172 18293 6173 18357
rect 5628 18269 6173 18293
rect 5628 18205 5629 18269
rect 5693 18205 5725 18269
rect 5789 18205 5821 18269
rect 5885 18205 5917 18269
rect 5981 18205 6013 18269
rect 6077 18205 6108 18269
rect 6172 18205 6173 18269
rect 5628 18181 6173 18205
rect 5628 18117 5629 18181
rect 5693 18117 5725 18181
rect 5789 18117 5821 18181
rect 5885 18117 5917 18181
rect 5981 18117 6013 18181
rect 6077 18117 6108 18181
rect 6172 18117 6173 18181
rect 5628 18093 6173 18117
rect 5628 18029 5629 18093
rect 5693 18029 5725 18093
rect 5789 18029 5821 18093
rect 5885 18029 5917 18093
rect 5981 18029 6013 18093
rect 6077 18029 6108 18093
rect 6172 18029 6173 18093
rect 5628 18028 6173 18029
rect 7426 18445 7971 18446
rect 7426 18381 7427 18445
rect 7491 18381 7523 18445
rect 7587 18381 7619 18445
rect 7683 18381 7715 18445
rect 7779 18381 7811 18445
rect 7875 18381 7906 18445
rect 7970 18381 7971 18445
rect 7426 18357 7971 18381
rect 7426 18293 7427 18357
rect 7491 18293 7523 18357
rect 7587 18293 7619 18357
rect 7683 18293 7715 18357
rect 7779 18293 7811 18357
rect 7875 18293 7906 18357
rect 7970 18293 7971 18357
rect 7426 18269 7971 18293
rect 7426 18205 7427 18269
rect 7491 18205 7523 18269
rect 7587 18205 7619 18269
rect 7683 18205 7715 18269
rect 7779 18205 7811 18269
rect 7875 18205 7906 18269
rect 7970 18205 7971 18269
rect 7426 18181 7971 18205
rect 7426 18117 7427 18181
rect 7491 18117 7523 18181
rect 7587 18117 7619 18181
rect 7683 18117 7715 18181
rect 7779 18117 7811 18181
rect 7875 18117 7906 18181
rect 7970 18117 7971 18181
rect 7426 18093 7971 18117
rect 7426 18029 7427 18093
rect 7491 18029 7523 18093
rect 7587 18029 7619 18093
rect 7683 18029 7715 18093
rect 7779 18029 7811 18093
rect 7875 18029 7906 18093
rect 7970 18029 7971 18093
rect 7426 18028 7971 18029
rect 9236 18445 9781 18446
rect 9236 18381 9237 18445
rect 9301 18381 9333 18445
rect 9397 18381 9429 18445
rect 9493 18381 9525 18445
rect 9589 18381 9621 18445
rect 9685 18381 9716 18445
rect 9780 18381 9781 18445
rect 9236 18357 9781 18381
rect 9236 18293 9237 18357
rect 9301 18293 9333 18357
rect 9397 18293 9429 18357
rect 9493 18293 9525 18357
rect 9589 18293 9621 18357
rect 9685 18293 9716 18357
rect 9780 18293 9781 18357
rect 9236 18269 9781 18293
rect 9236 18205 9237 18269
rect 9301 18205 9333 18269
rect 9397 18205 9429 18269
rect 9493 18205 9525 18269
rect 9589 18205 9621 18269
rect 9685 18205 9716 18269
rect 9780 18205 9781 18269
rect 9236 18181 9781 18205
rect 9236 18117 9237 18181
rect 9301 18117 9333 18181
rect 9397 18117 9429 18181
rect 9493 18117 9525 18181
rect 9589 18117 9621 18181
rect 9685 18117 9716 18181
rect 9780 18117 9781 18181
rect 9236 18093 9781 18117
rect 9236 18029 9237 18093
rect 9301 18029 9333 18093
rect 9397 18029 9429 18093
rect 9493 18029 9525 18093
rect 9589 18029 9621 18093
rect 9685 18029 9716 18093
rect 9780 18029 9781 18093
rect 9236 18028 9781 18029
rect 11035 18371 11581 18372
rect 11035 17347 11036 18371
rect 11580 17347 11581 18371
rect 11035 17330 11581 17347
rect 11035 17266 11036 17330
rect 11100 17266 11116 17330
rect 11180 17266 11196 17330
rect 11260 17266 11276 17330
rect 11340 17266 11356 17330
rect 11420 17266 11436 17330
rect 11500 17266 11516 17330
rect 11580 17266 11581 17330
rect 11035 17265 11581 17266
rect 12836 18371 13382 18372
rect 12836 17987 12837 18371
rect 13381 17987 13382 18371
rect 12836 17970 13382 17987
rect 12836 17906 12837 17970
rect 12901 17906 12917 17970
rect 12981 17906 12997 17970
rect 13061 17906 13077 17970
rect 13141 17906 13157 17970
rect 13221 17906 13237 17970
rect 13301 17906 13317 17970
rect 13381 17906 13382 17970
rect 12836 17889 13382 17906
rect 12836 17825 12837 17889
rect 12901 17825 12917 17889
rect 12981 17825 12997 17889
rect 13061 17825 13077 17889
rect 13141 17825 13157 17889
rect 13221 17825 13237 17889
rect 13301 17825 13317 17889
rect 13381 17825 13382 17889
rect 12836 17808 13382 17825
rect 12836 17744 12837 17808
rect 12901 17744 12917 17808
rect 12981 17744 12997 17808
rect 13061 17744 13077 17808
rect 13141 17744 13157 17808
rect 13221 17744 13237 17808
rect 13301 17744 13317 17808
rect 13381 17744 13382 17808
rect 12836 17727 13382 17744
rect 12836 17663 12837 17727
rect 12901 17663 12917 17727
rect 12981 17663 12997 17727
rect 13061 17663 13077 17727
rect 13141 17663 13157 17727
rect 13221 17663 13237 17727
rect 13301 17663 13317 17727
rect 13381 17663 13382 17727
rect 12836 17646 13382 17663
rect 12836 17582 12837 17646
rect 12901 17582 12917 17646
rect 12981 17582 12997 17646
rect 13061 17582 13077 17646
rect 13141 17582 13157 17646
rect 13221 17582 13237 17646
rect 13301 17582 13317 17646
rect 13381 17582 13382 17646
rect 12836 17565 13382 17582
rect 12836 17501 12837 17565
rect 12901 17501 12917 17565
rect 12981 17501 12997 17565
rect 13061 17501 13077 17565
rect 13141 17501 13157 17565
rect 13221 17501 13237 17565
rect 13301 17501 13317 17565
rect 13381 17501 13382 17565
rect 12836 17484 13382 17501
rect 12836 17420 12837 17484
rect 12901 17420 12917 17484
rect 12981 17420 12997 17484
rect 13061 17420 13077 17484
rect 13141 17420 13157 17484
rect 13221 17420 13237 17484
rect 13301 17420 13317 17484
rect 13381 17420 13382 17484
rect 12836 17403 13382 17420
rect 12836 17339 12837 17403
rect 12901 17339 12917 17403
rect 12981 17339 12997 17403
rect 13061 17339 13077 17403
rect 13141 17339 13157 17403
rect 13221 17339 13237 17403
rect 13301 17339 13317 17403
rect 13381 17339 13382 17403
rect 12836 17322 13382 17339
rect 12836 17258 12837 17322
rect 12901 17258 12917 17322
rect 12981 17258 12997 17322
rect 13061 17258 13077 17322
rect 13141 17258 13157 17322
rect 13221 17258 13237 17322
rect 13301 17258 13317 17322
rect 13381 17258 13382 17322
rect 12836 17241 13382 17258
rect 12836 17177 12837 17241
rect 12901 17177 12917 17241
rect 12981 17177 12997 17241
rect 13061 17177 13077 17241
rect 13141 17177 13157 17241
rect 13221 17177 13237 17241
rect 13301 17177 13317 17241
rect 13381 17177 13382 17241
rect 12836 17160 13382 17177
rect 12836 17096 12837 17160
rect 12901 17096 12917 17160
rect 12981 17096 12997 17160
rect 13061 17096 13077 17160
rect 13141 17096 13157 17160
rect 13221 17096 13237 17160
rect 13301 17096 13317 17160
rect 13381 17096 13382 17160
rect 12836 17079 13382 17096
rect 12836 17015 12837 17079
rect 12901 17015 12917 17079
rect 12981 17015 12997 17079
rect 13061 17015 13077 17079
rect 13141 17015 13157 17079
rect 13221 17015 13237 17079
rect 13301 17015 13317 17079
rect 13381 17015 13382 17079
rect 12836 16998 13382 17015
rect 12836 16934 12837 16998
rect 12901 16934 12917 16998
rect 12981 16934 12997 16998
rect 13061 16934 13077 16998
rect 13141 16934 13157 16998
rect 13221 16934 13237 16998
rect 13301 16934 13317 16998
rect 13381 16934 13382 16998
rect 12836 16933 13382 16934
tri -1772 5018 -1278 5512 se
rect -1278 5018 -738 5512
tri -1812 4978 -1772 5018 se
rect -1772 4978 -738 5018
tri 11222 4978 11262 5018 se
rect 11262 4978 11676 5615
tri -2028 4762 -1812 4978 se
rect -1812 4762 -738 4978
rect -3406 3997 -738 4762
tri -738 3997 243 4978 sw
tri 10241 3997 11222 4978 se
rect 11222 3997 11676 4978
tri 11676 3997 12785 5106 sw
rect -3406 3531 12936 3997
rect 12970 3669 13251 3813
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1707688321
transform 0 1 3129 1 0 770
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_1
timestamp 1707688321
transform 0 -1 1093 1 0 770
box 0 0 1 1
use M1M2_CDNS_52468879185967  M1M2_CDNS_52468879185967_0
timestamp 1707688321
transform -1 0 14173 0 -1 613
box 0 0 448 116
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_0
timestamp 1707688321
transform 1 0 -4109 0 1 11991
box 0 0 320 180
use M1M2_CDNS_524688791851177  M1M2_CDNS_524688791851177_0
timestamp 1707688321
transform 1 0 86 0 -1 12973
box 0 0 384 116
use M1M2_CDNS_524688791851177  M1M2_CDNS_524688791851177_1
timestamp 1707688321
transform 1 0 14530 0 -1 12973
box 0 0 384 116
use M1M2_CDNS_524688791851513  M1M2_CDNS_524688791851513_0
timestamp 1707688321
transform 1 0 2898 0 1 11680
box 0 0 576 436
use M1M2_CDNS_524688791851513  M1M2_CDNS_524688791851513_1
timestamp 1707688321
transform 1 0 1094 0 1 11680
box 0 0 576 436
use M1M2_CDNS_524688791851513  M1M2_CDNS_524688791851513_2
timestamp 1707688321
transform 1 0 4699 0 1 11680
box 0 0 576 436
use M1M2_CDNS_524688791851513  M1M2_CDNS_524688791851513_3
timestamp 1707688321
transform 1 0 6506 0 1 11680
box 0 0 576 436
use M1M2_CDNS_524688791851513  M1M2_CDNS_524688791851513_4
timestamp 1707688321
transform 1 0 10116 0 1 11680
box 0 0 576 436
use M1M2_CDNS_524688791851514  M1M2_CDNS_524688791851514_0
timestamp 1707688321
transform 1 0 6506 0 1 5210
box 0 0 576 6132
use M1M2_CDNS_524688791851514  M1M2_CDNS_524688791851514_1
timestamp 1707688321
transform 1 0 2898 0 1 5210
box 0 0 576 6132
use M1M2_CDNS_524688791851514  M1M2_CDNS_524688791851514_2
timestamp 1707688321
transform 1 0 5607 0 1 5210
box 0 0 576 6132
use M1M2_CDNS_524688791851514  M1M2_CDNS_524688791851514_3
timestamp 1707688321
transform 1 0 195 0 1 5210
box 0 0 576 6132
use M1M2_CDNS_524688791851514  M1M2_CDNS_524688791851514_4
timestamp 1707688321
transform 1 0 3803 0 1 5210
box 0 0 576 6132
use M1M2_CDNS_524688791851514  M1M2_CDNS_524688791851514_5
timestamp 1707688321
transform 1 0 1999 0 1 5210
box 0 0 576 6132
use M1M2_CDNS_524688791851514  M1M2_CDNS_524688791851514_6
timestamp 1707688321
transform 1 0 1094 0 1 5210
box 0 0 576 6132
use M1M2_CDNS_524688791851514  M1M2_CDNS_524688791851514_7
timestamp 1707688321
transform 1 0 4699 0 1 5210
box 0 0 576 6132
use M1M2_CDNS_524688791851514  M1M2_CDNS_524688791851514_8
timestamp 1707688321
transform 1 0 10116 0 1 5210
box 0 0 576 6132
use M1M2_CDNS_524688791851514  M1M2_CDNS_524688791851514_9
timestamp 1707688321
transform 1 0 7410 0 1 5210
box 0 0 576 6132
use M1M2_CDNS_524688791851514  M1M2_CDNS_524688791851514_10
timestamp 1707688321
transform 1 0 9212 0 1 5210
box 0 0 576 6132
use M1M2_CDNS_524688791851514  M1M2_CDNS_524688791851514_11
timestamp 1707688321
transform 1 0 11021 0 1 5210
box 0 0 576 6132
use M1M2_CDNS_524688791851515  M1M2_CDNS_524688791851515_0
timestamp 1707688321
transform 1 0 -1567 0 -1 4739
box 0 0 512 1204
use M1M2_CDNS_524688791851516  M1M2_CDNS_524688791851516_0
timestamp 1707688321
transform 1 0 -3416 0 -1 4739
box 0 0 576 1204
use M1M2_CDNS_524688791851517  M1M2_CDNS_524688791851517_0
timestamp 1707688321
transform 1 0 -3731 0 1 11681
box 0 0 1792 500
use M1M2_CDNS_524688791851518  M1M2_CDNS_524688791851518_0
timestamp 1707688321
transform 1 0 -4311 0 1 5139
box 0 0 576 6836
use M1M2_CDNS_524688791851519  M1M2_CDNS_524688791851519_0
timestamp 1707688321
transform 1 0 12825 0 1 5139
box 0 0 576 6196
use M1M2_CDNS_524688791851519  M1M2_CDNS_524688791851519_1
timestamp 1707688321
transform 1 0 -1617 0 1 5139
box 0 0 576 6196
use M1M2_CDNS_524688791851519  M1M2_CDNS_524688791851519_2
timestamp 1707688321
transform 1 0 -2515 0 1 5139
box 0 0 576 6196
use M1M2_CDNS_524688791851519  M1M2_CDNS_524688791851519_3
timestamp 1707688321
transform 1 0 11919 0 1 5139
box 0 0 576 6196
use M1M2_CDNS_524688791851520  M1M2_CDNS_524688791851520_0
timestamp 1707688321
transform 1 0 13722 0 1 5139
box 0 0 576 6772
use M1M2_CDNS_524688791851521  M1M2_CDNS_524688791851521_0
timestamp 1707688321
transform -1 0 1682 0 -1 613
box 0 0 576 116
use M1M2_CDNS_524688791851521  M1M2_CDNS_524688791851521_1
timestamp 1707688321
transform -1 0 10690 0 -1 613
box 0 0 576 116
use M1M2_CDNS_524688791851521  M1M2_CDNS_524688791851521_2
timestamp 1707688321
transform -1 0 8886 0 -1 613
box 0 0 576 116
use M1M2_CDNS_524688791851521  M1M2_CDNS_524688791851521_3
timestamp 1707688321
transform -1 0 7082 0 -1 613
box 0 0 576 116
use M1M2_CDNS_524688791851521  M1M2_CDNS_524688791851521_4
timestamp 1707688321
transform -1 0 12495 0 -1 613
box 0 0 576 116
use M1M2_CDNS_524688791851521  M1M2_CDNS_524688791851521_5
timestamp 1707688321
transform -1 0 -134 0 -1 613
box 0 0 576 116
use M1M2_CDNS_524688791851521  M1M2_CDNS_524688791851521_6
timestamp 1707688321
transform -1 0 -3743 0 -1 613
box 0 0 576 116
use M1M2_CDNS_524688791851521  M1M2_CDNS_524688791851521_7
timestamp 1707688321
transform -1 0 -1942 0 -1 613
box 0 0 576 116
use M1M2_CDNS_524688791851521  M1M2_CDNS_524688791851521_8
timestamp 1707688321
transform -1 0 5266 0 -1 613
box 0 0 576 116
use M1M2_CDNS_524688791851521  M1M2_CDNS_524688791851521_9
timestamp 1707688321
transform -1 0 3476 0 -1 613
box 0 0 576 116
use M1M2_CDNS_524688791851522  M1M2_CDNS_524688791851522_0
timestamp 1707688321
transform 1 0 9218 0 -1 4009
box 0 0 576 500
use M1M2_CDNS_524688791851522  M1M2_CDNS_524688791851522_1
timestamp 1707688321
transform 1 0 7408 0 -1 4009
box 0 0 576 500
use M1M2_CDNS_524688791851522  M1M2_CDNS_524688791851522_2
timestamp 1707688321
transform 1 0 198 0 -1 4009
box 0 0 576 500
use M1M2_CDNS_524688791851522  M1M2_CDNS_524688791851522_3
timestamp 1707688321
transform 1 0 3800 0 -1 4009
box 0 0 576 500
use M1M2_CDNS_524688791851522  M1M2_CDNS_524688791851522_4
timestamp 1707688321
transform 1 0 5607 0 -1 4009
box 0 0 576 500
use M1M2_CDNS_524688791851522  M1M2_CDNS_524688791851522_5
timestamp 1707688321
transform 1 0 11019 0 -1 4009
box 0 0 576 500
use M1M2_CDNS_524688791851522  M1M2_CDNS_524688791851522_6
timestamp 1707688321
transform 1 0 12818 0 -1 4009
box 0 0 576 500
use M1M2_CDNS_524688791851522  M1M2_CDNS_524688791851522_7
timestamp 1707688321
transform 1 0 2000 0 -1 4009
box 0 0 576 500
use M1M2_CDNS_524688791851522  M1M2_CDNS_524688791851522_8
timestamp 1707688321
transform 1 0 11919 0 1 11680
box 0 0 576 500
use M1M2_CDNS_524688791851523  M1M2_CDNS_524688791851523_0
timestamp 1707688321
transform 1 0 -4318 0 1 1135
box 0 0 576 1780
use M1M2_CDNS_524688791851523  M1M2_CDNS_524688791851523_1
timestamp 1707688321
transform 1 0 -2514 0 1 1135
box 0 0 576 1780
use M1M2_CDNS_524688791851523  M1M2_CDNS_524688791851523_2
timestamp 1707688321
transform 1 0 -710 0 1 1135
box 0 0 576 1780
use M1M2_CDNS_524688791851523  M1M2_CDNS_524688791851523_3
timestamp 1707688321
transform 1 0 1094 0 1 1135
box 0 0 576 1780
use M1M2_CDNS_524688791851523  M1M2_CDNS_524688791851523_4
timestamp 1707688321
transform 1 0 2898 0 1 1135
box 0 0 576 1780
use M1M2_CDNS_524688791851523  M1M2_CDNS_524688791851523_5
timestamp 1707688321
transform 1 0 10114 0 1 1135
box 0 0 576 1780
use M1M2_CDNS_524688791851523  M1M2_CDNS_524688791851523_6
timestamp 1707688321
transform 1 0 6506 0 1 1135
box 0 0 576 1780
use M1M2_CDNS_524688791851523  M1M2_CDNS_524688791851523_7
timestamp 1707688321
transform 1 0 13722 0 1 1135
box 0 0 576 1780
use M1M2_CDNS_524688791851523  M1M2_CDNS_524688791851523_8
timestamp 1707688321
transform 1 0 4696 0 1 1135
box 0 0 576 1780
use M1M2_CDNS_524688791851523  M1M2_CDNS_524688791851523_9
timestamp 1707688321
transform 1 0 8310 0 1 1135
box 0 0 576 1780
use M1M2_CDNS_524688791851523  M1M2_CDNS_524688791851523_10
timestamp 1707688321
transform 1 0 11918 0 1 1135
box 0 0 576 1780
use M1M2_CDNS_524688791851524  M1M2_CDNS_524688791851524_0
timestamp 1707688321
transform 0 1 14942 -1 0 12825
box 0 0 8704 116
use M2M3_CDNS_524688791851525  M2M3_CDNS_524688791851525_0
timestamp 1707688321
transform 1 0 2917 0 1 5210
box -5 0 541 6874
use M2M3_CDNS_524688791851525  M2M3_CDNS_524688791851525_1
timestamp 1707688321
transform 1 0 1113 0 1 5210
box -5 0 541 6874
use M2M3_CDNS_524688791851525  M2M3_CDNS_524688791851525_2
timestamp 1707688321
transform 1 0 4720 0 1 5210
box -5 0 541 6874
use M2M3_CDNS_524688791851525  M2M3_CDNS_524688791851525_3
timestamp 1707688321
transform 1 0 6528 0 1 5210
box -5 0 541 6874
use M2M3_CDNS_524688791851525  M2M3_CDNS_524688791851525_4
timestamp 1707688321
transform 1 0 10133 0 1 5210
box -5 0 541 6874
use M2M3_CDNS_524688791851526  M2M3_CDNS_524688791851526_0
timestamp 1707688321
transform 1 0 -4286 0 1 2915
box -5 0 541 9034
use M2M3_CDNS_524688791851527  M2M3_CDNS_524688791851527_0
timestamp 1707688321
transform 1 0 -2512 0 1 2915
box -5 0 381 8394
use M2M3_CDNS_524688791851528  M2M3_CDNS_524688791851528_0
timestamp 1707688321
transform 1 0 -3400 0 1 3535
box -5 0 541 1194
use M2M3_CDNS_524688791851528  M2M3_CDNS_524688791851528_1
timestamp 1707688321
transform 1 0 -1582 0 1 3535
box -5 0 541 1194
use M2M3_CDNS_524688791851529  M2M3_CDNS_524688791851529_0
timestamp 1707688321
transform 1 0 5628 0 1 5188
box -5 0 541 6154
use M2M3_CDNS_524688791851529  M2M3_CDNS_524688791851529_1
timestamp 1707688321
transform 1 0 216 0 1 5188
box -5 0 541 6154
use M2M3_CDNS_524688791851529  M2M3_CDNS_524688791851529_2
timestamp 1707688321
transform 1 0 12848 0 1 5140
box -5 0 541 6154
use M2M3_CDNS_524688791851529  M2M3_CDNS_524688791851529_3
timestamp 1707688321
transform 1 0 3824 0 1 5188
box -5 0 541 6154
use M2M3_CDNS_524688791851529  M2M3_CDNS_524688791851529_4
timestamp 1707688321
transform 1 0 -1593 0 1 5140
box -5 0 541 6154
use M2M3_CDNS_524688791851529  M2M3_CDNS_524688791851529_5
timestamp 1707688321
transform 1 0 2020 0 1 5188
box -5 0 541 6154
use M2M3_CDNS_524688791851529  M2M3_CDNS_524688791851529_6
timestamp 1707688321
transform 1 0 7433 0 1 5188
box -5 0 541 6154
use M2M3_CDNS_524688791851529  M2M3_CDNS_524688791851529_7
timestamp 1707688321
transform 1 0 9234 0 1 5188
box -5 0 541 6154
use M2M3_CDNS_524688791851529  M2M3_CDNS_524688791851529_8
timestamp 1707688321
transform 1 0 11047 0 1 5188
box -5 0 541 6154
use M2M3_CDNS_524688791851530  M2M3_CDNS_524688791851530_0
timestamp 1707688321
transform 1 0 13744 0 1 5140
box -5 0 541 6714
use M2M3_CDNS_524688791851531  M2M3_CDNS_524688791851531_0
timestamp 1707688321
transform 1 0 11934 0 1 5140
box -5 0 541 6954
use M2M3_CDNS_524688791851532  M2M3_CDNS_524688791851532_0
timestamp 1707688321
transform 1 0 214 0 1 3527
box -5 0 541 474
use M2M3_CDNS_524688791851532  M2M3_CDNS_524688791851532_1
timestamp 1707688321
transform 1 0 3816 0 1 3527
box -5 0 541 474
use M2M3_CDNS_524688791851532  M2M3_CDNS_524688791851532_2
timestamp 1707688321
transform 1 0 5623 0 1 3527
box -5 0 541 474
use M2M3_CDNS_524688791851532  M2M3_CDNS_524688791851532_3
timestamp 1707688321
transform 1 0 2018 0 1 3527
box -5 0 541 474
use M2M3_CDNS_524688791851532  M2M3_CDNS_524688791851532_4
timestamp 1707688321
transform 1 0 11035 0 1 3527
box -5 0 541 474
use M2M3_CDNS_524688791851532  M2M3_CDNS_524688791851532_5
timestamp 1707688321
transform 1 0 12834 0 1 3527
box -5 0 541 474
use M2M3_CDNS_524688791851532  M2M3_CDNS_524688791851532_6
timestamp 1707688321
transform 1 0 7424 0 1 3527
box -5 0 541 474
use M2M3_CDNS_524688791851532  M2M3_CDNS_524688791851532_7
timestamp 1707688321
transform 1 0 9234 0 1 3527
box -5 0 541 474
use M2M3_CDNS_524688791851533  M2M3_CDNS_524688791851533_0
timestamp 1707688321
transform 1 0 6527 0 1 1147
box -5 0 541 1754
use M2M3_CDNS_524688791851533  M2M3_CDNS_524688791851533_1
timestamp 1707688321
transform 1 0 4717 0 1 1147
box -5 0 541 1754
use M2M3_CDNS_524688791851533  M2M3_CDNS_524688791851533_2
timestamp 1707688321
transform 1 0 -4303 0 1 1147
box -5 0 541 1754
use M2M3_CDNS_524688791851533  M2M3_CDNS_524688791851533_3
timestamp 1707688321
transform 1 0 -2499 0 1 1147
box -5 0 541 1754
use M2M3_CDNS_524688791851533  M2M3_CDNS_524688791851533_4
timestamp 1707688321
transform 1 0 -695 0 1 1147
box -5 0 541 1754
use M2M3_CDNS_524688791851533  M2M3_CDNS_524688791851533_5
timestamp 1707688321
transform 1 0 1109 0 1 1147
box -5 0 541 1754
use M2M3_CDNS_524688791851533  M2M3_CDNS_524688791851533_6
timestamp 1707688321
transform 1 0 2913 0 1 1147
box -5 0 541 1754
use M2M3_CDNS_524688791851533  M2M3_CDNS_524688791851533_7
timestamp 1707688321
transform 1 0 13746 0 1 1147
box -5 0 541 1754
use M2M3_CDNS_524688791851533  M2M3_CDNS_524688791851533_8
timestamp 1707688321
transform 1 0 11940 0 1 1147
box -5 0 541 1754
use M2M3_CDNS_524688791851533  M2M3_CDNS_524688791851533_9
timestamp 1707688321
transform 1 0 10134 0 1 1147
box -5 0 541 1754
use M2M3_CDNS_524688791851533  M2M3_CDNS_524688791851533_10
timestamp 1707688321
transform 1 0 8322 0 1 1147
box -5 0 541 1754
use M3M4_CDNS_524688791851511  M3M4_CDNS_524688791851511_0
timestamp 1707688321
transform 1 0 -1586 0 1 3543
box -1 0 545 1196
use M3M4_CDNS_524688791851511  M3M4_CDNS_524688791851511_1
timestamp 1707688321
transform 1 0 -3404 0 1 3543
box -1 0 545 1196
use M3M4_CDNS_524688791851512  M3M4_CDNS_524688791851512_0
timestamp 1707688321
transform 1 0 210 0 1 3526
box -1 0 545 476
use M3M4_CDNS_524688791851512  M3M4_CDNS_524688791851512_1
timestamp 1707688321
transform 1 0 3812 0 1 3526
box -1 0 545 476
use M3M4_CDNS_524688791851512  M3M4_CDNS_524688791851512_2
timestamp 1707688321
transform 1 0 5619 0 1 3526
box -1 0 545 476
use M3M4_CDNS_524688791851512  M3M4_CDNS_524688791851512_3
timestamp 1707688321
transform 1 0 12830 0 1 3526
box -1 0 545 476
use M3M4_CDNS_524688791851512  M3M4_CDNS_524688791851512_4
timestamp 1707688321
transform 1 0 11031 0 1 3526
box -1 0 545 476
use M3M4_CDNS_524688791851512  M3M4_CDNS_524688791851512_5
timestamp 1707688321
transform 1 0 9230 0 1 3526
box -1 0 545 476
use M3M4_CDNS_524688791851512  M3M4_CDNS_524688791851512_6
timestamp 1707688321
transform 1 0 7420 0 1 3526
box -1 0 545 476
use M3M4_CDNS_524688791851512  M3M4_CDNS_524688791851512_7
timestamp 1707688321
transform 1 0 2013 0 1 3526
box -1 0 545 476
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_0
timestamp 1707688321
transform -1 0 1107 0 1 753
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_1
timestamp 1707688321
transform 1 0 3115 0 1 753
box 0 0 1 1
use PYres_CDNS_524688791856  PYres_CDNS_524688791856_0
timestamp 1707688321
transform -1 0 3131 0 1 736
box -50 0 2090 100
use sky130_fd_io__esd_signal_50_sym_hv_2k_dnwl_aup1_b  sky130_fd_io__esd_signal_50_sym_hv_2k_dnwl_aup1_b_0
timestamp 1707688321
transform 1 0 -185 0 1 0
box -5020 0 15370 13100
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_0
timestamp 1707688321
transform -1 0 12291 0 1 981
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_1
timestamp 1707688321
transform -1 0 8618 0 1 981
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_0
timestamp 1707688321
transform -1 0 13208 0 1 981
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_1
timestamp 1707688321
transform -1 0 10487 0 1 981
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_2
timestamp 1707688321
transform -1 0 11321 0 1 981
box 0 0 1 1
use sky130_fd_io__tk_em2o_CDNS_52468879185636  sky130_fd_io__tk_em2o_CDNS_52468879185636_0
timestamp 1707688321
transform 0 1 11750 1 0 837
box 0 0 1 1
use sky130_fd_io__tk_em2o_CDNS_52468879185636  sky130_fd_io__tk_em2o_CDNS_52468879185636_1
timestamp 1707688321
transform 0 1 10781 1 0 837
box 0 0 1 1
use sky130_fd_io__tk_em2s_CDNS_52468879185635  sky130_fd_io__tk_em2s_CDNS_52468879185635_0
timestamp 1707688321
transform 0 1 9005 1 0 837
box 0 0 1 1
<< labels >>
flabel comment s 9434 1085 9434 1085 0 FreeSans 200 0 0 0 force_lo_h
flabel comment s 1690 1091 1690 1091 0 FreeSans 200 0 0 0 pd_h<2>
flabel comment s 6865 1091 6865 1091 0 FreeSans 200 0 0 0 pd_h<3>
flabel comment s 7455 681 7455 681 0 FreeSans 200 0 0 0 tie_lo_esd
flabel metal1 s 13482 892 13532 945 0 FreeSans 200 0 0 0 pd_h<3>
port 2 nsew
flabel metal1 s 13959 947 14009 999 7 FreeSans 400 0 0 0 pd_h<2>
port 4 nsew
flabel metal1 s 13479 648 13532 705 7 FreeSans 400 0 0 0 tie_lo_esd
port 3 nsew
flabel metal1 s 13482 733 13532 790 7 FreeSans 400 0 0 0 pd_h<4>
port 5 nsew
flabel metal4 s 11132 3657 11466 3855 0 FreeSans 200 0 0 0 pad
port 6 nsew
flabel metal4 s 12970 3669 13251 3813 0 FreeSans 200 0 0 0 pad
port 6 nsew
flabel metal2 s 14724 4086 14906 4160 0 FreeSans 400 0 0 0 vcc_io
port 7 nsew
flabel metal2 s 12091 0 12313 74 0 FreeSans 400 0 0 0 vgnd_io
port 8 nsew
flabel metal2 s 10286 40 10508 114 0 FreeSans 400 0 0 0 vgnd_io
port 8 nsew
flabel metal2 s 8483 0 8705 74 0 FreeSans 400 0 0 0 vgnd_io
port 8 nsew
flabel metal2 s 6679 0 6901 74 0 FreeSans 400 0 0 0 vgnd_io
port 8 nsew
flabel metal2 s 4875 497 5097 571 0 FreeSans 400 0 0 0 vgnd_io
port 8 nsew
flabel metal2 s 13895 0 14117 74 0 FreeSans 400 0 0 0 vgnd_io
port 8 nsew
flabel metal2 s 3071 0 3293 74 0 FreeSans 400 0 0 0 vgnd_io
port 8 nsew
flabel metal2 s 1267 0 1489 74 0 FreeSans 400 0 0 0 vgnd_io
port 8 nsew
flabel metal2 s -537 0 -315 74 0 FreeSans 400 0 0 0 vgnd_io
port 8 nsew
flabel metal2 s -2341 0 -2119 74 0 FreeSans 400 0 0 0 vgnd_io
port 8 nsew
flabel metal2 s -4145 0 -3923 74 0 FreeSans 400 0 0 0 vgnd_io
port 8 nsew
<< properties >>
string GDS_END 94168976
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 93932058
string path 327.725 423.325 327.725 459.300 
<< end >>
