magic
tech sky130B
timestamp 1707688321
<< properties >>
string GDS_END 24028
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 23704
<< end >>
