magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect 12562 6849 17453 7153
rect 61 4666 2365 5941
rect 669 4576 883 4666
rect 12562 3852 12866 6849
rect 13266 4267 16749 6449
rect 12562 3826 12603 3852
rect 12825 3826 12866 3852
rect 17149 3852 17453 6849
rect 17149 3826 17190 3852
rect 17412 3826 17453 3852
<< pwell >>
rect 2914 6580 3100 6695
rect 2845 5096 4223 5182
rect 1421 4428 1555 4516
rect 1800 3848 2186 4406
rect 13004 6510 17011 6712
rect 13072 4256 13206 6510
rect 13004 4195 13206 4256
rect 16809 4195 17011 6510
rect 13004 3993 17011 4195
rect 12603 3774 12825 3852
rect 17190 3774 17412 3852
rect 2845 3506 4223 3592
<< mvnmos >>
rect 1826 3927 1910 4127
rect 2076 3927 2160 4127
<< mvpmos >>
rect 514 5541 714 5625
rect 838 5541 1038 5625
<< mvndiff >>
rect 2940 6651 3074 6669
rect 2940 6617 2958 6651
rect 2992 6617 3026 6651
rect 3060 6617 3074 6651
rect 2940 6606 3074 6617
rect 1826 4372 1910 4380
rect 1826 4338 1838 4372
rect 1872 4338 1910 4372
rect 1826 4127 1910 4338
rect 2076 4372 2160 4380
rect 2076 4338 2114 4372
rect 2148 4338 2160 4372
rect 2076 4127 2160 4338
rect 1826 3916 1910 3927
rect 1826 3882 1838 3916
rect 1872 3882 1910 3916
rect 2076 3916 2160 3927
rect 1826 3874 1910 3882
rect 2076 3882 2114 3916
rect 2148 3882 2160 3916
rect 2076 3874 2160 3882
<< mvpdiff >>
rect 193 5837 261 5875
rect 193 5803 201 5837
rect 235 5803 261 5837
rect 193 5791 261 5803
rect 1291 5837 1359 5875
rect 1291 5803 1317 5837
rect 1351 5803 1359 5837
rect 1291 5791 1359 5803
rect 193 5587 514 5625
rect 193 5553 201 5587
rect 235 5553 269 5587
rect 303 5553 514 5587
rect 193 5541 514 5553
rect 714 5587 838 5625
rect 714 5553 725 5587
rect 759 5553 793 5587
rect 827 5553 838 5587
rect 714 5541 838 5553
rect 1038 5587 1359 5625
rect 1038 5553 1249 5587
rect 1283 5553 1317 5587
rect 1351 5553 1359 5587
rect 1038 5541 1359 5553
<< mvndiffc >>
rect 2958 6617 2992 6651
rect 3026 6617 3060 6651
rect 1838 4338 1872 4372
rect 2114 4338 2148 4372
rect 1838 3882 1872 3916
rect 2114 3882 2148 3916
<< mvpdiffc >>
rect 201 5803 235 5837
rect 1317 5803 1351 5837
rect 201 5553 235 5587
rect 269 5553 303 5587
rect 725 5553 759 5587
rect 793 5553 827 5587
rect 1249 5553 1283 5587
rect 1317 5553 1351 5587
<< psubdiff >>
rect 13030 6662 16985 6686
rect 13030 6628 13092 6662
rect 13126 6661 16985 6662
rect 13126 6628 16900 6661
rect 13030 6627 16900 6628
rect 16934 6627 16985 6661
rect 13030 6594 16985 6627
rect 13030 6560 13065 6594
rect 13099 6593 16985 6594
rect 13099 6560 16927 6593
rect 13030 6559 16927 6560
rect 16961 6559 16985 6593
rect 13030 6536 16985 6559
rect 13098 4230 13180 6536
rect 13030 4169 13180 4230
rect 16835 4169 16985 6536
rect 13030 4145 16985 4169
rect 13030 4111 13065 4145
rect 13099 4111 16927 4145
rect 16961 4111 16985 4145
rect 13030 4077 16985 4111
rect 13030 4043 13092 4077
rect 13126 4043 16900 4077
rect 16934 4043 16985 4077
rect 13030 4019 16985 4043
<< nsubdiff >>
rect 12629 6984 12697 7086
rect 17219 7052 17253 7086
rect 17287 7052 17386 7086
rect 17219 7018 17386 7052
rect 17219 6984 17284 7018
rect 12629 6954 12765 6984
rect 12663 6920 12765 6954
rect 12629 6916 12765 6920
rect 17151 6950 17284 6984
rect 17151 6916 17216 6950
rect 12629 6886 12799 6916
rect 12731 6818 12799 6886
rect 12629 3800 12799 3860
rect 17216 3800 17386 3924
<< mvpsubdiff >>
rect 2871 5122 2895 5156
rect 2929 5122 2964 5156
rect 2998 5122 3033 5156
rect 3067 5122 3102 5156
rect 3136 5122 3171 5156
rect 3205 5122 3240 5156
rect 3274 5122 3309 5156
rect 3343 5122 3378 5156
rect 3412 5122 3447 5156
rect 3481 5122 3516 5156
rect 3550 5122 3585 5156
rect 3619 5122 3654 5156
rect 3688 5122 3723 5156
rect 3757 5122 3792 5156
rect 3826 5122 3861 5156
rect 3895 5122 3930 5156
rect 3964 5122 3999 5156
rect 4033 5122 4069 5156
rect 4103 5122 4139 5156
rect 4173 5122 4197 5156
rect 1447 4488 1529 4490
rect 1447 4454 1471 4488
rect 1505 4454 1529 4488
rect 2871 3532 2895 3566
rect 2929 3532 2964 3566
rect 2998 3532 3033 3566
rect 3067 3532 3102 3566
rect 3136 3532 3171 3566
rect 3205 3532 3240 3566
rect 3274 3532 3309 3566
rect 3343 3532 3378 3566
rect 3412 3532 3447 3566
rect 3481 3532 3516 3566
rect 3550 3532 3585 3566
rect 3619 3532 3654 3566
rect 3688 3532 3723 3566
rect 3757 3532 3792 3566
rect 3826 3532 3861 3566
rect 3895 3532 3930 3566
rect 3964 3532 3999 3566
rect 4033 3532 4069 3566
rect 4103 3532 4139 3566
rect 4173 3532 4197 3566
<< mvnsubdiff >>
rect 735 4644 759 4678
rect 793 4644 817 4678
rect 735 4642 817 4644
rect 13332 6279 13366 6383
rect 13400 6349 13474 6383
rect 13508 6349 13556 6383
rect 13590 6349 13624 6383
rect 13658 6349 13692 6383
rect 13726 6349 13760 6383
rect 13794 6349 13828 6383
rect 13862 6349 13896 6383
rect 13930 6349 13964 6383
rect 13998 6349 14032 6383
rect 14066 6349 14100 6383
rect 14134 6349 14168 6383
rect 14202 6349 14236 6383
rect 14270 6349 14304 6383
rect 14338 6349 14372 6383
rect 14406 6349 14440 6383
rect 14474 6349 14508 6383
rect 14542 6349 14576 6383
rect 14610 6349 14644 6383
rect 14678 6349 14712 6383
rect 14746 6349 14780 6383
rect 14814 6349 14848 6383
rect 14882 6349 14916 6383
rect 14950 6349 14984 6383
rect 15018 6349 15053 6383
rect 15087 6349 15122 6383
rect 15156 6349 15191 6383
rect 15225 6349 15260 6383
rect 15294 6349 15329 6383
rect 15363 6349 15398 6383
rect 15432 6349 15467 6383
rect 15501 6349 15536 6383
rect 15570 6349 15605 6383
rect 15639 6349 15674 6383
rect 15708 6349 15743 6383
rect 15777 6349 15812 6383
rect 15846 6349 15881 6383
rect 15915 6349 15950 6383
rect 15984 6349 16019 6383
rect 16053 6349 16088 6383
rect 16122 6349 16157 6383
rect 16191 6349 16226 6383
rect 16260 6349 16295 6383
rect 16329 6349 16364 6383
rect 16398 6349 16433 6383
rect 16467 6349 16502 6383
rect 16536 6349 16683 6383
rect 16649 6279 16683 6315
rect 13332 6210 13366 6245
rect 13332 6141 13366 6176
rect 13332 6072 13366 6107
rect 13332 6003 13366 6038
rect 16649 6209 16683 6245
rect 16649 6139 16683 6175
rect 16649 6069 16683 6105
rect 16649 5999 16683 6035
rect 13332 5934 13366 5969
rect 13332 5879 13366 5900
rect 16649 5929 16683 5965
rect 16649 5879 16683 5895
rect 13332 5865 13407 5879
rect 13366 5845 13407 5865
rect 13441 5845 13475 5879
rect 13509 5845 13543 5879
rect 13577 5845 13611 5879
rect 13645 5845 13679 5879
rect 13713 5845 13747 5879
rect 13781 5845 13815 5879
rect 13849 5845 13883 5879
rect 13917 5845 13951 5879
rect 13985 5845 14019 5879
rect 14053 5845 14087 5879
rect 14121 5845 14155 5879
rect 14189 5845 14223 5879
rect 14257 5845 14291 5879
rect 14325 5845 14359 5879
rect 14393 5845 14427 5879
rect 14461 5845 14495 5879
rect 14529 5845 14563 5879
rect 14597 5845 14631 5879
rect 14665 5845 14699 5879
rect 14733 5845 14767 5879
rect 14801 5845 14835 5879
rect 14869 5845 14903 5879
rect 14937 5845 14971 5879
rect 15005 5845 15039 5879
rect 15073 5845 15107 5879
rect 15141 5845 15175 5879
rect 15209 5845 15243 5879
rect 15277 5845 15311 5879
rect 15345 5845 15379 5879
rect 15413 5845 15447 5879
rect 15481 5845 15515 5879
rect 15549 5845 15583 5879
rect 15617 5845 15651 5879
rect 15685 5845 15719 5879
rect 15753 5845 15787 5879
rect 15821 5845 15855 5879
rect 15889 5845 15923 5879
rect 15957 5845 15991 5879
rect 16025 5845 16059 5879
rect 16093 5845 16127 5879
rect 16161 5845 16195 5879
rect 16229 5845 16263 5879
rect 16297 5845 16332 5879
rect 16366 5845 16401 5879
rect 16435 5845 16470 5879
rect 16504 5845 16539 5879
rect 16573 5859 16683 5879
rect 16573 5845 16649 5859
rect 13332 5796 13366 5831
rect 13332 5727 13366 5762
rect 16649 5789 16683 5825
rect 13332 5658 13366 5693
rect 13332 5589 13366 5624
rect 13332 5520 13366 5555
rect 13332 5451 13366 5486
rect 16649 5719 16683 5755
rect 16649 5649 16683 5685
rect 16649 5579 16683 5615
rect 16649 5509 16683 5545
rect 13332 5381 13366 5417
rect 16649 5439 16683 5475
rect 16649 5375 16683 5405
rect 13366 5347 13407 5375
rect 13332 5341 13407 5347
rect 13441 5341 13475 5375
rect 13509 5341 13543 5375
rect 13577 5341 13611 5375
rect 13645 5341 13679 5375
rect 13713 5341 13747 5375
rect 13781 5341 13815 5375
rect 13849 5341 13883 5375
rect 13917 5341 13951 5375
rect 13985 5341 14019 5375
rect 14053 5341 14087 5375
rect 14121 5341 14155 5375
rect 14189 5341 14223 5375
rect 14257 5341 14291 5375
rect 14325 5341 14359 5375
rect 14393 5341 14427 5375
rect 14461 5341 14495 5375
rect 14529 5341 14563 5375
rect 14597 5341 14631 5375
rect 14665 5341 14699 5375
rect 14733 5341 14767 5375
rect 14801 5341 14835 5375
rect 14869 5341 14903 5375
rect 14937 5341 14971 5375
rect 15005 5341 15039 5375
rect 15073 5341 15107 5375
rect 15141 5341 15175 5375
rect 15209 5341 15243 5375
rect 15277 5341 15311 5375
rect 15345 5341 15379 5375
rect 15413 5341 15447 5375
rect 15481 5341 15515 5375
rect 15549 5341 15583 5375
rect 15617 5341 15651 5375
rect 15685 5341 15719 5375
rect 15753 5341 15787 5375
rect 15821 5341 15855 5375
rect 15889 5341 15923 5375
rect 15957 5341 15991 5375
rect 16025 5341 16059 5375
rect 16093 5341 16127 5375
rect 16161 5341 16195 5375
rect 16229 5341 16263 5375
rect 16297 5341 16332 5375
rect 16366 5341 16401 5375
rect 16435 5341 16470 5375
rect 16504 5341 16539 5375
rect 16573 5369 16683 5375
rect 16573 5341 16649 5369
rect 13332 5311 13366 5341
rect 13332 5241 13366 5277
rect 16649 5299 16683 5335
rect 13332 5171 13366 5207
rect 13332 5101 13366 5137
rect 13332 5031 13366 5067
rect 13332 4961 13366 4997
rect 16649 5230 16683 5265
rect 16649 5161 16683 5196
rect 16649 5092 16683 5127
rect 16649 5023 16683 5058
rect 13332 4891 13366 4927
rect 16649 4954 16683 4989
rect 16649 4885 16683 4920
rect 13366 4857 13407 4871
rect 13332 4837 13407 4857
rect 13441 4837 13475 4871
rect 13509 4837 13543 4871
rect 13577 4837 13611 4871
rect 13645 4837 13679 4871
rect 13713 4837 13747 4871
rect 13781 4837 13815 4871
rect 13849 4837 13883 4871
rect 13917 4837 13951 4871
rect 13985 4837 14019 4871
rect 14053 4837 14087 4871
rect 14121 4837 14155 4871
rect 14189 4837 14223 4871
rect 14257 4837 14291 4871
rect 14325 4837 14359 4871
rect 14393 4837 14427 4871
rect 14461 4837 14495 4871
rect 14529 4837 14563 4871
rect 14597 4837 14631 4871
rect 14665 4837 14699 4871
rect 14733 4837 14767 4871
rect 14801 4837 14835 4871
rect 14869 4837 14903 4871
rect 14937 4837 14971 4871
rect 15005 4837 15039 4871
rect 15073 4837 15107 4871
rect 15141 4837 15175 4871
rect 15209 4837 15243 4871
rect 15277 4837 15311 4871
rect 15345 4837 15379 4871
rect 15413 4837 15447 4871
rect 15481 4837 15515 4871
rect 15549 4837 15583 4871
rect 15617 4837 15651 4871
rect 15685 4837 15719 4871
rect 15753 4837 15787 4871
rect 15821 4837 15855 4871
rect 15889 4837 15923 4871
rect 15957 4837 15991 4871
rect 16025 4837 16059 4871
rect 16093 4837 16127 4871
rect 16161 4837 16195 4871
rect 16229 4837 16263 4871
rect 16297 4837 16332 4871
rect 16366 4837 16401 4871
rect 16435 4837 16470 4871
rect 16504 4837 16539 4871
rect 16573 4851 16649 4871
rect 16573 4837 16683 4851
rect 13332 4821 13366 4837
rect 13332 4751 13366 4787
rect 16649 4816 16683 4837
rect 16649 4747 16683 4782
rect 13332 4681 13366 4717
rect 13332 4611 13366 4647
rect 13332 4541 13366 4577
rect 13332 4471 13366 4507
rect 16649 4678 16683 4713
rect 16649 4609 16683 4644
rect 16649 4540 16683 4575
rect 16649 4471 16683 4506
rect 13332 4401 13366 4437
rect 13332 4333 13436 4367
rect 13470 4333 13505 4367
rect 13539 4333 13574 4367
rect 13608 4333 13643 4367
rect 13677 4333 13712 4367
rect 13746 4333 13781 4367
rect 13815 4333 13850 4367
rect 13884 4333 13919 4367
rect 13953 4333 13988 4367
rect 14022 4333 14057 4367
rect 14091 4333 14126 4367
rect 14160 4333 14195 4367
rect 14229 4333 14264 4367
rect 14298 4333 14333 4367
rect 14367 4333 14402 4367
rect 14436 4333 14471 4367
rect 14505 4333 14540 4367
rect 14574 4333 14609 4367
rect 14643 4333 14678 4367
rect 14712 4333 14747 4367
rect 14781 4333 14816 4367
rect 14850 4333 14885 4367
rect 14919 4333 14954 4367
rect 14988 4333 15023 4367
rect 15057 4333 15092 4367
rect 15126 4333 15161 4367
rect 15195 4333 15230 4367
rect 15264 4333 15299 4367
rect 15333 4333 15368 4367
rect 15402 4333 15437 4367
rect 15471 4333 15506 4367
rect 15540 4333 15575 4367
rect 15609 4333 15644 4367
rect 15678 4333 15713 4367
rect 15747 4333 15782 4367
rect 15816 4333 15851 4367
rect 15885 4333 15920 4367
rect 15954 4333 15989 4367
rect 16023 4333 16058 4367
rect 16092 4333 16127 4367
rect 16161 4333 16196 4367
rect 16230 4333 16265 4367
rect 16299 4333 16335 4367
rect 16369 4333 16405 4367
rect 16439 4333 16475 4367
rect 16509 4333 16545 4367
rect 16579 4333 16615 4367
rect 16649 4333 16683 4437
<< psubdiffcont >>
rect 13092 6628 13126 6662
rect 16900 6627 16934 6661
rect 13065 6560 13099 6594
rect 16927 6559 16961 6593
rect 13065 4111 13099 4145
rect 16927 4111 16961 4145
rect 13092 4043 13126 4077
rect 16900 4043 16934 4077
<< nsubdiffcont >>
rect 12697 6984 17219 7086
rect 17253 7052 17287 7086
rect 12629 6920 12663 6954
rect 12765 6916 17151 6984
rect 17284 6950 17386 7018
rect 12629 6818 12731 6886
rect 12629 3860 12799 6818
rect 17216 3924 17386 6950
<< mvpsubdiffcont >>
rect 2895 5122 2929 5156
rect 2964 5122 2998 5156
rect 3033 5122 3067 5156
rect 3102 5122 3136 5156
rect 3171 5122 3205 5156
rect 3240 5122 3274 5156
rect 3309 5122 3343 5156
rect 3378 5122 3412 5156
rect 3447 5122 3481 5156
rect 3516 5122 3550 5156
rect 3585 5122 3619 5156
rect 3654 5122 3688 5156
rect 3723 5122 3757 5156
rect 3792 5122 3826 5156
rect 3861 5122 3895 5156
rect 3930 5122 3964 5156
rect 3999 5122 4033 5156
rect 4069 5122 4103 5156
rect 4139 5122 4173 5156
rect 1471 4454 1505 4488
rect 2895 3532 2929 3566
rect 2964 3532 2998 3566
rect 3033 3532 3067 3566
rect 3102 3532 3136 3566
rect 3171 3532 3205 3566
rect 3240 3532 3274 3566
rect 3309 3532 3343 3566
rect 3378 3532 3412 3566
rect 3447 3532 3481 3566
rect 3516 3532 3550 3566
rect 3585 3532 3619 3566
rect 3654 3532 3688 3566
rect 3723 3532 3757 3566
rect 3792 3532 3826 3566
rect 3861 3532 3895 3566
rect 3930 3532 3964 3566
rect 3999 3532 4033 3566
rect 4069 3532 4103 3566
rect 4139 3532 4173 3566
<< mvnsubdiffcont >>
rect 759 4644 793 4678
rect 13366 6349 13400 6383
rect 13474 6349 13508 6383
rect 13556 6349 13590 6383
rect 13624 6349 13658 6383
rect 13692 6349 13726 6383
rect 13760 6349 13794 6383
rect 13828 6349 13862 6383
rect 13896 6349 13930 6383
rect 13964 6349 13998 6383
rect 14032 6349 14066 6383
rect 14100 6349 14134 6383
rect 14168 6349 14202 6383
rect 14236 6349 14270 6383
rect 14304 6349 14338 6383
rect 14372 6349 14406 6383
rect 14440 6349 14474 6383
rect 14508 6349 14542 6383
rect 14576 6349 14610 6383
rect 14644 6349 14678 6383
rect 14712 6349 14746 6383
rect 14780 6349 14814 6383
rect 14848 6349 14882 6383
rect 14916 6349 14950 6383
rect 14984 6349 15018 6383
rect 15053 6349 15087 6383
rect 15122 6349 15156 6383
rect 15191 6349 15225 6383
rect 15260 6349 15294 6383
rect 15329 6349 15363 6383
rect 15398 6349 15432 6383
rect 15467 6349 15501 6383
rect 15536 6349 15570 6383
rect 15605 6349 15639 6383
rect 15674 6349 15708 6383
rect 15743 6349 15777 6383
rect 15812 6349 15846 6383
rect 15881 6349 15915 6383
rect 15950 6349 15984 6383
rect 16019 6349 16053 6383
rect 16088 6349 16122 6383
rect 16157 6349 16191 6383
rect 16226 6349 16260 6383
rect 16295 6349 16329 6383
rect 16364 6349 16398 6383
rect 16433 6349 16467 6383
rect 16502 6349 16536 6383
rect 13332 6245 13366 6279
rect 16649 6315 16683 6349
rect 13332 6176 13366 6210
rect 13332 6107 13366 6141
rect 13332 6038 13366 6072
rect 13332 5969 13366 6003
rect 16649 6245 16683 6279
rect 16649 6175 16683 6209
rect 16649 6105 16683 6139
rect 16649 6035 16683 6069
rect 13332 5900 13366 5934
rect 16649 5965 16683 5999
rect 16649 5895 16683 5929
rect 13332 5831 13366 5865
rect 13407 5845 13441 5879
rect 13475 5845 13509 5879
rect 13543 5845 13577 5879
rect 13611 5845 13645 5879
rect 13679 5845 13713 5879
rect 13747 5845 13781 5879
rect 13815 5845 13849 5879
rect 13883 5845 13917 5879
rect 13951 5845 13985 5879
rect 14019 5845 14053 5879
rect 14087 5845 14121 5879
rect 14155 5845 14189 5879
rect 14223 5845 14257 5879
rect 14291 5845 14325 5879
rect 14359 5845 14393 5879
rect 14427 5845 14461 5879
rect 14495 5845 14529 5879
rect 14563 5845 14597 5879
rect 14631 5845 14665 5879
rect 14699 5845 14733 5879
rect 14767 5845 14801 5879
rect 14835 5845 14869 5879
rect 14903 5845 14937 5879
rect 14971 5845 15005 5879
rect 15039 5845 15073 5879
rect 15107 5845 15141 5879
rect 15175 5845 15209 5879
rect 15243 5845 15277 5879
rect 15311 5845 15345 5879
rect 15379 5845 15413 5879
rect 15447 5845 15481 5879
rect 15515 5845 15549 5879
rect 15583 5845 15617 5879
rect 15651 5845 15685 5879
rect 15719 5845 15753 5879
rect 15787 5845 15821 5879
rect 15855 5845 15889 5879
rect 15923 5845 15957 5879
rect 15991 5845 16025 5879
rect 16059 5845 16093 5879
rect 16127 5845 16161 5879
rect 16195 5845 16229 5879
rect 16263 5845 16297 5879
rect 16332 5845 16366 5879
rect 16401 5845 16435 5879
rect 16470 5845 16504 5879
rect 16539 5845 16573 5879
rect 13332 5762 13366 5796
rect 16649 5825 16683 5859
rect 16649 5755 16683 5789
rect 13332 5693 13366 5727
rect 13332 5624 13366 5658
rect 13332 5555 13366 5589
rect 13332 5486 13366 5520
rect 16649 5685 16683 5719
rect 16649 5615 16683 5649
rect 16649 5545 16683 5579
rect 16649 5475 16683 5509
rect 13332 5417 13366 5451
rect 13332 5347 13366 5381
rect 16649 5405 16683 5439
rect 13407 5341 13441 5375
rect 13475 5341 13509 5375
rect 13543 5341 13577 5375
rect 13611 5341 13645 5375
rect 13679 5341 13713 5375
rect 13747 5341 13781 5375
rect 13815 5341 13849 5375
rect 13883 5341 13917 5375
rect 13951 5341 13985 5375
rect 14019 5341 14053 5375
rect 14087 5341 14121 5375
rect 14155 5341 14189 5375
rect 14223 5341 14257 5375
rect 14291 5341 14325 5375
rect 14359 5341 14393 5375
rect 14427 5341 14461 5375
rect 14495 5341 14529 5375
rect 14563 5341 14597 5375
rect 14631 5341 14665 5375
rect 14699 5341 14733 5375
rect 14767 5341 14801 5375
rect 14835 5341 14869 5375
rect 14903 5341 14937 5375
rect 14971 5341 15005 5375
rect 15039 5341 15073 5375
rect 15107 5341 15141 5375
rect 15175 5341 15209 5375
rect 15243 5341 15277 5375
rect 15311 5341 15345 5375
rect 15379 5341 15413 5375
rect 15447 5341 15481 5375
rect 15515 5341 15549 5375
rect 15583 5341 15617 5375
rect 15651 5341 15685 5375
rect 15719 5341 15753 5375
rect 15787 5341 15821 5375
rect 15855 5341 15889 5375
rect 15923 5341 15957 5375
rect 15991 5341 16025 5375
rect 16059 5341 16093 5375
rect 16127 5341 16161 5375
rect 16195 5341 16229 5375
rect 16263 5341 16297 5375
rect 16332 5341 16366 5375
rect 16401 5341 16435 5375
rect 16470 5341 16504 5375
rect 16539 5341 16573 5375
rect 13332 5277 13366 5311
rect 16649 5335 16683 5369
rect 16649 5265 16683 5299
rect 13332 5207 13366 5241
rect 13332 5137 13366 5171
rect 13332 5067 13366 5101
rect 13332 4997 13366 5031
rect 16649 5196 16683 5230
rect 16649 5127 16683 5161
rect 16649 5058 16683 5092
rect 16649 4989 16683 5023
rect 13332 4927 13366 4961
rect 13332 4857 13366 4891
rect 16649 4920 16683 4954
rect 13407 4837 13441 4871
rect 13475 4837 13509 4871
rect 13543 4837 13577 4871
rect 13611 4837 13645 4871
rect 13679 4837 13713 4871
rect 13747 4837 13781 4871
rect 13815 4837 13849 4871
rect 13883 4837 13917 4871
rect 13951 4837 13985 4871
rect 14019 4837 14053 4871
rect 14087 4837 14121 4871
rect 14155 4837 14189 4871
rect 14223 4837 14257 4871
rect 14291 4837 14325 4871
rect 14359 4837 14393 4871
rect 14427 4837 14461 4871
rect 14495 4837 14529 4871
rect 14563 4837 14597 4871
rect 14631 4837 14665 4871
rect 14699 4837 14733 4871
rect 14767 4837 14801 4871
rect 14835 4837 14869 4871
rect 14903 4837 14937 4871
rect 14971 4837 15005 4871
rect 15039 4837 15073 4871
rect 15107 4837 15141 4871
rect 15175 4837 15209 4871
rect 15243 4837 15277 4871
rect 15311 4837 15345 4871
rect 15379 4837 15413 4871
rect 15447 4837 15481 4871
rect 15515 4837 15549 4871
rect 15583 4837 15617 4871
rect 15651 4837 15685 4871
rect 15719 4837 15753 4871
rect 15787 4837 15821 4871
rect 15855 4837 15889 4871
rect 15923 4837 15957 4871
rect 15991 4837 16025 4871
rect 16059 4837 16093 4871
rect 16127 4837 16161 4871
rect 16195 4837 16229 4871
rect 16263 4837 16297 4871
rect 16332 4837 16366 4871
rect 16401 4837 16435 4871
rect 16470 4837 16504 4871
rect 16539 4837 16573 4871
rect 16649 4851 16683 4885
rect 13332 4787 13366 4821
rect 13332 4717 13366 4751
rect 16649 4782 16683 4816
rect 13332 4647 13366 4681
rect 13332 4577 13366 4611
rect 13332 4507 13366 4541
rect 13332 4437 13366 4471
rect 16649 4713 16683 4747
rect 16649 4644 16683 4678
rect 16649 4575 16683 4609
rect 16649 4506 16683 4540
rect 13332 4367 13366 4401
rect 16649 4437 16683 4471
rect 13436 4333 13470 4367
rect 13505 4333 13539 4367
rect 13574 4333 13608 4367
rect 13643 4333 13677 4367
rect 13712 4333 13746 4367
rect 13781 4333 13815 4367
rect 13850 4333 13884 4367
rect 13919 4333 13953 4367
rect 13988 4333 14022 4367
rect 14057 4333 14091 4367
rect 14126 4333 14160 4367
rect 14195 4333 14229 4367
rect 14264 4333 14298 4367
rect 14333 4333 14367 4367
rect 14402 4333 14436 4367
rect 14471 4333 14505 4367
rect 14540 4333 14574 4367
rect 14609 4333 14643 4367
rect 14678 4333 14712 4367
rect 14747 4333 14781 4367
rect 14816 4333 14850 4367
rect 14885 4333 14919 4367
rect 14954 4333 14988 4367
rect 15023 4333 15057 4367
rect 15092 4333 15126 4367
rect 15161 4333 15195 4367
rect 15230 4333 15264 4367
rect 15299 4333 15333 4367
rect 15368 4333 15402 4367
rect 15437 4333 15471 4367
rect 15506 4333 15540 4367
rect 15575 4333 15609 4367
rect 15644 4333 15678 4367
rect 15713 4333 15747 4367
rect 15782 4333 15816 4367
rect 15851 4333 15885 4367
rect 15920 4333 15954 4367
rect 15989 4333 16023 4367
rect 16058 4333 16092 4367
rect 16127 4333 16161 4367
rect 16196 4333 16230 4367
rect 16265 4333 16299 4367
rect 16335 4333 16369 4367
rect 16405 4333 16439 4367
rect 16475 4333 16509 4367
rect 16545 4333 16579 4367
rect 16615 4333 16649 4367
<< poly >>
rect 314 5743 1238 5765
rect 314 5709 330 5743
rect 364 5709 398 5743
rect 432 5709 466 5743
rect 500 5709 1238 5743
rect 314 5693 1238 5709
rect 514 5625 714 5651
rect 838 5625 1038 5651
rect 514 5515 714 5541
rect 380 5493 714 5515
rect 380 5459 396 5493
rect 430 5459 464 5493
rect 498 5472 714 5493
rect 838 5515 1038 5541
rect 838 5493 1172 5515
rect 838 5472 1054 5493
rect 498 5459 565 5472
rect 380 5443 565 5459
rect 987 5459 1054 5472
rect 1088 5459 1122 5493
rect 1156 5459 1172 5493
rect 987 5443 1172 5459
rect 1994 5482 2060 5498
rect 1994 5448 2010 5482
rect 2044 5448 2060 5482
rect 607 5414 748 5430
rect 607 5401 623 5414
rect 492 5380 623 5401
rect 657 5380 691 5414
rect 725 5380 748 5414
rect 492 5364 748 5380
rect 492 5358 592 5364
rect 648 5358 748 5364
rect 804 5414 945 5430
rect 1994 5429 2060 5448
rect 804 5380 827 5414
rect 861 5380 895 5414
rect 929 5401 945 5414
rect 1428 5414 2060 5429
rect 929 5380 1060 5401
rect 804 5364 1060 5380
rect 804 5358 904 5364
rect 960 5358 1060 5364
rect 1428 5380 2010 5414
rect 2044 5380 2060 5414
rect 1428 5364 2060 5380
rect 1428 5358 1528 5364
rect 1584 5358 1684 5364
rect 1740 5358 1840 5364
rect 1896 5358 1996 5364
rect 2815 4979 2881 4995
rect 2815 4945 2831 4979
rect 2865 4945 2881 4979
rect 2815 4911 2881 4945
rect 2815 4877 2831 4911
rect 2865 4877 2881 4911
rect 2815 4843 2881 4877
rect 2815 4809 2831 4843
rect 2865 4809 2881 4843
rect 2815 4775 2881 4809
rect 2815 4741 2831 4775
rect 2865 4741 2881 4775
rect 2815 4707 2881 4741
rect 180 4694 280 4706
rect 139 4688 280 4694
rect 336 4688 436 4706
rect 1116 4688 1216 4706
rect 1272 4688 1372 4706
rect 139 4678 436 4688
rect 139 4644 155 4678
rect 189 4644 223 4678
rect 257 4644 436 4678
rect 139 4628 436 4644
rect 1099 4672 1372 4688
rect 1099 4638 1115 4672
rect 1149 4638 1183 4672
rect 1217 4638 1372 4672
rect 1099 4622 1372 4638
rect 2815 4673 2831 4707
rect 2865 4673 2881 4707
rect 2815 4639 2881 4673
rect 2815 4605 2831 4639
rect 2865 4605 2881 4639
rect 2815 4571 2881 4605
rect 281 4530 381 4546
rect 281 4496 304 4530
rect 338 4506 381 4530
rect 859 4530 959 4546
rect 338 4496 537 4506
rect 281 4462 537 4496
rect 281 4428 304 4462
rect 338 4428 537 4462
rect 281 4406 537 4428
rect 859 4496 909 4530
rect 943 4496 959 4530
rect 1171 4530 1271 4546
rect 1171 4506 1214 4530
rect 859 4462 959 4496
rect 859 4428 909 4462
rect 943 4428 959 4462
rect 859 4406 959 4428
rect 1015 4496 1214 4506
rect 1248 4496 1271 4530
rect 1015 4462 1271 4496
rect 1015 4428 1214 4462
rect 1248 4428 1271 4462
rect 1015 4406 1271 4428
rect 1327 4530 1427 4546
rect 1327 4496 1343 4530
rect 1377 4496 1427 4530
rect 1327 4462 1427 4496
rect 2815 4537 2831 4571
rect 2865 4537 2881 4571
rect 2815 4502 2881 4537
rect 1327 4428 1343 4462
rect 1377 4428 1427 4462
rect 1593 4462 1812 4478
rect 1327 4406 1427 4428
rect 1593 4428 1694 4462
rect 1728 4428 1762 4462
rect 1796 4428 1812 4462
rect 1593 4412 1812 4428
rect 2163 4462 2393 4478
rect 2163 4428 2179 4462
rect 2213 4428 2247 4462
rect 2281 4428 2393 4462
rect 2163 4412 2393 4428
rect 1593 4406 1713 4412
rect 2273 4406 2393 4412
rect 2815 4468 2831 4502
rect 2865 4468 2881 4502
rect 2815 4433 2881 4468
rect 2815 4399 2831 4433
rect 2865 4399 2881 4433
rect 1936 4311 2008 4327
rect 1936 4277 1958 4311
rect 1992 4277 2008 4311
rect 1936 4243 2008 4277
rect 1936 4209 1958 4243
rect 1992 4209 2008 4243
rect 1936 4127 2008 4209
rect 2815 4364 2881 4399
rect 2815 4330 2831 4364
rect 2865 4330 2881 4364
rect 2815 4295 2881 4330
rect 2815 4261 2831 4295
rect 2865 4261 2881 4295
rect 2815 4226 2881 4261
rect 2815 4192 2831 4226
rect 2865 4192 2881 4226
rect 2815 4157 2881 4192
rect 1800 3927 1826 4127
rect 1910 4079 2008 4127
rect 1910 3927 1936 4079
rect 2050 4037 2076 4127
rect 1978 4021 2076 4037
rect 1978 3987 1994 4021
rect 2028 3987 2076 4021
rect 1978 3953 2076 3987
rect 1978 3919 1994 3953
rect 2028 3927 2076 3953
rect 2160 3927 2186 4127
rect 2815 4123 2831 4157
rect 2865 4123 2881 4157
rect 2815 4088 2881 4123
rect 2815 4054 2831 4088
rect 2865 4054 2881 4088
rect 2815 4019 2881 4054
rect 2815 3985 2831 4019
rect 2865 3985 2881 4019
rect 2815 3950 2881 3985
rect 2028 3919 2050 3927
rect 1978 3903 2050 3919
rect 2815 3916 2831 3950
rect 2865 3916 2881 3950
rect 2815 3881 2881 3916
rect 2815 3847 2831 3881
rect 2865 3847 2881 3881
rect 2815 3812 2881 3847
rect 2815 3778 2831 3812
rect 2865 3778 2881 3812
rect 125 3748 225 3754
rect 91 3732 225 3748
rect 91 3698 107 3732
rect 141 3698 175 3732
rect 209 3698 225 3732
rect 91 3682 225 3698
rect 593 3748 693 3754
rect 593 3732 727 3748
rect 593 3698 609 3732
rect 643 3698 677 3732
rect 711 3698 727 3732
rect 2815 3743 2881 3778
rect 593 3682 727 3698
rect 1201 3646 1227 3712
rect 2367 3646 2393 3712
rect 2815 3709 2831 3743
rect 2865 3709 2881 3743
rect 2815 3693 2881 3709
rect 4219 4979 4285 4995
rect 4219 4945 4235 4979
rect 4269 4945 4285 4979
rect 4219 4911 4285 4945
rect 4219 4877 4235 4911
rect 4269 4877 4285 4911
rect 4219 4843 4285 4877
rect 4219 4809 4235 4843
rect 4269 4809 4285 4843
rect 4219 4775 4285 4809
rect 4219 4741 4235 4775
rect 4269 4741 4285 4775
rect 4219 4707 4285 4741
rect 4219 4673 4235 4707
rect 4269 4673 4285 4707
rect 4219 4639 4285 4673
rect 4219 4605 4235 4639
rect 4269 4605 4285 4639
rect 4219 4571 4285 4605
rect 4219 4537 4235 4571
rect 4269 4537 4285 4571
rect 4219 4502 4285 4537
rect 4219 4468 4235 4502
rect 4269 4468 4285 4502
rect 4219 4433 4285 4468
rect 4219 4399 4235 4433
rect 4269 4399 4285 4433
rect 4219 4364 4285 4399
rect 4219 4330 4235 4364
rect 4269 4330 4285 4364
rect 4219 4295 4285 4330
rect 4219 4261 4235 4295
rect 4269 4261 4285 4295
rect 4219 4226 4285 4261
rect 4219 4192 4235 4226
rect 4269 4192 4285 4226
rect 4219 4157 4285 4192
rect 4219 4123 4235 4157
rect 4269 4123 4285 4157
rect 4219 4088 4285 4123
rect 4219 4054 4235 4088
rect 4269 4054 4285 4088
rect 4219 4019 4285 4054
rect 4219 3985 4235 4019
rect 4269 3985 4285 4019
rect 4219 3950 4285 3985
rect 4219 3916 4235 3950
rect 4269 3916 4285 3950
rect 4219 3881 4285 3916
rect 4219 3847 4235 3881
rect 4269 3847 4285 3881
rect 4219 3812 4285 3847
rect 4219 3778 4235 3812
rect 4269 3778 4285 3812
rect 13434 6243 13500 6259
rect 13434 6209 13450 6243
rect 13484 6242 13500 6243
rect 13484 6209 13509 6242
rect 13434 6169 13509 6209
rect 13434 6135 13450 6169
rect 13484 6142 13509 6169
rect 13484 6135 13500 6142
rect 13434 6094 13500 6135
rect 13434 6060 13450 6094
rect 13484 6086 13500 6094
rect 13484 6060 13509 6086
rect 13434 6019 13509 6060
rect 13434 5985 13450 6019
rect 13484 5986 13509 6019
rect 13484 5985 13500 5986
rect 13434 5969 13500 5985
rect 13434 5739 13500 5755
rect 13434 5705 13450 5739
rect 13484 5738 13500 5739
rect 13484 5705 13509 5738
rect 13434 5665 13509 5705
rect 13434 5631 13450 5665
rect 13484 5638 13509 5665
rect 13484 5631 13500 5638
rect 13434 5590 13500 5631
rect 13434 5556 13450 5590
rect 13484 5582 13500 5590
rect 13484 5556 13509 5582
rect 13434 5515 13509 5556
rect 13434 5481 13450 5515
rect 13484 5482 13509 5515
rect 13484 5481 13500 5482
rect 13434 5465 13500 5481
rect 13434 5235 13500 5251
rect 13434 5201 13450 5235
rect 13484 5234 13500 5235
rect 13484 5201 13509 5234
rect 13434 5161 13509 5201
rect 13434 5127 13450 5161
rect 13484 5134 13509 5161
rect 13484 5127 13500 5134
rect 13434 5086 13500 5127
rect 13434 5052 13450 5086
rect 13484 5078 13500 5086
rect 13484 5052 13509 5078
rect 13434 5011 13509 5052
rect 13434 4977 13450 5011
rect 13484 4978 13509 5011
rect 13484 4977 13500 4978
rect 13434 4961 13500 4977
rect 13434 4731 13500 4747
rect 13434 4697 13450 4731
rect 13484 4730 13500 4731
rect 13484 4697 13509 4730
rect 13434 4657 13509 4697
rect 13434 4623 13450 4657
rect 13484 4630 13509 4657
rect 13484 4623 13500 4630
rect 13434 4582 13500 4623
rect 13434 4548 13450 4582
rect 13484 4574 13500 4582
rect 13484 4548 13509 4574
rect 13434 4507 13509 4548
rect 13434 4473 13450 4507
rect 13484 4474 13509 4507
rect 13484 4473 13500 4474
rect 13434 4457 13500 4473
rect 4219 3743 4285 3778
rect 4219 3709 4235 3743
rect 4269 3709 4285 3743
rect 4219 3693 4285 3709
rect 1201 3640 1301 3646
rect 1357 3640 1457 3646
rect 1513 3640 1613 3646
rect 1669 3640 1769 3646
rect 1825 3640 1925 3646
rect 1981 3640 2081 3646
rect 2137 3640 2237 3646
rect 2293 3640 2393 3646
rect 46 184 122 3508
rect 546 1908 554 3508
rect 546 184 554 1784
<< polycont >>
rect 330 5709 364 5743
rect 398 5709 432 5743
rect 466 5709 500 5743
rect 396 5459 430 5493
rect 464 5459 498 5493
rect 1054 5459 1088 5493
rect 1122 5459 1156 5493
rect 2010 5448 2044 5482
rect 623 5380 657 5414
rect 691 5380 725 5414
rect 827 5380 861 5414
rect 895 5380 929 5414
rect 2010 5380 2044 5414
rect 2831 4945 2865 4979
rect 2831 4877 2865 4911
rect 2831 4809 2865 4843
rect 2831 4741 2865 4775
rect 155 4644 189 4678
rect 223 4644 257 4678
rect 1115 4638 1149 4672
rect 1183 4638 1217 4672
rect 2831 4673 2865 4707
rect 2831 4605 2865 4639
rect 304 4496 338 4530
rect 304 4428 338 4462
rect 909 4496 943 4530
rect 909 4428 943 4462
rect 1214 4496 1248 4530
rect 1214 4428 1248 4462
rect 1343 4496 1377 4530
rect 2831 4537 2865 4571
rect 1343 4428 1377 4462
rect 1694 4428 1728 4462
rect 1762 4428 1796 4462
rect 2179 4428 2213 4462
rect 2247 4428 2281 4462
rect 2831 4468 2865 4502
rect 2831 4399 2865 4433
rect 1958 4277 1992 4311
rect 1958 4209 1992 4243
rect 2831 4330 2865 4364
rect 2831 4261 2865 4295
rect 2831 4192 2865 4226
rect 1994 3987 2028 4021
rect 1994 3919 2028 3953
rect 2831 4123 2865 4157
rect 2831 4054 2865 4088
rect 2831 3985 2865 4019
rect 2831 3916 2865 3950
rect 2831 3847 2865 3881
rect 2831 3778 2865 3812
rect 107 3698 141 3732
rect 175 3698 209 3732
rect 609 3698 643 3732
rect 677 3698 711 3732
rect 2831 3709 2865 3743
rect 4235 4945 4269 4979
rect 4235 4877 4269 4911
rect 4235 4809 4269 4843
rect 4235 4741 4269 4775
rect 4235 4673 4269 4707
rect 4235 4605 4269 4639
rect 4235 4537 4269 4571
rect 4235 4468 4269 4502
rect 4235 4399 4269 4433
rect 4235 4330 4269 4364
rect 4235 4261 4269 4295
rect 4235 4192 4269 4226
rect 4235 4123 4269 4157
rect 4235 4054 4269 4088
rect 4235 3985 4269 4019
rect 4235 3916 4269 3950
rect 4235 3847 4269 3881
rect 4235 3778 4269 3812
rect 13450 6209 13484 6243
rect 13450 6135 13484 6169
rect 13450 6060 13484 6094
rect 13450 5985 13484 6019
rect 13450 5705 13484 5739
rect 13450 5631 13484 5665
rect 13450 5556 13484 5590
rect 13450 5481 13484 5515
rect 13450 5201 13484 5235
rect 13450 5127 13484 5161
rect 13450 5052 13484 5086
rect 13450 4977 13484 5011
rect 13450 4697 13484 4731
rect 13450 4623 13484 4657
rect 13450 4548 13484 4582
rect 13450 4473 13484 4507
rect 4235 3709 4269 3743
<< locali >>
rect 2315 8153 2355 8165
rect 2315 8119 2318 8153
rect 2352 8119 2355 8153
rect 2315 8081 2355 8119
rect 2315 8047 2318 8081
rect 2352 8047 2355 8081
rect 0 7995 83 8007
rect 0 7961 49 7995
rect 0 7923 83 7961
rect 0 7889 49 7923
rect 0 4546 40 7889
rect 2241 7461 2275 7499
rect 299 7231 333 7277
rect 265 7219 333 7231
rect 761 7219 795 7277
rect 1047 7219 1081 7277
rect 1427 7219 1461 7277
rect 2241 7219 2275 7277
rect 265 7021 299 7219
rect 265 6987 279 7021
rect 383 6953 421 6987
rect 201 5837 269 5853
rect 235 5803 269 5837
rect 201 5787 269 5803
rect 303 5787 677 5853
rect 314 5709 325 5743
rect 364 5709 397 5743
rect 432 5709 466 5743
rect 503 5709 516 5743
rect 201 5587 303 5603
rect 235 5553 269 5587
rect 201 5537 303 5553
rect 135 5248 169 5286
rect 135 5176 169 5214
rect 203 5089 257 5537
rect 396 5493 563 5509
rect 430 5459 464 5493
rect 498 5459 563 5493
rect 396 5443 563 5459
rect 447 5248 481 5286
rect 447 5176 481 5214
rect 203 5055 213 5089
rect 247 5055 257 5089
rect 203 5017 257 5055
rect 203 4983 213 5017
rect 247 4983 257 5017
rect 203 4971 257 4983
rect 288 4802 322 4840
rect 529 4694 563 5443
rect 623 5430 677 5787
rect 725 5587 827 5965
rect 759 5553 793 5587
rect 725 5537 827 5553
rect 875 5787 1249 5853
rect 1283 5837 1351 5853
rect 1283 5803 1317 5837
rect 1283 5787 1351 5803
rect 623 5414 725 5430
rect 657 5380 691 5414
rect 623 5364 725 5380
rect 603 5017 637 5055
rect 146 4678 257 4694
rect 189 4644 218 4678
rect 146 4628 257 4644
rect 474 4660 563 4694
rect 372 4608 426 4624
rect 372 4574 381 4608
rect 415 4574 426 4608
rect 0 4530 338 4546
rect 0 4506 304 4530
rect 304 4462 338 4496
rect 304 4412 338 4428
rect 372 4536 426 4574
rect 372 4502 381 4536
rect 415 4502 426 4536
rect 80 3898 114 3936
rect 80 3826 114 3864
rect 372 3776 426 4502
rect 474 4309 508 4660
rect 474 4237 508 4275
rect 474 4056 508 4094
rect 91 3698 107 3732
rect 141 3698 175 3732
rect 209 3698 225 3732
rect 91 3678 225 3698
rect 259 3678 297 3712
rect 474 3553 508 4022
rect 677 3776 725 5364
rect 759 5320 793 5537
rect 875 5430 929 5787
rect 1249 5587 1351 5603
rect 1283 5553 1317 5587
rect 1249 5537 1351 5553
rect 759 5248 793 5286
rect 759 5176 793 5214
rect 827 5414 929 5430
rect 861 5380 895 5414
rect 827 5364 929 5380
rect 989 5493 1156 5509
rect 989 5459 1054 5493
rect 1088 5459 1122 5493
rect 989 5443 1156 5459
rect 759 4678 793 4728
rect 759 4628 793 4644
rect 827 4262 870 5364
rect 915 5017 949 5055
rect 989 4694 1023 5443
rect 1071 5248 1105 5286
rect 1071 5176 1105 5214
rect 1295 5089 1349 5537
rect 1994 5448 2010 5482
rect 2044 5448 2060 5482
rect 1994 5414 2060 5448
rect 1994 5380 2010 5414
rect 2044 5380 2060 5414
rect 1383 5248 1417 5286
rect 1383 5176 1417 5214
rect 1695 5248 1729 5286
rect 1695 5176 1729 5214
rect 2007 5248 2041 5286
rect 2007 5176 2041 5214
rect 1295 5055 1305 5089
rect 1339 5055 1349 5089
rect 1295 5017 1349 5055
rect 1295 4983 1305 5017
rect 1339 4983 1349 5017
rect 1295 4971 1349 4983
rect 1768 4961 1802 4999
rect 1227 4803 1261 4841
rect 1539 4803 1573 4841
rect 989 4660 1078 4694
rect 938 4564 976 4598
rect 909 4530 943 4564
rect 909 4462 943 4496
rect 909 4412 943 4428
rect 1044 4369 1078 4660
rect 1115 4678 1226 4688
rect 1149 4672 1187 4678
rect 1149 4638 1183 4672
rect 1221 4644 1226 4678
rect 1217 4638 1226 4644
rect 1115 4622 1226 4638
rect 1297 4564 1324 4598
rect 1358 4564 1396 4598
rect 1214 4542 1248 4546
rect 1176 4508 1214 4542
rect 1214 4462 1248 4496
rect 1214 4412 1248 4428
rect 1343 4530 1377 4564
rect 1343 4462 1377 4496
rect 1438 4488 1505 4504
rect 1438 4428 1471 4488
rect 1343 4412 1377 4428
rect 1044 4297 1078 4335
rect 827 3776 868 4262
rect 902 4112 936 4150
rect 593 3712 609 3732
rect 593 3678 605 3712
rect 643 3698 677 3732
rect 639 3678 677 3698
rect 711 3678 727 3732
rect 902 3553 936 4078
rect 1438 3970 1505 4380
rect 1472 3936 1505 3970
rect 1438 3898 1505 3936
rect 1472 3864 1505 3898
rect 1438 3826 1505 3864
rect 1472 3792 1505 3826
rect 1438 3776 1505 3792
rect 1539 3776 1573 4728
rect 1619 4564 1628 4598
rect 1662 4564 1700 4598
rect 1126 3706 1160 3776
rect 1619 3696 1659 4564
rect 1768 4478 1802 4927
rect 2089 5017 2123 5055
rect 1851 4803 1885 4841
rect 2089 4478 2123 4983
rect 2163 4598 2203 5471
rect 2237 5248 2271 5286
rect 2237 5176 2271 5214
rect 2197 4564 2235 4598
rect 2315 4592 2355 8047
rect 2349 4558 2355 4592
rect 2315 4520 2355 4558
rect 2349 4486 2355 4520
rect 2392 7895 2432 7907
rect 2392 7861 2395 7895
rect 2429 7861 2432 7895
rect 2392 7823 2432 7861
rect 2392 7789 2395 7823
rect 2429 7789 2432 7823
rect 1694 4462 1888 4478
rect 1728 4428 1762 4462
rect 1796 4428 1888 4462
rect 1694 4412 1888 4428
rect 2089 4462 2281 4478
rect 2089 4428 2179 4462
rect 2213 4428 2247 4462
rect 2392 4452 2432 7789
rect 3050 7732 3198 7766
rect 3232 7732 3250 7766
rect 3050 7694 3250 7732
rect 3050 7660 3198 7694
rect 3232 7660 3250 7694
rect 3080 7573 3118 7607
rect 3534 7606 3572 7640
rect 3606 7606 3644 7640
rect 3304 7107 3402 7234
rect 3304 7073 3368 7107
rect 3304 7035 3402 7073
rect 3304 7001 3368 7035
rect 3304 6963 3402 7001
rect 3304 6929 3368 6963
rect 12629 7081 12697 7086
rect 12629 7047 12643 7081
rect 12677 7047 12697 7081
rect 17219 7052 17253 7086
rect 17287 7052 17386 7086
rect 12629 6984 12697 7047
rect 17219 7018 17386 7052
rect 17219 6984 17284 7018
rect 12629 6955 12765 6984
rect 17151 6969 17284 6984
rect 17151 6955 17218 6969
rect 12629 6954 12643 6955
rect 12677 6921 12716 6955
rect 12750 6921 12765 6955
rect 17159 6950 17218 6955
rect 17252 6950 17284 6969
rect 17159 6921 17216 6950
rect 12663 6920 12765 6921
rect 12629 6916 12765 6920
rect 17151 6916 17216 6921
rect 12629 6886 12799 6916
rect 12731 6870 12799 6886
rect 12731 6836 12760 6870
rect 12794 6836 12799 6870
rect 12731 6818 12799 6836
rect 2842 6733 3318 6739
rect 2842 6699 2849 6733
rect 2883 6699 3318 6733
rect 2842 6685 3318 6699
rect 2842 6661 2908 6685
rect 2842 6627 2849 6661
rect 2883 6627 2908 6661
rect 2842 6589 2908 6627
rect 2992 6617 3014 6651
rect 3060 6617 3086 6651
rect 3120 6617 3162 6651
rect 3460 6623 3498 6657
rect 3532 6623 3570 6657
rect 3604 6623 3642 6657
rect 2842 6555 2849 6589
rect 2883 6555 2908 6589
rect 2842 6549 2908 6555
rect 3409 6549 3447 6583
rect 3375 6532 3481 6549
rect 2849 6406 2883 6444
rect 2879 5122 2895 5156
rect 2929 5122 2964 5156
rect 2998 5122 3033 5156
rect 3067 5122 3102 5156
rect 3136 5122 3171 5156
rect 3232 5146 3240 5156
rect 3205 5122 3240 5146
rect 3274 5122 3309 5156
rect 3343 5122 3378 5156
rect 3412 5122 3447 5156
rect 3481 5122 3516 5156
rect 3550 5122 3585 5156
rect 3619 5122 3654 5156
rect 3688 5122 3723 5156
rect 3757 5122 3792 5156
rect 3826 5122 3861 5156
rect 3895 5122 3930 5156
rect 3964 5122 3999 5156
rect 4033 5122 4069 5156
rect 4103 5122 4139 5156
rect 4173 5122 4189 5156
rect 3198 5108 3232 5122
rect 3008 5006 3046 5040
rect 3080 5006 3118 5040
rect 3747 5006 3796 5040
rect 3830 5006 3879 5040
rect 3913 5006 3962 5040
rect 3996 5006 4045 5040
rect 4079 5006 4127 5040
rect 2089 4412 2281 4428
rect 2327 4412 2432 4452
rect 2831 4979 2865 4995
rect 2831 4911 2865 4945
rect 4235 4979 4269 4995
rect 4235 4911 4269 4945
rect 2831 4843 2865 4877
rect 3507 4850 3659 4884
rect 3693 4850 3798 4884
rect 2831 4775 2865 4809
rect 2831 4707 2865 4741
rect 4235 4843 4269 4877
rect 4235 4775 4269 4809
rect 3008 4694 3046 4728
rect 3080 4694 3118 4728
rect 3747 4694 3796 4728
rect 3830 4694 3879 4728
rect 3913 4694 3962 4728
rect 3996 4694 4045 4728
rect 4079 4694 4127 4728
rect 4235 4708 4269 4741
rect 2831 4667 2837 4673
rect 2831 4639 2871 4667
rect 2865 4627 2871 4639
rect 4235 4639 4269 4673
rect 2831 4593 2837 4605
rect 2831 4571 2871 4593
rect 3008 4584 3046 4618
rect 3080 4584 3118 4618
rect 3946 4584 4020 4618
rect 4054 4584 4127 4618
rect 4235 4591 4269 4605
rect 2865 4552 2871 4571
rect 2831 4518 2837 4537
rect 2831 4502 2871 4518
rect 2865 4477 2871 4502
rect 2831 4443 2837 4468
rect 4235 4502 4269 4537
rect 2831 4433 2871 4443
rect 1822 4372 1888 4412
rect 1822 4369 1838 4372
rect 1822 4335 1832 4369
rect 1872 4338 1888 4372
rect 1866 4335 1888 4338
rect 1822 4297 1888 4335
rect 2026 4369 2060 4375
rect 1822 4263 1832 4297
rect 1866 4263 1888 4297
rect 1822 4245 1888 4263
rect 1926 4311 1992 4327
rect 1926 4309 1958 4311
rect 1960 4275 1992 4277
rect 1926 4243 1992 4275
rect 1926 4237 1958 4243
rect 1960 4203 1992 4209
rect 1926 4193 1992 4203
rect 2026 4297 2060 4335
rect 1770 4016 1808 4050
rect 2026 4037 2060 4263
rect 2098 4372 2164 4412
rect 2098 4338 2114 4372
rect 2148 4338 2164 4372
rect 2098 4309 2164 4338
rect 2098 4275 2114 4309
rect 2148 4275 2164 4309
rect 2098 4237 2164 4275
rect 2098 4203 2114 4237
rect 2148 4203 2164 4237
rect 2098 4191 2164 4203
rect 2178 4113 2216 4147
rect 1994 4021 2060 4037
rect 2028 3987 2060 4021
rect 1994 3953 2060 3987
rect 2028 3919 2060 3953
rect 1822 3882 1838 3916
rect 1872 3882 1888 3916
rect 1994 3903 2060 3919
rect 1822 3869 1888 3882
rect 2098 3882 2114 3916
rect 2148 3882 2164 3916
rect 2098 3869 2164 3882
rect 1822 3835 1832 3869
rect 1866 3835 1904 3869
rect 1938 3835 1976 3869
rect 2010 3835 2048 3869
rect 2082 3835 2120 3869
rect 2154 3835 2164 3869
rect 2327 3696 2367 4412
rect 2865 4402 2871 4433
rect 3507 4428 3654 4462
rect 3688 4428 3726 4462
rect 3760 4428 3798 4462
rect 4235 4433 4269 4468
rect 2831 4368 2837 4399
rect 2831 4364 2871 4368
rect 2865 4330 2871 4364
rect 2831 4327 2871 4330
rect 2831 4295 2837 4327
rect 2865 4261 2871 4293
rect 3008 4272 3046 4306
rect 3080 4272 3118 4306
rect 2831 4252 2871 4261
rect 2831 4226 2837 4252
rect 2865 4192 2871 4218
rect 2831 4177 2871 4192
rect 2831 4157 2837 4177
rect 3541 4150 3625 4428
rect 4235 4364 4269 4399
rect 3946 4272 4020 4306
rect 4054 4272 4127 4306
rect 4235 4295 4269 4303
rect 4235 4226 4269 4227
rect 4235 4185 4269 4192
rect 2865 4123 2871 4143
rect 2831 4102 2871 4123
rect 3507 4116 3654 4150
rect 3688 4116 3726 4150
rect 3760 4116 3798 4150
rect 2831 4088 2837 4102
rect 2865 4054 2871 4068
rect 2831 4027 2871 4054
rect 2831 4019 2837 4027
rect 2865 3985 2871 3993
rect 2831 3952 2871 3985
rect 3008 3960 3046 3994
rect 3080 3960 3118 3994
rect 2831 3950 2837 3952
rect 2865 3916 2871 3918
rect 2831 3881 2871 3916
rect 2865 3877 2871 3881
rect 2831 3843 2837 3847
rect 2831 3812 2871 3843
rect 3541 3838 3625 4116
rect 4235 4109 4269 4123
rect 4235 4033 4269 4054
rect 3946 3960 4020 3994
rect 4054 3960 4127 3994
rect 4235 3957 4269 3985
rect 4235 3881 4269 3916
rect 2865 3802 2871 3812
rect 3507 3804 3654 3838
rect 3688 3804 3726 3838
rect 3760 3804 3798 3838
rect 4235 3812 4269 3847
rect 1126 3634 1160 3672
rect 2404 3628 2438 3776
rect 2831 3768 2837 3778
rect 2831 3743 2871 3768
rect 2865 3727 2871 3743
rect 2831 3693 2837 3709
rect 13030 6685 16986 6686
rect 13030 6651 13038 6685
rect 13072 6662 13111 6685
rect 13072 6651 13092 6662
rect 13145 6651 13184 6685
rect 13218 6651 13257 6685
rect 13291 6651 13330 6685
rect 13364 6651 13403 6685
rect 13437 6651 13476 6685
rect 13510 6651 13549 6685
rect 13583 6651 13622 6685
rect 13656 6651 13695 6685
rect 13729 6651 13768 6685
rect 13802 6651 13841 6685
rect 13875 6651 13914 6685
rect 13948 6651 13987 6685
rect 14021 6651 14060 6685
rect 14094 6651 14133 6685
rect 14167 6651 14206 6685
rect 14240 6651 14279 6685
rect 14313 6651 14352 6685
rect 14386 6651 14425 6685
rect 14459 6651 14497 6685
rect 14531 6651 14569 6685
rect 14603 6651 14641 6685
rect 14675 6651 14713 6685
rect 14747 6651 14785 6685
rect 14819 6651 14857 6685
rect 14891 6651 14929 6685
rect 14963 6651 15001 6685
rect 15035 6651 15073 6685
rect 15107 6651 15145 6685
rect 15179 6651 15217 6685
rect 15251 6651 15289 6685
rect 15323 6651 15361 6685
rect 15395 6651 15433 6685
rect 15467 6651 15505 6685
rect 15539 6651 15577 6685
rect 15611 6651 15649 6685
rect 15683 6651 15721 6685
rect 15755 6651 15793 6685
rect 15827 6651 15865 6685
rect 15899 6651 15937 6685
rect 15971 6651 16009 6685
rect 16043 6651 16081 6685
rect 16115 6651 16153 6685
rect 16187 6651 16225 6685
rect 16259 6651 16297 6685
rect 16331 6651 16369 6685
rect 16403 6651 16441 6685
rect 16475 6651 16513 6685
rect 16547 6651 16585 6685
rect 16619 6651 16657 6685
rect 16691 6651 16729 6685
rect 16763 6651 16801 6685
rect 16835 6651 16873 6685
rect 16907 6661 16945 6685
rect 16934 6651 16945 6661
rect 16979 6651 16986 6685
rect 13030 6628 13092 6651
rect 13126 6628 16900 6651
rect 13030 6627 16900 6628
rect 16934 6627 16986 6651
rect 13030 6594 16986 6627
rect 13030 6571 13065 6594
rect 13099 6593 16986 6594
rect 13099 6571 16927 6593
rect 16961 6571 16986 6593
rect 13030 6537 13038 6571
rect 13099 6560 13111 6571
rect 13072 6537 13111 6560
rect 13145 6537 13184 6571
rect 13218 6537 13257 6571
rect 13291 6537 13330 6571
rect 13364 6537 13403 6571
rect 13437 6537 13476 6571
rect 13510 6537 13549 6571
rect 13583 6537 13622 6571
rect 13656 6537 13695 6571
rect 13729 6537 13768 6571
rect 13802 6537 13841 6571
rect 13875 6537 13914 6571
rect 13948 6537 13987 6571
rect 14021 6537 14060 6571
rect 14094 6537 14133 6571
rect 14167 6537 14206 6571
rect 14240 6537 14279 6571
rect 14313 6537 14352 6571
rect 14386 6537 14425 6571
rect 14459 6537 14497 6571
rect 14531 6537 14569 6571
rect 14603 6537 14641 6571
rect 14675 6537 14713 6571
rect 14747 6537 14785 6571
rect 14819 6537 14857 6571
rect 14891 6537 14929 6571
rect 14963 6537 15001 6571
rect 15035 6537 15073 6571
rect 15107 6537 15145 6571
rect 15179 6537 15217 6571
rect 15251 6537 15289 6571
rect 15323 6537 15361 6571
rect 15395 6537 15433 6571
rect 15467 6537 15505 6571
rect 15539 6537 15577 6571
rect 15611 6537 15649 6571
rect 15683 6537 15721 6571
rect 15755 6537 15793 6571
rect 15827 6537 15865 6571
rect 15899 6537 15937 6571
rect 15971 6537 16009 6571
rect 16043 6537 16081 6571
rect 16115 6537 16153 6571
rect 16187 6537 16225 6571
rect 16259 6537 16297 6571
rect 16331 6537 16369 6571
rect 16403 6537 16441 6571
rect 16475 6537 16513 6571
rect 16547 6537 16585 6571
rect 16619 6537 16657 6571
rect 16691 6537 16729 6571
rect 16763 6537 16801 6571
rect 16835 6537 16873 6571
rect 16907 6559 16927 6571
rect 16907 6537 16945 6559
rect 16979 6537 16986 6571
rect 13030 6536 16986 6537
rect 13030 6490 13180 6536
rect 13030 6456 13032 6490
rect 13066 6456 13146 6490
rect 13030 6418 13180 6456
rect 13030 6384 13032 6418
rect 13066 6384 13146 6418
rect 16835 6490 16986 6536
rect 16835 6456 16837 6490
rect 16871 6456 16951 6490
rect 16985 6456 16986 6490
rect 16835 6418 16986 6456
rect 13030 6346 13180 6384
rect 13030 6312 13032 6346
rect 13066 6312 13146 6346
rect 13030 6274 13180 6312
rect 13030 6240 13032 6274
rect 13066 6240 13146 6274
rect 13030 6202 13180 6240
rect 13030 6168 13032 6202
rect 13066 6168 13146 6202
rect 13030 6130 13180 6168
rect 13030 6096 13032 6130
rect 13066 6096 13146 6130
rect 13030 6058 13180 6096
rect 13030 6024 13032 6058
rect 13066 6024 13146 6058
rect 13030 5986 13180 6024
rect 13030 5952 13032 5986
rect 13066 5952 13146 5986
rect 13030 5914 13180 5952
rect 13030 5880 13032 5914
rect 13066 5880 13146 5914
rect 13030 5842 13180 5880
rect 13030 5808 13032 5842
rect 13066 5808 13146 5842
rect 13030 5770 13180 5808
rect 13030 5736 13032 5770
rect 13066 5736 13146 5770
rect 13030 5698 13180 5736
rect 13030 5664 13032 5698
rect 13066 5664 13146 5698
rect 13030 5626 13180 5664
rect 13030 5592 13032 5626
rect 13066 5592 13146 5626
rect 13030 5554 13180 5592
rect 13030 5520 13032 5554
rect 13066 5520 13146 5554
rect 13030 5482 13180 5520
rect 13030 5448 13032 5482
rect 13066 5448 13146 5482
rect 13030 5410 13180 5448
rect 13030 5376 13032 5410
rect 13066 5376 13146 5410
rect 13030 5338 13180 5376
rect 13030 5304 13032 5338
rect 13066 5304 13146 5338
rect 13030 5266 13180 5304
rect 13030 5232 13032 5266
rect 13066 5232 13146 5266
rect 13030 5194 13180 5232
rect 13030 5160 13032 5194
rect 13066 5160 13146 5194
rect 13030 5122 13180 5160
rect 13030 5088 13032 5122
rect 13066 5088 13146 5122
rect 13030 5050 13180 5088
rect 13030 5016 13032 5050
rect 13066 5016 13146 5050
rect 13030 4978 13180 5016
rect 13030 4944 13032 4978
rect 13066 4944 13146 4978
rect 13030 4906 13180 4944
rect 13030 4872 13032 4906
rect 13066 4872 13146 4906
rect 13030 4834 13180 4872
rect 13030 4800 13032 4834
rect 13066 4800 13146 4834
rect 13030 4762 13180 4800
rect 13030 4728 13032 4762
rect 13066 4728 13146 4762
rect 13030 4690 13180 4728
rect 13030 4656 13032 4690
rect 13066 4656 13146 4690
rect 13030 4618 13180 4656
rect 13030 4584 13032 4618
rect 13066 4584 13146 4618
rect 13030 4546 13180 4584
rect 13030 4512 13032 4546
rect 13066 4512 13146 4546
rect 13030 4474 13180 4512
rect 13030 4440 13032 4474
rect 13066 4440 13146 4474
rect 13030 4402 13180 4440
rect 13030 4368 13032 4402
rect 13066 4368 13146 4402
rect 13030 4330 13180 4368
rect 13332 6383 13404 6391
rect 13332 6319 13366 6383
rect 13400 6357 13404 6383
rect 13438 6383 13476 6391
rect 13438 6357 13474 6383
rect 13510 6357 13548 6391
rect 13582 6383 13620 6391
rect 13654 6383 13692 6391
rect 13726 6383 13764 6391
rect 13798 6383 13836 6391
rect 13870 6383 13908 6391
rect 13942 6383 13980 6391
rect 14014 6383 14052 6391
rect 14086 6383 14124 6391
rect 14158 6383 14196 6391
rect 14230 6383 14268 6391
rect 14302 6383 14340 6391
rect 14374 6383 14412 6391
rect 14446 6383 14484 6391
rect 14518 6383 14556 6391
rect 14590 6383 14628 6391
rect 14662 6383 14700 6391
rect 14734 6383 14772 6391
rect 14806 6383 14844 6391
rect 14878 6383 14916 6391
rect 14950 6383 14988 6391
rect 15022 6383 15060 6391
rect 15094 6383 15132 6391
rect 15166 6383 15204 6391
rect 15238 6383 15276 6391
rect 15310 6383 15348 6391
rect 15382 6383 15420 6391
rect 15454 6383 15492 6391
rect 15526 6383 15564 6391
rect 15598 6383 15636 6391
rect 15670 6383 15708 6391
rect 13590 6357 13620 6383
rect 13400 6349 13474 6357
rect 13508 6349 13556 6357
rect 13590 6349 13624 6357
rect 13658 6349 13692 6383
rect 13726 6349 13760 6383
rect 13798 6357 13828 6383
rect 13870 6357 13896 6383
rect 13942 6357 13964 6383
rect 14014 6357 14032 6383
rect 14086 6357 14100 6383
rect 14158 6357 14168 6383
rect 14230 6357 14236 6383
rect 14302 6357 14304 6383
rect 13794 6349 13828 6357
rect 13862 6349 13896 6357
rect 13930 6349 13964 6357
rect 13998 6349 14032 6357
rect 14066 6349 14100 6357
rect 14134 6349 14168 6357
rect 14202 6349 14236 6357
rect 14270 6349 14304 6357
rect 14338 6357 14340 6383
rect 14406 6357 14412 6383
rect 14474 6357 14484 6383
rect 14542 6357 14556 6383
rect 14610 6357 14628 6383
rect 14678 6357 14700 6383
rect 14746 6357 14772 6383
rect 14814 6357 14844 6383
rect 14338 6349 14372 6357
rect 14406 6349 14440 6357
rect 14474 6349 14508 6357
rect 14542 6349 14576 6357
rect 14610 6349 14644 6357
rect 14678 6349 14712 6357
rect 14746 6349 14780 6357
rect 14814 6349 14848 6357
rect 14882 6349 14916 6383
rect 14950 6349 14984 6383
rect 15022 6357 15053 6383
rect 15094 6357 15122 6383
rect 15166 6357 15191 6383
rect 15238 6357 15260 6383
rect 15310 6357 15329 6383
rect 15382 6357 15398 6383
rect 15454 6357 15467 6383
rect 15526 6357 15536 6383
rect 15598 6357 15605 6383
rect 15670 6357 15674 6383
rect 15018 6349 15053 6357
rect 15087 6349 15122 6357
rect 15156 6349 15191 6357
rect 15225 6349 15260 6357
rect 15294 6349 15329 6357
rect 15363 6349 15398 6357
rect 15432 6349 15467 6357
rect 15501 6349 15536 6357
rect 15570 6349 15605 6357
rect 15639 6349 15674 6357
rect 15742 6383 15780 6391
rect 15814 6383 15852 6391
rect 15886 6383 15924 6391
rect 15958 6383 15996 6391
rect 16030 6383 16068 6391
rect 16102 6383 16140 6391
rect 16174 6383 16213 6391
rect 16247 6383 16286 6391
rect 16320 6383 16359 6391
rect 16393 6383 16432 6391
rect 16466 6383 16505 6391
rect 15742 6357 15743 6383
rect 15708 6349 15743 6357
rect 15777 6357 15780 6383
rect 15846 6357 15852 6383
rect 15915 6357 15924 6383
rect 15984 6357 15996 6383
rect 16053 6357 16068 6383
rect 16122 6357 16140 6383
rect 16191 6357 16213 6383
rect 16260 6357 16286 6383
rect 16329 6357 16359 6383
rect 16398 6357 16432 6383
rect 15777 6349 15812 6357
rect 15846 6349 15881 6357
rect 15915 6349 15950 6357
rect 15984 6349 16019 6357
rect 16053 6349 16088 6357
rect 16122 6349 16157 6357
rect 16191 6349 16226 6357
rect 16260 6349 16295 6357
rect 16329 6349 16364 6357
rect 16398 6349 16433 6357
rect 16467 6349 16502 6383
rect 16539 6357 16578 6391
rect 16612 6357 16684 6391
rect 16536 6349 16684 6357
rect 16683 6319 16684 6349
rect 13332 6279 13366 6285
rect 13332 6210 13366 6212
rect 13332 6173 13366 6176
rect 13332 6100 13366 6107
rect 13332 6027 13366 6038
rect 13450 6247 13484 6259
rect 13564 6253 13603 6287
rect 13637 6253 13676 6287
rect 13710 6253 13749 6287
rect 13783 6253 13822 6287
rect 13856 6253 13895 6287
rect 13929 6253 13968 6287
rect 14002 6253 14041 6287
rect 14075 6253 14114 6287
rect 14148 6253 14187 6287
rect 14221 6253 14260 6287
rect 14294 6253 14333 6287
rect 14367 6253 14406 6287
rect 14440 6253 14479 6287
rect 14513 6253 14552 6287
rect 14586 6253 14625 6287
rect 14659 6253 14698 6287
rect 14732 6253 14771 6287
rect 14805 6253 14844 6287
rect 14878 6253 14917 6287
rect 14951 6253 14990 6287
rect 15024 6253 15063 6287
rect 15097 6253 15136 6287
rect 15170 6253 15209 6287
rect 15243 6253 15282 6287
rect 15316 6253 15355 6287
rect 15389 6253 15427 6287
rect 15461 6253 15499 6287
rect 15533 6253 15571 6287
rect 15605 6253 15643 6287
rect 15677 6253 15715 6287
rect 15749 6253 15787 6287
rect 15821 6253 15859 6287
rect 15893 6253 15931 6287
rect 15965 6253 16003 6287
rect 16037 6253 16075 6287
rect 16109 6253 16147 6287
rect 16181 6253 16219 6287
rect 16253 6253 16291 6287
rect 16649 6285 16650 6315
rect 16649 6279 16684 6285
rect 13450 6171 13484 6209
rect 13450 6095 13484 6135
rect 16683 6247 16684 6279
rect 16649 6213 16650 6245
rect 16649 6209 16684 6213
rect 16683 6175 16684 6209
rect 16649 6141 16650 6175
rect 16649 6139 16684 6141
rect 13804 6097 13844 6131
rect 13878 6097 13918 6131
rect 13952 6097 13992 6131
rect 14026 6097 14066 6131
rect 14100 6097 14140 6131
rect 14174 6097 14214 6131
rect 14248 6097 14288 6131
rect 14322 6097 14362 6131
rect 14396 6097 14436 6131
rect 14470 6097 14510 6131
rect 14544 6097 14584 6131
rect 14618 6097 14658 6131
rect 14692 6097 14732 6131
rect 14766 6097 14806 6131
rect 14840 6097 14880 6131
rect 14914 6097 14954 6131
rect 14988 6097 15028 6131
rect 15062 6097 15102 6131
rect 15136 6097 15176 6131
rect 15210 6097 15250 6131
rect 15284 6097 15323 6131
rect 15357 6097 15396 6131
rect 15430 6097 15469 6131
rect 15503 6097 15542 6131
rect 15576 6097 15615 6131
rect 15649 6097 15688 6131
rect 15722 6097 15761 6131
rect 15795 6097 15834 6131
rect 15868 6097 15907 6131
rect 15941 6097 15980 6131
rect 16014 6097 16053 6131
rect 16087 6097 16126 6131
rect 16160 6097 16199 6131
rect 16233 6097 16272 6131
rect 16306 6097 16345 6131
rect 16379 6097 16418 6131
rect 16683 6105 16684 6139
rect 16649 6103 16684 6105
rect 13450 6019 13484 6060
rect 13450 5969 13484 5984
rect 16649 6069 16650 6103
rect 16683 6035 16684 6069
rect 16649 6031 16684 6035
rect 16649 5999 16650 6031
rect 13332 5954 13366 5969
rect 13564 5941 13603 5975
rect 13637 5941 13676 5975
rect 13710 5941 13749 5975
rect 13783 5941 13822 5975
rect 13856 5941 13895 5975
rect 13929 5941 13968 5975
rect 14002 5941 14041 5975
rect 14075 5941 14114 5975
rect 14148 5941 14187 5975
rect 14221 5941 14260 5975
rect 14294 5941 14333 5975
rect 14367 5941 14406 5975
rect 14440 5941 14479 5975
rect 14513 5941 14552 5975
rect 14586 5941 14625 5975
rect 14659 5941 14698 5975
rect 14732 5941 14771 5975
rect 14805 5941 14844 5975
rect 14878 5941 14917 5975
rect 14951 5941 14990 5975
rect 15024 5941 15063 5975
rect 15097 5941 15136 5975
rect 15170 5941 15209 5975
rect 15243 5941 15282 5975
rect 15316 5941 15355 5975
rect 15389 5941 15427 5975
rect 15461 5941 15499 5975
rect 15533 5941 15571 5975
rect 15605 5941 15643 5975
rect 15677 5941 15715 5975
rect 15749 5941 15787 5975
rect 15821 5941 15859 5975
rect 15893 5941 15931 5975
rect 15965 5941 16003 5975
rect 16037 5941 16075 5975
rect 16109 5941 16147 5975
rect 16181 5941 16219 5975
rect 16253 5941 16291 5975
rect 16683 5965 16684 5997
rect 16649 5959 16684 5965
rect 13332 5881 13366 5900
rect 16649 5929 16650 5959
rect 16683 5895 16684 5925
rect 16649 5887 16684 5895
rect 16649 5879 16650 5887
rect 13366 5845 13407 5879
rect 13441 5845 13475 5879
rect 13509 5845 13543 5879
rect 13577 5845 13611 5879
rect 13645 5845 13679 5879
rect 13713 5845 13747 5879
rect 13781 5845 13815 5879
rect 13853 5845 13883 5879
rect 13926 5845 13951 5879
rect 13999 5845 14019 5879
rect 14072 5845 14087 5879
rect 14145 5845 14155 5879
rect 14218 5845 14223 5879
rect 14325 5845 14330 5879
rect 14393 5845 14403 5879
rect 14461 5845 14476 5879
rect 14529 5845 14549 5879
rect 14597 5845 14622 5879
rect 14665 5845 14695 5879
rect 14733 5845 14767 5879
rect 14802 5845 14835 5879
rect 14875 5845 14903 5879
rect 14948 5845 14971 5879
rect 15021 5845 15039 5879
rect 15094 5845 15107 5879
rect 15167 5845 15175 5879
rect 15240 5845 15243 5879
rect 15277 5845 15279 5879
rect 15345 5845 15352 5879
rect 15413 5845 15425 5879
rect 15481 5845 15498 5879
rect 15549 5845 15571 5879
rect 15617 5845 15644 5879
rect 15685 5845 15717 5879
rect 15753 5845 15787 5879
rect 15823 5845 15855 5879
rect 15895 5845 15923 5879
rect 15967 5845 15991 5879
rect 16039 5845 16059 5879
rect 16111 5845 16127 5879
rect 16183 5845 16195 5879
rect 16255 5845 16263 5879
rect 16327 5845 16332 5879
rect 16366 5845 16401 5879
rect 16435 5845 16470 5879
rect 16504 5845 16539 5879
rect 16573 5859 16650 5879
rect 16573 5845 16649 5859
rect 13332 5808 13366 5831
rect 16683 5825 16684 5853
rect 16649 5815 16684 5825
rect 16649 5789 16650 5815
rect 13332 5735 13366 5762
rect 13332 5662 13366 5693
rect 13332 5590 13366 5624
rect 13332 5520 13366 5555
rect 13332 5451 13366 5484
rect 13450 5743 13484 5755
rect 13564 5749 13603 5783
rect 13637 5749 13676 5783
rect 13710 5749 13749 5783
rect 13783 5749 13822 5783
rect 13856 5749 13895 5783
rect 13929 5749 13968 5783
rect 14002 5749 14041 5783
rect 14075 5749 14114 5783
rect 14148 5749 14187 5783
rect 14221 5749 14260 5783
rect 14294 5749 14333 5783
rect 14367 5749 14406 5783
rect 14440 5749 14479 5783
rect 14513 5749 14552 5783
rect 14586 5749 14625 5783
rect 14659 5749 14698 5783
rect 14732 5749 14771 5783
rect 14805 5749 14844 5783
rect 14878 5749 14917 5783
rect 14951 5749 14990 5783
rect 15024 5749 15063 5783
rect 15097 5749 15136 5783
rect 15170 5749 15209 5783
rect 15243 5749 15282 5783
rect 15316 5749 15355 5783
rect 15389 5749 15427 5783
rect 15461 5749 15499 5783
rect 15533 5749 15571 5783
rect 15605 5749 15643 5783
rect 15677 5749 15715 5783
rect 15749 5749 15787 5783
rect 15821 5749 15859 5783
rect 15893 5749 15931 5783
rect 15965 5749 16003 5783
rect 16037 5749 16075 5783
rect 16109 5749 16147 5783
rect 16181 5749 16219 5783
rect 16253 5749 16291 5783
rect 16683 5755 16684 5781
rect 13450 5667 13484 5705
rect 13450 5591 13484 5631
rect 16649 5743 16684 5755
rect 16649 5719 16650 5743
rect 16683 5685 16684 5709
rect 16649 5671 16684 5685
rect 16649 5649 16650 5671
rect 13804 5593 13844 5627
rect 13878 5593 13918 5627
rect 13952 5593 13992 5627
rect 14026 5593 14066 5627
rect 14100 5593 14140 5627
rect 14174 5593 14214 5627
rect 14248 5593 14288 5627
rect 14322 5593 14362 5627
rect 14396 5593 14436 5627
rect 14470 5593 14510 5627
rect 14544 5593 14584 5627
rect 14618 5593 14658 5627
rect 14692 5593 14732 5627
rect 14766 5593 14806 5627
rect 14840 5593 14880 5627
rect 14914 5593 14954 5627
rect 14988 5593 15028 5627
rect 15062 5593 15102 5627
rect 15136 5593 15176 5627
rect 15210 5593 15250 5627
rect 15284 5593 15323 5627
rect 15357 5593 15396 5627
rect 15430 5593 15469 5627
rect 15503 5593 15542 5627
rect 15576 5593 15615 5627
rect 15649 5593 15688 5627
rect 15722 5593 15761 5627
rect 15795 5593 15834 5627
rect 15868 5593 15907 5627
rect 15941 5593 15980 5627
rect 16014 5593 16053 5627
rect 16087 5593 16126 5627
rect 16160 5593 16199 5627
rect 16233 5593 16272 5627
rect 16306 5593 16345 5627
rect 16379 5593 16418 5627
rect 16683 5615 16684 5637
rect 16649 5599 16684 5615
rect 13450 5515 13484 5556
rect 13450 5465 13484 5480
rect 16649 5579 16650 5599
rect 16683 5545 16684 5565
rect 16649 5527 16684 5545
rect 16649 5509 16650 5527
rect 16683 5475 16684 5493
rect 13564 5437 13603 5471
rect 13637 5437 13676 5471
rect 13710 5437 13749 5471
rect 13783 5437 13822 5471
rect 13856 5437 13895 5471
rect 13929 5437 13968 5471
rect 14002 5437 14041 5471
rect 14075 5437 14114 5471
rect 14148 5437 14187 5471
rect 14221 5437 14260 5471
rect 14294 5437 14333 5471
rect 14367 5437 14406 5471
rect 14440 5437 14479 5471
rect 14513 5437 14552 5471
rect 14586 5437 14625 5471
rect 14659 5437 14698 5471
rect 14732 5437 14771 5471
rect 14805 5437 14844 5471
rect 14878 5437 14917 5471
rect 14951 5437 14990 5471
rect 15024 5437 15063 5471
rect 15097 5437 15136 5471
rect 15170 5437 15209 5471
rect 15243 5437 15282 5471
rect 15316 5437 15355 5471
rect 15389 5437 15427 5471
rect 15461 5437 15499 5471
rect 15533 5437 15571 5471
rect 15605 5437 15643 5471
rect 15677 5437 15715 5471
rect 15749 5437 15787 5471
rect 15821 5437 15859 5471
rect 15893 5437 15931 5471
rect 15965 5437 16003 5471
rect 16037 5437 16075 5471
rect 16109 5437 16147 5471
rect 16181 5437 16219 5471
rect 16253 5437 16291 5471
rect 16649 5455 16684 5475
rect 16649 5439 16650 5455
rect 13332 5381 13366 5412
rect 16683 5405 16684 5421
rect 16649 5383 16684 5405
rect 16649 5375 16650 5383
rect 13366 5341 13407 5375
rect 13441 5341 13475 5375
rect 13509 5341 13543 5375
rect 13577 5341 13611 5375
rect 13645 5341 13679 5375
rect 13713 5341 13747 5375
rect 13781 5341 13815 5375
rect 13853 5341 13883 5375
rect 13926 5341 13951 5375
rect 13999 5341 14019 5375
rect 14072 5341 14087 5375
rect 14145 5341 14155 5375
rect 14218 5341 14223 5375
rect 14325 5341 14330 5375
rect 14393 5341 14403 5375
rect 14461 5341 14476 5375
rect 14529 5341 14549 5375
rect 14597 5341 14622 5375
rect 14665 5341 14695 5375
rect 14733 5341 14767 5375
rect 14802 5341 14835 5375
rect 14875 5341 14903 5375
rect 14948 5341 14971 5375
rect 15021 5341 15039 5375
rect 15094 5341 15107 5375
rect 15167 5341 15175 5375
rect 15240 5341 15243 5375
rect 15277 5341 15279 5375
rect 15345 5341 15352 5375
rect 15413 5341 15425 5375
rect 15481 5341 15498 5375
rect 15549 5341 15571 5375
rect 15617 5341 15644 5375
rect 15685 5341 15717 5375
rect 15753 5341 15787 5375
rect 15823 5341 15855 5375
rect 15895 5341 15923 5375
rect 15967 5341 15991 5375
rect 16039 5341 16059 5375
rect 16111 5341 16127 5375
rect 16183 5341 16195 5375
rect 16255 5341 16263 5375
rect 16327 5341 16332 5375
rect 16366 5341 16401 5375
rect 16435 5341 16470 5375
rect 16504 5341 16539 5375
rect 16573 5369 16650 5375
rect 16573 5341 16649 5369
rect 13332 5311 13366 5340
rect 16683 5335 16684 5349
rect 16649 5311 16684 5335
rect 16649 5299 16650 5311
rect 13332 5241 13366 5268
rect 13332 5171 13366 5196
rect 13332 5101 13366 5124
rect 13332 5031 13366 5052
rect 13332 4961 13366 4980
rect 13450 5239 13484 5251
rect 13564 5245 13603 5279
rect 13637 5245 13676 5279
rect 13710 5245 13749 5279
rect 13783 5245 13822 5279
rect 13856 5245 13895 5279
rect 13929 5245 13968 5279
rect 14002 5245 14041 5279
rect 14075 5245 14114 5279
rect 14148 5245 14187 5279
rect 14221 5245 14260 5279
rect 14294 5245 14333 5279
rect 14367 5245 14406 5279
rect 14440 5245 14479 5279
rect 14513 5245 14552 5279
rect 14586 5245 14625 5279
rect 14659 5245 14698 5279
rect 14732 5245 14771 5279
rect 14805 5245 14844 5279
rect 14878 5245 14917 5279
rect 14951 5245 14990 5279
rect 15024 5245 15063 5279
rect 15097 5245 15136 5279
rect 15170 5245 15209 5279
rect 15243 5245 15282 5279
rect 15316 5245 15355 5279
rect 15389 5245 15428 5279
rect 15462 5245 15501 5279
rect 15535 5245 15573 5279
rect 15607 5245 15645 5279
rect 15679 5245 15717 5279
rect 15751 5245 15789 5279
rect 15823 5245 15861 5279
rect 15895 5245 15933 5279
rect 15967 5245 16005 5279
rect 16039 5245 16077 5279
rect 16111 5245 16149 5279
rect 16183 5245 16221 5279
rect 16255 5245 16293 5279
rect 16683 5265 16684 5277
rect 13450 5163 13484 5201
rect 13450 5087 13484 5127
rect 16649 5239 16684 5265
rect 16649 5230 16650 5239
rect 16683 5196 16684 5205
rect 16649 5167 16684 5196
rect 16649 5161 16650 5167
rect 16683 5127 16684 5133
rect 13804 5089 13844 5123
rect 13878 5089 13918 5123
rect 13952 5089 13992 5123
rect 14026 5089 14066 5123
rect 14100 5089 14140 5123
rect 14174 5089 14214 5123
rect 14248 5089 14288 5123
rect 14322 5089 14362 5123
rect 14396 5089 14436 5123
rect 14470 5089 14510 5123
rect 14544 5089 14583 5123
rect 14617 5089 14656 5123
rect 14690 5089 14729 5123
rect 14763 5089 14802 5123
rect 14836 5089 14875 5123
rect 14909 5089 14948 5123
rect 14982 5089 15021 5123
rect 15055 5089 15094 5123
rect 15128 5089 15167 5123
rect 15201 5089 15240 5123
rect 15274 5089 15313 5123
rect 15347 5089 15386 5123
rect 15420 5089 15459 5123
rect 15493 5089 15532 5123
rect 15566 5089 15605 5123
rect 15639 5089 15678 5123
rect 15712 5089 15751 5123
rect 15785 5089 15824 5123
rect 15858 5089 15897 5123
rect 15931 5089 15970 5123
rect 16004 5089 16043 5123
rect 16077 5089 16116 5123
rect 16150 5089 16189 5123
rect 16223 5089 16262 5123
rect 16296 5089 16335 5123
rect 16369 5089 16408 5123
rect 16649 5095 16684 5127
rect 16649 5092 16650 5095
rect 13450 5011 13484 5052
rect 13450 4961 13484 4976
rect 16683 5058 16684 5061
rect 16649 5023 16684 5058
rect 16683 5022 16684 5023
rect 16649 4988 16650 4989
rect 13564 4933 13603 4967
rect 13637 4933 13676 4967
rect 13710 4933 13749 4967
rect 13783 4933 13822 4967
rect 13856 4933 13895 4967
rect 13929 4933 13968 4967
rect 14002 4933 14041 4967
rect 14075 4933 14114 4967
rect 14148 4933 14187 4967
rect 14221 4933 14260 4967
rect 14294 4933 14333 4967
rect 14367 4933 14406 4967
rect 14440 4933 14479 4967
rect 14513 4933 14552 4967
rect 14586 4933 14625 4967
rect 14659 4933 14698 4967
rect 14732 4933 14771 4967
rect 14805 4933 14844 4967
rect 14878 4933 14917 4967
rect 14951 4933 14990 4967
rect 15024 4933 15063 4967
rect 15097 4933 15136 4967
rect 15170 4933 15209 4967
rect 15243 4933 15282 4967
rect 15316 4933 15355 4967
rect 15389 4933 15428 4967
rect 15462 4933 15501 4967
rect 15535 4933 15573 4967
rect 15607 4933 15645 4967
rect 15679 4933 15717 4967
rect 15751 4933 15789 4967
rect 15823 4933 15861 4967
rect 15895 4933 15933 4967
rect 15967 4933 16005 4967
rect 16039 4933 16077 4967
rect 16111 4933 16149 4967
rect 16183 4933 16221 4967
rect 16255 4933 16293 4967
rect 16649 4954 16684 4988
rect 16683 4949 16684 4954
rect 13332 4891 13366 4908
rect 16649 4915 16650 4920
rect 16649 4885 16684 4915
rect 16683 4876 16684 4885
rect 13366 4837 13407 4871
rect 13441 4837 13475 4871
rect 13509 4837 13543 4871
rect 13577 4837 13611 4871
rect 13645 4837 13679 4871
rect 13713 4837 13747 4871
rect 13781 4837 13815 4871
rect 13853 4837 13883 4871
rect 13926 4837 13951 4871
rect 13999 4837 14019 4871
rect 14072 4837 14087 4871
rect 14145 4837 14155 4871
rect 14218 4837 14223 4871
rect 14325 4837 14330 4871
rect 14393 4837 14403 4871
rect 14461 4837 14476 4871
rect 14529 4837 14549 4871
rect 14597 4837 14622 4871
rect 14665 4837 14695 4871
rect 14733 4837 14767 4871
rect 14802 4837 14835 4871
rect 14875 4837 14903 4871
rect 14948 4837 14971 4871
rect 15021 4837 15039 4871
rect 15094 4837 15107 4871
rect 15167 4837 15175 4871
rect 15240 4837 15243 4871
rect 15277 4837 15279 4871
rect 15345 4837 15352 4871
rect 15413 4837 15425 4871
rect 15481 4837 15498 4871
rect 15549 4837 15571 4871
rect 15617 4837 15644 4871
rect 15685 4837 15717 4871
rect 15753 4837 15787 4871
rect 15823 4837 15855 4871
rect 15895 4837 15923 4871
rect 15967 4837 15991 4871
rect 16039 4837 16059 4871
rect 16111 4837 16127 4871
rect 16183 4837 16195 4871
rect 16255 4837 16263 4871
rect 16327 4837 16332 4871
rect 16366 4837 16401 4871
rect 16435 4837 16470 4871
rect 16504 4837 16539 4871
rect 16573 4851 16649 4871
rect 16573 4842 16650 4851
rect 16573 4837 16684 4842
rect 13332 4821 13366 4836
rect 16649 4816 16684 4837
rect 16683 4803 16684 4816
rect 13332 4751 13366 4764
rect 13332 4681 13366 4692
rect 13332 4611 13366 4620
rect 13332 4541 13366 4548
rect 13332 4471 13366 4476
rect 13450 4735 13484 4747
rect 13564 4741 13603 4775
rect 13637 4741 13676 4775
rect 13710 4741 13749 4775
rect 13783 4741 13822 4775
rect 13856 4741 13895 4775
rect 13929 4741 13968 4775
rect 14002 4741 14041 4775
rect 14075 4741 14114 4775
rect 14148 4741 14187 4775
rect 14221 4741 14260 4775
rect 14294 4741 14333 4775
rect 14367 4741 14406 4775
rect 14440 4741 14479 4775
rect 14513 4741 14552 4775
rect 14586 4741 14625 4775
rect 14659 4741 14698 4775
rect 14732 4741 14771 4775
rect 14805 4741 14844 4775
rect 14878 4741 14917 4775
rect 14951 4741 14990 4775
rect 15024 4741 15063 4775
rect 15097 4741 15136 4775
rect 15170 4741 15209 4775
rect 15243 4741 15282 4775
rect 15316 4741 15355 4775
rect 15389 4741 15428 4775
rect 15462 4741 15501 4775
rect 15535 4741 15573 4775
rect 15607 4741 15645 4775
rect 15679 4741 15717 4775
rect 15751 4741 15789 4775
rect 15823 4741 15861 4775
rect 15895 4741 15933 4775
rect 15967 4741 16005 4775
rect 16039 4741 16077 4775
rect 16111 4741 16149 4775
rect 16183 4741 16221 4775
rect 16255 4741 16293 4775
rect 16649 4769 16650 4782
rect 16649 4747 16684 4769
rect 13450 4659 13484 4697
rect 13450 4582 13484 4623
rect 16683 4730 16684 4747
rect 16649 4696 16650 4713
rect 16649 4678 16684 4696
rect 16683 4657 16684 4678
rect 16649 4623 16650 4644
rect 13804 4585 13844 4619
rect 13878 4585 13918 4619
rect 13952 4585 13992 4619
rect 14026 4585 14066 4619
rect 14100 4585 14140 4619
rect 14174 4585 14214 4619
rect 14248 4585 14288 4619
rect 14322 4585 14362 4619
rect 14396 4585 14435 4619
rect 14469 4585 14508 4619
rect 14542 4585 14581 4619
rect 14615 4585 14654 4619
rect 14688 4585 14727 4619
rect 14761 4585 14800 4619
rect 14834 4585 14873 4619
rect 14907 4585 14946 4619
rect 14980 4585 15019 4619
rect 15053 4585 15092 4619
rect 15126 4585 15165 4619
rect 15199 4585 15238 4619
rect 15272 4585 15311 4619
rect 15345 4585 15384 4619
rect 15418 4585 15457 4619
rect 15491 4585 15530 4619
rect 15564 4585 15603 4619
rect 15637 4585 15676 4619
rect 15710 4585 15749 4619
rect 15783 4585 15822 4619
rect 15856 4585 15895 4619
rect 15929 4585 15968 4619
rect 16002 4585 16041 4619
rect 16075 4585 16114 4619
rect 16148 4585 16187 4619
rect 16221 4585 16260 4619
rect 16294 4585 16333 4619
rect 16367 4585 16406 4619
rect 16649 4609 16684 4623
rect 13450 4507 13484 4548
rect 13450 4457 13484 4471
rect 16683 4584 16684 4609
rect 16649 4550 16650 4575
rect 16649 4540 16684 4550
rect 16683 4511 16684 4540
rect 16649 4477 16650 4506
rect 16649 4471 16684 4477
rect 13564 4429 13603 4463
rect 13637 4429 13676 4463
rect 13710 4429 13749 4463
rect 13783 4429 13822 4463
rect 13856 4429 13895 4463
rect 13929 4429 13968 4463
rect 14002 4429 14041 4463
rect 14075 4429 14114 4463
rect 14148 4429 14187 4463
rect 14221 4429 14260 4463
rect 14294 4429 14333 4463
rect 14367 4429 14406 4463
rect 14440 4429 14479 4463
rect 14513 4429 14552 4463
rect 14586 4429 14625 4463
rect 14659 4429 14698 4463
rect 14732 4429 14771 4463
rect 14805 4429 14844 4463
rect 14878 4429 14917 4463
rect 14951 4429 14990 4463
rect 15024 4429 15063 4463
rect 15097 4429 15136 4463
rect 15170 4429 15209 4463
rect 15243 4429 15282 4463
rect 15316 4429 15355 4463
rect 15389 4429 15428 4463
rect 15462 4429 15501 4463
rect 15535 4429 15574 4463
rect 15608 4429 15646 4463
rect 15680 4429 15718 4463
rect 15752 4429 15790 4463
rect 15824 4429 15862 4463
rect 15896 4429 15934 4463
rect 15968 4429 16006 4463
rect 16040 4429 16078 4463
rect 16112 4429 16150 4463
rect 16184 4429 16222 4463
rect 16256 4429 16294 4463
rect 16683 4438 16684 4471
rect 13332 4401 13366 4404
rect 16649 4404 16650 4437
rect 13332 4366 13436 4367
rect 13470 4366 13505 4367
rect 13539 4366 13574 4367
rect 13608 4366 13643 4367
rect 13677 4366 13712 4367
rect 13746 4366 13781 4367
rect 13815 4366 13850 4367
rect 13884 4366 13919 4367
rect 13953 4366 13988 4367
rect 13332 4332 13356 4366
rect 13390 4333 13436 4366
rect 13473 4333 13505 4366
rect 13546 4333 13574 4366
rect 13619 4333 13643 4366
rect 13692 4333 13712 4366
rect 13765 4333 13781 4366
rect 13838 4333 13850 4366
rect 13911 4333 13919 4366
rect 13984 4333 13988 4366
rect 14022 4366 14057 4367
rect 14022 4333 14023 4366
rect 13390 4332 13439 4333
rect 13473 4332 13512 4333
rect 13546 4332 13585 4333
rect 13619 4332 13658 4333
rect 13692 4332 13731 4333
rect 13765 4332 13804 4333
rect 13838 4332 13877 4333
rect 13911 4332 13950 4333
rect 13984 4332 14023 4333
rect 14091 4366 14126 4367
rect 14160 4366 14195 4367
rect 14229 4366 14264 4367
rect 14298 4366 14333 4367
rect 14367 4366 14402 4367
rect 14436 4366 14471 4367
rect 14505 4366 14540 4367
rect 14574 4366 14609 4367
rect 14091 4333 14096 4366
rect 14160 4333 14169 4366
rect 14229 4333 14242 4366
rect 14298 4333 14315 4366
rect 14367 4333 14388 4366
rect 14436 4333 14461 4366
rect 14505 4333 14534 4366
rect 14574 4333 14607 4366
rect 14643 4333 14678 4367
rect 14712 4366 14747 4367
rect 14781 4366 14816 4367
rect 14850 4366 14885 4367
rect 14919 4366 14954 4367
rect 14988 4366 15023 4367
rect 15057 4366 15092 4367
rect 15126 4366 15161 4367
rect 15195 4366 15230 4367
rect 14714 4333 14747 4366
rect 14787 4333 14816 4366
rect 14860 4333 14885 4366
rect 14933 4333 14954 4366
rect 15006 4333 15023 4366
rect 15079 4333 15092 4366
rect 15152 4333 15161 4366
rect 15225 4333 15230 4366
rect 15264 4366 15299 4367
rect 14057 4332 14096 4333
rect 14130 4332 14169 4333
rect 14203 4332 14242 4333
rect 14276 4332 14315 4333
rect 14349 4332 14388 4333
rect 14422 4332 14461 4333
rect 14495 4332 14534 4333
rect 14568 4332 14607 4333
rect 14641 4332 14680 4333
rect 14714 4332 14753 4333
rect 14787 4332 14826 4333
rect 14860 4332 14899 4333
rect 14933 4332 14972 4333
rect 15006 4332 15045 4333
rect 15079 4332 15118 4333
rect 15152 4332 15191 4333
rect 15225 4332 15264 4333
rect 15298 4333 15299 4366
rect 15333 4366 15368 4367
rect 15402 4366 15437 4367
rect 15471 4366 15506 4367
rect 15540 4366 15575 4367
rect 15609 4366 15644 4367
rect 15678 4366 15713 4367
rect 15747 4366 15782 4367
rect 15816 4366 15851 4367
rect 15333 4333 15337 4366
rect 15402 4333 15410 4366
rect 15471 4333 15483 4366
rect 15540 4333 15556 4366
rect 15609 4333 15629 4366
rect 15678 4333 15702 4366
rect 15747 4333 15775 4366
rect 15816 4333 15848 4366
rect 15885 4333 15920 4367
rect 15954 4366 15989 4367
rect 16023 4366 16058 4367
rect 16092 4366 16127 4367
rect 16161 4366 16196 4367
rect 16230 4366 16265 4367
rect 16299 4366 16335 4367
rect 16369 4366 16405 4367
rect 16439 4366 16475 4367
rect 16509 4366 16545 4367
rect 16579 4366 16615 4367
rect 15955 4333 15989 4366
rect 16028 4333 16058 4366
rect 16101 4333 16127 4366
rect 16174 4333 16196 4366
rect 16247 4333 16265 4366
rect 16320 4333 16335 4366
rect 16393 4333 16405 4366
rect 16466 4333 16475 4366
rect 16539 4333 16545 4366
rect 16612 4333 16615 4366
rect 16649 4333 16684 4404
rect 15298 4332 15337 4333
rect 15371 4332 15410 4333
rect 15444 4332 15483 4333
rect 15517 4332 15556 4333
rect 15590 4332 15629 4333
rect 15663 4332 15702 4333
rect 15736 4332 15775 4333
rect 15809 4332 15848 4333
rect 15882 4332 15921 4333
rect 15955 4332 15994 4333
rect 16028 4332 16067 4333
rect 16101 4332 16140 4333
rect 16174 4332 16213 4333
rect 16247 4332 16286 4333
rect 16320 4332 16359 4333
rect 16393 4332 16432 4333
rect 16466 4332 16505 4333
rect 16539 4332 16578 4333
rect 16612 4332 16684 4333
rect 16835 6384 16837 6418
rect 16871 6384 16951 6418
rect 16985 6384 16986 6418
rect 16835 6346 16986 6384
rect 16835 6312 16837 6346
rect 16871 6312 16951 6346
rect 16985 6312 16986 6346
rect 16835 6274 16986 6312
rect 16835 6240 16837 6274
rect 16871 6240 16951 6274
rect 16985 6240 16986 6274
rect 16835 6202 16986 6240
rect 16835 6168 16837 6202
rect 16871 6168 16951 6202
rect 16985 6168 16986 6202
rect 16835 6130 16986 6168
rect 16835 6096 16837 6130
rect 16871 6096 16951 6130
rect 16985 6096 16986 6130
rect 16835 6058 16986 6096
rect 16835 6024 16837 6058
rect 16871 6024 16951 6058
rect 16985 6024 16986 6058
rect 16835 5986 16986 6024
rect 16835 5952 16837 5986
rect 16871 5952 16951 5986
rect 16985 5952 16986 5986
rect 16835 5914 16986 5952
rect 16835 5880 16837 5914
rect 16871 5880 16951 5914
rect 16985 5880 16986 5914
rect 16835 5842 16986 5880
rect 16835 5808 16837 5842
rect 16871 5808 16951 5842
rect 16985 5808 16986 5842
rect 16835 5770 16986 5808
rect 16835 5736 16837 5770
rect 16871 5736 16951 5770
rect 16985 5736 16986 5770
rect 16835 5698 16986 5736
rect 16835 5664 16837 5698
rect 16871 5664 16951 5698
rect 16985 5664 16986 5698
rect 16835 5626 16986 5664
rect 16835 5592 16837 5626
rect 16871 5592 16951 5626
rect 16985 5592 16986 5626
rect 16835 5554 16986 5592
rect 16835 5520 16837 5554
rect 16871 5520 16951 5554
rect 16985 5520 16986 5554
rect 16835 5482 16986 5520
rect 16835 5448 16837 5482
rect 16871 5448 16951 5482
rect 16985 5448 16986 5482
rect 16835 5410 16986 5448
rect 16835 5376 16837 5410
rect 16871 5376 16951 5410
rect 16985 5376 16986 5410
rect 16835 5338 16986 5376
rect 16835 5304 16837 5338
rect 16871 5304 16951 5338
rect 16985 5304 16986 5338
rect 16835 5266 16986 5304
rect 16835 5232 16837 5266
rect 16871 5232 16951 5266
rect 16985 5232 16986 5266
rect 16835 5194 16986 5232
rect 16835 5160 16837 5194
rect 16871 5160 16951 5194
rect 16985 5160 16986 5194
rect 16835 5122 16986 5160
rect 16835 5088 16837 5122
rect 16871 5088 16951 5122
rect 16985 5088 16986 5122
rect 16835 5050 16986 5088
rect 16835 5016 16837 5050
rect 16871 5016 16951 5050
rect 16985 5016 16986 5050
rect 16835 4978 16986 5016
rect 16835 4944 16837 4978
rect 16871 4944 16951 4978
rect 16985 4944 16986 4978
rect 16835 4906 16986 4944
rect 16835 4872 16837 4906
rect 16871 4872 16951 4906
rect 16985 4872 16986 4906
rect 16835 4834 16986 4872
rect 16835 4800 16837 4834
rect 16871 4800 16951 4834
rect 16985 4800 16986 4834
rect 16835 4762 16986 4800
rect 16835 4728 16837 4762
rect 16871 4728 16951 4762
rect 16985 4728 16986 4762
rect 16835 4690 16986 4728
rect 16835 4656 16837 4690
rect 16871 4656 16951 4690
rect 16985 4656 16986 4690
rect 16835 4618 16986 4656
rect 16835 4584 16837 4618
rect 16871 4584 16951 4618
rect 16985 4584 16986 4618
rect 16835 4546 16986 4584
rect 16835 4512 16837 4546
rect 16871 4512 16951 4546
rect 16985 4512 16986 4546
rect 16835 4474 16986 4512
rect 16835 4440 16837 4474
rect 16871 4440 16951 4474
rect 16985 4440 16986 4474
rect 16835 4402 16986 4440
rect 16835 4368 16837 4402
rect 16871 4368 16951 4402
rect 16985 4368 16986 4402
rect 13030 4296 13032 4330
rect 13066 4296 13146 4330
rect 13030 4257 13180 4296
rect 13030 4223 13032 4257
rect 13066 4223 13146 4257
rect 13030 4169 13180 4223
rect 16835 4330 16986 4368
rect 16835 4296 16837 4330
rect 16871 4296 16951 4330
rect 16985 4296 16986 4330
rect 16835 4257 16986 4296
rect 16835 4223 16837 4257
rect 16871 4223 16951 4257
rect 16985 4223 16986 4257
rect 16835 4169 16986 4223
rect 13030 4168 16986 4169
rect 13030 4134 13038 4168
rect 13072 4145 13111 4168
rect 13099 4134 13111 4145
rect 13145 4134 13184 4168
rect 13218 4134 13257 4168
rect 13291 4134 13330 4168
rect 13364 4134 13403 4168
rect 13437 4134 13476 4168
rect 13510 4134 13549 4168
rect 13583 4134 13622 4168
rect 13656 4134 13695 4168
rect 13729 4134 13768 4168
rect 13802 4134 13841 4168
rect 13875 4134 13914 4168
rect 13948 4134 13987 4168
rect 14021 4134 14060 4168
rect 14094 4134 14133 4168
rect 14167 4134 14206 4168
rect 14240 4134 14279 4168
rect 14313 4134 14352 4168
rect 14386 4134 14425 4168
rect 14459 4134 14497 4168
rect 14531 4134 14569 4168
rect 14603 4134 14641 4168
rect 14675 4134 14713 4168
rect 14747 4134 14785 4168
rect 14819 4134 14857 4168
rect 14891 4134 14929 4168
rect 14963 4134 15001 4168
rect 15035 4134 15073 4168
rect 15107 4134 15145 4168
rect 15179 4134 15217 4168
rect 15251 4134 15289 4168
rect 15323 4134 15361 4168
rect 15395 4134 15433 4168
rect 15467 4134 15505 4168
rect 15539 4134 15577 4168
rect 15611 4134 15649 4168
rect 15683 4134 15721 4168
rect 15755 4134 15793 4168
rect 15827 4134 15865 4168
rect 15899 4134 15937 4168
rect 15971 4134 16009 4168
rect 16043 4134 16081 4168
rect 16115 4134 16153 4168
rect 16187 4134 16225 4168
rect 16259 4134 16297 4168
rect 16331 4134 16369 4168
rect 16403 4134 16441 4168
rect 16475 4134 16513 4168
rect 16547 4134 16585 4168
rect 16619 4134 16657 4168
rect 16691 4134 16729 4168
rect 16763 4134 16801 4168
rect 16835 4134 16873 4168
rect 16907 4145 16945 4168
rect 16907 4134 16927 4145
rect 16979 4134 16986 4168
rect 13030 4111 13065 4134
rect 13099 4111 16927 4134
rect 16961 4111 16986 4134
rect 13030 4077 16986 4111
rect 13030 4054 13092 4077
rect 13126 4054 16900 4077
rect 16934 4054 16986 4077
rect 13030 4020 13038 4054
rect 13072 4043 13092 4054
rect 13072 4020 13111 4043
rect 13145 4020 13184 4054
rect 13218 4020 13257 4054
rect 13291 4020 13330 4054
rect 13364 4020 13403 4054
rect 13437 4020 13476 4054
rect 13510 4020 13549 4054
rect 13583 4020 13622 4054
rect 13656 4020 13695 4054
rect 13729 4020 13768 4054
rect 13802 4020 13841 4054
rect 13875 4020 13914 4054
rect 13948 4020 13987 4054
rect 14021 4020 14060 4054
rect 14094 4020 14133 4054
rect 14167 4020 14206 4054
rect 14240 4020 14279 4054
rect 14313 4020 14352 4054
rect 14386 4020 14425 4054
rect 14459 4020 14497 4054
rect 14531 4020 14569 4054
rect 14603 4020 14641 4054
rect 14675 4020 14713 4054
rect 14747 4020 14785 4054
rect 14819 4020 14857 4054
rect 14891 4020 14929 4054
rect 14963 4020 15001 4054
rect 15035 4020 15073 4054
rect 15107 4020 15145 4054
rect 15179 4020 15217 4054
rect 15251 4020 15289 4054
rect 15323 4020 15361 4054
rect 15395 4020 15433 4054
rect 15467 4020 15505 4054
rect 15539 4020 15577 4054
rect 15611 4020 15649 4054
rect 15683 4020 15721 4054
rect 15755 4020 15793 4054
rect 15827 4020 15865 4054
rect 15899 4020 15937 4054
rect 15971 4020 16009 4054
rect 16043 4020 16081 4054
rect 16115 4020 16153 4054
rect 16187 4020 16225 4054
rect 16259 4020 16297 4054
rect 16331 4020 16369 4054
rect 16403 4020 16441 4054
rect 16475 4020 16513 4054
rect 16547 4020 16585 4054
rect 16619 4020 16657 4054
rect 16691 4020 16729 4054
rect 16763 4020 16801 4054
rect 16835 4020 16873 4054
rect 16934 4043 16945 4054
rect 16907 4020 16945 4043
rect 16979 4020 16986 4054
rect 13030 4019 16986 4020
rect 12629 3836 12634 3860
rect 12668 3836 12760 3860
rect 12794 3836 12799 3860
rect 12629 3800 12799 3836
rect 17216 3898 17386 3924
rect 17216 3864 17218 3898
rect 17252 3864 17344 3898
rect 17378 3864 17386 3898
rect 17216 3800 17386 3864
rect 4235 3743 4269 3770
rect 3008 3648 3046 3682
rect 3080 3648 3118 3682
rect 3944 3648 3983 3682
rect 4017 3648 4055 3682
rect 4089 3648 4127 3682
rect 1310 3594 1348 3628
rect 1622 3594 1660 3628
rect 1934 3594 1972 3628
rect 2246 3594 2284 3628
rect 2318 3594 2438 3628
rect 1312 3552 1346 3594
rect 1624 3552 1658 3594
rect 1936 3552 1970 3594
rect 2248 3552 2282 3594
rect 3198 3566 3232 3580
rect 2092 3540 2208 3552
rect 62 217 126 3479
rect 1156 3468 1190 3506
rect 1156 3396 1190 3434
rect 1468 3468 1502 3506
rect 1468 3396 1502 3434
rect 1780 3468 1814 3506
rect 1780 3396 1814 3434
rect 2126 3506 2208 3540
rect 2092 3468 2208 3506
rect 2126 3434 2208 3468
rect 2092 3396 2208 3434
rect 2126 3362 2208 3396
rect 2092 3087 2208 3362
rect 1156 3015 1190 3053
rect 1156 2943 1190 2981
rect 1156 2871 1190 2909
rect 1156 2799 1190 2837
rect 1156 2727 1190 2765
rect 1468 3015 1502 3053
rect 1468 2943 1502 2981
rect 1468 2871 1502 2909
rect 1468 2799 1502 2837
rect 1468 2727 1502 2765
rect 1780 3015 1814 3053
rect 1780 2943 1814 2981
rect 1780 2871 1814 2909
rect 1780 2799 1814 2837
rect 1780 2727 1814 2765
rect 2126 3053 2208 3087
rect 2092 3015 2208 3053
rect 2126 2981 2208 3015
rect 2092 2970 2208 2981
rect 2322 2970 2478 3552
rect 2879 3532 2895 3566
rect 2929 3532 2964 3566
rect 2998 3532 3033 3566
rect 3067 3532 3102 3566
rect 3136 3532 3171 3566
rect 3205 3542 3240 3566
rect 3232 3532 3240 3542
rect 3274 3532 3309 3566
rect 3343 3532 3378 3566
rect 3412 3532 3447 3566
rect 3481 3532 3516 3566
rect 3550 3532 3585 3566
rect 3619 3532 3654 3566
rect 3688 3532 3723 3566
rect 3757 3532 3792 3566
rect 3826 3532 3861 3566
rect 3895 3532 3930 3566
rect 3964 3532 3999 3566
rect 4033 3532 4069 3566
rect 4103 3532 4139 3566
rect 4173 3532 4189 3566
rect 2092 2943 2478 2970
rect 2126 2909 2478 2943
rect 2092 2871 2478 2909
rect 2126 2837 2478 2871
rect 2092 2809 2478 2837
rect 2092 2799 2126 2809
rect 2092 2727 2126 2765
rect 186 178 220 216
rect 186 106 220 144
rect 618 178 652 216
rect 618 106 652 144
rect 170 -38 236 68
rect 602 -38 668 68
rect 164 -72 180 -38
rect 502 -72 596 -38
<< viali >>
rect 2318 8119 2352 8153
rect 2318 8047 2352 8081
rect 49 7961 83 7995
rect 49 7889 83 7923
rect 2241 7499 2275 7533
rect 2241 7427 2275 7461
rect 349 6953 383 6987
rect 421 6953 455 6987
rect 325 5709 330 5743
rect 330 5709 359 5743
rect 397 5709 398 5743
rect 398 5709 431 5743
rect 469 5709 500 5743
rect 500 5709 503 5743
rect 135 5286 169 5320
rect 135 5214 169 5248
rect 135 5142 169 5176
rect 447 5286 481 5320
rect 447 5214 481 5248
rect 447 5142 481 5176
rect 213 5055 247 5089
rect 213 4983 247 5017
rect 288 4840 322 4874
rect 288 4768 322 4802
rect 603 5055 637 5089
rect 603 4983 637 5017
rect 146 4644 155 4678
rect 155 4644 180 4678
rect 218 4644 223 4678
rect 223 4644 252 4678
rect 381 4574 415 4608
rect 381 4502 415 4536
rect 80 3936 114 3970
rect 80 3864 114 3898
rect 80 3792 114 3826
rect 474 4275 508 4309
rect 474 4203 508 4237
rect 474 4094 508 4128
rect 474 4022 508 4056
rect 225 3678 259 3712
rect 297 3678 331 3712
rect 759 5286 793 5320
rect 759 5214 793 5248
rect 759 5142 793 5176
rect 915 5055 949 5089
rect 915 4983 949 5017
rect 1071 5286 1105 5320
rect 1071 5214 1105 5248
rect 1071 5142 1105 5176
rect 1383 5286 1417 5320
rect 1383 5214 1417 5248
rect 1383 5142 1417 5176
rect 1695 5286 1729 5320
rect 1695 5214 1729 5248
rect 1695 5142 1729 5176
rect 2007 5286 2041 5320
rect 2007 5214 2041 5248
rect 2007 5142 2041 5176
rect 1305 5055 1339 5089
rect 2089 5055 2123 5089
rect 1305 4983 1339 5017
rect 1768 4999 1802 5033
rect 1768 4927 1802 4961
rect 1227 4841 1261 4875
rect 1227 4769 1261 4803
rect 1539 4841 1573 4875
rect 1539 4769 1573 4803
rect 904 4564 938 4598
rect 976 4564 1010 4598
rect 1115 4672 1149 4678
rect 1187 4672 1221 4678
rect 1115 4644 1149 4672
rect 1187 4644 1217 4672
rect 1217 4644 1221 4672
rect 1324 4564 1358 4598
rect 1396 4564 1430 4598
rect 1142 4508 1176 4542
rect 1214 4530 1248 4542
rect 1214 4508 1248 4530
rect 1471 4454 1505 4462
rect 1471 4428 1505 4454
rect 1044 4335 1078 4369
rect 1044 4263 1078 4297
rect 902 4150 936 4184
rect 902 4078 936 4112
rect 605 3698 609 3712
rect 609 3698 639 3712
rect 677 3698 711 3712
rect 605 3678 639 3698
rect 677 3678 711 3698
rect 1438 3936 1472 3970
rect 1438 3864 1472 3898
rect 1438 3792 1472 3826
rect 1628 4564 1662 4598
rect 1700 4564 1734 4598
rect 1126 3672 1160 3706
rect 2089 4983 2123 5017
rect 1851 4841 1885 4875
rect 1851 4769 1885 4803
rect 2237 5286 2271 5320
rect 2237 5214 2271 5248
rect 2237 5142 2271 5176
rect 2163 4564 2197 4598
rect 2235 4564 2269 4598
rect 2315 4558 2349 4592
rect 2315 4486 2349 4520
rect 2395 7861 2429 7895
rect 2395 7789 2429 7823
rect 3198 7732 3232 7766
rect 3198 7660 3232 7694
rect 3046 7573 3080 7607
rect 3118 7573 3152 7607
rect 3500 7606 3534 7640
rect 3572 7606 3606 7640
rect 3644 7606 3678 7640
rect 3368 7073 3402 7107
rect 3368 7001 3402 7035
rect 3368 6929 3402 6963
rect 12643 7047 12677 7081
rect 12716 7047 12750 7081
rect 12789 7047 12823 7081
rect 12862 7047 12896 7081
rect 12935 7047 12969 7081
rect 13008 7047 13042 7081
rect 13081 7047 13115 7081
rect 13154 7047 13188 7081
rect 13227 7047 13261 7081
rect 13300 7047 13334 7081
rect 13373 7047 13407 7081
rect 13446 7047 13480 7081
rect 13519 7047 13553 7081
rect 13592 7047 13626 7081
rect 13665 7047 13699 7081
rect 13738 7047 13772 7081
rect 13811 7047 13845 7081
rect 13884 7047 13918 7081
rect 13957 7047 13991 7081
rect 14029 7047 14063 7081
rect 14101 7047 14135 7081
rect 14173 7047 14207 7081
rect 14245 7047 14279 7081
rect 14317 7047 14351 7081
rect 14389 7047 14423 7081
rect 14461 7047 14495 7081
rect 14533 7047 14567 7081
rect 14605 7047 14639 7081
rect 14677 7047 14711 7081
rect 14749 7047 14783 7081
rect 14821 7047 14855 7081
rect 14893 7047 14927 7081
rect 14965 7047 14999 7081
rect 15037 7047 15071 7081
rect 15109 7047 15143 7081
rect 15181 7047 15215 7081
rect 15253 7047 15287 7081
rect 15325 7047 15359 7081
rect 15397 7047 15431 7081
rect 15469 7047 15503 7081
rect 15541 7047 15575 7081
rect 15613 7047 15647 7081
rect 15685 7047 15719 7081
rect 15757 7047 15791 7081
rect 15829 7047 15863 7081
rect 15901 7047 15935 7081
rect 15973 7047 16007 7081
rect 16045 7047 16079 7081
rect 16117 7047 16151 7081
rect 16189 7047 16223 7081
rect 16261 7047 16295 7081
rect 16333 7047 16367 7081
rect 16405 7047 16439 7081
rect 16477 7047 16511 7081
rect 16549 7047 16583 7081
rect 16621 7047 16655 7081
rect 16693 7047 16727 7081
rect 16765 7047 16799 7081
rect 16837 7047 16871 7081
rect 16909 7047 16943 7081
rect 16981 7047 17015 7081
rect 17053 7047 17087 7081
rect 17125 7047 17159 7081
rect 12643 6954 12677 6955
rect 12643 6921 12663 6954
rect 12663 6921 12677 6954
rect 12716 6921 12750 6955
rect 12789 6921 12823 6955
rect 12862 6921 12896 6955
rect 12935 6921 12969 6955
rect 13008 6921 13042 6955
rect 13081 6921 13115 6955
rect 13154 6921 13188 6955
rect 13227 6921 13261 6955
rect 13300 6921 13334 6955
rect 13373 6921 13407 6955
rect 13446 6921 13480 6955
rect 13519 6921 13553 6955
rect 13592 6921 13626 6955
rect 13665 6921 13699 6955
rect 13738 6921 13772 6955
rect 13811 6921 13845 6955
rect 13884 6921 13918 6955
rect 13957 6921 13991 6955
rect 14029 6921 14063 6955
rect 14101 6921 14135 6955
rect 14173 6921 14207 6955
rect 14245 6921 14279 6955
rect 14317 6921 14351 6955
rect 14389 6921 14423 6955
rect 14461 6921 14495 6955
rect 14533 6921 14567 6955
rect 14605 6921 14639 6955
rect 14677 6921 14711 6955
rect 14749 6921 14783 6955
rect 14821 6921 14855 6955
rect 14893 6921 14927 6955
rect 14965 6921 14999 6955
rect 15037 6921 15071 6955
rect 15109 6921 15143 6955
rect 15181 6921 15215 6955
rect 15253 6921 15287 6955
rect 15325 6921 15359 6955
rect 15397 6921 15431 6955
rect 15469 6921 15503 6955
rect 15541 6921 15575 6955
rect 15613 6921 15647 6955
rect 15685 6921 15719 6955
rect 15757 6921 15791 6955
rect 15829 6921 15863 6955
rect 15901 6921 15935 6955
rect 15973 6921 16007 6955
rect 16045 6921 16079 6955
rect 16117 6921 16151 6955
rect 16189 6921 16223 6955
rect 16261 6921 16295 6955
rect 16333 6921 16367 6955
rect 16405 6921 16439 6955
rect 16477 6921 16511 6955
rect 16549 6921 16583 6955
rect 16621 6921 16655 6955
rect 16693 6921 16727 6955
rect 16765 6921 16799 6955
rect 16837 6921 16871 6955
rect 16909 6921 16943 6955
rect 16981 6921 17015 6955
rect 17053 6921 17087 6955
rect 17125 6921 17151 6955
rect 17151 6921 17159 6955
rect 17218 6950 17252 6969
rect 17218 6935 17252 6950
rect 17344 6935 17378 6969
rect 12634 6836 12668 6870
rect 12760 6836 12794 6870
rect 12634 6763 12668 6797
rect 12760 6763 12794 6797
rect 2849 6699 2883 6733
rect 12634 6690 12668 6724
rect 12760 6690 12794 6724
rect 2849 6627 2883 6661
rect 2942 6617 2958 6651
rect 2958 6617 2976 6651
rect 3014 6617 3026 6651
rect 3026 6617 3048 6651
rect 3086 6617 3120 6651
rect 3426 6623 3460 6657
rect 3498 6623 3532 6657
rect 3570 6623 3604 6657
rect 3642 6623 3676 6657
rect 17218 6862 17252 6896
rect 17344 6862 17378 6896
rect 17218 6789 17252 6823
rect 17344 6789 17378 6823
rect 17218 6716 17252 6750
rect 17344 6716 17378 6750
rect 12634 6617 12668 6651
rect 12760 6617 12794 6651
rect 2849 6555 2883 6589
rect 3375 6549 3409 6583
rect 3447 6549 3481 6583
rect 12634 6544 12668 6578
rect 12760 6544 12794 6578
rect 2849 6444 2883 6478
rect 2849 6372 2883 6406
rect 12634 6471 12668 6505
rect 12760 6471 12794 6505
rect 12634 6398 12668 6432
rect 12760 6398 12794 6432
rect 12634 6325 12668 6359
rect 12760 6325 12794 6359
rect 12634 6252 12668 6286
rect 12760 6252 12794 6286
rect 12634 6179 12668 6213
rect 12760 6179 12794 6213
rect 12634 6106 12668 6140
rect 12760 6106 12794 6140
rect 12634 6033 12668 6067
rect 12760 6033 12794 6067
rect 12634 5960 12668 5994
rect 12760 5960 12794 5994
rect 12634 5887 12668 5921
rect 12760 5887 12794 5921
rect 12634 5814 12668 5848
rect 12760 5814 12794 5848
rect 12634 5741 12668 5775
rect 12760 5741 12794 5775
rect 12634 5668 12668 5702
rect 12760 5668 12794 5702
rect 12634 5595 12668 5629
rect 12760 5595 12794 5629
rect 12634 5522 12668 5556
rect 12760 5522 12794 5556
rect 12634 5449 12668 5483
rect 12760 5449 12794 5483
rect 12634 5376 12668 5410
rect 12760 5376 12794 5410
rect 12634 5303 12668 5337
rect 12760 5303 12794 5337
rect 12634 5230 12668 5264
rect 12760 5230 12794 5264
rect 3198 5156 3232 5180
rect 12634 5157 12668 5191
rect 12760 5157 12794 5191
rect 3198 5146 3205 5156
rect 3205 5146 3232 5156
rect 3198 5074 3232 5108
rect 12634 5084 12668 5118
rect 12760 5084 12794 5118
rect 2974 5006 3008 5040
rect 3046 5006 3080 5040
rect 3118 5006 3152 5040
rect 3713 5006 3747 5040
rect 3796 5006 3830 5040
rect 3879 5006 3913 5040
rect 3962 5006 3996 5040
rect 4045 5006 4079 5040
rect 4127 5006 4161 5040
rect 12634 5011 12668 5045
rect 12760 5011 12794 5045
rect 3659 4850 3693 4884
rect 3798 4850 3832 4884
rect 2837 4673 2865 4701
rect 2865 4673 2871 4701
rect 2974 4694 3008 4728
rect 3046 4694 3080 4728
rect 3118 4694 3152 4728
rect 3713 4694 3747 4728
rect 3796 4694 3830 4728
rect 3879 4694 3913 4728
rect 3962 4694 3996 4728
rect 4045 4694 4079 4728
rect 4127 4694 4161 4728
rect 4235 4707 4269 4708
rect 2837 4667 2871 4673
rect 2837 4605 2865 4627
rect 2865 4605 2871 4627
rect 4235 4674 4269 4707
rect 2837 4593 2871 4605
rect 2974 4584 3008 4618
rect 3046 4584 3080 4618
rect 3118 4584 3152 4618
rect 3912 4584 3946 4618
rect 4020 4584 4054 4618
rect 4127 4584 4161 4618
rect 2837 4537 2865 4552
rect 2865 4537 2871 4552
rect 2837 4518 2871 4537
rect 2837 4468 2865 4477
rect 2865 4468 2871 4477
rect 2837 4443 2871 4468
rect 4235 4571 4269 4591
rect 4235 4557 4269 4571
rect 1832 4338 1838 4369
rect 1838 4338 1866 4369
rect 1832 4335 1866 4338
rect 2026 4335 2060 4369
rect 1832 4263 1866 4297
rect 1926 4277 1958 4309
rect 1958 4277 1960 4309
rect 1926 4275 1960 4277
rect 1926 4209 1958 4237
rect 1958 4209 1960 4237
rect 1926 4203 1960 4209
rect 2026 4263 2060 4297
rect 1736 4016 1770 4050
rect 1808 4016 1842 4050
rect 2114 4275 2148 4309
rect 2114 4203 2148 4237
rect 2144 4113 2178 4147
rect 2216 4113 2250 4147
rect 1832 3835 1866 3869
rect 1904 3835 1938 3869
rect 1976 3835 2010 3869
rect 2048 3835 2082 3869
rect 2120 3835 2154 3869
rect 3654 4428 3688 4462
rect 3726 4428 3760 4462
rect 3798 4428 3832 4462
rect 2837 4399 2865 4402
rect 2865 4399 2871 4402
rect 2837 4368 2871 4399
rect 2837 4295 2871 4327
rect 2837 4293 2865 4295
rect 2865 4293 2871 4295
rect 2974 4272 3008 4306
rect 3046 4272 3080 4306
rect 3118 4272 3152 4306
rect 2837 4226 2871 4252
rect 2837 4218 2865 4226
rect 2865 4218 2871 4226
rect 2837 4157 2871 4177
rect 2837 4143 2865 4157
rect 2865 4143 2871 4157
rect 4235 4330 4269 4337
rect 3912 4272 3946 4306
rect 4020 4272 4054 4306
rect 4127 4272 4161 4306
rect 4235 4303 4269 4330
rect 4235 4227 4269 4261
rect 4235 4157 4269 4185
rect 4235 4151 4269 4157
rect 3654 4116 3688 4150
rect 3726 4116 3760 4150
rect 3798 4116 3832 4150
rect 2837 4088 2871 4102
rect 2837 4068 2865 4088
rect 2865 4068 2871 4088
rect 2837 4019 2871 4027
rect 2837 3993 2865 4019
rect 2865 3993 2871 4019
rect 2974 3960 3008 3994
rect 3046 3960 3080 3994
rect 3118 3960 3152 3994
rect 2837 3950 2871 3952
rect 2837 3918 2865 3950
rect 2865 3918 2871 3950
rect 2837 3847 2865 3877
rect 2865 3847 2871 3877
rect 2837 3843 2871 3847
rect 4235 4088 4269 4109
rect 4235 4075 4269 4088
rect 4235 4019 4269 4033
rect 4235 3999 4269 4019
rect 3912 3960 3946 3994
rect 4020 3960 4054 3994
rect 4127 3960 4161 3994
rect 4235 3950 4269 3957
rect 4235 3923 4269 3950
rect 4235 3847 4269 3881
rect 3654 3804 3688 3838
rect 3726 3804 3760 3838
rect 3798 3804 3832 3838
rect 2837 3778 2865 3802
rect 2865 3778 2871 3802
rect 1126 3600 1160 3634
rect 2837 3768 2871 3778
rect 2837 3709 2865 3727
rect 2865 3709 2871 3727
rect 2837 3693 2871 3709
rect 4235 3778 4269 3804
rect 12634 4938 12668 4972
rect 12760 4938 12794 4972
rect 12634 4865 12668 4899
rect 12760 4865 12794 4899
rect 12634 4792 12668 4826
rect 12760 4792 12794 4826
rect 12634 4719 12668 4753
rect 12760 4719 12794 4753
rect 12634 4646 12668 4680
rect 12760 4646 12794 4680
rect 12634 4573 12668 4607
rect 12760 4573 12794 4607
rect 12634 4500 12668 4534
rect 12760 4500 12794 4534
rect 12634 4427 12668 4461
rect 12760 4427 12794 4461
rect 12634 4354 12668 4388
rect 12760 4354 12794 4388
rect 12634 4280 12668 4314
rect 12760 4280 12794 4314
rect 12634 4206 12668 4240
rect 12760 4206 12794 4240
rect 12634 4132 12668 4166
rect 12760 4132 12794 4166
rect 12634 4058 12668 4092
rect 12760 4058 12794 4092
rect 13038 6651 13072 6685
rect 13111 6662 13145 6685
rect 13111 6651 13126 6662
rect 13126 6651 13145 6662
rect 13184 6651 13218 6685
rect 13257 6651 13291 6685
rect 13330 6651 13364 6685
rect 13403 6651 13437 6685
rect 13476 6651 13510 6685
rect 13549 6651 13583 6685
rect 13622 6651 13656 6685
rect 13695 6651 13729 6685
rect 13768 6651 13802 6685
rect 13841 6651 13875 6685
rect 13914 6651 13948 6685
rect 13987 6651 14021 6685
rect 14060 6651 14094 6685
rect 14133 6651 14167 6685
rect 14206 6651 14240 6685
rect 14279 6651 14313 6685
rect 14352 6651 14386 6685
rect 14425 6651 14459 6685
rect 14497 6651 14531 6685
rect 14569 6651 14603 6685
rect 14641 6651 14675 6685
rect 14713 6651 14747 6685
rect 14785 6651 14819 6685
rect 14857 6651 14891 6685
rect 14929 6651 14963 6685
rect 15001 6651 15035 6685
rect 15073 6651 15107 6685
rect 15145 6651 15179 6685
rect 15217 6651 15251 6685
rect 15289 6651 15323 6685
rect 15361 6651 15395 6685
rect 15433 6651 15467 6685
rect 15505 6651 15539 6685
rect 15577 6651 15611 6685
rect 15649 6651 15683 6685
rect 15721 6651 15755 6685
rect 15793 6651 15827 6685
rect 15865 6651 15899 6685
rect 15937 6651 15971 6685
rect 16009 6651 16043 6685
rect 16081 6651 16115 6685
rect 16153 6651 16187 6685
rect 16225 6651 16259 6685
rect 16297 6651 16331 6685
rect 16369 6651 16403 6685
rect 16441 6651 16475 6685
rect 16513 6651 16547 6685
rect 16585 6651 16619 6685
rect 16657 6651 16691 6685
rect 16729 6651 16763 6685
rect 16801 6651 16835 6685
rect 16873 6661 16907 6685
rect 16873 6651 16900 6661
rect 16900 6651 16907 6661
rect 16945 6651 16979 6685
rect 13038 6560 13065 6571
rect 13065 6560 13072 6571
rect 13038 6537 13072 6560
rect 13111 6537 13145 6571
rect 13184 6537 13218 6571
rect 13257 6537 13291 6571
rect 13330 6537 13364 6571
rect 13403 6537 13437 6571
rect 13476 6537 13510 6571
rect 13549 6537 13583 6571
rect 13622 6537 13656 6571
rect 13695 6537 13729 6571
rect 13768 6537 13802 6571
rect 13841 6537 13875 6571
rect 13914 6537 13948 6571
rect 13987 6537 14021 6571
rect 14060 6537 14094 6571
rect 14133 6537 14167 6571
rect 14206 6537 14240 6571
rect 14279 6537 14313 6571
rect 14352 6537 14386 6571
rect 14425 6537 14459 6571
rect 14497 6537 14531 6571
rect 14569 6537 14603 6571
rect 14641 6537 14675 6571
rect 14713 6537 14747 6571
rect 14785 6537 14819 6571
rect 14857 6537 14891 6571
rect 14929 6537 14963 6571
rect 15001 6537 15035 6571
rect 15073 6537 15107 6571
rect 15145 6537 15179 6571
rect 15217 6537 15251 6571
rect 15289 6537 15323 6571
rect 15361 6537 15395 6571
rect 15433 6537 15467 6571
rect 15505 6537 15539 6571
rect 15577 6537 15611 6571
rect 15649 6537 15683 6571
rect 15721 6537 15755 6571
rect 15793 6537 15827 6571
rect 15865 6537 15899 6571
rect 15937 6537 15971 6571
rect 16009 6537 16043 6571
rect 16081 6537 16115 6571
rect 16153 6537 16187 6571
rect 16225 6537 16259 6571
rect 16297 6537 16331 6571
rect 16369 6537 16403 6571
rect 16441 6537 16475 6571
rect 16513 6537 16547 6571
rect 16585 6537 16619 6571
rect 16657 6537 16691 6571
rect 16729 6537 16763 6571
rect 16801 6537 16835 6571
rect 16873 6537 16907 6571
rect 16945 6559 16961 6571
rect 16961 6559 16979 6571
rect 16945 6537 16979 6559
rect 13032 6456 13066 6490
rect 13146 6456 13180 6490
rect 13032 6384 13066 6418
rect 13146 6384 13180 6418
rect 16837 6456 16871 6490
rect 16951 6456 16985 6490
rect 13032 6312 13066 6346
rect 13146 6312 13180 6346
rect 13032 6240 13066 6274
rect 13146 6240 13180 6274
rect 13032 6168 13066 6202
rect 13146 6168 13180 6202
rect 13032 6096 13066 6130
rect 13146 6096 13180 6130
rect 13032 6024 13066 6058
rect 13146 6024 13180 6058
rect 13032 5952 13066 5986
rect 13146 5952 13180 5986
rect 13032 5880 13066 5914
rect 13146 5880 13180 5914
rect 13032 5808 13066 5842
rect 13146 5808 13180 5842
rect 13032 5736 13066 5770
rect 13146 5736 13180 5770
rect 13032 5664 13066 5698
rect 13146 5664 13180 5698
rect 13032 5592 13066 5626
rect 13146 5592 13180 5626
rect 13032 5520 13066 5554
rect 13146 5520 13180 5554
rect 13032 5448 13066 5482
rect 13146 5448 13180 5482
rect 13032 5376 13066 5410
rect 13146 5376 13180 5410
rect 13032 5304 13066 5338
rect 13146 5304 13180 5338
rect 13032 5232 13066 5266
rect 13146 5232 13180 5266
rect 13032 5160 13066 5194
rect 13146 5160 13180 5194
rect 13032 5088 13066 5122
rect 13146 5088 13180 5122
rect 13032 5016 13066 5050
rect 13146 5016 13180 5050
rect 13032 4944 13066 4978
rect 13146 4944 13180 4978
rect 13032 4872 13066 4906
rect 13146 4872 13180 4906
rect 13032 4800 13066 4834
rect 13146 4800 13180 4834
rect 13032 4728 13066 4762
rect 13146 4728 13180 4762
rect 13032 4656 13066 4690
rect 13146 4656 13180 4690
rect 13032 4584 13066 4618
rect 13146 4584 13180 4618
rect 13032 4512 13066 4546
rect 13146 4512 13180 4546
rect 13032 4440 13066 4474
rect 13146 4440 13180 4474
rect 13032 4368 13066 4402
rect 13146 4368 13180 4402
rect 13404 6357 13438 6391
rect 13476 6383 13510 6391
rect 13476 6357 13508 6383
rect 13508 6357 13510 6383
rect 13548 6383 13582 6391
rect 13620 6383 13654 6391
rect 13692 6383 13726 6391
rect 13764 6383 13798 6391
rect 13836 6383 13870 6391
rect 13908 6383 13942 6391
rect 13980 6383 14014 6391
rect 14052 6383 14086 6391
rect 14124 6383 14158 6391
rect 14196 6383 14230 6391
rect 14268 6383 14302 6391
rect 14340 6383 14374 6391
rect 14412 6383 14446 6391
rect 14484 6383 14518 6391
rect 14556 6383 14590 6391
rect 14628 6383 14662 6391
rect 14700 6383 14734 6391
rect 14772 6383 14806 6391
rect 14844 6383 14878 6391
rect 14916 6383 14950 6391
rect 14988 6383 15022 6391
rect 15060 6383 15094 6391
rect 15132 6383 15166 6391
rect 15204 6383 15238 6391
rect 15276 6383 15310 6391
rect 15348 6383 15382 6391
rect 15420 6383 15454 6391
rect 15492 6383 15526 6391
rect 15564 6383 15598 6391
rect 15636 6383 15670 6391
rect 13548 6357 13556 6383
rect 13556 6357 13582 6383
rect 13620 6357 13624 6383
rect 13624 6357 13654 6383
rect 13692 6357 13726 6383
rect 13764 6357 13794 6383
rect 13794 6357 13798 6383
rect 13836 6357 13862 6383
rect 13862 6357 13870 6383
rect 13908 6357 13930 6383
rect 13930 6357 13942 6383
rect 13980 6357 13998 6383
rect 13998 6357 14014 6383
rect 14052 6357 14066 6383
rect 14066 6357 14086 6383
rect 14124 6357 14134 6383
rect 14134 6357 14158 6383
rect 14196 6357 14202 6383
rect 14202 6357 14230 6383
rect 14268 6357 14270 6383
rect 14270 6357 14302 6383
rect 14340 6357 14372 6383
rect 14372 6357 14374 6383
rect 14412 6357 14440 6383
rect 14440 6357 14446 6383
rect 14484 6357 14508 6383
rect 14508 6357 14518 6383
rect 14556 6357 14576 6383
rect 14576 6357 14590 6383
rect 14628 6357 14644 6383
rect 14644 6357 14662 6383
rect 14700 6357 14712 6383
rect 14712 6357 14734 6383
rect 14772 6357 14780 6383
rect 14780 6357 14806 6383
rect 14844 6357 14848 6383
rect 14848 6357 14878 6383
rect 14916 6357 14950 6383
rect 14988 6357 15018 6383
rect 15018 6357 15022 6383
rect 15060 6357 15087 6383
rect 15087 6357 15094 6383
rect 15132 6357 15156 6383
rect 15156 6357 15166 6383
rect 15204 6357 15225 6383
rect 15225 6357 15238 6383
rect 15276 6357 15294 6383
rect 15294 6357 15310 6383
rect 15348 6357 15363 6383
rect 15363 6357 15382 6383
rect 15420 6357 15432 6383
rect 15432 6357 15454 6383
rect 15492 6357 15501 6383
rect 15501 6357 15526 6383
rect 15564 6357 15570 6383
rect 15570 6357 15598 6383
rect 15636 6357 15639 6383
rect 15639 6357 15670 6383
rect 15708 6357 15742 6391
rect 15780 6383 15814 6391
rect 15852 6383 15886 6391
rect 15924 6383 15958 6391
rect 15996 6383 16030 6391
rect 16068 6383 16102 6391
rect 16140 6383 16174 6391
rect 16213 6383 16247 6391
rect 16286 6383 16320 6391
rect 16359 6383 16393 6391
rect 16432 6383 16466 6391
rect 16505 6383 16539 6391
rect 15780 6357 15812 6383
rect 15812 6357 15814 6383
rect 15852 6357 15881 6383
rect 15881 6357 15886 6383
rect 15924 6357 15950 6383
rect 15950 6357 15958 6383
rect 15996 6357 16019 6383
rect 16019 6357 16030 6383
rect 16068 6357 16088 6383
rect 16088 6357 16102 6383
rect 16140 6357 16157 6383
rect 16157 6357 16174 6383
rect 16213 6357 16226 6383
rect 16226 6357 16247 6383
rect 16286 6357 16295 6383
rect 16295 6357 16320 6383
rect 16359 6357 16364 6383
rect 16364 6357 16393 6383
rect 16432 6357 16433 6383
rect 16433 6357 16466 6383
rect 16505 6357 16536 6383
rect 16536 6357 16539 6383
rect 16578 6357 16612 6391
rect 13332 6285 13366 6319
rect 16650 6315 16683 6319
rect 16683 6315 16684 6319
rect 13332 6245 13366 6246
rect 13332 6212 13366 6245
rect 13332 6141 13366 6173
rect 13332 6139 13366 6141
rect 13332 6072 13366 6100
rect 13332 6066 13366 6072
rect 13332 6003 13366 6027
rect 13332 5993 13366 6003
rect 13530 6253 13564 6287
rect 13603 6253 13637 6287
rect 13676 6253 13710 6287
rect 13749 6253 13783 6287
rect 13822 6253 13856 6287
rect 13895 6253 13929 6287
rect 13968 6253 14002 6287
rect 14041 6253 14075 6287
rect 14114 6253 14148 6287
rect 14187 6253 14221 6287
rect 14260 6253 14294 6287
rect 14333 6253 14367 6287
rect 14406 6253 14440 6287
rect 14479 6253 14513 6287
rect 14552 6253 14586 6287
rect 14625 6253 14659 6287
rect 14698 6253 14732 6287
rect 14771 6253 14805 6287
rect 14844 6253 14878 6287
rect 14917 6253 14951 6287
rect 14990 6253 15024 6287
rect 15063 6253 15097 6287
rect 15136 6253 15170 6287
rect 15209 6253 15243 6287
rect 15282 6253 15316 6287
rect 15355 6253 15389 6287
rect 15427 6253 15461 6287
rect 15499 6253 15533 6287
rect 15571 6253 15605 6287
rect 15643 6253 15677 6287
rect 15715 6253 15749 6287
rect 15787 6253 15821 6287
rect 15859 6253 15893 6287
rect 15931 6253 15965 6287
rect 16003 6253 16037 6287
rect 16075 6253 16109 6287
rect 16147 6253 16181 6287
rect 16219 6253 16253 6287
rect 16291 6253 16325 6287
rect 16650 6285 16684 6315
rect 13450 6243 13484 6247
rect 13450 6213 13484 6243
rect 13450 6169 13484 6171
rect 13450 6137 13484 6169
rect 16650 6245 16683 6247
rect 16683 6245 16684 6247
rect 16650 6213 16684 6245
rect 16650 6141 16684 6175
rect 13770 6097 13804 6131
rect 13844 6097 13878 6131
rect 13918 6097 13952 6131
rect 13992 6097 14026 6131
rect 14066 6097 14100 6131
rect 14140 6097 14174 6131
rect 14214 6097 14248 6131
rect 14288 6097 14322 6131
rect 14362 6097 14396 6131
rect 14436 6097 14470 6131
rect 14510 6097 14544 6131
rect 14584 6097 14618 6131
rect 14658 6097 14692 6131
rect 14732 6097 14766 6131
rect 14806 6097 14840 6131
rect 14880 6097 14914 6131
rect 14954 6097 14988 6131
rect 15028 6097 15062 6131
rect 15102 6097 15136 6131
rect 15176 6097 15210 6131
rect 15250 6097 15284 6131
rect 15323 6097 15357 6131
rect 15396 6097 15430 6131
rect 15469 6097 15503 6131
rect 15542 6097 15576 6131
rect 15615 6097 15649 6131
rect 15688 6097 15722 6131
rect 15761 6097 15795 6131
rect 15834 6097 15868 6131
rect 15907 6097 15941 6131
rect 15980 6097 16014 6131
rect 16053 6097 16087 6131
rect 16126 6097 16160 6131
rect 16199 6097 16233 6131
rect 16272 6097 16306 6131
rect 16345 6097 16379 6131
rect 16418 6097 16452 6131
rect 13450 6094 13484 6095
rect 13450 6061 13484 6094
rect 13450 5985 13484 6018
rect 13450 5984 13484 5985
rect 16650 6069 16684 6103
rect 16650 5999 16684 6031
rect 16650 5997 16683 5999
rect 16683 5997 16684 5999
rect 13332 5934 13366 5954
rect 13530 5941 13564 5975
rect 13603 5941 13637 5975
rect 13676 5941 13710 5975
rect 13749 5941 13783 5975
rect 13822 5941 13856 5975
rect 13895 5941 13929 5975
rect 13968 5941 14002 5975
rect 14041 5941 14075 5975
rect 14114 5941 14148 5975
rect 14187 5941 14221 5975
rect 14260 5941 14294 5975
rect 14333 5941 14367 5975
rect 14406 5941 14440 5975
rect 14479 5941 14513 5975
rect 14552 5941 14586 5975
rect 14625 5941 14659 5975
rect 14698 5941 14732 5975
rect 14771 5941 14805 5975
rect 14844 5941 14878 5975
rect 14917 5941 14951 5975
rect 14990 5941 15024 5975
rect 15063 5941 15097 5975
rect 15136 5941 15170 5975
rect 15209 5941 15243 5975
rect 15282 5941 15316 5975
rect 15355 5941 15389 5975
rect 15427 5941 15461 5975
rect 15499 5941 15533 5975
rect 15571 5941 15605 5975
rect 15643 5941 15677 5975
rect 15715 5941 15749 5975
rect 15787 5941 15821 5975
rect 15859 5941 15893 5975
rect 15931 5941 15965 5975
rect 16003 5941 16037 5975
rect 16075 5941 16109 5975
rect 16147 5941 16181 5975
rect 16219 5941 16253 5975
rect 16291 5941 16325 5975
rect 13332 5920 13366 5934
rect 13332 5865 13366 5881
rect 16650 5929 16684 5959
rect 16650 5925 16683 5929
rect 16683 5925 16684 5929
rect 13332 5847 13366 5865
rect 13819 5845 13849 5879
rect 13849 5845 13853 5879
rect 13892 5845 13917 5879
rect 13917 5845 13926 5879
rect 13965 5845 13985 5879
rect 13985 5845 13999 5879
rect 14038 5845 14053 5879
rect 14053 5845 14072 5879
rect 14111 5845 14121 5879
rect 14121 5845 14145 5879
rect 14184 5845 14189 5879
rect 14189 5845 14218 5879
rect 14257 5845 14291 5879
rect 14330 5845 14359 5879
rect 14359 5845 14364 5879
rect 14403 5845 14427 5879
rect 14427 5845 14437 5879
rect 14476 5845 14495 5879
rect 14495 5845 14510 5879
rect 14549 5845 14563 5879
rect 14563 5845 14583 5879
rect 14622 5845 14631 5879
rect 14631 5845 14656 5879
rect 14695 5845 14699 5879
rect 14699 5845 14729 5879
rect 14768 5845 14801 5879
rect 14801 5845 14802 5879
rect 14841 5845 14869 5879
rect 14869 5845 14875 5879
rect 14914 5845 14937 5879
rect 14937 5845 14948 5879
rect 14987 5845 15005 5879
rect 15005 5845 15021 5879
rect 15060 5845 15073 5879
rect 15073 5845 15094 5879
rect 15133 5845 15141 5879
rect 15141 5845 15167 5879
rect 15206 5845 15209 5879
rect 15209 5845 15240 5879
rect 15279 5845 15311 5879
rect 15311 5845 15313 5879
rect 15352 5845 15379 5879
rect 15379 5845 15386 5879
rect 15425 5845 15447 5879
rect 15447 5845 15459 5879
rect 15498 5845 15515 5879
rect 15515 5845 15532 5879
rect 15571 5845 15583 5879
rect 15583 5845 15605 5879
rect 15644 5845 15651 5879
rect 15651 5845 15678 5879
rect 15717 5845 15719 5879
rect 15719 5845 15751 5879
rect 15789 5845 15821 5879
rect 15821 5845 15823 5879
rect 15861 5845 15889 5879
rect 15889 5845 15895 5879
rect 15933 5845 15957 5879
rect 15957 5845 15967 5879
rect 16005 5845 16025 5879
rect 16025 5845 16039 5879
rect 16077 5845 16093 5879
rect 16093 5845 16111 5879
rect 16149 5845 16161 5879
rect 16161 5845 16183 5879
rect 16221 5845 16229 5879
rect 16229 5845 16255 5879
rect 16293 5845 16297 5879
rect 16297 5845 16327 5879
rect 16650 5859 16684 5887
rect 16650 5853 16683 5859
rect 16683 5853 16684 5859
rect 13332 5796 13366 5808
rect 13332 5774 13366 5796
rect 16650 5789 16684 5815
rect 13332 5727 13366 5735
rect 13332 5701 13366 5727
rect 13332 5658 13366 5662
rect 13332 5628 13366 5658
rect 13332 5589 13366 5590
rect 13332 5556 13366 5589
rect 13332 5486 13366 5518
rect 13332 5484 13366 5486
rect 13530 5749 13564 5783
rect 13603 5749 13637 5783
rect 13676 5749 13710 5783
rect 13749 5749 13783 5783
rect 13822 5749 13856 5783
rect 13895 5749 13929 5783
rect 13968 5749 14002 5783
rect 14041 5749 14075 5783
rect 14114 5749 14148 5783
rect 14187 5749 14221 5783
rect 14260 5749 14294 5783
rect 14333 5749 14367 5783
rect 14406 5749 14440 5783
rect 14479 5749 14513 5783
rect 14552 5749 14586 5783
rect 14625 5749 14659 5783
rect 14698 5749 14732 5783
rect 14771 5749 14805 5783
rect 14844 5749 14878 5783
rect 14917 5749 14951 5783
rect 14990 5749 15024 5783
rect 15063 5749 15097 5783
rect 15136 5749 15170 5783
rect 15209 5749 15243 5783
rect 15282 5749 15316 5783
rect 15355 5749 15389 5783
rect 15427 5749 15461 5783
rect 15499 5749 15533 5783
rect 15571 5749 15605 5783
rect 15643 5749 15677 5783
rect 15715 5749 15749 5783
rect 15787 5749 15821 5783
rect 15859 5749 15893 5783
rect 15931 5749 15965 5783
rect 16003 5749 16037 5783
rect 16075 5749 16109 5783
rect 16147 5749 16181 5783
rect 16219 5749 16253 5783
rect 16291 5749 16325 5783
rect 16650 5781 16683 5789
rect 16683 5781 16684 5789
rect 13450 5739 13484 5743
rect 13450 5709 13484 5739
rect 13450 5665 13484 5667
rect 13450 5633 13484 5665
rect 16650 5719 16684 5743
rect 16650 5709 16683 5719
rect 16683 5709 16684 5719
rect 16650 5649 16684 5671
rect 16650 5637 16683 5649
rect 16683 5637 16684 5649
rect 13770 5593 13804 5627
rect 13844 5593 13878 5627
rect 13918 5593 13952 5627
rect 13992 5593 14026 5627
rect 14066 5593 14100 5627
rect 14140 5593 14174 5627
rect 14214 5593 14248 5627
rect 14288 5593 14322 5627
rect 14362 5593 14396 5627
rect 14436 5593 14470 5627
rect 14510 5593 14544 5627
rect 14584 5593 14618 5627
rect 14658 5593 14692 5627
rect 14732 5593 14766 5627
rect 14806 5593 14840 5627
rect 14880 5593 14914 5627
rect 14954 5593 14988 5627
rect 15028 5593 15062 5627
rect 15102 5593 15136 5627
rect 15176 5593 15210 5627
rect 15250 5593 15284 5627
rect 15323 5593 15357 5627
rect 15396 5593 15430 5627
rect 15469 5593 15503 5627
rect 15542 5593 15576 5627
rect 15615 5593 15649 5627
rect 15688 5593 15722 5627
rect 15761 5593 15795 5627
rect 15834 5593 15868 5627
rect 15907 5593 15941 5627
rect 15980 5593 16014 5627
rect 16053 5593 16087 5627
rect 16126 5593 16160 5627
rect 16199 5593 16233 5627
rect 16272 5593 16306 5627
rect 16345 5593 16379 5627
rect 16418 5593 16452 5627
rect 13450 5590 13484 5591
rect 13450 5557 13484 5590
rect 13450 5481 13484 5514
rect 13450 5480 13484 5481
rect 16650 5579 16684 5599
rect 16650 5565 16683 5579
rect 16683 5565 16684 5579
rect 16650 5509 16684 5527
rect 16650 5493 16683 5509
rect 16683 5493 16684 5509
rect 13332 5417 13366 5446
rect 13530 5437 13564 5471
rect 13603 5437 13637 5471
rect 13676 5437 13710 5471
rect 13749 5437 13783 5471
rect 13822 5437 13856 5471
rect 13895 5437 13929 5471
rect 13968 5437 14002 5471
rect 14041 5437 14075 5471
rect 14114 5437 14148 5471
rect 14187 5437 14221 5471
rect 14260 5437 14294 5471
rect 14333 5437 14367 5471
rect 14406 5437 14440 5471
rect 14479 5437 14513 5471
rect 14552 5437 14586 5471
rect 14625 5437 14659 5471
rect 14698 5437 14732 5471
rect 14771 5437 14805 5471
rect 14844 5437 14878 5471
rect 14917 5437 14951 5471
rect 14990 5437 15024 5471
rect 15063 5437 15097 5471
rect 15136 5437 15170 5471
rect 15209 5437 15243 5471
rect 15282 5437 15316 5471
rect 15355 5437 15389 5471
rect 15427 5437 15461 5471
rect 15499 5437 15533 5471
rect 15571 5437 15605 5471
rect 15643 5437 15677 5471
rect 15715 5437 15749 5471
rect 15787 5437 15821 5471
rect 15859 5437 15893 5471
rect 15931 5437 15965 5471
rect 16003 5437 16037 5471
rect 16075 5437 16109 5471
rect 16147 5437 16181 5471
rect 16219 5437 16253 5471
rect 16291 5437 16325 5471
rect 16650 5439 16684 5455
rect 13332 5412 13366 5417
rect 16650 5421 16683 5439
rect 16683 5421 16684 5439
rect 13332 5347 13366 5374
rect 13332 5340 13366 5347
rect 13819 5341 13849 5375
rect 13849 5341 13853 5375
rect 13892 5341 13917 5375
rect 13917 5341 13926 5375
rect 13965 5341 13985 5375
rect 13985 5341 13999 5375
rect 14038 5341 14053 5375
rect 14053 5341 14072 5375
rect 14111 5341 14121 5375
rect 14121 5341 14145 5375
rect 14184 5341 14189 5375
rect 14189 5341 14218 5375
rect 14257 5341 14291 5375
rect 14330 5341 14359 5375
rect 14359 5341 14364 5375
rect 14403 5341 14427 5375
rect 14427 5341 14437 5375
rect 14476 5341 14495 5375
rect 14495 5341 14510 5375
rect 14549 5341 14563 5375
rect 14563 5341 14583 5375
rect 14622 5341 14631 5375
rect 14631 5341 14656 5375
rect 14695 5341 14699 5375
rect 14699 5341 14729 5375
rect 14768 5341 14801 5375
rect 14801 5341 14802 5375
rect 14841 5341 14869 5375
rect 14869 5341 14875 5375
rect 14914 5341 14937 5375
rect 14937 5341 14948 5375
rect 14987 5341 15005 5375
rect 15005 5341 15021 5375
rect 15060 5341 15073 5375
rect 15073 5341 15094 5375
rect 15133 5341 15141 5375
rect 15141 5341 15167 5375
rect 15206 5341 15209 5375
rect 15209 5341 15240 5375
rect 15279 5341 15311 5375
rect 15311 5341 15313 5375
rect 15352 5341 15379 5375
rect 15379 5341 15386 5375
rect 15425 5341 15447 5375
rect 15447 5341 15459 5375
rect 15498 5341 15515 5375
rect 15515 5341 15532 5375
rect 15571 5341 15583 5375
rect 15583 5341 15605 5375
rect 15644 5341 15651 5375
rect 15651 5341 15678 5375
rect 15717 5341 15719 5375
rect 15719 5341 15751 5375
rect 15789 5341 15821 5375
rect 15821 5341 15823 5375
rect 15861 5341 15889 5375
rect 15889 5341 15895 5375
rect 15933 5341 15957 5375
rect 15957 5341 15967 5375
rect 16005 5341 16025 5375
rect 16025 5341 16039 5375
rect 16077 5341 16093 5375
rect 16093 5341 16111 5375
rect 16149 5341 16161 5375
rect 16161 5341 16183 5375
rect 16221 5341 16229 5375
rect 16229 5341 16255 5375
rect 16293 5341 16297 5375
rect 16297 5341 16327 5375
rect 16650 5369 16684 5383
rect 16650 5349 16683 5369
rect 16683 5349 16684 5369
rect 13332 5277 13366 5302
rect 16650 5299 16684 5311
rect 13332 5268 13366 5277
rect 13332 5207 13366 5230
rect 13332 5196 13366 5207
rect 13332 5137 13366 5158
rect 13332 5124 13366 5137
rect 13332 5067 13366 5086
rect 13332 5052 13366 5067
rect 13332 4997 13366 5014
rect 13332 4980 13366 4997
rect 13530 5245 13564 5279
rect 13603 5245 13637 5279
rect 13676 5245 13710 5279
rect 13749 5245 13783 5279
rect 13822 5245 13856 5279
rect 13895 5245 13929 5279
rect 13968 5245 14002 5279
rect 14041 5245 14075 5279
rect 14114 5245 14148 5279
rect 14187 5245 14221 5279
rect 14260 5245 14294 5279
rect 14333 5245 14367 5279
rect 14406 5245 14440 5279
rect 14479 5245 14513 5279
rect 14552 5245 14586 5279
rect 14625 5245 14659 5279
rect 14698 5245 14732 5279
rect 14771 5245 14805 5279
rect 14844 5245 14878 5279
rect 14917 5245 14951 5279
rect 14990 5245 15024 5279
rect 15063 5245 15097 5279
rect 15136 5245 15170 5279
rect 15209 5245 15243 5279
rect 15282 5245 15316 5279
rect 15355 5245 15389 5279
rect 15428 5245 15462 5279
rect 15501 5245 15535 5279
rect 15573 5245 15607 5279
rect 15645 5245 15679 5279
rect 15717 5245 15751 5279
rect 15789 5245 15823 5279
rect 15861 5245 15895 5279
rect 15933 5245 15967 5279
rect 16005 5245 16039 5279
rect 16077 5245 16111 5279
rect 16149 5245 16183 5279
rect 16221 5245 16255 5279
rect 16293 5245 16327 5279
rect 16650 5277 16683 5299
rect 16683 5277 16684 5299
rect 13450 5235 13484 5239
rect 13450 5205 13484 5235
rect 13450 5161 13484 5163
rect 13450 5129 13484 5161
rect 16650 5230 16684 5239
rect 16650 5205 16683 5230
rect 16683 5205 16684 5230
rect 16650 5161 16684 5167
rect 16650 5133 16683 5161
rect 16683 5133 16684 5161
rect 13770 5089 13804 5123
rect 13844 5089 13878 5123
rect 13918 5089 13952 5123
rect 13992 5089 14026 5123
rect 14066 5089 14100 5123
rect 14140 5089 14174 5123
rect 14214 5089 14248 5123
rect 14288 5089 14322 5123
rect 14362 5089 14396 5123
rect 14436 5089 14470 5123
rect 14510 5089 14544 5123
rect 14583 5089 14617 5123
rect 14656 5089 14690 5123
rect 14729 5089 14763 5123
rect 14802 5089 14836 5123
rect 14875 5089 14909 5123
rect 14948 5089 14982 5123
rect 15021 5089 15055 5123
rect 15094 5089 15128 5123
rect 15167 5089 15201 5123
rect 15240 5089 15274 5123
rect 15313 5089 15347 5123
rect 15386 5089 15420 5123
rect 15459 5089 15493 5123
rect 15532 5089 15566 5123
rect 15605 5089 15639 5123
rect 15678 5089 15712 5123
rect 15751 5089 15785 5123
rect 15824 5089 15858 5123
rect 15897 5089 15931 5123
rect 15970 5089 16004 5123
rect 16043 5089 16077 5123
rect 16116 5089 16150 5123
rect 16189 5089 16223 5123
rect 16262 5089 16296 5123
rect 16335 5089 16369 5123
rect 16408 5089 16442 5123
rect 16650 5092 16684 5095
rect 13450 5086 13484 5087
rect 13450 5053 13484 5086
rect 13450 4977 13484 5010
rect 13450 4976 13484 4977
rect 16650 5061 16683 5092
rect 16683 5061 16684 5092
rect 16650 4989 16683 5022
rect 16683 4989 16684 5022
rect 16650 4988 16684 4989
rect 13332 4927 13366 4942
rect 13530 4933 13564 4967
rect 13603 4933 13637 4967
rect 13676 4933 13710 4967
rect 13749 4933 13783 4967
rect 13822 4933 13856 4967
rect 13895 4933 13929 4967
rect 13968 4933 14002 4967
rect 14041 4933 14075 4967
rect 14114 4933 14148 4967
rect 14187 4933 14221 4967
rect 14260 4933 14294 4967
rect 14333 4933 14367 4967
rect 14406 4933 14440 4967
rect 14479 4933 14513 4967
rect 14552 4933 14586 4967
rect 14625 4933 14659 4967
rect 14698 4933 14732 4967
rect 14771 4933 14805 4967
rect 14844 4933 14878 4967
rect 14917 4933 14951 4967
rect 14990 4933 15024 4967
rect 15063 4933 15097 4967
rect 15136 4933 15170 4967
rect 15209 4933 15243 4967
rect 15282 4933 15316 4967
rect 15355 4933 15389 4967
rect 15428 4933 15462 4967
rect 15501 4933 15535 4967
rect 15573 4933 15607 4967
rect 15645 4933 15679 4967
rect 15717 4933 15751 4967
rect 15789 4933 15823 4967
rect 15861 4933 15895 4967
rect 15933 4933 15967 4967
rect 16005 4933 16039 4967
rect 16077 4933 16111 4967
rect 16149 4933 16183 4967
rect 16221 4933 16255 4967
rect 16293 4933 16327 4967
rect 13332 4908 13366 4927
rect 16650 4920 16683 4949
rect 16683 4920 16684 4949
rect 16650 4915 16684 4920
rect 13332 4857 13366 4870
rect 13332 4836 13366 4857
rect 13819 4837 13849 4871
rect 13849 4837 13853 4871
rect 13892 4837 13917 4871
rect 13917 4837 13926 4871
rect 13965 4837 13985 4871
rect 13985 4837 13999 4871
rect 14038 4837 14053 4871
rect 14053 4837 14072 4871
rect 14111 4837 14121 4871
rect 14121 4837 14145 4871
rect 14184 4837 14189 4871
rect 14189 4837 14218 4871
rect 14257 4837 14291 4871
rect 14330 4837 14359 4871
rect 14359 4837 14364 4871
rect 14403 4837 14427 4871
rect 14427 4837 14437 4871
rect 14476 4837 14495 4871
rect 14495 4837 14510 4871
rect 14549 4837 14563 4871
rect 14563 4837 14583 4871
rect 14622 4837 14631 4871
rect 14631 4837 14656 4871
rect 14695 4837 14699 4871
rect 14699 4837 14729 4871
rect 14768 4837 14801 4871
rect 14801 4837 14802 4871
rect 14841 4837 14869 4871
rect 14869 4837 14875 4871
rect 14914 4837 14937 4871
rect 14937 4837 14948 4871
rect 14987 4837 15005 4871
rect 15005 4837 15021 4871
rect 15060 4837 15073 4871
rect 15073 4837 15094 4871
rect 15133 4837 15141 4871
rect 15141 4837 15167 4871
rect 15206 4837 15209 4871
rect 15209 4837 15240 4871
rect 15279 4837 15311 4871
rect 15311 4837 15313 4871
rect 15352 4837 15379 4871
rect 15379 4837 15386 4871
rect 15425 4837 15447 4871
rect 15447 4837 15459 4871
rect 15498 4837 15515 4871
rect 15515 4837 15532 4871
rect 15571 4837 15583 4871
rect 15583 4837 15605 4871
rect 15644 4837 15651 4871
rect 15651 4837 15678 4871
rect 15717 4837 15719 4871
rect 15719 4837 15751 4871
rect 15789 4837 15821 4871
rect 15821 4837 15823 4871
rect 15861 4837 15889 4871
rect 15889 4837 15895 4871
rect 15933 4837 15957 4871
rect 15957 4837 15967 4871
rect 16005 4837 16025 4871
rect 16025 4837 16039 4871
rect 16077 4837 16093 4871
rect 16093 4837 16111 4871
rect 16149 4837 16161 4871
rect 16161 4837 16183 4871
rect 16221 4837 16229 4871
rect 16229 4837 16255 4871
rect 16293 4837 16297 4871
rect 16297 4837 16327 4871
rect 16650 4851 16683 4876
rect 16683 4851 16684 4876
rect 16650 4842 16684 4851
rect 13332 4787 13366 4798
rect 13332 4764 13366 4787
rect 16650 4782 16683 4803
rect 16683 4782 16684 4803
rect 13332 4717 13366 4726
rect 13332 4692 13366 4717
rect 13332 4647 13366 4654
rect 13332 4620 13366 4647
rect 13332 4577 13366 4582
rect 13332 4548 13366 4577
rect 13332 4507 13366 4510
rect 13332 4476 13366 4507
rect 13530 4741 13564 4775
rect 13603 4741 13637 4775
rect 13676 4741 13710 4775
rect 13749 4741 13783 4775
rect 13822 4741 13856 4775
rect 13895 4741 13929 4775
rect 13968 4741 14002 4775
rect 14041 4741 14075 4775
rect 14114 4741 14148 4775
rect 14187 4741 14221 4775
rect 14260 4741 14294 4775
rect 14333 4741 14367 4775
rect 14406 4741 14440 4775
rect 14479 4741 14513 4775
rect 14552 4741 14586 4775
rect 14625 4741 14659 4775
rect 14698 4741 14732 4775
rect 14771 4741 14805 4775
rect 14844 4741 14878 4775
rect 14917 4741 14951 4775
rect 14990 4741 15024 4775
rect 15063 4741 15097 4775
rect 15136 4741 15170 4775
rect 15209 4741 15243 4775
rect 15282 4741 15316 4775
rect 15355 4741 15389 4775
rect 15428 4741 15462 4775
rect 15501 4741 15535 4775
rect 15573 4741 15607 4775
rect 15645 4741 15679 4775
rect 15717 4741 15751 4775
rect 15789 4741 15823 4775
rect 15861 4741 15895 4775
rect 15933 4741 15967 4775
rect 16005 4741 16039 4775
rect 16077 4741 16111 4775
rect 16149 4741 16183 4775
rect 16221 4741 16255 4775
rect 16293 4741 16327 4775
rect 16650 4769 16684 4782
rect 13450 4731 13484 4735
rect 13450 4701 13484 4731
rect 13450 4657 13484 4659
rect 13450 4625 13484 4657
rect 16650 4713 16683 4730
rect 16683 4713 16684 4730
rect 16650 4696 16684 4713
rect 16650 4644 16683 4657
rect 16683 4644 16684 4657
rect 16650 4623 16684 4644
rect 13770 4585 13804 4619
rect 13844 4585 13878 4619
rect 13918 4585 13952 4619
rect 13992 4585 14026 4619
rect 14066 4585 14100 4619
rect 14140 4585 14174 4619
rect 14214 4585 14248 4619
rect 14288 4585 14322 4619
rect 14362 4585 14396 4619
rect 14435 4585 14469 4619
rect 14508 4585 14542 4619
rect 14581 4585 14615 4619
rect 14654 4585 14688 4619
rect 14727 4585 14761 4619
rect 14800 4585 14834 4619
rect 14873 4585 14907 4619
rect 14946 4585 14980 4619
rect 15019 4585 15053 4619
rect 15092 4585 15126 4619
rect 15165 4585 15199 4619
rect 15238 4585 15272 4619
rect 15311 4585 15345 4619
rect 15384 4585 15418 4619
rect 15457 4585 15491 4619
rect 15530 4585 15564 4619
rect 15603 4585 15637 4619
rect 15676 4585 15710 4619
rect 15749 4585 15783 4619
rect 15822 4585 15856 4619
rect 15895 4585 15929 4619
rect 15968 4585 16002 4619
rect 16041 4585 16075 4619
rect 16114 4585 16148 4619
rect 16187 4585 16221 4619
rect 16260 4585 16294 4619
rect 16333 4585 16367 4619
rect 16406 4585 16440 4619
rect 13450 4548 13484 4582
rect 13450 4473 13484 4505
rect 13450 4471 13484 4473
rect 16650 4575 16683 4584
rect 16683 4575 16684 4584
rect 16650 4550 16684 4575
rect 16650 4506 16683 4511
rect 16683 4506 16684 4511
rect 16650 4477 16684 4506
rect 13332 4437 13366 4438
rect 13332 4404 13366 4437
rect 13530 4429 13564 4463
rect 13603 4429 13637 4463
rect 13676 4429 13710 4463
rect 13749 4429 13783 4463
rect 13822 4429 13856 4463
rect 13895 4429 13929 4463
rect 13968 4429 14002 4463
rect 14041 4429 14075 4463
rect 14114 4429 14148 4463
rect 14187 4429 14221 4463
rect 14260 4429 14294 4463
rect 14333 4429 14367 4463
rect 14406 4429 14440 4463
rect 14479 4429 14513 4463
rect 14552 4429 14586 4463
rect 14625 4429 14659 4463
rect 14698 4429 14732 4463
rect 14771 4429 14805 4463
rect 14844 4429 14878 4463
rect 14917 4429 14951 4463
rect 14990 4429 15024 4463
rect 15063 4429 15097 4463
rect 15136 4429 15170 4463
rect 15209 4429 15243 4463
rect 15282 4429 15316 4463
rect 15355 4429 15389 4463
rect 15428 4429 15462 4463
rect 15501 4429 15535 4463
rect 15574 4429 15608 4463
rect 15646 4429 15680 4463
rect 15718 4429 15752 4463
rect 15790 4429 15824 4463
rect 15862 4429 15896 4463
rect 15934 4429 15968 4463
rect 16006 4429 16040 4463
rect 16078 4429 16112 4463
rect 16150 4429 16184 4463
rect 16222 4429 16256 4463
rect 16294 4429 16328 4463
rect 16650 4437 16683 4438
rect 16683 4437 16684 4438
rect 16650 4404 16684 4437
rect 13356 4332 13390 4366
rect 13439 4333 13470 4366
rect 13470 4333 13473 4366
rect 13512 4333 13539 4366
rect 13539 4333 13546 4366
rect 13585 4333 13608 4366
rect 13608 4333 13619 4366
rect 13658 4333 13677 4366
rect 13677 4333 13692 4366
rect 13731 4333 13746 4366
rect 13746 4333 13765 4366
rect 13804 4333 13815 4366
rect 13815 4333 13838 4366
rect 13877 4333 13884 4366
rect 13884 4333 13911 4366
rect 13950 4333 13953 4366
rect 13953 4333 13984 4366
rect 13439 4332 13473 4333
rect 13512 4332 13546 4333
rect 13585 4332 13619 4333
rect 13658 4332 13692 4333
rect 13731 4332 13765 4333
rect 13804 4332 13838 4333
rect 13877 4332 13911 4333
rect 13950 4332 13984 4333
rect 14023 4332 14057 4366
rect 14096 4333 14126 4366
rect 14126 4333 14130 4366
rect 14169 4333 14195 4366
rect 14195 4333 14203 4366
rect 14242 4333 14264 4366
rect 14264 4333 14276 4366
rect 14315 4333 14333 4366
rect 14333 4333 14349 4366
rect 14388 4333 14402 4366
rect 14402 4333 14422 4366
rect 14461 4333 14471 4366
rect 14471 4333 14495 4366
rect 14534 4333 14540 4366
rect 14540 4333 14568 4366
rect 14607 4333 14609 4366
rect 14609 4333 14641 4366
rect 14680 4333 14712 4366
rect 14712 4333 14714 4366
rect 14753 4333 14781 4366
rect 14781 4333 14787 4366
rect 14826 4333 14850 4366
rect 14850 4333 14860 4366
rect 14899 4333 14919 4366
rect 14919 4333 14933 4366
rect 14972 4333 14988 4366
rect 14988 4333 15006 4366
rect 15045 4333 15057 4366
rect 15057 4333 15079 4366
rect 15118 4333 15126 4366
rect 15126 4333 15152 4366
rect 15191 4333 15195 4366
rect 15195 4333 15225 4366
rect 14096 4332 14130 4333
rect 14169 4332 14203 4333
rect 14242 4332 14276 4333
rect 14315 4332 14349 4333
rect 14388 4332 14422 4333
rect 14461 4332 14495 4333
rect 14534 4332 14568 4333
rect 14607 4332 14641 4333
rect 14680 4332 14714 4333
rect 14753 4332 14787 4333
rect 14826 4332 14860 4333
rect 14899 4332 14933 4333
rect 14972 4332 15006 4333
rect 15045 4332 15079 4333
rect 15118 4332 15152 4333
rect 15191 4332 15225 4333
rect 15264 4332 15298 4366
rect 15337 4333 15368 4366
rect 15368 4333 15371 4366
rect 15410 4333 15437 4366
rect 15437 4333 15444 4366
rect 15483 4333 15506 4366
rect 15506 4333 15517 4366
rect 15556 4333 15575 4366
rect 15575 4333 15590 4366
rect 15629 4333 15644 4366
rect 15644 4333 15663 4366
rect 15702 4333 15713 4366
rect 15713 4333 15736 4366
rect 15775 4333 15782 4366
rect 15782 4333 15809 4366
rect 15848 4333 15851 4366
rect 15851 4333 15882 4366
rect 15921 4333 15954 4366
rect 15954 4333 15955 4366
rect 15994 4333 16023 4366
rect 16023 4333 16028 4366
rect 16067 4333 16092 4366
rect 16092 4333 16101 4366
rect 16140 4333 16161 4366
rect 16161 4333 16174 4366
rect 16213 4333 16230 4366
rect 16230 4333 16247 4366
rect 16286 4333 16299 4366
rect 16299 4333 16320 4366
rect 16359 4333 16369 4366
rect 16369 4333 16393 4366
rect 16432 4333 16439 4366
rect 16439 4333 16466 4366
rect 16505 4333 16509 4366
rect 16509 4333 16539 4366
rect 16578 4333 16579 4366
rect 16579 4333 16612 4366
rect 15337 4332 15371 4333
rect 15410 4332 15444 4333
rect 15483 4332 15517 4333
rect 15556 4332 15590 4333
rect 15629 4332 15663 4333
rect 15702 4332 15736 4333
rect 15775 4332 15809 4333
rect 15848 4332 15882 4333
rect 15921 4332 15955 4333
rect 15994 4332 16028 4333
rect 16067 4332 16101 4333
rect 16140 4332 16174 4333
rect 16213 4332 16247 4333
rect 16286 4332 16320 4333
rect 16359 4332 16393 4333
rect 16432 4332 16466 4333
rect 16505 4332 16539 4333
rect 16578 4332 16612 4333
rect 16837 6384 16871 6418
rect 16951 6384 16985 6418
rect 16837 6312 16871 6346
rect 16951 6312 16985 6346
rect 16837 6240 16871 6274
rect 16951 6240 16985 6274
rect 16837 6168 16871 6202
rect 16951 6168 16985 6202
rect 16837 6096 16871 6130
rect 16951 6096 16985 6130
rect 16837 6024 16871 6058
rect 16951 6024 16985 6058
rect 16837 5952 16871 5986
rect 16951 5952 16985 5986
rect 16837 5880 16871 5914
rect 16951 5880 16985 5914
rect 16837 5808 16871 5842
rect 16951 5808 16985 5842
rect 16837 5736 16871 5770
rect 16951 5736 16985 5770
rect 16837 5664 16871 5698
rect 16951 5664 16985 5698
rect 16837 5592 16871 5626
rect 16951 5592 16985 5626
rect 16837 5520 16871 5554
rect 16951 5520 16985 5554
rect 16837 5448 16871 5482
rect 16951 5448 16985 5482
rect 16837 5376 16871 5410
rect 16951 5376 16985 5410
rect 16837 5304 16871 5338
rect 16951 5304 16985 5338
rect 16837 5232 16871 5266
rect 16951 5232 16985 5266
rect 16837 5160 16871 5194
rect 16951 5160 16985 5194
rect 16837 5088 16871 5122
rect 16951 5088 16985 5122
rect 16837 5016 16871 5050
rect 16951 5016 16985 5050
rect 16837 4944 16871 4978
rect 16951 4944 16985 4978
rect 16837 4872 16871 4906
rect 16951 4872 16985 4906
rect 16837 4800 16871 4834
rect 16951 4800 16985 4834
rect 16837 4728 16871 4762
rect 16951 4728 16985 4762
rect 16837 4656 16871 4690
rect 16951 4656 16985 4690
rect 16837 4584 16871 4618
rect 16951 4584 16985 4618
rect 16837 4512 16871 4546
rect 16951 4512 16985 4546
rect 16837 4440 16871 4474
rect 16951 4440 16985 4474
rect 16837 4368 16871 4402
rect 16951 4368 16985 4402
rect 13032 4296 13066 4330
rect 13146 4296 13180 4330
rect 13032 4223 13066 4257
rect 13146 4223 13180 4257
rect 16837 4296 16871 4330
rect 16951 4296 16985 4330
rect 16837 4223 16871 4257
rect 16951 4223 16985 4257
rect 13038 4145 13072 4168
rect 13038 4134 13065 4145
rect 13065 4134 13072 4145
rect 13111 4134 13145 4168
rect 13184 4134 13218 4168
rect 13257 4134 13291 4168
rect 13330 4134 13364 4168
rect 13403 4134 13437 4168
rect 13476 4134 13510 4168
rect 13549 4134 13583 4168
rect 13622 4134 13656 4168
rect 13695 4134 13729 4168
rect 13768 4134 13802 4168
rect 13841 4134 13875 4168
rect 13914 4134 13948 4168
rect 13987 4134 14021 4168
rect 14060 4134 14094 4168
rect 14133 4134 14167 4168
rect 14206 4134 14240 4168
rect 14279 4134 14313 4168
rect 14352 4134 14386 4168
rect 14425 4134 14459 4168
rect 14497 4134 14531 4168
rect 14569 4134 14603 4168
rect 14641 4134 14675 4168
rect 14713 4134 14747 4168
rect 14785 4134 14819 4168
rect 14857 4134 14891 4168
rect 14929 4134 14963 4168
rect 15001 4134 15035 4168
rect 15073 4134 15107 4168
rect 15145 4134 15179 4168
rect 15217 4134 15251 4168
rect 15289 4134 15323 4168
rect 15361 4134 15395 4168
rect 15433 4134 15467 4168
rect 15505 4134 15539 4168
rect 15577 4134 15611 4168
rect 15649 4134 15683 4168
rect 15721 4134 15755 4168
rect 15793 4134 15827 4168
rect 15865 4134 15899 4168
rect 15937 4134 15971 4168
rect 16009 4134 16043 4168
rect 16081 4134 16115 4168
rect 16153 4134 16187 4168
rect 16225 4134 16259 4168
rect 16297 4134 16331 4168
rect 16369 4134 16403 4168
rect 16441 4134 16475 4168
rect 16513 4134 16547 4168
rect 16585 4134 16619 4168
rect 16657 4134 16691 4168
rect 16729 4134 16763 4168
rect 16801 4134 16835 4168
rect 16873 4134 16907 4168
rect 16945 4145 16979 4168
rect 16945 4134 16961 4145
rect 16961 4134 16979 4145
rect 13038 4020 13072 4054
rect 13111 4043 13126 4054
rect 13126 4043 13145 4054
rect 13111 4020 13145 4043
rect 13184 4020 13218 4054
rect 13257 4020 13291 4054
rect 13330 4020 13364 4054
rect 13403 4020 13437 4054
rect 13476 4020 13510 4054
rect 13549 4020 13583 4054
rect 13622 4020 13656 4054
rect 13695 4020 13729 4054
rect 13768 4020 13802 4054
rect 13841 4020 13875 4054
rect 13914 4020 13948 4054
rect 13987 4020 14021 4054
rect 14060 4020 14094 4054
rect 14133 4020 14167 4054
rect 14206 4020 14240 4054
rect 14279 4020 14313 4054
rect 14352 4020 14386 4054
rect 14425 4020 14459 4054
rect 14497 4020 14531 4054
rect 14569 4020 14603 4054
rect 14641 4020 14675 4054
rect 14713 4020 14747 4054
rect 14785 4020 14819 4054
rect 14857 4020 14891 4054
rect 14929 4020 14963 4054
rect 15001 4020 15035 4054
rect 15073 4020 15107 4054
rect 15145 4020 15179 4054
rect 15217 4020 15251 4054
rect 15289 4020 15323 4054
rect 15361 4020 15395 4054
rect 15433 4020 15467 4054
rect 15505 4020 15539 4054
rect 15577 4020 15611 4054
rect 15649 4020 15683 4054
rect 15721 4020 15755 4054
rect 15793 4020 15827 4054
rect 15865 4020 15899 4054
rect 15937 4020 15971 4054
rect 16009 4020 16043 4054
rect 16081 4020 16115 4054
rect 16153 4020 16187 4054
rect 16225 4020 16259 4054
rect 16297 4020 16331 4054
rect 16369 4020 16403 4054
rect 16441 4020 16475 4054
rect 16513 4020 16547 4054
rect 16585 4020 16619 4054
rect 16657 4020 16691 4054
rect 16729 4020 16763 4054
rect 16801 4020 16835 4054
rect 16873 4043 16900 4054
rect 16900 4043 16907 4054
rect 16873 4020 16907 4043
rect 16945 4020 16979 4054
rect 17218 6643 17252 6677
rect 17344 6643 17378 6677
rect 17218 6570 17252 6604
rect 17344 6570 17378 6604
rect 17218 6497 17252 6531
rect 17344 6497 17378 6531
rect 17218 6424 17252 6458
rect 17344 6424 17378 6458
rect 17218 6351 17252 6385
rect 17344 6351 17378 6385
rect 17218 6278 17252 6312
rect 17344 6278 17378 6312
rect 17218 6205 17252 6239
rect 17344 6205 17378 6239
rect 17218 6132 17252 6166
rect 17344 6132 17378 6166
rect 17218 6059 17252 6093
rect 17344 6059 17378 6093
rect 17218 5986 17252 6020
rect 17344 5986 17378 6020
rect 17218 5913 17252 5947
rect 17344 5913 17378 5947
rect 17218 5840 17252 5874
rect 17344 5840 17378 5874
rect 17218 5767 17252 5801
rect 17344 5767 17378 5801
rect 17218 5694 17252 5728
rect 17344 5694 17378 5728
rect 17218 5621 17252 5655
rect 17344 5621 17378 5655
rect 17218 5548 17252 5582
rect 17344 5548 17378 5582
rect 17218 5475 17252 5509
rect 17344 5475 17378 5509
rect 17218 5402 17252 5436
rect 17344 5402 17378 5436
rect 17218 5329 17252 5363
rect 17344 5329 17378 5363
rect 17218 5256 17252 5290
rect 17344 5256 17378 5290
rect 17218 5183 17252 5217
rect 17344 5183 17378 5217
rect 17218 5110 17252 5144
rect 17344 5110 17378 5144
rect 17218 5037 17252 5071
rect 17344 5037 17378 5071
rect 17218 4964 17252 4998
rect 17344 4964 17378 4998
rect 17218 4891 17252 4925
rect 17344 4891 17378 4925
rect 17218 4818 17252 4852
rect 17344 4818 17378 4852
rect 17218 4745 17252 4779
rect 17344 4745 17378 4779
rect 17218 4672 17252 4706
rect 17344 4672 17378 4706
rect 17218 4599 17252 4633
rect 17344 4599 17378 4633
rect 17218 4526 17252 4560
rect 17344 4526 17378 4560
rect 17218 4453 17252 4487
rect 17344 4453 17378 4487
rect 17218 4380 17252 4414
rect 17344 4380 17378 4414
rect 17218 4307 17252 4341
rect 17344 4307 17378 4341
rect 17218 4234 17252 4268
rect 17344 4234 17378 4268
rect 17218 4160 17252 4194
rect 17344 4160 17378 4194
rect 17218 4086 17252 4120
rect 17344 4086 17378 4120
rect 12634 3984 12668 4018
rect 12760 3984 12794 4018
rect 12634 3910 12668 3944
rect 12760 3910 12794 3944
rect 12634 3860 12668 3870
rect 12760 3860 12794 3870
rect 12634 3836 12668 3860
rect 12760 3836 12794 3860
rect 17218 4012 17252 4046
rect 17344 4012 17378 4046
rect 17218 3938 17252 3972
rect 17344 3938 17378 3972
rect 17218 3864 17252 3898
rect 17344 3864 17378 3898
rect 4235 3770 4269 3778
rect 4235 3709 4269 3727
rect 4235 3693 4269 3709
rect 2974 3648 3008 3682
rect 3046 3648 3080 3682
rect 3118 3648 3152 3682
rect 3910 3648 3944 3682
rect 3983 3648 4017 3682
rect 4055 3648 4089 3682
rect 4127 3648 4161 3682
rect 1276 3594 1310 3628
rect 1348 3594 1382 3628
rect 1588 3594 1622 3628
rect 1660 3594 1694 3628
rect 1900 3594 1934 3628
rect 1972 3594 2006 3628
rect 2212 3594 2246 3628
rect 2284 3594 2318 3628
rect 3198 3580 3232 3614
rect 1156 3506 1190 3540
rect 1156 3434 1190 3468
rect 1156 3362 1190 3396
rect 1468 3506 1502 3540
rect 1468 3434 1502 3468
rect 1468 3362 1502 3396
rect 1780 3506 1814 3540
rect 1780 3434 1814 3468
rect 1780 3362 1814 3396
rect 2092 3506 2126 3540
rect 2092 3434 2126 3468
rect 2092 3362 2126 3396
rect 1156 3053 1190 3087
rect 1156 2981 1190 3015
rect 1156 2909 1190 2943
rect 1156 2837 1190 2871
rect 1156 2765 1190 2799
rect 1156 2693 1190 2727
rect 1468 3053 1502 3087
rect 1468 2981 1502 3015
rect 1468 2909 1502 2943
rect 1468 2837 1502 2871
rect 1468 2765 1502 2799
rect 1468 2693 1502 2727
rect 1780 3053 1814 3087
rect 1780 2981 1814 3015
rect 1780 2909 1814 2943
rect 1780 2837 1814 2871
rect 1780 2765 1814 2799
rect 1780 2693 1814 2727
rect 2092 3053 2126 3087
rect 2092 2981 2126 3015
rect 3198 3532 3205 3542
rect 3205 3532 3232 3542
rect 3198 3508 3232 3532
rect 2491 3168 2597 3346
rect 2092 2909 2126 2943
rect 2092 2837 2126 2871
rect 2092 2765 2126 2799
rect 2092 2693 2126 2727
rect 186 216 220 250
rect 186 144 220 178
rect 186 72 220 106
rect 618 216 652 250
rect 618 144 652 178
rect 618 72 652 106
<< metal1 >>
rect 2312 8153 2358 8165
rect 2312 8119 2318 8153
rect 2352 8119 2358 8153
tri 2287 8087 2312 8112 se
rect 2312 8087 2358 8119
rect 2287 8081 2358 8087
rect 2287 8047 2318 8081
rect 2352 8047 2358 8081
rect 2287 8035 2358 8047
rect 43 7995 287 8007
rect 43 7961 49 7995
rect 83 7961 287 7995
rect 43 7955 287 7961
rect 43 7923 89 7955
tri 89 7930 114 7955 nw
rect 43 7889 49 7923
rect 83 7889 89 7923
rect 43 7877 89 7889
rect 2389 7895 2435 7907
tri 2376 7861 2389 7874 se
rect 2389 7861 2395 7895
rect 2429 7861 2435 7895
tri 2364 7849 2376 7861 se
rect 2376 7849 2435 7861
rect 2287 7823 2435 7849
rect 2287 7797 2395 7823
tri 2369 7789 2377 7797 ne
rect 2377 7789 2395 7797
rect 2429 7789 2435 7823
tri 2377 7777 2389 7789 ne
rect 2389 7777 2435 7789
rect 140 7567 169 7769
rect 140 7539 345 7567
rect 2210 7545 2269 7769
rect 3192 7766 3238 7778
tri 2287 7732 2304 7749 sw
rect 3192 7732 3198 7766
rect 3232 7732 3238 7766
rect 2287 7694 2304 7732
tri 2304 7694 2342 7732 sw
rect 3192 7694 3238 7732
rect 2287 7660 2342 7694
tri 2342 7660 2376 7694 sw
rect 3192 7660 3198 7694
rect 3232 7660 3238 7694
rect 2287 7648 2376 7660
tri 2376 7648 2388 7660 sw
rect 2287 7646 2388 7648
tri 2388 7646 2390 7648 sw
rect 2287 7640 2390 7646
tri 2390 7640 2396 7646 sw
rect 2287 7638 2396 7640
tri 2396 7638 2398 7640 sw
rect 2287 7613 2398 7638
tri 2398 7613 2423 7638 sw
tri 3167 7613 3192 7638 se
rect 3192 7613 3238 7660
tri 4395 7658 4420 7683 se
rect 2287 7607 2423 7613
tri 2423 7607 2429 7613 sw
rect 2923 7607 3238 7613
rect 2287 7594 2429 7607
tri 2429 7594 2442 7607 sw
rect 140 7493 169 7539
rect 2210 7533 2281 7545
rect 2210 7499 2241 7533
rect 2275 7499 2281 7533
rect 2210 7493 2281 7499
rect 2287 7493 2442 7594
tri 2157 7461 2189 7493 ne
rect 2189 7461 2442 7493
tri 2189 7427 2223 7461 ne
rect 2223 7427 2241 7461
rect 2275 7427 2442 7461
tri 2223 7415 2235 7427 ne
rect 2235 7415 2442 7427
tri 2235 7335 2315 7415 ne
tri 142 7317 148 7323 se
rect -132 7271 140 7317
rect 148 7271 154 7323
rect 206 7271 218 7323
rect 270 7271 282 7323
rect 334 7271 346 7323
rect 398 7271 404 7323
tri 404 7317 410 7323 sw
rect -133 7243 345 7271
tri 345 7247 369 7271 nw
rect -104 7041 140 7243
rect -104 7035 -4 7041
tri -4 7035 2 7041 nw
rect -104 7001 -38 7035
tri -38 7001 -4 7035 nw
rect -104 6999 -40 7001
tri -40 6999 -38 7001 nw
rect -104 6998 -41 6999
tri -41 6998 -40 6999 nw
rect 337 6998 465 6999
rect -104 6987 -52 6998
tri -52 6987 -41 6998 nw
rect -104 6953 -86 6987
tri -86 6953 -52 6987 nw
rect -104 6946 -93 6953
tri -93 6946 -86 6953 nw
rect 337 6946 343 6998
rect 395 6946 407 6998
rect 459 6946 465 6998
rect -104 6941 -98 6946
tri -98 6941 -93 6946 nw
rect 337 6941 465 6946
tri -104 6935 -98 6941 nw
tri -104 6836 -100 6840 sw
rect -104 6823 -100 6836
tri -100 6823 -87 6836 sw
rect -104 6797 -87 6823
tri -87 6797 -61 6823 sw
rect -104 6782 -61 6797
tri -61 6782 -46 6797 sw
rect -104 6763 -46 6782
tri -46 6763 -27 6782 sw
rect -104 6750 -27 6763
tri -27 6750 -14 6763 sw
rect -104 6739 -14 6750
tri -14 6739 -3 6750 sw
rect -104 6733 -3 6739
tri -3 6733 3 6739 sw
rect -104 6709 3 6733
tri 3 6709 27 6733 sw
rect -104 6703 27 6709
rect -104 6651 -40 6703
rect 12 6699 27 6703
tri 27 6699 37 6709 sw
rect 12 6651 73 6699
rect -104 6639 73 6651
rect -104 6587 -40 6639
rect 12 6587 73 6639
rect -104 6575 73 6587
rect -104 6523 -40 6575
rect 12 6523 73 6575
rect -104 6511 73 6523
rect -104 6459 -40 6511
rect 12 6497 73 6511
rect 12 6469 2287 6497
rect 12 6459 221 6469
rect -104 6447 221 6459
rect -104 6395 -40 6447
rect 12 6417 221 6447
rect 12 6406 210 6417
tri 210 6406 221 6417 nw
rect 12 6395 176 6406
rect -104 6383 176 6395
rect -104 6331 -40 6383
rect 12 6372 176 6383
tri 176 6372 210 6406 nw
rect 12 6359 163 6372
tri 163 6359 176 6372 nw
rect 12 6331 129 6359
rect -104 6325 129 6331
tri 129 6325 163 6359 nw
rect -104 6319 117 6325
rect -104 6267 -40 6319
rect 12 6313 117 6319
tri 117 6313 129 6325 nw
rect 12 6312 116 6313
tri 116 6312 117 6313 nw
tri 2314 6312 2315 6313 se
rect 2315 6312 2442 7415
rect 2923 7573 3046 7607
rect 3080 7573 3118 7607
rect 3152 7573 3238 7607
rect 2831 7096 2895 7102
rect 2831 7044 2837 7096
rect 2889 7044 2895 7096
rect 2831 7032 2895 7044
rect 2831 6980 2837 7032
rect 2889 6980 2895 7032
rect 2831 6968 2895 6980
rect 2831 6916 2837 6968
rect 2889 6916 2895 6968
rect 2831 6904 2895 6916
rect 2831 6852 2837 6904
rect 2889 6852 2895 6904
rect 2831 6840 2895 6852
rect 2831 6788 2837 6840
rect 2889 6788 2895 6840
rect 2831 6782 2895 6788
rect 12 6286 90 6312
tri 90 6286 116 6312 nw
tri 2288 6286 2314 6312 se
rect 2314 6286 2442 6312
rect 12 6267 73 6286
tri 73 6269 90 6286 nw
tri 2271 6269 2288 6286 se
rect 2288 6269 2442 6286
rect -104 5814 73 6267
tri 2263 6261 2271 6269 se
rect 2271 6261 2442 6269
tri 2254 6252 2263 6261 se
rect 2263 6252 2442 6261
tri 2249 6247 2254 6252 se
rect 2254 6247 2442 6252
rect 2287 6168 2442 6247
rect 2831 6733 2895 6739
rect 2831 6699 2849 6733
rect 2883 6699 2895 6733
rect 2831 6661 2895 6699
rect 2831 6627 2849 6661
rect 2883 6627 2895 6661
rect 2831 6589 2895 6627
rect 2831 6555 2849 6589
rect 2883 6555 2895 6589
rect 2831 6478 2895 6555
rect 2831 6444 2849 6478
rect 2883 6444 2895 6478
rect 2831 6406 2895 6444
rect 2831 6372 2849 6406
rect 2883 6372 2895 6406
tri 2442 6168 2451 6177 sw
rect 2287 6140 2451 6168
tri 2451 6140 2479 6168 sw
rect 2287 6106 2479 6140
tri 2479 6106 2513 6140 sw
rect 2287 6096 2513 6106
tri 2513 6096 2523 6106 sw
rect 2287 6067 2523 6096
tri 2523 6067 2552 6096 sw
rect 2287 6033 2552 6067
tri 2552 6033 2586 6067 sw
rect 2287 6024 2586 6033
tri 2586 6024 2595 6033 sw
rect 2287 6014 2595 6024
tri 2595 6014 2605 6024 sw
rect 2287 5971 2605 6014
tri 2339 5960 2350 5971 ne
rect 2350 5960 2605 5971
tri 2350 5952 2358 5960 ne
rect 2358 5952 2605 5960
tri 2358 5921 2389 5952 ne
rect 2389 5921 2605 5952
tri 2389 5887 2423 5921 ne
rect 2423 5887 2605 5921
tri 2423 5880 2430 5887 ne
rect 2430 5880 2605 5887
tri 2430 5848 2462 5880 ne
rect 2462 5848 2605 5880
tri 2462 5833 2477 5848 ne
tri 73 5814 92 5833 sw
rect -104 5808 92 5814
tri 92 5808 98 5814 sw
rect -104 5775 98 5808
tri 98 5775 131 5808 sw
rect -104 5749 131 5775
tri 131 5749 157 5775 sw
rect -104 5743 515 5749
rect -104 5709 325 5743
rect 359 5709 397 5743
rect 431 5709 469 5743
rect 503 5709 515 5743
rect -104 5703 515 5709
rect -104 5702 156 5703
tri 156 5702 157 5703 nw
rect -104 5668 122 5702
tri 122 5668 156 5702 nw
rect -104 5664 118 5668
tri 118 5664 122 5668 nw
rect -104 5662 116 5664
tri 116 5662 118 5664 nw
rect -104 5629 83 5662
tri 83 5629 116 5662 nw
rect -104 4203 73 5629
tri 73 5619 83 5629 nw
tri 2460 5340 2477 5357 se
rect 2477 5340 2605 5848
tri 2458 5338 2460 5340 se
rect 2460 5338 2605 5340
tri 2457 5337 2458 5338 se
rect 2458 5337 2605 5338
tri 2452 5332 2457 5337 se
rect 2457 5332 2605 5337
rect 129 5320 2605 5332
rect 129 5286 135 5320
rect 169 5286 447 5320
rect 481 5286 759 5320
rect 793 5286 1071 5320
rect 1105 5286 1383 5320
rect 1417 5286 1695 5320
rect 1729 5286 2007 5320
rect 2041 5286 2237 5320
rect 2271 5286 2605 5320
rect 129 5248 2605 5286
rect 129 5214 135 5248
rect 169 5214 447 5248
rect 481 5214 759 5248
rect 793 5214 1071 5248
rect 1105 5214 1383 5248
rect 1417 5214 1695 5248
rect 1729 5214 2007 5248
rect 2041 5214 2237 5248
rect 2271 5214 2605 5248
rect 129 5176 2605 5214
rect 129 5142 135 5176
rect 169 5142 447 5176
rect 481 5142 759 5176
rect 793 5142 1071 5176
rect 1105 5142 1383 5176
rect 1417 5142 1695 5176
rect 1729 5142 2007 5176
rect 2041 5142 2237 5176
rect 2271 5142 2605 5176
rect 129 5130 2605 5142
tri 2452 5124 2458 5130 ne
rect 2458 5124 2605 5130
tri 2458 5123 2459 5124 ne
rect 2459 5123 2605 5124
tri 2459 5122 2460 5123 ne
rect 2460 5122 2605 5123
tri 2460 5118 2464 5122 ne
rect 2464 5118 2605 5122
tri 2464 5108 2474 5118 ne
rect 2474 5108 2605 5118
tri 2474 5105 2477 5108 ne
rect 207 5089 253 5101
rect 207 5055 213 5089
rect 247 5055 253 5089
rect 207 5017 253 5055
rect 597 5089 643 5101
rect 597 5055 603 5089
rect 637 5055 643 5089
tri 253 5017 260 5024 sw
tri 590 5017 597 5024 se
rect 597 5017 643 5055
rect 207 4983 213 5017
rect 247 4999 260 5017
tri 260 4999 278 5017 sw
tri 572 4999 590 5017 se
rect 590 4999 603 5017
rect 247 4983 603 4999
rect 637 4983 643 5017
rect 207 4971 643 4983
rect 909 5089 955 5101
rect 909 5055 915 5089
rect 949 5055 955 5089
rect 909 5017 955 5055
rect 1299 5089 2129 5101
rect 1299 5055 1305 5089
rect 1339 5073 2089 5089
rect 1339 5055 1352 5073
tri 1352 5055 1370 5073 nw
tri 2058 5055 2076 5073 ne
rect 2076 5055 2089 5073
rect 2123 5055 2129 5089
rect 1299 5052 1349 5055
tri 1349 5052 1352 5055 nw
tri 2076 5052 2079 5055 ne
rect 2079 5052 2129 5055
rect 1299 5050 1347 5052
tri 1347 5050 1349 5052 nw
tri 2079 5050 2081 5052 ne
rect 2081 5050 2129 5052
tri 955 5017 962 5024 sw
tri 1292 5017 1299 5024 se
rect 1299 5017 1345 5050
tri 1345 5048 1347 5050 nw
tri 2081 5048 2083 5050 ne
rect 909 4983 915 5017
rect 949 4999 962 5017
tri 962 4999 980 5017 sw
tri 1274 4999 1292 5017 se
rect 1292 4999 1305 5017
rect 949 4983 1305 4999
rect 1339 4983 1345 5017
rect 909 4971 1345 4983
rect 1762 5033 1826 5045
rect 1762 4979 1768 5033
rect 1802 5031 1826 5033
rect 1820 4979 1826 5031
tri 572 4968 575 4971 ne
rect 575 4968 643 4971
tri 575 4961 582 4968 ne
rect 582 4961 643 4968
tri 643 4961 650 4968 sw
tri 1755 4961 1762 4968 se
rect 1762 4967 1826 4979
rect 2083 5017 2129 5050
rect 2083 4983 2089 5017
rect 2123 4983 2129 5017
rect 2083 4971 2129 4983
rect 1762 4961 1768 4967
tri 582 4946 597 4961 ne
rect 597 4943 650 4961
tri 650 4943 668 4961 sw
tri 1737 4943 1755 4961 se
rect 1755 4943 1768 4961
rect 597 4915 1768 4943
rect 1820 4915 1826 4967
rect 282 4881 334 4887
rect 282 4817 334 4829
rect 282 4756 334 4765
rect 1221 4881 1273 4887
rect 1508 4875 1851 4887
rect 1508 4859 1539 4875
tri 1508 4841 1526 4859 ne
rect 1526 4841 1539 4859
rect 1573 4859 1851 4875
rect 1573 4841 1586 4859
tri 1586 4841 1604 4859 nw
tri 1820 4841 1838 4859 ne
rect 1838 4841 1851 4859
tri 1526 4836 1531 4841 ne
rect 1531 4836 1581 4841
tri 1581 4836 1586 4841 nw
tri 1838 4836 1843 4841 ne
rect 1843 4836 1851 4841
tri 1531 4834 1533 4836 ne
rect 1221 4817 1273 4829
rect 1221 4757 1273 4765
rect 1533 4803 1579 4836
tri 1579 4834 1581 4836 nw
tri 1843 4834 1845 4836 ne
rect 1845 4835 1851 4836
rect 1903 4835 1909 4887
rect 1533 4769 1539 4803
rect 1573 4769 1579 4803
rect 1533 4757 1579 4769
rect 1845 4823 1909 4835
rect 1845 4769 1851 4823
rect 1903 4771 1909 4823
rect 1885 4769 1909 4771
rect 1845 4757 1909 4769
tri 312 4701 334 4723 se
rect 334 4716 489 4723
tri 489 4716 496 4723 sw
rect 334 4701 496 4716
tri 496 4701 511 4716 sw
tri 1247 4701 1262 4716 se
rect 1262 4701 1525 4716
tri 1525 4701 1540 4716 sw
tri 301 4690 312 4701 se
rect 312 4690 511 4701
tri 511 4690 522 4701 sw
tri 1236 4690 1247 4701 se
rect 1247 4690 1540 4701
tri 1540 4690 1551 4701 sw
rect 140 4686 2367 4690
rect 140 4678 2283 4686
rect 140 4644 146 4678
rect 180 4644 218 4678
rect 252 4654 1115 4678
rect 252 4644 345 4654
tri 345 4644 355 4654 nw
tri 460 4644 470 4654 ne
rect 470 4644 1115 4654
rect 1149 4644 1187 4678
rect 1221 4655 2283 4678
rect 1221 4646 1271 4655
tri 1271 4646 1280 4655 nw
tri 1488 4646 1497 4655 ne
rect 1497 4646 2283 4655
rect 1221 4644 1259 4646
rect 140 4632 333 4644
tri 333 4632 345 4644 nw
tri 470 4632 482 4644 ne
rect 482 4634 1259 4644
tri 1259 4634 1271 4646 nw
tri 1497 4634 1509 4646 ne
rect 1509 4634 2283 4646
rect 2335 4634 2347 4686
rect 2399 4634 2405 4686
rect 482 4632 1257 4634
tri 1257 4632 1259 4634 nw
tri 1509 4632 1511 4634 ne
rect 1511 4632 2367 4634
rect 369 4614 427 4624
tri 427 4614 437 4624 sw
rect 369 4610 437 4614
tri 437 4610 441 4614 sw
rect 369 4608 441 4610
rect 369 4574 381 4608
rect 415 4604 441 4608
tri 441 4604 447 4610 sw
tri 1306 4604 1312 4610 se
rect 1312 4604 1318 4610
rect 415 4598 1318 4604
rect 415 4574 904 4598
rect 369 4564 904 4574
rect 938 4564 976 4598
rect 1010 4576 1318 4598
rect 1010 4564 1028 4576
tri 1028 4564 1040 4576 nw
tri 1294 4564 1306 4576 ne
rect 1306 4564 1318 4576
rect 369 4558 1022 4564
tri 1022 4558 1028 4564 nw
tri 1306 4558 1312 4564 ne
rect 1312 4558 1318 4564
rect 1370 4558 1382 4610
rect 1434 4558 1442 4610
rect 1616 4598 2281 4604
rect 1616 4564 1628 4598
rect 1662 4564 1700 4598
rect 1734 4564 2163 4598
rect 2197 4564 2235 4598
rect 2269 4564 2281 4598
rect 1616 4558 2281 4564
rect 2309 4592 2355 4604
rect 2309 4558 2315 4592
rect 2349 4558 2355 4592
rect 369 4557 460 4558
tri 460 4557 461 4558 nw
rect 369 4552 455 4557
tri 455 4552 460 4557 nw
rect 369 4548 451 4552
tri 451 4548 455 4552 nw
rect 369 4542 445 4548
tri 445 4542 451 4548 nw
rect 1130 4542 1260 4548
tri 1260 4542 1266 4548 sw
rect 369 4536 427 4542
rect 369 4502 381 4536
rect 415 4502 427 4536
tri 427 4524 445 4542 nw
rect 1130 4508 1142 4542
rect 1176 4508 1214 4542
rect 1248 4530 1266 4542
tri 1266 4530 1278 4542 sw
tri 2297 4530 2309 4542 se
rect 2309 4530 2355 4558
rect 1248 4520 2222 4530
tri 2222 4520 2232 4530 sw
tri 2287 4520 2297 4530 se
rect 2297 4520 2355 4530
rect 1248 4517 2232 4520
tri 2232 4517 2235 4520 sw
tri 2284 4517 2287 4520 se
rect 2287 4517 2315 4520
rect 1248 4508 2233 4517
rect 1130 4502 2233 4508
rect 369 4496 427 4502
tri 2190 4496 2196 4502 ne
rect 2196 4496 2233 4502
tri 2196 4486 2206 4496 ne
rect 2206 4486 2233 4496
tri 2206 4477 2215 4486 ne
rect 2215 4477 2233 4486
tri 2215 4472 2220 4477 ne
rect 2220 4472 2233 4477
tri 277 4468 281 4472 sw
tri 2220 4468 2224 4472 ne
rect 2224 4468 2233 4472
rect 149 4462 1517 4468
tri 2224 4465 2227 4468 ne
rect 2227 4465 2233 4468
rect 2285 4465 2297 4517
rect 2349 4465 2355 4520
rect 149 4428 1471 4462
rect 1505 4428 1517 4462
rect 149 4422 1517 4428
tri 277 4420 279 4422 nw
rect 1032 4369 2072 4375
rect 1032 4335 1044 4369
rect 1078 4347 1832 4369
rect 1078 4335 1103 4347
tri 1103 4335 1115 4347 nw
tri 1795 4335 1807 4347 ne
rect 1807 4335 1832 4347
rect 1866 4347 2026 4369
rect 1866 4335 1891 4347
tri 1891 4335 1903 4347 nw
tri 1989 4335 2001 4347 ne
rect 2001 4335 2026 4347
rect 2060 4335 2072 4369
rect 1032 4327 1095 4335
tri 1095 4327 1103 4335 nw
tri 1807 4327 1815 4335 ne
rect 1815 4327 1883 4335
tri 1883 4327 1891 4335 nw
tri 2001 4327 2009 4335 ne
rect 2009 4327 2072 4335
rect 468 4309 514 4321
rect 468 4275 474 4309
rect 508 4275 514 4309
rect 468 4237 514 4275
rect 1032 4297 1090 4327
tri 1090 4322 1095 4327 nw
tri 1815 4322 1820 4327 ne
rect 1032 4263 1044 4297
rect 1078 4263 1090 4297
rect 1032 4257 1090 4263
rect 1820 4297 1878 4327
tri 1878 4322 1883 4327 nw
tri 2009 4322 2014 4327 ne
rect 1820 4263 1832 4297
rect 1866 4263 1878 4297
rect 1820 4257 1878 4263
rect 1914 4309 1972 4315
rect 1914 4275 1926 4309
rect 1960 4275 1972 4309
tri 861 4244 869 4252 se
rect 869 4244 977 4252
tri 977 4244 985 4252 sw
tri 514 4237 521 4244 sw
tri 854 4237 861 4244 se
rect 861 4237 985 4244
tri 985 4237 992 4244 sw
tri 1907 4237 1914 4244 se
rect 1914 4237 1972 4275
rect 2014 4297 2072 4327
rect 2477 4355 2605 5108
rect 2831 5031 2895 6372
rect 2831 4979 2837 5031
rect 2889 4979 2895 5031
rect 2831 4967 2895 4979
rect 2831 4915 2837 4967
rect 2889 4915 2895 4967
rect 2923 6651 3238 7573
rect 3488 7640 3690 7646
rect 3488 7606 3500 7640
rect 3534 7606 3572 7640
rect 3606 7606 3644 7640
rect 3678 7606 3690 7640
rect 3488 7464 3690 7606
tri 3505 7439 3530 7464 ne
rect 3266 7109 3322 7119
rect 3324 7118 3360 7119
rect 3266 7057 3270 7109
rect 3266 7045 3322 7057
rect 3266 6993 3270 7045
rect 3266 6981 3322 6993
rect 3266 6929 3270 6981
rect 3266 6917 3322 6929
rect 3266 6865 3270 6917
rect 3266 6859 3322 6865
rect 3323 6860 3361 7118
rect 3362 7107 3408 7119
rect 3362 7073 3368 7107
rect 3402 7073 3408 7107
rect 3362 7035 3408 7073
rect 3362 7001 3368 7035
rect 3402 7001 3408 7035
rect 3362 6963 3408 7001
rect 3362 6929 3368 6963
rect 3402 6929 3408 6963
rect 3324 6859 3360 6860
rect 3362 6859 3408 6929
rect 3266 6836 3300 6859
tri 3300 6836 3323 6859 nw
rect 3266 6790 3298 6836
tri 3298 6834 3300 6836 nw
tri 3298 6790 3302 6794 sw
rect 3266 6744 3302 6790
rect 3267 6742 3301 6743
rect 2923 6617 2942 6651
rect 2976 6617 3014 6651
rect 3048 6617 3086 6651
rect 3120 6617 3238 6651
rect 2923 6515 3238 6617
rect 3267 6705 3301 6706
rect 3266 6658 3302 6704
tri 3527 6685 3530 6688 se
rect 3530 6685 3690 7464
tri 3505 6663 3527 6685 se
rect 3527 6663 3690 6685
rect 3266 6657 3301 6658
tri 3301 6657 3302 6658 nw
rect 3414 6657 3690 6663
rect 3266 6611 3298 6657
tri 3298 6654 3301 6657 nw
rect 3414 6623 3426 6657
rect 3460 6623 3498 6657
rect 3532 6623 3570 6657
rect 3604 6623 3642 6657
rect 3676 6623 3690 6657
rect 4392 6648 4420 7658
rect 3414 6617 3690 6623
tri 4346 6617 4377 6648 ne
rect 4377 6617 4420 6648
tri 3505 6614 3508 6617 ne
rect 3508 6614 3690 6617
tri 3298 6611 3301 6614 sw
tri 3508 6611 3511 6614 ne
rect 3511 6611 3690 6614
tri 4377 6611 4383 6617 ne
rect 4383 6611 4420 6617
rect 3266 6604 3301 6611
tri 3301 6604 3308 6611 sw
tri 3511 6604 3518 6611 ne
rect 3518 6604 3690 6611
tri 4383 6604 4390 6611 ne
rect 4390 6604 4420 6611
rect 3266 6589 3308 6604
tri 3308 6589 3323 6604 sw
tri 3518 6592 3530 6604 ne
rect 3266 6543 3322 6589
rect 3324 6588 3360 6589
rect 3323 6544 3361 6588
rect 3362 6583 3493 6589
rect 3362 6549 3375 6583
rect 3409 6549 3447 6583
rect 3481 6549 3493 6583
rect 3324 6543 3360 6544
rect 3362 6543 3493 6549
rect 3266 6537 3317 6543
tri 3317 6537 3323 6543 nw
tri 3527 6537 3530 6540 se
rect 3530 6537 3690 6604
tri 4390 6589 4405 6604 ne
rect 4405 6589 4420 6604
tri 4405 6578 4416 6589 ne
rect 4416 6578 4420 6589
tri 4416 6574 4420 6578 ne
rect 12628 7081 17278 7087
rect 12628 7047 12643 7081
rect 12677 7047 12716 7081
rect 12750 7047 12789 7081
rect 12823 7047 12862 7081
rect 12896 7047 12935 7081
rect 12969 7047 13008 7081
rect 13042 7047 13081 7081
rect 13115 7047 13154 7081
rect 13188 7047 13227 7081
rect 13261 7047 13300 7081
rect 13334 7047 13373 7081
rect 13407 7047 13446 7081
rect 13480 7047 13519 7081
rect 13553 7047 13592 7081
rect 13626 7047 13665 7081
rect 13699 7047 13738 7081
rect 13772 7047 13811 7081
rect 13845 7047 13884 7081
rect 13918 7047 13957 7081
rect 13991 7047 14029 7081
rect 14063 7047 14101 7081
rect 14135 7047 14173 7081
rect 14207 7047 14245 7081
rect 14279 7047 14317 7081
rect 14351 7047 14389 7081
rect 14423 7047 14461 7081
rect 14495 7047 14533 7081
rect 14567 7047 14605 7081
rect 14639 7047 14677 7081
rect 14711 7047 14749 7081
rect 14783 7047 14821 7081
rect 14855 7047 14893 7081
rect 14927 7047 14965 7081
rect 14999 7047 15037 7081
rect 15071 7047 15109 7081
rect 15143 7047 15181 7081
rect 15215 7047 15253 7081
rect 15287 7047 15325 7081
rect 15359 7047 15397 7081
rect 15431 7047 15469 7081
rect 15503 7047 15541 7081
rect 15575 7047 15613 7081
rect 15647 7047 15685 7081
rect 15719 7047 15757 7081
rect 15791 7047 15829 7081
rect 15863 7047 15901 7081
rect 15935 7047 15973 7081
rect 16007 7047 16045 7081
rect 16079 7047 16117 7081
rect 16151 7047 16189 7081
rect 16223 7047 16261 7081
rect 16295 7047 16333 7081
rect 16367 7047 16405 7081
rect 16439 7047 16477 7081
rect 16511 7047 16549 7081
rect 16583 7047 16621 7081
rect 16655 7047 16693 7081
rect 16727 7047 16765 7081
rect 16799 7047 16837 7081
rect 16871 7047 16909 7081
rect 16943 7047 16981 7081
rect 17015 7047 17053 7081
rect 17087 7047 17125 7081
rect 17159 7047 17278 7081
rect 12628 6981 17278 7047
tri 17278 6981 17384 7087 sw
rect 12628 6969 17384 6981
rect 12628 6955 17218 6969
rect 12628 6921 12643 6955
rect 12677 6921 12716 6955
rect 12750 6921 12789 6955
rect 12823 6921 12862 6955
rect 12896 6921 12935 6955
rect 12969 6921 13008 6955
rect 13042 6921 13081 6955
rect 13115 6921 13154 6955
rect 13188 6921 13227 6955
rect 13261 6921 13300 6955
rect 13334 6921 13373 6955
rect 13407 6921 13446 6955
rect 13480 6921 13519 6955
rect 13553 6921 13592 6955
rect 13626 6921 13665 6955
rect 13699 6921 13738 6955
rect 13772 6921 13811 6955
rect 13845 6921 13884 6955
rect 13918 6921 13957 6955
rect 13991 6921 14029 6955
rect 14063 6921 14101 6955
rect 14135 6921 14173 6955
rect 14207 6921 14245 6955
rect 14279 6921 14317 6955
rect 14351 6921 14389 6955
rect 14423 6921 14461 6955
rect 14495 6921 14533 6955
rect 14567 6921 14605 6955
rect 14639 6921 14677 6955
rect 14711 6921 14749 6955
rect 14783 6921 14821 6955
rect 14855 6921 14893 6955
rect 14927 6921 14965 6955
rect 14999 6921 15037 6955
rect 15071 6921 15109 6955
rect 15143 6921 15181 6955
rect 15215 6921 15253 6955
rect 15287 6921 15325 6955
rect 15359 6921 15397 6955
rect 15431 6921 15469 6955
rect 15503 6921 15541 6955
rect 15575 6921 15613 6955
rect 15647 6921 15685 6955
rect 15719 6921 15757 6955
rect 15791 6921 15829 6955
rect 15863 6921 15901 6955
rect 15935 6921 15973 6955
rect 16007 6921 16045 6955
rect 16079 6921 16117 6955
rect 16151 6921 16189 6955
rect 16223 6921 16261 6955
rect 16295 6921 16333 6955
rect 16367 6921 16405 6955
rect 16439 6921 16477 6955
rect 16511 6921 16549 6955
rect 16583 6921 16621 6955
rect 16655 6921 16693 6955
rect 16727 6921 16765 6955
rect 16799 6921 16837 6955
rect 16871 6921 16909 6955
rect 16943 6921 16981 6955
rect 17015 6921 17053 6955
rect 17087 6921 17125 6955
rect 17159 6935 17218 6955
rect 17252 6935 17344 6969
rect 17378 6935 17384 6969
rect 17159 6921 17384 6935
rect 12628 6915 17384 6921
rect 12628 6896 12860 6915
tri 12860 6896 12879 6915 nw
tri 17164 6896 17183 6915 ne
rect 17183 6896 17384 6915
rect 12628 6882 12846 6896
tri 12846 6882 12860 6896 nw
tri 17183 6882 17197 6896 ne
rect 17197 6882 17218 6896
rect 12628 6870 12826 6882
rect 12628 6836 12634 6870
rect 12668 6836 12760 6870
rect 12794 6862 12826 6870
tri 12826 6862 12846 6882 nw
tri 17197 6867 17212 6882 ne
rect 17212 6862 17218 6882
rect 17252 6862 17344 6896
rect 17378 6862 17384 6896
rect 12794 6836 12800 6862
tri 12800 6836 12826 6862 nw
rect 12628 6797 12800 6836
rect 12628 6763 12634 6797
rect 12668 6763 12760 6797
rect 12794 6763 12800 6797
rect 12628 6724 12800 6763
rect 12628 6690 12634 6724
rect 12668 6690 12760 6724
rect 12794 6690 12800 6724
rect 17212 6823 17384 6862
rect 17212 6789 17218 6823
rect 17252 6789 17344 6823
rect 17378 6789 17384 6823
rect 17212 6750 17384 6789
rect 17212 6716 17218 6750
rect 17252 6716 17344 6750
rect 17378 6716 17384 6750
rect 12628 6651 12800 6690
rect 12628 6617 12634 6651
rect 12668 6617 12760 6651
rect 12794 6617 12800 6651
rect 12628 6578 12800 6617
rect 3266 6531 3311 6537
tri 3311 6531 3317 6537 nw
tri 3521 6531 3527 6537 se
rect 3527 6531 3690 6537
rect 2923 6351 3192 6515
rect 3266 6498 3298 6531
tri 3298 6518 3311 6531 nw
tri 3508 6518 3521 6531 se
rect 3521 6518 3690 6531
tri 3505 6515 3508 6518 se
rect 3508 6515 3690 6518
rect 12628 6544 12634 6578
rect 12668 6544 12760 6578
rect 12794 6544 12800 6578
rect 3460 6368 3488 6515
rect 12628 6505 12800 6544
rect 12628 6471 12634 6505
rect 12668 6471 12760 6505
rect 12794 6471 12800 6505
rect 12628 6432 12800 6471
rect 12628 6398 12634 6432
rect 12668 6398 12760 6432
rect 12794 6398 12800 6432
rect 2923 6339 3238 6351
rect 3414 6339 3690 6368
rect 12628 6359 12800 6398
rect 2923 6310 3192 6339
rect 3460 6310 3488 6339
rect 12628 6325 12634 6359
rect 12668 6325 12760 6359
rect 12794 6325 12800 6359
rect 2923 5180 3238 6310
rect 12628 6286 12800 6325
rect 12628 6252 12634 6286
rect 12668 6252 12760 6286
rect 12794 6252 12800 6286
rect 12628 6213 12800 6252
rect 12628 6179 12634 6213
rect 12668 6179 12760 6213
rect 12794 6179 12800 6213
rect 12628 6140 12800 6179
rect 12628 6106 12634 6140
rect 12668 6106 12760 6140
rect 12794 6106 12800 6140
rect 12628 6067 12800 6106
rect 12628 6033 12634 6067
rect 12668 6033 12760 6067
rect 12794 6033 12800 6067
rect 12628 5994 12800 6033
rect 12628 5960 12634 5994
rect 12668 5960 12760 5994
rect 12794 5960 12800 5994
rect 12628 5930 12800 5960
rect 11263 5909 11435 5915
rect 11315 5857 11383 5909
rect 11263 5845 11435 5857
rect 11315 5793 11383 5845
rect 11263 5780 11435 5793
rect 11315 5728 11383 5780
rect 11263 5715 11435 5728
rect 11315 5663 11383 5715
rect 11263 5650 11435 5663
rect 11315 5598 11383 5650
rect 11263 5585 11435 5598
rect 11315 5533 11383 5585
rect 11263 5527 11435 5533
rect 12680 5878 12748 5930
rect 12628 5859 12800 5878
rect 12680 5807 12748 5859
rect 12628 5787 12800 5807
rect 12680 5735 12748 5787
rect 12628 5702 12800 5735
rect 12628 5668 12634 5702
rect 12668 5668 12760 5702
rect 12794 5668 12800 5702
rect 12628 5629 12800 5668
rect 12628 5595 12634 5629
rect 12668 5595 12760 5629
rect 12794 5595 12800 5629
rect 12628 5556 12800 5595
rect 2923 5146 3198 5180
rect 3232 5146 3238 5180
rect 2923 5108 3238 5146
rect 2923 5074 3198 5108
rect 3232 5074 3238 5108
rect 2923 5040 3238 5074
rect 12628 5522 12634 5556
rect 12668 5522 12760 5556
rect 12794 5522 12800 5556
rect 12628 5483 12800 5522
rect 12628 5449 12634 5483
rect 12668 5449 12760 5483
rect 12794 5449 12800 5483
rect 12628 5410 12800 5449
rect 12628 5376 12634 5410
rect 12668 5376 12760 5410
rect 12794 5376 12800 5410
rect 12628 5337 12800 5376
rect 12628 5303 12634 5337
rect 12668 5303 12760 5337
rect 12794 5303 12800 5337
rect 12628 5264 12800 5303
rect 12628 5230 12634 5264
rect 12668 5230 12760 5264
rect 12794 5230 12800 5264
rect 12628 5191 12800 5230
rect 12628 5157 12634 5191
rect 12668 5157 12760 5191
rect 12794 5157 12800 5191
rect 12628 5118 12800 5157
rect 12628 5084 12634 5118
rect 12668 5084 12760 5118
rect 12794 5084 12800 5118
rect 2923 5006 2974 5040
rect 3008 5006 3046 5040
rect 3080 5006 3118 5040
rect 3152 5006 3238 5040
rect 2923 4887 3238 5006
rect 2014 4263 2026 4297
rect 2060 4263 2072 4297
rect 2014 4257 2072 4263
rect 2108 4309 2154 4321
rect 2108 4275 2114 4309
rect 2148 4275 2154 4309
tri 1972 4237 1979 4244 sw
tri 2101 4237 2108 4244 se
rect 2108 4237 2154 4275
tri 73 4203 76 4206 sw
rect 468 4203 474 4237
rect 508 4219 521 4237
tri 521 4219 539 4237 sw
tri 836 4219 854 4237 se
rect 854 4224 992 4237
rect 854 4219 879 4224
tri 879 4219 884 4224 nw
tri 962 4219 967 4224 ne
rect 967 4219 992 4224
tri 992 4219 1010 4237 sw
tri 1889 4219 1907 4237 se
rect 1907 4219 1926 4237
rect 508 4203 863 4219
tri 863 4203 879 4219 nw
tri 967 4209 977 4219 ne
rect 977 4209 1926 4219
tri 977 4203 983 4209 ne
rect 983 4203 1926 4209
rect 1960 4219 1979 4237
tri 1979 4219 1997 4237 sw
tri 2083 4219 2101 4237 se
rect 2101 4219 2114 4237
rect 1960 4203 2114 4219
rect 2148 4203 2154 4237
rect -104 4194 76 4203
tri 76 4194 85 4203 sw
rect 468 4197 857 4203
tri 857 4197 863 4203 nw
tri 983 4197 989 4203 ne
rect 989 4197 2154 4203
rect 468 4196 856 4197
tri 856 4196 857 4197 nw
tri 989 4196 990 4197 ne
rect 990 4196 2154 4197
rect 468 4194 854 4196
tri 854 4194 856 4196 nw
rect 896 4194 942 4196
tri 942 4194 944 4196 sw
tri 990 4194 992 4196 ne
rect 992 4194 2154 4196
rect -104 4191 85 4194
tri 85 4191 88 4194 sw
rect 468 4191 851 4194
tri 851 4191 854 4194 nw
rect 896 4191 944 4194
tri 944 4191 947 4194 sw
tri 992 4191 995 4194 ne
rect 995 4191 2154 4194
rect -104 4185 88 4191
tri 88 4185 94 4191 sw
rect 896 4185 947 4191
tri 947 4185 953 4191 sw
rect -104 4184 94 4185
tri 94 4184 95 4185 sw
rect 896 4184 953 4185
rect -104 4150 95 4184
tri 95 4150 129 4184 sw
rect 896 4150 902 4184
rect 936 4177 953 4184
tri 953 4177 961 4185 sw
rect 936 4175 961 4177
tri 961 4175 963 4177 sw
rect 2477 4175 2483 4355
rect 2599 4175 2605 4355
rect 2831 4835 2837 4887
rect 2889 4835 2895 4887
rect 2831 4823 2895 4835
rect 2831 4771 2837 4823
rect 2889 4771 2895 4823
rect 2831 4753 2895 4771
rect 2832 4751 2894 4752
rect 2831 4715 2895 4751
rect 2832 4714 2894 4715
rect 2831 4701 2895 4713
rect 2831 4667 2837 4701
rect 2871 4667 2895 4701
rect 2831 4627 2895 4667
rect 2831 4593 2837 4627
rect 2871 4593 2895 4627
rect 2831 4552 2895 4593
rect 2831 4518 2837 4552
rect 2871 4518 2895 4552
rect 2831 4477 2895 4518
rect 2831 4443 2837 4477
rect 2871 4443 2895 4477
rect 2831 4402 2895 4443
rect 2831 4368 2837 4402
rect 2871 4368 2895 4402
rect 2831 4327 2895 4368
rect 2831 4293 2837 4327
rect 2871 4293 2895 4327
rect 2831 4252 2895 4293
rect 2831 4218 2837 4252
rect 2871 4218 2895 4252
rect 2831 4177 2895 4218
rect 936 4153 963 4175
tri 963 4153 985 4175 sw
rect 936 4150 2262 4153
rect -104 4147 129 4150
tri 129 4147 132 4150 sw
rect 896 4147 2262 4150
rect -104 4140 132 4147
tri 132 4140 139 4147 sw
rect -104 4128 139 4140
tri 139 4128 151 4140 sw
rect 468 4128 514 4140
rect -104 4094 151 4128
tri 151 4094 185 4128 sw
rect 468 4094 474 4128
rect 508 4094 514 4128
rect -104 4078 185 4094
tri 185 4078 201 4094 sw
rect -104 4068 201 4078
tri 201 4068 211 4078 sw
rect -104 4058 211 4068
tri 211 4058 221 4068 sw
rect 468 4058 514 4094
rect 896 4113 2144 4147
rect 2178 4113 2216 4147
rect 2250 4113 2262 4147
rect 896 4112 2262 4113
rect 896 4078 902 4112
rect 936 4107 2262 4112
rect 2831 4143 2837 4177
rect 2871 4143 2895 4177
rect 936 4102 978 4107
tri 978 4102 983 4107 nw
rect 2831 4102 2895 4143
rect 936 4078 944 4102
rect 896 4068 944 4078
tri 944 4068 978 4102 nw
rect 2831 4068 2837 4102
rect 2871 4068 2895 4102
rect 896 4066 942 4068
tri 942 4066 944 4068 nw
tri 514 4058 519 4063 sw
rect -104 4056 221 4058
tri 221 4056 223 4058 sw
rect 468 4056 519 4058
tri 519 4056 521 4058 sw
rect -104 4022 223 4056
tri 223 4022 257 4056 sw
rect 468 4022 474 4056
rect 508 4054 521 4056
tri 521 4054 523 4056 sw
tri 1722 4054 1724 4056 se
rect 1724 4054 1854 4056
rect 508 4050 523 4054
tri 523 4050 527 4054 sw
tri 1718 4050 1722 4054 se
rect 1722 4050 1854 4054
rect 508 4038 527 4050
tri 527 4038 539 4050 sw
tri 1706 4038 1718 4050 se
rect 1718 4038 1736 4050
rect 508 4022 1736 4038
rect -104 4016 257 4022
tri 257 4016 263 4022 sw
rect 468 4016 1736 4022
rect 1770 4016 1808 4050
rect 1842 4016 1854 4050
rect -104 4010 263 4016
tri 263 4010 269 4016 sw
rect 468 4010 1854 4016
rect 2831 4027 2895 4068
rect -104 3993 269 4010
tri 269 3993 286 4010 sw
rect 2831 3993 2837 4027
rect 2871 3993 2895 4027
rect -104 3982 286 3993
tri 286 3982 297 3993 sw
rect -104 3970 2166 3982
rect -104 3936 80 3970
rect 114 3936 1438 3970
rect 1472 3936 2166 3970
rect -104 3898 2166 3936
rect -104 3864 80 3898
rect 114 3864 1438 3898
rect 1472 3869 2166 3898
rect 1472 3864 1832 3869
rect -104 3835 1832 3864
rect 1866 3835 1904 3869
rect 1938 3835 1976 3869
rect 2010 3835 2048 3869
rect 2082 3835 2120 3869
rect 2154 3835 2166 3869
rect -104 3826 2166 3835
rect -104 3792 80 3826
rect 114 3792 1438 3826
rect 1472 3792 2166 3826
rect -104 3780 2166 3792
rect 2831 3952 2895 3993
rect 2831 3918 2837 3952
rect 2871 3918 2895 3952
rect 2831 3877 2895 3918
rect 2831 3843 2837 3877
rect 2871 3843 2895 3877
rect 2831 3802 2895 3843
rect -104 3768 -59 3780
tri -59 3768 -47 3780 nw
rect 2831 3768 2837 3802
rect 2871 3768 2895 3802
rect -104 3727 -100 3768
tri -100 3727 -59 3768 nw
tri 1372 3727 1385 3740 se
rect 1385 3727 2162 3740
tri 2162 3727 2175 3740 sw
rect 2831 3727 2895 3768
tri -104 3723 -100 3727 nw
tri 1368 3723 1372 3727 se
rect 1372 3723 2175 3727
tri 2175 3723 2179 3727 sw
tri 1363 3718 1368 3723 se
rect 1368 3718 2179 3723
tri 2179 3718 2184 3723 sw
rect 213 3716 2305 3718
tri 2305 3716 2307 3718 sw
rect 213 3712 1582 3716
rect 213 3678 225 3712
rect 259 3678 297 3712
rect 331 3678 605 3712
rect 639 3678 677 3712
rect 711 3706 1582 3712
rect 711 3678 1126 3706
rect 213 3672 1126 3678
rect 1160 3672 1582 3706
rect 213 3664 1582 3672
rect 1634 3664 1646 3716
rect 1698 3664 1894 3716
rect 1946 3664 1958 3716
rect 2010 3693 2307 3716
tri 2307 3693 2330 3716 sw
rect 2831 3693 2837 3727
rect 2871 3693 2895 3727
rect 2010 3682 2330 3693
tri 2330 3682 2341 3693 sw
rect 2010 3679 2341 3682
tri 2341 3679 2344 3682 sw
rect 2831 3681 2895 3693
rect 2832 3679 2894 3680
rect 2923 4771 2971 4887
rect 3151 4771 3238 4887
rect 2923 4728 3238 4771
rect 2923 4694 2974 4728
rect 3008 4694 3046 4728
rect 3080 4694 3118 4728
rect 3152 4694 3238 4728
rect 2923 4618 3238 4694
rect 2923 4584 2974 4618
rect 3008 4584 3046 4618
rect 3080 4584 3118 4618
rect 3152 4584 3238 4618
rect 2923 4306 3238 4584
rect 2923 4272 2974 4306
rect 3008 4272 3046 4306
rect 3080 4272 3118 4306
rect 3152 4272 3238 4306
rect 2923 3994 3238 4272
rect 2923 3960 2974 3994
rect 3008 3960 3046 3994
rect 3080 3960 3118 3994
rect 3152 3960 3238 3994
rect 2923 3682 3238 3960
rect 2010 3667 2344 3679
tri 2344 3667 2356 3679 sw
rect 2010 3664 2356 3667
rect 213 3648 1540 3664
tri 1540 3648 1556 3664 nw
tri 2038 3648 2054 3664 ne
rect 2054 3648 2356 3664
rect 213 3643 1535 3648
tri 1535 3643 1540 3648 nw
tri 2054 3643 2059 3648 ne
rect 2059 3643 2356 3648
rect 2923 3648 2974 3682
rect 3008 3648 3046 3682
rect 3080 3648 3118 3682
rect 3152 3648 3238 3682
rect 213 3634 1526 3643
tri 1526 3634 1535 3643 nw
tri 2059 3634 2068 3643 ne
rect 2068 3634 2356 3643
tri -104 3600 -95 3609 sw
rect 213 3600 1126 3634
rect 1160 3628 1520 3634
tri 1520 3628 1526 3634 nw
rect 1160 3600 1276 3628
rect -104 3594 -95 3600
tri -95 3594 -89 3600 sw
rect 213 3594 1276 3600
rect 1310 3594 1348 3628
rect 1382 3594 1486 3628
tri 1486 3594 1520 3628 nw
rect -104 3588 -89 3594
tri -89 3588 -83 3594 sw
rect -104 3582 -83 3588
tri -83 3582 -77 3588 sw
rect 213 3582 1474 3594
tri 1474 3582 1486 3594 nw
rect 1576 3582 1582 3634
rect 1634 3582 1646 3634
rect 1698 3582 1706 3634
rect 1888 3582 1894 3634
rect 1946 3582 1958 3634
rect 2010 3582 2018 3634
tri 2068 3628 2074 3634 ne
rect 2074 3628 2356 3634
tri 2074 3594 2108 3628 ne
rect 2108 3594 2212 3628
rect 2246 3594 2284 3628
rect 2318 3594 2356 3628
tri 2108 3588 2114 3594 ne
rect 2114 3588 2356 3594
rect 2832 3642 2894 3643
rect 2923 3642 3238 3648
rect -104 3580 -77 3582
tri -77 3580 -75 3582 sw
rect -104 3552 -75 3580
tri -75 3552 -47 3580 sw
rect -104 3540 1582 3552
rect -104 3506 1156 3540
rect 1190 3506 1468 3540
rect 1502 3506 1582 3540
rect -104 3500 1582 3506
rect 1634 3500 1646 3552
rect 1698 3540 1894 3552
rect 1698 3506 1780 3540
rect 1814 3506 1894 3540
rect 1698 3500 1894 3506
rect 1946 3500 1958 3552
rect 2010 3540 2132 3552
rect 2010 3506 2092 3540
rect 2126 3506 2132 3540
rect 2010 3500 2132 3506
rect -104 3468 2132 3500
rect -104 3434 1156 3468
rect 1190 3434 1468 3468
rect 1502 3434 1780 3468
rect 1814 3434 2092 3468
rect 2126 3434 2132 3468
rect -104 3396 2132 3434
rect -104 3362 1156 3396
rect 1190 3362 1468 3396
rect 1502 3362 1780 3396
rect 1814 3362 2092 3396
rect 2126 3362 2132 3396
rect -104 3354 2132 3362
rect -104 3350 1147 3354
rect -104 3346 353 3350
tri 353 3346 357 3350 nw
tri 1107 3346 1111 3350 ne
rect 1111 3346 1147 3350
rect -104 3310 317 3346
tri 317 3310 353 3346 nw
tri 1111 3310 1147 3346 ne
rect -104 3168 175 3310
tri 175 3168 317 3310 nw
rect 1199 3350 1459 3354
rect 1199 3346 1235 3350
tri 1235 3346 1239 3350 nw
tri 1419 3346 1423 3350 ne
rect 1423 3346 1459 3350
tri 1199 3310 1235 3346 nw
tri 1423 3310 1459 3346 ne
rect 1147 3290 1199 3302
rect 1147 3226 1199 3238
rect -104 3087 94 3168
tri 94 3087 175 3168 nw
rect 1147 3093 1199 3174
rect -104 845 73 3087
tri 73 3066 94 3087 nw
rect 1147 3029 1199 3041
rect 1147 2965 1199 2977
rect 1147 2909 1156 2913
rect 1190 2909 1199 2913
rect 1147 2901 1199 2909
rect 1147 2837 1156 2849
rect 1190 2837 1199 2849
rect 1147 2799 1199 2837
rect 1147 2765 1156 2799
rect 1190 2765 1199 2799
rect 1147 2727 1199 2765
rect 1147 2693 1156 2727
rect 1190 2693 1199 2727
rect 1147 2681 1199 2693
rect 1511 3350 1771 3354
rect 1511 3346 1547 3350
tri 1547 3346 1551 3350 nw
tri 1731 3346 1735 3350 ne
rect 1735 3346 1771 3350
tri 1511 3310 1547 3346 nw
tri 1735 3310 1771 3346 ne
rect 1459 3290 1511 3302
rect 1459 3226 1511 3238
rect 1459 3093 1511 3174
rect 1459 3029 1511 3041
rect 1459 2965 1511 2977
rect 1459 2909 1468 2913
rect 1502 2909 1511 2913
rect 1459 2901 1511 2909
rect 1459 2837 1468 2849
rect 1502 2837 1511 2849
rect 1459 2799 1511 2837
rect 1459 2765 1468 2799
rect 1502 2765 1511 2799
rect 1459 2727 1511 2765
rect 1459 2693 1468 2727
rect 1502 2693 1511 2727
rect 1459 2681 1511 2693
rect 1823 3350 2080 3354
rect 1823 3346 1859 3350
tri 1859 3346 1863 3350 nw
tri 2040 3346 2044 3350 ne
rect 2044 3346 2080 3350
tri 1823 3310 1859 3346 nw
tri 2044 3310 2080 3346 ne
rect 1771 3290 1823 3302
rect 1771 3226 1823 3238
rect 1771 3093 1823 3174
rect 1771 3029 1823 3041
rect 1771 2965 1823 2977
rect 1771 2909 1780 2913
rect 1814 2909 1823 2913
rect 1771 2901 1823 2909
rect 1771 2837 1780 2849
rect 1814 2837 1823 2849
rect 1771 2799 1823 2837
rect 1771 2765 1780 2799
rect 1814 2765 1823 2799
rect 1771 2727 1823 2765
rect 1771 2693 1780 2727
rect 1814 2693 1823 2727
rect 1771 2681 1823 2693
rect 2080 3290 2132 3302
rect 2080 3226 2132 3238
rect 2080 3093 2132 3174
rect 2485 3358 2487 3383
rect 2485 3346 2603 3358
rect 2485 3168 2491 3346
rect 2597 3168 2603 3346
rect 2485 3156 2603 3168
rect 2831 3308 2895 3641
rect 3164 3614 3238 3642
rect 3164 3580 3198 3614
rect 3232 3580 3238 3614
rect 3164 3542 3238 3580
rect 3164 3508 3198 3542
rect 3232 3508 3238 3542
rect 3164 3496 3238 3508
rect 3164 3441 3183 3496
tri 3183 3441 3238 3496 nw
rect 3416 4946 3661 5046
rect 3662 4947 3663 5045
rect 3699 4947 3700 5045
rect 3701 5040 4173 5046
rect 3701 5006 3713 5040
rect 3747 5006 3796 5040
rect 3830 5006 3879 5040
rect 3913 5006 3962 5040
rect 3996 5006 4045 5040
rect 4079 5006 4127 5040
rect 4161 5006 4173 5040
rect 3701 4946 4173 5006
rect 3416 4938 3649 4946
tri 3649 4938 3657 4946 nw
tri 3857 4938 3865 4946 ne
rect 3865 4938 4173 4946
rect 3416 4908 3619 4938
tri 3619 4908 3649 4938 nw
tri 3865 4908 3895 4938 ne
rect 3895 4908 4173 4938
rect 3416 4906 3617 4908
tri 3617 4906 3619 4908 nw
tri 3895 4906 3897 4908 ne
rect 3897 4906 4173 4908
rect 3416 3727 3614 4906
tri 3614 4903 3617 4906 nw
tri 3897 4903 3900 4906 ne
rect 3647 4884 3844 4890
rect 3647 4850 3659 4884
rect 3693 4850 3798 4884
rect 3832 4850 3844 4884
rect 3647 4844 3844 4850
tri 3887 4764 3900 4777 se
rect 3900 4764 4173 4906
rect 12628 5045 12800 5084
rect 12628 5011 12634 5045
rect 12668 5011 12760 5045
rect 12794 5011 12800 5045
rect 12628 4972 12800 5011
rect 12628 4938 12634 4972
rect 12668 4938 12760 4972
rect 12794 4938 12800 4972
rect 12628 4899 12800 4938
tri 3885 4762 3887 4764 se
rect 3887 4762 4173 4764
tri 3881 4758 3885 4762 se
rect 3885 4758 4173 4762
rect 4229 4835 4235 4887
rect 4287 4835 4293 4887
rect 4229 4823 4293 4835
rect 4229 4771 4235 4823
rect 4287 4771 4293 4823
rect 4229 4764 4286 4771
tri 4286 4764 4293 4771 nw
rect 12628 4865 12634 4899
rect 12668 4865 12760 4899
rect 12794 4865 12800 4899
rect 12628 4826 12800 4865
rect 12628 4792 12634 4826
rect 12668 4792 12760 4826
rect 12794 4792 12800 4826
rect 4229 4762 4284 4764
tri 4284 4762 4286 4764 nw
rect 4229 4760 4282 4762
tri 4282 4760 4284 4762 nw
tri 4281 4759 4282 4760 nw
rect 4230 4758 4280 4759
tri 3876 4753 3881 4758 se
rect 3881 4753 4173 4758
tri 3857 4734 3876 4753 se
rect 3876 4734 4173 4753
rect 3701 4728 4173 4734
rect 3701 4694 3713 4728
rect 3747 4694 3796 4728
rect 3830 4694 3879 4728
rect 3913 4694 3962 4728
rect 3996 4694 4045 4728
rect 4079 4694 4127 4728
rect 4161 4694 4173 4728
rect 12628 4753 12800 4792
rect 3701 4688 4173 4694
rect 4230 4721 4280 4722
rect 4229 4708 4281 4720
rect 4229 4674 4235 4708
rect 4269 4674 4281 4708
rect 3900 4618 4173 4624
rect 3900 4584 3912 4618
rect 3946 4584 4020 4618
rect 4054 4584 4127 4618
rect 4161 4584 4173 4618
rect 3642 4462 3844 4468
rect 3642 4428 3654 4462
rect 3688 4428 3726 4462
rect 3760 4428 3798 4462
rect 3832 4428 3844 4462
rect 3642 4150 3844 4428
rect 3642 4116 3654 4150
rect 3688 4116 3726 4150
rect 3760 4116 3798 4150
rect 3832 4116 3844 4150
rect 3642 3838 3844 4116
rect 3642 3804 3654 3838
rect 3688 3804 3726 3838
rect 3760 3804 3798 3838
rect 3832 3804 3844 3838
rect 3642 3798 3844 3804
rect 3900 4306 4173 4584
rect 4229 4591 4281 4674
rect 4229 4557 4235 4591
rect 4269 4557 4281 4591
rect 4229 4545 4281 4557
rect 12628 4719 12634 4753
rect 12668 4719 12760 4753
rect 12794 4719 12800 4753
rect 12628 4680 12800 4719
rect 12628 4646 12634 4680
rect 12668 4646 12760 4680
rect 12794 4646 12800 4680
rect 12628 4607 12800 4646
rect 12628 4573 12634 4607
rect 12668 4573 12760 4607
rect 12794 4573 12800 4607
rect 12628 4534 12800 4573
rect 3900 4272 3912 4306
rect 3946 4272 4020 4306
rect 4054 4272 4127 4306
rect 4161 4272 4173 4306
rect 3900 3994 4173 4272
rect 3900 3960 3912 3994
rect 3946 3960 4020 3994
rect 4054 3960 4127 3994
rect 4161 3960 4173 3994
tri 3884 3770 3900 3786 se
rect 3900 3770 4173 3960
tri 3849 3735 3884 3770 se
rect 3884 3735 4173 3770
tri 3614 3727 3622 3735 sw
tri 3841 3727 3849 3735 se
rect 3849 3727 4173 3735
rect 3416 3693 3622 3727
tri 3622 3693 3656 3727 sw
tri 3807 3693 3841 3727 se
rect 3841 3693 4173 3727
rect 3416 3688 3656 3693
tri 3656 3688 3661 3693 sw
tri 3802 3688 3807 3693 se
rect 3807 3688 4173 3693
rect 3416 3682 3661 3688
tri 3661 3682 3667 3688 sw
tri 3796 3682 3802 3688 se
rect 3802 3682 4173 3688
rect 3416 3648 3667 3682
tri 3667 3648 3701 3682 sw
tri 3762 3648 3796 3682 se
rect 3796 3648 3910 3682
rect 3944 3648 3983 3682
rect 4017 3648 4055 3682
rect 4089 3648 4127 3682
rect 4161 3648 4173 3682
rect 4229 4511 4281 4517
rect 4229 4447 4281 4459
rect 12628 4500 12634 4534
rect 12668 4500 12760 4534
rect 12794 4500 12800 4534
rect 12628 4461 12800 4500
rect 4229 4389 4281 4395
rect 11189 4445 11394 4450
rect 11189 4393 11195 4445
rect 11247 4393 11266 4445
rect 11318 4393 11336 4445
rect 11388 4393 11394 4445
rect 11189 4388 11394 4393
rect 12628 4427 12634 4461
rect 12668 4427 12760 4461
rect 12794 4427 12800 4461
rect 12628 4388 12800 4427
rect 4230 4387 4280 4388
rect 4229 4351 4281 4387
rect 4230 4350 4280 4351
rect 4229 4337 4281 4349
rect 4229 4303 4235 4337
rect 4269 4303 4281 4337
rect 4229 4297 4281 4303
rect 4229 4261 4275 4297
tri 4275 4291 4281 4297 nw
rect 12628 4354 12634 4388
rect 12668 4354 12760 4388
rect 12794 4354 12800 4388
rect 12628 4314 12800 4354
rect 4229 4227 4235 4261
rect 4269 4227 4275 4261
rect 4229 4185 4275 4227
rect 4229 4151 4235 4185
rect 4269 4151 4275 4185
rect 4229 4109 4275 4151
rect 4229 4075 4235 4109
rect 4269 4075 4275 4109
rect 4229 4033 4275 4075
rect 4229 3999 4235 4033
rect 4269 3999 4275 4033
rect 4229 3957 4275 3999
rect 4229 3923 4235 3957
rect 4269 3923 4275 3957
rect 4229 3881 4275 3923
rect 12628 4280 12634 4314
rect 12668 4280 12760 4314
rect 12794 4280 12800 4314
rect 12628 4240 12800 4280
rect 12628 4206 12634 4240
rect 12668 4206 12760 4240
rect 12794 4206 12800 4240
rect 12628 4166 12800 4206
rect 12628 4132 12634 4166
rect 12668 4132 12760 4166
rect 12794 4132 12800 4166
rect 12628 4092 12800 4132
rect 12628 4058 12634 4092
rect 12668 4058 12760 4092
rect 12794 4058 12800 4092
rect 12628 4018 12800 4058
rect 12628 3984 12634 4018
rect 12668 3984 12760 4018
rect 12794 3984 12800 4018
rect 13026 6685 16991 6691
rect 13026 6651 13038 6685
rect 13072 6651 13111 6685
rect 13145 6651 13184 6685
rect 13218 6651 13257 6685
rect 13291 6651 13330 6685
rect 13364 6651 13403 6685
rect 13437 6651 13476 6685
rect 13510 6651 13549 6685
rect 13583 6651 13622 6685
rect 13656 6651 13695 6685
rect 13729 6651 13768 6685
rect 13802 6651 13841 6685
rect 13875 6651 13914 6685
rect 13948 6651 13987 6685
rect 14021 6651 14060 6685
rect 14094 6651 14133 6685
rect 14167 6651 14206 6685
rect 14240 6651 14279 6685
rect 14313 6651 14352 6685
rect 14386 6651 14425 6685
rect 14459 6651 14497 6685
rect 14531 6651 14569 6685
rect 14603 6651 14641 6685
rect 14675 6651 14713 6685
rect 14747 6651 14785 6685
rect 14819 6651 14857 6685
rect 14891 6651 14929 6685
rect 14963 6651 15001 6685
rect 15035 6651 15073 6685
rect 15107 6651 15145 6685
rect 15179 6651 15217 6685
rect 15251 6651 15289 6685
rect 15323 6651 15361 6685
rect 15395 6651 15433 6685
rect 15467 6651 15505 6685
rect 15539 6651 15577 6685
rect 15611 6651 15649 6685
rect 15683 6651 15721 6685
rect 15755 6651 15793 6685
rect 15827 6651 15865 6685
rect 15899 6651 15937 6685
rect 15971 6651 16009 6685
rect 16043 6651 16081 6685
rect 16115 6651 16153 6685
rect 16187 6651 16225 6685
rect 16259 6651 16297 6685
rect 16331 6651 16369 6685
rect 16403 6651 16441 6685
rect 16475 6651 16513 6685
rect 16547 6651 16585 6685
rect 16619 6651 16657 6685
rect 16691 6651 16729 6685
rect 16763 6651 16801 6685
rect 16835 6651 16873 6685
rect 16907 6651 16945 6685
rect 16979 6651 16991 6685
rect 13026 6571 16991 6651
rect 13026 6537 13038 6571
rect 13072 6537 13111 6571
rect 13145 6537 13184 6571
rect 13218 6537 13257 6571
rect 13291 6537 13330 6571
rect 13364 6537 13403 6571
rect 13437 6537 13476 6571
rect 13510 6537 13549 6571
rect 13583 6537 13622 6571
rect 13656 6537 13695 6571
rect 13729 6537 13768 6571
rect 13802 6537 13841 6571
rect 13875 6537 13914 6571
rect 13948 6537 13987 6571
rect 14021 6537 14060 6571
rect 14094 6537 14133 6571
rect 14167 6537 14206 6571
rect 14240 6537 14279 6571
rect 14313 6537 14352 6571
rect 14386 6537 14425 6571
rect 14459 6537 14497 6571
rect 14531 6537 14569 6571
rect 14603 6537 14641 6571
rect 14675 6537 14713 6571
rect 14747 6537 14785 6571
rect 14819 6537 14857 6571
rect 14891 6537 14929 6571
rect 14963 6537 15001 6571
rect 15035 6537 15073 6571
rect 15107 6537 15145 6571
rect 15179 6537 15217 6571
rect 15251 6537 15289 6571
rect 15323 6537 15361 6571
rect 15395 6537 15433 6571
rect 15467 6537 15505 6571
rect 15539 6537 15577 6571
rect 15611 6537 15649 6571
rect 15683 6537 15721 6571
rect 15755 6537 15793 6571
rect 15827 6537 15865 6571
rect 15899 6537 15937 6571
rect 15971 6537 16009 6571
rect 16043 6537 16081 6571
rect 16115 6537 16153 6571
rect 16187 6537 16225 6571
rect 16259 6537 16297 6571
rect 16331 6537 16369 6571
rect 16403 6537 16441 6571
rect 16475 6537 16513 6571
rect 16547 6537 16585 6571
rect 16619 6537 16657 6571
rect 16691 6537 16729 6571
rect 16763 6537 16801 6571
rect 16835 6537 16873 6571
rect 16907 6537 16945 6571
rect 16979 6537 16991 6571
rect 13026 6531 16991 6537
rect 13026 6502 13202 6531
tri 13202 6502 13231 6531 nw
tri 16789 6502 16818 6531 ne
rect 16818 6502 16991 6531
rect 13026 6497 13197 6502
tri 13197 6497 13202 6502 nw
tri 16818 6497 16823 6502 ne
rect 16823 6497 16991 6502
rect 13026 6490 13190 6497
tri 13190 6490 13197 6497 nw
tri 16823 6490 16830 6497 ne
rect 16830 6490 16991 6497
rect 13026 6456 13032 6490
rect 13066 6456 13146 6490
rect 13180 6489 13189 6490
tri 13189 6489 13190 6490 nw
tri 16830 6489 16831 6490 ne
rect 13180 6456 13186 6489
tri 13186 6486 13189 6489 nw
rect 13026 6418 13186 6456
rect 13026 6384 13032 6418
rect 13066 6384 13146 6418
rect 13180 6384 13186 6418
rect 16831 6456 16837 6490
rect 16871 6456 16951 6490
rect 16985 6456 16991 6490
rect 16831 6418 16991 6456
rect 13026 6346 13186 6384
rect 13026 6312 13032 6346
rect 13066 6312 13146 6346
rect 13180 6312 13186 6346
rect 13026 6274 13186 6312
rect 13026 6240 13032 6274
rect 13066 6240 13146 6274
rect 13180 6240 13186 6274
rect 13026 6202 13186 6240
rect 13026 6168 13032 6202
rect 13066 6168 13146 6202
rect 13180 6168 13186 6202
rect 13026 6130 13186 6168
rect 13026 6096 13032 6130
rect 13066 6096 13146 6130
rect 13180 6096 13186 6130
rect 13026 6058 13186 6096
rect 13026 6024 13032 6058
rect 13066 6024 13146 6058
rect 13180 6024 13186 6058
rect 13026 5986 13186 6024
rect 13026 5952 13032 5986
rect 13066 5952 13146 5986
rect 13180 5952 13186 5986
rect 13026 5914 13186 5952
rect 13026 5880 13032 5914
rect 13066 5880 13146 5914
rect 13180 5880 13186 5914
rect 13026 5842 13186 5880
rect 13026 5808 13032 5842
rect 13066 5808 13146 5842
rect 13180 5808 13186 5842
rect 13026 5770 13186 5808
rect 13026 5736 13032 5770
rect 13066 5736 13146 5770
rect 13180 5736 13186 5770
rect 13026 5698 13186 5736
rect 13026 5664 13032 5698
rect 13066 5664 13146 5698
rect 13180 5664 13186 5698
rect 13026 5626 13186 5664
rect 13026 5592 13032 5626
rect 13066 5592 13146 5626
rect 13180 5592 13186 5626
rect 13026 5554 13186 5592
rect 13026 5520 13032 5554
rect 13066 5520 13146 5554
rect 13180 5520 13186 5554
rect 13026 5482 13186 5520
rect 13026 5448 13032 5482
rect 13066 5448 13146 5482
rect 13180 5448 13186 5482
rect 13026 5410 13186 5448
rect 13026 5376 13032 5410
rect 13066 5376 13146 5410
rect 13180 5376 13186 5410
rect 13026 5338 13186 5376
rect 13026 5304 13032 5338
rect 13066 5304 13146 5338
rect 13180 5304 13186 5338
rect 13026 5266 13186 5304
rect 13026 5232 13032 5266
rect 13066 5232 13146 5266
rect 13180 5232 13186 5266
rect 13026 5194 13186 5232
rect 13026 5160 13032 5194
rect 13066 5160 13146 5194
rect 13180 5160 13186 5194
rect 13026 5122 13186 5160
rect 13026 5088 13032 5122
rect 13066 5088 13146 5122
rect 13180 5088 13186 5122
rect 13026 5050 13186 5088
rect 13026 5016 13032 5050
rect 13066 5016 13146 5050
rect 13180 5016 13186 5050
rect 13026 4978 13186 5016
rect 13026 4944 13032 4978
rect 13066 4944 13146 4978
rect 13180 4944 13186 4978
rect 13026 4906 13186 4944
rect 13026 4872 13032 4906
rect 13066 4872 13146 4906
rect 13180 4872 13186 4906
rect 13026 4834 13186 4872
rect 13026 4800 13032 4834
rect 13066 4800 13146 4834
rect 13180 4800 13186 4834
rect 13026 4762 13186 4800
rect 13026 4728 13032 4762
rect 13066 4728 13146 4762
rect 13180 4728 13186 4762
rect 13026 4690 13186 4728
rect 13026 4656 13032 4690
rect 13066 4656 13146 4690
rect 13180 4656 13186 4690
rect 13026 4618 13186 4656
rect 13026 4584 13032 4618
rect 13066 4584 13146 4618
rect 13180 4584 13186 4618
rect 13026 4546 13186 4584
rect 13026 4512 13032 4546
rect 13066 4512 13146 4546
rect 13180 4512 13186 4546
rect 13026 4474 13186 4512
rect 13026 4440 13032 4474
rect 13066 4440 13146 4474
rect 13180 4440 13186 4474
rect 13026 4402 13186 4440
rect 13026 4368 13032 4402
rect 13066 4368 13146 4402
rect 13180 4368 13186 4402
rect 13026 4330 13186 4368
rect 13026 4296 13032 4330
rect 13066 4296 13146 4330
rect 13180 4296 13186 4330
rect 13326 6392 16690 6397
rect 13326 6391 13976 6392
rect 13326 6357 13404 6391
rect 13438 6357 13476 6391
rect 13510 6357 13548 6391
rect 13582 6357 13620 6391
rect 13654 6357 13692 6391
rect 13726 6357 13764 6391
rect 13798 6357 13836 6391
rect 13870 6357 13908 6391
rect 13942 6357 13976 6391
rect 13326 6351 13976 6357
rect 13326 6346 13401 6351
tri 13401 6346 13406 6351 nw
tri 13917 6346 13922 6351 ne
rect 13922 6346 13976 6351
rect 13326 6340 13395 6346
tri 13395 6340 13401 6346 nw
tri 13922 6340 13928 6346 ne
rect 13928 6340 13976 6346
rect 14028 6340 14040 6392
rect 14092 6340 14104 6392
rect 14156 6391 16690 6392
rect 14158 6357 14196 6391
rect 14230 6357 14268 6391
rect 14302 6357 14340 6391
rect 14374 6357 14412 6391
rect 14446 6357 14484 6391
rect 14518 6357 14556 6391
rect 14590 6357 14628 6391
rect 14662 6357 14700 6391
rect 14734 6357 14772 6391
rect 14806 6357 14844 6391
rect 14878 6357 14916 6391
rect 14950 6357 14988 6391
rect 15022 6357 15060 6391
rect 15094 6357 15132 6391
rect 15166 6357 15204 6391
rect 15238 6357 15276 6391
rect 15310 6357 15348 6391
rect 15382 6357 15420 6391
rect 15454 6357 15492 6391
rect 15526 6357 15564 6391
rect 15598 6357 15636 6391
rect 15670 6357 15708 6391
rect 15742 6357 15780 6391
rect 15814 6357 15852 6391
rect 15886 6357 15924 6391
rect 15958 6357 15996 6391
rect 16030 6357 16068 6391
rect 16102 6357 16140 6391
rect 16174 6357 16213 6391
rect 16247 6357 16286 6391
rect 16320 6357 16359 6391
rect 16393 6357 16432 6391
rect 16466 6357 16505 6391
rect 16539 6357 16578 6391
rect 16612 6357 16690 6391
rect 14156 6351 16690 6357
rect 14156 6346 14168 6351
tri 14168 6346 14173 6351 nw
tri 16610 6346 16615 6351 ne
rect 16615 6346 16690 6351
rect 14156 6340 14162 6346
tri 14162 6340 14168 6346 nw
tri 16615 6340 16621 6346 ne
rect 16621 6340 16690 6346
rect 13326 6319 13374 6340
tri 13374 6319 13395 6340 nw
tri 16621 6319 16642 6340 ne
rect 16642 6319 16690 6340
rect 13326 6285 13332 6319
rect 13366 6318 13373 6319
tri 13373 6318 13374 6319 nw
tri 16642 6318 16643 6319 ne
rect 16643 6318 16650 6319
rect 13366 6285 13372 6318
tri 13372 6317 13373 6318 nw
rect 13326 6246 13372 6285
rect 13518 6296 13730 6318
tri 13730 6296 13752 6318 sw
tri 16643 6317 16644 6318 ne
rect 13518 6293 13752 6296
tri 13752 6293 13755 6296 sw
tri 14385 6293 14388 6296 se
rect 14388 6293 14451 6296
rect 13518 6287 14451 6293
rect 14503 6287 14515 6296
rect 14567 6287 14579 6296
rect 14631 6293 14637 6296
tri 14637 6293 14640 6296 sw
rect 14631 6287 16337 6293
rect 13326 6212 13332 6246
rect 13366 6212 13372 6246
rect 13326 6173 13372 6212
rect 13326 6139 13332 6173
rect 13366 6139 13372 6173
rect 13326 6100 13372 6139
rect 13326 6066 13332 6100
rect 13366 6066 13372 6100
rect 13326 6027 13372 6066
rect 13326 5993 13332 6027
rect 13366 5993 13372 6027
rect 13326 5954 13372 5993
rect 13326 5920 13332 5954
rect 13366 5920 13372 5954
rect 13326 5881 13372 5920
rect 13326 5847 13332 5881
rect 13366 5847 13372 5881
rect 13326 5808 13372 5847
rect 13326 5774 13332 5808
rect 13366 5774 13372 5808
rect 13326 5735 13372 5774
rect 13326 5701 13332 5735
rect 13366 5701 13372 5735
rect 13326 5662 13372 5701
rect 13326 5628 13332 5662
rect 13366 5628 13372 5662
rect 13326 5590 13372 5628
rect 13326 5556 13332 5590
rect 13366 5556 13372 5590
rect 13326 5518 13372 5556
rect 13326 5484 13332 5518
rect 13366 5484 13372 5518
rect 13326 5446 13372 5484
rect 13326 5412 13332 5446
rect 13366 5412 13372 5446
rect 13326 5374 13372 5412
rect 13326 5340 13332 5374
rect 13366 5340 13372 5374
rect 13326 5302 13372 5340
rect 13326 5268 13332 5302
rect 13366 5268 13372 5302
rect 13326 5230 13372 5268
rect 13326 5196 13332 5230
rect 13366 5196 13372 5230
rect 13326 5158 13372 5196
rect 13326 5124 13332 5158
rect 13366 5124 13372 5158
rect 13326 5086 13372 5124
rect 13326 5052 13332 5086
rect 13366 5052 13372 5086
rect 13326 5014 13372 5052
rect 13326 4980 13332 5014
rect 13366 4980 13372 5014
rect 13326 4942 13372 4980
rect 13326 4908 13332 4942
rect 13366 4908 13372 4942
rect 13326 4870 13372 4908
rect 13326 4836 13332 4870
rect 13366 4836 13372 4870
rect 13326 4798 13372 4836
rect 13326 4764 13332 4798
rect 13366 4764 13372 4798
rect 13326 4726 13372 4764
rect 13326 4692 13332 4726
rect 13366 4692 13372 4726
rect 13326 4654 13372 4692
rect 13444 6247 13490 6259
rect 13444 6213 13450 6247
rect 13484 6213 13490 6247
rect 13444 6171 13490 6213
rect 13444 6137 13450 6171
rect 13484 6137 13490 6171
rect 13444 6095 13490 6137
rect 13444 6061 13450 6095
rect 13484 6061 13490 6095
rect 13444 6018 13490 6061
rect 13444 5984 13450 6018
rect 13484 5984 13490 6018
rect 13444 5743 13490 5984
rect 13444 5709 13450 5743
rect 13484 5709 13490 5743
rect 13444 5667 13490 5709
rect 13444 5633 13450 5667
rect 13484 5633 13490 5667
rect 13444 5591 13490 5633
rect 13444 5557 13450 5591
rect 13484 5557 13490 5591
rect 13444 5514 13490 5557
rect 13444 5480 13450 5514
rect 13484 5480 13490 5514
rect 13444 5239 13490 5480
rect 13444 5205 13450 5239
rect 13484 5205 13490 5239
rect 13444 5163 13490 5205
rect 13444 5129 13450 5163
rect 13484 5129 13490 5163
rect 13444 5087 13490 5129
rect 13444 5053 13450 5087
rect 13484 5053 13490 5087
rect 13444 5010 13490 5053
rect 13444 4976 13450 5010
rect 13484 4976 13490 5010
rect 13444 4735 13490 4976
rect 13518 6253 13530 6287
rect 13564 6253 13603 6287
rect 13637 6253 13676 6287
rect 13710 6253 13749 6287
rect 13783 6253 13822 6287
rect 13856 6253 13895 6287
rect 13929 6253 13968 6287
rect 14002 6253 14041 6287
rect 14075 6253 14114 6287
rect 14148 6253 14187 6287
rect 14221 6253 14260 6287
rect 14294 6253 14333 6287
rect 14367 6253 14406 6287
rect 14440 6253 14451 6287
rect 14513 6253 14515 6287
rect 14659 6253 14698 6287
rect 14732 6253 14771 6287
rect 14805 6253 14844 6287
rect 14878 6253 14917 6287
rect 14951 6253 14990 6287
rect 15024 6253 15063 6287
rect 15097 6253 15136 6287
rect 15170 6253 15209 6287
rect 15243 6253 15282 6287
rect 15316 6253 15355 6287
rect 15389 6253 15427 6287
rect 15461 6253 15499 6287
rect 15533 6253 15571 6287
rect 15605 6253 15643 6287
rect 15677 6253 15715 6287
rect 15749 6253 15787 6287
rect 15821 6253 15859 6287
rect 15893 6253 15931 6287
rect 15965 6253 16003 6287
rect 16037 6253 16075 6287
rect 16109 6253 16147 6287
rect 16181 6253 16219 6287
rect 16253 6253 16291 6287
rect 16325 6253 16337 6287
rect 13518 6247 14451 6253
rect 13518 6245 13753 6247
tri 13753 6245 13755 6247 nw
tri 14386 6245 14388 6247 ne
rect 13518 6244 13752 6245
tri 13752 6244 13753 6245 nw
rect 14388 6244 14451 6247
rect 14503 6244 14515 6253
rect 14567 6244 14579 6253
rect 14631 6247 16337 6253
rect 14631 6244 14637 6247
tri 14637 6245 14639 6247 nw
rect 13518 5997 13730 6244
tri 13730 6222 13752 6244 nw
tri 16383 6141 16407 6165 se
rect 16407 6141 16543 6312
tri 14387 6140 14388 6141 se
rect 14388 6140 14451 6141
rect 13758 6137 13896 6140
tri 13896 6137 13899 6140 sw
tri 14384 6137 14387 6140 se
rect 14387 6137 14451 6140
rect 13758 6131 14451 6137
rect 14503 6131 14515 6141
rect 13758 6097 13770 6131
rect 13804 6097 13844 6131
rect 13878 6097 13918 6131
rect 13952 6097 13992 6131
rect 14026 6097 14066 6131
rect 14100 6097 14140 6131
rect 14174 6097 14214 6131
rect 14248 6097 14288 6131
rect 14322 6097 14362 6131
rect 14396 6097 14436 6131
rect 14503 6097 14510 6131
rect 13758 6091 14451 6097
rect 13758 6089 13897 6091
tri 13897 6089 13899 6091 nw
tri 14386 6089 14388 6091 ne
rect 14388 6089 14451 6091
rect 14503 6089 14515 6097
rect 14567 6089 14579 6141
rect 14631 6137 14637 6141
tri 14637 6137 14641 6141 sw
tri 16379 6137 16383 6141 se
rect 16383 6137 16543 6141
rect 14631 6131 16543 6137
rect 14631 6097 14658 6131
rect 14692 6097 14732 6131
rect 14766 6097 14806 6131
rect 14840 6097 14880 6131
rect 14914 6097 14954 6131
rect 14988 6097 15028 6131
rect 15062 6097 15102 6131
rect 15136 6097 15176 6131
rect 15210 6097 15250 6131
rect 15284 6097 15323 6131
rect 15357 6097 15396 6131
rect 15430 6097 15469 6131
rect 15503 6097 15542 6131
rect 15576 6097 15615 6131
rect 15649 6097 15688 6131
rect 15722 6097 15761 6131
rect 15795 6097 15834 6131
rect 15868 6097 15907 6131
rect 15941 6097 15980 6131
rect 16014 6097 16053 6131
rect 16087 6097 16126 6131
rect 16160 6097 16199 6131
rect 16233 6097 16272 6131
rect 16306 6097 16345 6131
rect 16379 6097 16418 6131
rect 16452 6097 16543 6131
rect 14631 6091 16543 6097
rect 14631 6089 14637 6091
tri 14637 6089 14639 6091 nw
tri 16370 6089 16372 6091 ne
rect 16372 6089 16543 6091
rect 13758 6088 13896 6089
tri 13896 6088 13897 6089 nw
tri 16372 6088 16373 6089 ne
rect 16373 6088 16543 6089
tri 16373 6069 16392 6088 ne
rect 16392 6069 16543 6088
tri 16392 6059 16402 6069 ne
rect 16402 6059 16543 6069
tri 16402 6058 16403 6059 ne
rect 16403 6058 16543 6059
tri 16403 6057 16404 6058 ne
tri 13730 5997 13739 6006 sw
rect 13518 5986 13739 5997
tri 13739 5986 13750 5997 sw
rect 13518 5981 13750 5986
tri 13750 5981 13755 5986 sw
rect 13518 5975 16337 5981
rect 13518 5941 13530 5975
rect 13564 5941 13603 5975
rect 13637 5941 13676 5975
rect 13710 5941 13749 5975
rect 13783 5941 13822 5975
rect 13856 5941 13895 5975
rect 13929 5941 13968 5975
rect 14002 5941 14041 5975
rect 14075 5941 14114 5975
rect 14148 5941 14187 5975
rect 14221 5941 14260 5975
rect 14294 5941 14333 5975
rect 14367 5941 14406 5975
rect 14440 5941 14479 5975
rect 14513 5941 14552 5975
rect 14586 5941 14625 5975
rect 14659 5941 14698 5975
rect 14732 5941 14771 5975
rect 14805 5941 14844 5975
rect 14878 5941 14917 5975
rect 14951 5941 14990 5975
rect 15024 5941 15063 5975
rect 15097 5941 15136 5975
rect 15170 5941 15209 5975
rect 15243 5941 15282 5975
rect 15316 5941 15355 5975
rect 15389 5941 15427 5975
rect 15461 5941 15499 5975
rect 15533 5941 15571 5975
rect 15605 5941 15643 5975
rect 15677 5941 15715 5975
rect 15749 5941 15787 5975
rect 15821 5941 15859 5975
rect 15893 5941 15931 5975
rect 15965 5941 16003 5975
rect 16037 5941 16075 5975
rect 16109 5941 16147 5975
rect 16181 5941 16219 5975
rect 16253 5941 16291 5975
rect 16325 5941 16337 5975
rect 13518 5935 16337 5941
rect 13518 5925 13745 5935
tri 13745 5925 13755 5935 nw
rect 13518 5914 13734 5925
tri 13734 5914 13745 5925 nw
rect 13518 5789 13730 5914
tri 13730 5910 13734 5914 nw
tri 13927 5887 13928 5888 se
rect 13928 5887 13991 5888
tri 13925 5885 13927 5887 se
rect 13927 5885 13991 5887
rect 13807 5879 13991 5885
rect 14043 5879 14055 5888
rect 14107 5879 14119 5888
rect 14171 5887 14177 5888
tri 14177 5887 14178 5888 sw
rect 14171 5885 14178 5887
tri 14178 5885 14180 5887 sw
rect 14171 5879 16339 5885
rect 13807 5845 13819 5879
rect 13853 5845 13892 5879
rect 13926 5845 13965 5879
rect 14107 5845 14111 5879
rect 14171 5845 14184 5879
rect 14218 5845 14257 5879
rect 14291 5845 14330 5879
rect 14364 5845 14403 5879
rect 14437 5845 14476 5879
rect 14510 5845 14549 5879
rect 14583 5845 14622 5879
rect 14656 5845 14695 5879
rect 14729 5845 14768 5879
rect 14802 5845 14841 5879
rect 14875 5845 14914 5879
rect 14948 5845 14987 5879
rect 15021 5845 15060 5879
rect 15094 5845 15133 5879
rect 15167 5845 15206 5879
rect 15240 5845 15279 5879
rect 15313 5845 15352 5879
rect 15386 5845 15425 5879
rect 15459 5845 15498 5879
rect 15532 5845 15571 5879
rect 15605 5845 15644 5879
rect 15678 5845 15717 5879
rect 15751 5845 15789 5879
rect 15823 5845 15861 5879
rect 15895 5845 15933 5879
rect 15967 5845 16005 5879
rect 16039 5845 16077 5879
rect 16111 5845 16149 5879
rect 16183 5845 16221 5879
rect 16255 5845 16293 5879
rect 16327 5845 16339 5879
rect 13807 5839 13991 5845
tri 13925 5836 13928 5839 ne
rect 13928 5836 13991 5839
rect 14043 5836 14055 5845
rect 14107 5836 14119 5845
rect 14171 5839 16339 5845
rect 14171 5836 14177 5839
tri 14177 5836 14180 5839 nw
tri 13730 5789 13755 5814 sw
rect 13518 5783 16337 5789
rect 13518 5749 13530 5783
rect 13564 5749 13603 5783
rect 13637 5749 13676 5783
rect 13710 5749 13749 5783
rect 13783 5749 13822 5783
rect 13856 5749 13895 5783
rect 13929 5749 13968 5783
rect 14002 5749 14041 5783
rect 14075 5749 14114 5783
rect 14148 5749 14187 5783
rect 14221 5749 14260 5783
rect 14294 5749 14333 5783
rect 14367 5749 14406 5783
rect 14440 5749 14479 5783
rect 14513 5749 14552 5783
rect 14586 5749 14625 5783
rect 14659 5749 14698 5783
rect 14732 5749 14771 5783
rect 14805 5749 14844 5783
rect 14878 5749 14917 5783
rect 14951 5749 14990 5783
rect 15024 5749 15063 5783
rect 15097 5749 15136 5783
rect 15170 5749 15209 5783
rect 15243 5749 15282 5783
rect 15316 5749 15355 5783
rect 15389 5749 15427 5783
rect 15461 5749 15499 5783
rect 15533 5749 15571 5783
rect 15605 5749 15643 5783
rect 15677 5749 15715 5783
rect 15749 5749 15787 5783
rect 15821 5749 15859 5783
rect 15893 5749 15931 5783
rect 15965 5749 16003 5783
rect 16037 5749 16075 5783
rect 16109 5749 16147 5783
rect 16181 5749 16219 5783
rect 16253 5749 16291 5783
rect 16325 5749 16337 5783
rect 13518 5743 16337 5749
rect 13518 5493 13730 5743
tri 13730 5718 13755 5743 nw
tri 16383 5637 16404 5658 se
rect 16404 5637 16543 6058
tri 16382 5636 16383 5637 se
rect 16383 5636 16543 5637
tri 14385 5633 14388 5636 se
rect 14388 5633 14451 5636
rect 13758 5627 14451 5633
rect 14503 5627 14515 5636
rect 13758 5593 13770 5627
rect 13804 5593 13844 5627
rect 13878 5593 13918 5627
rect 13952 5593 13992 5627
rect 14026 5593 14066 5627
rect 14100 5593 14140 5627
rect 14174 5593 14214 5627
rect 14248 5593 14288 5627
rect 14322 5593 14362 5627
rect 14396 5593 14436 5627
rect 14503 5593 14510 5627
rect 13758 5587 14451 5593
tri 14385 5584 14388 5587 ne
rect 14388 5584 14451 5587
rect 14503 5584 14515 5593
rect 14567 5584 14579 5636
rect 14631 5633 14637 5636
tri 14637 5633 14640 5636 sw
tri 16379 5633 16382 5636 se
rect 16382 5633 16543 5636
rect 14631 5627 16543 5633
rect 14631 5593 14658 5627
rect 14692 5593 14732 5627
rect 14766 5593 14806 5627
rect 14840 5593 14880 5627
rect 14914 5593 14954 5627
rect 14988 5593 15028 5627
rect 15062 5593 15102 5627
rect 15136 5593 15176 5627
rect 15210 5593 15250 5627
rect 15284 5593 15323 5627
rect 15357 5593 15396 5627
rect 15430 5593 15469 5627
rect 15503 5593 15542 5627
rect 15576 5593 15615 5627
rect 15649 5593 15688 5627
rect 15722 5593 15761 5627
rect 15795 5593 15834 5627
rect 15868 5593 15907 5627
rect 15941 5593 15980 5627
rect 16014 5593 16053 5627
rect 16087 5593 16126 5627
rect 16160 5593 16199 5627
rect 16233 5593 16272 5627
rect 16306 5593 16345 5627
rect 16379 5593 16418 5627
rect 16452 5593 16543 5627
rect 14631 5587 16543 5593
rect 14631 5584 14637 5587
tri 14637 5584 14640 5587 nw
tri 16379 5584 16382 5587 ne
rect 16382 5584 16543 5587
tri 16382 5565 16401 5584 ne
rect 16401 5565 16543 5584
tri 16401 5562 16404 5565 ne
tri 13730 5493 13739 5502 sw
rect 13518 5482 13739 5493
tri 13739 5482 13750 5493 sw
rect 13518 5477 13750 5482
tri 13750 5477 13755 5482 sw
rect 13518 5471 16337 5477
rect 13518 5437 13530 5471
rect 13564 5437 13603 5471
rect 13637 5437 13676 5471
rect 13710 5437 13749 5471
rect 13783 5437 13822 5471
rect 13856 5437 13895 5471
rect 13929 5437 13968 5471
rect 14002 5437 14041 5471
rect 14075 5437 14114 5471
rect 14148 5437 14187 5471
rect 14221 5437 14260 5471
rect 14294 5437 14333 5471
rect 14367 5437 14406 5471
rect 14440 5437 14479 5471
rect 14513 5437 14552 5471
rect 14586 5437 14625 5471
rect 14659 5437 14698 5471
rect 14732 5437 14771 5471
rect 14805 5437 14844 5471
rect 14878 5437 14917 5471
rect 14951 5437 14990 5471
rect 15024 5437 15063 5471
rect 15097 5437 15136 5471
rect 15170 5437 15209 5471
rect 15243 5437 15282 5471
rect 15316 5437 15355 5471
rect 15389 5437 15427 5471
rect 15461 5437 15499 5471
rect 15533 5437 15571 5471
rect 15605 5437 15643 5471
rect 15677 5437 15715 5471
rect 15749 5437 15787 5471
rect 15821 5437 15859 5471
rect 15893 5437 15931 5471
rect 15965 5437 16003 5471
rect 16037 5437 16075 5471
rect 16109 5437 16147 5471
rect 16181 5437 16219 5471
rect 16253 5437 16291 5471
rect 16325 5437 16337 5471
rect 13518 5431 16337 5437
rect 13518 5421 13745 5431
tri 13745 5421 13755 5431 nw
rect 13518 5410 13734 5421
tri 13734 5410 13745 5421 nw
rect 13518 5285 13730 5410
tri 13730 5406 13734 5410 nw
tri 13927 5383 13928 5384 se
rect 13928 5383 13976 5384
tri 13925 5381 13927 5383 se
rect 13927 5381 13976 5383
rect 13807 5375 13976 5381
rect 14028 5375 14040 5384
rect 13807 5341 13819 5375
rect 13853 5341 13892 5375
rect 13926 5341 13965 5375
rect 14028 5341 14038 5375
rect 13807 5335 13976 5341
tri 13925 5332 13928 5335 ne
rect 13928 5332 13976 5335
rect 14028 5332 14040 5341
rect 14092 5332 14104 5384
rect 14156 5383 14162 5384
tri 14162 5383 14163 5384 sw
rect 14156 5381 14163 5383
tri 14163 5381 14165 5383 sw
rect 14156 5375 16339 5381
rect 14156 5341 14184 5375
rect 14218 5341 14257 5375
rect 14291 5341 14330 5375
rect 14364 5341 14403 5375
rect 14437 5341 14476 5375
rect 14510 5341 14549 5375
rect 14583 5341 14622 5375
rect 14656 5341 14695 5375
rect 14729 5341 14768 5375
rect 14802 5341 14841 5375
rect 14875 5341 14914 5375
rect 14948 5341 14987 5375
rect 15021 5341 15060 5375
rect 15094 5341 15133 5375
rect 15167 5341 15206 5375
rect 15240 5341 15279 5375
rect 15313 5341 15352 5375
rect 15386 5341 15425 5375
rect 15459 5341 15498 5375
rect 15532 5341 15571 5375
rect 15605 5341 15644 5375
rect 15678 5341 15717 5375
rect 15751 5341 15789 5375
rect 15823 5341 15861 5375
rect 15895 5341 15933 5375
rect 15967 5341 16005 5375
rect 16039 5341 16077 5375
rect 16111 5341 16149 5375
rect 16183 5341 16221 5375
rect 16255 5341 16293 5375
rect 16327 5341 16339 5375
rect 14156 5335 16339 5341
rect 14156 5332 14162 5335
tri 14162 5332 14165 5335 nw
tri 13730 5285 13755 5310 sw
rect 13518 5279 16339 5285
rect 13518 5245 13530 5279
rect 13564 5245 13603 5279
rect 13637 5245 13676 5279
rect 13710 5245 13749 5279
rect 13783 5245 13822 5279
rect 13856 5245 13895 5279
rect 13929 5245 13968 5279
rect 14002 5245 14041 5279
rect 14075 5245 14114 5279
rect 14148 5245 14187 5279
rect 14221 5245 14260 5279
rect 14294 5245 14333 5279
rect 14367 5245 14406 5279
rect 14440 5245 14479 5279
rect 14513 5245 14552 5279
rect 14586 5245 14625 5279
rect 14659 5245 14698 5279
rect 14732 5245 14771 5279
rect 14805 5245 14844 5279
rect 14878 5245 14917 5279
rect 14951 5245 14990 5279
rect 15024 5245 15063 5279
rect 15097 5245 15136 5279
rect 15170 5245 15209 5279
rect 15243 5245 15282 5279
rect 15316 5245 15355 5279
rect 15389 5245 15428 5279
rect 15462 5245 15501 5279
rect 15535 5245 15573 5279
rect 15607 5245 15645 5279
rect 15679 5245 15717 5279
rect 15751 5245 15789 5279
rect 15823 5245 15861 5279
rect 15895 5245 15933 5279
rect 15967 5245 16005 5279
rect 16039 5245 16077 5279
rect 16111 5245 16149 5279
rect 16183 5245 16221 5279
rect 16255 5245 16293 5279
rect 16327 5245 16339 5279
rect 13518 5239 16339 5245
rect 13518 4988 13730 5239
tri 13730 5214 13755 5239 nw
tri 16383 5133 16404 5154 se
rect 16404 5133 16543 5565
tri 14384 5129 14388 5133 se
rect 14388 5129 14451 5133
rect 13758 5123 14451 5129
rect 14503 5123 14515 5133
rect 13758 5089 13770 5123
rect 13804 5089 13844 5123
rect 13878 5089 13918 5123
rect 13952 5089 13992 5123
rect 14026 5089 14066 5123
rect 14100 5089 14140 5123
rect 14174 5089 14214 5123
rect 14248 5089 14288 5123
rect 14322 5089 14362 5123
rect 14396 5089 14436 5123
rect 14503 5089 14510 5123
rect 13758 5083 14451 5089
tri 14386 5081 14388 5083 ne
rect 14388 5081 14451 5083
rect 14503 5081 14515 5089
rect 14567 5081 14579 5133
rect 14631 5129 14637 5133
tri 14637 5129 14641 5133 sw
tri 16379 5129 16383 5133 se
rect 16383 5129 16543 5133
rect 14631 5123 16543 5129
rect 14631 5089 14656 5123
rect 14690 5089 14729 5123
rect 14763 5089 14802 5123
rect 14836 5089 14875 5123
rect 14909 5089 14948 5123
rect 14982 5089 15021 5123
rect 15055 5089 15094 5123
rect 15128 5089 15167 5123
rect 15201 5089 15240 5123
rect 15274 5089 15313 5123
rect 15347 5089 15386 5123
rect 15420 5089 15459 5123
rect 15493 5089 15532 5123
rect 15566 5089 15605 5123
rect 15639 5089 15678 5123
rect 15712 5089 15751 5123
rect 15785 5089 15824 5123
rect 15858 5089 15897 5123
rect 15931 5089 15970 5123
rect 16004 5089 16043 5123
rect 16077 5089 16116 5123
rect 16150 5089 16189 5123
rect 16223 5089 16262 5123
rect 16296 5089 16335 5123
rect 16369 5089 16408 5123
rect 16442 5089 16543 5123
rect 14631 5083 16543 5089
rect 14631 5081 14637 5083
tri 14637 5081 14639 5083 nw
tri 16379 5081 16381 5083 ne
rect 16381 5081 16543 5083
tri 16381 5061 16401 5081 ne
rect 16401 5061 16543 5081
tri 16401 5058 16404 5061 ne
tri 13730 4988 13740 4998 sw
rect 13518 4978 13740 4988
tri 13740 4978 13750 4988 sw
rect 13518 4973 13750 4978
tri 13750 4973 13755 4978 sw
rect 13518 4967 16339 4973
rect 13518 4933 13530 4967
rect 13564 4933 13603 4967
rect 13637 4933 13676 4967
rect 13710 4933 13749 4967
rect 13783 4933 13822 4967
rect 13856 4933 13895 4967
rect 13929 4933 13968 4967
rect 14002 4933 14041 4967
rect 14075 4933 14114 4967
rect 14148 4933 14187 4967
rect 14221 4933 14260 4967
rect 14294 4933 14333 4967
rect 14367 4933 14406 4967
rect 14440 4933 14479 4967
rect 14513 4933 14552 4967
rect 14586 4933 14625 4967
rect 14659 4933 14698 4967
rect 14732 4933 14771 4967
rect 14805 4933 14844 4967
rect 14878 4933 14917 4967
rect 14951 4933 14990 4967
rect 15024 4933 15063 4967
rect 15097 4933 15136 4967
rect 15170 4933 15209 4967
rect 15243 4933 15282 4967
rect 15316 4933 15355 4967
rect 15389 4933 15428 4967
rect 15462 4933 15501 4967
rect 15535 4933 15573 4967
rect 15607 4933 15645 4967
rect 15679 4933 15717 4967
rect 15751 4933 15789 4967
rect 15823 4933 15861 4967
rect 15895 4933 15933 4967
rect 15967 4933 16005 4967
rect 16039 4933 16077 4967
rect 16111 4933 16149 4967
rect 16183 4933 16221 4967
rect 16255 4933 16293 4967
rect 16327 4933 16339 4967
rect 13518 4927 16339 4933
rect 13518 4915 13743 4927
tri 13743 4915 13755 4927 nw
rect 13518 4906 13734 4915
tri 13734 4906 13743 4915 nw
rect 13518 4902 13730 4906
tri 13730 4902 13734 4906 nw
tri 13925 4877 13928 4880 se
rect 13928 4877 13991 4880
rect 13807 4871 13991 4877
rect 14043 4871 14055 4880
rect 14107 4871 14119 4880
rect 14171 4877 14177 4880
tri 14177 4877 14180 4880 sw
rect 14171 4871 16339 4877
rect 13807 4837 13819 4871
rect 13853 4837 13892 4871
rect 13926 4837 13965 4871
rect 14107 4837 14111 4871
rect 14171 4837 14184 4871
rect 14218 4837 14257 4871
rect 14291 4837 14330 4871
rect 14364 4837 14403 4871
rect 14437 4837 14476 4871
rect 14510 4837 14549 4871
rect 14583 4837 14622 4871
rect 14656 4837 14695 4871
rect 14729 4837 14768 4871
rect 14802 4837 14841 4871
rect 14875 4837 14914 4871
rect 14948 4837 14987 4871
rect 15021 4837 15060 4871
rect 15094 4837 15133 4871
rect 15167 4837 15206 4871
rect 15240 4837 15279 4871
rect 15313 4837 15352 4871
rect 15386 4837 15425 4871
rect 15459 4837 15498 4871
rect 15532 4837 15571 4871
rect 15605 4837 15644 4871
rect 15678 4837 15717 4871
rect 15751 4837 15789 4871
rect 15823 4837 15861 4871
rect 15895 4837 15933 4871
rect 15967 4837 16005 4871
rect 16039 4837 16077 4871
rect 16111 4837 16149 4871
rect 16183 4837 16221 4871
rect 16255 4837 16293 4871
rect 16327 4837 16339 4871
rect 13807 4831 13991 4837
tri 13925 4828 13928 4831 ne
rect 13928 4828 13991 4831
rect 14043 4828 14055 4837
rect 14107 4828 14119 4837
rect 14171 4831 16339 4837
rect 14171 4828 14177 4831
tri 14177 4828 14180 4831 nw
rect 13444 4701 13450 4735
rect 13484 4701 13490 4735
rect 13326 4620 13332 4654
rect 13366 4620 13372 4654
rect 13326 4582 13372 4620
rect 13326 4548 13332 4582
rect 13366 4548 13372 4582
rect 13326 4510 13372 4548
rect 13326 4476 13332 4510
rect 13366 4476 13372 4510
rect 13326 4438 13372 4476
tri 13438 4669 13444 4675 se
rect 13444 4669 13490 4701
rect 13438 4659 13490 4669
rect 13438 4641 13450 4659
rect 13484 4641 13490 4659
rect 13438 4582 13490 4589
rect 13438 4577 13450 4582
rect 13484 4577 13490 4582
rect 13438 4513 13490 4525
rect 13438 4455 13490 4461
rect 13518 4803 13730 4806
tri 13730 4803 13733 4806 sw
rect 13518 4781 13733 4803
tri 13733 4781 13755 4803 sw
rect 13518 4775 16339 4781
rect 13518 4741 13530 4775
rect 13564 4741 13603 4775
rect 13637 4741 13676 4775
rect 13710 4741 13749 4775
rect 13783 4741 13822 4775
rect 13856 4741 13895 4775
rect 13929 4741 13968 4775
rect 14002 4741 14041 4775
rect 14075 4741 14114 4775
rect 14148 4741 14187 4775
rect 14221 4741 14260 4775
rect 14294 4741 14333 4775
rect 14367 4741 14406 4775
rect 14440 4741 14479 4775
rect 14513 4741 14552 4775
rect 14586 4741 14625 4775
rect 14659 4741 14698 4775
rect 14732 4741 14771 4775
rect 14805 4741 14844 4775
rect 14878 4741 14917 4775
rect 14951 4741 14990 4775
rect 15024 4741 15063 4775
rect 15097 4741 15136 4775
rect 15170 4741 15209 4775
rect 15243 4741 15282 4775
rect 15316 4741 15355 4775
rect 15389 4741 15428 4775
rect 15462 4741 15501 4775
rect 15535 4741 15573 4775
rect 15607 4741 15645 4775
rect 15679 4741 15717 4775
rect 15751 4741 15789 4775
rect 15823 4741 15861 4775
rect 15895 4741 15933 4775
rect 15967 4741 16005 4775
rect 16039 4741 16077 4775
rect 16111 4741 16149 4775
rect 16183 4741 16221 4775
rect 16255 4741 16293 4775
rect 16327 4741 16339 4775
rect 13518 4735 16339 4741
rect 13518 4730 13750 4735
tri 13750 4730 13755 4735 nw
rect 13518 4477 13730 4730
tri 13730 4710 13750 4730 nw
tri 16382 4628 16404 4650 se
rect 16404 4628 16543 5061
tri 14385 4625 14388 4628 se
rect 14388 4625 14451 4628
rect 13758 4619 14451 4625
rect 14503 4619 14515 4628
rect 13758 4585 13770 4619
rect 13804 4585 13844 4619
rect 13878 4585 13918 4619
rect 13952 4585 13992 4619
rect 14026 4585 14066 4619
rect 14100 4585 14140 4619
rect 14174 4585 14214 4619
rect 14248 4585 14288 4619
rect 14322 4585 14362 4619
rect 14396 4585 14435 4619
rect 14503 4585 14508 4619
rect 13758 4579 14451 4585
tri 14385 4576 14388 4579 ne
rect 14388 4576 14451 4579
rect 14503 4576 14515 4585
rect 14567 4576 14579 4628
rect 14631 4625 14637 4628
tri 14637 4625 14640 4628 sw
tri 16379 4625 16382 4628 se
rect 16382 4625 16543 4628
rect 14631 4619 16543 4625
rect 14631 4585 14654 4619
rect 14688 4585 14727 4619
rect 14761 4585 14800 4619
rect 14834 4585 14873 4619
rect 14907 4585 14946 4619
rect 14980 4585 15019 4619
rect 15053 4585 15092 4619
rect 15126 4585 15165 4619
rect 15199 4585 15238 4619
rect 15272 4585 15311 4619
rect 15345 4585 15384 4619
rect 15418 4585 15457 4619
rect 15491 4585 15530 4619
rect 15564 4585 15603 4619
rect 15637 4585 15676 4619
rect 15710 4585 15749 4619
rect 15783 4585 15822 4619
rect 15856 4585 15895 4619
rect 15929 4585 15968 4619
rect 16002 4585 16041 4619
rect 16075 4585 16114 4619
rect 16148 4585 16187 4619
rect 16221 4585 16260 4619
rect 16294 4585 16333 4619
rect 16367 4585 16406 4619
rect 16440 4585 16543 4619
rect 14631 4579 16543 4585
rect 16644 6285 16650 6318
rect 16684 6285 16690 6319
rect 16644 6247 16690 6285
rect 16644 6213 16650 6247
rect 16684 6213 16690 6247
rect 16644 6175 16690 6213
rect 16644 6141 16650 6175
rect 16684 6141 16690 6175
rect 16644 6103 16690 6141
rect 16644 6069 16650 6103
rect 16684 6069 16690 6103
rect 16644 6031 16690 6069
rect 16644 5997 16650 6031
rect 16684 5997 16690 6031
rect 16644 5959 16690 5997
rect 16644 5925 16650 5959
rect 16684 5925 16690 5959
rect 16644 5887 16690 5925
rect 16644 5853 16650 5887
rect 16684 5853 16690 5887
rect 16644 5815 16690 5853
rect 16644 5781 16650 5815
rect 16684 5781 16690 5815
rect 16644 5743 16690 5781
rect 16644 5709 16650 5743
rect 16684 5709 16690 5743
rect 16644 5671 16690 5709
rect 16644 5637 16650 5671
rect 16684 5637 16690 5671
rect 16644 5599 16690 5637
rect 16644 5565 16650 5599
rect 16684 5565 16690 5599
rect 16644 5527 16690 5565
rect 16644 5493 16650 5527
rect 16684 5493 16690 5527
rect 16644 5455 16690 5493
rect 16644 5421 16650 5455
rect 16684 5421 16690 5455
rect 16644 5383 16690 5421
rect 16644 5349 16650 5383
rect 16684 5349 16690 5383
rect 16644 5311 16690 5349
rect 16644 5277 16650 5311
rect 16684 5277 16690 5311
rect 16644 5239 16690 5277
rect 16644 5205 16650 5239
rect 16684 5205 16690 5239
rect 16644 5167 16690 5205
rect 16644 5133 16650 5167
rect 16684 5133 16690 5167
rect 16644 5095 16690 5133
rect 16644 5061 16650 5095
rect 16684 5061 16690 5095
rect 16644 5022 16690 5061
rect 16644 4988 16650 5022
rect 16684 4988 16690 5022
rect 16644 4949 16690 4988
rect 16644 4915 16650 4949
rect 16684 4915 16690 4949
rect 16644 4876 16690 4915
rect 16644 4842 16650 4876
rect 16684 4842 16690 4876
rect 16644 4803 16690 4842
rect 16644 4769 16650 4803
rect 16684 4769 16690 4803
rect 16644 4730 16690 4769
rect 16644 4696 16650 4730
rect 16684 4696 16690 4730
rect 16644 4657 16690 4696
rect 16644 4623 16650 4657
rect 16684 4623 16690 4657
rect 16644 4584 16690 4623
rect 14631 4576 14637 4579
tri 14637 4576 14640 4579 nw
rect 16644 4550 16650 4584
rect 16684 4550 16690 4584
rect 16644 4511 16690 4550
tri 13730 4477 13747 4494 sw
rect 16644 4477 16650 4511
rect 16684 4477 16690 4511
rect 13518 4474 13747 4477
tri 13747 4474 13750 4477 sw
rect 13518 4469 13750 4474
tri 13750 4469 13755 4474 sw
rect 13518 4463 16340 4469
rect 13326 4404 13332 4438
rect 13366 4404 13372 4438
rect 13518 4429 13530 4463
rect 13564 4429 13603 4463
rect 13637 4429 13676 4463
rect 13710 4429 13749 4463
rect 13783 4429 13822 4463
rect 13856 4429 13895 4463
rect 13929 4429 13968 4463
rect 14002 4429 14041 4463
rect 14075 4429 14114 4463
rect 14148 4429 14187 4463
rect 14221 4429 14260 4463
rect 14294 4429 14333 4463
rect 14367 4429 14406 4463
rect 14440 4429 14479 4463
rect 14513 4429 14552 4463
rect 14586 4429 14625 4463
rect 14659 4429 14698 4463
rect 14732 4429 14771 4463
rect 14805 4429 14844 4463
rect 14878 4429 14917 4463
rect 14951 4429 14990 4463
rect 15024 4429 15063 4463
rect 15097 4429 15136 4463
rect 15170 4429 15209 4463
rect 15243 4429 15282 4463
rect 15316 4429 15355 4463
rect 15389 4429 15428 4463
rect 15462 4429 15501 4463
rect 15535 4429 15574 4463
rect 15608 4429 15646 4463
rect 15680 4429 15718 4463
rect 15752 4429 15790 4463
rect 15824 4429 15862 4463
rect 15896 4429 15934 4463
rect 15968 4429 16006 4463
rect 16040 4429 16078 4463
rect 16112 4429 16150 4463
rect 16184 4429 16222 4463
rect 16256 4429 16294 4463
rect 16328 4429 16340 4463
rect 13518 4423 16340 4429
rect 16644 4438 16690 4477
tri 13372 4404 13374 4406 sw
tri 16642 4404 16644 4406 se
rect 16644 4404 16650 4438
rect 16684 4404 16690 4438
rect 13326 4402 13374 4404
tri 13374 4402 13376 4404 sw
tri 16640 4402 16642 4404 se
rect 16642 4402 16690 4404
rect 13326 4375 13376 4402
tri 13376 4375 13403 4402 sw
tri 16613 4375 16640 4402 se
rect 16640 4375 16690 4402
rect 13326 4372 13403 4375
tri 13403 4372 13406 4375 sw
tri 13925 4372 13928 4375 se
rect 13928 4372 13991 4375
rect 13326 4366 13991 4372
rect 14043 4366 14055 4375
rect 14107 4366 14119 4375
rect 14171 4372 14177 4375
tri 14177 4372 14180 4375 sw
tri 16610 4372 16613 4375 se
rect 16613 4372 16690 4375
rect 14171 4366 16690 4372
rect 13326 4332 13356 4366
rect 13390 4332 13439 4366
rect 13473 4332 13512 4366
rect 13546 4332 13585 4366
rect 13619 4332 13658 4366
rect 13692 4332 13731 4366
rect 13765 4332 13804 4366
rect 13838 4332 13877 4366
rect 13911 4332 13950 4366
rect 13984 4332 13991 4366
rect 14203 4332 14242 4366
rect 14276 4332 14315 4366
rect 14349 4332 14388 4366
rect 14422 4332 14461 4366
rect 14495 4332 14534 4366
rect 14568 4332 14607 4366
rect 14641 4332 14680 4366
rect 14714 4332 14753 4366
rect 14787 4332 14826 4366
rect 14860 4332 14899 4366
rect 14933 4332 14972 4366
rect 15006 4332 15045 4366
rect 15079 4332 15118 4366
rect 15152 4332 15191 4366
rect 15225 4332 15264 4366
rect 15298 4332 15337 4366
rect 15371 4332 15410 4366
rect 15444 4332 15483 4366
rect 15517 4332 15556 4366
rect 15590 4332 15629 4366
rect 15663 4332 15702 4366
rect 15736 4332 15775 4366
rect 15809 4332 15848 4366
rect 15882 4332 15921 4366
rect 15955 4332 15994 4366
rect 16028 4332 16067 4366
rect 16101 4332 16140 4366
rect 16174 4332 16213 4366
rect 16247 4332 16286 4366
rect 16320 4332 16359 4366
rect 16393 4332 16432 4366
rect 16466 4332 16505 4366
rect 16539 4332 16578 4366
rect 16612 4332 16690 4366
rect 13326 4326 13991 4332
tri 13925 4323 13928 4326 ne
rect 13928 4323 13991 4326
rect 14043 4323 14055 4332
rect 14107 4323 14119 4332
rect 14171 4326 16690 4332
rect 16831 6384 16837 6418
rect 16871 6384 16951 6418
rect 16985 6384 16991 6418
rect 16831 6346 16991 6384
rect 16831 6312 16837 6346
rect 16871 6312 16951 6346
rect 16985 6312 16991 6346
rect 16831 6274 16991 6312
rect 16831 6240 16837 6274
rect 16871 6240 16951 6274
rect 16985 6240 16991 6274
rect 16831 6202 16991 6240
rect 16831 6168 16837 6202
rect 16871 6168 16951 6202
rect 16985 6168 16991 6202
rect 16831 6130 16991 6168
rect 16831 6096 16837 6130
rect 16871 6096 16951 6130
rect 16985 6096 16991 6130
rect 16831 6058 16991 6096
rect 16831 6024 16837 6058
rect 16871 6024 16951 6058
rect 16985 6024 16991 6058
rect 16831 5986 16991 6024
rect 16831 5952 16837 5986
rect 16871 5952 16951 5986
rect 16985 5952 16991 5986
rect 16831 5914 16991 5952
rect 16831 5880 16837 5914
rect 16871 5880 16951 5914
rect 16985 5880 16991 5914
rect 16831 5842 16991 5880
rect 16831 5808 16837 5842
rect 16871 5808 16951 5842
rect 16985 5808 16991 5842
rect 16831 5770 16991 5808
rect 16831 5736 16837 5770
rect 16871 5736 16951 5770
rect 16985 5736 16991 5770
rect 16831 5698 16991 5736
rect 16831 5664 16837 5698
rect 16871 5664 16951 5698
rect 16985 5664 16991 5698
rect 16831 5626 16991 5664
rect 16831 5592 16837 5626
rect 16871 5592 16951 5626
rect 16985 5592 16991 5626
rect 16831 5554 16991 5592
rect 16831 5520 16837 5554
rect 16871 5520 16951 5554
rect 16985 5520 16991 5554
rect 16831 5482 16991 5520
rect 16831 5448 16837 5482
rect 16871 5448 16951 5482
rect 16985 5448 16991 5482
rect 16831 5410 16991 5448
rect 16831 5376 16837 5410
rect 16871 5376 16951 5410
rect 16985 5376 16991 5410
rect 16831 5338 16991 5376
rect 16831 5304 16837 5338
rect 16871 5304 16951 5338
rect 16985 5304 16991 5338
rect 16831 5266 16991 5304
rect 16831 5232 16837 5266
rect 16871 5232 16951 5266
rect 16985 5232 16991 5266
rect 16831 5194 16991 5232
rect 16831 5160 16837 5194
rect 16871 5160 16951 5194
rect 16985 5160 16991 5194
rect 16831 5122 16991 5160
rect 16831 5088 16837 5122
rect 16871 5088 16951 5122
rect 16985 5088 16991 5122
rect 16831 5050 16991 5088
rect 16831 5016 16837 5050
rect 16871 5016 16951 5050
rect 16985 5016 16991 5050
rect 16831 4978 16991 5016
rect 16831 4944 16837 4978
rect 16871 4944 16951 4978
rect 16985 4944 16991 4978
rect 16831 4906 16991 4944
rect 16831 4872 16837 4906
rect 16871 4872 16951 4906
rect 16985 4872 16991 4906
rect 16831 4834 16991 4872
rect 16831 4800 16837 4834
rect 16871 4800 16951 4834
rect 16985 4800 16991 4834
rect 16831 4762 16991 4800
rect 16831 4728 16837 4762
rect 16871 4728 16951 4762
rect 16985 4728 16991 4762
rect 16831 4690 16991 4728
rect 16831 4656 16837 4690
rect 16871 4656 16951 4690
rect 16985 4656 16991 4690
rect 16831 4618 16991 4656
rect 16831 4584 16837 4618
rect 16871 4584 16951 4618
rect 16985 4584 16991 4618
rect 16831 4546 16991 4584
rect 16831 4512 16837 4546
rect 16871 4512 16951 4546
rect 16985 4512 16991 4546
rect 16831 4474 16991 4512
rect 16831 4440 16837 4474
rect 16871 4440 16951 4474
rect 16985 4440 16991 4474
rect 16831 4402 16991 4440
rect 16831 4368 16837 4402
rect 16871 4368 16951 4402
rect 16985 4368 16991 4402
rect 16831 4330 16991 4368
rect 14171 4323 14177 4326
tri 14177 4323 14180 4326 nw
rect 13026 4257 13186 4296
rect 16831 4296 16837 4330
rect 16871 4296 16951 4330
rect 16985 4296 16991 4330
tri 13186 4257 13195 4266 sw
rect 16831 4257 16991 4296
rect 13026 4223 13032 4257
rect 13066 4223 13146 4257
rect 13180 4223 13195 4257
tri 13195 4223 13229 4257 sw
rect 16831 4223 16837 4257
rect 16871 4223 16951 4257
rect 16985 4223 16991 4257
rect 13026 4194 13229 4223
tri 13229 4194 13258 4223 sw
tri 16803 4194 16831 4222 se
rect 16831 4194 16991 4223
rect 13026 4174 13258 4194
tri 13258 4174 13278 4194 sw
tri 16783 4174 16803 4194 se
rect 16803 4174 16991 4194
rect 13026 4168 16991 4174
rect 13026 4134 13038 4168
rect 13072 4134 13111 4168
rect 13145 4134 13184 4168
rect 13218 4134 13257 4168
rect 13291 4134 13330 4168
rect 13364 4134 13403 4168
rect 13437 4134 13476 4168
rect 13510 4134 13549 4168
rect 13583 4134 13622 4168
rect 13656 4134 13695 4168
rect 13729 4134 13768 4168
rect 13802 4134 13841 4168
rect 13875 4134 13914 4168
rect 13948 4134 13987 4168
rect 14021 4134 14060 4168
rect 14094 4134 14133 4168
rect 14167 4134 14206 4168
rect 14240 4134 14279 4168
rect 14313 4134 14352 4168
rect 14386 4134 14425 4168
rect 14459 4134 14497 4168
rect 14531 4134 14569 4168
rect 14603 4134 14641 4168
rect 14675 4134 14713 4168
rect 14747 4134 14785 4168
rect 14819 4134 14857 4168
rect 14891 4134 14929 4168
rect 14963 4134 15001 4168
rect 15035 4134 15073 4168
rect 15107 4134 15145 4168
rect 15179 4134 15217 4168
rect 15251 4134 15289 4168
rect 15323 4134 15361 4168
rect 15395 4134 15433 4168
rect 15467 4134 15505 4168
rect 15539 4134 15577 4168
rect 15611 4134 15649 4168
rect 15683 4134 15721 4168
rect 15755 4134 15793 4168
rect 15827 4134 15865 4168
rect 15899 4134 15937 4168
rect 15971 4134 16009 4168
rect 16043 4134 16081 4168
rect 16115 4134 16153 4168
rect 16187 4134 16225 4168
rect 16259 4134 16297 4168
rect 16331 4134 16369 4168
rect 16403 4134 16441 4168
rect 16475 4134 16513 4168
rect 16547 4134 16585 4168
rect 16619 4134 16657 4168
rect 16691 4134 16729 4168
rect 16763 4134 16801 4168
rect 16835 4134 16873 4168
rect 16907 4134 16945 4168
rect 16979 4134 16991 4168
rect 13026 4054 16991 4134
rect 13026 4020 13038 4054
rect 13072 4020 13111 4054
rect 13145 4020 13184 4054
rect 13218 4020 13257 4054
rect 13291 4020 13330 4054
rect 13364 4020 13403 4054
rect 13437 4020 13476 4054
rect 13510 4020 13549 4054
rect 13583 4020 13622 4054
rect 13656 4020 13695 4054
rect 13729 4020 13768 4054
rect 13802 4020 13841 4054
rect 13875 4020 13914 4054
rect 13948 4020 13987 4054
rect 14021 4020 14060 4054
rect 14094 4020 14133 4054
rect 14167 4020 14206 4054
rect 14240 4020 14279 4054
rect 14313 4020 14352 4054
rect 14386 4020 14425 4054
rect 14459 4020 14497 4054
rect 14531 4020 14569 4054
rect 14603 4020 14641 4054
rect 14675 4020 14713 4054
rect 14747 4020 14785 4054
rect 14819 4020 14857 4054
rect 14891 4020 14929 4054
rect 14963 4020 15001 4054
rect 15035 4020 15073 4054
rect 15107 4020 15145 4054
rect 15179 4020 15217 4054
rect 15251 4020 15289 4054
rect 15323 4020 15361 4054
rect 15395 4020 15433 4054
rect 15467 4020 15505 4054
rect 15539 4020 15577 4054
rect 15611 4020 15649 4054
rect 15683 4020 15721 4054
rect 15755 4020 15793 4054
rect 15827 4020 15865 4054
rect 15899 4020 15937 4054
rect 15971 4020 16009 4054
rect 16043 4020 16081 4054
rect 16115 4020 16153 4054
rect 16187 4020 16225 4054
rect 16259 4020 16297 4054
rect 16331 4020 16369 4054
rect 16403 4020 16441 4054
rect 16475 4020 16513 4054
rect 16547 4020 16585 4054
rect 16619 4020 16657 4054
rect 16691 4020 16729 4054
rect 16763 4020 16801 4054
rect 16835 4020 16873 4054
rect 16907 4020 16945 4054
rect 16979 4020 16991 4054
rect 13026 4014 16991 4020
rect 17212 6677 17384 6716
rect 17212 6643 17218 6677
rect 17252 6643 17344 6677
rect 17378 6643 17384 6677
rect 17212 6604 17384 6643
rect 17212 6570 17218 6604
rect 17252 6570 17344 6604
rect 17378 6570 17384 6604
rect 17212 6531 17384 6570
rect 17212 6497 17218 6531
rect 17252 6497 17344 6531
rect 17378 6497 17384 6531
rect 17212 6458 17384 6497
rect 17212 6424 17218 6458
rect 17252 6424 17344 6458
rect 17378 6424 17384 6458
rect 17212 6385 17384 6424
rect 17212 6351 17218 6385
rect 17252 6351 17344 6385
rect 17378 6351 17384 6385
rect 17212 6312 17384 6351
rect 17212 6278 17218 6312
rect 17252 6278 17344 6312
rect 17378 6278 17384 6312
rect 17212 6239 17384 6278
rect 17212 6205 17218 6239
rect 17252 6205 17344 6239
rect 17378 6205 17384 6239
rect 17212 6166 17384 6205
rect 17212 6132 17218 6166
rect 17252 6132 17344 6166
rect 17378 6132 17384 6166
rect 17212 6093 17384 6132
rect 17212 6059 17218 6093
rect 17252 6059 17344 6093
rect 17378 6059 17384 6093
rect 17212 6020 17384 6059
rect 17212 5986 17218 6020
rect 17252 5986 17344 6020
rect 17378 5986 17384 6020
rect 17212 5947 17384 5986
rect 17212 5913 17218 5947
rect 17252 5913 17344 5947
rect 17378 5913 17384 5947
rect 17212 5874 17384 5913
rect 17212 5840 17218 5874
rect 17252 5840 17344 5874
rect 17378 5840 17384 5874
rect 17212 5801 17384 5840
rect 17212 5767 17218 5801
rect 17252 5767 17344 5801
rect 17378 5767 17384 5801
rect 17212 5728 17384 5767
rect 17212 5694 17218 5728
rect 17252 5694 17344 5728
rect 17378 5694 17384 5728
rect 17212 5655 17384 5694
rect 17212 5621 17218 5655
rect 17252 5621 17344 5655
rect 17378 5621 17384 5655
rect 17212 5582 17384 5621
rect 17212 5548 17218 5582
rect 17252 5548 17344 5582
rect 17378 5548 17384 5582
rect 17212 5509 17384 5548
rect 17212 5475 17218 5509
rect 17252 5475 17344 5509
rect 17378 5475 17384 5509
rect 17212 5436 17384 5475
rect 17212 5402 17218 5436
rect 17252 5402 17344 5436
rect 17378 5402 17384 5436
rect 17212 5363 17384 5402
rect 17212 5329 17218 5363
rect 17252 5329 17344 5363
rect 17378 5329 17384 5363
rect 17212 5290 17384 5329
rect 17212 5256 17218 5290
rect 17252 5256 17344 5290
rect 17378 5256 17384 5290
rect 17212 5217 17384 5256
rect 17212 5183 17218 5217
rect 17252 5183 17344 5217
rect 17378 5183 17384 5217
rect 17212 5144 17384 5183
rect 17212 5110 17218 5144
rect 17252 5110 17344 5144
rect 17378 5110 17384 5144
rect 17212 5071 17384 5110
rect 17212 5037 17218 5071
rect 17252 5037 17344 5071
rect 17378 5037 17384 5071
rect 17212 4998 17384 5037
rect 17212 4964 17218 4998
rect 17252 4964 17344 4998
rect 17378 4964 17384 4998
rect 17212 4925 17384 4964
rect 17212 4891 17218 4925
rect 17252 4891 17344 4925
rect 17378 4891 17384 4925
rect 17212 4852 17384 4891
rect 17212 4818 17218 4852
rect 17252 4818 17344 4852
rect 17378 4818 17384 4852
rect 17212 4779 17384 4818
rect 17212 4745 17218 4779
rect 17252 4745 17344 4779
rect 17378 4745 17384 4779
rect 17212 4706 17384 4745
rect 17212 4672 17218 4706
rect 17252 4672 17344 4706
rect 17378 4672 17384 4706
rect 17212 4633 17384 4672
rect 17212 4599 17218 4633
rect 17252 4599 17344 4633
rect 17378 4599 17384 4633
rect 17212 4560 17384 4599
rect 17212 4526 17218 4560
rect 17252 4526 17344 4560
rect 17378 4526 17384 4560
rect 17212 4487 17384 4526
rect 17212 4453 17218 4487
rect 17252 4453 17344 4487
rect 17378 4453 17384 4487
rect 17212 4414 17384 4453
rect 17212 4380 17218 4414
rect 17252 4380 17344 4414
rect 17378 4380 17384 4414
rect 17212 4341 17384 4380
rect 17212 4307 17218 4341
rect 17252 4307 17344 4341
rect 17378 4307 17384 4341
rect 17212 4268 17384 4307
rect 17212 4234 17218 4268
rect 17252 4234 17344 4268
rect 17378 4234 17384 4268
rect 17212 4194 17384 4234
rect 17212 4160 17218 4194
rect 17252 4160 17344 4194
rect 17378 4160 17384 4194
rect 17212 4120 17384 4160
rect 17212 4086 17218 4120
rect 17252 4086 17344 4120
rect 17378 4086 17384 4120
rect 17212 4046 17384 4086
rect 12628 3944 12800 3984
rect 17212 4012 17218 4046
rect 17252 4012 17344 4046
rect 17378 4012 17384 4046
rect 17212 3972 17384 4012
rect 4229 3847 4235 3881
rect 4269 3847 4275 3881
rect 11186 3911 12470 3916
rect 11186 3859 11195 3911
rect 11247 3859 11266 3911
rect 11318 3859 11336 3911
rect 11388 3859 12339 3911
rect 12391 3859 12412 3911
rect 12464 3859 12470 3911
rect 11186 3854 12470 3859
rect 12628 3910 12634 3944
rect 12668 3910 12760 3944
rect 12794 3910 12800 3944
rect 12628 3870 12800 3910
rect 4229 3804 4275 3847
rect 12628 3836 12634 3870
rect 12668 3836 12760 3870
rect 12794 3836 12800 3870
rect 13928 3907 13934 3959
rect 13986 3907 13999 3959
rect 13928 3895 13999 3907
rect 13928 3843 13934 3895
rect 13986 3843 13999 3895
rect 14179 3843 14185 3959
rect 14388 3913 14394 3965
rect 14446 3913 14487 3965
rect 14539 3913 14579 3965
rect 14631 3913 14637 3965
rect 14388 3901 14637 3913
rect 14388 3849 14394 3901
rect 14446 3849 14487 3901
rect 14539 3849 14579 3901
rect 14631 3849 14637 3901
rect 17212 3938 17218 3972
rect 17252 3938 17344 3972
rect 17378 3938 17384 3972
rect 17212 3898 17384 3938
rect 17212 3864 17218 3898
rect 17252 3864 17344 3898
rect 17378 3864 17384 3898
rect 4229 3770 4235 3804
rect 4269 3770 4275 3804
tri 12600 3780 12628 3808 se
rect 12628 3780 12800 3836
tri 12594 3774 12600 3780 se
rect 12600 3774 12800 3780
tri 12800 3774 12834 3808 sw
tri 17178 3774 17212 3808 se
rect 17212 3780 17384 3864
tri 17384 3780 17412 3808 sw
rect 17212 3774 17412 3780
tri 17412 3774 17418 3780 sw
rect 4229 3727 4275 3770
rect 4229 3693 4235 3727
rect 4269 3693 4275 3727
rect 4229 3681 4275 3693
rect 14388 3722 14394 3774
rect 14446 3722 14487 3774
rect 14539 3722 14579 3774
rect 14631 3722 14637 3774
rect 14388 3710 14637 3722
rect 14388 3658 14394 3710
rect 14446 3658 14487 3710
rect 14539 3658 14579 3710
rect 14631 3658 14637 3710
rect 3416 3644 3701 3648
tri 3701 3644 3705 3648 sw
tri 3758 3644 3762 3648 se
rect 3762 3644 4173 3648
rect 3416 3441 3705 3644
rect 3707 3643 3743 3644
rect 3706 3442 3744 3643
rect 3707 3441 3743 3442
rect 3745 3441 4173 3644
tri 3164 3422 3183 3441 nw
rect 3416 3422 3686 3441
tri 3686 3422 3705 3441 nw
rect 2831 3256 2837 3308
rect 2889 3256 2895 3308
rect 2831 3244 2895 3256
rect 2831 3192 2837 3244
rect 2889 3192 2895 3244
rect 2831 3180 2895 3192
rect 2485 3127 2487 3156
rect 2831 3128 2837 3180
rect 2889 3128 2895 3180
rect 2831 3116 2895 3128
rect 2831 3064 2837 3116
rect 2889 3064 2895 3116
rect 2831 3058 2895 3064
rect 2080 3029 2132 3041
rect 2080 2965 2132 2977
rect 2080 2909 2092 2913
rect 2126 2909 2132 2913
rect 2080 2901 2132 2909
rect 2080 2837 2092 2849
rect 2126 2837 2132 2849
rect 2080 2799 2132 2837
rect 3416 2803 3614 3422
tri 3614 3350 3686 3422 nw
rect 2080 2765 2092 2799
rect 2126 2765 2132 2799
rect 2080 2727 2132 2765
rect 2080 2693 2092 2727
rect 2126 2693 2132 2727
rect 2080 2681 2132 2693
rect -104 262 68 845
tri 68 840 73 845 nw
tri 68 262 219 413 sw
rect -104 250 988 262
rect -104 216 186 250
rect 220 216 618 250
rect 652 216 988 250
rect -104 178 988 216
rect -104 144 186 178
rect 220 144 618 178
rect 652 144 988 178
rect -104 140 988 144
tri -104 106 -70 140 ne
rect -70 106 988 140
tri -70 72 -36 106 ne
rect -36 72 186 106
rect 220 72 618 106
rect 652 72 988 106
tri -36 60 -24 72 ne
rect -24 60 988 72
tri -24 0 36 60 ne
rect 36 0 988 60
<< rmetal1 >>
rect 3322 7118 3324 7119
rect 3360 7118 3362 7119
rect 3322 6860 3323 7118
rect 3361 6860 3362 7118
rect 3322 6859 3324 6860
rect 3360 6859 3362 6860
rect 3266 6743 3302 6744
rect 3266 6742 3267 6743
rect 3301 6742 3302 6743
rect 3266 6705 3267 6706
rect 3301 6705 3302 6706
rect 3266 6704 3302 6705
rect 3322 6588 3324 6589
rect 3360 6588 3362 6589
rect 3322 6544 3323 6588
rect 3361 6544 3362 6588
rect 3322 6543 3324 6544
rect 3360 6543 3362 6544
rect 2831 4752 2895 4753
rect 2831 4751 2832 4752
rect 2894 4751 2895 4752
rect 2831 4714 2832 4715
rect 2894 4714 2895 4715
rect 2831 4713 2895 4714
rect 2831 3680 2895 3681
rect 2831 3679 2832 3680
rect 2894 3679 2895 3680
rect 2831 3642 2832 3643
rect 2894 3642 2895 3643
rect 2831 3641 2895 3642
rect 3661 5045 3663 5046
rect 3661 4947 3662 5045
rect 3661 4946 3663 4947
rect 3699 5045 3701 5046
rect 3700 4947 3701 5045
rect 3699 4946 3701 4947
rect 4229 4759 4281 4760
rect 4229 4758 4230 4759
rect 4280 4758 4281 4759
rect 4229 4721 4230 4722
rect 4280 4721 4281 4722
rect 4229 4720 4281 4721
rect 4229 4388 4281 4389
rect 4229 4387 4230 4388
rect 4280 4387 4281 4388
rect 4229 4350 4230 4351
rect 4280 4350 4281 4351
rect 4229 4349 4281 4350
rect 3705 3643 3707 3644
rect 3743 3643 3745 3644
rect 3705 3442 3706 3643
rect 3744 3442 3745 3643
rect 3705 3441 3707 3442
rect 3743 3441 3745 3442
<< via1 >>
rect 154 7271 206 7323
rect 218 7271 270 7323
rect 282 7271 334 7323
rect 346 7271 398 7323
rect 343 6987 395 6998
rect 343 6953 349 6987
rect 349 6953 383 6987
rect 383 6953 395 6987
rect 343 6946 395 6953
rect 407 6987 459 6998
rect 407 6953 421 6987
rect 421 6953 455 6987
rect 455 6953 459 6987
rect 407 6946 459 6953
rect -40 6651 12 6703
rect -40 6587 12 6639
rect -40 6523 12 6575
rect -40 6459 12 6511
rect -40 6395 12 6447
rect -40 6331 12 6383
rect -40 6267 12 6319
rect 2837 7044 2889 7096
rect 2837 6980 2889 7032
rect 2837 6916 2889 6968
rect 2837 6852 2889 6904
rect 2837 6788 2889 6840
rect 1768 4999 1802 5031
rect 1802 4999 1820 5031
rect 1768 4979 1820 4999
rect 1768 4961 1820 4967
rect 1768 4927 1802 4961
rect 1802 4927 1820 4961
rect 1768 4915 1820 4927
rect 282 4874 334 4881
rect 282 4840 288 4874
rect 288 4840 322 4874
rect 322 4840 334 4874
rect 282 4829 334 4840
rect 282 4802 334 4817
rect 282 4768 288 4802
rect 288 4768 322 4802
rect 322 4768 334 4802
rect 282 4765 334 4768
rect 1221 4875 1273 4881
rect 1221 4841 1227 4875
rect 1227 4841 1261 4875
rect 1261 4841 1273 4875
rect 1851 4875 1903 4887
rect 1851 4841 1885 4875
rect 1885 4841 1903 4875
rect 1221 4829 1273 4841
rect 1221 4803 1273 4817
rect 1221 4769 1227 4803
rect 1227 4769 1261 4803
rect 1261 4769 1273 4803
rect 1221 4765 1273 4769
rect 1851 4835 1903 4841
rect 1851 4803 1903 4823
rect 1851 4771 1885 4803
rect 1885 4771 1903 4803
rect 2283 4634 2335 4686
rect 2347 4634 2399 4686
rect 1318 4598 1370 4610
rect 1318 4564 1324 4598
rect 1324 4564 1358 4598
rect 1358 4564 1370 4598
rect 1318 4558 1370 4564
rect 1382 4598 1434 4610
rect 1382 4564 1396 4598
rect 1396 4564 1430 4598
rect 1430 4564 1434 4598
rect 1382 4558 1434 4564
rect 2233 4465 2285 4517
rect 2297 4486 2315 4517
rect 2315 4486 2349 4517
rect 2297 4465 2349 4486
rect 2837 4979 2889 5031
rect 2837 4915 2889 4967
rect 3270 7057 3322 7109
rect 3270 6993 3322 7045
rect 3270 6929 3322 6981
rect 3270 6865 3322 6917
rect 12628 5921 12680 5930
rect 11263 5857 11315 5909
rect 11383 5857 11435 5909
rect 11263 5793 11315 5845
rect 11383 5793 11435 5845
rect 11263 5728 11315 5780
rect 11383 5728 11435 5780
rect 11263 5663 11315 5715
rect 11383 5663 11435 5715
rect 11263 5598 11315 5650
rect 11383 5598 11435 5650
rect 11263 5533 11315 5585
rect 11383 5533 11435 5585
rect 12628 5887 12634 5921
rect 12634 5887 12668 5921
rect 12668 5887 12680 5921
rect 12628 5878 12680 5887
rect 12748 5921 12800 5930
rect 12748 5887 12760 5921
rect 12760 5887 12794 5921
rect 12794 5887 12800 5921
rect 12748 5878 12800 5887
rect 12628 5848 12680 5859
rect 12628 5814 12634 5848
rect 12634 5814 12668 5848
rect 12668 5814 12680 5848
rect 12628 5807 12680 5814
rect 12748 5848 12800 5859
rect 12748 5814 12760 5848
rect 12760 5814 12794 5848
rect 12794 5814 12800 5848
rect 12748 5807 12800 5814
rect 12628 5775 12680 5787
rect 12628 5741 12634 5775
rect 12634 5741 12668 5775
rect 12668 5741 12680 5775
rect 12628 5735 12680 5741
rect 12748 5775 12800 5787
rect 12748 5741 12760 5775
rect 12760 5741 12794 5775
rect 12794 5741 12800 5775
rect 12748 5735 12800 5741
rect 2483 4175 2599 4355
rect 2837 4835 2889 4887
rect 2837 4771 2889 4823
rect 1582 3664 1634 3716
rect 1646 3664 1698 3716
rect 1894 3664 1946 3716
rect 1958 3664 2010 3716
rect 2971 4771 3151 4887
rect 1582 3628 1634 3634
rect 1582 3594 1588 3628
rect 1588 3594 1622 3628
rect 1622 3594 1634 3628
rect 1582 3582 1634 3594
rect 1646 3628 1698 3634
rect 1646 3594 1660 3628
rect 1660 3594 1694 3628
rect 1694 3594 1698 3628
rect 1646 3582 1698 3594
rect 1894 3628 1946 3634
rect 1894 3594 1900 3628
rect 1900 3594 1934 3628
rect 1934 3594 1946 3628
rect 1894 3582 1946 3594
rect 1958 3628 2010 3634
rect 1958 3594 1972 3628
rect 1972 3594 2006 3628
rect 2006 3594 2010 3628
rect 1958 3582 2010 3594
rect 1582 3500 1634 3552
rect 1646 3500 1698 3552
rect 1894 3500 1946 3552
rect 1958 3500 2010 3552
rect 1147 3302 1199 3354
rect 1147 3238 1199 3290
rect 1147 3174 1199 3226
rect 1147 3087 1199 3093
rect 1147 3053 1156 3087
rect 1156 3053 1190 3087
rect 1190 3053 1199 3087
rect 1147 3041 1199 3053
rect 1147 3015 1199 3029
rect 1147 2981 1156 3015
rect 1156 2981 1190 3015
rect 1190 2981 1199 3015
rect 1147 2977 1199 2981
rect 1147 2943 1199 2965
rect 1147 2913 1156 2943
rect 1156 2913 1190 2943
rect 1190 2913 1199 2943
rect 1147 2871 1199 2901
rect 1147 2849 1156 2871
rect 1156 2849 1190 2871
rect 1190 2849 1199 2871
rect 1459 3302 1511 3354
rect 1459 3238 1511 3290
rect 1459 3174 1511 3226
rect 1459 3087 1511 3093
rect 1459 3053 1468 3087
rect 1468 3053 1502 3087
rect 1502 3053 1511 3087
rect 1459 3041 1511 3053
rect 1459 3015 1511 3029
rect 1459 2981 1468 3015
rect 1468 2981 1502 3015
rect 1502 2981 1511 3015
rect 1459 2977 1511 2981
rect 1459 2943 1511 2965
rect 1459 2913 1468 2943
rect 1468 2913 1502 2943
rect 1502 2913 1511 2943
rect 1459 2871 1511 2901
rect 1459 2849 1468 2871
rect 1468 2849 1502 2871
rect 1502 2849 1511 2871
rect 1771 3302 1823 3354
rect 1771 3238 1823 3290
rect 1771 3174 1823 3226
rect 1771 3087 1823 3093
rect 1771 3053 1780 3087
rect 1780 3053 1814 3087
rect 1814 3053 1823 3087
rect 1771 3041 1823 3053
rect 1771 3015 1823 3029
rect 1771 2981 1780 3015
rect 1780 2981 1814 3015
rect 1814 2981 1823 3015
rect 1771 2977 1823 2981
rect 1771 2943 1823 2965
rect 1771 2913 1780 2943
rect 1780 2913 1814 2943
rect 1814 2913 1823 2943
rect 1771 2871 1823 2901
rect 1771 2849 1780 2871
rect 1780 2849 1814 2871
rect 1814 2849 1823 2871
rect 2080 3302 2132 3354
rect 2080 3238 2132 3290
rect 2080 3174 2132 3226
rect 4235 4835 4287 4887
rect 4235 4771 4287 4823
rect 4229 4459 4281 4511
rect 4229 4395 4281 4447
rect 11195 4393 11247 4445
rect 11266 4393 11318 4445
rect 11336 4393 11388 4445
rect 13976 6391 14028 6392
rect 13976 6357 13980 6391
rect 13980 6357 14014 6391
rect 14014 6357 14028 6391
rect 13976 6340 14028 6357
rect 14040 6391 14092 6392
rect 14040 6357 14052 6391
rect 14052 6357 14086 6391
rect 14086 6357 14092 6391
rect 14040 6340 14092 6357
rect 14104 6391 14156 6392
rect 14104 6357 14124 6391
rect 14124 6357 14156 6391
rect 14104 6340 14156 6357
rect 14451 6287 14503 6296
rect 14515 6287 14567 6296
rect 14579 6287 14631 6296
rect 14451 6253 14479 6287
rect 14479 6253 14503 6287
rect 14515 6253 14552 6287
rect 14552 6253 14567 6287
rect 14579 6253 14586 6287
rect 14586 6253 14625 6287
rect 14625 6253 14631 6287
rect 14451 6244 14503 6253
rect 14515 6244 14567 6253
rect 14579 6244 14631 6253
rect 14451 6131 14503 6141
rect 14515 6131 14567 6141
rect 14451 6097 14470 6131
rect 14470 6097 14503 6131
rect 14515 6097 14544 6131
rect 14544 6097 14567 6131
rect 14451 6089 14503 6097
rect 14515 6089 14567 6097
rect 14579 6131 14631 6141
rect 14579 6097 14584 6131
rect 14584 6097 14618 6131
rect 14618 6097 14631 6131
rect 14579 6089 14631 6097
rect 13991 5879 14043 5888
rect 14055 5879 14107 5888
rect 14119 5879 14171 5888
rect 13991 5845 13999 5879
rect 13999 5845 14038 5879
rect 14038 5845 14043 5879
rect 14055 5845 14072 5879
rect 14072 5845 14107 5879
rect 14119 5845 14145 5879
rect 14145 5845 14171 5879
rect 13991 5836 14043 5845
rect 14055 5836 14107 5845
rect 14119 5836 14171 5845
rect 14451 5627 14503 5636
rect 14515 5627 14567 5636
rect 14451 5593 14470 5627
rect 14470 5593 14503 5627
rect 14515 5593 14544 5627
rect 14544 5593 14567 5627
rect 14451 5584 14503 5593
rect 14515 5584 14567 5593
rect 14579 5627 14631 5636
rect 14579 5593 14584 5627
rect 14584 5593 14618 5627
rect 14618 5593 14631 5627
rect 14579 5584 14631 5593
rect 13976 5375 14028 5384
rect 14040 5375 14092 5384
rect 13976 5341 13999 5375
rect 13999 5341 14028 5375
rect 14040 5341 14072 5375
rect 14072 5341 14092 5375
rect 13976 5332 14028 5341
rect 14040 5332 14092 5341
rect 14104 5375 14156 5384
rect 14104 5341 14111 5375
rect 14111 5341 14145 5375
rect 14145 5341 14156 5375
rect 14104 5332 14156 5341
rect 14451 5123 14503 5133
rect 14515 5123 14567 5133
rect 14451 5089 14470 5123
rect 14470 5089 14503 5123
rect 14515 5089 14544 5123
rect 14544 5089 14567 5123
rect 14451 5081 14503 5089
rect 14515 5081 14567 5089
rect 14579 5123 14631 5133
rect 14579 5089 14583 5123
rect 14583 5089 14617 5123
rect 14617 5089 14631 5123
rect 14579 5081 14631 5089
rect 13991 4871 14043 4880
rect 14055 4871 14107 4880
rect 14119 4871 14171 4880
rect 13991 4837 13999 4871
rect 13999 4837 14038 4871
rect 14038 4837 14043 4871
rect 14055 4837 14072 4871
rect 14072 4837 14107 4871
rect 14119 4837 14145 4871
rect 14145 4837 14171 4871
rect 13991 4828 14043 4837
rect 14055 4828 14107 4837
rect 14119 4828 14171 4837
rect 13438 4625 13450 4641
rect 13450 4625 13484 4641
rect 13484 4625 13490 4641
rect 13438 4589 13490 4625
rect 13438 4548 13450 4577
rect 13450 4548 13484 4577
rect 13484 4548 13490 4577
rect 13438 4525 13490 4548
rect 13438 4505 13490 4513
rect 13438 4471 13450 4505
rect 13450 4471 13484 4505
rect 13484 4471 13490 4505
rect 13438 4461 13490 4471
rect 14451 4619 14503 4628
rect 14515 4619 14567 4628
rect 14451 4585 14469 4619
rect 14469 4585 14503 4619
rect 14515 4585 14542 4619
rect 14542 4585 14567 4619
rect 14451 4576 14503 4585
rect 14515 4576 14567 4585
rect 14579 4619 14631 4628
rect 14579 4585 14581 4619
rect 14581 4585 14615 4619
rect 14615 4585 14631 4619
rect 14579 4576 14631 4585
rect 13991 4366 14043 4375
rect 14055 4366 14107 4375
rect 14119 4366 14171 4375
rect 13991 4332 14023 4366
rect 14023 4332 14043 4366
rect 14055 4332 14057 4366
rect 14057 4332 14096 4366
rect 14096 4332 14107 4366
rect 14119 4332 14130 4366
rect 14130 4332 14169 4366
rect 14169 4332 14171 4366
rect 13991 4323 14043 4332
rect 14055 4323 14107 4332
rect 14119 4323 14171 4332
rect 11195 3859 11247 3911
rect 11266 3859 11318 3911
rect 11336 3859 11388 3911
rect 12339 3859 12391 3911
rect 12412 3859 12464 3911
rect 13934 3907 13986 3959
rect 13934 3843 13986 3895
rect 13999 3843 14179 3959
rect 14394 3913 14446 3965
rect 14487 3913 14539 3965
rect 14579 3913 14631 3965
rect 14394 3849 14446 3901
rect 14487 3849 14539 3901
rect 14579 3849 14631 3901
rect 14394 3722 14446 3774
rect 14487 3722 14539 3774
rect 14579 3722 14631 3774
rect 14394 3658 14446 3710
rect 14487 3658 14539 3710
rect 14579 3658 14631 3710
rect 2837 3256 2889 3308
rect 2837 3192 2889 3244
rect 2837 3128 2889 3180
rect 2080 3087 2132 3093
rect 2080 3053 2092 3087
rect 2092 3053 2126 3087
rect 2126 3053 2132 3087
rect 2837 3064 2889 3116
rect 2080 3041 2132 3053
rect 2080 3015 2132 3029
rect 2080 2981 2092 3015
rect 2092 2981 2126 3015
rect 2126 2981 2132 3015
rect 2080 2977 2132 2981
rect 2080 2943 2132 2965
rect 2080 2913 2092 2943
rect 2092 2913 2126 2943
rect 2126 2913 2132 2943
rect 2080 2871 2132 2901
rect 2080 2849 2092 2871
rect 2092 2849 2126 2871
rect 2126 2849 2132 2871
<< metal2 >>
rect 148 7271 154 7323
rect 206 7271 218 7323
rect 270 7271 282 7323
rect 334 7271 346 7323
rect 398 7271 747 7323
tri 747 7271 799 7323 sw
tri 148 7244 175 7271 ne
rect 175 7115 799 7271
tri 799 7115 955 7271 sw
rect 175 7109 955 7115
tri 955 7109 961 7115 sw
rect 3267 7109 3331 7115
rect 175 7102 961 7109
tri 961 7102 968 7109 sw
rect 2837 7096 2889 7102
rect 2837 7032 2889 7044
rect 337 6946 343 6998
rect 395 6946 407 6998
rect 459 6946 465 6998
rect 2837 6968 2889 6980
tri 465 6946 474 6955 sw
rect 337 6917 474 6946
tri 474 6917 503 6946 sw
rect 337 6916 503 6917
tri 503 6916 504 6917 sw
rect 337 6904 504 6916
tri 504 6904 516 6916 sw
rect 2837 6904 2889 6916
rect 337 6891 516 6904
tri 439 6852 478 6891 ne
rect 478 6852 516 6891
tri 516 6852 568 6904 sw
tri 478 6840 490 6852 ne
rect 490 6840 568 6852
tri 568 6840 580 6852 sw
rect 2837 6840 2889 6852
tri 490 6827 503 6840 ne
rect 503 6827 580 6840
tri 580 6827 593 6840 sw
tri 503 6788 542 6827 ne
rect 542 6788 593 6827
tri 593 6788 632 6827 sw
tri 542 6737 593 6788 ne
rect 593 6782 632 6788
tri 632 6782 638 6788 sw
rect 2837 6782 2889 6788
rect 3267 7057 3270 7109
rect 3322 7057 3331 7109
rect 3267 7045 3331 7057
rect 3267 6993 3270 7045
rect 3322 6993 3331 7045
rect 3267 6981 3331 6993
rect 3267 6929 3270 6981
rect 3322 6929 3331 6981
rect 3267 6917 3331 6929
rect 3267 6865 3270 6917
rect 3322 6865 3331 6917
tri 3266 6782 3267 6783 se
rect 3267 6782 3331 6865
rect 593 6737 638 6782
tri 638 6737 683 6782 sw
tri 3221 6737 3266 6782 se
rect 3266 6757 3331 6782
rect 3266 6737 3311 6757
tri 3311 6737 3331 6757 nw
tri 593 6709 621 6737 ne
rect 621 6709 3247 6737
rect -40 6703 12 6709
tri 621 6673 657 6709 ne
rect 657 6673 3247 6709
tri 3247 6673 3311 6737 nw
rect 13029 6668 13413 7271
rect -40 6639 12 6651
rect -40 6575 12 6587
rect -40 6511 12 6523
rect -40 6447 12 6459
rect -40 6383 12 6395
rect -40 6319 12 6331
rect -40 6261 12 6267
rect 13928 6392 14185 6407
rect 13928 6340 13976 6392
rect 14028 6340 14040 6392
rect 14092 6340 14104 6392
rect 14156 6340 14185 6392
rect 12628 5930 12800 5936
rect 11263 5909 11653 5915
rect 11315 5857 11383 5909
rect 11435 5878 11653 5909
tri 11653 5878 11690 5915 sw
rect 12680 5878 12748 5930
rect 11435 5859 11690 5878
tri 11690 5859 11709 5878 sw
rect 12628 5859 12800 5878
rect 13928 5888 14185 6340
rect 14388 6244 14451 6296
rect 14503 6244 14515 6296
rect 14567 6244 14579 6296
rect 14631 6244 14637 6296
rect 11435 5857 11709 5859
rect 11263 5845 11709 5857
rect 11315 5793 11383 5845
rect 11435 5807 11709 5845
tri 11709 5807 11761 5859 sw
rect 12680 5807 12748 5859
tri 13904 5836 13928 5860 se
rect 13928 5836 13991 5888
rect 14043 5836 14055 5888
rect 14107 5836 14119 5888
rect 14171 5836 14185 5888
rect 11435 5793 11761 5807
rect 11263 5787 11761 5793
tri 11761 5787 11781 5807 sw
rect 12628 5787 12800 5807
rect 11263 5780 11781 5787
rect 11315 5728 11383 5780
rect 11435 5735 11781 5780
tri 11781 5735 11833 5787 sw
rect 12680 5735 12748 5787
rect 11435 5729 11833 5735
tri 11833 5729 11839 5735 sw
rect 12628 5729 12800 5735
tri 13797 5729 13904 5836 se
rect 13904 5729 14185 5836
rect 11435 5728 11839 5729
rect 11263 5715 11839 5728
rect 11315 5663 11383 5715
rect 11435 5689 11839 5715
tri 11839 5689 11879 5729 sw
tri 13757 5689 13797 5729 se
rect 13797 5689 14185 5729
rect 11435 5663 14185 5689
rect 11263 5650 14185 5663
rect 11315 5598 11383 5650
rect 11435 5598 14185 5650
rect 11263 5585 14185 5598
rect 11315 5533 11383 5585
rect 11435 5533 14185 5585
rect 11263 5527 14185 5533
tri 11537 5384 11680 5527 ne
rect 11680 5384 14185 5527
tri 11680 5332 11732 5384 ne
rect 11732 5332 13976 5384
rect 14028 5332 14040 5384
rect 14092 5332 14104 5384
rect 14156 5332 14185 5384
tri 11732 5253 11811 5332 ne
rect 11811 5253 14185 5332
tri 13752 5133 13872 5253 ne
rect 13872 5133 14185 5253
tri 13872 5081 13924 5133 ne
rect 13924 5081 14185 5133
tri 13924 5077 13928 5081 ne
rect 1762 4979 1768 5031
rect 1820 4979 2837 5031
rect 2889 4979 2895 5031
rect 1762 4967 2895 4979
rect 1762 4915 1768 4967
rect 1820 4915 2837 4967
rect 2889 4915 2895 4967
rect 282 4881 334 4887
tri 334 4881 339 4886 sw
tri 1216 4881 1221 4886 se
rect 1221 4881 1273 4887
rect 334 4852 339 4881
tri 339 4852 368 4881 sw
tri 1187 4852 1216 4881 se
rect 1216 4852 1221 4881
rect 334 4829 1221 4852
tri 1273 4852 1308 4887 sw
tri 1810 4852 1845 4887 se
rect 1845 4852 1851 4887
rect 1273 4835 1851 4852
rect 1903 4835 2837 4887
rect 2889 4835 2895 4887
rect 1273 4829 2895 4835
rect 282 4823 2895 4829
rect 282 4817 1851 4823
rect 334 4797 1221 4817
rect 334 4765 336 4797
tri 336 4765 368 4797 nw
tri 1187 4765 1219 4797 ne
rect 1219 4765 1221 4797
rect 1273 4797 1851 4817
rect 1273 4771 1285 4797
tri 1285 4771 1311 4797 nw
tri 1811 4771 1837 4797 ne
rect 1837 4771 1851 4797
rect 1903 4771 2837 4823
rect 2889 4771 2895 4823
rect 2962 4771 2971 4887
rect 3151 4835 4235 4887
rect 4287 4835 4293 4887
rect 3151 4823 4293 4835
tri 13515 4828 13524 4837 se
rect 13524 4828 13716 4902
rect 3151 4771 4235 4823
rect 4287 4771 4293 4823
tri 13490 4803 13515 4828 se
rect 13515 4803 13716 4828
rect 13928 4880 14185 5081
rect 13928 4828 13991 4880
rect 14043 4828 14055 4880
rect 14107 4828 14119 4880
rect 14171 4828 14185 4880
rect 1273 4768 1282 4771
tri 1282 4768 1285 4771 nw
tri 1837 4768 1840 4771 ne
rect 1840 4768 1940 4771
tri 1940 4768 1943 4771 nw
tri 2797 4768 2800 4771 ne
rect 2800 4768 2895 4771
rect 282 4759 334 4765
tri 334 4763 336 4765 nw
tri 1219 4763 1221 4765 ne
rect 1221 4759 1273 4765
tri 1273 4759 1282 4768 nw
tri 1840 4763 1845 4768 ne
rect 1845 4763 1935 4768
tri 1935 4763 1940 4768 nw
tri 2800 4763 2805 4768 ne
rect 2805 4763 2895 4768
rect 1845 4759 1931 4763
tri 1931 4759 1935 4763 nw
tri 2805 4759 2809 4763 ne
rect 2809 4759 2895 4763
tri 2895 4759 2904 4768 sw
tri 1820 4634 1845 4659 se
rect 1845 4634 1909 4759
tri 1909 4737 1931 4759 nw
tri 2809 4737 2831 4759 ne
rect 2831 4737 2904 4759
tri 2831 4725 2843 4737 ne
rect 2843 4725 2904 4737
tri 2904 4725 2938 4759 sw
rect 12208 4741 13524 4803
rect 12208 4725 12326 4741
tri 12326 4725 12342 4741 nw
tri 13490 4725 13506 4741 ne
rect 13506 4725 13524 4741
tri 2843 4686 2882 4725 ne
rect 2882 4686 5001 4725
tri 5001 4686 5040 4725 sw
rect 2277 4634 2283 4686
rect 2335 4634 2347 4686
rect 2399 4641 2405 4686
tri 2405 4641 2450 4686 sw
tri 2882 4685 2883 4686 ne
rect 2883 4685 5040 4686
tri 5040 4685 5041 4686 sw
tri 2883 4673 2895 4685 ne
rect 2895 4673 5041 4685
tri 2895 4647 2921 4673 ne
rect 2921 4647 5041 4673
tri 4962 4641 4968 4647 ne
rect 4968 4641 5041 4647
tri 5041 4641 5085 4685 sw
rect 12208 4667 12288 4725
tri 12288 4687 12326 4725 nw
tri 13506 4707 13524 4725 ne
rect 13438 4641 13490 4669
tri 1796 4610 1820 4634 se
rect 1820 4610 1909 4634
tri 2375 4610 2399 4634 ne
rect 2399 4610 2450 4641
tri 2450 4610 2481 4641 sw
tri 4968 4610 4999 4641 ne
rect 4999 4610 5085 4641
tri 5085 4610 5116 4641 sw
rect 1312 4558 1318 4610
rect 1370 4558 1382 4610
rect 1434 4590 1909 4610
tri 2399 4607 2402 4610 ne
rect 2402 4607 2481 4610
tri 2481 4607 2484 4610 sw
tri 4999 4607 5002 4610 ne
rect 5002 4607 5116 4610
tri 5116 4607 5119 4610 sw
tri 2402 4604 2405 4607 ne
rect 2405 4604 4908 4607
rect 1434 4589 1908 4590
tri 1908 4589 1909 4590 nw
tri 2405 4589 2420 4604 ne
rect 2420 4589 4908 4604
tri 4908 4589 4926 4607 sw
tri 5002 4589 5020 4607 ne
rect 5020 4589 5119 4607
tri 5119 4589 5137 4607 sw
rect 1434 4588 1907 4589
tri 1907 4588 1908 4589 nw
tri 2420 4588 2421 4589 ne
rect 2421 4588 4926 4589
tri 4926 4588 4927 4589 sw
tri 5020 4588 5021 4589 ne
rect 5021 4588 5137 4589
tri 5137 4588 5138 4589 sw
rect 1434 4577 1896 4588
tri 1896 4577 1907 4588 nw
tri 2421 4577 2432 4588 ne
rect 2432 4577 4927 4588
tri 4927 4577 4938 4588 sw
tri 5021 4577 5032 4588 ne
rect 5032 4577 5138 4588
tri 5138 4577 5149 4588 sw
rect 13438 4577 13490 4589
rect 1434 4558 1877 4577
tri 1877 4558 1896 4577 nw
tri 2432 4558 2451 4577 ne
rect 2451 4558 4938 4577
tri 4938 4558 4957 4577 sw
tri 5032 4568 5041 4577 ne
rect 5041 4568 5149 4577
tri 5149 4568 5158 4577 sw
tri 5041 4558 5051 4568 ne
rect 5051 4558 5158 4568
tri 5158 4558 5168 4568 sw
tri 2451 4549 2460 4558 ne
rect 2460 4549 4957 4558
tri 4854 4525 4878 4549 ne
rect 4878 4525 4957 4549
tri 4957 4525 4990 4558 sw
tri 5051 4525 5084 4558 ne
rect 5084 4525 5168 4558
tri 5168 4525 5201 4558 sw
tri 13412 4525 13438 4551 se
tri 4878 4517 4886 4525 ne
rect 4886 4517 4990 4525
tri 4990 4517 4998 4525 sw
tri 5084 4517 5092 4525 ne
rect 5092 4517 5201 4525
tri 5201 4517 5209 4525 sw
tri 13404 4517 13412 4525 se
rect 13412 4517 13490 4525
rect 2227 4465 2233 4517
rect 2285 4465 2297 4517
rect 2349 4511 4281 4517
tri 4886 4513 4890 4517 ne
rect 4890 4513 4998 4517
tri 4998 4513 5002 4517 sw
tri 5092 4513 5096 4517 ne
rect 5096 4513 5209 4517
tri 5209 4513 5213 4517 sw
tri 12760 4513 12764 4517 se
rect 12764 4513 13490 4517
rect 2349 4465 4229 4511
tri 4204 4459 4210 4465 ne
rect 4210 4459 4229 4465
tri 4890 4476 4927 4513 ne
rect 4927 4476 5002 4513
tri 5002 4476 5039 4513 sw
tri 5096 4476 5133 4513 ne
rect 5133 4476 5213 4513
tri 5213 4476 5250 4513 sw
tri 12723 4476 12760 4513 se
rect 12760 4476 13438 4513
tri 4927 4461 4942 4476 ne
rect 4942 4474 5039 4476
tri 5039 4474 5041 4476 sw
tri 5133 4474 5135 4476 ne
rect 5135 4474 5250 4476
rect 4942 4461 5041 4474
tri 5041 4461 5054 4474 sw
tri 5135 4461 5148 4474 ne
rect 5148 4461 5250 4474
tri 5250 4461 5265 4476 sw
tri 12708 4461 12723 4476 se
rect 12723 4461 13438 4476
tri 4210 4447 4222 4459 ne
rect 4222 4447 4281 4459
tri 4222 4440 4229 4447 ne
tri 4942 4445 4958 4461 ne
rect 4958 4451 5054 4461
tri 5054 4451 5064 4461 sw
tri 5148 4451 5158 4461 ne
rect 5158 4451 5265 4461
tri 5265 4451 5275 4461 sw
tri 12702 4455 12708 4461 se
rect 12708 4455 13490 4461
tri 12698 4451 12702 4455 se
rect 12702 4451 12764 4455
rect 4958 4445 5064 4451
tri 5064 4445 5070 4451 sw
tri 5158 4445 5164 4451 ne
rect 5164 4445 11394 4451
rect 4229 4389 4281 4395
tri 4958 4393 5010 4445 ne
rect 5010 4393 5070 4445
tri 5070 4393 5122 4445 sw
tri 5164 4393 5216 4445 ne
rect 5216 4393 11195 4445
rect 11247 4393 11266 4445
rect 11318 4393 11336 4445
rect 11388 4393 11394 4445
tri 12678 4431 12698 4451 se
rect 12698 4431 12764 4451
tri 12764 4431 12788 4455 nw
tri 5010 4389 5014 4393 ne
rect 5014 4389 5122 4393
tri 5122 4389 5126 4393 sw
tri 5216 4389 5220 4393 ne
rect 5220 4389 11394 4393
tri 5014 4375 5028 4389 ne
rect 5028 4375 5126 4389
tri 5126 4375 5140 4389 sw
tri 5220 4388 5221 4389 ne
rect 5221 4388 11394 4389
tri 12635 4388 12678 4431 se
rect 12678 4388 12708 4431
tri 12622 4375 12635 4388 se
rect 12635 4375 12708 4388
tri 12708 4375 12764 4431 nw
rect 13928 4375 14185 4828
tri 5028 4364 5039 4375 ne
rect 5039 4364 5140 4375
tri 5140 4364 5151 4375 sw
tri 12611 4364 12622 4375 se
rect 12622 4364 12678 4375
tri 5039 4361 5042 4364 ne
rect 5042 4361 5151 4364
rect 72 4355 2535 4361
tri 5042 4355 5048 4361 ne
rect 5048 4355 5151 4361
tri 5151 4355 5160 4364 sw
tri 12602 4355 12611 4364 se
rect 12611 4355 12678 4364
rect 72 4175 2483 4355
rect 2599 4175 2605 4355
tri 5048 4323 5080 4355 ne
rect 5080 4323 5160 4355
tri 5160 4323 5192 4355 sw
tri 12592 4345 12602 4355 se
rect 12602 4345 12678 4355
tri 12678 4345 12708 4375 nw
tri 12571 4324 12592 4345 se
rect 12592 4324 12657 4345
tri 12657 4324 12678 4345 nw
rect 12571 4323 12656 4324
tri 12656 4323 12657 4324 nw
rect 13928 4323 13991 4375
rect 14043 4323 14055 4375
rect 14107 4323 14119 4375
rect 14171 4323 14185 4375
tri 5080 4252 5151 4323 ne
rect 5151 4252 5192 4323
tri 5192 4252 5263 4323 sw
tri 5151 4175 5228 4252 ne
rect 5228 4175 5263 4252
tri 5263 4175 5340 4252 sw
rect 72 4168 2535 4175
tri 5228 4168 5235 4175 ne
rect 5235 4168 5340 4175
tri 5235 4140 5263 4168 ne
rect 5263 4140 5340 4168
tri 5340 4140 5375 4175 sw
tri 5263 4028 5375 4140 ne
tri 5375 4028 5487 4140 sw
tri 5375 3965 5438 4028 ne
rect 5438 3965 5487 4028
tri 5487 3965 5550 4028 sw
tri 12519 3965 12571 4017 se
rect 12571 3965 12623 4323
tri 12623 4290 12656 4323 nw
tri 5438 3959 5444 3965 ne
rect 5444 3959 5550 3965
tri 5550 3959 5556 3965 sw
tri 12513 3959 12519 3965 se
rect 12519 3959 12623 3965
tri 5444 3916 5487 3959 ne
rect 5487 3916 5556 3959
tri 5556 3916 5599 3959 sw
tri 12470 3916 12513 3959 se
rect 12513 3930 12623 3959
rect 12513 3916 12609 3930
tri 12609 3916 12623 3930 nw
rect 13928 3959 14185 4323
tri 5487 3911 5492 3916 ne
rect 5492 3911 11394 3916
tri 5492 3859 5544 3911 ne
rect 5544 3859 11195 3911
rect 11247 3859 11266 3911
rect 11318 3859 11336 3911
rect 11388 3859 11394 3911
tri 5544 3855 5548 3859 ne
rect 5548 3855 11394 3859
rect 12333 3911 12600 3916
rect 12333 3859 12339 3911
rect 12391 3859 12412 3911
rect 12464 3907 12600 3911
tri 12600 3907 12609 3916 nw
rect 13928 3907 13934 3959
rect 13986 3907 13999 3959
rect 12464 3895 12588 3907
tri 12588 3895 12600 3907 nw
rect 13928 3895 13999 3907
rect 12464 3859 12547 3895
rect 12333 3854 12547 3859
tri 12547 3854 12588 3895 nw
rect 13928 3843 13934 3895
rect 13986 3843 13999 3895
rect 14179 3843 14185 3959
rect 1576 3664 1582 3716
rect 1634 3664 1646 3716
rect 1698 3664 1704 3716
rect 1888 3664 1894 3716
rect 1946 3664 1958 3716
rect 2010 3664 2016 3716
rect 1576 3582 1582 3634
rect 1634 3582 1646 3634
rect 1698 3582 1704 3634
rect 1576 3552 1704 3582
rect 1576 3500 1582 3552
rect 1634 3500 1646 3552
rect 1698 3500 1704 3552
rect 1888 3582 1894 3634
rect 1946 3582 1958 3634
rect 2010 3582 2016 3634
rect 1888 3552 2016 3582
rect 1888 3500 1894 3552
rect 1946 3500 1958 3552
rect 2010 3500 2016 3552
rect 1147 3354 1199 3360
rect 1147 3290 1199 3302
rect 1147 3226 1199 3238
rect 1147 3168 1199 3174
rect 1459 3354 1511 3360
rect 1459 3290 1511 3302
rect 1459 3226 1511 3238
rect 1459 3168 1511 3174
rect 1771 3354 1823 3360
rect 1771 3290 1823 3302
rect 1771 3226 1823 3238
rect 1771 3168 1823 3174
rect 2080 3354 2132 3360
rect 2080 3290 2132 3302
rect 2080 3226 2132 3238
rect 2080 3168 2132 3174
rect 2837 3308 2889 3314
rect 2837 3244 2889 3256
rect 2837 3180 2889 3192
rect 2837 3116 2889 3128
rect 1147 3093 1199 3099
rect 1147 3029 1199 3041
rect 1147 2965 1199 2977
rect 1147 2901 1199 2913
rect 1147 2843 1199 2849
rect 1459 3093 1511 3099
rect 1459 3029 1511 3041
rect 1459 2965 1511 2977
rect 1459 2901 1511 2913
rect 1459 2843 1511 2849
rect 1771 3093 1823 3099
rect 1771 3029 1823 3041
rect 1771 2965 1823 2977
rect 1771 2901 1823 2913
rect 1771 2843 1823 2849
rect 2080 3093 2132 3099
rect 2837 3058 2889 3064
rect 2080 3029 2132 3041
rect 2080 2965 2132 2977
rect 2080 2901 2132 2913
rect 2080 2843 2132 2849
rect 13928 2183 14185 3843
rect 14388 6089 14451 6141
rect 14503 6089 14515 6141
rect 14567 6089 14579 6141
rect 14631 6089 14637 6141
rect 14388 5636 14637 6089
rect 14388 5584 14451 5636
rect 14503 5584 14515 5636
rect 14567 5584 14579 5636
rect 14631 5584 14637 5636
rect 14388 5133 14637 5584
rect 14388 5081 14451 5133
rect 14503 5081 14515 5133
rect 14567 5081 14579 5133
rect 14631 5081 14637 5133
rect 14388 4628 14637 5081
rect 14388 4576 14451 4628
rect 14503 4576 14515 4628
rect 14567 4576 14579 4628
rect 14631 4576 14637 4628
rect 14388 3965 14637 4576
rect 14388 3913 14394 3965
rect 14446 3913 14487 3965
rect 14539 3913 14579 3965
rect 14631 3913 14637 3965
rect 14388 3901 14637 3913
rect 14388 3849 14394 3901
rect 14446 3849 14487 3901
rect 14539 3849 14579 3901
rect 14631 3849 14637 3901
rect 14388 3774 14637 3849
rect 14388 3722 14394 3774
rect 14446 3722 14487 3774
rect 14539 3722 14579 3774
rect 14631 3722 14637 3774
rect 14388 3710 14637 3722
rect 14388 3658 14394 3710
rect 14446 3658 14487 3710
rect 14539 3658 14579 3710
rect 14631 3658 14637 3710
rect 14388 3637 14637 3658
<< comment >>
rect 2831 6739 2895 6782
rect 2831 6484 2895 6547
rect 2821 6163 4211 6339
rect 2821 5349 4211 6053
use DFL1_CDNS_524688791851160  DFL1_CDNS_524688791851160_0
timestamp 1707688321
transform -1 0 243 0 -1 5849
box 0 0 1 1
use DFL1_CDNS_524688791851160  DFL1_CDNS_524688791851160_1
timestamp 1707688321
transform -1 0 243 0 -1 5599
box 0 0 1 1
use DFL1_CDNS_524688791851160  DFL1_CDNS_524688791851160_2
timestamp 1707688321
transform 1 0 1309 0 -1 5849
box 0 0 1 1
use DFL1_CDNS_524688791851160  DFL1_CDNS_524688791851160_3
timestamp 1707688321
transform 1 0 1309 0 -1 5599
box 0 0 1 1
use hvDFL1sd_CDNS_52468879185349  hvDFL1sd_CDNS_52468879185349_0
timestamp 1707688321
transform 0 -1 2160 -1 0 3927
box 0 0 1 1
use hvDFL1sd_CDNS_52468879185349  hvDFL1sd_CDNS_52468879185349_1
timestamp 1707688321
transform 0 1 1826 -1 0 3927
box 0 0 1 1
use hvDFL1sd_CDNS_52468879185349  hvDFL1sd_CDNS_52468879185349_2
timestamp 1707688321
transform 0 1 1826 1 0 4327
box 0 0 1 1
use hvDFL1sd_CDNS_52468879185349  hvDFL1sd_CDNS_52468879185349_3
timestamp 1707688321
transform 0 -1 2160 1 0 4327
box 0 0 1 1
use hvDFL1sd_CDNS_52468879185354  hvDFL1sd_CDNS_52468879185354_0
timestamp 1707688321
transform -1 0 838 0 1 5541
box 0 0 1 1
use hvDFL1sd_CDNS_52468879185354  hvDFL1sd_CDNS_52468879185354_1
timestamp 1707688321
transform -1 0 314 0 1 5541
box 0 0 1 1
use hvDFL1sd_CDNS_52468879185354  hvDFL1sd_CDNS_52468879185354_2
timestamp 1707688321
transform 1 0 1238 0 1 5541
box 0 0 1 1
use hvDFL1sd_CDNS_52468879185354  hvDFL1sd_CDNS_52468879185354_3
timestamp 1707688321
transform 1 0 714 0 1 5541
box 0 0 1 1
use hvnTran_CDNS_524688791851481  hvnTran_CDNS_524688791851481_0
timestamp 1707688321
transform 0 -1 4197 1 0 4739
box -79 -26 335 626
use hvnTran_CDNS_524688791851481  hvnTran_CDNS_524688791851481_1
timestamp 1707688321
transform 0 -1 3503 1 0 4739
box -79 -26 335 626
use hvnTran_CDNS_524688791851482  hvnTran_CDNS_524688791851482_0
timestamp 1707688321
transform 0 -1 3503 1 0 3693
box -79 -26 959 626
use hvnTran_CDNS_524688791851482  hvnTran_CDNS_524688791851482_1
timestamp 1707688321
transform 0 -1 4197 1 0 3693
box -79 -26 959 626
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1707688321
transform 0 1 349 -1 0 6987
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_1
timestamp 1707688321
transform -1 0 1078 0 1 4263
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_2
timestamp 1707688321
transform -1 0 1960 0 1 4203
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_3
timestamp 1707688321
transform -1 0 2060 0 1 4263
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_4
timestamp 1707688321
transform -1 0 1866 0 1 4263
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_5
timestamp 1707688321
transform 0 1 1115 1 0 4644
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_6
timestamp 1707688321
transform 0 -1 252 1 0 4644
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_7
timestamp 1707688321
transform 1 0 2849 0 1 6372
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_8
timestamp 1707688321
transform 1 0 381 0 1 4502
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1707688321
transform 0 -1 1261 -1 0 4875
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1707688321
transform 0 -1 1160 -1 0 3706
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1707688321
transform 0 -1 2352 -1 0 8153
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1707688321
transform 0 -1 2429 -1 0 7895
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1707688321
transform 0 -1 508 -1 0 4128
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1707688321
transform 0 -1 2275 -1 0 7533
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1707688321
transform 0 -1 3232 -1 0 7766
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1707688321
transform 0 -1 322 -1 0 4874
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1707688321
transform -1 0 1694 0 1 3594
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_9
timestamp 1707688321
transform -1 0 2006 0 1 3594
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_10
timestamp 1707688321
transform -1 0 2318 0 1 3594
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_11
timestamp 1707688321
transform -1 0 1382 0 1 3594
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_12
timestamp 1707688321
transform -1 0 1248 0 1 4508
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_13
timestamp 1707688321
transform -1 0 1430 0 1 4564
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_14
timestamp 1707688321
transform -1 0 2269 0 1 4564
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_15
timestamp 1707688321
transform -1 0 1734 0 1 4564
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_16
timestamp 1707688321
transform -1 0 1010 0 1 4564
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_17
timestamp 1707688321
transform -1 0 1842 0 1 4016
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_18
timestamp 1707688321
transform -1 0 2250 0 1 4113
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_19
timestamp 1707688321
transform 0 1 1305 1 0 4983
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_20
timestamp 1707688321
transform 0 1 2089 1 0 4983
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_21
timestamp 1707688321
transform 0 1 474 1 0 4203
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_22
timestamp 1707688321
transform 0 1 2315 1 0 4486
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_23
timestamp 1707688321
transform 0 1 49 1 0 7889
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_24
timestamp 1707688321
transform 0 -1 637 1 0 4983
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_25
timestamp 1707688321
transform 0 -1 949 1 0 4983
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_26
timestamp 1707688321
transform 0 -1 247 1 0 4983
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_27
timestamp 1707688321
transform 0 -1 1802 1 0 4927
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_28
timestamp 1707688321
transform 0 -1 1573 1 0 4769
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_29
timestamp 1707688321
transform 0 -1 1885 1 0 4769
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_30
timestamp 1707688321
transform 0 -1 936 1 0 4078
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_31
timestamp 1707688321
transform 0 -1 2148 1 0 4203
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_32
timestamp 1707688321
transform 1 0 225 0 -1 3712
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_33
timestamp 1707688321
transform 1 0 605 0 -1 3712
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_34
timestamp 1707688321
transform 1 0 3375 0 -1 6583
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_35
timestamp 1707688321
transform 1 0 3046 0 -1 7607
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1707688321
transform 0 -1 793 -1 0 5320
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1707688321
transform 0 -1 220 -1 0 250
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_2
timestamp 1707688321
transform 0 -1 481 -1 0 5320
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_3
timestamp 1707688321
transform 0 -1 169 -1 0 5320
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_4
timestamp 1707688321
transform 0 -1 1105 -1 0 5320
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_5
timestamp 1707688321
transform 0 -1 1729 -1 0 5320
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_6
timestamp 1707688321
transform 0 -1 2041 -1 0 5320
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_7
timestamp 1707688321
transform 0 -1 1472 -1 0 3970
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_8
timestamp 1707688321
transform 0 -1 114 -1 0 3970
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_9
timestamp 1707688321
transform 0 -1 652 -1 0 250
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_10
timestamp 1707688321
transform 0 -1 2126 -1 0 3540
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_11
timestamp 1707688321
transform 0 -1 1814 -1 0 3540
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_12
timestamp 1707688321
transform 0 -1 1502 -1 0 3540
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_13
timestamp 1707688321
transform 0 -1 1190 -1 0 3540
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_14
timestamp 1707688321
transform 0 -1 2271 -1 0 5320
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_15
timestamp 1707688321
transform 0 -1 1417 -1 0 5320
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_16
timestamp 1707688321
transform 0 1 3368 -1 0 7107
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_17
timestamp 1707688321
transform 1 0 325 0 -1 5743
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_18
timestamp 1707688321
transform 1 0 2942 0 -1 6651
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_19
timestamp 1707688321
transform 1 0 3500 0 -1 7640
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_0
timestamp 1707688321
transform 1 0 2849 0 1 6555
box 0 0 1 1
use L1M1_CDNS_52468879185193  L1M1_CDNS_52468879185193_0
timestamp 1707688321
transform 1 0 1832 0 -1 3869
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_0
timestamp 1707688321
transform 1 0 3426 0 -1 6657
box 0 0 1 1
use L1M1_CDNS_52468879185308  L1M1_CDNS_52468879185308_0
timestamp 1707688321
transform 0 1 2092 1 0 2693
box 0 0 1 1
use L1M1_CDNS_52468879185308  L1M1_CDNS_52468879185308_1
timestamp 1707688321
transform 0 1 1780 1 0 2693
box 0 0 1 1
use L1M1_CDNS_52468879185308  L1M1_CDNS_52468879185308_2
timestamp 1707688321
transform 0 1 1468 1 0 2693
box 0 0 1 1
use L1M1_CDNS_52468879185308  L1M1_CDNS_52468879185308_3
timestamp 1707688321
transform 0 1 1156 1 0 2693
box 0 0 1 1
use L1M1_CDNS_52468879185334  L1M1_CDNS_52468879185334_0
timestamp 1707688321
transform 0 1 2491 1 0 3168
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_0
timestamp 1707688321
transform -1 0 1505 0 1 4428
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1707688321
transform 0 -1 4281 -1 0 4517
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1707688321
transform 0 1 282 -1 0 4887
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1707688321
transform 0 1 1221 -1 0 4887
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1707688321
transform -1 0 465 0 1 6946
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1707688321
transform -1 0 1440 0 -1 4610
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_5
timestamp 1707688321
transform 1 0 2227 0 -1 4517
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_6
timestamp 1707688321
transform 1 0 1888 0 1 3664
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_7
timestamp 1707688321
transform 1 0 1888 0 1 3582
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_8
timestamp 1707688321
transform 1 0 1888 0 1 3500
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_9
timestamp 1707688321
transform 1 0 1576 0 1 3664
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_10
timestamp 1707688321
transform 1 0 1576 0 1 3582
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_11
timestamp 1707688321
transform 1 0 1576 0 1 3500
box 0 0 1 1
use M1M2_CDNS_52468879185197  M1M2_CDNS_52468879185197_0
timestamp 1707688321
transform 0 1 -248 1 0 3476
box 0 0 256 116
use M1M2_CDNS_52468879185197  M1M2_CDNS_52468879185197_1
timestamp 1707688321
transform 0 1 -248 1 0 2589
box 0 0 256 116
use M1M2_CDNS_52468879185197  M1M2_CDNS_52468879185197_2
timestamp 1707688321
transform 0 1 -104 1 0 889
box 0 0 256 116
use M1M2_CDNS_52468879185197  M1M2_CDNS_52468879185197_3
timestamp 1707688321
transform 0 1 -104 1 0 3127
box 0 0 256 116
use M1M2_CDNS_52468879185197  M1M2_CDNS_52468879185197_4
timestamp 1707688321
transform 0 1 2487 1 0 3127
box 0 0 256 116
use M1M2_CDNS_52468879185197  M1M2_CDNS_52468879185197_5
timestamp 1707688321
transform 1 0 13929 0 1 2202
box 0 0 256 116
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_0
timestamp 1707688321
transform 1 0 2965 0 1 4771
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_0
timestamp 1707688321
transform 1 0 2477 0 1 4175
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_0
timestamp 1707688321
transform 0 -1 2889 1 0 6782
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_0
timestamp 1707688321
transform 0 1 1147 1 0 3168
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_1
timestamp 1707688321
transform 0 1 1459 1 0 3168
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_2
timestamp 1707688321
transform 0 1 1771 1 0 3168
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_3
timestamp 1707688321
transform 0 1 2080 1 0 3168
box 0 0 1 1
use M1M2_CDNS_52468879185208  M1M2_CDNS_52468879185208_0
timestamp 1707688321
transform 1 0 13524 0 -1 4803
box 0 0 192 244
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_0
timestamp 1707688321
transform 0 -1 3322 -1 0 7115
box 0 0 1 1
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_1
timestamp 1707688321
transform 0 -1 2889 -1 0 3314
box 0 0 1 1
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_2
timestamp 1707688321
transform 0 1 1147 1 0 2843
box 0 0 1 1
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_3
timestamp 1707688321
transform 0 1 1459 1 0 2843
box 0 0 1 1
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_4
timestamp 1707688321
transform 0 1 1771 1 0 2843
box 0 0 1 1
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_5
timestamp 1707688321
transform 0 1 2080 1 0 2843
box 0 0 1 1
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_6
timestamp 1707688321
transform 1 0 148 0 -1 7323
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_0
timestamp 1707688321
transform 1 0 1762 0 1 4915
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_1
timestamp 1707688321
transform 1 0 2831 0 1 4915
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_2
timestamp 1707688321
transform 1 0 1845 0 1 4771
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_3
timestamp 1707688321
transform 1 0 2831 0 1 4771
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_4
timestamp 1707688321
transform 1 0 4229 0 1 4771
box 0 0 1 1
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_0
timestamp 1707688321
transform 1 0 13524 0 -1 5082
box 0 0 192 180
use M1M2_CDNS_524688791851084  M1M2_CDNS_524688791851084_0
timestamp 1707688321
transform 0 1 -104 1 0 6261
box 0 0 512 52
use M1M2_CDNS_524688791851113  M1M2_CDNS_524688791851113_0
timestamp 1707688321
transform 0 1 -40 1 0 6261
box 0 0 1 1
use M1M2_CDNS_524688791851177  M1M2_CDNS_524688791851177_0
timestamp 1707688321
transform 1 0 13029 0 1 7271
box 0 0 384 116
use M1M2_CDNS_524688791851177  M1M2_CDNS_524688791851177_1
timestamp 1707688321
transform 1 0 13029 0 1 6552
box 0 0 384 116
use nfet_CDNS_52468879185310  nfet_CDNS_52468879185310_0
timestamp 1707688321
transform -1 0 1713 0 1 3780
box -79 -26 199 626
use nfet_CDNS_52468879185310  nfet_CDNS_52468879185310_1
timestamp 1707688321
transform 1 0 2273 0 1 3780
box -79 -26 199 626
use nfet_CDNS_52468879185344  nfet_CDNS_52468879185344_0
timestamp 1707688321
transform -1 0 1427 0 1 3780
box -79 -26 179 626
use nfet_CDNS_52468879185344  nfet_CDNS_52468879185344_1
timestamp 1707688321
transform -1 0 1271 0 1 3780
box -79 -26 179 626
use nfet_CDNS_52468879185344  nfet_CDNS_52468879185344_2
timestamp 1707688321
transform -1 0 959 0 1 3780
box -79 -26 179 626
use nfet_CDNS_52468879185344  nfet_CDNS_52468879185344_3
timestamp 1707688321
transform -1 0 1115 0 1 3780
box -79 -26 179 626
use nfet_CDNS_52468879185344  nfet_CDNS_52468879185344_4
timestamp 1707688321
transform 1 0 125 0 1 3780
box -79 -26 179 626
use nfet_CDNS_52468879185344  nfet_CDNS_52468879185344_5
timestamp 1707688321
transform 1 0 281 0 1 3780
box -79 -26 179 626
use nfet_CDNS_52468879185344  nfet_CDNS_52468879185344_6
timestamp 1707688321
transform 1 0 437 0 1 3780
box -79 -26 179 626
use nfet_CDNS_52468879185344  nfet_CDNS_52468879185344_7
timestamp 1707688321
transform 1 0 593 0 1 3780
box -79 -26 179 626
use nfet_CDNS_524688791851483  nfet_CDNS_524688791851483_0
timestamp 1707688321
transform 1 0 1825 0 1 3014
box -79 -26 647 626
use nfet_CDNS_524688791851483  nfet_CDNS_524688791851483_1
timestamp 1707688321
transform 1 0 1201 0 1 3014
box -79 -26 647 626
use pfet_CDNS_52468879185324  pfet_CDNS_52468879185324_0
timestamp 1707688321
transform 1 0 180 0 1 4732
box -119 -66 375 666
use pfet_CDNS_52468879185324  pfet_CDNS_52468879185324_1
timestamp 1707688321
transform 1 0 1116 0 1 4732
box -119 -66 375 666
use pfet_CDNS_52468879185368  pfet_CDNS_52468879185368_0
timestamp 1707688321
transform -1 0 748 0 1 4732
box -119 -66 375 666
use pfet_CDNS_52468879185368  pfet_CDNS_52468879185368_1
timestamp 1707688321
transform -1 0 1060 0 1 4732
box -119 -66 375 666
use pfet_CDNS_524688791851484  pfet_CDNS_524688791851484_0
timestamp 1707688321
transform 0 -1 16532 1 0 5482
box -119 -66 375 3066
use pfet_CDNS_524688791851484  pfet_CDNS_524688791851484_1
timestamp 1707688321
transform 0 -1 16532 1 0 4978
box -119 -66 375 3066
use pfet_CDNS_524688791851484  pfet_CDNS_524688791851484_2
timestamp 1707688321
transform 0 -1 16532 1 0 4474
box -119 -66 375 3066
use pfet_CDNS_524688791851484  pfet_CDNS_524688791851484_3
timestamp 1707688321
transform 0 -1 16532 1 0 5986
box -119 -66 375 3066
use pfet_CDNS_524688791851485  pfet_CDNS_524688791851485_0
timestamp 1707688321
transform -1 0 714 0 1 5791
box -119 -66 519 150
use pfet_CDNS_524688791851485  pfet_CDNS_524688791851485_1
timestamp 1707688321
transform 1 0 838 0 1 5791
box -119 -66 519 150
use pfet_CDNS_524688791851486  pfet_CDNS_524688791851486_0
timestamp 1707688321
transform 1 0 1428 0 1 4732
box -119 -66 687 666
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_0
timestamp 1707688321
transform 0 -1 2060 -1 0 5498
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_1
timestamp 1707688321
transform -1 0 741 0 1 5364
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_2
timestamp 1707688321
transform -1 0 1172 0 1 5443
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_3
timestamp 1707688321
transform -1 0 2297 0 1 4412
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_4
timestamp 1707688321
transform -1 0 273 0 1 4628
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_5
timestamp 1707688321
transform -1 0 1233 0 1 4622
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_6
timestamp 1707688321
transform 1 0 380 0 1 5443
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_7
timestamp 1707688321
transform 1 0 811 0 1 5364
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_8
timestamp 1707688321
transform 1 0 1678 0 1 4412
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1707688321
transform 0 -1 225 -1 0 3748
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_1
timestamp 1707688321
transform 0 1 593 -1 0 3748
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_2
timestamp 1707688321
transform -1 0 959 0 1 4412
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_3
timestamp 1707688321
transform -1 0 1264 0 1 4412
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_4
timestamp 1707688321
transform 1 0 1978 0 1 3903
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_5
timestamp 1707688321
transform 1 0 1942 0 1 4193
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_6
timestamp 1707688321
transform 1 0 288 0 1 4412
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_7
timestamp 1707688321
transform 1 0 1327 0 1 4412
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_0
timestamp 1707688321
transform 0 1 314 1 0 5693
box 0 0 1 1
use PYL1_CDNS_52468879185318  PYL1_CDNS_52468879185318_0
timestamp 1707688321
transform 0 1 1227 1 0 3646
box 0 0 66 542
use PYL1_CDNS_52468879185318  PYL1_CDNS_52468879185318_1
timestamp 1707688321
transform 0 -1 2367 1 0 3646
box 0 0 66 542
use PYL1_CDNS_524688791851468  PYL1_CDNS_524688791851468_0
timestamp 1707688321
transform 1 0 46 0 -1 3479
box 0 0 66 3262
use sky130_fd_io__sio_hotswap_hys  sky130_fd_io__sio_hotswap_hys_0
timestamp 1707688321
transform 0 1 3100 1 0 6543
box 0 -76 1215 674
use sky130_fd_io__sio_hotswap_wpd  sky130_fd_io__sio_hotswap_wpd_0
timestamp 1707688321
transform 0 -1 520 1 0 63
box -161 -62 3595 434
use sky130_fd_io__sio_hotswap_wpd  sky130_fd_io__sio_hotswap_wpd_1
timestamp 1707688321
transform 0 -1 952 1 0 63
box -161 -62 3595 434
use sky130_fd_io__sio_hvsbt_inv_x1  sky130_fd_io__sio_hvsbt_inv_x1_0
timestamp 1707688321
transform -1 0 316 0 1 6900
box -107 21 267 1369
use sky130_fd_io__sio_hvsbt_inv_x1  sky130_fd_io__sio_hvsbt_inv_x1_1
timestamp 1707688321
transform 0 1 2821 1 0 6339
box -107 21 267 1369
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_0
timestamp 1707688321
transform 0 1 4229 1 0 4668
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_524688791851476  sky130_fd_io__tk_em1o_CDNS_524688791851476_0
timestamp 1707688321
transform 0 1 3266 -1 0 6796
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_524688791851477  sky130_fd_io__tk_em1o_CDNS_524688791851477_0
timestamp 1707688321
transform -1 0 3753 0 -1 5046
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_524688791851478  sky130_fd_io__tk_em1o_CDNS_524688791851478_0
timestamp 1707688321
transform 0 1 2831 -1 0 3733
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_0
timestamp 1707688321
transform 0 1 4229 -1 0 4441
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185341  sky130_fd_io__tk_em1s_CDNS_52468879185341_0
timestamp 1707688321
transform -1 0 3414 0 -1 6589
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851473  sky130_fd_io__tk_em1s_CDNS_524688791851473_0
timestamp 1707688321
transform -1 0 3797 0 -1 3644
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851474  sky130_fd_io__tk_em1s_CDNS_524688791851474_0
timestamp 1707688321
transform 0 1 2831 -1 0 4805
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851475  sky130_fd_io__tk_em1s_CDNS_524688791851475_0
timestamp 1707688321
transform 1 0 3270 0 1 6859
box 0 0 1 1
use TPL1_CDNS_524688791851469  TPL1_CDNS_524688791851469_0
timestamp 1707688321
transform -1 0 13180 0 -1 6545
box -26 -26 108 2412
use TPL1_CDNS_524688791851469  TPL1_CDNS_524688791851469_1
timestamp 1707688321
transform -1 0 13112 0 -1 6545
box -26 -26 108 2412
use TPL1_CDNS_524688791851470  TPL1_CDNS_524688791851470_0
timestamp 1707688321
transform 0 1 13136 -1 0 6618
box -26 -26 108 3780
use TPL1_CDNS_524688791851470  TPL1_CDNS_524688791851470_1
timestamp 1707688321
transform 0 1 13136 -1 0 4101
box -26 -26 108 3780
use TPL1_CDNS_524688791851470  TPL1_CDNS_524688791851470_2
timestamp 1707688321
transform 0 1 13136 -1 0 6686
box -26 -26 108 3780
use TPL1_CDNS_524688791851470  TPL1_CDNS_524688791851470_3
timestamp 1707688321
transform 0 1 13136 -1 0 4169
box -26 -26 108 3780
use TPL1_CDNS_524688791851471  TPL1_CDNS_524688791851471_0
timestamp 1707688321
transform -1 0 16985 0 -1 6549
box -26 -26 108 2420
use TPL1_CDNS_524688791851471  TPL1_CDNS_524688791851471_1
timestamp 1707688321
transform -1 0 16917 0 -1 6549
box -26 -26 108 2420
use TPL1_CDNS_524688791851472  TPL1_CDNS_524688791851472_0
timestamp 1707688321
transform 1 0 2213 0 -1 5332
box -36 -36 118 594
<< labels >>
flabel comment s 2831 6739 2895 6782 0 FreeSans 50 180 0 0 optional to vgnd
port 1 nsew
flabel comment s 1855 3899 1855 3899 0 FreeSans 300 90 0 0 S
flabel comment s 1855 4355 1855 4355 0 FreeSans 300 90 0 0 D
flabel comment s 2131 3899 2131 3899 0 FreeSans 300 90 0 0 S
flabel comment s 2131 4355 2131 4355 0 FreeSans 300 90 0 0 D
flabel comment s 742 5570 742 5570 0 FreeSans 300 180 0 0 S
flabel comment s 286 5570 286 5570 0 FreeSans 300 180 0 0 D
flabel comment s 810 5570 810 5570 0 FreeSans 300 0 0 0 S
flabel comment s 1266 5570 1266 5570 0 FreeSans 300 0 0 0 D
flabel metal1 s 2831 7090 2895 7102 3 FreeSans 200 270 0 0 vgnd
port 3 nsew
flabel metal1 s 2831 3058 2895 3070 3 FreeSans 200 90 0 0 vgnd
port 3 nsew
flabel metal1 s 1656 4517 1656 4517 0 FreeSans 100 0 0 0 enhs_h
flabel metal1 s 1637 4931 1637 4931 0 FreeSans 100 0 0 0 n6
flabel metal1 s 1637 4878 1637 4878 0 FreeSans 100 0 0 0 n2
flabel metal1 s 3192 6339 3238 6351 3 FreeSans 200 90 0 0 vgnd
port 3 nsew
flabel metal1 s 2923 6339 3164 6351 3 FreeSans 200 90 0 0 vgnd
port 3 nsew
flabel metal1 s -132 7271 -104 7317 0 FreeSans 200 0 0 0 vgnd
port 3 nsew
flabel metal1 s 3416 2803 3614 2841 7 FreeSans 200 270 0 0 pghs_h
port 4 nsew
flabel metal1 s 3414 6339 3690 6368 3 FreeSans 200 90 0 0 vcc_io
port 5 nsew
flabel metal1 s 3266 6498 3298 6532 7 FreeSans 200 270 0 0 enhs_lat_h_n
port 6 nsew
flabel metal1 s 2226 3588 2356 3626 0 FreeSans 200 270 0 0 pghs_h
port 4 nsew
flabel metal1 s 140 7493 169 7769 0 FreeSans 200 0 0 0 vcc_io
port 5 nsew
flabel metal1 s 73 7041 101 7243 0 FreeSans 200 0 0 0 vgnd
port 3 nsew
flabel metal1 s 2355 4632 2367 4690 0 FreeSans 200 0 0 0 pad_esd
port 7 nsew
flabel metal1 s 2260 5130 2287 5332 0 FreeSans 200 0 0 0 vcc_io
port 5 nsew
flabel locali s 164 -72 180 -38 0 FreeSans 200 0 0 0 vgnd
port 3 nsew
flabel locali s 349 6953 455 6987 0 FreeSans 200 270 0 0 enhs_lathys_h_n
port 8 nsew
flabel locali s 62 217 96 3479 0 FreeSans 200 180 0 0 vpwr_ka
port 9 nsew
flabel locali s 2315 5439 2355 5471 0 FreeSans 200 0 0 0 enhs_h
port 10 nsew
flabel locali s 2163 5439 2203 5471 0 FreeSans 200 0 0 0 dishs_h
port 11 nsew
flabel locali s 1994 5443 2060 5472 0 FreeSans 200 0 0 0 dishs_h_n
port 12 nsew
flabel locali s 2392 5439 2432 5472 0 FreeSans 200 0 0 0 exiths_h
port 13 nsew
flabel metal2 s 1656 6722 1656 6722 0 FreeSans 100 0 0 0 enhs_lathys_h_n
<< properties >>
string GDS_END 88805792
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 88596482
string path 365.925 140.250 359.700 140.250 
<< end >>
