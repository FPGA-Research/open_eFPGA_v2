magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -38 261 1602 582
<< pwell >>
rect 833 157 1563 203
rect 1 21 1563 157
rect 30 -17 64 21
<< locali >>
rect 17 197 65 325
rect 292 191 358 265
rect 890 199 1087 265
rect 1212 51 1282 493
rect 1495 357 1547 493
rect 1513 119 1547 357
rect 1495 51 1547 119
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 17 393 69 493
rect 103 427 169 527
rect 17 359 156 393
rect 122 280 156 359
rect 203 337 248 493
rect 122 214 168 280
rect 122 161 156 214
rect 17 127 156 161
rect 17 69 69 127
rect 103 17 169 93
rect 203 69 237 337
rect 291 333 357 483
rect 391 367 454 527
rect 549 451 717 485
rect 654 425 717 451
rect 751 427 918 527
rect 661 415 717 425
rect 679 409 717 415
rect 679 403 721 409
rect 585 381 626 399
rect 683 398 721 403
rect 684 395 721 398
rect 686 392 721 395
rect 291 299 428 333
rect 394 219 428 299
rect 494 271 551 337
rect 585 315 653 381
rect 394 157 468 219
rect 585 207 619 315
rect 687 265 721 392
rect 956 373 990 487
rect 1024 387 1178 527
rect 768 353 990 373
rect 768 307 1178 353
rect 687 233 840 265
rect 307 153 468 157
rect 520 153 619 207
rect 666 199 840 233
rect 307 123 428 153
rect 307 69 341 123
rect 666 107 700 199
rect 1131 165 1178 307
rect 375 17 441 89
rect 554 73 700 107
rect 848 131 1178 165
rect 747 17 814 106
rect 848 51 908 131
rect 1024 17 1178 97
rect 1316 265 1366 493
rect 1402 367 1461 527
rect 1316 199 1479 265
rect 1316 51 1361 199
rect 1395 17 1461 93
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
<< metal1 >>
rect 0 561 1564 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 0 496 1564 527
rect 0 17 1564 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
rect 0 -48 1564 -17
<< obsm1 >>
rect 202 388 260 397
rect 573 388 631 397
rect 202 360 631 388
rect 202 351 260 360
rect 573 351 631 360
rect 110 320 168 329
rect 482 320 540 329
rect 110 292 540 320
rect 110 283 168 292
rect 482 283 540 292
<< labels >>
rlabel locali s 292 191 358 265 6 D
port 1 nsew signal input
rlabel locali s 17 197 65 325 6 GATE
port 2 nsew clock input
rlabel locali s 890 199 1087 265 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 0 -48 1564 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 1563 157 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 833 157 1563 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 1602 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 1564 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1212 51 1282 493 6 Q
port 8 nsew signal output
rlabel locali s 1495 51 1547 119 6 Q_N
port 9 nsew signal output
rlabel locali s 1513 119 1547 357 6 Q_N
port 9 nsew signal output
rlabel locali s 1495 357 1547 493 6 Q_N
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1564 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2696512
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2683288
<< end >>
