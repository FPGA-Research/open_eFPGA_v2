magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -119 -66 375 366
<< mvpmos >>
rect 0 0 100 300
rect 156 0 256 300
<< mvpdiff >>
rect -50 0 0 300
rect 100 250 156 300
rect 100 216 111 250
rect 145 216 156 250
rect 100 182 156 216
rect 100 148 111 182
rect 145 148 156 182
rect 100 114 156 148
rect 100 80 111 114
rect 145 80 156 114
rect 100 46 156 80
rect 100 12 111 46
rect 145 12 156 46
rect 100 0 156 12
rect 256 0 306 300
<< mvpdiffc >>
rect 111 216 145 250
rect 111 148 145 182
rect 111 80 145 114
rect 111 12 145 46
<< poly >>
rect 0 300 100 326
rect 156 300 256 326
rect 0 -26 100 0
rect 156 -26 256 0
<< locali >>
rect 111 250 145 266
rect 111 182 145 216
rect 111 114 145 148
rect 111 46 145 80
rect 111 -4 145 12
<< metal1 >>
rect -51 -16 -5 258
rect 261 -16 307 258
use hvDFL1sd2_CDNS_52468879185277  hvDFL1sd2_CDNS_52468879185277_0
timestamp 1707688321
transform 1 0 100 0 1 0
box 0 0 1 1
use hvDFM1sd_CDNS_52468879185274  hvDFM1sd_CDNS_52468879185274_0
timestamp 1707688321
transform -1 0 0 0 1 0
box -36 -36 89 336
use hvDFM1sd_CDNS_52468879185274  hvDFM1sd_CDNS_52468879185274_1
timestamp 1707688321
transform 1 0 256 0 1 0
box -36 -36 89 336
<< labels >>
flabel comment s -28 121 -28 121 0 FreeSans 300 0 0 0 S
flabel comment s 128 131 128 131 0 FreeSans 300 0 0 0 D
flabel comment s 284 121 284 121 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 86837476
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86835958
<< end >>
