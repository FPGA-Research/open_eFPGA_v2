magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -76 -26 176 1026
<< mvnmos >>
rect 0 0 100 1000
<< mvndiff >>
rect -50 0 0 1000
rect 100 0 150 1000
<< poly >>
rect 0 1000 100 1032
rect 0 -32 100 0
<< locali >>
rect -45 -4 -11 946
rect 111 -4 145 946
use DFL1sd_CDNS_5246887918593  DFL1sd_CDNS_5246887918593_0
timestamp 1707688321
transform 1 0 100 0 1 0
box -26 -26 79 1026
use hvDFL1sd_CDNS_5246887918592  hvDFL1sd_CDNS_5246887918592_0
timestamp 1707688321
transform -1 0 0 0 1 0
box -26 -26 79 1026
<< labels >>
flabel comment s -28 471 -28 471 0 FreeSans 300 0 0 0 S
flabel comment s 128 471 128 471 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 80568090
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 80567202
<< end >>
