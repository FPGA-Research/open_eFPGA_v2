magic
tech sky130A
magscale 1 2
timestamp 1707688321
use sky130_fd_pr__nfet_01v8__example_55959141808248  sky130_fd_pr__nfet_01v8__example_55959141808248_0
timestamp 1707688321
transform 1 0 754 0 1 228
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808445  sky130_fd_pr__nfet_01v8__example_55959141808445_0
timestamp 1707688321
transform 1 0 286 0 1 228
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808446  sky130_fd_pr__nfet_01v8__example_55959141808446_0
timestamp 1707688321
transform -1 0 212 0 -1 1102
box -19 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808447  sky130_fd_pr__nfet_01v8__example_55959141808447_0
timestamp 1707688321
transform 1 0 442 0 1 228
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808447  sky130_fd_pr__nfet_01v8__example_55959141808447_1
timestamp 1707688321
transform 1 0 598 0 1 228
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808585  sky130_fd_pr__nfet_01v8__example_55959141808585_0
timestamp 1707688321
transform -1 0 212 0 1 685
box 100 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808450  sky130_fd_pr__pfet_01v8__example_55959141808450_0
timestamp 1707688321
transform -1 0 705 0 -1 1650
box -1 0 297 1
use sky130_fd_pr__pfet_01v8__example_55959141808451  sky130_fd_pr__pfet_01v8__example_55959141808451_0
timestamp 1707688321
transform 1 0 779 0 -1 1650
box -19 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808457  sky130_fd_pr__pfet_01v8__example_55959141808457_0
timestamp 1707688321
transform 1 0 57 0 -1 1650
box -1 0 297 1
<< properties >>
string GDS_END 22105450
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 22091072
<< end >>
