magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -68 -26 4410 106
<< ndiff >>
rect -42 57 0 80
rect -42 23 -34 57
rect -42 0 0 23
rect 4342 57 4384 80
rect 4376 23 4384 57
rect 4342 0 4384 23
<< ndiffc >>
rect -34 23 0 57
rect 4342 23 4376 57
<< ndiffres >>
rect 0 0 4342 80
<< locali >>
rect -34 57 0 73
rect -34 7 0 23
rect 4342 57 4376 73
rect 4342 7 4376 23
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_0
timestamp 1707688321
transform -1 0 8 0 1 11
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_1
timestamp 1707688321
transform 1 0 4334 0 1 11
box 0 0 1 1
<< properties >>
string GDS_END 78948580
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 78948078
<< end >>
