magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -26 -26 286 2026
<< ndiff >>
rect 0 1950 60 2000
rect 200 1950 260 2000
rect 0 1916 11 1950
rect 45 1916 60 1950
rect 200 1916 215 1950
rect 249 1916 260 1950
rect 0 1882 60 1916
rect 200 1882 260 1916
rect 0 1848 11 1882
rect 45 1848 60 1882
rect 200 1848 215 1882
rect 249 1848 260 1882
rect 0 1814 60 1848
rect 200 1814 260 1848
rect 0 1780 11 1814
rect 45 1780 60 1814
rect 200 1780 215 1814
rect 249 1780 260 1814
rect 0 1746 60 1780
rect 200 1746 260 1780
rect 0 1712 11 1746
rect 45 1712 60 1746
rect 200 1712 215 1746
rect 249 1712 260 1746
rect 0 1678 60 1712
rect 200 1678 260 1712
rect 0 1644 11 1678
rect 45 1644 60 1678
rect 200 1644 215 1678
rect 249 1644 260 1678
rect 0 1610 60 1644
rect 200 1610 260 1644
rect 0 1576 11 1610
rect 45 1576 60 1610
rect 200 1576 215 1610
rect 249 1576 260 1610
rect 0 1542 60 1576
rect 200 1542 260 1576
rect 0 1508 11 1542
rect 45 1508 60 1542
rect 200 1508 215 1542
rect 249 1508 260 1542
rect 0 1474 60 1508
rect 200 1474 260 1508
rect 0 1440 11 1474
rect 45 1440 60 1474
rect 200 1440 215 1474
rect 249 1440 260 1474
rect 0 1406 60 1440
rect 200 1406 260 1440
rect 0 1372 11 1406
rect 45 1372 60 1406
rect 200 1372 215 1406
rect 249 1372 260 1406
rect 0 1338 60 1372
rect 200 1338 260 1372
rect 0 1304 11 1338
rect 45 1304 60 1338
rect 200 1304 215 1338
rect 249 1304 260 1338
rect 0 1270 60 1304
rect 200 1270 260 1304
rect 0 1236 11 1270
rect 45 1236 60 1270
rect 200 1236 215 1270
rect 249 1236 260 1270
rect 0 1202 60 1236
rect 200 1202 260 1236
rect 0 1168 11 1202
rect 45 1168 60 1202
rect 200 1168 215 1202
rect 249 1168 260 1202
rect 0 1134 60 1168
rect 200 1134 260 1168
rect 0 1100 11 1134
rect 45 1100 60 1134
rect 200 1100 215 1134
rect 249 1100 260 1134
rect 0 1066 60 1100
rect 200 1066 260 1100
rect 0 1032 11 1066
rect 45 1032 60 1066
rect 200 1032 215 1066
rect 249 1032 260 1066
rect 0 998 60 1032
rect 200 998 260 1032
rect 0 964 11 998
rect 45 964 60 998
rect 200 964 215 998
rect 249 964 260 998
rect 0 930 60 964
rect 200 930 260 964
rect 0 896 11 930
rect 45 896 60 930
rect 200 896 215 930
rect 249 896 260 930
rect 0 862 60 896
rect 200 862 260 896
rect 0 828 11 862
rect 45 828 60 862
rect 200 828 215 862
rect 249 828 260 862
rect 0 794 60 828
rect 200 794 260 828
rect 0 760 11 794
rect 45 760 60 794
rect 200 760 215 794
rect 249 760 260 794
rect 0 726 60 760
rect 200 726 260 760
rect 0 692 11 726
rect 45 692 60 726
rect 200 692 215 726
rect 249 692 260 726
rect 0 658 60 692
rect 200 658 260 692
rect 0 624 11 658
rect 45 624 60 658
rect 200 624 215 658
rect 249 624 260 658
rect 0 590 60 624
rect 200 590 260 624
rect 0 556 11 590
rect 45 556 60 590
rect 200 556 215 590
rect 249 556 260 590
rect 0 522 60 556
rect 200 522 260 556
rect 0 488 11 522
rect 45 488 60 522
rect 200 488 215 522
rect 249 488 260 522
rect 0 454 60 488
rect 200 454 260 488
rect 0 420 11 454
rect 45 420 60 454
rect 200 420 215 454
rect 249 420 260 454
rect 0 386 60 420
rect 200 386 260 420
rect 0 352 11 386
rect 45 352 60 386
rect 200 352 215 386
rect 249 352 260 386
rect 0 318 60 352
rect 200 318 260 352
rect 0 284 11 318
rect 45 284 60 318
rect 200 284 215 318
rect 249 284 260 318
rect 0 250 60 284
rect 200 250 260 284
rect 0 216 11 250
rect 45 216 60 250
rect 200 216 215 250
rect 249 216 260 250
rect 0 182 60 216
rect 200 182 260 216
rect 0 148 11 182
rect 45 148 60 182
rect 200 148 215 182
rect 249 148 260 182
rect 0 114 60 148
rect 200 114 260 148
rect 0 80 11 114
rect 45 80 60 114
rect 200 80 215 114
rect 249 80 260 114
rect 0 46 60 80
rect 200 46 260 80
rect 0 12 11 46
rect 45 12 60 46
rect 200 12 215 46
rect 249 12 260 46
rect 0 0 60 12
rect 200 0 260 12
<< ndiffc >>
rect 11 1916 45 1950
rect 215 1916 249 1950
rect 11 1848 45 1882
rect 215 1848 249 1882
rect 11 1780 45 1814
rect 215 1780 249 1814
rect 11 1712 45 1746
rect 215 1712 249 1746
rect 11 1644 45 1678
rect 215 1644 249 1678
rect 11 1576 45 1610
rect 215 1576 249 1610
rect 11 1508 45 1542
rect 215 1508 249 1542
rect 11 1440 45 1474
rect 215 1440 249 1474
rect 11 1372 45 1406
rect 215 1372 249 1406
rect 11 1304 45 1338
rect 215 1304 249 1338
rect 11 1236 45 1270
rect 215 1236 249 1270
rect 11 1168 45 1202
rect 215 1168 249 1202
rect 11 1100 45 1134
rect 215 1100 249 1134
rect 11 1032 45 1066
rect 215 1032 249 1066
rect 11 964 45 998
rect 215 964 249 998
rect 11 896 45 930
rect 215 896 249 930
rect 11 828 45 862
rect 215 828 249 862
rect 11 760 45 794
rect 215 760 249 794
rect 11 692 45 726
rect 215 692 249 726
rect 11 624 45 658
rect 215 624 249 658
rect 11 556 45 590
rect 215 556 249 590
rect 11 488 45 522
rect 215 488 249 522
rect 11 420 45 454
rect 215 420 249 454
rect 11 352 45 386
rect 215 352 249 386
rect 11 284 45 318
rect 215 284 249 318
rect 11 216 45 250
rect 215 216 249 250
rect 11 148 45 182
rect 215 148 249 182
rect 11 80 45 114
rect 215 80 249 114
rect 11 12 45 46
rect 215 12 249 46
<< psubdiff >>
rect 60 1950 200 2000
rect 60 1916 113 1950
rect 147 1916 200 1950
rect 60 1882 200 1916
rect 60 1848 113 1882
rect 147 1848 200 1882
rect 60 1814 200 1848
rect 60 1780 113 1814
rect 147 1780 200 1814
rect 60 1746 200 1780
rect 60 1712 113 1746
rect 147 1712 200 1746
rect 60 1678 200 1712
rect 60 1644 113 1678
rect 147 1644 200 1678
rect 60 1610 200 1644
rect 60 1576 113 1610
rect 147 1576 200 1610
rect 60 1542 200 1576
rect 60 1508 113 1542
rect 147 1508 200 1542
rect 60 1474 200 1508
rect 60 1440 113 1474
rect 147 1440 200 1474
rect 60 1406 200 1440
rect 60 1372 113 1406
rect 147 1372 200 1406
rect 60 1338 200 1372
rect 60 1304 113 1338
rect 147 1304 200 1338
rect 60 1270 200 1304
rect 60 1236 113 1270
rect 147 1236 200 1270
rect 60 1202 200 1236
rect 60 1168 113 1202
rect 147 1168 200 1202
rect 60 1134 200 1168
rect 60 1100 113 1134
rect 147 1100 200 1134
rect 60 1066 200 1100
rect 60 1032 113 1066
rect 147 1032 200 1066
rect 60 998 200 1032
rect 60 964 113 998
rect 147 964 200 998
rect 60 930 200 964
rect 60 896 113 930
rect 147 896 200 930
rect 60 862 200 896
rect 60 828 113 862
rect 147 828 200 862
rect 60 794 200 828
rect 60 760 113 794
rect 147 760 200 794
rect 60 726 200 760
rect 60 692 113 726
rect 147 692 200 726
rect 60 658 200 692
rect 60 624 113 658
rect 147 624 200 658
rect 60 590 200 624
rect 60 556 113 590
rect 147 556 200 590
rect 60 522 200 556
rect 60 488 113 522
rect 147 488 200 522
rect 60 454 200 488
rect 60 420 113 454
rect 147 420 200 454
rect 60 386 200 420
rect 60 352 113 386
rect 147 352 200 386
rect 60 318 200 352
rect 60 284 113 318
rect 147 284 200 318
rect 60 250 200 284
rect 60 216 113 250
rect 147 216 200 250
rect 60 182 200 216
rect 60 148 113 182
rect 147 148 200 182
rect 60 114 200 148
rect 60 80 113 114
rect 147 80 200 114
rect 60 46 200 80
rect 60 12 113 46
rect 147 12 200 46
rect 60 0 200 12
<< psubdiffcont >>
rect 113 1916 147 1950
rect 113 1848 147 1882
rect 113 1780 147 1814
rect 113 1712 147 1746
rect 113 1644 147 1678
rect 113 1576 147 1610
rect 113 1508 147 1542
rect 113 1440 147 1474
rect 113 1372 147 1406
rect 113 1304 147 1338
rect 113 1236 147 1270
rect 113 1168 147 1202
rect 113 1100 147 1134
rect 113 1032 147 1066
rect 113 964 147 998
rect 113 896 147 930
rect 113 828 147 862
rect 113 760 147 794
rect 113 692 147 726
rect 113 624 147 658
rect 113 556 147 590
rect 113 488 147 522
rect 113 420 147 454
rect 113 352 147 386
rect 113 284 147 318
rect 113 216 147 250
rect 113 148 147 182
rect 113 80 147 114
rect 113 12 147 46
<< locali >>
rect 11 1950 249 1966
rect 45 1916 113 1950
rect 147 1916 215 1950
rect 11 1882 249 1916
rect 45 1848 113 1882
rect 147 1848 215 1882
rect 11 1814 249 1848
rect 45 1780 113 1814
rect 147 1780 215 1814
rect 11 1746 249 1780
rect 45 1712 113 1746
rect 147 1712 215 1746
rect 11 1678 249 1712
rect 45 1644 113 1678
rect 147 1644 215 1678
rect 11 1610 249 1644
rect 45 1576 113 1610
rect 147 1576 215 1610
rect 11 1542 249 1576
rect 45 1508 113 1542
rect 147 1508 215 1542
rect 11 1474 249 1508
rect 45 1440 113 1474
rect 147 1440 215 1474
rect 11 1406 249 1440
rect 45 1372 113 1406
rect 147 1372 215 1406
rect 11 1338 249 1372
rect 45 1304 113 1338
rect 147 1304 215 1338
rect 11 1270 249 1304
rect 45 1236 113 1270
rect 147 1236 215 1270
rect 11 1202 249 1236
rect 45 1168 113 1202
rect 147 1168 215 1202
rect 11 1134 249 1168
rect 45 1100 113 1134
rect 147 1100 215 1134
rect 11 1066 249 1100
rect 45 1032 113 1066
rect 147 1032 215 1066
rect 11 998 249 1032
rect 45 964 113 998
rect 147 964 215 998
rect 11 930 249 964
rect 45 896 113 930
rect 147 896 215 930
rect 11 862 249 896
rect 45 828 113 862
rect 147 828 215 862
rect 11 794 249 828
rect 45 760 113 794
rect 147 760 215 794
rect 11 726 249 760
rect 45 692 113 726
rect 147 692 215 726
rect 11 658 249 692
rect 45 624 113 658
rect 147 624 215 658
rect 11 590 249 624
rect 45 556 113 590
rect 147 556 215 590
rect 11 522 249 556
rect 45 488 113 522
rect 147 488 215 522
rect 11 454 249 488
rect 45 420 113 454
rect 147 420 215 454
rect 11 386 249 420
rect 45 352 113 386
rect 147 352 215 386
rect 11 318 249 352
rect 45 284 113 318
rect 147 284 215 318
rect 11 250 249 284
rect 45 216 113 250
rect 147 216 215 250
rect 11 182 249 216
rect 45 148 113 182
rect 147 148 215 182
rect 11 114 249 148
rect 45 80 113 114
rect 147 80 215 114
rect 11 46 249 80
rect 45 12 113 46
rect 147 12 215 46
rect 11 -4 249 12
<< properties >>
string GDS_END 34396924
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 34390776
<< end >>
