magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect 5489 1660 7123 1893
rect 9693 1660 11327 1890
<< pwell >>
rect 10427 690 10521 778
rect 1432 243 2189 294
rect 3113 243 11360 294
rect 1432 72 11360 243
<< pdiff >>
rect 285 4080 493 4109
rect 545 1164 571 1200
rect 1221 1164 1247 1200
rect 545 1066 571 1102
rect 1221 1066 1247 1102
<< psubdiff >>
rect 3615 265 3765 268
rect 1458 217 2163 265
rect 3139 234 3765 265
rect 3799 234 3834 268
rect 3868 234 3903 268
rect 3937 234 3972 268
rect 4006 234 4041 268
rect 4075 234 4110 268
rect 4144 234 4179 268
rect 4213 234 4248 268
rect 4282 234 4317 268
rect 4351 234 4386 268
rect 4420 234 4455 268
rect 4489 234 4524 268
rect 4558 234 4593 268
rect 4627 234 4662 268
rect 4696 234 4731 268
rect 4765 234 4800 268
rect 4834 234 4869 268
rect 4903 234 4938 268
rect 4972 234 5007 268
rect 5041 234 5076 268
rect 5110 234 5145 268
rect 5179 234 5214 268
rect 5248 234 5283 268
rect 5317 234 5352 268
rect 5386 234 5421 268
rect 5455 234 5490 268
rect 5524 234 5559 268
rect 5593 234 5628 268
rect 5662 234 5697 268
rect 5731 234 5766 268
rect 5800 234 5835 268
rect 5869 234 5904 268
rect 3139 217 5904 234
rect 1458 200 5904 217
rect 1458 166 3765 200
rect 3799 166 3834 200
rect 3868 166 3903 200
rect 3937 166 3972 200
rect 4006 166 4041 200
rect 4075 166 4110 200
rect 4144 166 4179 200
rect 4213 166 4248 200
rect 4282 166 4317 200
rect 4351 166 4386 200
rect 4420 166 4455 200
rect 4489 166 4524 200
rect 4558 166 4593 200
rect 4627 166 4662 200
rect 4696 166 4731 200
rect 4765 166 4800 200
rect 4834 166 4869 200
rect 4903 166 4938 200
rect 4972 166 5007 200
rect 5041 166 5076 200
rect 5110 166 5145 200
rect 5179 166 5214 200
rect 5248 166 5283 200
rect 5317 166 5352 200
rect 5386 166 5421 200
rect 5455 166 5490 200
rect 5524 166 5559 200
rect 5593 166 5628 200
rect 5662 166 5697 200
rect 5731 166 5766 200
rect 5800 166 5835 200
rect 5869 166 5904 200
rect 1458 132 5904 166
rect 1458 98 1482 132
rect 1516 98 1550 132
rect 1584 98 1618 132
rect 1652 98 1686 132
rect 1720 98 1754 132
rect 1788 98 1822 132
rect 1856 98 1890 132
rect 1924 98 1958 132
rect 1992 98 2026 132
rect 2060 98 2094 132
rect 2128 98 2162 132
rect 2196 98 2230 132
rect 2264 98 2298 132
rect 2332 98 2366 132
rect 2400 98 2434 132
rect 2468 98 2502 132
rect 2536 98 2570 132
rect 2604 98 2638 132
rect 2672 98 2707 132
rect 2741 98 2776 132
rect 2810 98 2845 132
rect 2879 98 2914 132
rect 2948 98 2983 132
rect 3017 98 3052 132
rect 3086 98 3121 132
rect 3155 98 3190 132
rect 3224 98 3259 132
rect 3293 98 3328 132
rect 3362 98 3397 132
rect 3431 98 3466 132
rect 3500 98 3535 132
rect 3569 98 3604 132
rect 3638 98 3673 132
rect 3707 98 3765 132
rect 3799 98 3834 132
rect 3868 98 3903 132
rect 3937 98 3972 132
rect 4006 98 4041 132
rect 4075 98 4110 132
rect 4144 98 4179 132
rect 4213 98 4248 132
rect 4282 98 4317 132
rect 4351 98 4386 132
rect 4420 98 4455 132
rect 4489 98 4524 132
rect 4558 98 4593 132
rect 4627 98 4662 132
rect 4696 98 4731 132
rect 4765 98 4800 132
rect 4834 98 4869 132
rect 4903 98 4938 132
rect 4972 98 5007 132
rect 5041 98 5076 132
rect 5110 98 5145 132
rect 5179 98 5214 132
rect 5248 98 5283 132
rect 5317 98 5352 132
rect 5386 98 5421 132
rect 5455 98 5490 132
rect 5524 98 5559 132
rect 5593 98 5628 132
rect 5662 98 5697 132
rect 5731 98 5766 132
rect 5800 98 5835 132
rect 5869 98 5904 132
rect 11310 98 11334 268
<< psubdiffcont >>
rect 3765 234 3799 268
rect 3834 234 3868 268
rect 3903 234 3937 268
rect 3972 234 4006 268
rect 4041 234 4075 268
rect 4110 234 4144 268
rect 4179 234 4213 268
rect 4248 234 4282 268
rect 4317 234 4351 268
rect 4386 234 4420 268
rect 4455 234 4489 268
rect 4524 234 4558 268
rect 4593 234 4627 268
rect 4662 234 4696 268
rect 4731 234 4765 268
rect 4800 234 4834 268
rect 4869 234 4903 268
rect 4938 234 4972 268
rect 5007 234 5041 268
rect 5076 234 5110 268
rect 5145 234 5179 268
rect 5214 234 5248 268
rect 5283 234 5317 268
rect 5352 234 5386 268
rect 5421 234 5455 268
rect 5490 234 5524 268
rect 5559 234 5593 268
rect 5628 234 5662 268
rect 5697 234 5731 268
rect 5766 234 5800 268
rect 5835 234 5869 268
rect 3765 166 3799 200
rect 3834 166 3868 200
rect 3903 166 3937 200
rect 3972 166 4006 200
rect 4041 166 4075 200
rect 4110 166 4144 200
rect 4179 166 4213 200
rect 4248 166 4282 200
rect 4317 166 4351 200
rect 4386 166 4420 200
rect 4455 166 4489 200
rect 4524 166 4558 200
rect 4593 166 4627 200
rect 4662 166 4696 200
rect 4731 166 4765 200
rect 4800 166 4834 200
rect 4869 166 4903 200
rect 4938 166 4972 200
rect 5007 166 5041 200
rect 5076 166 5110 200
rect 5145 166 5179 200
rect 5214 166 5248 200
rect 5283 166 5317 200
rect 5352 166 5386 200
rect 5421 166 5455 200
rect 5490 166 5524 200
rect 5559 166 5593 200
rect 5628 166 5662 200
rect 5697 166 5731 200
rect 5766 166 5800 200
rect 5835 166 5869 200
rect 1482 98 1516 132
rect 1550 98 1584 132
rect 1618 98 1652 132
rect 1686 98 1720 132
rect 1754 98 1788 132
rect 1822 98 1856 132
rect 1890 98 1924 132
rect 1958 98 1992 132
rect 2026 98 2060 132
rect 2094 98 2128 132
rect 2162 98 2196 132
rect 2230 98 2264 132
rect 2298 98 2332 132
rect 2366 98 2400 132
rect 2434 98 2468 132
rect 2502 98 2536 132
rect 2570 98 2604 132
rect 2638 98 2672 132
rect 2707 98 2741 132
rect 2776 98 2810 132
rect 2845 98 2879 132
rect 2914 98 2948 132
rect 2983 98 3017 132
rect 3052 98 3086 132
rect 3121 98 3155 132
rect 3190 98 3224 132
rect 3259 98 3293 132
rect 3328 98 3362 132
rect 3397 98 3431 132
rect 3466 98 3500 132
rect 3535 98 3569 132
rect 3604 98 3638 132
rect 3673 98 3707 132
rect 3765 98 3799 132
rect 3834 98 3868 132
rect 3903 98 3937 132
rect 3972 98 4006 132
rect 4041 98 4075 132
rect 4110 98 4144 132
rect 4179 98 4213 132
rect 4248 98 4282 132
rect 4317 98 4351 132
rect 4386 98 4420 132
rect 4455 98 4489 132
rect 4524 98 4558 132
rect 4593 98 4627 132
rect 4662 98 4696 132
rect 4731 98 4765 132
rect 4800 98 4834 132
rect 4869 98 4903 132
rect 4938 98 4972 132
rect 5007 98 5041 132
rect 5076 98 5110 132
rect 5145 98 5179 132
rect 5214 98 5248 132
rect 5283 98 5317 132
rect 5352 98 5386 132
rect 5421 98 5455 132
rect 5490 98 5524 132
rect 5559 98 5593 132
rect 5628 98 5662 132
rect 5697 98 5731 132
rect 5766 98 5800 132
rect 5835 98 5869 132
rect 5904 98 11310 268
<< locali >>
rect -17 3195 17 3233
rect -17 3123 17 3161
rect 615 3195 649 3233
rect 615 3123 649 3161
rect 1579 3195 1613 3233
rect 1579 3123 1613 3161
rect 2591 3195 2625 3233
rect 2591 3123 2625 3161
rect 3555 3195 3589 3233
rect 3555 3123 3589 3161
rect 4819 3195 4853 3233
rect 4819 3123 4853 3161
rect 5783 3195 5817 3233
rect 5783 3123 5817 3161
rect 6795 3195 6829 3233
rect 6795 3123 6829 3161
rect 7759 3195 7793 3233
rect 7759 3123 7793 3161
rect 8391 3195 8425 3233
rect 8391 3123 8425 3161
rect 9023 3195 9057 3233
rect 9023 3123 9057 3161
rect 9987 3195 10021 3233
rect 9987 3123 10021 3161
rect 10999 3195 11033 3233
rect 10999 3123 11033 3161
rect 11963 3195 11997 3233
rect 11963 3123 11997 3161
rect 14983 3195 15017 3233
rect 14983 3123 15017 3161
rect 342 2204 376 2242
rect 3842 2204 3876 2242
rect 4532 2204 4566 2242
rect 8046 2204 8080 2242
rect 8736 2204 8770 2242
rect 12250 2204 12284 2242
rect 8041 1722 8079 1756
rect 8007 1626 8113 1722
rect 8458 1644 8573 1682
rect 765 1586 803 1620
rect 837 1586 875 1620
rect 909 1586 947 1620
rect 981 1586 1019 1620
rect 1053 1586 1055 1620
rect 737 1540 771 1586
rect 1021 1540 1055 1586
rect 8231 1594 8265 1644
rect 519 814 629 1050
rect 879 1000 913 1066
rect 1163 814 1273 1050
rect 1628 734 1803 944
rect 3483 734 3629 944
rect 4044 890 4183 1532
rect 8231 1510 8265 1560
rect 8231 1426 8265 1476
rect 4501 956 4535 990
rect 4853 956 4887 990
rect 5205 956 5239 990
rect 5557 956 5591 990
rect 5909 956 5943 990
rect 6261 956 6295 990
rect 6613 956 6647 990
rect 6965 956 6999 990
rect 7317 956 7351 990
rect 7669 956 7703 990
rect 8307 956 8341 990
rect 1628 426 1871 734
rect 2233 416 2349 734
rect 2971 416 3053 734
rect 3415 426 3629 734
rect 4044 444 4183 746
rect 4501 654 4535 700
rect 4853 654 4887 700
rect 5205 654 5239 700
rect 5557 654 5591 700
rect 5909 654 5943 700
rect 6261 654 6295 700
rect 6613 654 6647 700
rect 7317 654 7351 700
rect 7669 654 7703 700
rect 3674 234 3765 268
rect 3799 234 3834 268
rect 3868 234 3903 268
rect 3937 234 3972 268
rect 4006 234 4041 268
rect 4075 234 4110 268
rect 4144 234 4179 268
rect 4213 234 4248 268
rect 4282 234 4317 268
rect 4351 234 4386 268
rect 4420 234 4455 268
rect 4489 234 4524 268
rect 4558 234 4593 268
rect 4627 234 4662 268
rect 4696 234 4731 268
rect 4765 234 4800 268
rect 4834 234 4869 268
rect 4903 234 4938 268
rect 4972 234 5007 268
rect 5041 234 5076 268
rect 5110 234 5145 268
rect 5179 234 5214 268
rect 5248 234 5283 268
rect 5317 234 5352 268
rect 5386 234 5421 268
rect 5455 234 5490 268
rect 5524 234 5559 268
rect 5593 234 5628 268
rect 5662 234 5697 268
rect 5731 234 5766 268
rect 5800 234 5835 268
rect 5869 234 5904 268
rect 3674 225 5904 234
rect 1458 200 5904 225
rect 1458 166 3765 200
rect 3799 166 3834 200
rect 3868 166 3903 200
rect 3937 166 3972 200
rect 4006 166 4041 200
rect 4075 166 4110 200
rect 4144 166 4179 200
rect 4213 166 4248 200
rect 4282 166 4317 200
rect 4351 166 4386 200
rect 4420 166 4455 200
rect 4489 166 4524 200
rect 4558 166 4593 200
rect 4627 166 4662 200
rect 4696 166 4731 200
rect 4765 166 4800 200
rect 4834 166 4869 200
rect 4903 166 4938 200
rect 4972 166 5007 200
rect 5041 166 5076 200
rect 5110 166 5145 200
rect 5179 166 5214 200
rect 5248 166 5283 200
rect 5317 166 5352 200
rect 5386 166 5421 200
rect 5455 166 5490 200
rect 5524 166 5559 200
rect 5593 166 5628 200
rect 5662 166 5697 200
rect 5731 166 5766 200
rect 5800 166 5835 200
rect 5869 166 5904 200
rect 1458 132 5904 166
rect 1458 98 1482 132
rect 1516 98 1550 132
rect 1584 98 1618 132
rect 1652 98 1686 132
rect 1720 98 1754 132
rect 1788 98 1822 132
rect 1856 98 1890 132
rect 1924 98 1958 132
rect 1992 98 2026 132
rect 2060 98 2094 132
rect 2128 98 2162 132
rect 2196 98 2230 132
rect 2264 98 2298 132
rect 2332 98 2366 132
rect 2400 98 2434 132
rect 2468 98 2502 132
rect 2536 98 2570 132
rect 2604 98 2638 132
rect 2672 98 2707 132
rect 2741 98 2776 132
rect 2810 98 2845 132
rect 2879 98 2914 132
rect 2948 98 2983 132
rect 3017 98 3052 132
rect 3086 98 3121 132
rect 3155 98 3190 132
rect 3224 98 3259 132
rect 3293 98 3328 132
rect 3362 98 3397 132
rect 3431 98 3466 132
rect 3500 98 3535 132
rect 3569 98 3604 132
rect 3638 98 3673 132
rect 3707 98 3765 132
rect 3799 98 3834 132
rect 3868 98 3903 132
rect 3937 98 3972 132
rect 4006 98 4041 132
rect 4075 98 4110 132
rect 4144 98 4179 132
rect 4213 98 4248 132
rect 4282 98 4317 132
rect 4351 98 4386 132
rect 4420 98 4455 132
rect 4489 98 4524 132
rect 4558 98 4593 132
rect 4627 98 4662 132
rect 4696 98 4731 132
rect 4765 98 4800 132
rect 4834 98 4869 132
rect 4903 98 4938 132
rect 4972 98 5007 132
rect 5041 98 5076 132
rect 5110 98 5145 132
rect 5179 98 5214 132
rect 5248 98 5283 132
rect 5317 98 5352 132
rect 5386 98 5421 132
rect 5455 98 5490 132
rect 5524 98 5559 132
rect 5593 98 5628 132
rect 5662 98 5697 132
rect 5731 98 5766 132
rect 5800 98 5835 132
rect 5869 98 5904 132
rect 11310 98 11334 268
<< viali >>
rect -17 3233 17 3267
rect -17 3161 17 3195
rect -17 3089 17 3123
rect 615 3233 649 3267
rect 615 3161 649 3195
rect 615 3089 649 3123
rect 1579 3233 1613 3267
rect 1579 3161 1613 3195
rect 1579 3089 1613 3123
rect 2591 3233 2625 3267
rect 2591 3161 2625 3195
rect 2591 3089 2625 3123
rect 3555 3233 3589 3267
rect 3555 3161 3589 3195
rect 3555 3089 3589 3123
rect 4819 3233 4853 3267
rect 4819 3161 4853 3195
rect 4819 3089 4853 3123
rect 5783 3233 5817 3267
rect 5783 3161 5817 3195
rect 5783 3089 5817 3123
rect 6795 3233 6829 3267
rect 6795 3161 6829 3195
rect 6795 3089 6829 3123
rect 7759 3233 7793 3267
rect 7759 3161 7793 3195
rect 7759 3089 7793 3123
rect 8391 3233 8425 3267
rect 8391 3161 8425 3195
rect 8391 3089 8425 3123
rect 9023 3233 9057 3267
rect 9023 3161 9057 3195
rect 9023 3089 9057 3123
rect 9987 3233 10021 3267
rect 9987 3161 10021 3195
rect 9987 3089 10021 3123
rect 10999 3233 11033 3267
rect 10999 3161 11033 3195
rect 10999 3089 11033 3123
rect 11963 3233 11997 3267
rect 11963 3161 11997 3195
rect 11963 3089 11997 3123
rect 14983 3233 15017 3267
rect 14983 3161 15017 3195
rect 14983 3089 15017 3123
rect 342 2242 376 2276
rect 342 2170 376 2204
rect 3842 2242 3876 2276
rect 3842 2170 3876 2204
rect 4532 2242 4566 2276
rect 4532 2170 4566 2204
rect 8046 2242 8080 2276
rect 8046 2170 8080 2204
rect 8736 2242 8770 2276
rect 8736 2170 8770 2204
rect 12250 2242 12284 2276
rect 12250 2170 12284 2204
rect 8007 1722 8041 1756
rect 8079 1722 8113 1756
rect 8231 1644 8265 1678
rect 731 1586 765 1620
rect 803 1586 837 1620
rect 875 1586 909 1620
rect 947 1586 981 1620
rect 1019 1586 1053 1620
rect 8231 1560 8265 1594
rect 8231 1476 8265 1510
rect 8231 1392 8265 1426
<< metal1 >>
rect 126 3954 132 4070
rect 312 3954 318 4070
rect 6244 4018 6250 4070
rect 6302 4018 6328 4070
rect 6380 4018 6405 4070
rect 6457 4018 6482 4070
rect 6534 4018 6559 4070
rect 6611 4018 6617 4070
rect 6244 3996 6617 4018
rect 6244 3944 6250 3996
rect 6302 3944 6328 3996
rect 6380 3944 6405 3996
rect 6457 3944 6482 3996
rect 6534 3944 6559 3996
rect 6611 3944 6617 3996
rect 10451 4069 10767 4070
rect 10451 4017 10457 4069
rect 10509 4017 10541 4069
rect 10593 4017 10625 4069
rect 10677 4017 10709 4069
rect 10761 4017 10767 4069
rect 10451 4005 10767 4017
rect 10451 3953 10457 4005
rect 10509 3953 10541 4005
rect 10593 3953 10625 4005
rect 10677 3953 10709 4005
rect 10761 3953 10767 4005
rect 10451 3952 10767 3953
rect 10951 4069 11267 4070
rect 10951 4017 10957 4069
rect 11009 4017 11041 4069
rect 11093 4017 11125 4069
rect 11177 4017 11209 4069
rect 11261 4017 11267 4069
rect 10951 4005 11267 4017
rect 10951 3953 10957 4005
rect 11009 3953 11041 4005
rect 11093 3953 11125 4005
rect 11177 3953 11209 4005
rect 11261 3953 11267 4005
rect 10951 3952 11267 3953
rect 6244 3922 6617 3944
rect 6244 3870 6250 3922
rect 6302 3870 6328 3922
rect 6380 3870 6405 3922
rect 6457 3870 6482 3922
rect 6534 3870 6559 3922
rect 6611 3870 6617 3922
rect 6244 3848 6617 3870
rect 6244 3796 6250 3848
rect 6302 3796 6328 3848
rect 6380 3796 6405 3848
rect 6457 3796 6482 3848
rect 6534 3796 6559 3848
rect 6611 3796 6617 3848
rect 6244 3774 6617 3796
rect 6244 3722 6250 3774
rect 6302 3722 6328 3774
rect 6380 3722 6405 3774
rect 6457 3722 6482 3774
rect 6534 3722 6559 3774
rect 6611 3722 6617 3774
rect 1364 3608 5620 3614
rect 1416 3577 5620 3608
rect 1416 3556 1419 3577
rect 1364 3554 1419 3556
tri 1419 3554 1442 3577 nw
tri 5543 3554 5566 3577 ne
rect 5566 3554 5620 3577
rect 1364 3544 1416 3554
tri 1416 3551 1419 3554 nw
tri 5566 3552 5568 3554 ne
rect 5568 3548 5620 3554
rect 5648 3502 5654 3554
rect 5706 3502 5718 3554
rect 5770 3517 10886 3554
rect 5770 3502 5776 3517
tri 5776 3502 5791 3517 nw
tri 10865 3502 10880 3517 ne
rect 10880 3502 10886 3517
rect 10938 3502 10950 3554
rect 11002 3502 11008 3554
rect 1364 3486 1416 3492
rect 132 3429 223 3435
rect 132 3377 171 3429
rect 2003 3429 2055 3435
rect 132 3365 223 3377
rect 132 3336 171 3365
tri 223 3353 248 3378 sw
tri 1978 3353 2003 3378 se
rect 2003 3365 2055 3377
rect 171 3307 223 3313
tri 2055 3359 2080 3384 sw
rect 2003 3307 2055 3313
rect -48 3267 34 3279
rect 609 3273 655 3279
rect -48 3233 -17 3267
rect 17 3233 34 3267
rect -48 3195 34 3233
rect -48 3161 -17 3195
rect 17 3161 34 3195
rect -48 3123 34 3161
rect -48 3089 -17 3123
rect 17 3089 34 3123
rect -48 3077 34 3089
rect 436 3267 552 3273
rect 436 3081 552 3087
rect 597 3267 655 3273
rect 649 3215 655 3267
rect 597 3203 655 3215
rect 649 3151 655 3203
rect 597 3139 655 3151
rect 649 3087 655 3139
rect 597 3081 655 3087
rect 609 3077 655 3081
rect 1573 3267 1619 3279
rect 1573 3233 1579 3267
rect 1613 3233 1619 3267
rect 1573 3195 1619 3233
rect 1573 3161 1579 3195
rect 1613 3161 1619 3195
rect 1573 3123 1619 3161
rect 1573 3089 1579 3123
rect 1613 3089 1619 3123
rect 1573 3077 1619 3089
rect 2585 3267 2631 3279
rect 2585 3233 2591 3267
rect 2625 3233 2631 3267
rect 2585 3195 2631 3233
rect 2585 3161 2591 3195
rect 2625 3161 2631 3195
rect 2585 3123 2631 3161
rect 2585 3089 2591 3123
rect 2625 3089 2631 3123
rect 2585 3077 2631 3089
rect 3549 3267 3595 3279
rect 3549 3233 3555 3267
rect 3589 3233 3595 3267
rect 3549 3195 3595 3233
rect 3549 3161 3555 3195
rect 3589 3161 3595 3195
rect 3549 3123 3595 3161
rect 3549 3089 3555 3123
rect 3589 3089 3595 3123
rect 3549 3077 3595 3089
rect 4416 3268 4532 3274
rect 4416 3082 4532 3088
rect 4813 3267 4859 3279
rect 4813 3233 4819 3267
rect 4853 3233 4859 3267
rect 4813 3195 4859 3233
rect 4813 3161 4819 3195
rect 4853 3161 4859 3195
rect 4813 3123 4859 3161
rect 4813 3089 4819 3123
rect 4853 3089 4859 3123
rect 4813 3077 4859 3089
rect 5777 3267 5823 3279
rect 5777 3233 5783 3267
rect 5817 3233 5823 3267
rect 5777 3195 5823 3233
rect 5777 3161 5783 3195
rect 5817 3161 5823 3195
rect 5777 3123 5823 3161
rect 5777 3089 5783 3123
rect 5817 3089 5823 3123
rect 5777 3077 5823 3089
rect 6789 3267 6835 3279
rect 6789 3233 6795 3267
rect 6829 3233 6835 3267
rect 6789 3195 6835 3233
rect 6789 3161 6795 3195
rect 6829 3161 6835 3195
rect 6789 3123 6835 3161
rect 6789 3089 6795 3123
rect 6829 3089 6835 3123
rect 6789 3077 6835 3089
rect 7753 3267 7799 3279
rect 7753 3233 7759 3267
rect 7793 3233 7799 3267
rect 7753 3195 7799 3233
rect 7753 3161 7759 3195
rect 7793 3161 7799 3195
rect 7753 3123 7799 3161
rect 7753 3089 7759 3123
rect 7793 3089 7799 3123
rect 7753 3077 7799 3089
rect 8385 3267 8431 3279
rect 8385 3233 8391 3267
rect 8425 3233 8431 3267
rect 8385 3195 8431 3233
rect 8385 3161 8391 3195
rect 8425 3161 8431 3195
rect 8385 3123 8431 3161
rect 8385 3089 8391 3123
rect 8425 3089 8431 3123
rect 8385 3077 8431 3089
rect 9017 3267 9063 3279
rect 9017 3233 9023 3267
rect 9057 3233 9063 3267
rect 9017 3195 9063 3233
rect 9017 3161 9023 3195
rect 9057 3161 9063 3195
rect 9017 3123 9063 3161
rect 9017 3089 9023 3123
rect 9057 3089 9063 3123
rect 9017 3077 9063 3089
rect 9981 3267 10027 3279
rect 9981 3233 9987 3267
rect 10021 3233 10027 3267
rect 9981 3195 10027 3233
rect 9981 3161 9987 3195
rect 10021 3161 10027 3195
rect 9981 3123 10027 3161
rect 9981 3089 9987 3123
rect 10021 3089 10027 3123
rect 9981 3077 10027 3089
rect 10993 3267 11039 3279
rect 10993 3233 10999 3267
rect 11033 3233 11039 3267
rect 10993 3195 11039 3233
rect 10993 3161 10999 3195
rect 11033 3161 11039 3195
rect 10993 3123 11039 3161
rect 10993 3089 10999 3123
rect 11033 3089 11039 3123
rect 10993 3077 11039 3089
rect 11957 3267 12003 3279
rect 11957 3233 11963 3267
rect 11997 3233 12003 3267
rect 11957 3195 12003 3233
rect 11957 3161 11963 3195
rect 11997 3161 12003 3195
rect 11957 3123 12003 3161
rect 11957 3089 11963 3123
rect 11997 3089 12003 3123
rect 11957 3077 12003 3089
rect 12612 3077 12646 3279
rect 13766 3273 14010 3279
rect 13818 3221 13830 3273
rect 13882 3221 13894 3273
rect 13946 3221 13958 3273
rect 13766 3201 14010 3221
rect 13818 3149 13830 3201
rect 13882 3149 13894 3201
rect 13946 3149 13958 3201
rect 13766 3128 14010 3149
rect -48 3076 13766 3077
rect 13818 3076 13830 3128
rect 13882 3076 13894 3128
rect 13946 3076 13958 3128
rect 14680 3077 14714 3279
rect 14739 3267 15048 3279
rect 14739 3233 14983 3267
rect 15017 3233 15048 3267
rect 14739 3195 15048 3233
rect 14739 3161 14983 3195
rect 15017 3161 15048 3195
rect 14739 3123 15048 3161
rect 14739 3089 14983 3123
rect 15017 3089 15048 3123
rect 14739 3077 15048 3089
rect 14010 3076 15048 3077
rect -48 3055 15048 3076
rect -48 3049 13766 3055
rect 3981 2997 3987 3049
rect 4039 2997 4051 3049
rect 4103 2997 4115 3049
rect 4167 2997 4179 3049
rect 4231 2997 4243 3049
rect 4295 2997 4301 3049
rect 11148 2997 11154 3049
rect 11206 2997 11218 3049
rect 11270 2997 11276 3049
rect 12464 2997 12470 3049
rect 12522 2997 12534 3049
rect 12586 2997 12598 3049
rect 12650 2997 12662 3049
rect 12714 2997 12726 3049
rect 12778 2997 12784 3049
rect 13818 3003 13830 3055
rect 13882 3003 13894 3055
rect 13946 3003 13958 3055
rect 14010 3049 15048 3055
rect 13766 2997 14010 3003
rect 54 2929 175 2935
rect 54 2877 91 2929
rect 143 2877 175 2929
rect 3555 2917 3561 2969
rect 3613 2917 3625 2969
rect 3677 2940 4113 2969
rect 3677 2935 3701 2940
tri 3701 2935 3706 2940 nw
tri 4004 2935 4009 2940 ne
rect 4009 2935 4113 2940
tri 4113 2935 4147 2969 sw
rect 3677 2917 3683 2935
tri 3683 2917 3701 2935 nw
tri 4009 2917 4027 2935 ne
rect 4027 2931 4147 2935
tri 4261 2941 4289 2969 se
rect 4289 2963 4379 2969
rect 4289 2941 4327 2963
rect 4027 2917 4029 2931
tri 4027 2915 4029 2917 ne
rect 54 2865 175 2877
rect 54 2813 91 2865
rect 143 2813 175 2865
rect 4261 2911 4327 2941
tri 8465 2935 8499 2969 se
rect 8499 2940 9373 2969
rect 8499 2935 8603 2940
tri 8603 2935 8608 2940 nw
tri 9344 2935 9349 2940 ne
rect 9349 2935 9373 2940
rect 4261 2899 4379 2911
rect 4261 2847 4327 2899
rect 6596 2881 6602 2933
rect 6654 2881 6666 2933
rect 6718 2881 6724 2933
rect 8264 2929 8316 2935
rect 8583 2917 8585 2935
tri 8585 2917 8603 2935 nw
tri 9349 2917 9367 2935 ne
rect 9367 2917 9373 2935
rect 9425 2917 9437 2969
rect 9489 2917 9495 2969
rect 11614 2917 11620 2969
rect 11672 2917 11684 2969
rect 11736 2954 12540 2969
tri 12540 2954 12555 2969 sw
rect 11736 2940 12555 2954
rect 11736 2935 11760 2940
tri 11760 2935 11765 2940 nw
tri 12412 2935 12417 2940 ne
rect 12417 2935 12555 2940
tri 12669 2954 12684 2969 se
rect 12684 2954 13552 2969
rect 12669 2940 13552 2954
rect 12669 2935 12789 2940
rect 11736 2917 11742 2935
tri 11742 2917 11760 2935 nw
tri 12417 2917 12435 2935 ne
rect 12435 2917 12437 2935
tri 8583 2915 8585 2917 nw
tri 12435 2915 12437 2917 ne
rect 12479 2887 12513 2921
rect 12695 2890 12764 2925
rect 12787 2917 12789 2935
tri 12789 2917 12812 2940 nw
tri 13523 2917 13546 2940 ne
rect 13546 2917 13552 2940
rect 13604 2917 13616 2969
rect 13668 2917 13674 2969
tri 12787 2915 12789 2917 nw
tri 8239 2852 8264 2877 ne
rect 8264 2865 8316 2877
rect 4261 2841 4379 2847
rect 54 2807 175 2813
tri 8316 2852 8341 2877 nw
rect 8264 2807 8316 2813
rect 12464 2727 12470 2779
rect 12522 2727 12534 2779
rect 12586 2727 12598 2779
rect 12650 2727 12662 2779
rect 12714 2727 12726 2779
rect 12778 2727 12784 2779
rect 1680 2617 1732 2623
rect 2316 2617 2368 2623
rect 1680 2553 1732 2565
tri 1732 2541 1757 2566 sw
rect 2760 2619 2920 2625
rect 2760 2567 2868 2619
rect 2316 2553 2368 2565
rect 1680 2495 1732 2501
tri 2368 2541 2393 2566 sw
rect 2760 2555 2920 2567
rect 2368 2501 2373 2541
rect 2316 2495 2373 2501
rect 2760 2503 2868 2555
rect 2760 2494 2920 2503
rect 5884 2617 5936 2623
rect 6676 2617 6728 2623
rect 5884 2553 5936 2565
tri 5936 2541 5961 2566 sw
tri 6651 2541 6676 2566 se
rect 6676 2553 6728 2565
rect 5884 2495 5936 2501
rect 6676 2495 6728 2501
rect 10088 2617 10140 2623
rect 10662 2617 10714 2623
rect 10088 2553 10140 2565
tri 10140 2541 10165 2566 sw
rect 11180 2617 11356 2625
rect 10662 2553 10714 2565
rect 10088 2495 10140 2501
tri 10714 2541 10756 2583 sw
rect 11180 2565 11304 2617
rect 11180 2553 11356 2565
rect 10714 2501 10781 2541
rect 10831 2501 10865 2535
rect 11180 2501 11304 2553
rect 10662 2495 10781 2501
rect 11180 2494 11356 2501
rect 11418 2541 11470 2547
rect 11418 2477 11470 2489
tri 9357 2465 9363 2471 se
rect 9363 2419 9369 2471
rect 9421 2419 9433 2471
rect 9485 2419 9491 2471
tri 9491 2465 9497 2471 sw
rect 11418 2419 11470 2425
rect 2792 2328 2798 2380
rect 2850 2328 2862 2380
rect 2914 2328 11393 2380
rect 11445 2328 11457 2380
rect 11509 2328 11515 2380
rect 0 2158 34 2288
rect 336 2287 382 2288
rect 336 2281 398 2287
rect 336 2276 346 2281
rect 336 2242 342 2276
rect 336 2229 346 2242
rect 336 2217 398 2229
rect 336 2204 346 2217
rect 336 2170 342 2204
rect 336 2165 346 2170
rect 336 2159 398 2165
rect 597 2281 649 2287
rect 2552 2280 2668 2286
rect 597 2217 649 2229
rect 597 2159 649 2165
rect 1444 2161 1450 2277
rect 1566 2161 1572 2277
rect 336 2158 382 2159
rect 2552 2158 2668 2164
rect 3836 2276 3882 2288
rect 3836 2242 3842 2276
rect 3876 2242 3882 2276
rect 3836 2204 3882 2242
rect 3836 2170 3842 2204
rect 3876 2170 3882 2204
rect 3836 2158 3882 2170
rect 4526 2276 4572 2288
rect 4526 2242 4532 2276
rect 4566 2242 4572 2276
rect 4526 2204 4572 2242
rect 4526 2170 4532 2204
rect 4566 2170 4572 2204
rect 4526 2158 4572 2170
rect 4805 2166 4811 2282
rect 4927 2166 4933 2282
rect 5348 2166 5354 2282
rect 5534 2166 5540 2282
rect 8040 2276 8086 2288
rect 8730 2287 8776 2288
rect 8730 2281 8806 2287
rect 8040 2242 8046 2276
rect 8080 2242 8086 2276
rect 8040 2204 8086 2242
rect 8040 2170 8046 2204
rect 8080 2170 8086 2204
rect 8040 2158 8086 2170
rect 8344 2165 8350 2281
rect 8466 2165 8472 2281
rect 8730 2276 8754 2281
rect 8730 2242 8736 2276
rect 8730 2229 8754 2242
rect 8730 2217 8806 2229
rect 8730 2204 8754 2217
rect 8730 2170 8736 2204
rect 8730 2165 8754 2170
rect 8730 2159 8806 2165
rect 9599 2281 9715 2287
rect 9599 2159 9715 2165
rect 12244 2276 12290 2288
rect 12244 2242 12250 2276
rect 12284 2242 12290 2276
rect 12244 2204 12290 2242
rect 12244 2170 12250 2204
rect 12284 2170 12290 2204
rect 8730 2158 8776 2159
rect 12244 2158 12290 2170
rect 12850 2158 12898 2288
rect 13428 2172 13434 2288
rect 13550 2172 13556 2288
rect 13790 2165 13796 2281
rect 13976 2165 13982 2281
rect 14680 2158 14714 2288
rect 14966 2158 15000 2288
rect 0 1928 34 2130
rect 5660 2114 5776 2120
rect 5660 1928 5776 1934
rect 6756 2114 6872 2120
rect 6756 1928 6872 1934
rect 9110 2114 9226 2120
rect 9110 1928 9226 1934
rect 11040 2114 11156 2120
rect 11040 1928 11156 1934
rect 14737 1928 15000 2130
rect 926 1894 978 1900
rect 1680 1894 1732 1900
tri 978 1853 1003 1878 sw
tri 1655 1853 1680 1878 se
rect 978 1842 1680 1853
rect 926 1830 1732 1842
rect 978 1778 1680 1830
rect 926 1772 1732 1778
rect 11211 1894 11463 1900
rect 11263 1842 11411 1894
rect 11211 1830 11463 1842
rect 11263 1778 11411 1830
rect 7976 1725 7982 1777
rect 8034 1756 8046 1777
rect 8098 1756 8125 1777
rect 11211 1772 11463 1778
rect 8041 1725 8046 1756
rect 7976 1722 8007 1725
rect 8041 1722 8079 1725
rect 8113 1722 8125 1756
rect 7976 1716 8125 1722
rect 2316 1699 2368 1705
tri 5437 1678 5447 1688 se
rect 5447 1678 7826 1688
rect 2316 1636 2368 1647
tri 5403 1644 5437 1678 se
rect 5437 1644 7826 1678
tri 5398 1639 5403 1644 se
rect 5403 1639 7826 1644
tri 2368 1636 2371 1639 sw
tri 5395 1636 5398 1639 se
rect 5398 1636 7826 1639
rect 7878 1636 7890 1688
rect 7942 1636 7948 1688
rect 8225 1678 8271 1690
rect 8225 1644 8231 1678
rect 8265 1644 8271 1678
rect 2316 1635 2371 1636
rect 171 1574 177 1626
rect 229 1574 241 1626
rect 293 1620 1065 1626
rect 293 1586 731 1620
rect 765 1586 803 1620
rect 837 1586 875 1620
rect 909 1586 947 1620
rect 981 1586 1019 1620
rect 1053 1586 1065 1620
rect 1602 1616 1652 1618
rect 293 1574 1065 1586
rect 1600 1610 1652 1616
rect 2368 1614 2371 1635
tri 2371 1614 2393 1636 sw
tri 5373 1614 5395 1636 se
rect 5395 1614 5447 1636
tri 5447 1614 5469 1636 nw
rect 2368 1594 5427 1614
tri 5427 1594 5447 1614 nw
rect 8225 1594 8271 1644
rect 10662 1609 10714 1615
rect 2368 1583 5410 1594
rect 2316 1577 5410 1583
tri 5410 1577 5427 1594 nw
rect 2316 1571 5404 1577
tri 5404 1571 5410 1577 nw
rect 1600 1546 1652 1558
rect 8225 1560 8231 1594
rect 8265 1560 8271 1594
tri 4342 1540 4345 1543 se
rect 4345 1540 4525 1543
rect 1600 1488 1652 1494
rect 2236 1488 2242 1540
rect 2294 1488 2306 1540
rect 2358 1510 3566 1540
tri 3566 1510 3596 1540 sw
tri 4312 1510 4342 1540 se
rect 4342 1537 4525 1540
rect 4342 1510 4409 1537
rect 2358 1501 3596 1510
tri 3596 1501 3605 1510 sw
tri 4303 1501 4312 1510 se
rect 4312 1501 4409 1510
rect 2358 1488 4409 1501
tri 3555 1479 3564 1488 ne
rect 3564 1485 4409 1488
rect 4461 1485 4473 1537
rect 3564 1479 4525 1485
rect 8225 1510 8271 1560
tri 3564 1476 3567 1479 ne
rect 3567 1476 4352 1479
tri 4352 1476 4355 1479 nw
rect 8225 1476 8231 1510
rect 8265 1476 8271 1510
tri 3567 1460 3583 1476 ne
rect 3583 1460 4325 1476
rect 1767 1408 1779 1460
rect 1831 1408 1843 1460
rect 1895 1408 1907 1460
rect 1959 1408 3198 1460
tri 3583 1449 3594 1460 ne
rect 3594 1449 4325 1460
tri 4325 1449 4352 1476 nw
rect 8225 1426 8271 1476
rect 8592 1592 8644 1598
tri 8644 1560 8682 1598 sw
rect 8644 1545 9271 1560
tri 9271 1545 9286 1560 sw
tri 10714 1569 10745 1600 sw
rect 10714 1563 12932 1569
rect 10714 1557 12880 1563
rect 10662 1545 12880 1557
rect 8644 1540 9286 1545
rect 8592 1528 9286 1540
rect 8644 1527 9286 1528
tri 9286 1527 9304 1545 sw
rect 9439 1539 9491 1545
rect 8644 1508 9304 1527
tri 9304 1508 9323 1527 sw
rect 8592 1470 8644 1476
tri 8644 1470 8682 1508 nw
tri 9249 1470 9287 1508 ne
rect 9287 1475 9323 1508
tri 9323 1475 9356 1508 sw
rect 9287 1470 9356 1475
tri 9287 1453 9304 1470 ne
tri 8212 1392 8225 1405 se
rect 8225 1392 8231 1426
rect 8265 1392 8271 1426
tri 8196 1376 8212 1392 se
rect 8212 1376 8271 1392
rect 4409 1372 8271 1376
rect 4409 1370 8254 1372
rect 4461 1355 8254 1370
tri 8254 1355 8271 1372 nw
rect 9304 1355 9356 1470
rect 10714 1517 12880 1545
rect 10662 1487 10714 1493
tri 10714 1487 10744 1517 nw
rect 12880 1499 12932 1511
rect 9439 1473 9491 1487
rect 12880 1441 12932 1447
rect 9439 1415 9491 1421
tri 9356 1355 9359 1358 sw
rect 4461 1349 8248 1355
tri 8248 1349 8254 1355 nw
rect 9304 1349 9359 1355
tri 9359 1349 9365 1355 sw
tri 13266 1349 13272 1355 ne
rect 4461 1344 8243 1349
tri 8243 1344 8248 1349 nw
rect 9304 1344 9365 1349
tri 9365 1344 9370 1349 sw
rect 4461 1343 4516 1344
rect 9304 1343 9370 1344
tri 9370 1343 9371 1344 sw
rect 4461 1318 4470 1343
rect 4409 1313 4470 1318
tri 4470 1313 4500 1343 nw
rect 9304 1336 9371 1343
tri 9371 1336 9378 1343 sw
tri 9304 1313 9327 1336 ne
rect 9327 1314 9378 1336
tri 9378 1314 9400 1336 sw
rect 9327 1313 10199 1314
rect 4409 1306 4461 1313
tri 4461 1304 4470 1313 nw
tri 9327 1304 9336 1313 ne
rect 9336 1304 10199 1313
tri 9336 1262 9378 1304 ne
rect 9378 1262 10199 1304
rect 10249 1261 10368 1311
rect 11736 1261 11742 1313
rect 11794 1261 11806 1313
rect 11858 1261 13278 1313
rect 13330 1261 13342 1313
rect 13394 1261 13400 1313
rect 4409 1248 4461 1254
rect 5660 1175 5776 1181
rect 3631 1148 3947 1154
rect 346 1113 1652 1119
rect 346 1061 1600 1113
rect 346 1049 1652 1061
rect 346 1029 1600 1049
rect 398 977 438 1029
rect 346 965 438 977
rect 398 913 438 965
rect 554 977 597 1029
rect 649 997 1600 1029
rect 3683 1096 3895 1148
rect 3631 1084 3947 1096
rect 3683 1081 3895 1084
tri 3683 1056 3708 1081 nw
tri 3870 1056 3895 1081 ne
rect 3631 1026 3683 1032
rect 3895 1026 3947 1032
rect 649 985 1652 997
rect 649 977 1600 985
rect 554 965 1600 977
rect 554 913 597 965
rect 649 933 1600 965
rect 3815 1000 3867 1006
rect 649 913 1652 933
tri 3790 930 3815 955 se
rect 5660 989 5776 995
rect 6756 1175 6872 1181
rect 6756 989 6872 995
rect 3815 936 3867 948
rect 346 904 1652 913
rect 2396 878 2402 930
rect 2454 878 2466 930
rect 2518 884 3815 930
rect 8500 916 8607 1192
rect 10945 916 11156 1192
rect 2518 878 3867 884
tri 4968 814 4974 820 se
rect 4974 768 4980 820
rect 5032 768 5044 820
rect 5096 768 5102 820
tri 5102 814 5108 820 sw
tri 8331 752 8344 765 se
rect 8344 752 8350 810
tri 1438 746 1444 752 se
tri 8325 746 8331 752 se
rect 8331 746 8350 752
tri 1386 694 1438 746 se
rect 1438 694 1444 746
tri 4016 740 4022 746 se
rect 4022 694 4028 746
rect 4080 694 4092 746
rect 4144 694 4156 746
rect 4208 694 4220 746
rect 4272 694 4278 746
tri 4278 740 4284 746 sw
tri 8319 740 8325 746 se
rect 8325 740 8350 746
rect 8344 694 8350 740
rect 8466 746 8472 810
rect 9687 777 9846 806
tri 8472 746 8491 765 sw
rect 8466 740 8491 746
tri 8491 740 8497 746 sw
tri 9067 740 9073 746 se
rect 9073 740 9081 746
rect 8466 694 8472 740
rect 8500 694 8606 740
rect 9075 694 9081 740
rect 9133 694 9145 746
rect 9197 694 9209 746
rect 9261 694 9273 746
rect 9325 740 9333 746
tri 9333 740 9339 746 sw
rect 9325 694 9331 740
rect 9599 694 9605 740
tri 1358 666 1386 694 se
rect 1386 688 9605 694
rect 9657 688 9669 740
rect 9721 694 9727 740
rect 10008 725 10060 731
rect 9721 688 10008 694
rect 1386 673 10008 688
rect 10060 673 11084 694
rect 1386 666 11084 673
rect -11 653 1125 666
rect -11 601 346 653
rect 398 601 437 653
rect -11 589 437 601
rect -11 537 346 589
rect 398 537 437 589
rect -11 525 437 537
rect -11 473 346 525
rect 398 473 437 525
rect 553 601 597 653
rect 649 601 1125 653
rect 553 589 1125 601
rect 553 537 597 589
rect 649 537 1125 589
rect 553 525 1125 537
rect 553 473 597 525
rect 649 473 1125 525
rect 2552 665 2668 666
rect 2552 479 2668 485
rect 3735 654 3787 660
rect 3735 590 3787 602
rect 3735 526 3787 538
rect -11 464 1125 473
rect 3735 468 3787 474
rect 4553 658 4605 664
rect 4553 594 4605 606
rect 4553 530 4605 542
rect 4553 472 4605 478
rect 8310 464 8327 666
rect 8500 464 8636 666
rect 9605 665 9721 666
rect 9605 479 9721 485
rect 10008 661 10060 666
rect 10008 597 10060 609
rect 10008 533 10060 545
rect 10008 475 10060 481
rect 91 384 97 436
rect 149 384 161 436
rect 213 384 2402 436
rect 2454 384 2466 436
rect 2518 384 2524 436
rect 8264 384 8270 436
rect 8322 384 8334 436
rect 8386 384 10379 436
rect 1444 261 1450 313
rect 1502 261 1514 313
rect 1566 307 1652 313
rect 1566 261 1600 307
rect 1444 255 1600 261
tri 1652 268 1697 313 sw
rect 1652 255 1697 268
rect 1444 243 1697 255
rect 1444 191 1600 243
rect 1652 237 1697 243
tri 1697 237 1728 268 sw
rect 1652 225 1728 237
tri 1728 225 1740 237 sw
rect 1652 191 1740 225
rect 1444 185 1740 191
rect 3130 185 3987 237
rect 4039 185 4051 237
rect 4103 185 4115 237
rect 4167 185 4179 237
rect 4231 185 4243 237
rect 4295 185 4811 237
rect 4863 185 4875 237
rect 4927 185 5354 237
rect 5406 185 5418 237
rect 5470 185 5482 237
rect 5534 185 5658 237
rect 5710 185 5722 237
rect 5774 185 5780 237
rect 5808 216 5814 268
rect 5866 216 5878 268
rect 5930 216 8561 268
rect 8613 216 8625 268
rect 8677 216 8683 268
rect 8728 185 9081 237
rect 9133 185 9145 237
rect 9197 185 9209 237
rect 9261 185 9273 237
rect 9325 185 9605 237
rect 9657 185 9669 237
rect 9721 185 9938 237
rect 9990 185 10002 237
rect 10054 185 10586 237
rect 13606 162 13658 168
tri 13546 92 13606 152 se
rect 13606 98 13658 110
rect 11304 40 11310 92
rect 11362 40 11374 92
rect 11426 46 13606 92
rect 11426 40 13658 46
rect 13348 -1988 13658 -1982
rect 13400 -2040 13606 -1988
rect 13348 -2052 13658 -2040
rect 13400 -2104 13606 -2052
rect 13348 -2110 13658 -2104
tri 12924 -5144 12963 -5105 se
rect 12963 -5144 13709 -5105
rect 6816 -5196 6822 -5144
rect 6874 -5196 6886 -5144
rect 6938 -5157 13709 -5144
rect 13761 -5157 13776 -5105
rect 13828 -5157 13834 -5105
rect 6938 -5196 12946 -5157
tri 12946 -5196 12985 -5157 nw
<< via1 >>
rect 132 3954 312 4070
rect 6250 4018 6302 4070
rect 6328 4018 6380 4070
rect 6405 4018 6457 4070
rect 6482 4018 6534 4070
rect 6559 4018 6611 4070
rect 6250 3944 6302 3996
rect 6328 3944 6380 3996
rect 6405 3944 6457 3996
rect 6482 3944 6534 3996
rect 6559 3944 6611 3996
rect 10457 4017 10509 4069
rect 10541 4017 10593 4069
rect 10625 4017 10677 4069
rect 10709 4017 10761 4069
rect 10457 3953 10509 4005
rect 10541 3953 10593 4005
rect 10625 3953 10677 4005
rect 10709 3953 10761 4005
rect 10957 4017 11009 4069
rect 11041 4017 11093 4069
rect 11125 4017 11177 4069
rect 11209 4017 11261 4069
rect 10957 3953 11009 4005
rect 11041 3953 11093 4005
rect 11125 3953 11177 4005
rect 11209 3953 11261 4005
rect 6250 3870 6302 3922
rect 6328 3870 6380 3922
rect 6405 3870 6457 3922
rect 6482 3870 6534 3922
rect 6559 3870 6611 3922
rect 6250 3796 6302 3848
rect 6328 3796 6380 3848
rect 6405 3796 6457 3848
rect 6482 3796 6534 3848
rect 6559 3796 6611 3848
rect 6250 3722 6302 3774
rect 6328 3722 6380 3774
rect 6405 3722 6457 3774
rect 6482 3722 6534 3774
rect 6559 3722 6611 3774
rect 1364 3556 1416 3608
rect 1364 3492 1416 3544
rect 5654 3502 5706 3554
rect 5718 3502 5770 3554
rect 10886 3502 10938 3554
rect 10950 3502 11002 3554
rect 171 3377 223 3429
rect 171 3313 223 3365
rect 2003 3377 2055 3429
rect 2003 3313 2055 3365
rect 436 3087 552 3267
rect 597 3233 615 3267
rect 615 3233 649 3267
rect 597 3215 649 3233
rect 597 3195 649 3203
rect 597 3161 615 3195
rect 615 3161 649 3195
rect 597 3151 649 3161
rect 597 3123 649 3139
rect 597 3089 615 3123
rect 615 3089 649 3123
rect 597 3087 649 3089
rect 4416 3088 4532 3268
rect 13766 3221 13818 3273
rect 13830 3221 13882 3273
rect 13894 3221 13946 3273
rect 13958 3221 14010 3273
rect 13766 3149 13818 3201
rect 13830 3149 13882 3201
rect 13894 3149 13946 3201
rect 13958 3149 14010 3201
rect 13766 3076 13818 3128
rect 13830 3076 13882 3128
rect 13894 3076 13946 3128
rect 13958 3076 14010 3128
rect 3987 2997 4039 3049
rect 4051 2997 4103 3049
rect 4115 2997 4167 3049
rect 4179 2997 4231 3049
rect 4243 2997 4295 3049
rect 11154 2997 11206 3049
rect 11218 2997 11270 3049
rect 12470 2997 12522 3049
rect 12534 2997 12586 3049
rect 12598 2997 12650 3049
rect 12662 2997 12714 3049
rect 12726 2997 12778 3049
rect 13766 3003 13818 3055
rect 13830 3003 13882 3055
rect 13894 3003 13946 3055
rect 13958 3003 14010 3055
rect 91 2877 143 2929
rect 3561 2917 3613 2969
rect 3625 2917 3677 2969
rect 91 2813 143 2865
rect 4327 2911 4379 2963
rect 4327 2847 4379 2899
rect 6602 2881 6654 2933
rect 6666 2881 6718 2933
rect 8264 2877 8316 2929
rect 9373 2917 9425 2969
rect 9437 2917 9489 2969
rect 11620 2917 11672 2969
rect 11684 2917 11736 2969
rect 13552 2917 13604 2969
rect 13616 2917 13668 2969
rect 8264 2813 8316 2865
rect 12470 2727 12522 2779
rect 12534 2727 12586 2779
rect 12598 2727 12650 2779
rect 12662 2727 12714 2779
rect 12726 2727 12778 2779
rect 1680 2565 1732 2617
rect 1680 2501 1732 2553
rect 2316 2565 2368 2617
rect 2868 2567 2920 2619
rect 2316 2501 2368 2553
rect 2868 2503 2920 2555
rect 5884 2565 5936 2617
rect 5884 2501 5936 2553
rect 6676 2565 6728 2617
rect 6676 2501 6728 2553
rect 10088 2565 10140 2617
rect 10088 2501 10140 2553
rect 10662 2565 10714 2617
rect 10662 2501 10714 2553
rect 11304 2565 11356 2617
rect 11304 2501 11356 2553
rect 11418 2489 11470 2541
rect 9369 2419 9421 2471
rect 9433 2419 9485 2471
rect 11418 2425 11470 2477
rect 2798 2328 2850 2380
rect 2862 2328 2914 2380
rect 11393 2328 11445 2380
rect 11457 2328 11509 2380
rect 346 2276 398 2281
rect 346 2242 376 2276
rect 376 2242 398 2276
rect 346 2229 398 2242
rect 346 2204 398 2217
rect 346 2170 376 2204
rect 376 2170 398 2204
rect 346 2165 398 2170
rect 597 2229 649 2281
rect 597 2165 649 2217
rect 1450 2161 1566 2277
rect 2552 2164 2668 2280
rect 4811 2166 4927 2282
rect 5354 2166 5534 2282
rect 8350 2165 8466 2281
rect 8754 2276 8806 2281
rect 8754 2242 8770 2276
rect 8770 2242 8806 2276
rect 8754 2229 8806 2242
rect 8754 2204 8806 2217
rect 8754 2170 8770 2204
rect 8770 2170 8806 2204
rect 8754 2165 8806 2170
rect 9599 2165 9715 2281
rect 13434 2172 13550 2288
rect 13796 2165 13976 2281
rect 5660 1934 5776 2114
rect 6756 1934 6872 2114
rect 9110 1934 9226 2114
rect 11040 1934 11156 2114
rect 926 1842 978 1894
rect 1680 1842 1732 1894
rect 926 1778 978 1830
rect 1680 1778 1732 1830
rect 11211 1842 11263 1894
rect 11411 1842 11463 1894
rect 11211 1778 11263 1830
rect 11411 1778 11463 1830
rect 7982 1756 8034 1777
rect 8046 1756 8098 1777
rect 7982 1725 8007 1756
rect 8007 1725 8034 1756
rect 8046 1725 8079 1756
rect 8079 1725 8098 1756
rect 2316 1647 2368 1699
rect 7826 1636 7878 1688
rect 7890 1636 7942 1688
rect 177 1574 229 1626
rect 241 1574 293 1626
rect 1600 1558 1652 1610
rect 2316 1583 2368 1635
rect 1600 1494 1652 1546
rect 2242 1488 2294 1540
rect 2306 1488 2358 1540
rect 4409 1485 4461 1537
rect 4473 1485 4525 1537
rect 1779 1408 1831 1460
rect 1843 1408 1895 1460
rect 1907 1408 1959 1460
rect 8592 1540 8644 1592
rect 10662 1557 10714 1609
rect 8592 1476 8644 1528
rect 4409 1318 4461 1370
rect 9439 1487 9491 1539
rect 10662 1493 10714 1545
rect 12880 1511 12932 1563
rect 9439 1421 9491 1473
rect 12880 1447 12932 1499
rect 4409 1254 4461 1306
rect 11742 1261 11794 1313
rect 11806 1261 11858 1313
rect 13278 1261 13330 1313
rect 13342 1261 13394 1313
rect 1600 1061 1652 1113
rect 346 977 398 1029
rect 346 913 398 965
rect 438 913 554 1029
rect 597 977 649 1029
rect 1600 997 1652 1049
rect 3631 1096 3683 1148
rect 3895 1096 3947 1148
rect 3631 1032 3683 1084
rect 3895 1032 3947 1084
rect 597 913 649 965
rect 1600 933 1652 985
rect 3815 948 3867 1000
rect 5660 995 5776 1175
rect 6756 995 6872 1175
rect 2402 878 2454 930
rect 2466 878 2518 930
rect 3815 884 3867 936
rect 4980 768 5032 820
rect 5044 768 5096 820
rect 4028 694 4080 746
rect 4092 694 4144 746
rect 4156 694 4208 746
rect 4220 694 4272 746
rect 8350 694 8466 810
rect 9081 694 9133 746
rect 9145 694 9197 746
rect 9209 694 9261 746
rect 9273 694 9325 746
rect 9605 688 9657 740
rect 9669 688 9721 740
rect 10008 673 10060 725
rect 346 601 398 653
rect 346 537 398 589
rect 346 473 398 525
rect 437 473 553 653
rect 597 601 649 653
rect 597 537 649 589
rect 597 473 649 525
rect 2552 485 2668 665
rect 3735 602 3787 654
rect 3735 538 3787 590
rect 3735 474 3787 526
rect 4553 606 4605 658
rect 4553 542 4605 594
rect 4553 478 4605 530
rect 9605 485 9721 665
rect 10008 609 10060 661
rect 10008 545 10060 597
rect 10008 481 10060 533
rect 97 384 149 436
rect 161 384 213 436
rect 2402 384 2454 436
rect 2466 384 2518 436
rect 8270 384 8322 436
rect 8334 384 8386 436
rect 1450 261 1502 313
rect 1514 261 1566 313
rect 1600 255 1652 307
rect 1600 191 1652 243
rect 3987 185 4039 237
rect 4051 185 4103 237
rect 4115 185 4167 237
rect 4179 185 4231 237
rect 4243 185 4295 237
rect 4811 185 4863 237
rect 4875 185 4927 237
rect 5354 185 5406 237
rect 5418 185 5470 237
rect 5482 185 5534 237
rect 5658 185 5710 237
rect 5722 185 5774 237
rect 5814 216 5866 268
rect 5878 216 5930 268
rect 8561 216 8613 268
rect 8625 216 8677 268
rect 9081 185 9133 237
rect 9145 185 9197 237
rect 9209 185 9261 237
rect 9273 185 9325 237
rect 9605 185 9657 237
rect 9669 185 9721 237
rect 9938 185 9990 237
rect 10002 185 10054 237
rect 13606 110 13658 162
rect 11310 40 11362 92
rect 11374 40 11426 92
rect 13606 46 13658 98
rect 13348 -2040 13400 -1988
rect 13606 -2040 13658 -1988
rect 13348 -2104 13400 -2052
rect 13606 -2104 13658 -2052
rect 6822 -5196 6874 -5144
rect 6886 -5196 6938 -5144
rect 13709 -5157 13761 -5105
rect 13776 -5157 13828 -5105
<< metal2 >>
rect 126 4070 318 4141
rect 126 3954 132 4070
rect 312 3954 318 4070
rect 126 3952 318 3954
rect 346 3540 582 4141
rect 346 3446 552 3540
tri 552 3510 582 3540 nw
tri 346 3435 357 3446 ne
rect 357 3435 552 3446
rect 171 3429 223 3435
tri 357 3429 363 3435 ne
rect 363 3429 552 3435
tri 363 3377 415 3429 ne
rect 415 3377 552 3429
rect 171 3365 223 3377
tri 415 3365 427 3377 ne
rect 427 3365 552 3377
tri 427 3356 436 3365 ne
rect 91 2929 143 2935
rect 91 2865 143 2877
rect 91 436 143 2813
rect 171 1647 223 3313
rect 436 3267 552 3365
rect 436 3081 552 3087
rect 597 3267 649 3273
rect 597 3203 649 3215
rect 597 3139 649 3151
rect 346 2281 398 2497
rect 346 2217 398 2229
tri 223 1647 227 1651 sw
rect 171 1636 227 1647
tri 227 1636 238 1647 sw
rect 171 1635 238 1636
tri 238 1635 239 1636 sw
rect 171 1626 239 1635
tri 239 1626 248 1635 sw
rect 171 1574 177 1626
rect 229 1574 241 1626
rect 293 1574 299 1626
rect 346 1476 398 2165
rect 597 2281 649 3087
rect 597 2217 649 2229
tri 398 1476 407 1485 sw
tri 588 1476 597 1485 se
rect 597 1476 649 2165
rect 926 1894 978 4141
rect 926 1830 978 1842
rect 926 1772 978 1778
rect 346 1473 407 1476
tri 407 1473 410 1476 sw
tri 585 1473 588 1476 se
rect 588 1473 649 1476
rect 346 1460 410 1473
tri 410 1460 423 1473 sw
tri 572 1460 585 1473 se
rect 585 1460 649 1473
tri 333 1447 346 1460 se
rect 346 1447 649 1460
rect 333 1175 649 1447
rect 1006 1228 1336 4141
rect 1364 3608 1416 4141
rect 1364 3544 1416 3556
rect 1364 3486 1416 3492
rect 1444 2933 1496 4141
rect 1524 3318 1975 4456
tri 11304 4195 11317 4208 se
rect 11317 4195 11369 4273
tri 8567 4181 8570 4184 ne
rect 8570 4181 8652 4184
tri 8652 4181 8655 4184 nw
rect 9932 4181 10073 4191
rect 11304 4186 11369 4195
rect 11304 4181 11364 4186
tri 11364 4181 11369 4186 nw
tri 8570 4159 8592 4181 ne
tri 1524 3313 1529 3318 ne
rect 1529 3313 1975 3318
tri 1529 3307 1535 3313 ne
rect 1535 3307 1975 3313
rect 2003 3429 2055 4156
rect 2003 3365 2055 3377
rect 2003 3307 2055 3313
tri 1535 3273 1569 3307 ne
rect 1569 3273 1975 3307
tri 1569 3268 1574 3273 ne
rect 1574 3268 1975 3273
tri 1574 3088 1754 3268 ne
rect 1754 3088 1975 3268
tri 1754 3082 1760 3088 ne
tri 1496 2933 1521 2958 sw
rect 1680 2617 1732 2623
rect 1680 2553 1732 2565
tri 1584 2350 1600 2366 se
tri 1562 2328 1584 2350 se
rect 1584 2328 1600 2350
tri 1522 2288 1562 2328 se
rect 1562 2288 1600 2328
tri 1516 2282 1522 2288 se
rect 1522 2282 1600 2288
tri 1514 2280 1516 2282 se
rect 1516 2280 1600 2282
tri 1511 2277 1514 2280 se
rect 1514 2277 1600 2280
rect 1444 2161 1450 2277
rect 1566 2161 1652 2277
rect 1444 1610 1652 2161
rect 1444 1558 1600 1610
rect 1444 1546 1652 1558
rect 1444 1494 1600 1546
tri 649 1175 653 1179 sw
rect 333 1148 653 1175
tri 653 1148 680 1175 sw
rect 333 1113 680 1148
tri 680 1113 715 1148 sw
rect 1444 1113 1652 1494
rect 333 1061 715 1113
tri 715 1061 767 1113 sw
rect 1444 1061 1600 1113
rect 333 1049 767 1061
tri 767 1049 779 1061 sw
rect 1444 1049 1652 1061
rect 333 1035 779 1049
tri 779 1035 793 1049 sw
rect 333 1029 793 1035
rect 333 977 346 1029
rect 398 977 438 1029
rect 333 965 438 977
rect 333 913 346 965
rect 398 913 438 965
rect 554 977 597 1029
rect 649 977 793 1029
rect 554 965 793 977
rect 554 913 597 965
rect 649 913 793 965
rect 333 653 793 913
rect 333 601 346 653
rect 398 601 437 653
rect 333 589 437 601
rect 333 537 346 589
rect 398 537 437 589
rect 333 525 437 537
rect 333 473 346 525
rect 398 473 437 525
rect 553 601 597 653
rect 649 601 793 653
rect 553 589 793 601
rect 553 537 597 589
rect 649 537 793 589
rect 553 525 793 537
rect 553 473 597 525
rect 649 473 793 525
rect 333 467 793 473
rect 1444 997 1600 1049
rect 1444 985 1652 997
rect 1444 933 1600 985
tri 143 436 168 461 sw
rect 91 384 97 436
rect 149 384 161 436
rect 213 384 219 436
rect 1444 313 1652 933
rect 1444 261 1450 313
rect 1502 261 1514 313
rect 1566 307 1652 313
rect 1566 261 1600 307
rect 1444 255 1600 261
rect 1444 243 1652 255
rect 1444 191 1600 243
rect 1444 185 1652 191
rect 1680 1894 1732 2501
rect 1680 1830 1732 1842
rect 1680 0 1732 1778
rect 1760 1460 1975 3088
rect 1760 1408 1779 1460
rect 1831 1408 1843 1460
rect 1895 1408 1907 1460
rect 1959 1408 1975 1460
rect 2088 0 2208 4141
rect 2236 1540 2288 4141
rect 2316 2617 2368 4141
rect 2552 3138 2604 4141
tri 2604 3138 2629 3163 sw
rect 2552 3120 2712 3138
tri 2552 3090 2582 3120 ne
rect 2582 3090 2712 3120
tri 2712 3090 2760 3138 sw
tri 2582 3088 2584 3090 ne
rect 2584 3088 2760 3090
tri 2584 3086 2586 3088 ne
rect 2586 3086 2760 3088
tri 2683 3076 2693 3086 ne
rect 2693 3076 2760 3086
tri 2693 3061 2708 3076 ne
tri 2683 2933 2708 2958 se
rect 2708 2928 2760 3076
rect 2316 2553 2368 2565
rect 2316 1699 2368 2501
rect 2868 2619 2920 2625
rect 2868 2555 2920 2567
tri 2831 2419 2868 2456 se
rect 2868 2419 2920 2503
tri 2792 2380 2831 2419 se
rect 2831 2380 2920 2419
rect 2316 1635 2368 1647
rect 2316 1577 2368 1583
rect 2552 2328 2604 2350
tri 2604 2328 2626 2350 sw
rect 2792 2328 2798 2380
rect 2850 2328 2862 2380
rect 2914 2328 2920 2380
rect 2552 2288 2626 2328
tri 2626 2288 2666 2328 sw
rect 2552 2287 2666 2288
tri 2666 2287 2667 2288 sw
rect 2552 2286 2667 2287
tri 2667 2286 2668 2287 sw
rect 2552 2280 2668 2286
tri 2288 1540 2313 1565 sw
rect 2236 1488 2242 1540
rect 2294 1488 2306 1540
rect 2358 1488 2364 1540
rect 2396 878 2402 930
rect 2454 878 2466 930
rect 2518 878 2524 930
rect 2396 436 2524 878
rect 2552 704 2668 2164
rect 2948 1171 3192 4141
rect 3745 3375 3797 4122
tri 3745 3336 3784 3375 ne
rect 3784 3336 3797 3375
tri 3797 3336 3858 3397 sw
tri 3784 3323 3797 3336 ne
rect 3797 3323 3858 3336
tri 3797 3314 3806 3323 ne
rect 3806 3273 3858 3323
rect 3981 3049 4301 4122
rect 5050 4103 5102 4141
rect 5648 3554 5700 4141
tri 5700 3554 5725 3579 sw
rect 5648 3502 5654 3554
rect 5706 3502 5718 3554
rect 5770 3502 5776 3554
rect 4416 3268 4602 3274
rect 4532 3088 4602 3268
rect 4416 3078 4602 3088
tri 4449 3076 4451 3078 ne
rect 4451 3076 4550 3078
tri 4451 3055 4472 3076 ne
rect 4472 3055 4550 3076
tri 4472 3049 4478 3055 ne
rect 4478 3049 4550 3055
rect 3981 2997 3987 3049
rect 4039 2997 4051 3049
rect 4103 2997 4115 3049
rect 4167 2997 4179 3049
rect 4231 2997 4243 3049
rect 4295 2997 4301 3049
tri 4478 2997 4530 3049 ne
rect 4530 2997 4550 3049
rect 3981 2983 4301 2997
rect 3555 2917 3561 2969
rect 3613 2917 3625 2969
rect 3677 2917 3683 2969
tri 3606 2911 3612 2917 ne
rect 3612 2911 3683 2917
tri 3612 2899 3624 2911 ne
rect 3624 2899 3683 2911
tri 3624 2892 3631 2899 ne
rect 3631 1148 3683 2899
rect 3981 2772 4299 2983
tri 4299 2981 4301 2983 nw
tri 4530 2981 4546 2997 ne
rect 4546 2981 4550 2997
tri 4546 2977 4550 2981 ne
rect 4327 2963 4379 2969
rect 4327 2899 4379 2911
rect 5648 2935 5700 3502
tri 5700 3477 5725 3502 nw
tri 5700 2935 5723 2958 sw
rect 5648 2933 5723 2935
tri 5723 2933 5725 2935 sw
rect 5648 2876 5700 2933
rect 4327 2807 4379 2847
tri 4379 2807 4380 2808 sw
rect 4327 2806 4380 2807
tri 4380 2806 4381 2807 sw
rect 4327 2786 4381 2806
tri 4327 2784 4329 2786 ne
tri 4299 2772 4301 2774 sw
tri 3766 1725 3806 1765 se
rect 3806 1743 3858 2508
rect 3806 1725 3840 1743
tri 3840 1725 3858 1743 nw
rect 3631 1084 3683 1096
rect 3631 1026 3683 1032
tri 3735 1694 3766 1725 se
rect 3766 1694 3809 1725
tri 3809 1694 3840 1725 nw
rect 3735 1688 3803 1694
tri 3803 1688 3809 1694 nw
rect 2552 665 2668 671
rect 2552 479 2668 485
rect 3735 654 3787 1688
tri 3787 1672 3803 1688 nw
rect 3895 1148 3947 1154
rect 3895 1084 3947 1096
rect 3735 590 3787 602
rect 3735 526 3787 538
rect 3735 468 3787 474
rect 3815 1000 3867 1006
rect 3815 936 3867 948
rect 2396 384 2402 436
rect 2454 384 2466 436
rect 2518 384 2524 436
rect 3815 0 3867 884
rect 3895 0 3947 1032
rect 3981 746 4301 2772
rect 3981 694 4028 746
rect 4080 694 4092 746
rect 4144 694 4156 746
rect 4208 694 4220 746
rect 4272 694 4301 746
rect 3981 237 4301 694
rect 3981 185 3987 237
rect 4039 185 4051 237
rect 4103 185 4115 237
rect 4167 185 4179 237
rect 4231 185 4243 237
rect 4295 185 4301 237
rect 3981 0 4301 185
rect 4329 0 4381 2786
rect 5884 2617 5936 4141
rect 6244 4018 6250 4070
rect 6302 4068 6328 4070
rect 6380 4068 6405 4070
rect 6457 4068 6482 4070
rect 6534 4068 6559 4070
rect 6309 4018 6328 4068
rect 6534 4018 6552 4068
rect 6611 4018 6617 4070
rect 6244 4012 6253 4018
rect 6309 4012 6353 4018
rect 6409 4012 6453 4018
rect 6509 4012 6552 4018
rect 6608 4012 6617 4018
rect 6244 3996 6617 4012
rect 6244 3944 6250 3996
rect 6302 3972 6328 3996
rect 6380 3972 6405 3996
rect 6457 3972 6482 3996
rect 6534 3972 6559 3996
rect 6309 3944 6328 3972
rect 6534 3944 6552 3972
rect 6611 3944 6617 3996
rect 6244 3922 6253 3944
rect 6309 3922 6353 3944
rect 6409 3922 6453 3944
rect 6509 3922 6552 3944
rect 6608 3922 6617 3944
rect 6244 3870 6250 3922
rect 6309 3916 6328 3922
rect 6534 3916 6552 3922
rect 6302 3876 6328 3916
rect 6380 3876 6405 3916
rect 6457 3876 6482 3916
rect 6534 3876 6559 3916
rect 6309 3870 6328 3876
rect 6534 3870 6552 3876
rect 6611 3870 6617 3922
rect 6244 3848 6253 3870
rect 6309 3848 6353 3870
rect 6409 3848 6453 3870
rect 6509 3848 6552 3870
rect 6608 3848 6617 3870
rect 6244 3796 6250 3848
rect 6309 3820 6328 3848
rect 6534 3820 6552 3848
rect 6302 3796 6328 3820
rect 6380 3796 6405 3820
rect 6457 3796 6482 3820
rect 6534 3796 6559 3820
rect 6611 3796 6617 3848
rect 6244 3780 6617 3796
rect 6244 3774 6253 3780
rect 6309 3774 6353 3780
rect 6409 3774 6453 3780
rect 6509 3774 6552 3780
rect 6608 3774 6617 3780
rect 6244 3722 6250 3774
rect 6309 3724 6328 3774
rect 6534 3724 6552 3774
rect 6302 3722 6328 3724
rect 6380 3722 6405 3724
rect 6457 3722 6482 3724
rect 6534 3722 6559 3724
rect 6611 3722 6617 3774
rect 6980 2958 7307 4122
rect 8010 3081 8382 4122
rect 8427 3307 8491 4122
tri 8491 3307 8516 3332 sw
rect 8427 3306 8516 3307
tri 8427 3274 8459 3306 ne
rect 8459 3279 8516 3306
tri 8516 3279 8544 3307 sw
rect 8459 3274 8544 3279
tri 8544 3274 8549 3279 sw
tri 8459 3273 8460 3274 ne
rect 8460 3273 8549 3274
tri 8549 3273 8550 3274 sw
tri 8460 3259 8474 3273 ne
rect 8474 3259 8550 3273
tri 8550 3259 8564 3273 sw
tri 8474 3242 8491 3259 ne
rect 8491 3242 8564 3259
tri 8491 3233 8500 3242 ne
tri 6980 2946 6992 2958 ne
rect 6596 2881 6602 2933
rect 6654 2881 6666 2933
rect 6718 2881 6724 2933
rect 6596 2877 6669 2881
tri 6669 2877 6673 2881 nw
rect 6596 2865 6657 2877
tri 6657 2865 6669 2877 nw
rect 5884 2553 5936 2565
rect 4550 1662 4602 2497
rect 4805 2166 4811 2282
rect 4927 2166 4933 2282
tri 4602 1662 4605 1665 sw
rect 4550 1613 4605 1662
tri 4550 1610 4553 1613 ne
rect 4409 1537 4525 1543
rect 4461 1485 4473 1537
rect 4409 1479 4525 1485
rect 4409 1370 4461 1376
rect 4409 1306 4461 1318
rect 4409 0 4461 1254
rect 4553 658 4605 1613
rect 4553 594 4605 606
rect 4553 530 4605 542
rect 4553 0 4605 478
rect 4805 237 4933 2166
rect 5348 2166 5354 2282
rect 5534 2166 5540 2282
tri 5025 820 5050 845 se
rect 5050 820 5102 1794
rect 4974 768 4980 820
rect 5032 768 5044 820
rect 5096 768 5102 820
rect 4805 185 4811 237
rect 4863 185 4875 237
rect 4927 185 4933 237
rect 5348 237 5540 2166
rect 5660 2114 5776 2120
rect 5660 1175 5776 1934
rect 5660 989 5776 995
tri 5736 878 5804 946 se
rect 5804 924 5856 2158
tri 5730 872 5736 878 se
rect 5736 872 5804 878
tri 5804 872 5856 924 nw
tri 5678 820 5730 872 se
rect 5730 820 5780 872
tri 5780 848 5804 872 nw
tri 5668 810 5678 820 se
rect 5678 810 5780 820
rect 5348 185 5354 237
rect 5406 185 5418 237
rect 5470 185 5482 237
rect 5534 185 5540 237
tri 5652 794 5668 810 se
rect 5668 794 5780 810
rect 5652 237 5780 794
tri 5859 268 5884 293 se
rect 5884 268 5936 2501
rect 5652 185 5658 237
rect 5710 185 5722 237
rect 5774 185 5780 237
rect 5808 216 5814 268
rect 5866 216 5878 268
rect 5930 216 5936 268
rect 6225 0 6545 2813
rect 6596 0 6648 2865
tri 6648 2856 6657 2865 nw
rect 6676 2617 6728 2623
rect 6676 2553 6728 2565
rect 6676 0 6728 2501
tri 6986 2489 6992 2495 se
rect 6992 2489 7307 2958
rect 8062 3078 8266 3081
tri 8266 3078 8269 3081 nw
rect 8062 3076 8264 3078
tri 8264 3076 8266 3078 nw
rect 8062 3055 8243 3076
tri 8243 3055 8264 3076 nw
rect 8062 3049 8237 3055
tri 8237 3049 8243 3055 nw
rect 8062 2997 8185 3049
tri 8185 2997 8237 3049 nw
rect 8062 2977 8165 2997
tri 8165 2977 8185 2997 nw
rect 8062 2969 8157 2977
tri 8157 2969 8165 2977 nw
rect 8062 2958 8146 2969
tri 8146 2958 8157 2969 nw
rect 8062 2935 8123 2958
tri 8123 2935 8146 2958 nw
rect 8062 2933 8121 2935
tri 8121 2933 8123 2935 nw
rect 8062 2929 8117 2933
tri 8117 2929 8121 2933 nw
rect 8264 2929 8316 2935
rect 8062 2881 8069 2929
tri 8069 2881 8117 2929 nw
rect 8062 2877 8065 2881
tri 8065 2877 8069 2881 nw
tri 8062 2874 8065 2877 nw
tri 6982 2485 6986 2489 se
rect 6986 2485 7307 2489
rect 6756 2114 6872 2120
rect 6756 1175 6872 1934
rect 6756 989 6872 995
rect 6982 1778 7307 2485
rect 8264 2865 8316 2877
tri 7307 1778 7342 1813 sw
rect 6982 1777 7342 1778
tri 7342 1777 7343 1778 sw
rect 6982 1725 7343 1777
tri 7343 1725 7395 1777 sw
rect 7976 1725 7982 1777
rect 8034 1725 8046 1777
rect 8098 1725 8104 1777
rect 6982 1688 7395 1725
tri 7395 1688 7432 1725 sw
rect 6982 1636 7432 1688
tri 7432 1636 7484 1688 sw
rect 7820 1636 7826 1688
rect 7878 1636 7890 1688
rect 7942 1636 7948 1688
rect 6982 1611 7484 1636
tri 7484 1611 7509 1636 sw
tri 7871 1611 7896 1636 ne
rect 6982 1609 7509 1611
tri 7509 1609 7511 1611 sw
rect 6982 1592 7511 1609
tri 7511 1592 7528 1609 sw
rect 6982 1540 7528 1592
tri 7528 1540 7580 1592 sw
rect 6982 1539 7580 1540
tri 7580 1539 7581 1540 sw
rect 6982 1528 7581 1539
tri 7581 1528 7592 1539 sw
rect 6982 1490 7592 1528
tri 7592 1490 7630 1528 sw
rect 6982 1481 7630 1490
rect 6982 1425 7353 1481
rect 7409 1425 7433 1481
rect 7489 1476 7630 1481
tri 7630 1476 7644 1490 sw
rect 7489 1473 7644 1476
tri 7644 1473 7647 1476 sw
rect 7489 1436 7647 1473
tri 7647 1436 7684 1473 sw
rect 7489 1425 7795 1436
rect 6982 1395 7795 1425
rect 6982 1339 7353 1395
rect 7409 1339 7433 1395
rect 7489 1339 7795 1395
rect 6982 1308 7795 1339
rect 6982 1252 7353 1308
rect 7409 1252 7433 1308
rect 7489 1252 7585 1308
rect 7641 1252 7795 1308
rect 6982 1221 7795 1252
rect 6982 1165 7353 1221
rect 7409 1165 7433 1221
rect 7489 1165 7585 1221
rect 7641 1165 7795 1221
rect 6982 1134 7795 1165
rect 6982 1078 7353 1134
rect 7409 1078 7433 1134
rect 7489 1078 7585 1134
rect 7641 1078 7795 1134
rect 6982 0 7795 1078
rect 7896 0 7948 1636
rect 7976 0 8028 1725
tri 8028 1700 8053 1725 nw
rect 8264 436 8316 2813
rect 8344 2165 8350 2281
rect 8466 2165 8472 2281
rect 8344 810 8472 2165
rect 8344 694 8350 810
rect 8466 694 8472 810
rect 8500 568 8564 3242
rect 8592 1598 8631 4181
tri 8631 4160 8652 4181 nw
rect 8754 3273 8806 4122
rect 10451 4069 10767 4070
rect 10451 4017 10457 4069
rect 10509 4017 10541 4069
rect 10593 4017 10625 4069
rect 10677 4017 10709 4069
rect 10761 4017 10767 4069
rect 10451 4005 10767 4017
rect 10451 3953 10457 4005
rect 10509 3953 10541 4005
rect 10593 3953 10625 4005
rect 10677 3953 10709 4005
rect 10761 3953 10767 4005
rect 10451 3952 10767 3953
rect 10951 4069 11267 4070
rect 10951 4017 10957 4069
rect 11009 4017 11041 4069
rect 11093 4017 11125 4069
rect 11177 4017 11209 4069
rect 11261 4017 11267 4069
rect 10951 4005 11267 4017
rect 10951 3953 10957 4005
rect 11009 3953 11041 4005
rect 11093 3953 11125 4005
rect 11177 3953 11209 4005
rect 11261 3953 11267 4005
rect 10951 3952 11267 3953
rect 10880 3502 10886 3554
rect 10938 3502 10950 3554
rect 11002 3502 11008 3554
rect 9367 2917 9373 2969
rect 9425 2917 9437 2969
rect 9489 2917 9571 2969
tri 9494 2892 9519 2917 ne
rect 8754 2281 8806 2497
rect 9363 2419 9369 2471
rect 9421 2419 9433 2471
rect 9485 2419 9491 2471
rect 8754 2217 8806 2229
rect 8592 1592 8644 1598
rect 8592 1528 8644 1540
rect 8592 1470 8644 1476
rect 8754 694 8806 2165
rect 9110 2114 9226 2120
rect 9110 989 9226 1934
rect 9439 1539 9491 2419
rect 9439 1473 9491 1487
rect 9439 1415 9491 1421
tri 8806 694 8857 745 sw
rect 9075 694 9081 746
rect 9133 694 9145 746
rect 9197 694 9209 746
rect 9261 694 9273 746
rect 9325 694 9331 746
rect 8754 688 8857 694
tri 8857 688 8863 694 sw
rect 8754 673 8863 688
tri 8863 673 8878 688 sw
rect 8754 665 8878 673
tri 8878 665 8886 673 sw
tri 8500 563 8505 568 ne
rect 8505 563 8564 568
tri 8564 563 8595 594 sw
tri 8505 504 8564 563 ne
rect 8564 504 8595 563
tri 8564 485 8583 504 ne
rect 8583 485 8595 504
tri 8595 485 8673 563 sw
tri 8583 481 8587 485 ne
rect 8587 481 8673 485
tri 8673 481 8677 485 sw
tri 8587 473 8595 481 ne
rect 8595 473 8677 481
tri 8677 473 8685 481 sw
tri 8595 461 8607 473 ne
rect 8607 461 8685 473
tri 8316 436 8341 461 sw
tri 8607 436 8632 461 ne
rect 8632 436 8685 461
tri 8685 436 8722 473 sw
rect 8754 467 9047 665
tri 8754 436 8785 467 ne
rect 8785 436 9047 467
rect 8264 384 8270 436
rect 8322 384 8334 436
rect 8386 384 8392 436
tri 8632 384 8684 436 ne
rect 8684 418 8722 436
tri 8722 418 8740 436 sw
tri 8785 418 8803 436 ne
rect 8684 384 8740 418
tri 8740 384 8774 418 sw
tri 8684 383 8685 384 ne
rect 8685 383 8774 384
tri 8774 383 8775 384 sw
tri 8685 357 8711 383 ne
rect 8555 216 8561 268
rect 8613 216 8625 268
rect 8677 216 8683 268
tri 8606 191 8631 216 ne
rect 8631 0 8683 216
rect 8711 0 8775 383
rect 8803 0 9047 436
rect 9075 237 9331 694
rect 9075 185 9081 237
rect 9133 185 9145 237
rect 9197 185 9209 237
rect 9261 185 9273 237
rect 9325 185 9331 237
rect 9519 0 9571 2917
rect 9833 2509 9885 2933
rect 10088 2617 10140 2623
rect 10088 2553 10140 2565
rect 9833 2501 9902 2509
tri 9902 2501 9910 2509 nw
rect 9833 2489 9890 2501
tri 9890 2489 9902 2501 nw
rect 9599 2281 9725 2287
rect 9715 2165 9725 2281
rect 9599 1758 9725 2165
tri 9725 1758 9727 1760 sw
rect 9599 740 9727 1758
rect 9599 688 9605 740
rect 9657 688 9669 740
rect 9721 688 9727 740
rect 9599 665 9727 688
rect 9599 485 9605 665
rect 9721 485 9727 665
rect 9599 237 9727 485
rect 9599 185 9605 237
rect 9657 185 9669 237
rect 9721 185 9727 237
rect 9833 0 9885 2489
tri 9885 2484 9890 2489 nw
rect 10008 725 10060 2169
rect 10008 661 10060 673
rect 10008 597 10060 609
rect 10008 533 10060 545
tri 10005 268 10008 271 se
rect 10008 268 10060 481
tri 9988 251 10005 268 se
rect 10005 251 10060 268
tri 9974 237 9988 251 se
rect 9988 237 10060 251
rect 9932 185 9938 237
rect 9990 185 10002 237
rect 10054 185 10060 237
rect 10088 0 10140 2501
rect 10296 0 10612 2794
rect 10662 2617 10714 2623
rect 10662 2553 10714 2565
rect 10662 1609 10714 2501
rect 10662 1545 10714 1557
rect 10662 1487 10714 1493
rect 10880 0 10932 3502
tri 10932 3477 10957 3502 nw
rect 11032 2997 11154 3049
rect 11206 2997 11218 3049
rect 11270 2997 11276 3049
tri 11171 2972 11196 2997 ne
tri 11012 2288 11035 2311 sw
tri 11173 2288 11196 2311 se
rect 11196 2288 11276 2997
rect 11304 2824 11356 4181
tri 11356 4173 11364 4181 nw
rect 11418 3953 11930 4122
rect 12464 3049 12784 4122
rect 12464 2997 12470 3049
rect 12522 2997 12534 3049
rect 12586 2997 12598 3049
rect 12650 2997 12662 3049
rect 12714 2997 12726 3049
rect 12778 2997 12784 3049
rect 11614 2917 11620 2969
rect 11672 2917 11684 2969
rect 11736 2917 11742 2969
tri 11356 2824 11378 2846 sw
tri 11304 2807 11321 2824 ne
rect 11321 2807 11378 2824
tri 11321 2779 11349 2807 ne
rect 11349 2784 11378 2807
tri 11378 2784 11418 2824 sw
rect 11349 2779 11418 2784
tri 11418 2779 11423 2784 sw
tri 11349 2750 11378 2779 ne
rect 11378 2750 11423 2779
tri 11423 2750 11452 2779 sw
tri 11378 2727 11401 2750 ne
rect 11401 2732 11452 2750
tri 11452 2732 11470 2750 sw
rect 11401 2727 11470 2732
tri 11401 2710 11418 2727 ne
rect 11012 2287 11035 2288
tri 11035 2287 11036 2288 sw
tri 11172 2287 11173 2288 se
rect 11173 2287 11276 2288
rect 11012 2286 11036 2287
tri 11036 2286 11037 2287 sw
tri 11171 2286 11172 2287 se
rect 11172 2286 11276 2287
rect 10960 2158 11032 2286
rect 11196 2175 11276 2286
rect 11304 2617 11356 2629
rect 11304 2553 11356 2565
rect 11040 2114 11156 2120
rect 11040 989 11156 1934
rect 11211 1894 11263 1900
rect 11211 1830 11263 1842
tri 11196 384 11211 399 se
rect 11211 384 11263 1778
tri 11137 325 11196 384 se
rect 11196 377 11263 384
rect 11196 325 11211 377
tri 11211 325 11263 377 nw
tri 11125 313 11137 325 se
tri 11080 268 11125 313 se
rect 11125 268 11137 313
tri 11063 251 11080 268 se
rect 11080 251 11137 268
tri 11137 251 11211 325 nw
tri 11049 237 11063 251 se
tri 10997 185 11049 237 se
rect 11049 185 11063 237
tri 10989 177 10997 185 se
rect 10997 177 11063 185
tri 11063 177 11137 251 nw
tri 10974 162 10989 177 se
rect 10989 162 11048 177
tri 11048 162 11063 177 nw
tri 10960 148 10974 162 se
rect 10974 148 11034 162
tri 11034 148 11048 162 nw
rect 10960 -17 11012 148
tri 11012 126 11034 148 nw
rect 11304 126 11356 2501
rect 11418 2541 11470 2727
rect 11418 2477 11470 2489
rect 11418 2418 11470 2425
rect 11652 2380 11704 2917
rect 12464 2779 12784 2997
rect 13766 3273 14011 4122
rect 14495 3722 14815 4122
rect 13818 3221 13830 3273
rect 13882 3221 13894 3273
rect 13946 3221 13958 3273
rect 14010 3221 14011 3273
rect 13766 3201 14011 3221
rect 13818 3149 13830 3201
rect 13882 3149 13894 3201
rect 13946 3149 13958 3201
rect 14010 3149 14011 3201
rect 13766 3128 14011 3149
rect 13818 3076 13830 3128
rect 13882 3076 13894 3128
rect 13946 3076 13958 3128
rect 14010 3076 14011 3128
rect 13766 3055 14011 3076
rect 13818 3003 13830 3055
rect 13882 3003 13894 3055
rect 13946 3003 13958 3055
rect 14010 3003 14011 3055
rect 13546 2917 13552 2969
rect 13604 2917 13616 2969
rect 13668 2917 13674 2969
tri 13546 2879 13584 2917 ne
rect 12464 2727 12470 2779
rect 12522 2727 12534 2779
rect 12586 2727 12598 2779
rect 12650 2727 12662 2779
rect 12714 2727 12726 2779
rect 12778 2727 12784 2779
tri 11704 2380 11721 2397 sw
rect 11387 2328 11393 2380
rect 11445 2328 11457 2380
rect 11509 2328 11515 2380
rect 11652 2375 11721 2380
tri 11721 2375 11726 2380 sw
tri 11652 2328 11699 2375 ne
rect 11699 2328 11726 2375
tri 11387 2304 11411 2328 ne
rect 11411 2304 11491 2328
tri 11491 2304 11515 2328 nw
tri 11699 2304 11723 2328 ne
rect 11723 2313 11726 2328
tri 11726 2313 11788 2375 sw
rect 11723 2304 11788 2313
rect 11411 2301 11488 2304
tri 11488 2301 11491 2304 nw
tri 11723 2301 11726 2304 ne
rect 11726 2301 11788 2304
rect 11411 2291 11478 2301
tri 11478 2291 11488 2301 nw
tri 11726 2291 11736 2301 ne
rect 11411 2288 11475 2291
tri 11475 2288 11478 2291 nw
rect 11411 2287 11474 2288
tri 11474 2287 11475 2288 nw
rect 11411 1894 11463 2287
tri 11463 2276 11474 2287 nw
rect 11411 1830 11463 1842
rect 11411 1772 11463 1778
rect 11492 437 11672 1928
rect 11736 1313 11788 2301
tri 11788 1313 11846 1371 sw
rect 11736 1261 11742 1313
rect 11794 1261 11806 1313
rect 11858 1261 11864 1313
rect 12214 1060 12266 2497
rect 12464 1098 12784 2727
rect 13428 2172 13434 2288
rect 13550 2172 13556 2288
rect 12880 1563 12932 1569
rect 12880 1499 12932 1511
rect 12880 1070 12932 1447
rect 13272 1261 13278 1313
rect 13330 1261 13342 1313
rect 13394 1261 13400 1313
tri 13272 1185 13348 1261 ne
tri 12932 1070 12944 1082 sw
rect 12880 1060 12944 1070
tri 12880 1048 12892 1060 ne
tri 11672 437 11850 615 sw
tri 11356 126 11377 147 sw
rect 11304 110 11377 126
tri 11377 110 11393 126 sw
rect 11304 98 11393 110
tri 11393 98 11405 110 sw
rect 11304 92 11405 98
tri 11405 92 11411 98 sw
rect 11304 40 11310 92
rect 11362 40 11374 92
rect 11426 40 11432 92
rect 11492 -103 11850 437
rect 12892 0 12944 1060
rect 13348 -1988 13400 1261
rect 13428 0 13556 2172
rect 13584 1058 13636 2917
tri 13636 2879 13674 2917 nw
rect 13766 2281 14011 3003
rect 13766 2165 13796 2281
rect 13976 2165 14011 2281
tri 13695 1898 13766 1969 se
rect 13766 1552 14011 2165
tri 14011 1552 14149 1690 sw
rect 13766 1523 14149 1552
tri 13766 1460 13829 1523 ne
rect 13829 1088 14149 1523
tri 13695 1080 13703 1088 ne
rect 13703 1080 14149 1088
tri 13584 1035 13607 1058 ne
rect 13607 1035 13636 1058
tri 13636 1035 13681 1080 sw
tri 13703 1035 13748 1080 ne
rect 13748 1035 14149 1080
tri 13607 1006 13636 1035 ne
rect 13636 1021 13681 1035
tri 13681 1021 13695 1035 sw
tri 13748 1021 13762 1035 ne
rect 13762 1021 14149 1035
rect 13636 1006 13695 1021
tri 13636 989 13653 1006 ne
rect 13653 989 13695 1006
tri 13695 989 13727 1021 sw
tri 13762 989 13794 1021 ne
rect 13794 989 14149 1021
tri 13653 961 13681 989 ne
rect 13681 961 13727 989
tri 13727 961 13755 989 sw
tri 13681 954 13688 961 ne
rect 13688 954 13755 961
tri 13794 954 13829 989 ne
tri 13688 939 13703 954 ne
rect 13606 162 13658 168
rect 13606 98 13658 110
rect 13606 40 13658 46
rect 13348 -2052 13400 -2040
rect 13348 -2110 13400 -2104
rect 13606 -1988 13658 -1982
rect 13606 -2052 13658 -2040
rect 6816 -5196 6822 -5144
rect 6874 -5196 6886 -5144
rect 6938 -5196 6944 -5144
rect 13606 -5222 13658 -2104
rect 13703 -5105 13755 954
rect 13829 17 14149 989
rect 13703 -5157 13709 -5105
rect 13761 -5157 13776 -5105
rect 13828 -5157 13834 -5105
tri 13658 -5222 13680 -5200 sw
tri 13606 -5296 13680 -5222 ne
tri 13680 -5291 13749 -5222 sw
rect 13680 -5296 13749 -5291
tri 13749 -5296 13754 -5291 sw
tri 13680 -5365 13749 -5296 ne
rect 13749 -5343 13754 -5296
tri 13754 -5343 13801 -5296 sw
rect 13749 -5613 13801 -5343
<< via2 >>
rect 6253 4018 6302 4068
rect 6302 4018 6309 4068
rect 6353 4018 6380 4068
rect 6380 4018 6405 4068
rect 6405 4018 6409 4068
rect 6453 4018 6457 4068
rect 6457 4018 6482 4068
rect 6482 4018 6509 4068
rect 6552 4018 6559 4068
rect 6559 4018 6608 4068
rect 6253 4012 6309 4018
rect 6353 4012 6409 4018
rect 6453 4012 6509 4018
rect 6552 4012 6608 4018
rect 6253 3944 6302 3972
rect 6302 3944 6309 3972
rect 6353 3944 6380 3972
rect 6380 3944 6405 3972
rect 6405 3944 6409 3972
rect 6453 3944 6457 3972
rect 6457 3944 6482 3972
rect 6482 3944 6509 3972
rect 6552 3944 6559 3972
rect 6559 3944 6608 3972
rect 6253 3922 6309 3944
rect 6353 3922 6409 3944
rect 6453 3922 6509 3944
rect 6552 3922 6608 3944
rect 6253 3916 6302 3922
rect 6302 3916 6309 3922
rect 6353 3916 6380 3922
rect 6380 3916 6405 3922
rect 6405 3916 6409 3922
rect 6453 3916 6457 3922
rect 6457 3916 6482 3922
rect 6482 3916 6509 3922
rect 6552 3916 6559 3922
rect 6559 3916 6608 3922
rect 6253 3870 6302 3876
rect 6302 3870 6309 3876
rect 6353 3870 6380 3876
rect 6380 3870 6405 3876
rect 6405 3870 6409 3876
rect 6453 3870 6457 3876
rect 6457 3870 6482 3876
rect 6482 3870 6509 3876
rect 6552 3870 6559 3876
rect 6559 3870 6608 3876
rect 6253 3848 6309 3870
rect 6353 3848 6409 3870
rect 6453 3848 6509 3870
rect 6552 3848 6608 3870
rect 6253 3820 6302 3848
rect 6302 3820 6309 3848
rect 6353 3820 6380 3848
rect 6380 3820 6405 3848
rect 6405 3820 6409 3848
rect 6453 3820 6457 3848
rect 6457 3820 6482 3848
rect 6482 3820 6509 3848
rect 6552 3820 6559 3848
rect 6559 3820 6608 3848
rect 6253 3774 6309 3780
rect 6353 3774 6409 3780
rect 6453 3774 6509 3780
rect 6552 3774 6608 3780
rect 6253 3724 6302 3774
rect 6302 3724 6309 3774
rect 6353 3724 6380 3774
rect 6380 3724 6405 3774
rect 6405 3724 6409 3774
rect 6453 3724 6457 3774
rect 6457 3724 6482 3774
rect 6482 3724 6509 3774
rect 6552 3724 6559 3774
rect 6559 3724 6608 3774
rect 7353 1425 7409 1481
rect 7433 1425 7489 1481
rect 7353 1339 7409 1395
rect 7433 1339 7489 1395
rect 7353 1252 7409 1308
rect 7433 1252 7489 1308
rect 7585 1252 7641 1308
rect 7353 1165 7409 1221
rect 7433 1165 7489 1221
rect 7585 1165 7641 1221
rect 7353 1078 7409 1134
rect 7433 1078 7489 1134
rect 7585 1078 7641 1134
<< metal3 >>
rect 6248 4068 6613 4075
rect 6248 4012 6253 4068
rect 6309 4012 6353 4068
rect 6409 4012 6453 4068
rect 6509 4012 6552 4068
rect 6608 4012 6613 4068
rect 6248 3972 6613 4012
rect 6248 3916 6253 3972
rect 6309 3916 6353 3972
rect 6409 3916 6453 3972
rect 6509 3916 6552 3972
rect 6608 3916 6613 3972
rect 6248 3876 6613 3916
rect 6248 3820 6253 3876
rect 6309 3820 6353 3876
rect 6409 3820 6453 3876
rect 6509 3820 6552 3876
rect 6608 3820 6613 3876
rect 6248 3780 6613 3820
rect 6248 3724 6253 3780
rect 6309 3724 6353 3780
rect 6409 3724 6453 3780
rect 6509 3724 6552 3780
rect 6608 3724 6613 3780
rect 6248 3717 6613 3724
rect 7328 1481 7514 1486
rect 7328 1425 7353 1481
rect 7409 1425 7433 1481
rect 7489 1425 7514 1481
rect 7328 1395 7514 1425
rect 7328 1339 7353 1395
rect 7409 1339 7433 1395
rect 7489 1339 7514 1395
rect 7328 1308 7514 1339
rect 7328 1252 7353 1308
rect 7409 1252 7433 1308
rect 7489 1252 7514 1308
rect 7328 1221 7514 1252
rect 7328 1165 7353 1221
rect 7409 1165 7433 1221
rect 7489 1165 7514 1221
rect 7328 1134 7514 1165
rect 7328 1078 7353 1134
rect 7409 1078 7433 1134
rect 7489 1078 7514 1134
rect 7328 1073 7514 1078
rect 7545 1308 7681 1313
rect 7545 1252 7585 1308
rect 7641 1252 7681 1308
rect 7545 1221 7681 1252
rect 7545 1165 7585 1221
rect 7641 1165 7681 1221
rect 7545 1134 7681 1165
rect 7545 1078 7585 1134
rect 7641 1078 7681 1134
rect 7545 1073 7681 1078
<< comment >>
rect 0 814 3503 1104
tri 3503 814 3793 1104 sw
tri 14307 814 14597 1104 se
rect 14597 814 15000 1104
rect 0 112 4367 814
tri 4367 112 5069 814 sw
rect 0 0 5069 112
tri 13895 402 14307 814 se
rect 14307 402 15000 814
rect 13895 0 15000 402
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1707688321
transform -1 0 8113 0 1 1722
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1707688321
transform 0 -1 12284 1 0 2170
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1707688321
transform 0 -1 8770 1 0 2170
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1707688321
transform 0 -1 8080 1 0 2170
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1707688321
transform 0 -1 4566 1 0 2170
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1707688321
transform 0 -1 3876 1 0 2170
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1707688321
transform 0 -1 376 1 0 2170
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1707688321
transform 0 -1 17 1 0 3089
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1707688321
transform 0 -1 1613 1 0 3089
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_2
timestamp 1707688321
transform 0 -1 2625 1 0 3089
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_3
timestamp 1707688321
transform 0 -1 3589 1 0 3089
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_4
timestamp 1707688321
transform 0 -1 4853 1 0 3089
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_5
timestamp 1707688321
transform 0 -1 5817 1 0 3089
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_6
timestamp 1707688321
transform 0 -1 6829 1 0 3089
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_7
timestamp 1707688321
transform 0 -1 8425 1 0 3089
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_8
timestamp 1707688321
transform 0 -1 7793 1 0 3089
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_9
timestamp 1707688321
transform 0 -1 9057 1 0 3089
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_10
timestamp 1707688321
transform 0 -1 10021 1 0 3089
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_11
timestamp 1707688321
transform 0 -1 11033 1 0 3089
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_12
timestamp 1707688321
transform 0 -1 11997 1 0 3089
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_13
timestamp 1707688321
transform 0 -1 649 1 0 3089
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_14
timestamp 1707688321
transform 0 -1 15017 1 0 3089
box 0 0 1 1
use L1M1_CDNS_52468879185193  L1M1_CDNS_52468879185193_0
timestamp 1707688321
transform 1 0 731 0 1 1586
box 0 0 1 1
use L1M1_CDNS_52468879185941  L1M1_CDNS_52468879185941_0
timestamp 1707688321
transform 1 0 3790 0 1 191
box -12 -6 1990 40
use L1M1_CDNS_52468879185945  L1M1_CDNS_52468879185945_0
timestamp 1707688321
transform 1 0 8740 0 1 191
box -12 -6 1846 40
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1707688321
transform 0 -1 6728 -1 0 2623
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1707688321
transform 0 -1 10140 -1 0 2623
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1707688321
transform 0 -1 2920 -1 0 2625
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1707688321
transform 0 -1 8316 -1 0 2935
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1707688321
transform 0 -1 978 -1 0 1900
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_5
timestamp 1707688321
transform 0 -1 1732 -1 0 1900
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_6
timestamp 1707688321
transform 0 -1 649 -1 0 1035
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_7
timestamp 1707688321
transform 0 -1 3867 -1 0 1006
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_8
timestamp 1707688321
transform 0 -1 4379 -1 0 2969
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_9
timestamp 1707688321
transform 0 -1 4461 -1 0 1376
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_10
timestamp 1707688321
transform -1 0 5102 0 1 768
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_11
timestamp 1707688321
transform -1 0 299 0 1 1574
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_12
timestamp 1707688321
transform -1 0 5776 0 1 3502
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_13
timestamp 1707688321
transform -1 0 5936 0 1 216
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_14
timestamp 1707688321
transform -1 0 3683 0 1 2917
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_15
timestamp 1707688321
transform -1 0 5780 0 1 185
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_16
timestamp 1707688321
transform -1 0 10060 0 1 185
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_17
timestamp 1707688321
transform -1 0 6724 0 -1 2933
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_18
timestamp 1707688321
transform -1 0 7948 0 -1 1688
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_19
timestamp 1707688321
transform -1 0 8683 0 -1 268
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_20
timestamp 1707688321
transform -1 0 1572 0 -1 313
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_21
timestamp 1707688321
transform -1 0 8104 0 -1 1777
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_22
timestamp 1707688321
transform 0 1 1680 1 0 2495
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_23
timestamp 1707688321
transform 0 1 1364 1 0 3486
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_24
timestamp 1707688321
transform 0 -1 398 1 0 907
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_25
timestamp 1707688321
transform 0 -1 223 1 0 3307
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_26
timestamp 1707688321
transform 0 -1 2055 1 0 3307
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_27
timestamp 1707688321
transform 0 -1 8806 1 0 2159
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_28
timestamp 1707688321
transform 0 -1 11470 1 0 2419
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_29
timestamp 1707688321
transform 0 -1 11356 1 0 2495
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_30
timestamp 1707688321
transform 0 -1 2368 1 0 2495
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_31
timestamp 1707688321
transform 0 -1 2368 1 0 1577
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_32
timestamp 1707688321
transform 0 -1 5936 1 0 2495
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_33
timestamp 1707688321
transform 0 -1 143 1 0 2807
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_34
timestamp 1707688321
transform 0 -1 1652 1 0 1488
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_35
timestamp 1707688321
transform 0 -1 1652 1 0 185
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_36
timestamp 1707688321
transform 0 -1 3683 1 0 1026
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_37
timestamp 1707688321
transform 0 -1 3947 1 0 1026
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_38
timestamp 1707688321
transform 0 -1 649 1 0 2159
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_39
timestamp 1707688321
transform 0 -1 398 1 0 2159
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_40
timestamp 1707688321
transform 1 0 10880 0 -1 3554
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_41
timestamp 1707688321
transform 1 0 2236 0 -1 1540
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_42
timestamp 1707688321
transform 1 0 2792 0 -1 2380
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_43
timestamp 1707688321
transform 1 0 9599 0 1 688
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_44
timestamp 1707688321
transform 1 0 2396 0 1 878
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_45
timestamp 1707688321
transform 1 0 8264 0 1 384
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_46
timestamp 1707688321
transform 1 0 9367 0 1 2917
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_47
timestamp 1707688321
transform 1 0 11148 0 1 2997
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_48
timestamp 1707688321
transform 1 0 2396 0 1 384
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_49
timestamp 1707688321
transform 1 0 91 0 1 384
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_50
timestamp 1707688321
transform 1 0 9599 0 1 185
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_51
timestamp 1707688321
transform 1 0 4805 0 1 185
box 0 0 1 1
use M1M2_CDNS_52468879185197  M1M2_CDNS_52468879185197_0
timestamp 1707688321
transform 0 1 9110 -1 0 1181
box 0 0 256 116
use M1M2_CDNS_52468879185197  M1M2_CDNS_52468879185197_1
timestamp 1707688321
transform 0 1 11040 -1 0 1181
box 0 0 256 116
use M1M2_CDNS_52468879185197  M1M2_CDNS_52468879185197_2
timestamp 1707688321
transform 0 -1 4927 1 0 479
box 0 0 256 116
use M1M2_CDNS_52468879185197  M1M2_CDNS_52468879185197_3
timestamp 1707688321
transform 1 0 13457 0 -1 4069
box 0 0 256 116
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_0
timestamp 1707688321
transform 0 -1 5776 -1 0 2120
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_1
timestamp 1707688321
transform 0 -1 5776 -1 0 1181
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_2
timestamp 1707688321
transform 0 1 6756 -1 0 2120
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_3
timestamp 1707688321
transform 0 1 6756 -1 0 1181
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_4
timestamp 1707688321
transform 0 1 9110 -1 0 2120
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_5
timestamp 1707688321
transform 0 1 11040 -1 0 2120
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_6
timestamp 1707688321
transform 0 1 4416 -1 0 3274
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_7
timestamp 1707688321
transform 0 1 437 -1 0 659
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_8
timestamp 1707688321
transform 0 1 436 -1 0 3273
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_9
timestamp 1707688321
transform 0 -1 2668 1 0 479
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_10
timestamp 1707688321
transform 0 -1 9721 1 0 479
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_11
timestamp 1707688321
transform 1 0 126 0 -1 4070
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_12
timestamp 1707688321
transform 1 0 5348 0 -1 2282
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_13
timestamp 1707688321
transform 1 0 13790 0 1 2165
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_0
timestamp 1707688321
transform 0 -1 554 -1 0 1035
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_1
timestamp 1707688321
transform -1 0 1572 0 1 2161
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_2
timestamp 1707688321
transform 0 1 2552 1 0 2158
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_3
timestamp 1707688321
transform 0 1 9599 1 0 2159
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_4
timestamp 1707688321
transform 1 0 4805 0 -1 2282
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_5
timestamp 1707688321
transform 1 0 8344 0 1 2165
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_6
timestamp 1707688321
transform 1 0 8344 0 1 694
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_7
timestamp 1707688321
transform 1 0 13428 0 1 2172
box 0 0 1 1
use M1M2_CDNS_52468879185201  M1M2_CDNS_52468879185201_0
timestamp 1707688321
transform 1 0 1010 0 -1 1355
box 0 0 320 116
use M1M2_CDNS_52468879185201  M1M2_CDNS_52468879185201_1
timestamp 1707688321
transform 1 0 3981 0 1 2165
box 0 0 320 116
use M1M2_CDNS_52468879185201  M1M2_CDNS_52468879185201_2
timestamp 1707688321
transform 1 0 12464 0 1 2165
box 0 0 320 116
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_0
timestamp 1707688321
transform -1 0 4301 0 1 185
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_1
timestamp 1707688321
transform 1 0 3981 0 -1 3049
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_2
timestamp 1707688321
transform 1 0 12464 0 -1 2779
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_3
timestamp 1707688321
transform 1 0 12464 0 -1 3049
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_0
timestamp 1707688321
transform 0 -1 398 -1 0 659
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_1
timestamp 1707688321
transform 0 -1 1652 -1 0 1119
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_2
timestamp 1707688321
transform 0 -1 649 -1 0 659
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_3
timestamp 1707688321
transform 0 -1 4605 1 0 472
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_4
timestamp 1707688321
transform 0 -1 649 1 0 3081
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_5
timestamp 1707688321
transform 0 -1 3787 1 0 468
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_6
timestamp 1707688321
transform 1 0 1773 0 1 1408
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_7
timestamp 1707688321
transform 1 0 5348 0 1 185
box 0 0 1 1
use M1M2_CDNS_52468879185208  M1M2_CDNS_52468879185208_0
timestamp 1707688321
transform 0 -1 9028 -1 0 659
box 0 0 192 244
use M1M2_CDNS_52468879185208  M1M2_CDNS_52468879185208_1
timestamp 1707688321
transform 0 1 2948 -1 0 1345
box 0 0 192 244
use M1M2_CDNS_52468879185208  M1M2_CDNS_52468879185208_2
timestamp 1707688321
transform 0 1 2948 -1 0 3921
box 0 0 192 244
use M1M2_CDNS_52468879185208  M1M2_CDNS_52468879185208_3
timestamp 1707688321
transform 0 -1 9325 1 0 479
box 0 0 192 244
use M1M2_CDNS_52468879185209  M1M2_CDNS_52468879185209_0
timestamp 1707688321
transform 0 1 11032 -1 0 2286
box 0 0 128 244
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_0
timestamp 1707688321
transform 0 -1 10060 1 0 475
box 0 0 1 1
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_1
timestamp 1707688321
transform 1 0 4022 0 1 694
box 0 0 1 1
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_2
timestamp 1707688321
transform 1 0 9075 0 1 694
box 0 0 1 1
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_3
timestamp 1707688321
transform 1 0 9075 0 1 185
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_0
timestamp 1707688321
transform 0 1 4409 1 0 1479
box 0 0 1 1
use M1M2_CDNS_52468879185967  M1M2_CDNS_52468879185967_0
timestamp 1707688321
transform 1 0 1525 0 -1 4069
box 0 0 448 116
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_0
timestamp 1707688321
transform 0 -1 11672 -1 0 2120
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_1
timestamp 1707688321
transform 0 -1 1635 1 0 479
box 0 0 192 180
use M1M2_CDNS_524688791851032  M1M2_CDNS_524688791851032_0
timestamp 1707688321
transform 0 1 8010 -1 0 3273
box 0 0 192 372
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_0
timestamp 1707688321
transform 1 0 6983 0 -1 3267
box 0 0 320 180
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_1
timestamp 1707688321
transform 1 0 1011 0 -1 3914
box 0 0 320 180
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_2
timestamp 1707688321
transform 1 0 12464 0 1 3085
box 0 0 320 180
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_3
timestamp 1707688321
transform 1 0 6225 0 1 1938
box 0 0 320 180
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_4
timestamp 1707688321
transform 1 0 3981 0 1 3089
box 0 0 320 180
use M1M2_CDNS_524688791851081  M1M2_CDNS_524688791851081_0
timestamp 1707688321
transform 0 -1 5534 1 0 479
box 0 0 256 180
use M1M2_CDNS_524688791851175  M1M2_CDNS_524688791851175_0
timestamp 1707688321
transform 0 -1 7299 1 0 2159
box 0 0 128 308
use M1M2_CDNS_524688791851176  M1M2_CDNS_524688791851176_0
timestamp 1707688321
transform 0 1 10296 -1 0 1181
box 0 0 256 308
use M1M2_CDNS_524688791851185  M1M2_CDNS_524688791851185_0
timestamp 1707688321
transform 1 0 6225 0 -1 1177
box 0 0 320 244
use M1M2_CDNS_524688791851186  M1M2_CDNS_524688791851186_0
timestamp 1707688321
transform 0 -1 10767 -1 0 3921
box 0 0 192 308
use M1M2_CDNS_524688791851186  M1M2_CDNS_524688791851186_1
timestamp 1707688321
transform 0 -1 14808 -1 0 3921
box 0 0 192 308
use M1M2_CDNS_524688791851186  M1M2_CDNS_524688791851186_2
timestamp 1707688321
transform 0 1 10296 -1 0 2126
box 0 0 192 308
use M1M2_CDNS_524688791851186  M1M2_CDNS_524688791851186_3
timestamp 1707688321
transform 0 -1 4294 1 0 479
box 0 0 192 308
use M1M2_CDNS_524688791851187  M1M2_CDNS_524688791851187_0
timestamp 1707688321
transform 1 0 7008 0 -1 652
box 0 0 768 180
use M1M2_CDNS_524688791851188  M1M2_CDNS_524688791851188_0
timestamp 1707688321
transform 1 0 11418 0 -1 4069
box 0 0 512 116
use M2M3_CDNS_524688791851179  M2M3_CDNS_524688791851179_0
timestamp 1707688321
transform 1 0 347 0 1 1098
box -5 0 301 314
use M2M3_CDNS_524688791851180  M2M3_CDNS_524688791851180_0
timestamp 1707688321
transform 1 0 3993 0 1 1054
box -5 0 301 714
use M2M3_CDNS_524688791851181  M2M3_CDNS_524688791851181_0
timestamp 1707688321
transform 1 0 12214 0 1 1060
box -5 0 61 634
use M2M3_CDNS_524688791851181  M2M3_CDNS_524688791851181_1
timestamp 1707688321
transform 1 0 8754 0 1 1060
box -5 0 61 634
use M2M3_CDNS_524688791851181  M2M3_CDNS_524688791851181_2
timestamp 1707688321
transform 1 0 4553 0 1 1060
box -5 0 61 634
use M2M3_CDNS_524688791851181  M2M3_CDNS_524688791851181_3
timestamp 1707688321
transform 1 0 3735 0 1 1060
box -5 0 61 634
use M2M3_CDNS_524688791851182  M2M3_CDNS_524688791851182_0
timestamp 1707688321
transform 1 0 12475 0 1 1098
box -5 0 301 794
use M2M3_CDNS_524688791851183  M2M3_CDNS_524688791851183_0
timestamp 1707688321
transform 1 0 13466 0 1 1098
box -5 0 61 794
use M2M3_CDNS_524688791851183  M2M3_CDNS_524688791851183_1
timestamp 1707688321
transform 1 0 9637 0 1 1098
box -5 0 61 794
use M2M3_CDNS_524688791851183  M2M3_CDNS_524688791851183_2
timestamp 1707688321
transform 1 0 8382 0 1 1098
box -5 0 61 794
use M2M3_CDNS_524688791851183  M2M3_CDNS_524688791851183_3
timestamp 1707688321
transform 1 0 4843 0 1 1098
box -5 0 61 794
use M2M3_CDNS_524688791851183  M2M3_CDNS_524688791851183_4
timestamp 1707688321
transform 1 0 2585 0 1 1098
box -5 0 61 794
use M2M3_CDNS_524688791851184  M2M3_CDNS_524688791851184_0
timestamp 1707688321
transform 1 0 5380 0 1 1098
box -5 0 141 794
use M2M3_CDNS_524688791851184  M2M3_CDNS_524688791851184_1
timestamp 1707688321
transform 1 0 1480 0 1 1098
box -5 0 141 794
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_0
timestamp 1707688321
transform 1 0 987 0 1 3780
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_1
timestamp 1707688321
transform 1 0 6203 0 1 2422
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_2
timestamp 1707688321
transform 1 0 14447 0 1 3780
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_3
timestamp 1707688321
transform 1 0 13671 0 1 1064
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_4
timestamp 1707688321
transform 1 0 10927 0 1 3780
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_5
timestamp 1707688321
transform 1 0 10427 0 1 3780
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_6
timestamp 1707688321
transform 1 0 10272 0 1 2422
box 0 0 364 858
use sky130_fd_io__sio_com_m2m3_strap  sky130_fd_io__sio_com_m2m3_strap_7
timestamp 1707688321
transform 1 0 6961 0 1 1064
box 0 0 364 858
use sky130_fd_io__sio_ctl_hld  sky130_fd_io__sio_ctl_hld_0
timestamp 1707688321
transform -1 0 8654 0 -1 1717
box -6668 -2440 8211 1555
use sky130_fd_io__sio_ctl_lsbank  sky130_fd_io__sio_ctl_lsbank_0
timestamp 1707688321
transform 1 0 0 0 1 1838
box -53 -96 15043 2388
use sky130_fd_io__sio_hvsbt_endcap  sky130_fd_io__sio_hvsbt_endcap_0
timestamp 1707688321
transform -1 0 11055 0 1 323
box -84 93 164 1337
<< labels >>
flabel comment s 11325 69 11325 69 0 FreeSans 200 90 0 0 vpwr_ka
flabel comment s 11325 4080 11325 4080 0 FreeSans 200 90 0 0 vpwr_ka
flabel comment s 12832 4080 12832 4080 0 FreeSans 200 90 0 0 vpb_ka
flabel comment s 12832 64 12832 64 0 FreeSans 200 90 0 0 vpb_ka
flabel comment s 6411 17 6411 17 0 FreeSans 200 0 0 0 vccio
flabel comment s 1384 4084 1384 4084 0 FreeSans 200 90 0 0 slow
flabel comment s 2258 4076 2258 4076 0 FreeSans 200 90 0 0 od_h
flabel comment s 8744 81 8744 81 0 FreeSans 200 90 0 0 dm_h<0>
flabel comment s 8529 4048 8529 4048 0 FreeSans 200 90 0 0 dm_h<0>
flabel comment s 14090 4078 14090 4078 0 FreeSans 200 0 0 0 vgnd
flabel comment s 13741 4078 13741 4078 0 FreeSans 200 0 0 0 vgnd
flabel comment s 2141 19 2141 19 0 FreeSans 200 180 0 0 pad
flabel comment s 2141 4107 2141 4107 0 FreeSans 200 180 0 0 pad
flabel comment s 3982 3598 3982 3598 0 FreeSans 200 0 0 0 slow
flabel comment s 257 1600 257 1600 0 FreeSans 200 0 0 0 hld_i_vpwr
flabel comment s 14453 186 14453 186 0 FreeSans 1000 0 0 0 Well Keepout
flabel comment s 920 494 920 494 0 FreeSans 1000 0 0 0 Well Keepout
flabel metal1 s 14680 3077 14714 3279 3 FreeSans 400 180 0 0 vgnd
port 2 nsew
flabel metal1 s 12612 3077 12646 3279 7 FreeSans 400 180 0 0 vgnd
port 2 nsew
flabel metal1 s 14680 2158 14714 2288 3 FreeSans 400 180 0 0 vgnd
port 2 nsew
flabel metal1 s 14697 3178 14697 3178 3 FreeSans 400 180 0 0 vgnd
flabel metal1 s 8310 464 8327 666 3 FreeSans 400 180 0 0 vgnd
port 2 nsew
flabel metal1 s 14697 3178 14697 3178 3 FreeSans 400 180 0 0 vgnd
flabel metal1 s 12629 3178 12629 3178 7 FreeSans 400 180 0 0 vgnd
flabel metal1 s 10831 2501 10865 2535 0 FreeSans 400 0 0 0 inp_dis_h_n
port 3 nsew
flabel metal1 s 14697 2223 14697 2223 3 FreeSans 400 180 0 0 vgnd
flabel metal1 s 8318 565 8318 565 3 FreeSans 400 180 0 0 vgnd
flabel metal1 s 0 2158 34 2288 3 FreeSans 400 0 0 0 vgnd
port 2 nsew
flabel metal1 s 14697 2223 14697 2223 3 FreeSans 400 180 0 0 vgnd
flabel metal1 s 12629 3178 12629 3178 7 FreeSans 400 180 0 0 vgnd
flabel metal1 s 0 3077 34 3279 3 FreeSans 400 0 0 0 vgnd
port 2 nsew
flabel metal1 s 17 3178 17 3178 3 FreeSans 400 0 0 0 vgnd
flabel metal1 s 14966 2158 15000 2288 3 FreeSans 400 180 0 0 vgnd
port 2 nsew
flabel metal1 s 12629 3178 12629 3178 7 FreeSans 400 180 0 0 vgnd
flabel metal1 s 14697 3178 14697 3178 3 FreeSans 400 180 0 0 vgnd
flabel metal1 s 14697 2223 14697 2223 3 FreeSans 400 180 0 0 vgnd
flabel metal1 s 17 2223 17 2223 3 FreeSans 400 0 0 0 vgnd
flabel metal1 s 9687 777 9846 806 3 FreeSans 520 180 0 0 od_i_h
port 7 nsew
flabel metal1 s 12695 2890 12764 2925 3 FreeSans 520 180 0 0 hld_ovr
port 9 nsew
flabel metal1 s 10249 1261 10368 1311 3 FreeSans 520 180 0 0 hld_i_ovr_h
port 5 nsew
flabel metal1 s 14983 2223 14983 2223 3 FreeSans 400 180 0 0 vgnd
flabel metal1 s 11268 2540 11336 2602 3 FreeSans 520 0 0 0 inp_dis_h
port 6 nsew
flabel metal1 s 12479 2887 12513 2921 0 FreeSans 400 0 0 0 inp_dis
port 10 nsew
flabel metal1 s 14966 3077 15000 3279 7 FreeSans 400 0 0 0 vgnd
port 2 nsew
flabel metal1 s 14966 1928 15000 2130 7 FreeSans 400 0 0 0 vcc_io
port 4 nsew
flabel metal1 s 17 3183 17 3183 3 FreeSans 400 0 0 0 vgnd
flabel metal1 s 0 1928 34 2130 3 FreeSans 400 0 0 0 vcc_io
port 4 nsew
flabel metal1 s 10344 384 10379 436 7 FreeSans 200 0 0 0 ibuf_sel
port 8 nsew
flabel locali s 8458 1644 8573 1682 3 FreeSans 520 180 0 0 enable_h
port 11 nsew
flabel metal2 s 7976 0 8028 43 3 FreeSans 200 90 0 0 hld_h_n
port 12 nsew
flabel metal2 s 1680 0 1732 46 3 FreeSans 200 90 0 0 dm_h_n<0>
port 13 nsew
flabel metal2 s 8631 0 8683 46 7 FreeSans 200 270 0 0 dm_h_n<2>
port 14 nsew
flabel metal2 s 7896 0 7948 43 8 FreeSans 200 270 0 0 dm_h_n<1>
port 15 nsew
flabel metal2 s 926 4052 978 4098 3 FreeSans 200 270 0 0 dm_h_n<0>
port 13 nsew
flabel metal2 s 10088 0 10140 46 3 FreeSans 200 90 0 0 vtrip_sel_h_n
port 16 nsew
flabel metal2 s 9519 0 9571 46 3 FreeSans 200 90 0 0 vtrip_sel
port 17 nsew
flabel metal2 s 1006 4096 1336 4141 0 FreeSans 200 0 0 0 vpwr
port 18 nsew
flabel metal2 s 6676 0 6728 46 3 FreeSans 200 90 0 0 ibuf_sel_h_n
port 19 nsew
flabel metal2 s 6596 0 6648 46 3 FreeSans 200 90 0 0 ibuf_sel_h
port 20 nsew
flabel metal2 s 2003 4115 2055 4156 7 FreeSans 200 90 0 0 hld_i_vpwr
port 21 nsew
flabel metal2 s 5884 4095 5936 4141 7 FreeSans 200 90 0 0 dm_h_n<2>
port 14 nsew
flabel metal2 s 2316 4098 2368 4141 8 FreeSans 200 90 0 0 dm_h_n<1>
port 15 nsew
flabel metal2 s 4329 0 4381 43 3 FreeSans 200 90 0 0 dm<2>
port 22 nsew
flabel metal2 s 3895 0 3947 43 3 FreeSans 200 90 0 0 dm<1>
port 23 nsew
flabel metal2 s 3815 0 3867 43 3 FreeSans 200 90 0 0 dm<0>
port 24 nsew
flabel metal2 s 5648 4095 5700 4141 7 FreeSans 200 90 0 0 dm_h<2>
port 25 nsew
flabel metal2 s 2868 2328 2920 2371 7 FreeSans 200 270 0 0 dm_h<1>
port 26 nsew
flabel metal2 s 9833 0 9885 46 3 FreeSans 200 90 0 0 vtrip_sel_h
port 27 nsew
flabel metal2 s 5050 4103 5102 4141 3 FreeSans 400 270 0 0 hld_i_h_n
port 28 nsew
flabel metal2 s 10880 0 10932 46 3 FreeSans 200 90 0 0 dm_h<2>
port 25 nsew
flabel metal2 s 2552 4098 2604 4141 3 FreeSans 200 270 0 0 dm_h<1>
port 26 nsew
flabel metal2 s 1444 4098 1496 4141 7 FreeSans 200 90 0 0 dm_h<0>
port 29 nsew
<< properties >>
string GDS_END 85498572
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85426428
string path 156.200 97.400 165.325 97.400 
<< end >>
