magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -26 -26 82 2026
<< ndiff >>
rect 0 1950 56 2000
rect 0 1916 11 1950
rect 45 1916 56 1950
rect 0 1882 56 1916
rect 0 1848 11 1882
rect 45 1848 56 1882
rect 0 1814 56 1848
rect 0 1780 11 1814
rect 45 1780 56 1814
rect 0 1746 56 1780
rect 0 1712 11 1746
rect 45 1712 56 1746
rect 0 1678 56 1712
rect 0 1644 11 1678
rect 45 1644 56 1678
rect 0 1610 56 1644
rect 0 1576 11 1610
rect 45 1576 56 1610
rect 0 1542 56 1576
rect 0 1508 11 1542
rect 45 1508 56 1542
rect 0 1474 56 1508
rect 0 1440 11 1474
rect 45 1440 56 1474
rect 0 1406 56 1440
rect 0 1372 11 1406
rect 45 1372 56 1406
rect 0 1338 56 1372
rect 0 1304 11 1338
rect 45 1304 56 1338
rect 0 1270 56 1304
rect 0 1236 11 1270
rect 45 1236 56 1270
rect 0 1202 56 1236
rect 0 1168 11 1202
rect 45 1168 56 1202
rect 0 1134 56 1168
rect 0 1100 11 1134
rect 45 1100 56 1134
rect 0 1066 56 1100
rect 0 1032 11 1066
rect 45 1032 56 1066
rect 0 998 56 1032
rect 0 964 11 998
rect 45 964 56 998
rect 0 930 56 964
rect 0 896 11 930
rect 45 896 56 930
rect 0 862 56 896
rect 0 828 11 862
rect 45 828 56 862
rect 0 794 56 828
rect 0 760 11 794
rect 45 760 56 794
rect 0 726 56 760
rect 0 692 11 726
rect 45 692 56 726
rect 0 658 56 692
rect 0 624 11 658
rect 45 624 56 658
rect 0 590 56 624
rect 0 556 11 590
rect 45 556 56 590
rect 0 522 56 556
rect 0 488 11 522
rect 45 488 56 522
rect 0 454 56 488
rect 0 420 11 454
rect 45 420 56 454
rect 0 386 56 420
rect 0 352 11 386
rect 45 352 56 386
rect 0 318 56 352
rect 0 284 11 318
rect 45 284 56 318
rect 0 250 56 284
rect 0 216 11 250
rect 45 216 56 250
rect 0 182 56 216
rect 0 148 11 182
rect 45 148 56 182
rect 0 114 56 148
rect 0 80 11 114
rect 45 80 56 114
rect 0 46 56 80
rect 0 12 11 46
rect 45 12 56 46
rect 0 0 56 12
<< ndiffc >>
rect 11 1916 45 1950
rect 11 1848 45 1882
rect 11 1780 45 1814
rect 11 1712 45 1746
rect 11 1644 45 1678
rect 11 1576 45 1610
rect 11 1508 45 1542
rect 11 1440 45 1474
rect 11 1372 45 1406
rect 11 1304 45 1338
rect 11 1236 45 1270
rect 11 1168 45 1202
rect 11 1100 45 1134
rect 11 1032 45 1066
rect 11 964 45 998
rect 11 896 45 930
rect 11 828 45 862
rect 11 760 45 794
rect 11 692 45 726
rect 11 624 45 658
rect 11 556 45 590
rect 11 488 45 522
rect 11 420 45 454
rect 11 352 45 386
rect 11 284 45 318
rect 11 216 45 250
rect 11 148 45 182
rect 11 80 45 114
rect 11 12 45 46
<< locali >>
rect 11 1902 45 1916
rect 11 1830 45 1848
rect 11 1758 45 1780
rect 11 1686 45 1712
rect 11 1614 45 1644
rect 11 1542 45 1576
rect 11 1474 45 1508
rect 11 1406 45 1436
rect 11 1338 45 1364
rect 11 1270 45 1292
rect 11 1202 45 1220
rect 11 1134 45 1148
rect 11 1066 45 1076
rect 11 998 45 1004
rect 11 930 45 932
rect 11 894 45 896
rect 11 822 45 828
rect 11 750 45 760
rect 11 678 45 692
rect 11 606 45 624
rect 11 534 45 556
rect 11 462 45 488
rect 11 390 45 420
rect 11 318 45 352
rect 11 250 45 284
rect 11 182 45 212
rect 11 114 45 140
rect 11 46 45 68
<< viali >>
rect 11 1950 45 1974
rect 11 1940 45 1950
rect 11 1882 45 1902
rect 11 1868 45 1882
rect 11 1814 45 1830
rect 11 1796 45 1814
rect 11 1746 45 1758
rect 11 1724 45 1746
rect 11 1678 45 1686
rect 11 1652 45 1678
rect 11 1610 45 1614
rect 11 1580 45 1610
rect 11 1508 45 1542
rect 11 1440 45 1470
rect 11 1436 45 1440
rect 11 1372 45 1398
rect 11 1364 45 1372
rect 11 1304 45 1326
rect 11 1292 45 1304
rect 11 1236 45 1254
rect 11 1220 45 1236
rect 11 1168 45 1182
rect 11 1148 45 1168
rect 11 1100 45 1110
rect 11 1076 45 1100
rect 11 1032 45 1038
rect 11 1004 45 1032
rect 11 964 45 966
rect 11 932 45 964
rect 11 862 45 894
rect 11 860 45 862
rect 11 794 45 822
rect 11 788 45 794
rect 11 726 45 750
rect 11 716 45 726
rect 11 658 45 678
rect 11 644 45 658
rect 11 590 45 606
rect 11 572 45 590
rect 11 522 45 534
rect 11 500 45 522
rect 11 454 45 462
rect 11 428 45 454
rect 11 386 45 390
rect 11 356 45 386
rect 11 284 45 318
rect 11 216 45 246
rect 11 212 45 216
rect 11 148 45 174
rect 11 140 45 148
rect 11 80 45 102
rect 11 68 45 80
rect 11 12 45 30
rect 11 -4 45 12
<< metal1 >>
rect 5 1974 51 1986
rect 5 1940 11 1974
rect 45 1940 51 1974
rect 5 1902 51 1940
rect 5 1868 11 1902
rect 45 1868 51 1902
rect 5 1830 51 1868
rect 5 1796 11 1830
rect 45 1796 51 1830
rect 5 1758 51 1796
rect 5 1724 11 1758
rect 45 1724 51 1758
rect 5 1686 51 1724
rect 5 1652 11 1686
rect 45 1652 51 1686
rect 5 1614 51 1652
rect 5 1580 11 1614
rect 45 1580 51 1614
rect 5 1542 51 1580
rect 5 1508 11 1542
rect 45 1508 51 1542
rect 5 1470 51 1508
rect 5 1436 11 1470
rect 45 1436 51 1470
rect 5 1398 51 1436
rect 5 1364 11 1398
rect 45 1364 51 1398
rect 5 1326 51 1364
rect 5 1292 11 1326
rect 45 1292 51 1326
rect 5 1254 51 1292
rect 5 1220 11 1254
rect 45 1220 51 1254
rect 5 1182 51 1220
rect 5 1148 11 1182
rect 45 1148 51 1182
rect 5 1110 51 1148
rect 5 1076 11 1110
rect 45 1076 51 1110
rect 5 1038 51 1076
rect 5 1004 11 1038
rect 45 1004 51 1038
rect 5 966 51 1004
rect 5 932 11 966
rect 45 932 51 966
rect 5 894 51 932
rect 5 860 11 894
rect 45 860 51 894
rect 5 822 51 860
rect 5 788 11 822
rect 45 788 51 822
rect 5 750 51 788
rect 5 716 11 750
rect 45 716 51 750
rect 5 678 51 716
rect 5 644 11 678
rect 45 644 51 678
rect 5 606 51 644
rect 5 572 11 606
rect 45 572 51 606
rect 5 534 51 572
rect 5 500 11 534
rect 45 500 51 534
rect 5 462 51 500
rect 5 428 11 462
rect 45 428 51 462
rect 5 390 51 428
rect 5 356 11 390
rect 45 356 51 390
rect 5 318 51 356
rect 5 284 11 318
rect 45 284 51 318
rect 5 246 51 284
rect 5 212 11 246
rect 45 212 51 246
rect 5 174 51 212
rect 5 140 11 174
rect 45 140 51 174
rect 5 102 51 140
rect 5 68 11 102
rect 45 68 51 102
rect 5 30 51 68
rect 5 -4 11 30
rect 45 -4 51 30
rect 5 -16 51 -4
<< properties >>
string GDS_END 21448
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 17540
<< end >>
