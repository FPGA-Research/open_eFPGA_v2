magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -76 -26 1732 2026
<< mvnnmos >>
rect 0 0 800 2000
rect 856 0 1656 2000
<< mvndiff >>
rect -50 0 0 2000
rect 1656 0 1706 2000
<< poly >>
rect 0 2000 800 2026
rect 0 -26 800 0
rect 856 2000 1656 2026
rect 856 -26 1656 0
<< locali >>
rect -45 -4 -11 1966
rect 811 -4 845 1966
rect 1667 -4 1701 1966
use hvDFL1sd2_CDNS_52468879185991  hvDFL1sd2_CDNS_52468879185991_0
timestamp 1707688321
transform 1 0 800 0 1 0
box -26 -26 82 2026
use hvDFL1sd_CDNS_52468879185990  hvDFL1sd_CDNS_52468879185990_0
timestamp 1707688321
transform -1 0 0 0 1 0
box -26 -26 79 2026
use hvDFL1sd_CDNS_52468879185990  hvDFL1sd_CDNS_52468879185990_1
timestamp 1707688321
transform 1 0 1656 0 1 0
box -26 -26 79 2026
<< labels >>
flabel comment s -28 981 -28 981 0 FreeSans 300 0 0 0 S
flabel comment s 828 981 828 981 0 FreeSans 300 0 0 0 D
flabel comment s 1684 981 1684 981 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 97520888
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 97519434
<< end >>
