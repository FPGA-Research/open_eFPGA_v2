magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -76 -26 532 626
<< mvnmos >>
rect 0 0 200 600
rect 256 0 456 600
<< mvndiff >>
rect -50 0 0 600
rect 456 0 506 600
<< poly >>
rect 0 600 200 626
rect 0 -26 200 0
rect 256 600 456 626
rect 256 -26 456 0
<< metal1 >>
rect -51 -16 -5 546
rect 205 -16 251 546
rect 461 -16 507 546
use hvDFM1sd2_CDNS_52468879185154  hvDFM1sd2_CDNS_52468879185154_0
timestamp 1707688321
transform 1 0 200 0 1 0
box -26 -26 82 626
use hvDFM1sd_CDNS_52468879185149  hvDFM1sd_CDNS_52468879185149_0
timestamp 1707688321
transform -1 0 0 0 1 0
box -26 -26 79 626
use hvDFM1sd_CDNS_52468879185149  hvDFM1sd_CDNS_52468879185149_1
timestamp 1707688321
transform 1 0 456 0 1 0
box -26 -26 79 626
<< labels >>
flabel comment s -28 265 -28 265 0 FreeSans 300 0 0 0 S
flabel comment s 228 265 228 265 0 FreeSans 300 0 0 0 D
flabel comment s 484 265 484 265 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 86617622
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86616232
<< end >>
