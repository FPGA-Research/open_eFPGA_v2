magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -68 -26 374 162
<< ndiff >>
rect -42 119 0 136
rect -42 85 -34 119
rect -42 51 0 85
rect -42 17 -34 51
rect -42 0 0 17
rect 306 119 348 136
rect 340 85 348 119
rect 306 51 348 85
rect 340 17 348 51
rect 306 0 348 17
<< ndiffc >>
rect -34 85 0 119
rect -34 17 0 51
rect 306 85 340 119
rect 306 17 340 51
<< ndiffres >>
rect 0 0 306 136
<< locali >>
rect -34 119 0 135
rect -34 51 0 85
rect -34 1 0 17
rect 306 119 340 135
rect 306 51 340 85
rect 306 1 340 17
use DFL1_CDNS_524688791851252  DFL1_CDNS_524688791851252_0
timestamp 1707688321
transform -1 0 8 0 1 5
box 0 0 1 1
use DFL1_CDNS_524688791851252  DFL1_CDNS_524688791851252_1
timestamp 1707688321
transform 1 0 298 0 1 5
box 0 0 1 1
<< properties >>
string GDS_END 86903432
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86902926
<< end >>
