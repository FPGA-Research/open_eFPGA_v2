magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< metal2 >>
rect 0 6145 536 6154
rect 0 0 536 9
<< via2 >>
rect 0 9 536 6145
<< metal3 >>
rect -5 6145 541 6150
rect -5 9 0 6145
rect 536 9 541 6145
rect -5 4 541 9
<< properties >>
string GDS_END 93487290
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 93452662
<< end >>
