magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< metal3 >>
rect 0 470 944 476
rect 0 0 944 6
<< via3 >>
rect 0 6 944 470
<< metal4 >>
rect -1 470 945 471
rect -1 6 0 470
rect 944 6 945 470
rect -1 5 945 6
<< properties >>
string GDS_END 87517180
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87512440
<< end >>
