magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< poly >>
rect -50 50 0 66
rect -50 16 -34 50
rect -50 0 0 16
rect 11896 -598 11946 -582
rect 11930 -632 11946 -598
rect 11896 -648 11946 -632
<< polycont >>
rect -34 16 0 50
rect 11896 -632 11930 -598
<< npolyres >>
rect 0 0 11946 66
rect 11880 -96 11946 0
rect -50 -162 11946 -96
rect -50 -258 16 -162
rect -50 -324 11946 -258
rect 11880 -420 11946 -324
rect -50 -486 11946 -420
rect -50 -582 16 -486
rect -50 -648 11896 -582
<< locali >>
rect -34 50 0 66
rect -34 0 0 16
rect 11896 -598 11930 -582
rect 11896 -648 11930 -632
use PYL1_CDNS_5595914180839  PYL1_CDNS_5595914180839_0
timestamp 1707688321
transform 1 0 -50 0 1 0
box 0 0 1 1
use PYL1_CDNS_5595914180839  PYL1_CDNS_5595914180839_1
timestamp 1707688321
transform 1 0 11880 0 1 -648
box 0 0 1 1
<< properties >>
string GDS_END 42935772
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 42934200
<< end >>
