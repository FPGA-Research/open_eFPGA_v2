magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -38 261 1602 582
<< pwell >>
rect 5 21 1558 203
rect 29 -17 63 21
<< locali >>
rect 1154 339 1188 493
rect 1322 339 1356 493
rect 1490 339 1547 493
rect 755 289 1547 339
rect 18 211 356 285
rect 390 211 721 285
rect 755 211 1188 255
rect 1222 177 1259 289
rect 1293 211 1547 255
rect 1222 129 1456 177
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 18 379 89 493
rect 123 413 157 527
rect 191 379 257 493
rect 291 413 325 527
rect 359 441 777 493
rect 359 379 425 441
rect 18 319 425 379
rect 459 353 493 407
rect 527 387 593 441
rect 816 407 1120 493
rect 627 373 1120 407
rect 627 353 721 373
rect 459 319 721 353
rect 1222 378 1288 527
rect 1390 378 1456 527
rect 18 143 1188 177
rect 18 51 89 143
rect 123 17 157 109
rect 191 51 257 143
rect 291 17 325 109
rect 359 51 425 143
rect 459 17 493 109
rect 527 51 593 143
rect 627 17 661 109
rect 695 51 761 143
rect 799 17 928 109
rect 962 79 996 143
rect 1030 17 1120 109
rect 1154 95 1188 143
rect 1490 95 1547 177
rect 1154 51 1547 95
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
<< metal1 >>
rect 0 561 1564 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 0 496 1564 527
rect 0 17 1564 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
rect 0 -48 1564 -17
<< labels >>
rlabel locali s 18 211 356 285 6 A1
port 1 nsew signal input
rlabel locali s 390 211 721 285 6 A2
port 2 nsew signal input
rlabel locali s 755 211 1188 255 6 A3
port 3 nsew signal input
rlabel locali s 1293 211 1547 255 6 B1
port 4 nsew signal input
rlabel metal1 s 0 -48 1564 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 5 21 1558 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 1602 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 1564 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1222 129 1456 177 6 Y
port 9 nsew signal output
rlabel locali s 1222 177 1259 289 6 Y
port 9 nsew signal output
rlabel locali s 755 289 1547 339 6 Y
port 9 nsew signal output
rlabel locali s 1490 339 1547 493 6 Y
port 9 nsew signal output
rlabel locali s 1322 339 1356 493 6 Y
port 9 nsew signal output
rlabel locali s 1154 339 1188 493 6 Y
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1564 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1448880
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1434396
<< end >>
