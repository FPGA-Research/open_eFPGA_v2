magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -79 -26 879 226
<< mvnmos >>
rect 0 0 800 200
<< mvndiff >>
rect -53 182 0 200
rect -53 148 -45 182
rect -11 148 0 182
rect -53 114 0 148
rect -53 80 -45 114
rect -11 80 0 114
rect -53 46 0 80
rect -53 12 -45 46
rect -11 12 0 46
rect -53 0 0 12
rect 800 182 853 200
rect 800 148 811 182
rect 845 148 853 182
rect 800 114 853 148
rect 800 80 811 114
rect 845 80 853 114
rect 800 46 853 80
rect 800 12 811 46
rect 845 12 853 46
rect 800 0 853 12
<< mvndiffc >>
rect -45 148 -11 182
rect -45 80 -11 114
rect -45 12 -11 46
rect 811 148 845 182
rect 811 80 845 114
rect 811 12 845 46
<< poly >>
rect 0 200 800 232
rect 0 -32 800 0
<< locali >>
rect -45 182 -11 198
rect -45 114 -11 148
rect -45 46 -11 80
rect -45 -4 -11 12
rect 811 182 845 198
rect 811 114 845 148
rect 811 46 845 80
rect 811 -4 845 12
use DFL1sd_CDNS_5246887918538  DFL1sd_CDNS_5246887918538_0
timestamp 1707688321
transform -1 0 0 0 1 0
box 0 0 1 1
use DFL1sd_CDNS_5246887918538  DFL1sd_CDNS_5246887918538_1
timestamp 1707688321
transform 1 0 800 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 97 -28 97 0 FreeSans 300 0 0 0 S
flabel comment s 828 97 828 97 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 89251798
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 89250912
<< end >>
