magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< dnwell >>
rect 2376 6058 7066 11061
<< nwell >>
rect 0 27767 2436 27937
rect 0 25624 170 27767
rect 2266 11146 2436 27767
rect 2266 10976 7146 11146
rect 2266 6338 2656 10976
rect 6786 6338 7146 10976
rect 2266 5978 7146 6338
rect 5742 5791 7146 5978
rect 3274 170 3444 966
rect 675 144 3444 170
rect 675 -385 3707 144
rect 675 -561 845 -385
rect 1613 -467 3707 -385
rect 1613 -561 1783 -467
rect 675 -731 1783 -561
<< pwell >>
rect 230 27477 2206 27707
rect 230 23830 318 27477
rect 2118 23830 2206 27477
rect 230 23582 2206 23830
rect 230 19935 318 23582
rect 2118 22359 2206 23582
rect 1348 19935 2206 22359
rect 230 19687 2206 19935
rect 230 16040 318 19687
rect 2118 16040 2206 19687
rect 230 15792 2206 16040
rect 230 12145 318 15792
rect 2118 12145 2206 15792
rect 230 11897 2206 12145
rect 230 8250 318 11897
rect 2118 8250 2206 11897
rect 230 8002 2206 8250
rect 230 6816 318 8002
rect 205 4355 318 6816
rect 1978 5601 2206 8002
rect 2716 10828 6726 10916
rect 2716 6486 2804 10828
rect 4677 6486 4765 10828
rect 6638 6486 6726 10828
rect 2716 6398 6726 6486
rect 1978 5371 3214 5601
rect 205 4351 1970 4355
rect 230 4101 1970 4351
rect 230 460 318 4101
rect 1852 4066 1970 4101
rect 3126 460 3214 5371
rect 3504 5514 5682 5602
rect 3504 4362 3592 5514
rect 5594 4362 5682 5514
rect 3504 4274 5682 4362
rect 230 230 3214 460
rect 2122 -615 3524 -527
rect 2122 -968 2210 -615
rect 3436 -968 3524 -615
rect 2122 -1056 3524 -968
<< mvndiff >>
rect 366 27563 432 27571
rect 366 27529 382 27563
rect 416 27529 432 27563
rect 366 27503 432 27529
rect 492 27563 558 27571
rect 492 27529 508 27563
rect 542 27529 558 27563
rect 492 27503 558 27529
rect 618 27563 684 27571
rect 618 27529 634 27563
rect 668 27529 684 27563
rect 618 27503 684 27529
rect 744 27563 810 27571
rect 744 27529 760 27563
rect 794 27529 810 27563
rect 744 27503 810 27529
rect 870 27563 936 27571
rect 870 27529 886 27563
rect 920 27529 936 27563
rect 870 27503 936 27529
rect 996 27563 1062 27571
rect 996 27529 1012 27563
rect 1046 27529 1062 27563
rect 996 27503 1062 27529
rect 1122 27563 1188 27571
rect 1122 27529 1138 27563
rect 1172 27529 1188 27563
rect 1122 27503 1188 27529
rect 1248 27563 1314 27571
rect 1248 27529 1264 27563
rect 1298 27529 1314 27563
rect 1248 27503 1314 27529
rect 1374 27563 1440 27571
rect 1374 27529 1390 27563
rect 1424 27529 1440 27563
rect 1374 27503 1440 27529
rect 1500 27563 1566 27571
rect 1500 27529 1516 27563
rect 1550 27529 1566 27563
rect 1500 27503 1566 27529
rect 1626 27563 1692 27571
rect 1626 27529 1642 27563
rect 1676 27529 1692 27563
rect 1626 27503 1692 27529
rect 1752 27563 1818 27571
rect 1752 27529 1768 27563
rect 1802 27529 1818 27563
rect 1752 27503 1818 27529
rect 1878 27563 1944 27571
rect 1878 27529 1894 27563
rect 1928 27529 1944 27563
rect 1878 27503 1944 27529
rect 2004 27563 2070 27571
rect 2004 27529 2020 27563
rect 2054 27529 2070 27563
rect 2004 27503 2070 27529
rect 366 23778 432 23804
rect 366 23744 382 23778
rect 416 23744 432 23778
rect 366 23736 432 23744
rect 492 23778 558 23804
rect 492 23744 508 23778
rect 542 23744 558 23778
rect 492 23736 558 23744
rect 618 23778 684 23804
rect 618 23744 634 23778
rect 668 23744 684 23778
rect 618 23736 684 23744
rect 744 23778 810 23804
rect 744 23744 760 23778
rect 794 23744 810 23778
rect 744 23736 810 23744
rect 870 23778 936 23804
rect 870 23744 886 23778
rect 920 23744 936 23778
rect 870 23736 936 23744
rect 996 23778 1062 23804
rect 996 23744 1012 23778
rect 1046 23744 1062 23778
rect 996 23736 1062 23744
rect 1122 23778 1188 23804
rect 1122 23744 1138 23778
rect 1172 23744 1188 23778
rect 1122 23736 1188 23744
rect 1248 23778 1314 23804
rect 1248 23744 1264 23778
rect 1298 23744 1314 23778
rect 1248 23736 1314 23744
rect 1374 23778 1440 23804
rect 1374 23744 1390 23778
rect 1424 23744 1440 23778
rect 1374 23736 1440 23744
rect 1500 23778 1566 23804
rect 1500 23744 1516 23778
rect 1550 23744 1566 23778
rect 1500 23736 1566 23744
rect 1626 23778 1692 23804
rect 1626 23744 1642 23778
rect 1676 23744 1692 23778
rect 1626 23736 1692 23744
rect 1752 23778 1818 23804
rect 1752 23744 1768 23778
rect 1802 23744 1818 23778
rect 1752 23736 1818 23744
rect 1878 23778 1944 23804
rect 1878 23744 1894 23778
rect 1928 23744 1944 23778
rect 1878 23736 1944 23744
rect 2004 23778 2070 23804
rect 2004 23744 2020 23778
rect 2054 23744 2070 23778
rect 2004 23736 2070 23744
rect 366 23668 432 23676
rect 366 23634 382 23668
rect 416 23634 432 23668
rect 366 23608 432 23634
rect 492 23668 558 23676
rect 492 23634 508 23668
rect 542 23634 558 23668
rect 492 23608 558 23634
rect 618 23668 684 23676
rect 618 23634 634 23668
rect 668 23634 684 23668
rect 618 23608 684 23634
rect 744 23668 810 23676
rect 744 23634 760 23668
rect 794 23634 810 23668
rect 744 23608 810 23634
rect 870 23668 936 23676
rect 870 23634 886 23668
rect 920 23634 936 23668
rect 870 23608 936 23634
rect 996 23668 1062 23676
rect 996 23634 1012 23668
rect 1046 23634 1062 23668
rect 996 23608 1062 23634
rect 1122 23668 1188 23676
rect 1122 23634 1138 23668
rect 1172 23634 1188 23668
rect 1122 23608 1188 23634
rect 1248 23668 1314 23676
rect 1248 23634 1264 23668
rect 1298 23634 1314 23668
rect 1248 23608 1314 23634
rect 1374 23668 1440 23676
rect 1374 23634 1390 23668
rect 1424 23634 1440 23668
rect 1374 23608 1440 23634
rect 1500 23668 1566 23676
rect 1500 23634 1516 23668
rect 1550 23634 1566 23668
rect 1500 23608 1566 23634
rect 1626 23668 1692 23676
rect 1626 23634 1642 23668
rect 1676 23634 1692 23668
rect 1626 23608 1692 23634
rect 1752 23668 1818 23676
rect 1752 23634 1768 23668
rect 1802 23634 1818 23668
rect 1752 23608 1818 23634
rect 1878 23668 1944 23676
rect 1878 23634 1894 23668
rect 1928 23634 1944 23668
rect 1878 23608 1944 23634
rect 2004 23668 2070 23676
rect 2004 23634 2020 23668
rect 2054 23634 2070 23668
rect 2004 23608 2070 23634
rect 1374 22307 1440 22333
rect 1374 22273 1390 22307
rect 1424 22273 1440 22307
rect 366 19883 432 19909
rect 366 19849 382 19883
rect 416 19849 432 19883
rect 366 19841 432 19849
rect 492 19883 558 19909
rect 492 19849 508 19883
rect 542 19849 558 19883
rect 492 19841 558 19849
rect 618 19883 684 19909
rect 618 19849 634 19883
rect 668 19849 684 19883
rect 618 19841 684 19849
rect 744 19883 810 19909
rect 744 19849 760 19883
rect 794 19849 810 19883
rect 744 19841 810 19849
rect 870 19883 936 19909
rect 870 19849 886 19883
rect 920 19849 936 19883
rect 870 19841 936 19849
rect 996 19883 1062 19909
rect 996 19849 1012 19883
rect 1046 19849 1062 19883
rect 996 19841 1062 19849
rect 1122 19883 1188 19909
rect 1122 19849 1138 19883
rect 1172 19849 1188 19883
rect 1122 19841 1188 19849
rect 1248 19883 1314 19909
rect 1248 19849 1264 19883
rect 1298 19849 1314 19883
rect 1248 19841 1314 19849
rect 1374 19841 1440 22273
rect 1626 22307 1692 22333
rect 1626 22273 1642 22307
rect 1676 22273 1692 22307
rect 1500 19883 1566 19909
rect 1500 19849 1516 19883
rect 1550 19849 1566 19883
rect 1500 19841 1566 19849
rect 1626 19841 1692 22273
rect 1878 22307 1944 22333
rect 1878 22273 1894 22307
rect 1928 22273 1944 22307
rect 1752 19883 1818 19909
rect 1752 19849 1768 19883
rect 1802 19849 1818 19883
rect 1752 19841 1818 19849
rect 1878 19841 1944 22273
rect 2004 19883 2070 19909
rect 2004 19849 2020 19883
rect 2054 19849 2070 19883
rect 2004 19841 2070 19849
rect 366 19773 432 19781
rect 366 19739 382 19773
rect 416 19739 432 19773
rect 366 19713 432 19739
rect 492 19773 558 19781
rect 492 19739 508 19773
rect 542 19739 558 19773
rect 492 19713 558 19739
rect 618 19773 684 19781
rect 618 19739 634 19773
rect 668 19739 684 19773
rect 618 19713 684 19739
rect 744 19773 810 19781
rect 744 19739 760 19773
rect 794 19739 810 19773
rect 744 19713 810 19739
rect 870 19773 936 19781
rect 870 19739 886 19773
rect 920 19739 936 19773
rect 870 19713 936 19739
rect 996 19773 1062 19781
rect 996 19739 1012 19773
rect 1046 19739 1062 19773
rect 996 19713 1062 19739
rect 1122 19773 1188 19781
rect 1122 19739 1138 19773
rect 1172 19739 1188 19773
rect 1122 19713 1188 19739
rect 1248 19773 1314 19781
rect 1248 19739 1264 19773
rect 1298 19739 1314 19773
rect 1248 19713 1314 19739
rect 1374 19773 1440 19781
rect 1374 19739 1390 19773
rect 1424 19739 1440 19773
rect 1374 19713 1440 19739
rect 1500 19773 1566 19781
rect 1500 19739 1516 19773
rect 1550 19739 1566 19773
rect 1500 19713 1566 19739
rect 1626 19773 1692 19781
rect 1626 19739 1642 19773
rect 1676 19739 1692 19773
rect 1626 19713 1692 19739
rect 1752 19773 1818 19781
rect 1752 19739 1768 19773
rect 1802 19739 1818 19773
rect 1752 19713 1818 19739
rect 1878 19773 1944 19781
rect 1878 19739 1894 19773
rect 1928 19739 1944 19773
rect 1878 19713 1944 19739
rect 2004 19773 2070 19781
rect 2004 19739 2020 19773
rect 2054 19739 2070 19773
rect 2004 19713 2070 19739
rect 366 15988 432 16014
rect 366 15954 382 15988
rect 416 15954 432 15988
rect 366 15946 432 15954
rect 492 15988 558 16014
rect 492 15954 508 15988
rect 542 15954 558 15988
rect 492 15946 558 15954
rect 618 15988 684 16014
rect 618 15954 634 15988
rect 668 15954 684 15988
rect 618 15946 684 15954
rect 744 15988 810 16014
rect 744 15954 760 15988
rect 794 15954 810 15988
rect 744 15946 810 15954
rect 870 15988 936 16014
rect 870 15954 886 15988
rect 920 15954 936 15988
rect 870 15946 936 15954
rect 996 15988 1062 16014
rect 996 15954 1012 15988
rect 1046 15954 1062 15988
rect 996 15946 1062 15954
rect 1122 15988 1188 16014
rect 1122 15954 1138 15988
rect 1172 15954 1188 15988
rect 1122 15946 1188 15954
rect 1248 15988 1314 16014
rect 1248 15954 1264 15988
rect 1298 15954 1314 15988
rect 1248 15946 1314 15954
rect 1374 15988 1440 16014
rect 1374 15954 1390 15988
rect 1424 15954 1440 15988
rect 1374 15946 1440 15954
rect 1500 15988 1566 16014
rect 1500 15954 1516 15988
rect 1550 15954 1566 15988
rect 1500 15946 1566 15954
rect 1626 15988 1692 16014
rect 1626 15954 1642 15988
rect 1676 15954 1692 15988
rect 1626 15946 1692 15954
rect 1752 15988 1818 16014
rect 1752 15954 1768 15988
rect 1802 15954 1818 15988
rect 1752 15946 1818 15954
rect 1878 15988 1944 16014
rect 1878 15954 1894 15988
rect 1928 15954 1944 15988
rect 1878 15946 1944 15954
rect 2004 15988 2070 16014
rect 2004 15954 2020 15988
rect 2054 15954 2070 15988
rect 2004 15946 2070 15954
rect 366 15878 432 15886
rect 366 15844 382 15878
rect 416 15844 432 15878
rect 366 15818 432 15844
rect 492 15878 558 15886
rect 492 15844 508 15878
rect 542 15844 558 15878
rect 492 15818 558 15844
rect 618 15878 684 15886
rect 618 15844 634 15878
rect 668 15844 684 15878
rect 618 15818 684 15844
rect 744 15878 810 15886
rect 744 15844 760 15878
rect 794 15844 810 15878
rect 744 15818 810 15844
rect 870 15878 936 15886
rect 870 15844 886 15878
rect 920 15844 936 15878
rect 870 15818 936 15844
rect 996 15878 1062 15886
rect 996 15844 1012 15878
rect 1046 15844 1062 15878
rect 996 15818 1062 15844
rect 1122 15878 1188 15886
rect 1122 15844 1138 15878
rect 1172 15844 1188 15878
rect 1122 15818 1188 15844
rect 1248 15878 1314 15886
rect 1248 15844 1264 15878
rect 1298 15844 1314 15878
rect 1248 15818 1314 15844
rect 1374 15878 1440 15886
rect 1374 15844 1390 15878
rect 1424 15844 1440 15878
rect 1374 15818 1440 15844
rect 1500 15878 1566 15886
rect 1500 15844 1516 15878
rect 1550 15844 1566 15878
rect 1500 15818 1566 15844
rect 1626 15878 1692 15886
rect 1626 15844 1642 15878
rect 1676 15844 1692 15878
rect 1626 15818 1692 15844
rect 1752 15878 1818 15886
rect 1752 15844 1768 15878
rect 1802 15844 1818 15878
rect 1752 15818 1818 15844
rect 1878 15878 1944 15886
rect 1878 15844 1894 15878
rect 1928 15844 1944 15878
rect 1878 15818 1944 15844
rect 2004 15878 2070 15886
rect 2004 15844 2020 15878
rect 2054 15844 2070 15878
rect 2004 15818 2070 15844
rect 366 12093 432 12119
rect 366 12059 382 12093
rect 416 12059 432 12093
rect 366 12051 432 12059
rect 492 12093 558 12119
rect 492 12059 508 12093
rect 542 12059 558 12093
rect 492 12051 558 12059
rect 618 12093 684 12119
rect 618 12059 634 12093
rect 668 12059 684 12093
rect 618 12051 684 12059
rect 744 12093 810 12119
rect 744 12059 760 12093
rect 794 12059 810 12093
rect 744 12051 810 12059
rect 870 12093 936 12119
rect 870 12059 886 12093
rect 920 12059 936 12093
rect 870 12051 936 12059
rect 996 12093 1062 12119
rect 996 12059 1012 12093
rect 1046 12059 1062 12093
rect 996 12051 1062 12059
rect 1122 12093 1188 12119
rect 1122 12059 1138 12093
rect 1172 12059 1188 12093
rect 1122 12051 1188 12059
rect 1248 12093 1314 12119
rect 1248 12059 1264 12093
rect 1298 12059 1314 12093
rect 1248 12051 1314 12059
rect 1374 12093 1440 12119
rect 1374 12059 1390 12093
rect 1424 12059 1440 12093
rect 1374 12051 1440 12059
rect 1500 12093 1566 12119
rect 1500 12059 1516 12093
rect 1550 12059 1566 12093
rect 1500 12051 1566 12059
rect 1626 12093 1692 12119
rect 1626 12059 1642 12093
rect 1676 12059 1692 12093
rect 1626 12051 1692 12059
rect 1752 12093 1818 12119
rect 1752 12059 1768 12093
rect 1802 12059 1818 12093
rect 1752 12051 1818 12059
rect 1878 12093 1944 12119
rect 1878 12059 1894 12093
rect 1928 12059 1944 12093
rect 1878 12051 1944 12059
rect 2004 12093 2070 12119
rect 2004 12059 2020 12093
rect 2054 12059 2070 12093
rect 2004 12051 2070 12059
rect 366 11983 432 11991
rect 366 11949 382 11983
rect 416 11949 432 11983
rect 366 11923 432 11949
rect 492 11983 558 11991
rect 492 11949 508 11983
rect 542 11949 558 11983
rect 492 11923 558 11949
rect 618 11983 684 11991
rect 618 11949 634 11983
rect 668 11949 684 11983
rect 618 11923 684 11949
rect 744 11983 810 11991
rect 744 11949 760 11983
rect 794 11949 810 11983
rect 744 11923 810 11949
rect 870 11983 936 11991
rect 870 11949 886 11983
rect 920 11949 936 11983
rect 870 11923 936 11949
rect 996 11983 1062 11991
rect 996 11949 1012 11983
rect 1046 11949 1062 11983
rect 996 11923 1062 11949
rect 1122 11983 1188 11991
rect 1122 11949 1138 11983
rect 1172 11949 1188 11983
rect 1122 11923 1188 11949
rect 1248 11983 1314 11991
rect 1248 11949 1264 11983
rect 1298 11949 1314 11983
rect 1248 11923 1314 11949
rect 1374 11983 1440 11991
rect 1374 11949 1390 11983
rect 1424 11949 1440 11983
rect 1374 11923 1440 11949
rect 1500 11983 1566 11991
rect 1500 11949 1516 11983
rect 1550 11949 1566 11983
rect 1500 11923 1566 11949
rect 1626 11983 1692 11991
rect 1626 11949 1642 11983
rect 1676 11949 1692 11983
rect 1626 11923 1692 11949
rect 1752 11983 1818 11991
rect 1752 11949 1768 11983
rect 1802 11949 1818 11983
rect 1752 11923 1818 11949
rect 1878 11983 1944 11991
rect 1878 11949 1894 11983
rect 1928 11949 1944 11983
rect 1878 11923 1944 11949
rect 2004 11983 2070 11991
rect 2004 11949 2020 11983
rect 2054 11949 2070 11983
rect 2004 11923 2070 11949
rect 366 8198 432 8224
rect 366 8164 382 8198
rect 416 8164 432 8198
rect 366 8156 432 8164
rect 492 8198 558 8224
rect 492 8164 508 8198
rect 542 8164 558 8198
rect 492 8156 558 8164
rect 618 8198 684 8224
rect 618 8164 634 8198
rect 668 8164 684 8198
rect 618 8156 684 8164
rect 744 8198 810 8224
rect 744 8164 760 8198
rect 794 8164 810 8198
rect 744 8156 810 8164
rect 870 8198 936 8224
rect 870 8164 886 8198
rect 920 8164 936 8198
rect 870 8156 936 8164
rect 996 8198 1062 8224
rect 996 8164 1012 8198
rect 1046 8164 1062 8198
rect 996 8156 1062 8164
rect 1122 8198 1188 8224
rect 1122 8164 1138 8198
rect 1172 8164 1188 8198
rect 1122 8156 1188 8164
rect 1248 8198 1314 8224
rect 1248 8164 1264 8198
rect 1298 8164 1314 8198
rect 1248 8156 1314 8164
rect 1374 8198 1440 8224
rect 1374 8164 1390 8198
rect 1424 8164 1440 8198
rect 1374 8156 1440 8164
rect 1500 8198 1566 8224
rect 1500 8164 1516 8198
rect 1550 8164 1566 8198
rect 1500 8156 1566 8164
rect 1626 8198 1692 8224
rect 1626 8164 1642 8198
rect 1676 8164 1692 8198
rect 1626 8156 1692 8164
rect 1752 8198 1818 8224
rect 1752 8164 1768 8198
rect 1802 8164 1818 8198
rect 1752 8156 1818 8164
rect 1878 8198 1944 8224
rect 1878 8164 1894 8198
rect 1928 8164 1944 8198
rect 1878 8156 1944 8164
rect 2004 8198 2070 8224
rect 2004 8164 2020 8198
rect 2054 8164 2070 8198
rect 366 8088 432 8096
rect 366 8054 382 8088
rect 416 8054 432 8088
rect 366 8028 432 8054
rect 492 8088 558 8096
rect 492 8054 508 8088
rect 542 8054 558 8088
rect 492 8028 558 8054
rect 618 8088 684 8096
rect 618 8054 634 8088
rect 668 8054 684 8088
rect 618 8028 684 8054
rect 744 8088 810 8096
rect 744 8054 760 8088
rect 794 8054 810 8088
rect 744 8028 810 8054
rect 870 8088 936 8096
rect 870 8054 886 8088
rect 920 8054 936 8088
rect 870 8028 936 8054
rect 996 8088 1062 8096
rect 996 8054 1012 8088
rect 1046 8054 1062 8088
rect 996 8028 1062 8054
rect 1122 8088 1188 8096
rect 1122 8054 1138 8088
rect 1172 8054 1188 8088
rect 1122 8028 1188 8054
rect 1248 8088 1314 8096
rect 1248 8054 1264 8088
rect 1298 8054 1314 8088
rect 1248 8028 1314 8054
rect 1374 8088 1440 8096
rect 1374 8054 1390 8088
rect 1424 8054 1440 8088
rect 1374 8028 1440 8054
rect 1500 8088 1566 8096
rect 1500 8054 1516 8088
rect 1550 8054 1566 8088
rect 1500 8028 1566 8054
rect 1626 8088 1692 8096
rect 1626 8054 1642 8088
rect 1676 8054 1692 8088
rect 1626 8028 1692 8054
rect 1752 8088 1818 8096
rect 1752 8054 1768 8088
rect 1802 8054 1818 8088
rect 1752 8028 1818 8054
rect 1878 8088 1944 8096
rect 1878 8054 1894 8088
rect 1928 8054 1944 8088
rect 1878 8028 1944 8054
rect 2004 5525 2070 8164
rect 2004 5457 2070 5465
rect 2004 5423 2020 5457
rect 2054 5423 2070 5457
rect 2004 5397 2070 5423
rect 2130 5457 2196 5465
rect 2130 5423 2146 5457
rect 2180 5423 2196 5457
rect 2130 5397 2196 5423
rect 2256 5457 2322 5465
rect 2256 5423 2272 5457
rect 2306 5423 2322 5457
rect 2256 5397 2322 5423
rect 2382 5457 2448 5465
rect 2382 5423 2398 5457
rect 2432 5423 2448 5457
rect 2382 5397 2448 5423
rect 2508 5457 2574 5465
rect 2508 5423 2524 5457
rect 2558 5423 2574 5457
rect 2508 5397 2574 5423
rect 2634 5457 2700 5465
rect 2634 5423 2650 5457
rect 2684 5423 2700 5457
rect 2634 5397 2700 5423
rect 2760 5457 2826 5465
rect 2760 5423 2776 5457
rect 2810 5423 2826 5457
rect 2760 5397 2826 5423
rect 2886 5457 2952 5465
rect 2886 5423 2902 5457
rect 2936 5423 2952 5457
rect 2886 5397 2952 5423
rect 3012 5457 3078 5465
rect 3012 5423 3028 5457
rect 3062 5423 3078 5457
rect 3012 5397 3078 5423
rect 366 4303 432 4329
rect 366 4269 382 4303
rect 416 4269 432 4303
rect 366 4261 432 4269
rect 492 4303 558 4329
rect 492 4269 508 4303
rect 542 4269 558 4303
rect 492 4261 558 4269
rect 618 4303 684 4329
rect 618 4269 634 4303
rect 668 4269 684 4303
rect 618 4261 684 4269
rect 744 4303 810 4329
rect 744 4269 760 4303
rect 794 4269 810 4303
rect 744 4261 810 4269
rect 870 4303 936 4329
rect 870 4269 886 4303
rect 920 4269 936 4303
rect 870 4261 936 4269
rect 996 4303 1062 4329
rect 996 4269 1012 4303
rect 1046 4269 1062 4303
rect 996 4261 1062 4269
rect 1122 4303 1188 4329
rect 1122 4269 1138 4303
rect 1172 4269 1188 4303
rect 1122 4261 1188 4269
rect 1248 4303 1314 4329
rect 1248 4269 1264 4303
rect 1298 4269 1314 4303
rect 1248 4261 1314 4269
rect 1374 4303 1440 4329
rect 1374 4269 1390 4303
rect 1424 4269 1440 4303
rect 1374 4261 1440 4269
rect 1500 4303 1566 4329
rect 1500 4269 1516 4303
rect 1550 4269 1566 4303
rect 1500 4261 1566 4269
rect 1626 4303 1692 4329
rect 1626 4269 1642 4303
rect 1676 4269 1692 4303
rect 1626 4261 1692 4269
rect 1752 4303 1818 4329
rect 1752 4269 1768 4303
rect 1802 4269 1818 4303
rect 1752 4261 1818 4269
rect 1878 4303 1944 4329
rect 1878 4269 1894 4303
rect 1928 4269 1944 4303
rect 1878 4261 1944 4269
rect 366 4193 432 4201
rect 366 4159 382 4193
rect 416 4159 432 4193
rect 366 4127 432 4159
rect 492 4193 558 4201
rect 492 4159 508 4193
rect 542 4159 558 4193
rect 492 4127 558 4159
rect 618 4193 684 4201
rect 618 4159 634 4193
rect 668 4159 684 4193
rect 618 4127 684 4159
rect 744 4193 810 4201
rect 744 4159 760 4193
rect 794 4159 810 4193
rect 744 4127 810 4159
rect 870 4193 936 4201
rect 870 4159 886 4193
rect 920 4159 936 4193
rect 870 4127 936 4159
rect 996 4193 1062 4201
rect 996 4159 1012 4193
rect 1046 4159 1062 4193
rect 996 4127 1062 4159
rect 1122 4193 1188 4201
rect 1122 4159 1138 4193
rect 1172 4159 1188 4193
rect 1122 4127 1188 4159
rect 1248 4193 1314 4201
rect 1248 4159 1264 4193
rect 1298 4159 1314 4193
rect 1248 4127 1314 4159
rect 1374 4193 1440 4201
rect 1374 4159 1390 4193
rect 1424 4159 1440 4193
rect 1374 4127 1440 4159
rect 1500 4193 1566 4201
rect 1500 4159 1516 4193
rect 1550 4159 1566 4193
rect 1500 4127 1566 4159
rect 1626 4193 1692 4201
rect 1626 4159 1642 4193
rect 1676 4159 1692 4193
rect 1626 4127 1692 4159
rect 1752 4193 1818 4201
rect 1752 4159 1768 4193
rect 1802 4159 1818 4193
rect 1752 4127 1818 4159
rect 1878 4193 1944 4201
rect 1878 4159 1894 4193
rect 1928 4159 1944 4193
rect 1878 4092 1944 4159
rect 366 408 432 434
rect 366 374 382 408
rect 416 374 432 408
rect 366 366 432 374
rect 492 408 558 434
rect 492 374 508 408
rect 542 374 558 408
rect 492 366 558 374
rect 618 408 684 434
rect 618 374 634 408
rect 668 374 684 408
rect 618 366 684 374
rect 744 408 810 434
rect 744 374 760 408
rect 794 374 810 408
rect 744 366 810 374
rect 870 408 936 434
rect 870 374 886 408
rect 920 374 936 408
rect 870 366 936 374
rect 996 408 1062 434
rect 996 374 1012 408
rect 1046 374 1062 408
rect 996 366 1062 374
rect 1122 408 1188 434
rect 1122 374 1138 408
rect 1172 374 1188 408
rect 1122 366 1188 374
rect 1248 408 1314 434
rect 1248 374 1264 408
rect 1298 374 1314 408
rect 1248 366 1314 374
rect 1374 408 1440 434
rect 1374 374 1390 408
rect 1424 374 1440 408
rect 1374 366 1440 374
rect 1500 408 1566 434
rect 1500 374 1516 408
rect 1550 374 1566 408
rect 1500 366 1566 374
rect 1626 408 1692 434
rect 1626 374 1642 408
rect 1676 374 1692 408
rect 1626 366 1692 374
rect 1752 408 1818 434
rect 1752 374 1768 408
rect 1802 374 1818 408
rect 1752 366 1818 374
rect 1878 408 1944 434
rect 1878 374 1894 408
rect 1928 374 1944 408
rect 1878 366 1944 374
rect 2004 408 2070 434
rect 2004 374 2020 408
rect 2054 374 2070 408
rect 2004 366 2070 374
rect 2130 408 2196 434
rect 2130 374 2146 408
rect 2180 374 2196 408
rect 2130 366 2196 374
rect 2256 408 2322 434
rect 2256 374 2272 408
rect 2306 374 2322 408
rect 2256 366 2322 374
rect 2382 408 2448 434
rect 2382 374 2398 408
rect 2432 374 2448 408
rect 2382 366 2448 374
rect 2508 408 2574 434
rect 2508 374 2524 408
rect 2558 374 2574 408
rect 2508 366 2574 374
rect 2634 408 2700 434
rect 2634 374 2650 408
rect 2684 374 2700 408
rect 2634 366 2700 374
rect 2760 408 2826 434
rect 2760 374 2776 408
rect 2810 374 2826 408
rect 2760 366 2826 374
rect 2886 408 2952 434
rect 2886 374 2902 408
rect 2936 374 2952 408
rect 2886 366 2952 374
rect 3012 408 3078 434
rect 3012 374 3028 408
rect 3062 374 3078 408
rect 3012 366 3078 374
<< mvndiffc >>
rect 382 27529 416 27563
rect 508 27529 542 27563
rect 634 27529 668 27563
rect 760 27529 794 27563
rect 886 27529 920 27563
rect 1012 27529 1046 27563
rect 1138 27529 1172 27563
rect 1264 27529 1298 27563
rect 1390 27529 1424 27563
rect 1516 27529 1550 27563
rect 1642 27529 1676 27563
rect 1768 27529 1802 27563
rect 1894 27529 1928 27563
rect 2020 27529 2054 27563
rect 382 23744 416 23778
rect 508 23744 542 23778
rect 634 23744 668 23778
rect 760 23744 794 23778
rect 886 23744 920 23778
rect 1012 23744 1046 23778
rect 1138 23744 1172 23778
rect 1264 23744 1298 23778
rect 1390 23744 1424 23778
rect 1516 23744 1550 23778
rect 1642 23744 1676 23778
rect 1768 23744 1802 23778
rect 1894 23744 1928 23778
rect 2020 23744 2054 23778
rect 382 23634 416 23668
rect 508 23634 542 23668
rect 634 23634 668 23668
rect 760 23634 794 23668
rect 886 23634 920 23668
rect 1012 23634 1046 23668
rect 1138 23634 1172 23668
rect 1264 23634 1298 23668
rect 1390 23634 1424 23668
rect 1516 23634 1550 23668
rect 1642 23634 1676 23668
rect 1768 23634 1802 23668
rect 1894 23634 1928 23668
rect 2020 23634 2054 23668
rect 1390 22273 1424 22307
rect 382 19849 416 19883
rect 508 19849 542 19883
rect 634 19849 668 19883
rect 760 19849 794 19883
rect 886 19849 920 19883
rect 1012 19849 1046 19883
rect 1138 19849 1172 19883
rect 1264 19849 1298 19883
rect 1642 22273 1676 22307
rect 1516 19849 1550 19883
rect 1894 22273 1928 22307
rect 1768 19849 1802 19883
rect 2020 19849 2054 19883
rect 382 19739 416 19773
rect 508 19739 542 19773
rect 634 19739 668 19773
rect 760 19739 794 19773
rect 886 19739 920 19773
rect 1012 19739 1046 19773
rect 1138 19739 1172 19773
rect 1264 19739 1298 19773
rect 1390 19739 1424 19773
rect 1516 19739 1550 19773
rect 1642 19739 1676 19773
rect 1768 19739 1802 19773
rect 1894 19739 1928 19773
rect 2020 19739 2054 19773
rect 382 15954 416 15988
rect 508 15954 542 15988
rect 634 15954 668 15988
rect 760 15954 794 15988
rect 886 15954 920 15988
rect 1012 15954 1046 15988
rect 1138 15954 1172 15988
rect 1264 15954 1298 15988
rect 1390 15954 1424 15988
rect 1516 15954 1550 15988
rect 1642 15954 1676 15988
rect 1768 15954 1802 15988
rect 1894 15954 1928 15988
rect 2020 15954 2054 15988
rect 382 15844 416 15878
rect 508 15844 542 15878
rect 634 15844 668 15878
rect 760 15844 794 15878
rect 886 15844 920 15878
rect 1012 15844 1046 15878
rect 1138 15844 1172 15878
rect 1264 15844 1298 15878
rect 1390 15844 1424 15878
rect 1516 15844 1550 15878
rect 1642 15844 1676 15878
rect 1768 15844 1802 15878
rect 1894 15844 1928 15878
rect 2020 15844 2054 15878
rect 382 12059 416 12093
rect 508 12059 542 12093
rect 634 12059 668 12093
rect 760 12059 794 12093
rect 886 12059 920 12093
rect 1012 12059 1046 12093
rect 1138 12059 1172 12093
rect 1264 12059 1298 12093
rect 1390 12059 1424 12093
rect 1516 12059 1550 12093
rect 1642 12059 1676 12093
rect 1768 12059 1802 12093
rect 1894 12059 1928 12093
rect 2020 12059 2054 12093
rect 382 11949 416 11983
rect 508 11949 542 11983
rect 634 11949 668 11983
rect 760 11949 794 11983
rect 886 11949 920 11983
rect 1012 11949 1046 11983
rect 1138 11949 1172 11983
rect 1264 11949 1298 11983
rect 1390 11949 1424 11983
rect 1516 11949 1550 11983
rect 1642 11949 1676 11983
rect 1768 11949 1802 11983
rect 1894 11949 1928 11983
rect 2020 11949 2054 11983
rect 382 8164 416 8198
rect 508 8164 542 8198
rect 634 8164 668 8198
rect 760 8164 794 8198
rect 886 8164 920 8198
rect 1012 8164 1046 8198
rect 1138 8164 1172 8198
rect 1264 8164 1298 8198
rect 1390 8164 1424 8198
rect 1516 8164 1550 8198
rect 1642 8164 1676 8198
rect 1768 8164 1802 8198
rect 1894 8164 1928 8198
rect 2020 8164 2054 8198
rect 382 8054 416 8088
rect 508 8054 542 8088
rect 634 8054 668 8088
rect 760 8054 794 8088
rect 886 8054 920 8088
rect 1012 8054 1046 8088
rect 1138 8054 1172 8088
rect 1264 8054 1298 8088
rect 1390 8054 1424 8088
rect 1516 8054 1550 8088
rect 1642 8054 1676 8088
rect 1768 8054 1802 8088
rect 1894 8054 1928 8088
rect 2020 5423 2054 5457
rect 2146 5423 2180 5457
rect 2272 5423 2306 5457
rect 2398 5423 2432 5457
rect 2524 5423 2558 5457
rect 2650 5423 2684 5457
rect 2776 5423 2810 5457
rect 2902 5423 2936 5457
rect 3028 5423 3062 5457
rect 382 4269 416 4303
rect 508 4269 542 4303
rect 634 4269 668 4303
rect 760 4269 794 4303
rect 886 4269 920 4303
rect 1012 4269 1046 4303
rect 1138 4269 1172 4303
rect 1264 4269 1298 4303
rect 1390 4269 1424 4303
rect 1516 4269 1550 4303
rect 1642 4269 1676 4303
rect 1768 4269 1802 4303
rect 1894 4269 1928 4303
rect 382 4159 416 4193
rect 508 4159 542 4193
rect 634 4159 668 4193
rect 760 4159 794 4193
rect 886 4159 920 4193
rect 1012 4159 1046 4193
rect 1138 4159 1172 4193
rect 1264 4159 1298 4193
rect 1390 4159 1424 4193
rect 1516 4159 1550 4193
rect 1642 4159 1676 4193
rect 1768 4159 1802 4193
rect 1894 4159 1928 4193
rect 382 374 416 408
rect 508 374 542 408
rect 634 374 668 408
rect 760 374 794 408
rect 886 374 920 408
rect 1012 374 1046 408
rect 1138 374 1172 408
rect 1264 374 1298 408
rect 1390 374 1424 408
rect 1516 374 1550 408
rect 1642 374 1676 408
rect 1768 374 1802 408
rect 1894 374 1928 408
rect 2020 374 2054 408
rect 2146 374 2180 408
rect 2272 374 2306 408
rect 2398 374 2432 408
rect 2524 374 2558 408
rect 2650 374 2684 408
rect 2776 374 2810 408
rect 2902 374 2936 408
rect 3028 374 3062 408
<< psubdiff >>
rect 2148 -554 3498 -553
rect 2148 -587 2274 -554
rect 2148 -621 2149 -587
rect 2183 -588 2274 -587
rect 2308 -588 2342 -554
rect 2376 -588 2410 -554
rect 2444 -588 2478 -554
rect 2512 -588 2546 -554
rect 2580 -588 2614 -554
rect 2648 -588 2682 -554
rect 2716 -588 2750 -554
rect 2784 -588 2818 -554
rect 2852 -588 2886 -554
rect 2920 -588 2954 -554
rect 2988 -588 3022 -554
rect 3056 -588 3090 -554
rect 3124 -588 3158 -554
rect 3192 -588 3226 -554
rect 3260 -588 3294 -554
rect 3328 -588 3362 -554
rect 3396 -588 3430 -554
rect 3464 -588 3498 -554
rect 2183 -589 3498 -588
rect 2183 -621 2184 -589
rect 2148 -655 2184 -621
rect 3462 -622 3498 -589
rect 2148 -689 2149 -655
rect 2183 -689 2184 -655
rect 2148 -723 2184 -689
rect 3462 -656 3463 -622
rect 3497 -656 3498 -622
rect 3462 -690 3498 -656
rect 2148 -757 2149 -723
rect 2183 -757 2184 -723
rect 2148 -791 2184 -757
rect 2148 -825 2149 -791
rect 2183 -825 2184 -791
rect 2148 -859 2184 -825
rect 2148 -893 2149 -859
rect 2183 -893 2184 -859
rect 2148 -994 2184 -893
rect 3462 -724 3463 -690
rect 3497 -724 3498 -690
rect 3462 -758 3498 -724
rect 3462 -792 3463 -758
rect 3497 -792 3498 -758
rect 3462 -826 3498 -792
rect 3462 -860 3463 -826
rect 3497 -860 3498 -826
rect 3462 -894 3498 -860
rect 3462 -928 3463 -894
rect 3497 -928 3498 -894
rect 3462 -962 3498 -928
rect 3462 -994 3463 -962
rect 2148 -995 3463 -994
rect 2148 -1029 2182 -995
rect 2216 -1029 2250 -995
rect 2284 -1029 2318 -995
rect 2352 -1029 2386 -995
rect 2420 -1029 2454 -995
rect 2488 -1029 2522 -995
rect 2556 -1029 2590 -995
rect 2624 -1029 2658 -995
rect 2692 -1029 2726 -995
rect 2760 -1029 2794 -995
rect 2828 -1029 2862 -995
rect 2896 -1029 2930 -995
rect 2964 -1029 2998 -995
rect 3032 -1029 3066 -995
rect 3100 -1029 3134 -995
rect 3168 -1029 3202 -995
rect 3236 -1029 3270 -995
rect 3304 -1029 3338 -995
rect 3372 -996 3463 -995
rect 3497 -996 3498 -962
rect 3372 -1029 3498 -996
rect 2148 -1030 3498 -1029
<< mvpsubdiff >>
rect 256 27680 2180 27681
rect 256 27647 344 27680
rect 256 27613 257 27647
rect 291 27646 344 27647
rect 378 27646 412 27680
rect 446 27646 480 27680
rect 514 27646 548 27680
rect 582 27646 616 27680
rect 650 27646 684 27680
rect 718 27646 752 27680
rect 786 27646 820 27680
rect 854 27646 888 27680
rect 922 27646 956 27680
rect 990 27646 1024 27680
rect 1058 27646 1092 27680
rect 1126 27646 1160 27680
rect 1194 27646 1228 27680
rect 1262 27646 1296 27680
rect 1330 27646 1364 27680
rect 1398 27646 1432 27680
rect 1466 27646 1500 27680
rect 1534 27646 1568 27680
rect 1602 27646 1636 27680
rect 1670 27646 1704 27680
rect 1738 27646 1772 27680
rect 1806 27646 1840 27680
rect 1874 27646 1908 27680
rect 1942 27646 1976 27680
rect 2010 27646 2044 27680
rect 2078 27646 2112 27680
rect 2146 27646 2180 27680
rect 291 27645 2180 27646
rect 291 27613 292 27645
rect 256 27579 292 27613
rect 256 27545 257 27579
rect 291 27545 292 27579
rect 2144 27571 2180 27645
rect 256 27511 292 27545
rect 256 27477 257 27511
rect 291 27477 292 27511
rect 2144 27537 2145 27571
rect 2179 27537 2180 27571
rect 2144 27503 2180 27537
rect 256 27443 292 27477
rect 256 27409 257 27443
rect 291 27409 292 27443
rect 256 27375 292 27409
rect 256 27341 257 27375
rect 291 27341 292 27375
rect 256 27307 292 27341
rect 256 27273 257 27307
rect 291 27273 292 27307
rect 256 27239 292 27273
rect 256 27205 257 27239
rect 291 27205 292 27239
rect 256 27171 292 27205
rect 256 27137 257 27171
rect 291 27137 292 27171
rect 256 27103 292 27137
rect 256 27069 257 27103
rect 291 27069 292 27103
rect 256 27035 292 27069
rect 256 27001 257 27035
rect 291 27001 292 27035
rect 256 26967 292 27001
rect 256 26933 257 26967
rect 291 26933 292 26967
rect 256 26899 292 26933
rect 256 26865 257 26899
rect 291 26865 292 26899
rect 256 26831 292 26865
rect 256 26797 257 26831
rect 291 26797 292 26831
rect 256 26763 292 26797
rect 256 26729 257 26763
rect 291 26729 292 26763
rect 256 26695 292 26729
rect 256 26661 257 26695
rect 291 26661 292 26695
rect 256 26627 292 26661
rect 256 26593 257 26627
rect 291 26593 292 26627
rect 256 26559 292 26593
rect 256 26525 257 26559
rect 291 26525 292 26559
rect 256 26491 292 26525
rect 256 26457 257 26491
rect 291 26457 292 26491
rect 256 26423 292 26457
rect 256 26389 257 26423
rect 291 26389 292 26423
rect 256 26355 292 26389
rect 256 26321 257 26355
rect 291 26321 292 26355
rect 256 26287 292 26321
rect 256 26253 257 26287
rect 291 26253 292 26287
rect 256 26219 292 26253
rect 256 26185 257 26219
rect 291 26185 292 26219
rect 256 26151 292 26185
rect 256 26117 257 26151
rect 291 26117 292 26151
rect 256 26083 292 26117
rect 256 26049 257 26083
rect 291 26049 292 26083
rect 256 26015 292 26049
rect 256 25981 257 26015
rect 291 25981 292 26015
rect 256 25947 292 25981
rect 256 25913 257 25947
rect 291 25913 292 25947
rect 256 25879 292 25913
rect 256 25845 257 25879
rect 291 25845 292 25879
rect 256 25811 292 25845
rect 256 25777 257 25811
rect 291 25777 292 25811
rect 256 25743 292 25777
rect 256 25709 257 25743
rect 291 25709 292 25743
rect 256 25675 292 25709
rect 256 25641 257 25675
rect 291 25641 292 25675
rect 256 25607 292 25641
rect 256 25573 257 25607
rect 291 25573 292 25607
rect 256 25539 292 25573
rect 256 25505 257 25539
rect 291 25505 292 25539
rect 256 25471 292 25505
rect 256 25437 257 25471
rect 291 25437 292 25471
rect 256 25403 292 25437
rect 256 25369 257 25403
rect 291 25369 292 25403
rect 256 25335 292 25369
rect 256 25301 257 25335
rect 291 25301 292 25335
rect 256 25267 292 25301
rect 256 25233 257 25267
rect 291 25233 292 25267
rect 256 25199 292 25233
rect 256 25165 257 25199
rect 291 25165 292 25199
rect 256 25131 292 25165
rect 256 25097 257 25131
rect 291 25097 292 25131
rect 256 25063 292 25097
rect 256 25029 257 25063
rect 291 25029 292 25063
rect 256 24995 292 25029
rect 256 24961 257 24995
rect 291 24961 292 24995
rect 256 24927 292 24961
rect 256 24893 257 24927
rect 291 24893 292 24927
rect 256 24859 292 24893
rect 256 24825 257 24859
rect 291 24825 292 24859
rect 256 24791 292 24825
rect 256 24757 257 24791
rect 291 24757 292 24791
rect 256 24723 292 24757
rect 256 24689 257 24723
rect 291 24689 292 24723
rect 256 24655 292 24689
rect 256 24621 257 24655
rect 291 24621 292 24655
rect 256 24587 292 24621
rect 256 24553 257 24587
rect 291 24553 292 24587
rect 256 24519 292 24553
rect 256 24485 257 24519
rect 291 24485 292 24519
rect 256 24451 292 24485
rect 256 24417 257 24451
rect 291 24417 292 24451
rect 256 24383 292 24417
rect 256 24349 257 24383
rect 291 24349 292 24383
rect 256 24315 292 24349
rect 256 24281 257 24315
rect 291 24281 292 24315
rect 256 24247 292 24281
rect 256 24213 257 24247
rect 291 24213 292 24247
rect 256 24179 292 24213
rect 256 24145 257 24179
rect 291 24145 292 24179
rect 256 24111 292 24145
rect 256 24077 257 24111
rect 291 24077 292 24111
rect 256 24043 292 24077
rect 256 24009 257 24043
rect 291 24009 292 24043
rect 256 23975 292 24009
rect 256 23941 257 23975
rect 291 23941 292 23975
rect 256 23907 292 23941
rect 256 23873 257 23907
rect 291 23873 292 23907
rect 256 23839 292 23873
rect 256 23805 257 23839
rect 291 23805 292 23839
rect 256 23771 292 23805
rect 2144 27469 2145 27503
rect 2179 27469 2180 27503
rect 2144 27435 2180 27469
rect 2144 27401 2145 27435
rect 2179 27401 2180 27435
rect 2144 27367 2180 27401
rect 2144 27333 2145 27367
rect 2179 27333 2180 27367
rect 2144 27299 2180 27333
rect 2144 27265 2145 27299
rect 2179 27265 2180 27299
rect 2144 27231 2180 27265
rect 2144 27197 2145 27231
rect 2179 27197 2180 27231
rect 2144 27163 2180 27197
rect 2144 27129 2145 27163
rect 2179 27129 2180 27163
rect 2144 27095 2180 27129
rect 2144 27061 2145 27095
rect 2179 27061 2180 27095
rect 2144 27027 2180 27061
rect 2144 26993 2145 27027
rect 2179 26993 2180 27027
rect 2144 26959 2180 26993
rect 2144 26925 2145 26959
rect 2179 26925 2180 26959
rect 2144 26891 2180 26925
rect 2144 26857 2145 26891
rect 2179 26857 2180 26891
rect 2144 26823 2180 26857
rect 2144 26789 2145 26823
rect 2179 26789 2180 26823
rect 2144 26755 2180 26789
rect 2144 26721 2145 26755
rect 2179 26721 2180 26755
rect 2144 26687 2180 26721
rect 2144 26653 2145 26687
rect 2179 26653 2180 26687
rect 2144 26619 2180 26653
rect 2144 26585 2145 26619
rect 2179 26585 2180 26619
rect 2144 26551 2180 26585
rect 2144 26517 2145 26551
rect 2179 26517 2180 26551
rect 2144 26483 2180 26517
rect 2144 26449 2145 26483
rect 2179 26449 2180 26483
rect 2144 26415 2180 26449
rect 2144 26381 2145 26415
rect 2179 26381 2180 26415
rect 2144 26347 2180 26381
rect 2144 26313 2145 26347
rect 2179 26313 2180 26347
rect 2144 26279 2180 26313
rect 2144 26245 2145 26279
rect 2179 26245 2180 26279
rect 2144 26211 2180 26245
rect 2144 26177 2145 26211
rect 2179 26177 2180 26211
rect 2144 26143 2180 26177
rect 2144 26109 2145 26143
rect 2179 26109 2180 26143
rect 2144 26075 2180 26109
rect 2144 26041 2145 26075
rect 2179 26041 2180 26075
rect 2144 26007 2180 26041
rect 2144 25973 2145 26007
rect 2179 25973 2180 26007
rect 2144 25939 2180 25973
rect 2144 25905 2145 25939
rect 2179 25905 2180 25939
rect 2144 25871 2180 25905
rect 2144 25837 2145 25871
rect 2179 25837 2180 25871
rect 2144 25803 2180 25837
rect 2144 25769 2145 25803
rect 2179 25769 2180 25803
rect 2144 25735 2180 25769
rect 2144 25701 2145 25735
rect 2179 25701 2180 25735
rect 2144 25667 2180 25701
rect 2144 25633 2145 25667
rect 2179 25633 2180 25667
rect 2144 25599 2180 25633
rect 2144 25565 2145 25599
rect 2179 25565 2180 25599
rect 2144 25531 2180 25565
rect 2144 25497 2145 25531
rect 2179 25497 2180 25531
rect 2144 25463 2180 25497
rect 2144 25429 2145 25463
rect 2179 25429 2180 25463
rect 2144 25395 2180 25429
rect 2144 25361 2145 25395
rect 2179 25361 2180 25395
rect 2144 25327 2180 25361
rect 2144 25293 2145 25327
rect 2179 25293 2180 25327
rect 2144 25259 2180 25293
rect 2144 25225 2145 25259
rect 2179 25225 2180 25259
rect 2144 25191 2180 25225
rect 2144 25157 2145 25191
rect 2179 25157 2180 25191
rect 2144 25123 2180 25157
rect 2144 25089 2145 25123
rect 2179 25089 2180 25123
rect 2144 25055 2180 25089
rect 2144 25021 2145 25055
rect 2179 25021 2180 25055
rect 2144 24987 2180 25021
rect 2144 24953 2145 24987
rect 2179 24953 2180 24987
rect 2144 24919 2180 24953
rect 2144 24885 2145 24919
rect 2179 24885 2180 24919
rect 2144 24851 2180 24885
rect 2144 24817 2145 24851
rect 2179 24817 2180 24851
rect 2144 24783 2180 24817
rect 2144 24749 2145 24783
rect 2179 24749 2180 24783
rect 2144 24715 2180 24749
rect 2144 24681 2145 24715
rect 2179 24681 2180 24715
rect 2144 24647 2180 24681
rect 2144 24613 2145 24647
rect 2179 24613 2180 24647
rect 2144 24579 2180 24613
rect 2144 24545 2145 24579
rect 2179 24545 2180 24579
rect 2144 24511 2180 24545
rect 2144 24477 2145 24511
rect 2179 24477 2180 24511
rect 2144 24443 2180 24477
rect 2144 24409 2145 24443
rect 2179 24409 2180 24443
rect 2144 24375 2180 24409
rect 2144 24341 2145 24375
rect 2179 24341 2180 24375
rect 2144 24307 2180 24341
rect 2144 24273 2145 24307
rect 2179 24273 2180 24307
rect 2144 24239 2180 24273
rect 2144 24205 2145 24239
rect 2179 24205 2180 24239
rect 2144 24171 2180 24205
rect 2144 24137 2145 24171
rect 2179 24137 2180 24171
rect 2144 24103 2180 24137
rect 2144 24069 2145 24103
rect 2179 24069 2180 24103
rect 2144 24035 2180 24069
rect 2144 24001 2145 24035
rect 2179 24001 2180 24035
rect 2144 23967 2180 24001
rect 2144 23933 2145 23967
rect 2179 23933 2180 23967
rect 2144 23899 2180 23933
rect 2144 23865 2145 23899
rect 2179 23865 2180 23899
rect 2144 23831 2180 23865
rect 256 23737 257 23771
rect 291 23737 292 23771
rect 256 23703 292 23737
rect 2144 23797 2145 23831
rect 2179 23797 2180 23831
rect 2144 23763 2180 23797
rect 256 23669 257 23703
rect 291 23669 292 23703
rect 2144 23729 2145 23763
rect 2179 23729 2180 23763
rect 2144 23695 2180 23729
rect 256 23635 292 23669
rect 256 23601 257 23635
rect 291 23601 292 23635
rect 2144 23661 2145 23695
rect 2179 23661 2180 23695
rect 2144 23627 2180 23661
rect 256 23567 292 23601
rect 256 23533 257 23567
rect 291 23533 292 23567
rect 256 23499 292 23533
rect 256 23465 257 23499
rect 291 23465 292 23499
rect 256 23431 292 23465
rect 256 23397 257 23431
rect 291 23397 292 23431
rect 256 23363 292 23397
rect 256 23329 257 23363
rect 291 23329 292 23363
rect 256 23295 292 23329
rect 256 23261 257 23295
rect 291 23261 292 23295
rect 256 23227 292 23261
rect 256 23193 257 23227
rect 291 23193 292 23227
rect 256 23159 292 23193
rect 256 23125 257 23159
rect 291 23125 292 23159
rect 256 23091 292 23125
rect 256 23057 257 23091
rect 291 23057 292 23091
rect 256 23023 292 23057
rect 256 22989 257 23023
rect 291 22989 292 23023
rect 256 22955 292 22989
rect 256 22921 257 22955
rect 291 22921 292 22955
rect 256 22887 292 22921
rect 256 22853 257 22887
rect 291 22853 292 22887
rect 256 22819 292 22853
rect 256 22785 257 22819
rect 291 22785 292 22819
rect 256 22751 292 22785
rect 256 22717 257 22751
rect 291 22717 292 22751
rect 256 22683 292 22717
rect 256 22649 257 22683
rect 291 22649 292 22683
rect 256 22615 292 22649
rect 256 22581 257 22615
rect 291 22581 292 22615
rect 256 22547 292 22581
rect 256 22513 257 22547
rect 291 22513 292 22547
rect 256 22479 292 22513
rect 256 22445 257 22479
rect 291 22445 292 22479
rect 256 22411 292 22445
rect 256 22377 257 22411
rect 291 22377 292 22411
rect 256 22343 292 22377
rect 256 22309 257 22343
rect 291 22309 292 22343
rect 2144 23593 2145 23627
rect 2179 23593 2180 23627
rect 2144 23559 2180 23593
rect 2144 23525 2145 23559
rect 2179 23525 2180 23559
rect 2144 23491 2180 23525
rect 2144 23457 2145 23491
rect 2179 23457 2180 23491
rect 2144 23423 2180 23457
rect 2144 23389 2145 23423
rect 2179 23389 2180 23423
rect 2144 23355 2180 23389
rect 2144 23321 2145 23355
rect 2179 23321 2180 23355
rect 2144 23287 2180 23321
rect 2144 23253 2145 23287
rect 2179 23253 2180 23287
rect 2144 23219 2180 23253
rect 2144 23185 2145 23219
rect 2179 23185 2180 23219
rect 2144 23151 2180 23185
rect 2144 23117 2145 23151
rect 2179 23117 2180 23151
rect 2144 23083 2180 23117
rect 2144 23049 2145 23083
rect 2179 23049 2180 23083
rect 2144 23015 2180 23049
rect 2144 22981 2145 23015
rect 2179 22981 2180 23015
rect 2144 22947 2180 22981
rect 2144 22913 2145 22947
rect 2179 22913 2180 22947
rect 2144 22879 2180 22913
rect 2144 22845 2145 22879
rect 2179 22845 2180 22879
rect 2144 22811 2180 22845
rect 2144 22777 2145 22811
rect 2179 22777 2180 22811
rect 2144 22743 2180 22777
rect 2144 22709 2145 22743
rect 2179 22709 2180 22743
rect 2144 22675 2180 22709
rect 2144 22641 2145 22675
rect 2179 22641 2180 22675
rect 2144 22607 2180 22641
rect 2144 22573 2145 22607
rect 2179 22573 2180 22607
rect 2144 22539 2180 22573
rect 2144 22505 2145 22539
rect 2179 22505 2180 22539
rect 2144 22471 2180 22505
rect 2144 22437 2145 22471
rect 2179 22437 2180 22471
rect 2144 22403 2180 22437
rect 2144 22369 2145 22403
rect 2179 22369 2180 22403
rect 2144 22335 2180 22369
rect 256 22275 292 22309
rect 256 22241 257 22275
rect 291 22241 292 22275
rect 256 22207 292 22241
rect 256 22173 257 22207
rect 291 22173 292 22207
rect 256 22139 292 22173
rect 256 22105 257 22139
rect 291 22105 292 22139
rect 256 22071 292 22105
rect 256 22037 257 22071
rect 291 22037 292 22071
rect 256 22003 292 22037
rect 256 21969 257 22003
rect 291 21969 292 22003
rect 256 21935 292 21969
rect 256 21901 257 21935
rect 291 21901 292 21935
rect 256 21867 292 21901
rect 256 21833 257 21867
rect 291 21833 292 21867
rect 256 21799 292 21833
rect 256 21765 257 21799
rect 291 21765 292 21799
rect 256 21731 292 21765
rect 256 21697 257 21731
rect 291 21697 292 21731
rect 256 21663 292 21697
rect 256 21629 257 21663
rect 291 21629 292 21663
rect 256 21595 292 21629
rect 256 21561 257 21595
rect 291 21561 292 21595
rect 256 21527 292 21561
rect 256 21493 257 21527
rect 291 21493 292 21527
rect 256 21459 292 21493
rect 256 21425 257 21459
rect 291 21425 292 21459
rect 256 21391 292 21425
rect 256 21357 257 21391
rect 291 21357 292 21391
rect 256 21323 292 21357
rect 256 21289 257 21323
rect 291 21289 292 21323
rect 256 21255 292 21289
rect 256 21221 257 21255
rect 291 21221 292 21255
rect 256 21187 292 21221
rect 256 21153 257 21187
rect 291 21153 292 21187
rect 256 21119 292 21153
rect 256 21085 257 21119
rect 291 21085 292 21119
rect 256 21051 292 21085
rect 256 21017 257 21051
rect 291 21017 292 21051
rect 256 20983 292 21017
rect 256 20949 257 20983
rect 291 20949 292 20983
rect 256 20915 292 20949
rect 256 20881 257 20915
rect 291 20881 292 20915
rect 256 20847 292 20881
rect 256 20813 257 20847
rect 291 20813 292 20847
rect 256 20779 292 20813
rect 256 20745 257 20779
rect 291 20745 292 20779
rect 256 20711 292 20745
rect 256 20677 257 20711
rect 291 20677 292 20711
rect 256 20643 292 20677
rect 256 20609 257 20643
rect 291 20609 292 20643
rect 256 20575 292 20609
rect 256 20541 257 20575
rect 291 20541 292 20575
rect 256 20507 292 20541
rect 256 20473 257 20507
rect 291 20473 292 20507
rect 256 20439 292 20473
rect 256 20405 257 20439
rect 291 20405 292 20439
rect 256 20371 292 20405
rect 256 20337 257 20371
rect 291 20337 292 20371
rect 256 20303 292 20337
rect 256 20269 257 20303
rect 291 20269 292 20303
rect 256 20235 292 20269
rect 256 20201 257 20235
rect 291 20201 292 20235
rect 256 20167 292 20201
rect 256 20133 257 20167
rect 291 20133 292 20167
rect 256 20099 292 20133
rect 256 20065 257 20099
rect 291 20065 292 20099
rect 256 20031 292 20065
rect 256 19997 257 20031
rect 291 19997 292 20031
rect 256 19963 292 19997
rect 256 19929 257 19963
rect 291 19929 292 19963
rect 256 19895 292 19929
rect 256 19861 257 19895
rect 291 19861 292 19895
rect 256 19827 292 19861
rect 2144 22301 2145 22335
rect 2179 22301 2180 22335
rect 2144 22267 2180 22301
rect 2144 22233 2145 22267
rect 2179 22233 2180 22267
rect 2144 22199 2180 22233
rect 2144 22165 2145 22199
rect 2179 22165 2180 22199
rect 2144 22131 2180 22165
rect 2144 22097 2145 22131
rect 2179 22097 2180 22131
rect 2144 22063 2180 22097
rect 2144 22029 2145 22063
rect 2179 22029 2180 22063
rect 2144 21995 2180 22029
rect 2144 21961 2145 21995
rect 2179 21961 2180 21995
rect 2144 21927 2180 21961
rect 2144 21893 2145 21927
rect 2179 21893 2180 21927
rect 2144 21859 2180 21893
rect 2144 21825 2145 21859
rect 2179 21825 2180 21859
rect 2144 21791 2180 21825
rect 2144 21757 2145 21791
rect 2179 21757 2180 21791
rect 2144 21723 2180 21757
rect 2144 21689 2145 21723
rect 2179 21689 2180 21723
rect 2144 21655 2180 21689
rect 2144 21621 2145 21655
rect 2179 21621 2180 21655
rect 2144 21587 2180 21621
rect 2144 21553 2145 21587
rect 2179 21553 2180 21587
rect 2144 21519 2180 21553
rect 2144 21485 2145 21519
rect 2179 21485 2180 21519
rect 2144 21451 2180 21485
rect 2144 21417 2145 21451
rect 2179 21417 2180 21451
rect 2144 21383 2180 21417
rect 2144 21349 2145 21383
rect 2179 21349 2180 21383
rect 2144 21315 2180 21349
rect 2144 21281 2145 21315
rect 2179 21281 2180 21315
rect 2144 21247 2180 21281
rect 2144 21213 2145 21247
rect 2179 21213 2180 21247
rect 2144 21179 2180 21213
rect 2144 21145 2145 21179
rect 2179 21145 2180 21179
rect 2144 21111 2180 21145
rect 2144 21077 2145 21111
rect 2179 21077 2180 21111
rect 2144 21043 2180 21077
rect 2144 21009 2145 21043
rect 2179 21009 2180 21043
rect 2144 20975 2180 21009
rect 2144 20941 2145 20975
rect 2179 20941 2180 20975
rect 2144 20907 2180 20941
rect 2144 20873 2145 20907
rect 2179 20873 2180 20907
rect 2144 20839 2180 20873
rect 2144 20805 2145 20839
rect 2179 20805 2180 20839
rect 2144 20771 2180 20805
rect 2144 20737 2145 20771
rect 2179 20737 2180 20771
rect 2144 20703 2180 20737
rect 2144 20669 2145 20703
rect 2179 20669 2180 20703
rect 2144 20635 2180 20669
rect 2144 20601 2145 20635
rect 2179 20601 2180 20635
rect 2144 20567 2180 20601
rect 2144 20533 2145 20567
rect 2179 20533 2180 20567
rect 2144 20499 2180 20533
rect 2144 20465 2145 20499
rect 2179 20465 2180 20499
rect 2144 20431 2180 20465
rect 2144 20397 2145 20431
rect 2179 20397 2180 20431
rect 2144 20363 2180 20397
rect 2144 20329 2145 20363
rect 2179 20329 2180 20363
rect 2144 20295 2180 20329
rect 2144 20261 2145 20295
rect 2179 20261 2180 20295
rect 2144 20227 2180 20261
rect 2144 20193 2145 20227
rect 2179 20193 2180 20227
rect 2144 20159 2180 20193
rect 2144 20125 2145 20159
rect 2179 20125 2180 20159
rect 2144 20091 2180 20125
rect 2144 20057 2145 20091
rect 2179 20057 2180 20091
rect 2144 20023 2180 20057
rect 2144 19989 2145 20023
rect 2179 19989 2180 20023
rect 2144 19955 2180 19989
rect 2144 19921 2145 19955
rect 2179 19921 2180 19955
rect 2144 19887 2180 19921
rect 2144 19853 2145 19887
rect 2179 19853 2180 19887
rect 256 19793 257 19827
rect 291 19793 292 19827
rect 256 19759 292 19793
rect 2144 19819 2180 19853
rect 2144 19785 2145 19819
rect 2179 19785 2180 19819
rect 256 19725 257 19759
rect 291 19725 292 19759
rect 256 19691 292 19725
rect 2144 19751 2180 19785
rect 2144 19717 2145 19751
rect 2179 19717 2180 19751
rect 256 19657 257 19691
rect 291 19657 292 19691
rect 256 19623 292 19657
rect 256 19589 257 19623
rect 291 19589 292 19623
rect 256 19555 292 19589
rect 256 19521 257 19555
rect 291 19521 292 19555
rect 256 19487 292 19521
rect 256 19453 257 19487
rect 291 19453 292 19487
rect 256 19419 292 19453
rect 256 19385 257 19419
rect 291 19385 292 19419
rect 256 19351 292 19385
rect 256 19317 257 19351
rect 291 19317 292 19351
rect 256 19283 292 19317
rect 256 19249 257 19283
rect 291 19249 292 19283
rect 256 19215 292 19249
rect 256 19181 257 19215
rect 291 19181 292 19215
rect 256 19147 292 19181
rect 256 19113 257 19147
rect 291 19113 292 19147
rect 256 19079 292 19113
rect 256 19045 257 19079
rect 291 19045 292 19079
rect 256 19011 292 19045
rect 256 18977 257 19011
rect 291 18977 292 19011
rect 256 18943 292 18977
rect 256 18909 257 18943
rect 291 18909 292 18943
rect 256 18875 292 18909
rect 256 18841 257 18875
rect 291 18841 292 18875
rect 256 18807 292 18841
rect 256 18773 257 18807
rect 291 18773 292 18807
rect 256 18739 292 18773
rect 256 18705 257 18739
rect 291 18705 292 18739
rect 256 18671 292 18705
rect 256 18637 257 18671
rect 291 18637 292 18671
rect 256 18603 292 18637
rect 256 18569 257 18603
rect 291 18569 292 18603
rect 256 18535 292 18569
rect 256 18501 257 18535
rect 291 18501 292 18535
rect 256 18467 292 18501
rect 256 18433 257 18467
rect 291 18433 292 18467
rect 256 18399 292 18433
rect 256 18365 257 18399
rect 291 18365 292 18399
rect 256 18331 292 18365
rect 256 18297 257 18331
rect 291 18297 292 18331
rect 256 18263 292 18297
rect 256 18229 257 18263
rect 291 18229 292 18263
rect 256 18195 292 18229
rect 256 18161 257 18195
rect 291 18161 292 18195
rect 256 18127 292 18161
rect 256 18093 257 18127
rect 291 18093 292 18127
rect 256 18059 292 18093
rect 256 18025 257 18059
rect 291 18025 292 18059
rect 256 17991 292 18025
rect 256 17957 257 17991
rect 291 17957 292 17991
rect 256 17923 292 17957
rect 256 17889 257 17923
rect 291 17889 292 17923
rect 256 17855 292 17889
rect 256 17821 257 17855
rect 291 17821 292 17855
rect 256 17787 292 17821
rect 256 17753 257 17787
rect 291 17753 292 17787
rect 256 17719 292 17753
rect 256 17685 257 17719
rect 291 17685 292 17719
rect 256 17651 292 17685
rect 256 17617 257 17651
rect 291 17617 292 17651
rect 256 17583 292 17617
rect 256 17549 257 17583
rect 291 17549 292 17583
rect 256 17515 292 17549
rect 256 17481 257 17515
rect 291 17481 292 17515
rect 256 17447 292 17481
rect 256 17413 257 17447
rect 291 17413 292 17447
rect 256 17379 292 17413
rect 256 17345 257 17379
rect 291 17345 292 17379
rect 256 17311 292 17345
rect 256 17277 257 17311
rect 291 17277 292 17311
rect 256 17243 292 17277
rect 256 17209 257 17243
rect 291 17209 292 17243
rect 256 17175 292 17209
rect 256 17141 257 17175
rect 291 17141 292 17175
rect 256 17107 292 17141
rect 256 17073 257 17107
rect 291 17073 292 17107
rect 256 17039 292 17073
rect 256 17005 257 17039
rect 291 17005 292 17039
rect 256 16971 292 17005
rect 256 16937 257 16971
rect 291 16937 292 16971
rect 256 16903 292 16937
rect 256 16869 257 16903
rect 291 16869 292 16903
rect 256 16835 292 16869
rect 256 16801 257 16835
rect 291 16801 292 16835
rect 256 16767 292 16801
rect 256 16733 257 16767
rect 291 16733 292 16767
rect 256 16699 292 16733
rect 256 16665 257 16699
rect 291 16665 292 16699
rect 256 16631 292 16665
rect 256 16597 257 16631
rect 291 16597 292 16631
rect 256 16563 292 16597
rect 256 16529 257 16563
rect 291 16529 292 16563
rect 256 16495 292 16529
rect 256 16461 257 16495
rect 291 16461 292 16495
rect 256 16427 292 16461
rect 256 16393 257 16427
rect 291 16393 292 16427
rect 256 16359 292 16393
rect 256 16325 257 16359
rect 291 16325 292 16359
rect 256 16291 292 16325
rect 256 16257 257 16291
rect 291 16257 292 16291
rect 256 16223 292 16257
rect 256 16189 257 16223
rect 291 16189 292 16223
rect 256 16155 292 16189
rect 256 16121 257 16155
rect 291 16121 292 16155
rect 256 16087 292 16121
rect 256 16053 257 16087
rect 291 16053 292 16087
rect 256 16019 292 16053
rect 256 15985 257 16019
rect 291 15985 292 16019
rect 2144 19683 2180 19717
rect 2144 19649 2145 19683
rect 2179 19649 2180 19683
rect 2144 19615 2180 19649
rect 2144 19581 2145 19615
rect 2179 19581 2180 19615
rect 2144 19547 2180 19581
rect 2144 19513 2145 19547
rect 2179 19513 2180 19547
rect 2144 19479 2180 19513
rect 2144 19445 2145 19479
rect 2179 19445 2180 19479
rect 2144 19411 2180 19445
rect 2144 19377 2145 19411
rect 2179 19377 2180 19411
rect 2144 19343 2180 19377
rect 2144 19309 2145 19343
rect 2179 19309 2180 19343
rect 2144 19275 2180 19309
rect 2144 19241 2145 19275
rect 2179 19241 2180 19275
rect 2144 19207 2180 19241
rect 2144 19173 2145 19207
rect 2179 19173 2180 19207
rect 2144 19139 2180 19173
rect 2144 19105 2145 19139
rect 2179 19105 2180 19139
rect 2144 19071 2180 19105
rect 2144 19037 2145 19071
rect 2179 19037 2180 19071
rect 2144 19003 2180 19037
rect 2144 18969 2145 19003
rect 2179 18969 2180 19003
rect 2144 18935 2180 18969
rect 2144 18901 2145 18935
rect 2179 18901 2180 18935
rect 2144 18867 2180 18901
rect 2144 18833 2145 18867
rect 2179 18833 2180 18867
rect 2144 18799 2180 18833
rect 2144 18765 2145 18799
rect 2179 18765 2180 18799
rect 2144 18731 2180 18765
rect 2144 18697 2145 18731
rect 2179 18697 2180 18731
rect 2144 18663 2180 18697
rect 2144 18629 2145 18663
rect 2179 18629 2180 18663
rect 2144 18595 2180 18629
rect 2144 18561 2145 18595
rect 2179 18561 2180 18595
rect 2144 18527 2180 18561
rect 2144 18493 2145 18527
rect 2179 18493 2180 18527
rect 2144 18459 2180 18493
rect 2144 18425 2145 18459
rect 2179 18425 2180 18459
rect 2144 18391 2180 18425
rect 2144 18357 2145 18391
rect 2179 18357 2180 18391
rect 2144 18323 2180 18357
rect 2144 18289 2145 18323
rect 2179 18289 2180 18323
rect 2144 18255 2180 18289
rect 2144 18221 2145 18255
rect 2179 18221 2180 18255
rect 2144 18187 2180 18221
rect 2144 18153 2145 18187
rect 2179 18153 2180 18187
rect 2144 18119 2180 18153
rect 2144 18085 2145 18119
rect 2179 18085 2180 18119
rect 2144 18051 2180 18085
rect 2144 18017 2145 18051
rect 2179 18017 2180 18051
rect 2144 17983 2180 18017
rect 2144 17949 2145 17983
rect 2179 17949 2180 17983
rect 2144 17915 2180 17949
rect 2144 17881 2145 17915
rect 2179 17881 2180 17915
rect 2144 17847 2180 17881
rect 2144 17813 2145 17847
rect 2179 17813 2180 17847
rect 2144 17779 2180 17813
rect 2144 17745 2145 17779
rect 2179 17745 2180 17779
rect 2144 17711 2180 17745
rect 2144 17677 2145 17711
rect 2179 17677 2180 17711
rect 2144 17643 2180 17677
rect 2144 17609 2145 17643
rect 2179 17609 2180 17643
rect 2144 17575 2180 17609
rect 2144 17541 2145 17575
rect 2179 17541 2180 17575
rect 2144 17507 2180 17541
rect 2144 17473 2145 17507
rect 2179 17473 2180 17507
rect 2144 17439 2180 17473
rect 2144 17405 2145 17439
rect 2179 17405 2180 17439
rect 2144 17371 2180 17405
rect 2144 17337 2145 17371
rect 2179 17337 2180 17371
rect 2144 17303 2180 17337
rect 2144 17269 2145 17303
rect 2179 17269 2180 17303
rect 2144 17235 2180 17269
rect 2144 17201 2145 17235
rect 2179 17201 2180 17235
rect 2144 17167 2180 17201
rect 2144 17133 2145 17167
rect 2179 17133 2180 17167
rect 2144 17099 2180 17133
rect 2144 17065 2145 17099
rect 2179 17065 2180 17099
rect 2144 17031 2180 17065
rect 2144 16997 2145 17031
rect 2179 16997 2180 17031
rect 2144 16963 2180 16997
rect 2144 16929 2145 16963
rect 2179 16929 2180 16963
rect 2144 16895 2180 16929
rect 2144 16861 2145 16895
rect 2179 16861 2180 16895
rect 2144 16827 2180 16861
rect 2144 16793 2145 16827
rect 2179 16793 2180 16827
rect 2144 16759 2180 16793
rect 2144 16725 2145 16759
rect 2179 16725 2180 16759
rect 2144 16691 2180 16725
rect 2144 16657 2145 16691
rect 2179 16657 2180 16691
rect 2144 16623 2180 16657
rect 2144 16589 2145 16623
rect 2179 16589 2180 16623
rect 2144 16555 2180 16589
rect 2144 16521 2145 16555
rect 2179 16521 2180 16555
rect 2144 16487 2180 16521
rect 2144 16453 2145 16487
rect 2179 16453 2180 16487
rect 2144 16419 2180 16453
rect 2144 16385 2145 16419
rect 2179 16385 2180 16419
rect 2144 16351 2180 16385
rect 2144 16317 2145 16351
rect 2179 16317 2180 16351
rect 2144 16283 2180 16317
rect 2144 16249 2145 16283
rect 2179 16249 2180 16283
rect 2144 16215 2180 16249
rect 2144 16181 2145 16215
rect 2179 16181 2180 16215
rect 2144 16147 2180 16181
rect 2144 16113 2145 16147
rect 2179 16113 2180 16147
rect 2144 16079 2180 16113
rect 2144 16045 2145 16079
rect 2179 16045 2180 16079
rect 256 15951 292 15985
rect 256 15917 257 15951
rect 291 15917 292 15951
rect 2144 16011 2180 16045
rect 2144 15977 2145 16011
rect 2179 15977 2180 16011
rect 256 15883 292 15917
rect 2144 15943 2180 15977
rect 2144 15909 2145 15943
rect 2179 15909 2180 15943
rect 256 15849 257 15883
rect 291 15849 292 15883
rect 256 15815 292 15849
rect 2144 15875 2180 15909
rect 2144 15841 2145 15875
rect 2179 15841 2180 15875
rect 256 15781 257 15815
rect 291 15781 292 15815
rect 256 15747 292 15781
rect 256 15713 257 15747
rect 291 15713 292 15747
rect 256 15679 292 15713
rect 256 15645 257 15679
rect 291 15645 292 15679
rect 256 15611 292 15645
rect 256 15577 257 15611
rect 291 15577 292 15611
rect 256 15543 292 15577
rect 256 15509 257 15543
rect 291 15509 292 15543
rect 256 15475 292 15509
rect 256 15441 257 15475
rect 291 15441 292 15475
rect 256 15407 292 15441
rect 256 15373 257 15407
rect 291 15373 292 15407
rect 256 15339 292 15373
rect 256 15305 257 15339
rect 291 15305 292 15339
rect 256 15271 292 15305
rect 256 15237 257 15271
rect 291 15237 292 15271
rect 256 15203 292 15237
rect 256 15169 257 15203
rect 291 15169 292 15203
rect 256 15135 292 15169
rect 256 15101 257 15135
rect 291 15101 292 15135
rect 256 15067 292 15101
rect 256 15033 257 15067
rect 291 15033 292 15067
rect 256 14999 292 15033
rect 256 14965 257 14999
rect 291 14965 292 14999
rect 256 14931 292 14965
rect 256 14897 257 14931
rect 291 14897 292 14931
rect 256 14863 292 14897
rect 256 14829 257 14863
rect 291 14829 292 14863
rect 256 14795 292 14829
rect 256 14761 257 14795
rect 291 14761 292 14795
rect 256 14727 292 14761
rect 256 14693 257 14727
rect 291 14693 292 14727
rect 256 14659 292 14693
rect 256 14625 257 14659
rect 291 14625 292 14659
rect 256 14591 292 14625
rect 256 14557 257 14591
rect 291 14557 292 14591
rect 256 14523 292 14557
rect 256 14489 257 14523
rect 291 14489 292 14523
rect 256 14455 292 14489
rect 256 14421 257 14455
rect 291 14421 292 14455
rect 256 14387 292 14421
rect 256 14353 257 14387
rect 291 14353 292 14387
rect 256 14319 292 14353
rect 256 14285 257 14319
rect 291 14285 292 14319
rect 256 14251 292 14285
rect 256 14217 257 14251
rect 291 14217 292 14251
rect 256 14183 292 14217
rect 256 14149 257 14183
rect 291 14149 292 14183
rect 256 14115 292 14149
rect 256 14081 257 14115
rect 291 14081 292 14115
rect 256 14047 292 14081
rect 256 14013 257 14047
rect 291 14013 292 14047
rect 256 13979 292 14013
rect 256 13945 257 13979
rect 291 13945 292 13979
rect 256 13911 292 13945
rect 256 13877 257 13911
rect 291 13877 292 13911
rect 256 13843 292 13877
rect 256 13809 257 13843
rect 291 13809 292 13843
rect 256 13775 292 13809
rect 256 13741 257 13775
rect 291 13741 292 13775
rect 256 13707 292 13741
rect 256 13673 257 13707
rect 291 13673 292 13707
rect 256 13639 292 13673
rect 256 13605 257 13639
rect 291 13605 292 13639
rect 256 13571 292 13605
rect 256 13537 257 13571
rect 291 13537 292 13571
rect 256 13503 292 13537
rect 256 13469 257 13503
rect 291 13469 292 13503
rect 256 13435 292 13469
rect 256 13401 257 13435
rect 291 13401 292 13435
rect 256 13367 292 13401
rect 256 13333 257 13367
rect 291 13333 292 13367
rect 256 13299 292 13333
rect 256 13265 257 13299
rect 291 13265 292 13299
rect 256 13231 292 13265
rect 256 13197 257 13231
rect 291 13197 292 13231
rect 256 13163 292 13197
rect 256 13129 257 13163
rect 291 13129 292 13163
rect 256 13095 292 13129
rect 256 13061 257 13095
rect 291 13061 292 13095
rect 256 13027 292 13061
rect 256 12993 257 13027
rect 291 12993 292 13027
rect 256 12959 292 12993
rect 256 12925 257 12959
rect 291 12925 292 12959
rect 256 12891 292 12925
rect 256 12857 257 12891
rect 291 12857 292 12891
rect 256 12823 292 12857
rect 256 12789 257 12823
rect 291 12789 292 12823
rect 256 12755 292 12789
rect 256 12721 257 12755
rect 291 12721 292 12755
rect 256 12687 292 12721
rect 256 12653 257 12687
rect 291 12653 292 12687
rect 256 12619 292 12653
rect 256 12585 257 12619
rect 291 12585 292 12619
rect 256 12551 292 12585
rect 256 12517 257 12551
rect 291 12517 292 12551
rect 256 12483 292 12517
rect 256 12449 257 12483
rect 291 12449 292 12483
rect 256 12415 292 12449
rect 256 12381 257 12415
rect 291 12381 292 12415
rect 256 12347 292 12381
rect 256 12313 257 12347
rect 291 12313 292 12347
rect 256 12279 292 12313
rect 256 12245 257 12279
rect 291 12245 292 12279
rect 256 12211 292 12245
rect 256 12177 257 12211
rect 291 12177 292 12211
rect 256 12143 292 12177
rect 256 12109 257 12143
rect 291 12109 292 12143
rect 2144 15807 2180 15841
rect 2144 15773 2145 15807
rect 2179 15773 2180 15807
rect 2144 15739 2180 15773
rect 2144 15705 2145 15739
rect 2179 15705 2180 15739
rect 2144 15671 2180 15705
rect 2144 15637 2145 15671
rect 2179 15637 2180 15671
rect 2144 15603 2180 15637
rect 2144 15569 2145 15603
rect 2179 15569 2180 15603
rect 2144 15535 2180 15569
rect 2144 15501 2145 15535
rect 2179 15501 2180 15535
rect 2144 15467 2180 15501
rect 2144 15433 2145 15467
rect 2179 15433 2180 15467
rect 2144 15399 2180 15433
rect 2144 15365 2145 15399
rect 2179 15365 2180 15399
rect 2144 15331 2180 15365
rect 2144 15297 2145 15331
rect 2179 15297 2180 15331
rect 2144 15263 2180 15297
rect 2144 15229 2145 15263
rect 2179 15229 2180 15263
rect 2144 15195 2180 15229
rect 2144 15161 2145 15195
rect 2179 15161 2180 15195
rect 2144 15127 2180 15161
rect 2144 15093 2145 15127
rect 2179 15093 2180 15127
rect 2144 15059 2180 15093
rect 2144 15025 2145 15059
rect 2179 15025 2180 15059
rect 2144 14991 2180 15025
rect 2144 14957 2145 14991
rect 2179 14957 2180 14991
rect 2144 14923 2180 14957
rect 2144 14889 2145 14923
rect 2179 14889 2180 14923
rect 2144 14855 2180 14889
rect 2144 14821 2145 14855
rect 2179 14821 2180 14855
rect 2144 14787 2180 14821
rect 2144 14753 2145 14787
rect 2179 14753 2180 14787
rect 2144 14719 2180 14753
rect 2144 14685 2145 14719
rect 2179 14685 2180 14719
rect 2144 14651 2180 14685
rect 2144 14617 2145 14651
rect 2179 14617 2180 14651
rect 2144 14583 2180 14617
rect 2144 14549 2145 14583
rect 2179 14549 2180 14583
rect 2144 14515 2180 14549
rect 2144 14481 2145 14515
rect 2179 14481 2180 14515
rect 2144 14447 2180 14481
rect 2144 14413 2145 14447
rect 2179 14413 2180 14447
rect 2144 14379 2180 14413
rect 2144 14345 2145 14379
rect 2179 14345 2180 14379
rect 2144 14311 2180 14345
rect 2144 14277 2145 14311
rect 2179 14277 2180 14311
rect 2144 14243 2180 14277
rect 2144 14209 2145 14243
rect 2179 14209 2180 14243
rect 2144 14175 2180 14209
rect 2144 14141 2145 14175
rect 2179 14141 2180 14175
rect 2144 14107 2180 14141
rect 2144 14073 2145 14107
rect 2179 14073 2180 14107
rect 2144 14039 2180 14073
rect 2144 14005 2145 14039
rect 2179 14005 2180 14039
rect 2144 13971 2180 14005
rect 2144 13937 2145 13971
rect 2179 13937 2180 13971
rect 2144 13903 2180 13937
rect 2144 13869 2145 13903
rect 2179 13869 2180 13903
rect 2144 13835 2180 13869
rect 2144 13801 2145 13835
rect 2179 13801 2180 13835
rect 2144 13767 2180 13801
rect 2144 13733 2145 13767
rect 2179 13733 2180 13767
rect 2144 13699 2180 13733
rect 2144 13665 2145 13699
rect 2179 13665 2180 13699
rect 2144 13631 2180 13665
rect 2144 13597 2145 13631
rect 2179 13597 2180 13631
rect 2144 13563 2180 13597
rect 2144 13529 2145 13563
rect 2179 13529 2180 13563
rect 2144 13495 2180 13529
rect 2144 13461 2145 13495
rect 2179 13461 2180 13495
rect 2144 13427 2180 13461
rect 2144 13393 2145 13427
rect 2179 13393 2180 13427
rect 2144 13359 2180 13393
rect 2144 13325 2145 13359
rect 2179 13325 2180 13359
rect 2144 13291 2180 13325
rect 2144 13257 2145 13291
rect 2179 13257 2180 13291
rect 2144 13223 2180 13257
rect 2144 13189 2145 13223
rect 2179 13189 2180 13223
rect 2144 13155 2180 13189
rect 2144 13121 2145 13155
rect 2179 13121 2180 13155
rect 2144 13087 2180 13121
rect 2144 13053 2145 13087
rect 2179 13053 2180 13087
rect 2144 13019 2180 13053
rect 2144 12985 2145 13019
rect 2179 12985 2180 13019
rect 2144 12951 2180 12985
rect 2144 12917 2145 12951
rect 2179 12917 2180 12951
rect 2144 12883 2180 12917
rect 2144 12849 2145 12883
rect 2179 12849 2180 12883
rect 2144 12815 2180 12849
rect 2144 12781 2145 12815
rect 2179 12781 2180 12815
rect 2144 12747 2180 12781
rect 2144 12713 2145 12747
rect 2179 12713 2180 12747
rect 2144 12679 2180 12713
rect 2144 12645 2145 12679
rect 2179 12645 2180 12679
rect 2144 12611 2180 12645
rect 2144 12577 2145 12611
rect 2179 12577 2180 12611
rect 2144 12543 2180 12577
rect 2144 12509 2145 12543
rect 2179 12509 2180 12543
rect 2144 12475 2180 12509
rect 2144 12441 2145 12475
rect 2179 12441 2180 12475
rect 2144 12407 2180 12441
rect 2144 12373 2145 12407
rect 2179 12373 2180 12407
rect 2144 12339 2180 12373
rect 2144 12305 2145 12339
rect 2179 12305 2180 12339
rect 2144 12271 2180 12305
rect 2144 12237 2145 12271
rect 2179 12237 2180 12271
rect 2144 12203 2180 12237
rect 2144 12169 2145 12203
rect 2179 12169 2180 12203
rect 2144 12135 2180 12169
rect 256 12075 292 12109
rect 256 12041 257 12075
rect 291 12041 292 12075
rect 2144 12101 2145 12135
rect 2179 12101 2180 12135
rect 2144 12067 2180 12101
rect 256 12007 292 12041
rect 256 11973 257 12007
rect 291 11973 292 12007
rect 2144 12033 2145 12067
rect 2179 12033 2180 12067
rect 2144 11999 2180 12033
rect 256 11939 292 11973
rect 256 11905 257 11939
rect 291 11905 292 11939
rect 2144 11965 2145 11999
rect 2179 11965 2180 11999
rect 2144 11931 2180 11965
rect 256 11871 292 11905
rect 256 11837 257 11871
rect 291 11837 292 11871
rect 256 11803 292 11837
rect 256 11769 257 11803
rect 291 11769 292 11803
rect 256 11735 292 11769
rect 256 11701 257 11735
rect 291 11701 292 11735
rect 256 11667 292 11701
rect 256 11633 257 11667
rect 291 11633 292 11667
rect 256 11599 292 11633
rect 256 11565 257 11599
rect 291 11565 292 11599
rect 256 11531 292 11565
rect 256 11497 257 11531
rect 291 11497 292 11531
rect 256 11463 292 11497
rect 256 11429 257 11463
rect 291 11429 292 11463
rect 256 11395 292 11429
rect 256 11361 257 11395
rect 291 11361 292 11395
rect 256 11327 292 11361
rect 256 11293 257 11327
rect 291 11293 292 11327
rect 256 11259 292 11293
rect 256 11225 257 11259
rect 291 11225 292 11259
rect 256 11191 292 11225
rect 256 11157 257 11191
rect 291 11157 292 11191
rect 256 11123 292 11157
rect 256 11089 257 11123
rect 291 11089 292 11123
rect 256 11055 292 11089
rect 256 11021 257 11055
rect 291 11021 292 11055
rect 256 10987 292 11021
rect 256 10953 257 10987
rect 291 10953 292 10987
rect 256 10919 292 10953
rect 256 10885 257 10919
rect 291 10885 292 10919
rect 256 10851 292 10885
rect 256 10817 257 10851
rect 291 10817 292 10851
rect 256 10783 292 10817
rect 256 10749 257 10783
rect 291 10749 292 10783
rect 256 10715 292 10749
rect 256 10681 257 10715
rect 291 10681 292 10715
rect 256 10647 292 10681
rect 256 10613 257 10647
rect 291 10613 292 10647
rect 256 10579 292 10613
rect 256 10545 257 10579
rect 291 10545 292 10579
rect 256 10511 292 10545
rect 256 10477 257 10511
rect 291 10477 292 10511
rect 256 10443 292 10477
rect 256 10409 257 10443
rect 291 10409 292 10443
rect 256 10375 292 10409
rect 256 10341 257 10375
rect 291 10341 292 10375
rect 256 10307 292 10341
rect 256 10273 257 10307
rect 291 10273 292 10307
rect 256 10239 292 10273
rect 256 10205 257 10239
rect 291 10205 292 10239
rect 256 10171 292 10205
rect 256 10137 257 10171
rect 291 10137 292 10171
rect 256 10103 292 10137
rect 256 10069 257 10103
rect 291 10069 292 10103
rect 256 10035 292 10069
rect 256 10001 257 10035
rect 291 10001 292 10035
rect 256 9967 292 10001
rect 256 9933 257 9967
rect 291 9933 292 9967
rect 256 9899 292 9933
rect 256 9865 257 9899
rect 291 9865 292 9899
rect 256 9831 292 9865
rect 256 9797 257 9831
rect 291 9797 292 9831
rect 256 9763 292 9797
rect 256 9729 257 9763
rect 291 9729 292 9763
rect 256 9695 292 9729
rect 256 9661 257 9695
rect 291 9661 292 9695
rect 256 9627 292 9661
rect 256 9593 257 9627
rect 291 9593 292 9627
rect 256 9559 292 9593
rect 256 9525 257 9559
rect 291 9525 292 9559
rect 256 9491 292 9525
rect 256 9457 257 9491
rect 291 9457 292 9491
rect 256 9423 292 9457
rect 256 9389 257 9423
rect 291 9389 292 9423
rect 256 9355 292 9389
rect 256 9321 257 9355
rect 291 9321 292 9355
rect 256 9287 292 9321
rect 256 9253 257 9287
rect 291 9253 292 9287
rect 256 9219 292 9253
rect 256 9185 257 9219
rect 291 9185 292 9219
rect 256 9151 292 9185
rect 256 9117 257 9151
rect 291 9117 292 9151
rect 256 9083 292 9117
rect 256 9049 257 9083
rect 291 9049 292 9083
rect 256 9015 292 9049
rect 256 8981 257 9015
rect 291 8981 292 9015
rect 256 8947 292 8981
rect 256 8913 257 8947
rect 291 8913 292 8947
rect 256 8879 292 8913
rect 256 8845 257 8879
rect 291 8845 292 8879
rect 256 8811 292 8845
rect 256 8777 257 8811
rect 291 8777 292 8811
rect 256 8743 292 8777
rect 256 8709 257 8743
rect 291 8709 292 8743
rect 256 8675 292 8709
rect 256 8641 257 8675
rect 291 8641 292 8675
rect 256 8607 292 8641
rect 256 8573 257 8607
rect 291 8573 292 8607
rect 256 8539 292 8573
rect 256 8505 257 8539
rect 291 8505 292 8539
rect 256 8471 292 8505
rect 256 8437 257 8471
rect 291 8437 292 8471
rect 256 8403 292 8437
rect 256 8369 257 8403
rect 291 8369 292 8403
rect 256 8335 292 8369
rect 256 8301 257 8335
rect 291 8301 292 8335
rect 256 8267 292 8301
rect 256 8233 257 8267
rect 291 8233 292 8267
rect 256 8199 292 8233
rect 2144 11897 2145 11931
rect 2179 11897 2180 11931
rect 2144 11863 2180 11897
rect 2144 11829 2145 11863
rect 2179 11829 2180 11863
rect 2144 11795 2180 11829
rect 2144 11761 2145 11795
rect 2179 11761 2180 11795
rect 2144 11727 2180 11761
rect 2144 11693 2145 11727
rect 2179 11693 2180 11727
rect 2144 11659 2180 11693
rect 2144 11625 2145 11659
rect 2179 11625 2180 11659
rect 2144 11591 2180 11625
rect 2144 11557 2145 11591
rect 2179 11557 2180 11591
rect 2144 11523 2180 11557
rect 2144 11489 2145 11523
rect 2179 11489 2180 11523
rect 2144 11455 2180 11489
rect 2144 11421 2145 11455
rect 2179 11421 2180 11455
rect 2144 11387 2180 11421
rect 2144 11353 2145 11387
rect 2179 11353 2180 11387
rect 2144 11319 2180 11353
rect 2144 11285 2145 11319
rect 2179 11285 2180 11319
rect 2144 11251 2180 11285
rect 2144 11217 2145 11251
rect 2179 11217 2180 11251
rect 2144 11183 2180 11217
rect 2144 11149 2145 11183
rect 2179 11149 2180 11183
rect 2144 11115 2180 11149
rect 2144 11081 2145 11115
rect 2179 11081 2180 11115
rect 2144 11047 2180 11081
rect 2144 11013 2145 11047
rect 2179 11013 2180 11047
rect 2144 10979 2180 11013
rect 2144 10945 2145 10979
rect 2179 10945 2180 10979
rect 2144 10911 2180 10945
rect 2144 10877 2145 10911
rect 2179 10877 2180 10911
rect 2144 10843 2180 10877
rect 2144 10809 2145 10843
rect 2179 10809 2180 10843
rect 2144 10775 2180 10809
rect 2144 10741 2145 10775
rect 2179 10741 2180 10775
rect 2144 10707 2180 10741
rect 2144 10673 2145 10707
rect 2179 10673 2180 10707
rect 2144 10639 2180 10673
rect 2144 10605 2145 10639
rect 2179 10605 2180 10639
rect 2144 10571 2180 10605
rect 2144 10537 2145 10571
rect 2179 10537 2180 10571
rect 2144 10503 2180 10537
rect 2144 10469 2145 10503
rect 2179 10469 2180 10503
rect 2144 10435 2180 10469
rect 2144 10401 2145 10435
rect 2179 10401 2180 10435
rect 2144 10367 2180 10401
rect 2144 10333 2145 10367
rect 2179 10333 2180 10367
rect 2144 10299 2180 10333
rect 2144 10265 2145 10299
rect 2179 10265 2180 10299
rect 2144 10231 2180 10265
rect 2144 10197 2145 10231
rect 2179 10197 2180 10231
rect 2144 10163 2180 10197
rect 2144 10129 2145 10163
rect 2179 10129 2180 10163
rect 2144 10095 2180 10129
rect 2144 10061 2145 10095
rect 2179 10061 2180 10095
rect 2144 10027 2180 10061
rect 2144 9993 2145 10027
rect 2179 9993 2180 10027
rect 2144 9959 2180 9993
rect 2144 9925 2145 9959
rect 2179 9925 2180 9959
rect 2144 9891 2180 9925
rect 2144 9857 2145 9891
rect 2179 9857 2180 9891
rect 2144 9823 2180 9857
rect 2144 9789 2145 9823
rect 2179 9789 2180 9823
rect 2144 9755 2180 9789
rect 2144 9721 2145 9755
rect 2179 9721 2180 9755
rect 2144 9687 2180 9721
rect 2144 9653 2145 9687
rect 2179 9653 2180 9687
rect 2144 9619 2180 9653
rect 2144 9585 2145 9619
rect 2179 9585 2180 9619
rect 2144 9551 2180 9585
rect 2144 9517 2145 9551
rect 2179 9517 2180 9551
rect 2144 9483 2180 9517
rect 2144 9449 2145 9483
rect 2179 9449 2180 9483
rect 2144 9415 2180 9449
rect 2144 9381 2145 9415
rect 2179 9381 2180 9415
rect 2144 9347 2180 9381
rect 2144 9313 2145 9347
rect 2179 9313 2180 9347
rect 2144 9279 2180 9313
rect 2144 9245 2145 9279
rect 2179 9245 2180 9279
rect 2144 9211 2180 9245
rect 2144 9177 2145 9211
rect 2179 9177 2180 9211
rect 2144 9143 2180 9177
rect 2144 9109 2145 9143
rect 2179 9109 2180 9143
rect 2144 9075 2180 9109
rect 2144 9041 2145 9075
rect 2179 9041 2180 9075
rect 2144 9007 2180 9041
rect 2144 8973 2145 9007
rect 2179 8973 2180 9007
rect 2144 8939 2180 8973
rect 2144 8905 2145 8939
rect 2179 8905 2180 8939
rect 2144 8871 2180 8905
rect 2144 8837 2145 8871
rect 2179 8837 2180 8871
rect 2144 8803 2180 8837
rect 2144 8769 2145 8803
rect 2179 8769 2180 8803
rect 2144 8735 2180 8769
rect 2144 8701 2145 8735
rect 2179 8701 2180 8735
rect 2144 8667 2180 8701
rect 2144 8633 2145 8667
rect 2179 8633 2180 8667
rect 2144 8599 2180 8633
rect 2144 8565 2145 8599
rect 2179 8565 2180 8599
rect 2144 8531 2180 8565
rect 2144 8497 2145 8531
rect 2179 8497 2180 8531
rect 2144 8463 2180 8497
rect 2144 8429 2145 8463
rect 2179 8429 2180 8463
rect 2144 8395 2180 8429
rect 2144 8361 2145 8395
rect 2179 8361 2180 8395
rect 2144 8327 2180 8361
rect 2144 8293 2145 8327
rect 2179 8293 2180 8327
rect 2144 8259 2180 8293
rect 2144 8225 2145 8259
rect 2179 8225 2180 8259
rect 256 8165 257 8199
rect 291 8165 292 8199
rect 256 8131 292 8165
rect 256 8097 257 8131
rect 291 8097 292 8131
rect 256 8063 292 8097
rect 256 8029 257 8063
rect 291 8029 292 8063
rect 256 7995 292 8029
rect 256 7961 257 7995
rect 291 7961 292 7995
rect 256 7927 292 7961
rect 256 7893 257 7927
rect 291 7893 292 7927
rect 256 7859 292 7893
rect 256 7825 257 7859
rect 291 7825 292 7859
rect 256 7791 292 7825
rect 256 7757 257 7791
rect 291 7757 292 7791
rect 256 7723 292 7757
rect 256 7689 257 7723
rect 291 7689 292 7723
rect 256 7655 292 7689
rect 256 7621 257 7655
rect 291 7621 292 7655
rect 256 7587 292 7621
rect 256 7553 257 7587
rect 291 7553 292 7587
rect 256 7519 292 7553
rect 256 7485 257 7519
rect 291 7485 292 7519
rect 256 7451 292 7485
rect 256 7417 257 7451
rect 291 7417 292 7451
rect 256 7383 292 7417
rect 256 7349 257 7383
rect 291 7349 292 7383
rect 256 7315 292 7349
rect 256 7281 257 7315
rect 291 7281 292 7315
rect 256 7247 292 7281
rect 256 7213 257 7247
rect 291 7213 292 7247
rect 256 7179 292 7213
rect 256 7145 257 7179
rect 291 7145 292 7179
rect 256 7111 292 7145
rect 256 7077 257 7111
rect 291 7077 292 7111
rect 256 7043 292 7077
rect 256 7009 257 7043
rect 291 7009 292 7043
rect 256 6975 292 7009
rect 256 6941 257 6975
rect 291 6941 292 6975
rect 256 6907 292 6941
rect 256 6873 257 6907
rect 291 6873 292 6907
rect 256 6790 292 6873
rect 231 6766 292 6790
rect 265 6732 292 6766
rect 231 6694 292 6732
rect 265 6660 292 6694
rect 231 6623 292 6660
rect 265 6589 292 6623
rect 231 6552 292 6589
rect 265 6518 292 6552
rect 231 6481 292 6518
rect 265 6447 292 6481
rect 231 6410 292 6447
rect 265 6376 292 6410
rect 231 6339 292 6376
rect 265 6305 292 6339
rect 231 6268 292 6305
rect 265 6234 292 6268
rect 231 6197 292 6234
rect 265 6163 292 6197
rect 231 6126 292 6163
rect 265 6092 292 6126
rect 231 6055 292 6092
rect 265 6021 292 6055
rect 231 5984 292 6021
rect 265 5950 292 5984
rect 231 5913 292 5950
rect 265 5879 292 5913
rect 231 5842 292 5879
rect 265 5808 292 5842
rect 231 5706 292 5808
rect 231 5672 253 5706
rect 287 5672 292 5706
rect 231 5638 292 5672
rect 231 5604 253 5638
rect 287 5604 292 5638
rect 231 5570 292 5604
rect 231 5536 253 5570
rect 287 5536 292 5570
rect 231 5502 292 5536
rect 2144 8191 2180 8225
rect 2144 8157 2145 8191
rect 2179 8157 2180 8191
rect 2144 8123 2180 8157
rect 2144 8089 2145 8123
rect 2179 8089 2180 8123
rect 2144 8055 2180 8089
rect 2144 8021 2145 8055
rect 2179 8021 2180 8055
rect 2144 7987 2180 8021
rect 2144 7953 2145 7987
rect 2179 7953 2180 7987
rect 2144 7919 2180 7953
rect 2144 7885 2145 7919
rect 2179 7885 2180 7919
rect 2144 7851 2180 7885
rect 2144 7817 2145 7851
rect 2179 7817 2180 7851
rect 2144 7783 2180 7817
rect 2144 7749 2145 7783
rect 2179 7749 2180 7783
rect 2144 7715 2180 7749
rect 2144 7681 2145 7715
rect 2179 7681 2180 7715
rect 2144 7647 2180 7681
rect 2144 7613 2145 7647
rect 2179 7613 2180 7647
rect 2144 7579 2180 7613
rect 2144 7545 2145 7579
rect 2179 7545 2180 7579
rect 2144 7511 2180 7545
rect 2144 7477 2145 7511
rect 2179 7477 2180 7511
rect 2144 7443 2180 7477
rect 2144 7409 2145 7443
rect 2179 7409 2180 7443
rect 2144 7375 2180 7409
rect 2144 7341 2145 7375
rect 2179 7341 2180 7375
rect 2144 7307 2180 7341
rect 2144 7273 2145 7307
rect 2179 7273 2180 7307
rect 2144 7239 2180 7273
rect 2144 7205 2145 7239
rect 2179 7205 2180 7239
rect 2144 7171 2180 7205
rect 2144 7137 2145 7171
rect 2179 7137 2180 7171
rect 2144 7103 2180 7137
rect 2144 7069 2145 7103
rect 2179 7069 2180 7103
rect 2144 7035 2180 7069
rect 2144 7001 2145 7035
rect 2179 7001 2180 7035
rect 2144 6967 2180 7001
rect 2144 6933 2145 6967
rect 2179 6933 2180 6967
rect 2144 6899 2180 6933
rect 2144 6865 2145 6899
rect 2179 6865 2180 6899
rect 2144 6831 2180 6865
rect 2144 6797 2145 6831
rect 2179 6797 2180 6831
rect 2144 6763 2180 6797
rect 2144 6729 2145 6763
rect 2179 6729 2180 6763
rect 2144 6695 2180 6729
rect 2144 6661 2145 6695
rect 2179 6661 2180 6695
rect 2144 6627 2180 6661
rect 2144 6593 2145 6627
rect 2179 6593 2180 6627
rect 2144 6559 2180 6593
rect 2144 6525 2145 6559
rect 2179 6525 2180 6559
rect 2144 6491 2180 6525
rect 2144 6457 2145 6491
rect 2179 6457 2180 6491
rect 2144 6423 2180 6457
rect 2144 6389 2145 6423
rect 2179 6389 2180 6423
rect 2144 6355 2180 6389
rect 2144 6321 2145 6355
rect 2179 6321 2180 6355
rect 2144 6287 2180 6321
rect 2144 6253 2145 6287
rect 2179 6253 2180 6287
rect 2144 6219 2180 6253
rect 2144 6185 2145 6219
rect 2179 6185 2180 6219
rect 2144 6151 2180 6185
rect 2144 6117 2145 6151
rect 2179 6117 2180 6151
rect 2144 6083 2180 6117
rect 2144 6049 2145 6083
rect 2179 6049 2180 6083
rect 2742 10889 6700 10890
rect 2742 10856 2835 10889
rect 2742 10822 2743 10856
rect 2777 10855 2835 10856
rect 2869 10855 2903 10889
rect 2937 10855 2971 10889
rect 3005 10855 3039 10889
rect 3073 10855 3107 10889
rect 3141 10855 3175 10889
rect 3209 10855 3243 10889
rect 3277 10855 3311 10889
rect 3345 10855 3379 10889
rect 3413 10855 3447 10889
rect 3481 10855 3515 10889
rect 3549 10855 3583 10889
rect 3617 10855 3651 10889
rect 3685 10855 3719 10889
rect 3753 10855 3787 10889
rect 3821 10855 3855 10889
rect 3889 10855 3923 10889
rect 3957 10855 3991 10889
rect 4025 10855 4059 10889
rect 4093 10855 4127 10889
rect 4161 10855 4195 10889
rect 4229 10855 4263 10889
rect 4297 10855 4331 10889
rect 4365 10855 4399 10889
rect 4433 10855 4467 10889
rect 4501 10855 4535 10889
rect 4569 10855 4603 10889
rect 4637 10855 4671 10889
rect 4705 10855 4799 10889
rect 4833 10855 4867 10889
rect 4901 10855 4935 10889
rect 4969 10855 5003 10889
rect 5037 10855 5071 10889
rect 5105 10855 5139 10889
rect 5173 10855 5207 10889
rect 5241 10855 5275 10889
rect 5309 10855 5343 10889
rect 5377 10855 5411 10889
rect 5445 10855 5479 10889
rect 5513 10855 5547 10889
rect 5581 10855 5615 10889
rect 5649 10855 5683 10889
rect 5717 10855 5751 10889
rect 5785 10855 5819 10889
rect 5853 10855 5887 10889
rect 5921 10855 5955 10889
rect 5989 10855 6023 10889
rect 6057 10855 6091 10889
rect 6125 10855 6159 10889
rect 6193 10855 6227 10889
rect 6261 10855 6295 10889
rect 6329 10855 6363 10889
rect 6397 10855 6431 10889
rect 6465 10855 6499 10889
rect 6533 10855 6567 10889
rect 6601 10856 6700 10889
rect 6601 10855 6665 10856
rect 2777 10854 6665 10855
rect 2777 10822 2778 10854
rect 2742 10788 2778 10822
rect 2742 10754 2743 10788
rect 2777 10754 2778 10788
rect 2742 10720 2778 10754
rect 4703 10776 4739 10854
rect 6664 10822 6665 10854
rect 6699 10822 6700 10856
rect 2742 10686 2743 10720
rect 2777 10686 2778 10720
rect 2742 10652 2778 10686
rect 2742 10618 2743 10652
rect 2777 10618 2778 10652
rect 2742 10584 2778 10618
rect 2742 10550 2743 10584
rect 2777 10550 2778 10584
rect 2742 10516 2778 10550
rect 2742 10482 2743 10516
rect 2777 10482 2778 10516
rect 2742 10448 2778 10482
rect 2742 10414 2743 10448
rect 2777 10414 2778 10448
rect 2742 10380 2778 10414
rect 2742 10346 2743 10380
rect 2777 10346 2778 10380
rect 2742 10312 2778 10346
rect 2742 10278 2743 10312
rect 2777 10278 2778 10312
rect 2742 10244 2778 10278
rect 2742 10210 2743 10244
rect 2777 10210 2778 10244
rect 2742 10176 2778 10210
rect 2742 10142 2743 10176
rect 2777 10142 2778 10176
rect 2742 10108 2778 10142
rect 2742 10074 2743 10108
rect 2777 10074 2778 10108
rect 2742 10040 2778 10074
rect 2742 10006 2743 10040
rect 2777 10006 2778 10040
rect 2742 9972 2778 10006
rect 2742 9938 2743 9972
rect 2777 9938 2778 9972
rect 2742 9904 2778 9938
rect 2742 9870 2743 9904
rect 2777 9870 2778 9904
rect 2742 9836 2778 9870
rect 2742 9802 2743 9836
rect 2777 9802 2778 9836
rect 2742 9768 2778 9802
rect 2742 9734 2743 9768
rect 2777 9734 2778 9768
rect 2742 9700 2778 9734
rect 2742 9666 2743 9700
rect 2777 9666 2778 9700
rect 2742 9632 2778 9666
rect 2742 9598 2743 9632
rect 2777 9598 2778 9632
rect 2742 9564 2778 9598
rect 2742 9530 2743 9564
rect 2777 9530 2778 9564
rect 2742 9496 2778 9530
rect 2742 9462 2743 9496
rect 2777 9462 2778 9496
rect 2742 9428 2778 9462
rect 2742 9394 2743 9428
rect 2777 9394 2778 9428
rect 2742 9360 2778 9394
rect 2742 9326 2743 9360
rect 2777 9326 2778 9360
rect 2742 9292 2778 9326
rect 2742 9258 2743 9292
rect 2777 9258 2778 9292
rect 2742 9224 2778 9258
rect 2742 9190 2743 9224
rect 2777 9190 2778 9224
rect 2742 9156 2778 9190
rect 2742 9122 2743 9156
rect 2777 9122 2778 9156
rect 2742 9088 2778 9122
rect 2742 9054 2743 9088
rect 2777 9054 2778 9088
rect 2742 9020 2778 9054
rect 2742 8986 2743 9020
rect 2777 8986 2778 9020
rect 2742 8952 2778 8986
rect 2742 8918 2743 8952
rect 2777 8918 2778 8952
rect 2742 8884 2778 8918
rect 2742 8850 2743 8884
rect 2777 8850 2778 8884
rect 2742 8816 2778 8850
rect 2742 8782 2743 8816
rect 2777 8782 2778 8816
rect 2742 8748 2778 8782
rect 2742 8714 2743 8748
rect 2777 8714 2778 8748
rect 2742 8680 2778 8714
rect 2742 8646 2743 8680
rect 2777 8646 2778 8680
rect 2742 8612 2778 8646
rect 2742 8578 2743 8612
rect 2777 8578 2778 8612
rect 2742 8544 2778 8578
rect 2742 8510 2743 8544
rect 2777 8510 2778 8544
rect 2742 8476 2778 8510
rect 2742 8442 2743 8476
rect 2777 8442 2778 8476
rect 2742 8408 2778 8442
rect 2742 8374 2743 8408
rect 2777 8374 2778 8408
rect 2742 8340 2778 8374
rect 2742 8306 2743 8340
rect 2777 8306 2778 8340
rect 2742 8272 2778 8306
rect 2742 8238 2743 8272
rect 2777 8238 2778 8272
rect 2742 8204 2778 8238
rect 2742 8170 2743 8204
rect 2777 8170 2778 8204
rect 2742 8136 2778 8170
rect 2742 8102 2743 8136
rect 2777 8102 2778 8136
rect 2742 8068 2778 8102
rect 2742 8034 2743 8068
rect 2777 8034 2778 8068
rect 2742 8000 2778 8034
rect 2742 7966 2743 8000
rect 2777 7966 2778 8000
rect 2742 7932 2778 7966
rect 2742 7898 2743 7932
rect 2777 7898 2778 7932
rect 2742 7864 2778 7898
rect 2742 7830 2743 7864
rect 2777 7830 2778 7864
rect 2742 7796 2778 7830
rect 2742 7762 2743 7796
rect 2777 7762 2778 7796
rect 2742 7728 2778 7762
rect 2742 7694 2743 7728
rect 2777 7694 2778 7728
rect 2742 7660 2778 7694
rect 2742 7626 2743 7660
rect 2777 7626 2778 7660
rect 2742 7592 2778 7626
rect 2742 7558 2743 7592
rect 2777 7558 2778 7592
rect 2742 7524 2778 7558
rect 2742 7490 2743 7524
rect 2777 7490 2778 7524
rect 2742 7456 2778 7490
rect 2742 7422 2743 7456
rect 2777 7422 2778 7456
rect 2742 7388 2778 7422
rect 2742 7354 2743 7388
rect 2777 7354 2778 7388
rect 2742 7320 2778 7354
rect 2742 7286 2743 7320
rect 2777 7286 2778 7320
rect 2742 7252 2778 7286
rect 2742 7218 2743 7252
rect 2777 7218 2778 7252
rect 2742 7184 2778 7218
rect 2742 7150 2743 7184
rect 2777 7150 2778 7184
rect 2742 7116 2778 7150
rect 2742 7082 2743 7116
rect 2777 7082 2778 7116
rect 2742 7048 2778 7082
rect 2742 7014 2743 7048
rect 2777 7014 2778 7048
rect 2742 6980 2778 7014
rect 2742 6946 2743 6980
rect 2777 6946 2778 6980
rect 2742 6912 2778 6946
rect 2742 6878 2743 6912
rect 2777 6878 2778 6912
rect 2742 6844 2778 6878
rect 2742 6810 2743 6844
rect 2777 6810 2778 6844
rect 2742 6776 2778 6810
rect 2742 6742 2743 6776
rect 2777 6742 2778 6776
rect 2742 6708 2778 6742
rect 2742 6674 2743 6708
rect 2777 6674 2778 6708
rect 2742 6640 2778 6674
rect 2742 6606 2743 6640
rect 2777 6606 2778 6640
rect 2742 6572 2778 6606
rect 2742 6538 2743 6572
rect 2777 6538 2778 6572
rect 4703 10742 4704 10776
rect 4738 10742 4739 10776
rect 6664 10788 6700 10822
rect 6664 10754 6665 10788
rect 6699 10754 6700 10788
rect 4703 10708 4739 10742
rect 4703 10674 4704 10708
rect 4738 10674 4739 10708
rect 4703 10640 4739 10674
rect 4703 10606 4704 10640
rect 4738 10606 4739 10640
rect 4703 10572 4739 10606
rect 4703 10538 4704 10572
rect 4738 10538 4739 10572
rect 4703 10504 4739 10538
rect 4703 10470 4704 10504
rect 4738 10470 4739 10504
rect 4703 10436 4739 10470
rect 4703 10402 4704 10436
rect 4738 10402 4739 10436
rect 4703 10368 4739 10402
rect 4703 10334 4704 10368
rect 4738 10334 4739 10368
rect 4703 10300 4739 10334
rect 4703 10266 4704 10300
rect 4738 10266 4739 10300
rect 4703 10232 4739 10266
rect 4703 10198 4704 10232
rect 4738 10198 4739 10232
rect 4703 10164 4739 10198
rect 4703 10130 4704 10164
rect 4738 10130 4739 10164
rect 4703 10096 4739 10130
rect 4703 10062 4704 10096
rect 4738 10062 4739 10096
rect 4703 10028 4739 10062
rect 4703 9994 4704 10028
rect 4738 9994 4739 10028
rect 4703 9960 4739 9994
rect 4703 9926 4704 9960
rect 4738 9926 4739 9960
rect 4703 9892 4739 9926
rect 4703 9858 4704 9892
rect 4738 9858 4739 9892
rect 4703 9824 4739 9858
rect 4703 9790 4704 9824
rect 4738 9790 4739 9824
rect 4703 9756 4739 9790
rect 4703 9722 4704 9756
rect 4738 9722 4739 9756
rect 4703 9688 4739 9722
rect 4703 9654 4704 9688
rect 4738 9654 4739 9688
rect 4703 9620 4739 9654
rect 4703 9586 4704 9620
rect 4738 9586 4739 9620
rect 4703 9552 4739 9586
rect 4703 9518 4704 9552
rect 4738 9518 4739 9552
rect 4703 9484 4739 9518
rect 4703 9450 4704 9484
rect 4738 9450 4739 9484
rect 4703 9416 4739 9450
rect 4703 9382 4704 9416
rect 4738 9382 4739 9416
rect 4703 9348 4739 9382
rect 4703 9314 4704 9348
rect 4738 9314 4739 9348
rect 4703 9280 4739 9314
rect 4703 9246 4704 9280
rect 4738 9246 4739 9280
rect 4703 9212 4739 9246
rect 4703 9178 4704 9212
rect 4738 9178 4739 9212
rect 4703 9144 4739 9178
rect 4703 9110 4704 9144
rect 4738 9110 4739 9144
rect 4703 9076 4739 9110
rect 4703 9042 4704 9076
rect 4738 9042 4739 9076
rect 4703 9008 4739 9042
rect 4703 8974 4704 9008
rect 4738 8974 4739 9008
rect 4703 8940 4739 8974
rect 4703 8906 4704 8940
rect 4738 8906 4739 8940
rect 4703 8872 4739 8906
rect 4703 8838 4704 8872
rect 4738 8838 4739 8872
rect 4703 8804 4739 8838
rect 4703 8770 4704 8804
rect 4738 8770 4739 8804
rect 4703 8736 4739 8770
rect 4703 8702 4704 8736
rect 4738 8702 4739 8736
rect 4703 8668 4739 8702
rect 4703 8634 4704 8668
rect 4738 8634 4739 8668
rect 4703 8600 4739 8634
rect 4703 8566 4704 8600
rect 4738 8566 4739 8600
rect 4703 8532 4739 8566
rect 4703 8498 4704 8532
rect 4738 8498 4739 8532
rect 4703 8464 4739 8498
rect 4703 8430 4704 8464
rect 4738 8430 4739 8464
rect 4703 8396 4739 8430
rect 4703 8362 4704 8396
rect 4738 8362 4739 8396
rect 4703 8328 4739 8362
rect 4703 8294 4704 8328
rect 4738 8294 4739 8328
rect 4703 8260 4739 8294
rect 4703 8226 4704 8260
rect 4738 8226 4739 8260
rect 4703 8192 4739 8226
rect 4703 8158 4704 8192
rect 4738 8158 4739 8192
rect 4703 8124 4739 8158
rect 4703 8090 4704 8124
rect 4738 8090 4739 8124
rect 4703 8056 4739 8090
rect 4703 8022 4704 8056
rect 4738 8022 4739 8056
rect 4703 7988 4739 8022
rect 4703 7954 4704 7988
rect 4738 7954 4739 7988
rect 4703 7920 4739 7954
rect 4703 7886 4704 7920
rect 4738 7886 4739 7920
rect 4703 7852 4739 7886
rect 4703 7818 4704 7852
rect 4738 7818 4739 7852
rect 4703 7784 4739 7818
rect 4703 7750 4704 7784
rect 4738 7750 4739 7784
rect 4703 7716 4739 7750
rect 4703 7682 4704 7716
rect 4738 7682 4739 7716
rect 4703 7648 4739 7682
rect 4703 7614 4704 7648
rect 4738 7614 4739 7648
rect 4703 7580 4739 7614
rect 4703 7546 4704 7580
rect 4738 7546 4739 7580
rect 4703 7512 4739 7546
rect 4703 7478 4704 7512
rect 4738 7478 4739 7512
rect 4703 7444 4739 7478
rect 4703 7410 4704 7444
rect 4738 7410 4739 7444
rect 4703 7376 4739 7410
rect 4703 7342 4704 7376
rect 4738 7342 4739 7376
rect 4703 7308 4739 7342
rect 4703 7274 4704 7308
rect 4738 7274 4739 7308
rect 4703 7240 4739 7274
rect 4703 7206 4704 7240
rect 4738 7206 4739 7240
rect 4703 7172 4739 7206
rect 4703 7138 4704 7172
rect 4738 7138 4739 7172
rect 4703 7104 4739 7138
rect 4703 7070 4704 7104
rect 4738 7070 4739 7104
rect 4703 7036 4739 7070
rect 4703 7002 4704 7036
rect 4738 7002 4739 7036
rect 4703 6968 4739 7002
rect 4703 6934 4704 6968
rect 4738 6934 4739 6968
rect 4703 6900 4739 6934
rect 4703 6866 4704 6900
rect 4738 6866 4739 6900
rect 4703 6832 4739 6866
rect 4703 6798 4704 6832
rect 4738 6798 4739 6832
rect 4703 6764 4739 6798
rect 4703 6730 4704 6764
rect 4738 6730 4739 6764
rect 4703 6696 4739 6730
rect 4703 6662 4704 6696
rect 4738 6662 4739 6696
rect 4703 6628 4739 6662
rect 4703 6594 4704 6628
rect 4738 6594 4739 6628
rect 2742 6460 2778 6538
rect 4703 6560 4739 6594
rect 6664 10720 6700 10754
rect 6664 10686 6665 10720
rect 6699 10686 6700 10720
rect 6664 10652 6700 10686
rect 6664 10618 6665 10652
rect 6699 10618 6700 10652
rect 6664 10584 6700 10618
rect 6664 10550 6665 10584
rect 6699 10550 6700 10584
rect 6664 10516 6700 10550
rect 6664 10482 6665 10516
rect 6699 10482 6700 10516
rect 6664 10448 6700 10482
rect 6664 10414 6665 10448
rect 6699 10414 6700 10448
rect 6664 10380 6700 10414
rect 6664 10346 6665 10380
rect 6699 10346 6700 10380
rect 6664 10312 6700 10346
rect 6664 10278 6665 10312
rect 6699 10278 6700 10312
rect 6664 10244 6700 10278
rect 6664 10210 6665 10244
rect 6699 10210 6700 10244
rect 6664 10176 6700 10210
rect 6664 10142 6665 10176
rect 6699 10142 6700 10176
rect 6664 10108 6700 10142
rect 6664 10074 6665 10108
rect 6699 10074 6700 10108
rect 6664 10040 6700 10074
rect 6664 10006 6665 10040
rect 6699 10006 6700 10040
rect 6664 9972 6700 10006
rect 6664 9938 6665 9972
rect 6699 9938 6700 9972
rect 6664 9904 6700 9938
rect 6664 9870 6665 9904
rect 6699 9870 6700 9904
rect 6664 9836 6700 9870
rect 6664 9802 6665 9836
rect 6699 9802 6700 9836
rect 6664 9768 6700 9802
rect 6664 9734 6665 9768
rect 6699 9734 6700 9768
rect 6664 9700 6700 9734
rect 6664 9666 6665 9700
rect 6699 9666 6700 9700
rect 6664 9632 6700 9666
rect 6664 9598 6665 9632
rect 6699 9598 6700 9632
rect 6664 9564 6700 9598
rect 6664 9530 6665 9564
rect 6699 9530 6700 9564
rect 6664 9496 6700 9530
rect 6664 9462 6665 9496
rect 6699 9462 6700 9496
rect 6664 9428 6700 9462
rect 6664 9394 6665 9428
rect 6699 9394 6700 9428
rect 6664 9360 6700 9394
rect 6664 9326 6665 9360
rect 6699 9326 6700 9360
rect 6664 9292 6700 9326
rect 6664 9258 6665 9292
rect 6699 9258 6700 9292
rect 6664 9224 6700 9258
rect 6664 9190 6665 9224
rect 6699 9190 6700 9224
rect 6664 9156 6700 9190
rect 6664 9122 6665 9156
rect 6699 9122 6700 9156
rect 6664 9088 6700 9122
rect 6664 9054 6665 9088
rect 6699 9054 6700 9088
rect 6664 9020 6700 9054
rect 6664 8986 6665 9020
rect 6699 8986 6700 9020
rect 6664 8952 6700 8986
rect 6664 8918 6665 8952
rect 6699 8918 6700 8952
rect 6664 8884 6700 8918
rect 6664 8850 6665 8884
rect 6699 8850 6700 8884
rect 6664 8816 6700 8850
rect 6664 8782 6665 8816
rect 6699 8782 6700 8816
rect 6664 8748 6700 8782
rect 6664 8714 6665 8748
rect 6699 8714 6700 8748
rect 6664 8680 6700 8714
rect 6664 8646 6665 8680
rect 6699 8646 6700 8680
rect 6664 8612 6700 8646
rect 6664 8578 6665 8612
rect 6699 8578 6700 8612
rect 6664 8544 6700 8578
rect 6664 8510 6665 8544
rect 6699 8510 6700 8544
rect 6664 8476 6700 8510
rect 6664 8442 6665 8476
rect 6699 8442 6700 8476
rect 6664 8408 6700 8442
rect 6664 8374 6665 8408
rect 6699 8374 6700 8408
rect 6664 8340 6700 8374
rect 6664 8306 6665 8340
rect 6699 8306 6700 8340
rect 6664 8272 6700 8306
rect 6664 8238 6665 8272
rect 6699 8238 6700 8272
rect 6664 8204 6700 8238
rect 6664 8170 6665 8204
rect 6699 8170 6700 8204
rect 6664 8136 6700 8170
rect 6664 8102 6665 8136
rect 6699 8102 6700 8136
rect 6664 8068 6700 8102
rect 6664 8034 6665 8068
rect 6699 8034 6700 8068
rect 6664 8000 6700 8034
rect 6664 7966 6665 8000
rect 6699 7966 6700 8000
rect 6664 7932 6700 7966
rect 6664 7898 6665 7932
rect 6699 7898 6700 7932
rect 6664 7864 6700 7898
rect 6664 7830 6665 7864
rect 6699 7830 6700 7864
rect 6664 7796 6700 7830
rect 6664 7762 6665 7796
rect 6699 7762 6700 7796
rect 6664 7728 6700 7762
rect 6664 7694 6665 7728
rect 6699 7694 6700 7728
rect 6664 7660 6700 7694
rect 6664 7626 6665 7660
rect 6699 7626 6700 7660
rect 6664 7592 6700 7626
rect 6664 7558 6665 7592
rect 6699 7558 6700 7592
rect 6664 7524 6700 7558
rect 6664 7490 6665 7524
rect 6699 7490 6700 7524
rect 6664 7456 6700 7490
rect 6664 7422 6665 7456
rect 6699 7422 6700 7456
rect 6664 7388 6700 7422
rect 6664 7354 6665 7388
rect 6699 7354 6700 7388
rect 6664 7320 6700 7354
rect 6664 7286 6665 7320
rect 6699 7286 6700 7320
rect 6664 7252 6700 7286
rect 6664 7218 6665 7252
rect 6699 7218 6700 7252
rect 6664 7184 6700 7218
rect 6664 7150 6665 7184
rect 6699 7150 6700 7184
rect 6664 7116 6700 7150
rect 6664 7082 6665 7116
rect 6699 7082 6700 7116
rect 6664 7048 6700 7082
rect 6664 7014 6665 7048
rect 6699 7014 6700 7048
rect 6664 6980 6700 7014
rect 6664 6946 6665 6980
rect 6699 6946 6700 6980
rect 6664 6912 6700 6946
rect 6664 6878 6665 6912
rect 6699 6878 6700 6912
rect 6664 6844 6700 6878
rect 6664 6810 6665 6844
rect 6699 6810 6700 6844
rect 6664 6776 6700 6810
rect 6664 6742 6665 6776
rect 6699 6742 6700 6776
rect 6664 6708 6700 6742
rect 6664 6674 6665 6708
rect 6699 6674 6700 6708
rect 6664 6640 6700 6674
rect 6664 6606 6665 6640
rect 6699 6606 6700 6640
rect 6664 6572 6700 6606
rect 4703 6526 4704 6560
rect 4738 6526 4739 6560
rect 4703 6492 4739 6526
rect 4703 6460 4704 6492
rect 2742 6459 4704 6460
rect 2742 6425 2776 6459
rect 2810 6425 2844 6459
rect 2878 6425 2912 6459
rect 2946 6425 2980 6459
rect 3014 6425 3048 6459
rect 3082 6425 3116 6459
rect 3150 6425 3184 6459
rect 3218 6425 3252 6459
rect 3286 6425 3320 6459
rect 3354 6425 3388 6459
rect 3422 6425 3456 6459
rect 3490 6425 3524 6459
rect 3558 6425 3592 6459
rect 3626 6425 3660 6459
rect 3694 6425 3728 6459
rect 3762 6425 3796 6459
rect 3830 6425 3864 6459
rect 3898 6425 3932 6459
rect 3966 6425 4000 6459
rect 4034 6425 4068 6459
rect 4102 6425 4136 6459
rect 4170 6425 4204 6459
rect 4238 6425 4272 6459
rect 4306 6425 4340 6459
rect 4374 6425 4408 6459
rect 4442 6425 4476 6459
rect 4510 6425 4544 6459
rect 4578 6425 4612 6459
rect 4646 6458 4704 6459
rect 4738 6460 4739 6492
rect 6664 6538 6665 6572
rect 6699 6538 6700 6572
rect 6664 6460 6700 6538
rect 4738 6459 6700 6460
rect 4738 6458 4796 6459
rect 4646 6425 4796 6458
rect 4830 6425 4864 6459
rect 4898 6425 4932 6459
rect 4966 6425 5000 6459
rect 5034 6425 5068 6459
rect 5102 6425 5136 6459
rect 5170 6425 5204 6459
rect 5238 6425 5272 6459
rect 5306 6425 5340 6459
rect 5374 6425 5408 6459
rect 5442 6425 5476 6459
rect 5510 6425 5544 6459
rect 5578 6425 5612 6459
rect 5646 6425 5680 6459
rect 5714 6425 5748 6459
rect 5782 6425 5816 6459
rect 5850 6425 5884 6459
rect 5918 6425 5952 6459
rect 5986 6425 6020 6459
rect 6054 6425 6088 6459
rect 6122 6425 6156 6459
rect 6190 6425 6224 6459
rect 6258 6425 6292 6459
rect 6326 6425 6360 6459
rect 6394 6425 6428 6459
rect 6462 6425 6496 6459
rect 6530 6425 6564 6459
rect 6598 6425 6632 6459
rect 6666 6425 6700 6459
rect 2742 6424 6700 6425
rect 2144 6015 2180 6049
rect 2144 5981 2145 6015
rect 2179 5981 2180 6015
rect 2144 5947 2180 5981
rect 2144 5913 2145 5947
rect 2179 5913 2180 5947
rect 2144 5879 2180 5913
rect 2144 5845 2145 5879
rect 2179 5845 2180 5879
rect 2144 5811 2180 5845
rect 2144 5777 2145 5811
rect 2179 5777 2180 5811
rect 2144 5743 2180 5777
rect 2144 5709 2145 5743
rect 2179 5709 2180 5743
rect 2144 5675 2180 5709
rect 2144 5641 2145 5675
rect 2179 5641 2180 5675
rect 2144 5607 2180 5641
rect 2144 5573 2145 5607
rect 2179 5575 2180 5607
rect 3530 5575 5656 5576
rect 2179 5574 3188 5575
rect 2179 5573 2280 5574
rect 2144 5540 2280 5573
rect 2314 5540 2576 5574
rect 2610 5540 2644 5574
rect 2678 5540 2712 5574
rect 2746 5540 2780 5574
rect 2814 5540 2848 5574
rect 2882 5540 2916 5574
rect 2950 5540 2984 5574
rect 3018 5540 3052 5574
rect 3086 5540 3120 5574
rect 3154 5540 3188 5574
rect 2144 5539 3188 5540
rect 231 5468 253 5502
rect 287 5468 292 5502
rect 231 5402 292 5468
rect 3152 5492 3188 5539
rect 265 5368 292 5402
rect 3152 5458 3153 5492
rect 3187 5458 3188 5492
rect 3152 5424 3188 5458
rect 231 5329 292 5368
rect 265 5295 292 5329
rect 231 5256 292 5295
rect 265 5222 292 5256
rect 231 5183 292 5222
rect 265 5149 292 5183
rect 231 5110 292 5149
rect 265 5076 292 5110
rect 231 5037 292 5076
rect 265 5003 292 5037
rect 231 4965 292 5003
rect 265 4931 292 4965
rect 231 4893 292 4931
rect 265 4859 292 4893
rect 231 4821 292 4859
rect 265 4787 292 4821
rect 231 4749 292 4787
rect 265 4715 292 4749
rect 231 4677 292 4715
rect 265 4643 292 4677
rect 231 4605 292 4643
rect 265 4571 292 4605
rect 231 4533 292 4571
rect 265 4499 292 4533
rect 231 4461 292 4499
rect 265 4427 292 4461
rect 231 4377 292 4427
rect 256 4353 292 4377
rect 256 4319 257 4353
rect 291 4319 292 4353
rect 3152 5390 3153 5424
rect 3187 5390 3188 5424
rect 3152 5356 3188 5390
rect 3152 5322 3153 5356
rect 3187 5322 3188 5356
rect 3152 5288 3188 5322
rect 3152 5254 3153 5288
rect 3187 5254 3188 5288
rect 3152 5220 3188 5254
rect 3152 5186 3153 5220
rect 3187 5186 3188 5220
rect 3152 5152 3188 5186
rect 3152 5118 3153 5152
rect 3187 5118 3188 5152
rect 3152 5084 3188 5118
rect 3152 5050 3153 5084
rect 3187 5050 3188 5084
rect 3152 5016 3188 5050
rect 3152 4982 3153 5016
rect 3187 4982 3188 5016
rect 3152 4948 3188 4982
rect 3152 4914 3153 4948
rect 3187 4914 3188 4948
rect 3152 4880 3188 4914
rect 3152 4846 3153 4880
rect 3187 4846 3188 4880
rect 3152 4812 3188 4846
rect 3152 4778 3153 4812
rect 3187 4778 3188 4812
rect 3152 4744 3188 4778
rect 3152 4710 3153 4744
rect 3187 4710 3188 4744
rect 3152 4676 3188 4710
rect 3152 4642 3153 4676
rect 3187 4642 3188 4676
rect 3152 4608 3188 4642
rect 3152 4574 3153 4608
rect 3187 4574 3188 4608
rect 3152 4540 3188 4574
rect 3152 4506 3153 4540
rect 3187 4506 3188 4540
rect 3152 4472 3188 4506
rect 3152 4438 3153 4472
rect 3187 4438 3188 4472
rect 3152 4404 3188 4438
rect 3152 4370 3153 4404
rect 3187 4370 3188 4404
rect 3152 4336 3188 4370
rect 256 4284 292 4319
rect 256 4250 257 4284
rect 291 4250 292 4284
rect 3152 4302 3153 4336
rect 3187 4302 3188 4336
rect 3152 4268 3188 4302
rect 3530 5542 3651 5575
rect 3530 5508 3531 5542
rect 3565 5541 3651 5542
rect 3685 5541 3719 5575
rect 3753 5541 3787 5575
rect 3821 5541 3855 5575
rect 3889 5541 3923 5575
rect 3957 5541 3991 5575
rect 4025 5541 4059 5575
rect 4093 5541 4127 5575
rect 4161 5541 4195 5575
rect 4229 5541 4263 5575
rect 4297 5541 4331 5575
rect 4365 5541 4399 5575
rect 4433 5541 4467 5575
rect 4501 5541 4535 5575
rect 4569 5541 4603 5575
rect 4637 5541 4671 5575
rect 4705 5541 4739 5575
rect 4773 5541 4807 5575
rect 4841 5541 4875 5575
rect 4909 5541 4943 5575
rect 4977 5541 5011 5575
rect 5045 5541 5079 5575
rect 5113 5541 5147 5575
rect 5181 5541 5215 5575
rect 5249 5541 5283 5575
rect 5317 5541 5351 5575
rect 5385 5541 5588 5575
rect 5622 5541 5656 5575
rect 3565 5540 5656 5541
rect 3565 5508 3566 5540
rect 3530 5474 3566 5508
rect 3530 5440 3531 5474
rect 3565 5440 3566 5474
rect 3530 5406 3566 5440
rect 5620 5456 5656 5540
rect 3530 5372 3531 5406
rect 3565 5372 3566 5406
rect 3530 5338 3566 5372
rect 3530 5304 3531 5338
rect 3565 5304 3566 5338
rect 3530 5270 3566 5304
rect 3530 5236 3531 5270
rect 3565 5236 3566 5270
rect 3530 5202 3566 5236
rect 3530 5168 3531 5202
rect 3565 5168 3566 5202
rect 3530 5134 3566 5168
rect 3530 5100 3531 5134
rect 3565 5100 3566 5134
rect 3530 5066 3566 5100
rect 3530 5032 3531 5066
rect 3565 5032 3566 5066
rect 3530 4998 3566 5032
rect 3530 4964 3531 4998
rect 3565 4964 3566 4998
rect 3530 4930 3566 4964
rect 3530 4896 3531 4930
rect 3565 4896 3566 4930
rect 3530 4862 3566 4896
rect 3530 4828 3531 4862
rect 3565 4828 3566 4862
rect 3530 4794 3566 4828
rect 3530 4760 3531 4794
rect 3565 4760 3566 4794
rect 3530 4726 3566 4760
rect 3530 4692 3531 4726
rect 3565 4692 3566 4726
rect 3530 4658 3566 4692
rect 3530 4624 3531 4658
rect 3565 4624 3566 4658
rect 3530 4590 3566 4624
rect 3530 4556 3531 4590
rect 3565 4556 3566 4590
rect 3530 4522 3566 4556
rect 3530 4488 3531 4522
rect 3565 4488 3566 4522
rect 3530 4454 3566 4488
rect 3530 4420 3531 4454
rect 3565 4420 3566 4454
rect 3530 4336 3566 4420
rect 5620 5422 5621 5456
rect 5655 5422 5656 5456
rect 5620 5388 5656 5422
rect 5620 5354 5621 5388
rect 5655 5354 5656 5388
rect 5620 5320 5656 5354
rect 5620 5286 5621 5320
rect 5655 5286 5656 5320
rect 5620 5252 5656 5286
rect 5620 5218 5621 5252
rect 5655 5218 5656 5252
rect 5620 5184 5656 5218
rect 5620 5150 5621 5184
rect 5655 5150 5656 5184
rect 5620 5116 5656 5150
rect 5620 5082 5621 5116
rect 5655 5082 5656 5116
rect 5620 5048 5656 5082
rect 5620 5014 5621 5048
rect 5655 5014 5656 5048
rect 5620 4980 5656 5014
rect 5620 4946 5621 4980
rect 5655 4946 5656 4980
rect 5620 4912 5656 4946
rect 5620 4878 5621 4912
rect 5655 4878 5656 4912
rect 5620 4844 5656 4878
rect 5620 4810 5621 4844
rect 5655 4810 5656 4844
rect 5620 4776 5656 4810
rect 5620 4742 5621 4776
rect 5655 4742 5656 4776
rect 5620 4708 5656 4742
rect 5620 4674 5621 4708
rect 5655 4674 5656 4708
rect 5620 4640 5656 4674
rect 5620 4606 5621 4640
rect 5655 4606 5656 4640
rect 5620 4572 5656 4606
rect 5620 4538 5621 4572
rect 5655 4538 5656 4572
rect 5620 4504 5656 4538
rect 5620 4470 5621 4504
rect 5655 4470 5656 4504
rect 5620 4436 5656 4470
rect 5620 4402 5621 4436
rect 5655 4402 5656 4436
rect 5620 4368 5656 4402
rect 5620 4336 5621 4368
rect 3530 4335 5621 4336
rect 3530 4301 3564 4335
rect 3598 4301 3632 4335
rect 3666 4301 3700 4335
rect 3734 4301 3768 4335
rect 3802 4301 3836 4335
rect 3870 4301 3904 4335
rect 3938 4301 3972 4335
rect 4006 4301 4040 4335
rect 4074 4301 4108 4335
rect 4142 4301 4176 4335
rect 4210 4301 4244 4335
rect 4278 4301 4312 4335
rect 4346 4301 4380 4335
rect 4414 4301 4448 4335
rect 4482 4301 4516 4335
rect 4550 4301 4584 4335
rect 4618 4301 4652 4335
rect 4686 4301 4720 4335
rect 4754 4301 4788 4335
rect 4822 4301 4856 4335
rect 4890 4301 4924 4335
rect 4958 4301 4992 4335
rect 5026 4301 5060 4335
rect 5094 4301 5128 4335
rect 5162 4301 5196 4335
rect 5230 4301 5264 4335
rect 5298 4301 5332 4335
rect 5366 4301 5400 4335
rect 5434 4301 5468 4335
rect 5502 4301 5536 4335
rect 5570 4334 5621 4335
rect 5655 4334 5656 4368
rect 5570 4301 5656 4334
rect 3530 4300 5656 4301
rect 256 4215 292 4250
rect 256 4181 257 4215
rect 291 4181 292 4215
rect 3152 4234 3153 4268
rect 3187 4234 3188 4268
rect 256 4146 292 4181
rect 256 4112 257 4146
rect 291 4112 292 4146
rect 256 4077 292 4112
rect 3152 4200 3188 4234
rect 3152 4166 3153 4200
rect 3187 4166 3188 4200
rect 3152 4132 3188 4166
rect 3152 4098 3153 4132
rect 3187 4098 3188 4132
rect 256 4043 257 4077
rect 291 4043 292 4077
rect 256 4008 292 4043
rect 256 3974 257 4008
rect 291 3974 292 4008
rect 256 3939 292 3974
rect 256 3905 257 3939
rect 291 3905 292 3939
rect 256 3870 292 3905
rect 256 3836 257 3870
rect 291 3836 292 3870
rect 256 3801 292 3836
rect 256 3767 257 3801
rect 291 3767 292 3801
rect 256 3732 292 3767
rect 256 3698 257 3732
rect 291 3698 292 3732
rect 256 3663 292 3698
rect 256 3629 257 3663
rect 291 3629 292 3663
rect 256 3594 292 3629
rect 256 3560 257 3594
rect 291 3560 292 3594
rect 256 3525 292 3560
rect 256 3491 257 3525
rect 291 3491 292 3525
rect 256 3456 292 3491
rect 256 3422 257 3456
rect 291 3422 292 3456
rect 256 3387 292 3422
rect 256 3353 257 3387
rect 291 3353 292 3387
rect 256 3318 292 3353
rect 256 3284 257 3318
rect 291 3284 292 3318
rect 256 3249 292 3284
rect 256 3215 257 3249
rect 291 3215 292 3249
rect 256 3180 292 3215
rect 256 3146 257 3180
rect 291 3146 292 3180
rect 256 3111 292 3146
rect 256 3077 257 3111
rect 291 3077 292 3111
rect 256 3042 292 3077
rect 256 3008 257 3042
rect 291 3008 292 3042
rect 256 2973 292 3008
rect 256 2939 257 2973
rect 291 2939 292 2973
rect 256 2904 292 2939
rect 256 2870 257 2904
rect 291 2870 292 2904
rect 256 2835 292 2870
rect 256 2801 257 2835
rect 291 2801 292 2835
rect 256 2766 292 2801
rect 256 2732 257 2766
rect 291 2732 292 2766
rect 256 2697 292 2732
rect 256 2663 257 2697
rect 291 2663 292 2697
rect 256 2628 292 2663
rect 256 2594 257 2628
rect 291 2594 292 2628
rect 256 2559 292 2594
rect 256 2525 257 2559
rect 291 2525 292 2559
rect 256 2490 292 2525
rect 256 2456 257 2490
rect 291 2456 292 2490
rect 256 2421 292 2456
rect 256 2387 257 2421
rect 291 2387 292 2421
rect 256 2352 292 2387
rect 256 2318 257 2352
rect 291 2318 292 2352
rect 256 2283 292 2318
rect 256 2249 257 2283
rect 291 2249 292 2283
rect 256 2214 292 2249
rect 256 2180 257 2214
rect 291 2180 292 2214
rect 256 2145 292 2180
rect 256 2111 257 2145
rect 291 2111 292 2145
rect 256 2076 292 2111
rect 256 2042 257 2076
rect 291 2042 292 2076
rect 256 2007 292 2042
rect 256 1973 257 2007
rect 291 1973 292 2007
rect 256 1938 292 1973
rect 256 1904 257 1938
rect 291 1904 292 1938
rect 256 1869 292 1904
rect 256 1835 257 1869
rect 291 1835 292 1869
rect 256 1800 292 1835
rect 256 1766 257 1800
rect 291 1766 292 1800
rect 256 1731 292 1766
rect 256 1697 257 1731
rect 291 1697 292 1731
rect 256 1662 292 1697
rect 256 1628 257 1662
rect 291 1628 292 1662
rect 256 1593 292 1628
rect 256 1559 257 1593
rect 291 1559 292 1593
rect 256 1524 292 1559
rect 256 1490 257 1524
rect 291 1490 292 1524
rect 256 1456 292 1490
rect 256 1422 257 1456
rect 291 1422 292 1456
rect 256 1388 292 1422
rect 256 1354 257 1388
rect 291 1354 292 1388
rect 256 1320 292 1354
rect 256 1286 257 1320
rect 291 1286 292 1320
rect 256 1252 292 1286
rect 256 1218 257 1252
rect 291 1218 292 1252
rect 256 1184 292 1218
rect 256 1150 257 1184
rect 291 1150 292 1184
rect 256 1116 292 1150
rect 256 1082 257 1116
rect 291 1082 292 1116
rect 256 1048 292 1082
rect 256 1014 257 1048
rect 291 1014 292 1048
rect 256 980 292 1014
rect 256 946 257 980
rect 291 946 292 980
rect 256 912 292 946
rect 256 878 257 912
rect 291 878 292 912
rect 256 844 292 878
rect 256 810 257 844
rect 291 810 292 844
rect 256 776 292 810
rect 256 742 257 776
rect 291 742 292 776
rect 256 708 292 742
rect 256 674 257 708
rect 291 674 292 708
rect 256 640 292 674
rect 256 606 257 640
rect 291 606 292 640
rect 256 572 292 606
rect 256 538 257 572
rect 291 538 292 572
rect 256 504 292 538
rect 256 470 257 504
rect 291 470 292 504
rect 256 436 292 470
rect 256 402 257 436
rect 291 402 292 436
rect 3152 4064 3188 4098
rect 3152 4030 3153 4064
rect 3187 4030 3188 4064
rect 3152 3996 3188 4030
rect 3152 3962 3153 3996
rect 3187 3962 3188 3996
rect 3152 3928 3188 3962
rect 3152 3894 3153 3928
rect 3187 3894 3188 3928
rect 3152 3860 3188 3894
rect 3152 3826 3153 3860
rect 3187 3826 3188 3860
rect 3152 3792 3188 3826
rect 3152 3758 3153 3792
rect 3187 3758 3188 3792
rect 3152 3724 3188 3758
rect 3152 3690 3153 3724
rect 3187 3690 3188 3724
rect 3152 3656 3188 3690
rect 3152 3622 3153 3656
rect 3187 3622 3188 3656
rect 3152 3588 3188 3622
rect 3152 3554 3153 3588
rect 3187 3554 3188 3588
rect 3152 3520 3188 3554
rect 3152 3486 3153 3520
rect 3187 3486 3188 3520
rect 3152 3452 3188 3486
rect 3152 3418 3153 3452
rect 3187 3418 3188 3452
rect 3152 3384 3188 3418
rect 3152 3350 3153 3384
rect 3187 3350 3188 3384
rect 3152 3316 3188 3350
rect 3152 3282 3153 3316
rect 3187 3282 3188 3316
rect 3152 3248 3188 3282
rect 3152 3214 3153 3248
rect 3187 3214 3188 3248
rect 3152 3180 3188 3214
rect 3152 3146 3153 3180
rect 3187 3146 3188 3180
rect 3152 3112 3188 3146
rect 3152 3078 3153 3112
rect 3187 3078 3188 3112
rect 3152 3044 3188 3078
rect 3152 3010 3153 3044
rect 3187 3010 3188 3044
rect 3152 2976 3188 3010
rect 3152 2942 3153 2976
rect 3187 2942 3188 2976
rect 3152 2908 3188 2942
rect 3152 2874 3153 2908
rect 3187 2874 3188 2908
rect 3152 2840 3188 2874
rect 3152 2806 3153 2840
rect 3187 2806 3188 2840
rect 3152 2772 3188 2806
rect 3152 2738 3153 2772
rect 3187 2738 3188 2772
rect 3152 2704 3188 2738
rect 3152 2670 3153 2704
rect 3187 2670 3188 2704
rect 3152 2636 3188 2670
rect 3152 2602 3153 2636
rect 3187 2602 3188 2636
rect 3152 2568 3188 2602
rect 3152 2534 3153 2568
rect 3187 2534 3188 2568
rect 3152 2500 3188 2534
rect 3152 2466 3153 2500
rect 3187 2466 3188 2500
rect 3152 2432 3188 2466
rect 3152 2398 3153 2432
rect 3187 2398 3188 2432
rect 3152 2364 3188 2398
rect 3152 2330 3153 2364
rect 3187 2330 3188 2364
rect 3152 2296 3188 2330
rect 3152 2262 3153 2296
rect 3187 2262 3188 2296
rect 3152 2228 3188 2262
rect 3152 2194 3153 2228
rect 3187 2194 3188 2228
rect 3152 2160 3188 2194
rect 3152 2126 3153 2160
rect 3187 2126 3188 2160
rect 3152 2092 3188 2126
rect 3152 2058 3153 2092
rect 3187 2058 3188 2092
rect 3152 2024 3188 2058
rect 3152 1990 3153 2024
rect 3187 1990 3188 2024
rect 3152 1956 3188 1990
rect 3152 1922 3153 1956
rect 3187 1922 3188 1956
rect 3152 1888 3188 1922
rect 3152 1854 3153 1888
rect 3187 1854 3188 1888
rect 3152 1820 3188 1854
rect 3152 1786 3153 1820
rect 3187 1786 3188 1820
rect 3152 1752 3188 1786
rect 3152 1718 3153 1752
rect 3187 1718 3188 1752
rect 3152 1684 3188 1718
rect 3152 1650 3153 1684
rect 3187 1650 3188 1684
rect 3152 1616 3188 1650
rect 3152 1582 3153 1616
rect 3187 1582 3188 1616
rect 3152 1548 3188 1582
rect 3152 1514 3153 1548
rect 3187 1514 3188 1548
rect 3152 1480 3188 1514
rect 3152 1446 3153 1480
rect 3187 1446 3188 1480
rect 3152 1412 3188 1446
rect 3152 1378 3153 1412
rect 3187 1378 3188 1412
rect 3152 1344 3188 1378
rect 3152 1310 3153 1344
rect 3187 1310 3188 1344
rect 3152 1276 3188 1310
rect 3152 1242 3153 1276
rect 3187 1242 3188 1276
rect 3152 1208 3188 1242
rect 3152 1174 3153 1208
rect 3187 1174 3188 1208
rect 3152 1140 3188 1174
rect 3152 1106 3153 1140
rect 3187 1106 3188 1140
rect 3152 1072 3188 1106
rect 3152 1038 3153 1072
rect 3187 1038 3188 1072
rect 3152 1004 3188 1038
rect 3152 970 3153 1004
rect 3187 970 3188 1004
rect 3152 936 3188 970
rect 3152 902 3153 936
rect 3187 902 3188 936
rect 3152 868 3188 902
rect 3152 834 3153 868
rect 3187 834 3188 868
rect 3152 800 3188 834
rect 3152 766 3153 800
rect 3187 766 3188 800
rect 3152 732 3188 766
rect 3152 698 3153 732
rect 3187 698 3188 732
rect 3152 664 3188 698
rect 3152 630 3153 664
rect 3187 630 3188 664
rect 3152 596 3188 630
rect 3152 562 3153 596
rect 3187 562 3188 596
rect 3152 528 3188 562
rect 3152 494 3153 528
rect 3187 494 3188 528
rect 3152 460 3188 494
rect 256 292 292 402
rect 3152 426 3153 460
rect 3187 426 3188 460
rect 3152 392 3188 426
rect 3152 358 3153 392
rect 3187 358 3188 392
rect 3152 324 3188 358
rect 3152 292 3153 324
rect 256 291 3153 292
rect 256 257 290 291
rect 324 257 358 291
rect 392 257 426 291
rect 460 257 494 291
rect 528 257 562 291
rect 596 257 630 291
rect 664 257 698 291
rect 732 257 766 291
rect 800 257 834 291
rect 868 257 902 291
rect 936 257 970 291
rect 1004 257 1038 291
rect 1072 257 1106 291
rect 1140 257 1174 291
rect 1208 257 1242 291
rect 1276 257 1310 291
rect 1344 257 1378 291
rect 1412 257 1446 291
rect 1480 257 1514 291
rect 1548 257 1582 291
rect 1616 257 1650 291
rect 1684 257 1718 291
rect 1752 257 1786 291
rect 1820 257 1854 291
rect 1888 257 1922 291
rect 1956 257 1990 291
rect 2024 257 2058 291
rect 2092 257 2126 291
rect 2160 257 2194 291
rect 2228 257 2262 291
rect 2296 257 2330 291
rect 2364 257 2398 291
rect 2432 257 2466 291
rect 2500 257 2534 291
rect 2568 257 2602 291
rect 2636 257 2670 291
rect 2704 257 2738 291
rect 2772 257 2806 291
rect 2840 257 2874 291
rect 2908 257 2942 291
rect 2976 257 3010 291
rect 3044 257 3078 291
rect 3112 290 3153 291
rect 3187 290 3188 324
rect 3112 257 3188 290
rect 256 256 3188 257
<< mvnsubdiff >>
rect 67 27869 2369 27870
rect 67 27836 165 27869
rect 67 27802 68 27836
rect 102 27835 165 27836
rect 199 27835 233 27869
rect 267 27835 301 27869
rect 335 27835 369 27869
rect 403 27835 437 27869
rect 471 27835 505 27869
rect 539 27835 573 27869
rect 607 27835 641 27869
rect 675 27835 709 27869
rect 743 27835 777 27869
rect 811 27835 845 27869
rect 879 27835 913 27869
rect 947 27835 981 27869
rect 1015 27835 1049 27869
rect 1083 27835 1117 27869
rect 1151 27835 1185 27869
rect 1219 27835 1253 27869
rect 1287 27835 1321 27869
rect 1355 27835 1389 27869
rect 1423 27835 1457 27869
rect 1491 27835 1525 27869
rect 1559 27835 1593 27869
rect 1627 27835 1661 27869
rect 1695 27835 1729 27869
rect 1763 27835 1797 27869
rect 1831 27835 1865 27869
rect 1899 27835 1998 27869
rect 2032 27835 2066 27869
rect 2100 27835 2134 27869
rect 2168 27835 2202 27869
rect 2236 27835 2369 27869
rect 102 27834 2369 27835
rect 102 27802 103 27834
rect 67 27768 103 27802
rect 67 27734 68 27768
rect 102 27734 103 27768
rect 67 27700 103 27734
rect 67 27666 68 27700
rect 102 27666 103 27700
rect 2333 27797 2369 27834
rect 2333 27763 2334 27797
rect 2368 27763 2369 27797
rect 2333 27729 2369 27763
rect 2333 27695 2334 27729
rect 2368 27695 2369 27729
rect 67 27632 103 27666
rect 67 27598 68 27632
rect 102 27598 103 27632
rect 67 27564 103 27598
rect 67 27530 68 27564
rect 102 27530 103 27564
rect 67 27496 103 27530
rect 67 27462 68 27496
rect 102 27462 103 27496
rect 67 27428 103 27462
rect 67 27394 68 27428
rect 102 27394 103 27428
rect 67 27360 103 27394
rect 67 27326 68 27360
rect 102 27326 103 27360
rect 67 27292 103 27326
rect 67 27258 68 27292
rect 102 27258 103 27292
rect 67 27224 103 27258
rect 67 27190 68 27224
rect 102 27190 103 27224
rect 67 27156 103 27190
rect 67 27122 68 27156
rect 102 27122 103 27156
rect 67 27088 103 27122
rect 67 27054 68 27088
rect 102 27054 103 27088
rect 67 27020 103 27054
rect 67 26986 68 27020
rect 102 26986 103 27020
rect 67 26952 103 26986
rect 67 26918 68 26952
rect 102 26918 103 26952
rect 67 26884 103 26918
rect 67 26850 68 26884
rect 102 26850 103 26884
rect 67 26816 103 26850
rect 67 26782 68 26816
rect 102 26782 103 26816
rect 67 26748 103 26782
rect 67 26714 68 26748
rect 102 26714 103 26748
rect 67 26680 103 26714
rect 67 26646 68 26680
rect 102 26646 103 26680
rect 67 26612 103 26646
rect 67 26578 68 26612
rect 102 26578 103 26612
rect 67 26544 103 26578
rect 67 26510 68 26544
rect 102 26510 103 26544
rect 67 26476 103 26510
rect 67 26442 68 26476
rect 102 26442 103 26476
rect 67 26408 103 26442
rect 67 26374 68 26408
rect 102 26374 103 26408
rect 67 26340 103 26374
rect 67 26306 68 26340
rect 102 26306 103 26340
rect 67 26272 103 26306
rect 67 26238 68 26272
rect 102 26238 103 26272
rect 67 26204 103 26238
rect 67 26170 68 26204
rect 102 26170 103 26204
rect 67 26136 103 26170
rect 67 26102 68 26136
rect 102 26102 103 26136
rect 67 26068 103 26102
rect 67 26034 68 26068
rect 102 26034 103 26068
rect 67 26000 103 26034
rect 67 25966 68 26000
rect 102 25966 103 26000
rect 67 25932 103 25966
rect 67 25898 68 25932
rect 102 25898 103 25932
rect 67 25864 103 25898
rect 67 25830 68 25864
rect 102 25830 103 25864
rect 67 25796 103 25830
rect 67 25762 68 25796
rect 102 25762 103 25796
rect 67 25690 103 25762
rect 2333 27661 2369 27695
rect 2333 27627 2334 27661
rect 2368 27627 2369 27661
rect 2333 27593 2369 27627
rect 2333 27559 2334 27593
rect 2368 27559 2369 27593
rect 2333 27525 2369 27559
rect 2333 27491 2334 27525
rect 2368 27491 2369 27525
rect 2333 27457 2369 27491
rect 2333 27423 2334 27457
rect 2368 27423 2369 27457
rect 2333 27389 2369 27423
rect 2333 27355 2334 27389
rect 2368 27355 2369 27389
rect 2333 27321 2369 27355
rect 2333 27287 2334 27321
rect 2368 27287 2369 27321
rect 2333 27253 2369 27287
rect 2333 27219 2334 27253
rect 2368 27219 2369 27253
rect 2333 27185 2369 27219
rect 2333 27151 2334 27185
rect 2368 27151 2369 27185
rect 2333 27117 2369 27151
rect 2333 27083 2334 27117
rect 2368 27083 2369 27117
rect 2333 27049 2369 27083
rect 2333 27015 2334 27049
rect 2368 27015 2369 27049
rect 2333 26981 2369 27015
rect 2333 26947 2334 26981
rect 2368 26947 2369 26981
rect 2333 26913 2369 26947
rect 2333 26879 2334 26913
rect 2368 26879 2369 26913
rect 2333 26845 2369 26879
rect 2333 26811 2334 26845
rect 2368 26811 2369 26845
rect 2333 26777 2369 26811
rect 2333 26743 2334 26777
rect 2368 26743 2369 26777
rect 2333 26709 2369 26743
rect 2333 26675 2334 26709
rect 2368 26675 2369 26709
rect 2333 26641 2369 26675
rect 2333 26607 2334 26641
rect 2368 26607 2369 26641
rect 2333 26573 2369 26607
rect 2333 26539 2334 26573
rect 2368 26539 2369 26573
rect 2333 26505 2369 26539
rect 2333 26471 2334 26505
rect 2368 26471 2369 26505
rect 2333 26437 2369 26471
rect 2333 26403 2334 26437
rect 2368 26403 2369 26437
rect 2333 26369 2369 26403
rect 2333 26335 2334 26369
rect 2368 26335 2369 26369
rect 2333 26301 2369 26335
rect 2333 26267 2334 26301
rect 2368 26267 2369 26301
rect 2333 26233 2369 26267
rect 2333 26199 2334 26233
rect 2368 26199 2369 26233
rect 2333 26165 2369 26199
rect 2333 26131 2334 26165
rect 2368 26131 2369 26165
rect 2333 26097 2369 26131
rect 2333 26063 2334 26097
rect 2368 26063 2369 26097
rect 2333 26029 2369 26063
rect 2333 25995 2334 26029
rect 2368 25995 2369 26029
rect 2333 25961 2369 25995
rect 2333 25927 2334 25961
rect 2368 25927 2369 25961
rect 2333 25893 2369 25927
rect 2333 25859 2334 25893
rect 2368 25859 2369 25893
rect 2333 25825 2369 25859
rect 2333 25791 2334 25825
rect 2368 25791 2369 25825
rect 2333 25757 2369 25791
rect 2333 25723 2334 25757
rect 2368 25723 2369 25757
rect 2333 25689 2369 25723
rect 2333 25655 2334 25689
rect 2368 25655 2369 25689
rect 2333 25621 2369 25655
rect 2333 25587 2334 25621
rect 2368 25587 2369 25621
rect 2333 25553 2369 25587
rect 2333 25519 2334 25553
rect 2368 25519 2369 25553
rect 2333 25485 2369 25519
rect 2333 25451 2334 25485
rect 2368 25451 2369 25485
rect 2333 25417 2369 25451
rect 2333 25383 2334 25417
rect 2368 25383 2369 25417
rect 2333 25349 2369 25383
rect 2333 25315 2334 25349
rect 2368 25315 2369 25349
rect 2333 25281 2369 25315
rect 2333 25247 2334 25281
rect 2368 25247 2369 25281
rect 2333 25213 2369 25247
rect 2333 25179 2334 25213
rect 2368 25179 2369 25213
rect 2333 25145 2369 25179
rect 2333 25111 2334 25145
rect 2368 25111 2369 25145
rect 2333 25077 2369 25111
rect 2333 25043 2334 25077
rect 2368 25043 2369 25077
rect 2333 25009 2369 25043
rect 2333 24975 2334 25009
rect 2368 24975 2369 25009
rect 2333 24941 2369 24975
rect 2333 24907 2334 24941
rect 2368 24907 2369 24941
rect 2333 24873 2369 24907
rect 2333 24839 2334 24873
rect 2368 24839 2369 24873
rect 2333 24805 2369 24839
rect 2333 24771 2334 24805
rect 2368 24771 2369 24805
rect 2333 24737 2369 24771
rect 2333 24703 2334 24737
rect 2368 24703 2369 24737
rect 2333 24669 2369 24703
rect 2333 24635 2334 24669
rect 2368 24635 2369 24669
rect 2333 24601 2369 24635
rect 2333 24567 2334 24601
rect 2368 24567 2369 24601
rect 2333 24533 2369 24567
rect 2333 24499 2334 24533
rect 2368 24499 2369 24533
rect 2333 24465 2369 24499
rect 2333 24431 2334 24465
rect 2368 24431 2369 24465
rect 2333 24397 2369 24431
rect 2333 24363 2334 24397
rect 2368 24363 2369 24397
rect 2333 24329 2369 24363
rect 2333 24295 2334 24329
rect 2368 24295 2369 24329
rect 2333 24261 2369 24295
rect 2333 24227 2334 24261
rect 2368 24227 2369 24261
rect 2333 24193 2369 24227
rect 2333 24159 2334 24193
rect 2368 24159 2369 24193
rect 2333 24125 2369 24159
rect 2333 24091 2334 24125
rect 2368 24091 2369 24125
rect 2333 24057 2369 24091
rect 2333 24023 2334 24057
rect 2368 24023 2369 24057
rect 2333 23989 2369 24023
rect 2333 23955 2334 23989
rect 2368 23955 2369 23989
rect 2333 23921 2369 23955
rect 2333 23887 2334 23921
rect 2368 23887 2369 23921
rect 2333 23853 2369 23887
rect 2333 23819 2334 23853
rect 2368 23819 2369 23853
rect 2333 23785 2369 23819
rect 2333 23751 2334 23785
rect 2368 23751 2369 23785
rect 2333 23717 2369 23751
rect 2333 23683 2334 23717
rect 2368 23683 2369 23717
rect 2333 23649 2369 23683
rect 2333 23615 2334 23649
rect 2368 23615 2369 23649
rect 2333 23581 2369 23615
rect 2333 23547 2334 23581
rect 2368 23547 2369 23581
rect 2333 23513 2369 23547
rect 2333 23479 2334 23513
rect 2368 23479 2369 23513
rect 2333 23445 2369 23479
rect 2333 23411 2334 23445
rect 2368 23411 2369 23445
rect 2333 23377 2369 23411
rect 2333 23343 2334 23377
rect 2368 23343 2369 23377
rect 2333 23309 2369 23343
rect 2333 23275 2334 23309
rect 2368 23275 2369 23309
rect 2333 23241 2369 23275
rect 2333 23207 2334 23241
rect 2368 23207 2369 23241
rect 2333 23173 2369 23207
rect 2333 23139 2334 23173
rect 2368 23139 2369 23173
rect 2333 23105 2369 23139
rect 2333 23071 2334 23105
rect 2368 23071 2369 23105
rect 2333 23037 2369 23071
rect 2333 23003 2334 23037
rect 2368 23003 2369 23037
rect 2333 22969 2369 23003
rect 2333 22935 2334 22969
rect 2368 22935 2369 22969
rect 2333 22901 2369 22935
rect 2333 22867 2334 22901
rect 2368 22867 2369 22901
rect 2333 22833 2369 22867
rect 2333 22799 2334 22833
rect 2368 22799 2369 22833
rect 2333 22765 2369 22799
rect 2333 22731 2334 22765
rect 2368 22731 2369 22765
rect 2333 22697 2369 22731
rect 2333 22663 2334 22697
rect 2368 22663 2369 22697
rect 2333 22629 2369 22663
rect 2333 22595 2334 22629
rect 2368 22595 2369 22629
rect 2333 22561 2369 22595
rect 2333 22527 2334 22561
rect 2368 22527 2369 22561
rect 2333 22493 2369 22527
rect 2333 22459 2334 22493
rect 2368 22459 2369 22493
rect 2333 22425 2369 22459
rect 2333 22391 2334 22425
rect 2368 22391 2369 22425
rect 2333 22357 2369 22391
rect 2333 22323 2334 22357
rect 2368 22323 2369 22357
rect 2333 22289 2369 22323
rect 2333 22255 2334 22289
rect 2368 22255 2369 22289
rect 2333 22221 2369 22255
rect 2333 22187 2334 22221
rect 2368 22187 2369 22221
rect 2333 22153 2369 22187
rect 2333 22119 2334 22153
rect 2368 22119 2369 22153
rect 2333 22085 2369 22119
rect 2333 22051 2334 22085
rect 2368 22051 2369 22085
rect 2333 22017 2369 22051
rect 2333 21983 2334 22017
rect 2368 21983 2369 22017
rect 2333 21949 2369 21983
rect 2333 21915 2334 21949
rect 2368 21915 2369 21949
rect 2333 21881 2369 21915
rect 2333 21847 2334 21881
rect 2368 21847 2369 21881
rect 2333 21813 2369 21847
rect 2333 21779 2334 21813
rect 2368 21779 2369 21813
rect 2333 21745 2369 21779
rect 2333 21711 2334 21745
rect 2368 21711 2369 21745
rect 2333 21677 2369 21711
rect 2333 21643 2334 21677
rect 2368 21643 2369 21677
rect 2333 21609 2369 21643
rect 2333 21575 2334 21609
rect 2368 21575 2369 21609
rect 2333 21541 2369 21575
rect 2333 21507 2334 21541
rect 2368 21507 2369 21541
rect 2333 21473 2369 21507
rect 2333 21439 2334 21473
rect 2368 21439 2369 21473
rect 2333 21405 2369 21439
rect 2333 21371 2334 21405
rect 2368 21371 2369 21405
rect 2333 21337 2369 21371
rect 2333 21303 2334 21337
rect 2368 21303 2369 21337
rect 2333 21269 2369 21303
rect 2333 21235 2334 21269
rect 2368 21235 2369 21269
rect 2333 21201 2369 21235
rect 2333 21167 2334 21201
rect 2368 21167 2369 21201
rect 2333 21133 2369 21167
rect 2333 21099 2334 21133
rect 2368 21099 2369 21133
rect 2333 21065 2369 21099
rect 2333 21031 2334 21065
rect 2368 21031 2369 21065
rect 2333 20997 2369 21031
rect 2333 20963 2334 20997
rect 2368 20963 2369 20997
rect 2333 20929 2369 20963
rect 2333 20895 2334 20929
rect 2368 20895 2369 20929
rect 2333 20861 2369 20895
rect 2333 20827 2334 20861
rect 2368 20827 2369 20861
rect 2333 20793 2369 20827
rect 2333 20759 2334 20793
rect 2368 20759 2369 20793
rect 2333 20725 2369 20759
rect 2333 20691 2334 20725
rect 2368 20691 2369 20725
rect 2333 20657 2369 20691
rect 2333 20623 2334 20657
rect 2368 20623 2369 20657
rect 2333 20589 2369 20623
rect 2333 20555 2334 20589
rect 2368 20555 2369 20589
rect 2333 20521 2369 20555
rect 2333 20487 2334 20521
rect 2368 20487 2369 20521
rect 2333 20453 2369 20487
rect 2333 20419 2334 20453
rect 2368 20419 2369 20453
rect 2333 20385 2369 20419
rect 2333 20351 2334 20385
rect 2368 20351 2369 20385
rect 2333 20317 2369 20351
rect 2333 20283 2334 20317
rect 2368 20283 2369 20317
rect 2333 20249 2369 20283
rect 2333 20215 2334 20249
rect 2368 20215 2369 20249
rect 2333 20181 2369 20215
rect 2333 20147 2334 20181
rect 2368 20147 2369 20181
rect 2333 20113 2369 20147
rect 2333 20079 2334 20113
rect 2368 20079 2369 20113
rect 2333 20045 2369 20079
rect 2333 20011 2334 20045
rect 2368 20011 2369 20045
rect 2333 19977 2369 20011
rect 2333 19943 2334 19977
rect 2368 19943 2369 19977
rect 2333 19909 2369 19943
rect 2333 19875 2334 19909
rect 2368 19875 2369 19909
rect 2333 19841 2369 19875
rect 2333 19807 2334 19841
rect 2368 19807 2369 19841
rect 2333 19773 2369 19807
rect 2333 19739 2334 19773
rect 2368 19739 2369 19773
rect 2333 19705 2369 19739
rect 2333 19671 2334 19705
rect 2368 19671 2369 19705
rect 2333 19637 2369 19671
rect 2333 19603 2334 19637
rect 2368 19603 2369 19637
rect 2333 19569 2369 19603
rect 2333 19535 2334 19569
rect 2368 19535 2369 19569
rect 2333 19501 2369 19535
rect 2333 19467 2334 19501
rect 2368 19467 2369 19501
rect 2333 19433 2369 19467
rect 2333 19399 2334 19433
rect 2368 19399 2369 19433
rect 2333 19365 2369 19399
rect 2333 19331 2334 19365
rect 2368 19331 2369 19365
rect 2333 19297 2369 19331
rect 2333 19263 2334 19297
rect 2368 19263 2369 19297
rect 2333 19229 2369 19263
rect 2333 19195 2334 19229
rect 2368 19195 2369 19229
rect 2333 19161 2369 19195
rect 2333 19127 2334 19161
rect 2368 19127 2369 19161
rect 2333 19093 2369 19127
rect 2333 19059 2334 19093
rect 2368 19059 2369 19093
rect 2333 19025 2369 19059
rect 2333 18991 2334 19025
rect 2368 18991 2369 19025
rect 2333 18957 2369 18991
rect 2333 18923 2334 18957
rect 2368 18923 2369 18957
rect 2333 18889 2369 18923
rect 2333 18855 2334 18889
rect 2368 18855 2369 18889
rect 2333 18821 2369 18855
rect 2333 18787 2334 18821
rect 2368 18787 2369 18821
rect 2333 18753 2369 18787
rect 2333 18719 2334 18753
rect 2368 18719 2369 18753
rect 2333 18685 2369 18719
rect 2333 18651 2334 18685
rect 2368 18651 2369 18685
rect 2333 18617 2369 18651
rect 2333 18583 2334 18617
rect 2368 18583 2369 18617
rect 2333 18549 2369 18583
rect 2333 18515 2334 18549
rect 2368 18515 2369 18549
rect 2333 18481 2369 18515
rect 2333 18447 2334 18481
rect 2368 18447 2369 18481
rect 2333 18413 2369 18447
rect 2333 18379 2334 18413
rect 2368 18379 2369 18413
rect 2333 18345 2369 18379
rect 2333 18311 2334 18345
rect 2368 18311 2369 18345
rect 2333 18277 2369 18311
rect 2333 18243 2334 18277
rect 2368 18243 2369 18277
rect 2333 18209 2369 18243
rect 2333 18175 2334 18209
rect 2368 18175 2369 18209
rect 2333 18141 2369 18175
rect 2333 18107 2334 18141
rect 2368 18107 2369 18141
rect 2333 18073 2369 18107
rect 2333 18039 2334 18073
rect 2368 18039 2369 18073
rect 2333 18005 2369 18039
rect 2333 17971 2334 18005
rect 2368 17971 2369 18005
rect 2333 17937 2369 17971
rect 2333 17903 2334 17937
rect 2368 17903 2369 17937
rect 2333 17869 2369 17903
rect 2333 17835 2334 17869
rect 2368 17835 2369 17869
rect 2333 17801 2369 17835
rect 2333 17767 2334 17801
rect 2368 17767 2369 17801
rect 2333 17733 2369 17767
rect 2333 17699 2334 17733
rect 2368 17699 2369 17733
rect 2333 17665 2369 17699
rect 2333 17631 2334 17665
rect 2368 17631 2369 17665
rect 2333 17597 2369 17631
rect 2333 17563 2334 17597
rect 2368 17563 2369 17597
rect 2333 17529 2369 17563
rect 2333 17495 2334 17529
rect 2368 17495 2369 17529
rect 2333 17461 2369 17495
rect 2333 17427 2334 17461
rect 2368 17427 2369 17461
rect 2333 17393 2369 17427
rect 2333 17359 2334 17393
rect 2368 17359 2369 17393
rect 2333 17325 2369 17359
rect 2333 17291 2334 17325
rect 2368 17291 2369 17325
rect 2333 17257 2369 17291
rect 2333 17223 2334 17257
rect 2368 17223 2369 17257
rect 2333 17189 2369 17223
rect 2333 17155 2334 17189
rect 2368 17155 2369 17189
rect 2333 17121 2369 17155
rect 2333 17087 2334 17121
rect 2368 17087 2369 17121
rect 2333 17053 2369 17087
rect 2333 17019 2334 17053
rect 2368 17019 2369 17053
rect 2333 16985 2369 17019
rect 2333 16951 2334 16985
rect 2368 16951 2369 16985
rect 2333 16917 2369 16951
rect 2333 16883 2334 16917
rect 2368 16883 2369 16917
rect 2333 16849 2369 16883
rect 2333 16815 2334 16849
rect 2368 16815 2369 16849
rect 2333 16781 2369 16815
rect 2333 16747 2334 16781
rect 2368 16747 2369 16781
rect 2333 16713 2369 16747
rect 2333 16679 2334 16713
rect 2368 16679 2369 16713
rect 2333 16645 2369 16679
rect 2333 16611 2334 16645
rect 2368 16611 2369 16645
rect 2333 16577 2369 16611
rect 2333 16543 2334 16577
rect 2368 16543 2369 16577
rect 2333 16509 2369 16543
rect 2333 16475 2334 16509
rect 2368 16475 2369 16509
rect 2333 16441 2369 16475
rect 2333 16407 2334 16441
rect 2368 16407 2369 16441
rect 2333 16373 2369 16407
rect 2333 16339 2334 16373
rect 2368 16339 2369 16373
rect 2333 16305 2369 16339
rect 2333 16271 2334 16305
rect 2368 16271 2369 16305
rect 2333 16237 2369 16271
rect 2333 16203 2334 16237
rect 2368 16203 2369 16237
rect 2333 16169 2369 16203
rect 2333 16135 2334 16169
rect 2368 16135 2369 16169
rect 2333 16101 2369 16135
rect 2333 16067 2334 16101
rect 2368 16067 2369 16101
rect 2333 16033 2369 16067
rect 2333 15999 2334 16033
rect 2368 15999 2369 16033
rect 2333 15965 2369 15999
rect 2333 15931 2334 15965
rect 2368 15931 2369 15965
rect 2333 15897 2369 15931
rect 2333 15863 2334 15897
rect 2368 15863 2369 15897
rect 2333 15829 2369 15863
rect 2333 15795 2334 15829
rect 2368 15795 2369 15829
rect 2333 15761 2369 15795
rect 2333 15727 2334 15761
rect 2368 15727 2369 15761
rect 2333 15693 2369 15727
rect 2333 15659 2334 15693
rect 2368 15659 2369 15693
rect 2333 15625 2369 15659
rect 2333 15591 2334 15625
rect 2368 15591 2369 15625
rect 2333 15557 2369 15591
rect 2333 15523 2334 15557
rect 2368 15523 2369 15557
rect 2333 15489 2369 15523
rect 2333 15455 2334 15489
rect 2368 15455 2369 15489
rect 2333 15421 2369 15455
rect 2333 15387 2334 15421
rect 2368 15387 2369 15421
rect 2333 15353 2369 15387
rect 2333 15319 2334 15353
rect 2368 15319 2369 15353
rect 2333 15285 2369 15319
rect 2333 15251 2334 15285
rect 2368 15251 2369 15285
rect 2333 15217 2369 15251
rect 2333 15183 2334 15217
rect 2368 15183 2369 15217
rect 2333 15149 2369 15183
rect 2333 15115 2334 15149
rect 2368 15115 2369 15149
rect 2333 15081 2369 15115
rect 2333 15047 2334 15081
rect 2368 15047 2369 15081
rect 2333 15013 2369 15047
rect 2333 14979 2334 15013
rect 2368 14979 2369 15013
rect 2333 14945 2369 14979
rect 2333 14911 2334 14945
rect 2368 14911 2369 14945
rect 2333 14877 2369 14911
rect 2333 14843 2334 14877
rect 2368 14843 2369 14877
rect 2333 14809 2369 14843
rect 2333 14775 2334 14809
rect 2368 14775 2369 14809
rect 2333 14741 2369 14775
rect 2333 14707 2334 14741
rect 2368 14707 2369 14741
rect 2333 14673 2369 14707
rect 2333 14639 2334 14673
rect 2368 14639 2369 14673
rect 2333 14605 2369 14639
rect 2333 14571 2334 14605
rect 2368 14571 2369 14605
rect 2333 14537 2369 14571
rect 2333 14503 2334 14537
rect 2368 14503 2369 14537
rect 2333 14469 2369 14503
rect 2333 14435 2334 14469
rect 2368 14435 2369 14469
rect 2333 14401 2369 14435
rect 2333 14367 2334 14401
rect 2368 14367 2369 14401
rect 2333 14333 2369 14367
rect 2333 14299 2334 14333
rect 2368 14299 2369 14333
rect 2333 14265 2369 14299
rect 2333 14231 2334 14265
rect 2368 14231 2369 14265
rect 2333 14197 2369 14231
rect 2333 14163 2334 14197
rect 2368 14163 2369 14197
rect 2333 14129 2369 14163
rect 2333 14095 2334 14129
rect 2368 14095 2369 14129
rect 2333 14061 2369 14095
rect 2333 14027 2334 14061
rect 2368 14027 2369 14061
rect 2333 13993 2369 14027
rect 2333 13959 2334 13993
rect 2368 13959 2369 13993
rect 2333 13925 2369 13959
rect 2333 13891 2334 13925
rect 2368 13891 2369 13925
rect 2333 13857 2369 13891
rect 2333 13823 2334 13857
rect 2368 13823 2369 13857
rect 2333 13789 2369 13823
rect 2333 13755 2334 13789
rect 2368 13755 2369 13789
rect 2333 13721 2369 13755
rect 2333 13687 2334 13721
rect 2368 13687 2369 13721
rect 2333 13653 2369 13687
rect 2333 13619 2334 13653
rect 2368 13619 2369 13653
rect 2333 13585 2369 13619
rect 2333 13551 2334 13585
rect 2368 13551 2369 13585
rect 2333 13517 2369 13551
rect 2333 13483 2334 13517
rect 2368 13483 2369 13517
rect 2333 13449 2369 13483
rect 2333 13415 2334 13449
rect 2368 13415 2369 13449
rect 2333 13381 2369 13415
rect 2333 13347 2334 13381
rect 2368 13347 2369 13381
rect 2333 13313 2369 13347
rect 2333 13279 2334 13313
rect 2368 13279 2369 13313
rect 2333 13245 2369 13279
rect 2333 13211 2334 13245
rect 2368 13211 2369 13245
rect 2333 13177 2369 13211
rect 2333 13143 2334 13177
rect 2368 13143 2369 13177
rect 2333 13109 2369 13143
rect 2333 13075 2334 13109
rect 2368 13075 2369 13109
rect 2333 13041 2369 13075
rect 2333 13007 2334 13041
rect 2368 13007 2369 13041
rect 2333 12973 2369 13007
rect 2333 12939 2334 12973
rect 2368 12939 2369 12973
rect 2333 12905 2369 12939
rect 2333 12871 2334 12905
rect 2368 12871 2369 12905
rect 2333 12837 2369 12871
rect 2333 12803 2334 12837
rect 2368 12803 2369 12837
rect 2333 12769 2369 12803
rect 2333 12735 2334 12769
rect 2368 12735 2369 12769
rect 2333 12701 2369 12735
rect 2333 12667 2334 12701
rect 2368 12667 2369 12701
rect 2333 12633 2369 12667
rect 2333 12599 2334 12633
rect 2368 12599 2369 12633
rect 2333 12565 2369 12599
rect 2333 12531 2334 12565
rect 2368 12531 2369 12565
rect 2333 12497 2369 12531
rect 2333 12463 2334 12497
rect 2368 12463 2369 12497
rect 2333 12429 2369 12463
rect 2333 12395 2334 12429
rect 2368 12395 2369 12429
rect 2333 12361 2369 12395
rect 2333 12327 2334 12361
rect 2368 12327 2369 12361
rect 2333 12293 2369 12327
rect 2333 12259 2334 12293
rect 2368 12259 2369 12293
rect 2333 12225 2369 12259
rect 2333 12191 2334 12225
rect 2368 12191 2369 12225
rect 2333 12157 2369 12191
rect 2333 12123 2334 12157
rect 2368 12123 2369 12157
rect 2333 12089 2369 12123
rect 2333 12055 2334 12089
rect 2368 12055 2369 12089
rect 2333 12021 2369 12055
rect 2333 11987 2334 12021
rect 2368 11987 2369 12021
rect 2333 11953 2369 11987
rect 2333 11919 2334 11953
rect 2368 11919 2369 11953
rect 2333 11885 2369 11919
rect 2333 11851 2334 11885
rect 2368 11851 2369 11885
rect 2333 11817 2369 11851
rect 2333 11783 2334 11817
rect 2368 11783 2369 11817
rect 2333 11749 2369 11783
rect 2333 11715 2334 11749
rect 2368 11715 2369 11749
rect 2333 11681 2369 11715
rect 2333 11647 2334 11681
rect 2368 11647 2369 11681
rect 2333 11613 2369 11647
rect 2333 11579 2334 11613
rect 2368 11579 2369 11613
rect 2333 11545 2369 11579
rect 2333 11511 2334 11545
rect 2368 11511 2369 11545
rect 2333 11477 2369 11511
rect 2333 11443 2334 11477
rect 2368 11443 2369 11477
rect 2333 11409 2369 11443
rect 2333 11375 2334 11409
rect 2368 11375 2369 11409
rect 2333 11341 2369 11375
rect 2333 11307 2334 11341
rect 2368 11307 2369 11341
rect 2333 11273 2369 11307
rect 2333 11239 2334 11273
rect 2368 11239 2369 11273
rect 2333 11205 2369 11239
rect 2333 11171 2334 11205
rect 2368 11171 2369 11205
rect 2333 11137 2369 11171
rect 2333 11103 2334 11137
rect 2368 11103 2369 11137
rect 2333 11079 2369 11103
rect 2333 11069 6889 11079
rect 2333 11035 2334 11069
rect 2368 11043 6889 11069
rect 2368 11035 2369 11043
rect 2333 11001 2369 11035
rect 2333 10967 2334 11001
rect 2368 10967 2369 11001
rect 2333 10933 2369 10967
rect 2333 10899 2334 10933
rect 2368 10899 2369 10933
rect 2333 10865 2369 10899
rect 2333 10831 2334 10865
rect 2368 10831 2369 10865
rect 2333 10797 2369 10831
rect 2333 10763 2334 10797
rect 2368 10763 2369 10797
rect 2333 10729 2369 10763
rect 2333 10695 2334 10729
rect 2368 10695 2369 10729
rect 2333 10661 2369 10695
rect 2333 10627 2334 10661
rect 2368 10627 2369 10661
rect 2333 10593 2369 10627
rect 2333 10559 2334 10593
rect 2368 10559 2369 10593
rect 2333 10525 2369 10559
rect 2333 10491 2334 10525
rect 2368 10491 2369 10525
rect 2333 10457 2369 10491
rect 2333 10423 2334 10457
rect 2368 10423 2369 10457
rect 2333 10389 2369 10423
rect 2333 10355 2334 10389
rect 2368 10355 2369 10389
rect 2333 10321 2369 10355
rect 2333 10287 2334 10321
rect 2368 10287 2369 10321
rect 2333 10253 2369 10287
rect 2333 10219 2334 10253
rect 2368 10219 2369 10253
rect 2333 10185 2369 10219
rect 2333 10151 2334 10185
rect 2368 10151 2369 10185
rect 2333 10117 2369 10151
rect 2333 10083 2334 10117
rect 2368 10083 2369 10117
rect 2333 10049 2369 10083
rect 2333 10015 2334 10049
rect 2368 10015 2369 10049
rect 2333 9981 2369 10015
rect 2333 9947 2334 9981
rect 2368 9947 2369 9981
rect 2333 9913 2369 9947
rect 2333 9879 2334 9913
rect 2368 9879 2369 9913
rect 2333 9845 2369 9879
rect 2333 9811 2334 9845
rect 2368 9811 2369 9845
rect 2333 9777 2369 9811
rect 2333 9743 2334 9777
rect 2368 9743 2369 9777
rect 2333 9709 2369 9743
rect 2333 9675 2334 9709
rect 2368 9675 2369 9709
rect 2333 9641 2369 9675
rect 2333 9607 2334 9641
rect 2368 9607 2369 9641
rect 2333 9573 2369 9607
rect 2333 9539 2334 9573
rect 2368 9539 2369 9573
rect 2333 9505 2369 9539
rect 2333 9471 2334 9505
rect 2368 9471 2369 9505
rect 2333 9437 2369 9471
rect 2333 9403 2334 9437
rect 2368 9403 2369 9437
rect 2333 9369 2369 9403
rect 2333 9335 2334 9369
rect 2368 9335 2369 9369
rect 2333 9301 2369 9335
rect 2333 9267 2334 9301
rect 2368 9267 2369 9301
rect 2333 9233 2369 9267
rect 2333 9199 2334 9233
rect 2368 9199 2369 9233
rect 2333 9165 2369 9199
rect 2333 9131 2334 9165
rect 2368 9131 2369 9165
rect 2333 9097 2369 9131
rect 2333 9063 2334 9097
rect 2368 9063 2369 9097
rect 2333 9029 2369 9063
rect 2333 8995 2334 9029
rect 2368 8995 2369 9029
rect 2333 8961 2369 8995
rect 2333 8927 2334 8961
rect 2368 8927 2369 8961
rect 2333 8893 2369 8927
rect 2333 8859 2334 8893
rect 2368 8859 2369 8893
rect 2333 8825 2369 8859
rect 2333 8791 2334 8825
rect 2368 8791 2369 8825
rect 2333 8757 2369 8791
rect 2333 8723 2334 8757
rect 2368 8723 2369 8757
rect 2333 8689 2369 8723
rect 2333 8655 2334 8689
rect 2368 8655 2369 8689
rect 2333 8621 2369 8655
rect 2333 8587 2334 8621
rect 2368 8587 2369 8621
rect 2333 8553 2369 8587
rect 2333 8519 2334 8553
rect 2368 8519 2369 8553
rect 2333 8485 2369 8519
rect 2333 8451 2334 8485
rect 2368 8451 2369 8485
rect 2333 8417 2369 8451
rect 2333 8383 2334 8417
rect 2368 8383 2369 8417
rect 2333 8349 2369 8383
rect 2333 8315 2334 8349
rect 2368 8315 2369 8349
rect 2333 8281 2369 8315
rect 2333 8247 2334 8281
rect 2368 8247 2369 8281
rect 2333 8213 2369 8247
rect 2333 8179 2334 8213
rect 2368 8179 2369 8213
rect 2333 8145 2369 8179
rect 2333 8111 2334 8145
rect 2368 8111 2369 8145
rect 2333 8077 2369 8111
rect 2333 8043 2334 8077
rect 2368 8043 2369 8077
rect 2333 8009 2369 8043
rect 2333 7975 2334 8009
rect 2368 7975 2369 8009
rect 2333 7941 2369 7975
rect 2333 7907 2334 7941
rect 2368 7907 2369 7941
rect 2333 7873 2369 7907
rect 2333 7839 2334 7873
rect 2368 7839 2369 7873
rect 2333 7805 2369 7839
rect 2333 7771 2334 7805
rect 2368 7771 2369 7805
rect 2333 7737 2369 7771
rect 2333 7703 2334 7737
rect 2368 7703 2369 7737
rect 2333 7669 2369 7703
rect 2333 7635 2334 7669
rect 2368 7635 2369 7669
rect 2333 7601 2369 7635
rect 2333 7567 2334 7601
rect 2368 7567 2369 7601
rect 2333 7533 2369 7567
rect 2333 7499 2334 7533
rect 2368 7499 2369 7533
rect 2333 7465 2369 7499
rect 2333 7431 2334 7465
rect 2368 7431 2369 7465
rect 2333 7397 2369 7431
rect 2333 7363 2334 7397
rect 2368 7363 2369 7397
rect 2333 7329 2369 7363
rect 2333 7295 2334 7329
rect 2368 7295 2369 7329
rect 2333 7261 2369 7295
rect 2333 7227 2334 7261
rect 2368 7227 2369 7261
rect 2333 7193 2369 7227
rect 2333 7159 2334 7193
rect 2368 7159 2369 7193
rect 2333 7125 2369 7159
rect 2333 7091 2334 7125
rect 2368 7091 2369 7125
rect 2333 7057 2369 7091
rect 2333 7023 2334 7057
rect 2368 7023 2369 7057
rect 2333 6989 2369 7023
rect 2333 6955 2334 6989
rect 2368 6955 2369 6989
rect 2333 6921 2369 6955
rect 2333 6887 2334 6921
rect 2368 6887 2369 6921
rect 2333 6853 2369 6887
rect 2333 6819 2334 6853
rect 2368 6819 2369 6853
rect 2333 6785 2369 6819
rect 2333 6751 2334 6785
rect 2368 6751 2369 6785
rect 2333 6717 2369 6751
rect 2333 6683 2334 6717
rect 2368 6683 2369 6717
rect 2333 6649 2369 6683
rect 2333 6615 2334 6649
rect 2368 6615 2369 6649
rect 2333 6581 2369 6615
rect 2333 6547 2334 6581
rect 2368 6547 2369 6581
rect 2333 6513 2369 6547
rect 2333 6479 2334 6513
rect 2368 6479 2369 6513
rect 2333 6445 2369 6479
rect 2333 6411 2334 6445
rect 2368 6411 2369 6445
rect 2333 6377 2369 6411
rect 2333 6343 2334 6377
rect 2368 6343 2369 6377
rect 2333 6309 2369 6343
rect 2333 6275 2334 6309
rect 2368 6275 2369 6309
rect 2333 6241 2369 6275
rect 2333 6207 2334 6241
rect 2368 6207 2369 6241
rect 2553 11009 2589 11043
rect 2553 10975 2554 11009
rect 2588 10975 2589 11009
rect 2553 10941 2589 10975
rect 2553 10907 2554 10941
rect 2588 10907 2589 10941
rect 2553 10873 2589 10907
rect 6853 10995 6889 11043
rect 6853 10961 6854 10995
rect 6888 10961 6889 10995
rect 6853 10927 6889 10961
rect 6853 10893 6854 10927
rect 6888 10893 6889 10927
rect 2553 10839 2554 10873
rect 2588 10839 2589 10873
rect 2553 10805 2589 10839
rect 2553 10771 2554 10805
rect 2588 10771 2589 10805
rect 2553 10737 2589 10771
rect 2553 10703 2554 10737
rect 2588 10703 2589 10737
rect 2553 10669 2589 10703
rect 2553 10635 2554 10669
rect 2588 10635 2589 10669
rect 2553 10601 2589 10635
rect 2553 10567 2554 10601
rect 2588 10567 2589 10601
rect 2553 10533 2589 10567
rect 2553 10499 2554 10533
rect 2588 10499 2589 10533
rect 2553 10465 2589 10499
rect 2553 10431 2554 10465
rect 2588 10431 2589 10465
rect 2553 10397 2589 10431
rect 2553 10363 2554 10397
rect 2588 10363 2589 10397
rect 2553 10329 2589 10363
rect 2553 10295 2554 10329
rect 2588 10295 2589 10329
rect 2553 10261 2589 10295
rect 2553 10227 2554 10261
rect 2588 10227 2589 10261
rect 2553 10193 2589 10227
rect 2553 10159 2554 10193
rect 2588 10159 2589 10193
rect 2553 10125 2589 10159
rect 2553 10091 2554 10125
rect 2588 10091 2589 10125
rect 2553 10057 2589 10091
rect 2553 10023 2554 10057
rect 2588 10023 2589 10057
rect 2553 9989 2589 10023
rect 2553 9955 2554 9989
rect 2588 9955 2589 9989
rect 2553 9921 2589 9955
rect 2553 9887 2554 9921
rect 2588 9887 2589 9921
rect 2553 9853 2589 9887
rect 2553 9819 2554 9853
rect 2588 9819 2589 9853
rect 2553 9785 2589 9819
rect 2553 9751 2554 9785
rect 2588 9751 2589 9785
rect 2553 9717 2589 9751
rect 2553 9683 2554 9717
rect 2588 9683 2589 9717
rect 2553 9649 2589 9683
rect 2553 9615 2554 9649
rect 2588 9615 2589 9649
rect 2553 9581 2589 9615
rect 2553 9547 2554 9581
rect 2588 9547 2589 9581
rect 2553 9513 2589 9547
rect 2553 9479 2554 9513
rect 2588 9479 2589 9513
rect 2553 9445 2589 9479
rect 2553 9411 2554 9445
rect 2588 9411 2589 9445
rect 2553 9377 2589 9411
rect 2553 9343 2554 9377
rect 2588 9343 2589 9377
rect 2553 9309 2589 9343
rect 2553 9275 2554 9309
rect 2588 9275 2589 9309
rect 2553 9241 2589 9275
rect 2553 9207 2554 9241
rect 2588 9207 2589 9241
rect 2553 9173 2589 9207
rect 2553 9139 2554 9173
rect 2588 9139 2589 9173
rect 2553 9105 2589 9139
rect 2553 9071 2554 9105
rect 2588 9071 2589 9105
rect 2553 9037 2589 9071
rect 2553 9003 2554 9037
rect 2588 9003 2589 9037
rect 2553 8969 2589 9003
rect 2553 8935 2554 8969
rect 2588 8935 2589 8969
rect 2553 8901 2589 8935
rect 2553 8867 2554 8901
rect 2588 8867 2589 8901
rect 2553 8833 2589 8867
rect 2553 8799 2554 8833
rect 2588 8799 2589 8833
rect 2553 8765 2589 8799
rect 2553 8731 2554 8765
rect 2588 8731 2589 8765
rect 2553 8697 2589 8731
rect 2553 8663 2554 8697
rect 2588 8663 2589 8697
rect 2553 8629 2589 8663
rect 2553 8595 2554 8629
rect 2588 8595 2589 8629
rect 2553 8561 2589 8595
rect 2553 8527 2554 8561
rect 2588 8527 2589 8561
rect 2553 8493 2589 8527
rect 2553 8459 2554 8493
rect 2588 8459 2589 8493
rect 2553 8425 2589 8459
rect 2553 8391 2554 8425
rect 2588 8391 2589 8425
rect 2553 8357 2589 8391
rect 2553 8323 2554 8357
rect 2588 8323 2589 8357
rect 2553 8289 2589 8323
rect 2553 8255 2554 8289
rect 2588 8255 2589 8289
rect 2553 8221 2589 8255
rect 2553 8187 2554 8221
rect 2588 8187 2589 8221
rect 2553 8153 2589 8187
rect 2553 8119 2554 8153
rect 2588 8119 2589 8153
rect 2553 8085 2589 8119
rect 2553 8051 2554 8085
rect 2588 8051 2589 8085
rect 2553 8017 2589 8051
rect 2553 7983 2554 8017
rect 2588 7983 2589 8017
rect 2553 7949 2589 7983
rect 2553 7915 2554 7949
rect 2588 7915 2589 7949
rect 2553 7881 2589 7915
rect 2553 7847 2554 7881
rect 2588 7847 2589 7881
rect 2553 7813 2589 7847
rect 2553 7779 2554 7813
rect 2588 7779 2589 7813
rect 2553 7745 2589 7779
rect 2553 7711 2554 7745
rect 2588 7711 2589 7745
rect 2553 7677 2589 7711
rect 2553 7643 2554 7677
rect 2588 7643 2589 7677
rect 2553 7609 2589 7643
rect 2553 7575 2554 7609
rect 2588 7575 2589 7609
rect 2553 7541 2589 7575
rect 2553 7507 2554 7541
rect 2588 7507 2589 7541
rect 2553 7473 2589 7507
rect 2553 7439 2554 7473
rect 2588 7439 2589 7473
rect 2553 7405 2589 7439
rect 2553 7371 2554 7405
rect 2588 7371 2589 7405
rect 2553 7337 2589 7371
rect 2553 7303 2554 7337
rect 2588 7303 2589 7337
rect 2553 7269 2589 7303
rect 2553 7235 2554 7269
rect 2588 7235 2589 7269
rect 2553 7201 2589 7235
rect 2553 7167 2554 7201
rect 2588 7167 2589 7201
rect 2553 7133 2589 7167
rect 2553 7099 2554 7133
rect 2588 7099 2589 7133
rect 2553 7065 2589 7099
rect 2553 7031 2554 7065
rect 2588 7031 2589 7065
rect 2553 6997 2589 7031
rect 2553 6963 2554 6997
rect 2588 6963 2589 6997
rect 2553 6929 2589 6963
rect 2553 6895 2554 6929
rect 2588 6895 2589 6929
rect 2553 6861 2589 6895
rect 2553 6827 2554 6861
rect 2588 6827 2589 6861
rect 2553 6793 2589 6827
rect 2553 6759 2554 6793
rect 2588 6759 2589 6793
rect 2553 6725 2589 6759
rect 2553 6691 2554 6725
rect 2588 6691 2589 6725
rect 2553 6657 2589 6691
rect 2553 6623 2554 6657
rect 2588 6623 2589 6657
rect 2553 6589 2589 6623
rect 2553 6555 2554 6589
rect 2588 6555 2589 6589
rect 2553 6521 2589 6555
rect 2553 6487 2554 6521
rect 2588 6487 2589 6521
rect 2553 6453 2589 6487
rect 2553 6419 2554 6453
rect 2588 6419 2589 6453
rect 6853 10859 6889 10893
rect 6853 10825 6854 10859
rect 6888 10825 6889 10859
rect 6853 10791 6889 10825
rect 6853 10757 6854 10791
rect 6888 10757 6889 10791
rect 6853 10723 6889 10757
rect 6853 10689 6854 10723
rect 6888 10689 6889 10723
rect 6853 10655 6889 10689
rect 6853 10621 6854 10655
rect 6888 10621 6889 10655
rect 6853 10587 6889 10621
rect 6853 10553 6854 10587
rect 6888 10553 6889 10587
rect 6853 10519 6889 10553
rect 6853 10485 6854 10519
rect 6888 10485 6889 10519
rect 6853 10451 6889 10485
rect 6853 10417 6854 10451
rect 6888 10417 6889 10451
rect 6853 10383 6889 10417
rect 6853 10349 6854 10383
rect 6888 10349 6889 10383
rect 6853 10315 6889 10349
rect 6853 10281 6854 10315
rect 6888 10281 6889 10315
rect 6853 10247 6889 10281
rect 6853 10213 6854 10247
rect 6888 10213 6889 10247
rect 6853 10179 6889 10213
rect 6853 10145 6854 10179
rect 6888 10145 6889 10179
rect 6853 10111 6889 10145
rect 6853 10077 6854 10111
rect 6888 10077 6889 10111
rect 6853 10043 6889 10077
rect 6853 10009 6854 10043
rect 6888 10009 6889 10043
rect 6853 9975 6889 10009
rect 6853 9941 6854 9975
rect 6888 9941 6889 9975
rect 6853 9907 6889 9941
rect 6853 9873 6854 9907
rect 6888 9873 6889 9907
rect 6853 9839 6889 9873
rect 6853 9805 6854 9839
rect 6888 9805 6889 9839
rect 6853 9771 6889 9805
rect 6853 9737 6854 9771
rect 6888 9737 6889 9771
rect 6853 9703 6889 9737
rect 6853 9669 6854 9703
rect 6888 9669 6889 9703
rect 6853 9635 6889 9669
rect 6853 9601 6854 9635
rect 6888 9601 6889 9635
rect 6853 9567 6889 9601
rect 6853 9533 6854 9567
rect 6888 9533 6889 9567
rect 6853 9499 6889 9533
rect 6853 9465 6854 9499
rect 6888 9465 6889 9499
rect 6853 9431 6889 9465
rect 6853 9397 6854 9431
rect 6888 9397 6889 9431
rect 6853 9363 6889 9397
rect 6853 9329 6854 9363
rect 6888 9329 6889 9363
rect 6853 9295 6889 9329
rect 6853 9261 6854 9295
rect 6888 9261 6889 9295
rect 6853 9227 6889 9261
rect 6853 9193 6854 9227
rect 6888 9193 6889 9227
rect 6853 9159 6889 9193
rect 6853 9125 6854 9159
rect 6888 9125 6889 9159
rect 6853 9091 6889 9125
rect 6853 9057 6854 9091
rect 6888 9057 6889 9091
rect 6853 9023 6889 9057
rect 6853 8989 6854 9023
rect 6888 8989 6889 9023
rect 6853 8955 6889 8989
rect 6853 8921 6854 8955
rect 6888 8921 6889 8955
rect 6853 8887 6889 8921
rect 6853 8853 6854 8887
rect 6888 8853 6889 8887
rect 6853 8819 6889 8853
rect 6853 8785 6854 8819
rect 6888 8785 6889 8819
rect 6853 8751 6889 8785
rect 6853 8717 6854 8751
rect 6888 8717 6889 8751
rect 6853 8683 6889 8717
rect 6853 8649 6854 8683
rect 6888 8649 6889 8683
rect 6853 8615 6889 8649
rect 6853 8581 6854 8615
rect 6888 8581 6889 8615
rect 6853 8547 6889 8581
rect 6853 8513 6854 8547
rect 6888 8513 6889 8547
rect 6853 8479 6889 8513
rect 6853 8445 6854 8479
rect 6888 8445 6889 8479
rect 6853 8411 6889 8445
rect 6853 8377 6854 8411
rect 6888 8377 6889 8411
rect 6853 8343 6889 8377
rect 6853 8309 6854 8343
rect 6888 8309 6889 8343
rect 6853 8275 6889 8309
rect 6853 8241 6854 8275
rect 6888 8241 6889 8275
rect 6853 8207 6889 8241
rect 6853 8173 6854 8207
rect 6888 8173 6889 8207
rect 6853 8139 6889 8173
rect 6853 8105 6854 8139
rect 6888 8105 6889 8139
rect 6853 8071 6889 8105
rect 6853 8037 6854 8071
rect 6888 8037 6889 8071
rect 6853 8003 6889 8037
rect 6853 7969 6854 8003
rect 6888 7969 6889 8003
rect 6853 7935 6889 7969
rect 6853 7901 6854 7935
rect 6888 7901 6889 7935
rect 6853 7867 6889 7901
rect 6853 7833 6854 7867
rect 6888 7833 6889 7867
rect 6853 7799 6889 7833
rect 6853 7765 6854 7799
rect 6888 7765 6889 7799
rect 6853 7731 6889 7765
rect 6853 7697 6854 7731
rect 6888 7697 6889 7731
rect 6853 7663 6889 7697
rect 6853 7629 6854 7663
rect 6888 7629 6889 7663
rect 6853 7595 6889 7629
rect 6853 7561 6854 7595
rect 6888 7561 6889 7595
rect 6853 7527 6889 7561
rect 6853 7493 6854 7527
rect 6888 7493 6889 7527
rect 6853 7459 6889 7493
rect 6853 7425 6854 7459
rect 6888 7425 6889 7459
rect 6853 7391 6889 7425
rect 6853 7357 6854 7391
rect 6888 7357 6889 7391
rect 6853 7323 6889 7357
rect 6853 7289 6854 7323
rect 6888 7289 6889 7323
rect 6853 7255 6889 7289
rect 6853 7221 6854 7255
rect 6888 7221 6889 7255
rect 6853 7187 6889 7221
rect 6853 7153 6854 7187
rect 6888 7153 6889 7187
rect 6853 7119 6889 7153
rect 6853 7085 6854 7119
rect 6888 7085 6889 7119
rect 6853 7051 6889 7085
rect 6853 7017 6854 7051
rect 6888 7017 6889 7051
rect 6853 6983 6889 7017
rect 6853 6949 6854 6983
rect 6888 6949 6889 6983
rect 6853 6915 6889 6949
rect 6853 6881 6854 6915
rect 6888 6881 6889 6915
rect 6853 6847 6889 6881
rect 6853 6813 6854 6847
rect 6888 6813 6889 6847
rect 6853 6779 6889 6813
rect 6853 6745 6854 6779
rect 6888 6745 6889 6779
rect 6853 6711 6889 6745
rect 6853 6677 6854 6711
rect 6888 6677 6889 6711
rect 6853 6643 6889 6677
rect 6853 6609 6854 6643
rect 6888 6609 6889 6643
rect 6853 6575 6889 6609
rect 6853 6541 6854 6575
rect 6888 6541 6889 6575
rect 6853 6507 6889 6541
rect 6853 6473 6854 6507
rect 6888 6473 6889 6507
rect 6853 6439 6889 6473
rect 2553 6385 2589 6419
rect 2553 6351 2554 6385
rect 2588 6351 2589 6385
rect 2553 6271 2589 6351
rect 6853 6405 6854 6439
rect 6888 6405 6889 6439
rect 6853 6371 6889 6405
rect 6853 6337 6854 6371
rect 6888 6337 6889 6371
rect 6853 6303 6889 6337
rect 6853 6271 6854 6303
rect 2553 6270 6854 6271
rect 2553 6236 2587 6270
rect 2621 6236 2655 6270
rect 2689 6236 2723 6270
rect 2757 6236 2791 6270
rect 2825 6236 2859 6270
rect 2893 6236 2927 6270
rect 2961 6236 2995 6270
rect 3029 6236 3063 6270
rect 3097 6236 3131 6270
rect 3165 6236 3199 6270
rect 3233 6236 3267 6270
rect 3301 6236 3335 6270
rect 3369 6236 3403 6270
rect 3437 6236 3471 6270
rect 3505 6236 3539 6270
rect 3573 6236 3607 6270
rect 3641 6236 3675 6270
rect 3709 6236 3743 6270
rect 3777 6236 3811 6270
rect 3845 6236 3879 6270
rect 3913 6236 3947 6270
rect 3981 6236 4015 6270
rect 4049 6236 4083 6270
rect 4117 6236 4151 6270
rect 4185 6236 4219 6270
rect 4253 6236 4287 6270
rect 4321 6236 4355 6270
rect 4389 6236 4423 6270
rect 4457 6236 4491 6270
rect 4525 6236 4559 6270
rect 4593 6236 4627 6270
rect 4661 6236 4695 6270
rect 4729 6236 4763 6270
rect 4797 6236 4831 6270
rect 4865 6236 4899 6270
rect 4933 6236 4967 6270
rect 5001 6236 5035 6270
rect 5069 6236 5103 6270
rect 5137 6236 5171 6270
rect 5205 6236 5239 6270
rect 5273 6236 5307 6270
rect 5341 6236 5375 6270
rect 5409 6236 5443 6270
rect 5477 6236 5511 6270
rect 5545 6236 5579 6270
rect 5613 6236 5647 6270
rect 5681 6236 5715 6270
rect 5749 6236 5783 6270
rect 5817 6236 5851 6270
rect 5885 6236 5919 6270
rect 5953 6236 5987 6270
rect 6021 6236 6055 6270
rect 6089 6236 6123 6270
rect 6157 6236 6191 6270
rect 6225 6236 6259 6270
rect 6293 6236 6327 6270
rect 6361 6236 6395 6270
rect 6429 6236 6463 6270
rect 6497 6236 6531 6270
rect 6565 6236 6599 6270
rect 6633 6236 6667 6270
rect 6701 6236 6735 6270
rect 6769 6269 6854 6270
rect 6888 6269 6889 6303
rect 6769 6236 6889 6269
rect 2553 6235 6889 6236
rect 2333 6173 2369 6207
rect 2333 6139 2334 6173
rect 2368 6139 2369 6173
rect 2333 6105 2369 6139
rect 6854 6211 6888 6235
rect 6854 6139 6888 6177
rect 2333 6071 2357 6105
rect 2391 6071 2426 6105
rect 2460 6071 2495 6105
rect 2529 6071 2564 6105
rect 2598 6071 2633 6105
rect 2667 6071 2702 6105
rect 2736 6071 2771 6105
rect 2805 6071 2840 6105
rect 2874 6071 2909 6105
rect 2943 6071 2978 6105
rect 3012 6071 3047 6105
rect 3081 6071 3116 6105
rect 3150 6071 3185 6105
rect 3219 6071 3254 6105
rect 3288 6071 3323 6105
rect 3357 6071 3392 6105
rect 3426 6071 3461 6105
rect 3495 6071 3530 6105
rect 3564 6071 3599 6105
rect 3633 6071 3668 6105
rect 3702 6071 3737 6105
rect 3771 6071 3806 6105
rect 3840 6071 3875 6105
rect 3909 6071 3944 6105
rect 3978 6071 4013 6105
rect 4047 6071 4082 6105
rect 4116 6071 4151 6105
rect 4185 6071 4220 6105
rect 4254 6071 4289 6105
rect 4323 6071 4358 6105
rect 4392 6071 4427 6105
rect 4461 6071 4496 6105
rect 4530 6071 4565 6105
rect 4599 6071 4634 6105
rect 4668 6071 4703 6105
rect 4737 6071 4772 6105
rect 4806 6071 4841 6105
rect 4875 6071 4910 6105
rect 4944 6071 4979 6105
rect 5013 6071 5048 6105
rect 5082 6071 5117 6105
rect 5151 6071 5186 6105
rect 5220 6071 5255 6105
rect 5289 6071 5324 6105
rect 5358 6071 5392 6105
rect 5426 6071 5460 6105
rect 5494 6071 5528 6105
rect 5562 6071 5596 6105
rect 5630 6071 5664 6105
rect 5698 6071 5732 6105
rect 5766 6071 5800 6105
rect 5834 6071 5868 6105
rect 5902 6071 5936 6105
rect 5970 6071 6004 6105
rect 6038 6071 6072 6105
rect 6106 6071 6140 6105
rect 6174 6071 6208 6105
rect 6242 6071 6276 6105
rect 6310 6071 6344 6105
rect 6378 6071 6412 6105
rect 6446 6071 6480 6105
rect 6514 6071 6548 6105
rect 6582 6071 6616 6105
rect 6650 6071 6684 6105
rect 6718 6071 6752 6105
rect 6786 6071 6888 6105
rect 3341 815 3377 899
rect 3341 781 3342 815
rect 3376 781 3377 815
rect 3341 747 3377 781
rect 3341 713 3342 747
rect 3376 713 3377 747
rect 3341 679 3377 713
rect 3341 645 3342 679
rect 3376 645 3377 679
rect 3341 611 3377 645
rect 3341 577 3342 611
rect 3376 577 3377 611
rect 3341 543 3377 577
rect 3341 509 3342 543
rect 3376 509 3377 543
rect 3341 475 3377 509
rect 3341 441 3342 475
rect 3376 441 3377 475
rect 3341 407 3377 441
rect 3341 373 3342 407
rect 3376 373 3377 407
rect 3341 339 3377 373
rect 3341 305 3342 339
rect 3376 305 3377 339
rect 3341 271 3377 305
rect 3341 237 3342 271
rect 3376 237 3377 271
rect 3341 203 3377 237
rect 3341 169 3342 203
rect 3376 169 3377 203
rect 3341 135 3377 169
rect 3341 103 3342 135
rect 742 102 3342 103
rect 742 69 887 102
rect 742 35 743 69
rect 777 68 887 69
rect 921 68 955 102
rect 989 68 1023 102
rect 1057 68 1091 102
rect 1125 68 1159 102
rect 1193 68 1227 102
rect 1261 68 1295 102
rect 1329 68 1363 102
rect 1397 68 1431 102
rect 1465 68 1499 102
rect 1533 68 1567 102
rect 1601 68 1635 102
rect 1669 68 1703 102
rect 1737 68 1771 102
rect 1805 68 1839 102
rect 1873 68 1907 102
rect 1941 68 1975 102
rect 2009 68 2043 102
rect 2077 68 2111 102
rect 2145 68 2179 102
rect 2213 68 2247 102
rect 2281 68 2315 102
rect 2349 68 2383 102
rect 2417 68 2451 102
rect 2485 68 2519 102
rect 2553 68 2587 102
rect 2621 68 2655 102
rect 2689 68 2723 102
rect 2757 68 2791 102
rect 2825 68 2859 102
rect 2893 68 2927 102
rect 2961 68 2995 102
rect 3029 68 3063 102
rect 3097 68 3131 102
rect 3165 68 3199 102
rect 3233 68 3267 102
rect 3301 101 3342 102
rect 3376 101 3377 135
rect 3301 78 3377 101
rect 3301 68 3640 78
rect 777 67 3640 68
rect 777 35 778 67
rect 3341 44 3640 67
rect 742 1 778 35
rect 742 -33 743 1
rect 777 -33 778 1
rect 742 -67 778 -33
rect 742 -101 743 -67
rect 777 -101 778 -67
rect 742 -135 778 -101
rect 742 -169 743 -135
rect 777 -169 778 -135
rect 742 -203 778 -169
rect 742 -237 743 -203
rect 777 -237 778 -203
rect 742 -271 778 -237
rect 3604 8 3640 44
rect 3604 -26 3605 8
rect 3639 -26 3640 8
rect 3604 -60 3640 -26
rect 3604 -94 3605 -60
rect 3639 -94 3640 -60
rect 3604 -128 3640 -94
rect 3604 -162 3605 -128
rect 3639 -162 3640 -128
rect 3604 -196 3640 -162
rect 3604 -230 3605 -196
rect 3639 -230 3640 -196
rect 742 -305 743 -271
rect 777 -305 778 -271
rect 742 -339 778 -305
rect 3604 -264 3640 -230
rect 3604 -298 3605 -264
rect 3639 -298 3640 -264
rect 3604 -332 3640 -298
rect 742 -373 743 -339
rect 777 -373 778 -339
rect 3604 -364 3605 -332
rect 742 -407 778 -373
rect 742 -441 743 -407
rect 777 -441 778 -407
rect 742 -475 778 -441
rect 742 -509 743 -475
rect 777 -509 778 -475
rect 742 -543 778 -509
rect 742 -577 743 -543
rect 777 -577 778 -543
rect 742 -628 778 -577
rect 1680 -365 3605 -364
rect 1680 -399 1714 -365
rect 1748 -399 1861 -365
rect 1895 -399 1929 -365
rect 1963 -399 1997 -365
rect 2031 -399 2065 -365
rect 2099 -399 2133 -365
rect 2167 -399 2201 -365
rect 2235 -399 2269 -365
rect 2303 -399 2337 -365
rect 2371 -399 2405 -365
rect 2439 -399 2473 -365
rect 2507 -399 2541 -365
rect 2575 -399 2609 -365
rect 2643 -399 2677 -365
rect 2711 -399 2745 -365
rect 2779 -399 2813 -365
rect 2847 -399 2881 -365
rect 2915 -399 2949 -365
rect 2983 -399 3017 -365
rect 3051 -399 3085 -365
rect 3119 -399 3153 -365
rect 3187 -399 3221 -365
rect 3255 -399 3289 -365
rect 3323 -399 3357 -365
rect 3391 -399 3425 -365
rect 3459 -399 3493 -365
rect 3527 -366 3605 -365
rect 3639 -366 3640 -332
rect 3527 -399 3640 -366
rect 1680 -400 3640 -399
rect 1680 -460 1716 -400
rect 1680 -494 1681 -460
rect 1715 -494 1716 -460
rect 1680 -528 1716 -494
rect 1680 -562 1681 -528
rect 1715 -562 1716 -528
rect 1680 -596 1716 -562
rect 1680 -628 1681 -596
rect 742 -629 1681 -628
rect 742 -663 776 -629
rect 810 -663 844 -629
rect 878 -663 912 -629
rect 946 -663 980 -629
rect 1014 -663 1048 -629
rect 1082 -663 1116 -629
rect 1150 -663 1184 -629
rect 1218 -663 1252 -629
rect 1286 -663 1320 -629
rect 1354 -663 1388 -629
rect 1422 -663 1456 -629
rect 1490 -663 1524 -629
rect 1558 -663 1592 -629
rect 1626 -630 1681 -629
rect 1715 -630 1716 -596
rect 1626 -663 1716 -630
rect 742 -664 1716 -663
<< psubdiffcont >>
rect 2149 -621 2183 -587
rect 2274 -588 2308 -554
rect 2342 -588 2376 -554
rect 2410 -588 2444 -554
rect 2478 -588 2512 -554
rect 2546 -588 2580 -554
rect 2614 -588 2648 -554
rect 2682 -588 2716 -554
rect 2750 -588 2784 -554
rect 2818 -588 2852 -554
rect 2886 -588 2920 -554
rect 2954 -588 2988 -554
rect 3022 -588 3056 -554
rect 3090 -588 3124 -554
rect 3158 -588 3192 -554
rect 3226 -588 3260 -554
rect 3294 -588 3328 -554
rect 3362 -588 3396 -554
rect 3430 -588 3464 -554
rect 2149 -689 2183 -655
rect 3463 -656 3497 -622
rect 2149 -757 2183 -723
rect 2149 -825 2183 -791
rect 2149 -893 2183 -859
rect 3463 -724 3497 -690
rect 3463 -792 3497 -758
rect 3463 -860 3497 -826
rect 3463 -928 3497 -894
rect 2182 -1029 2216 -995
rect 2250 -1029 2284 -995
rect 2318 -1029 2352 -995
rect 2386 -1029 2420 -995
rect 2454 -1029 2488 -995
rect 2522 -1029 2556 -995
rect 2590 -1029 2624 -995
rect 2658 -1029 2692 -995
rect 2726 -1029 2760 -995
rect 2794 -1029 2828 -995
rect 2862 -1029 2896 -995
rect 2930 -1029 2964 -995
rect 2998 -1029 3032 -995
rect 3066 -1029 3100 -995
rect 3134 -1029 3168 -995
rect 3202 -1029 3236 -995
rect 3270 -1029 3304 -995
rect 3338 -1029 3372 -995
rect 3463 -996 3497 -962
<< mvpsubdiffcont >>
rect 257 27613 291 27647
rect 344 27646 378 27680
rect 412 27646 446 27680
rect 480 27646 514 27680
rect 548 27646 582 27680
rect 616 27646 650 27680
rect 684 27646 718 27680
rect 752 27646 786 27680
rect 820 27646 854 27680
rect 888 27646 922 27680
rect 956 27646 990 27680
rect 1024 27646 1058 27680
rect 1092 27646 1126 27680
rect 1160 27646 1194 27680
rect 1228 27646 1262 27680
rect 1296 27646 1330 27680
rect 1364 27646 1398 27680
rect 1432 27646 1466 27680
rect 1500 27646 1534 27680
rect 1568 27646 1602 27680
rect 1636 27646 1670 27680
rect 1704 27646 1738 27680
rect 1772 27646 1806 27680
rect 1840 27646 1874 27680
rect 1908 27646 1942 27680
rect 1976 27646 2010 27680
rect 2044 27646 2078 27680
rect 2112 27646 2146 27680
rect 257 27545 291 27579
rect 257 27477 291 27511
rect 2145 27537 2179 27571
rect 257 27409 291 27443
rect 257 27341 291 27375
rect 257 27273 291 27307
rect 257 27205 291 27239
rect 257 27137 291 27171
rect 257 27069 291 27103
rect 257 27001 291 27035
rect 257 26933 291 26967
rect 257 26865 291 26899
rect 257 26797 291 26831
rect 257 26729 291 26763
rect 257 26661 291 26695
rect 257 26593 291 26627
rect 257 26525 291 26559
rect 257 26457 291 26491
rect 257 26389 291 26423
rect 257 26321 291 26355
rect 257 26253 291 26287
rect 257 26185 291 26219
rect 257 26117 291 26151
rect 257 26049 291 26083
rect 257 25981 291 26015
rect 257 25913 291 25947
rect 257 25845 291 25879
rect 257 25777 291 25811
rect 257 25709 291 25743
rect 257 25641 291 25675
rect 257 25573 291 25607
rect 257 25505 291 25539
rect 257 25437 291 25471
rect 257 25369 291 25403
rect 257 25301 291 25335
rect 257 25233 291 25267
rect 257 25165 291 25199
rect 257 25097 291 25131
rect 257 25029 291 25063
rect 257 24961 291 24995
rect 257 24893 291 24927
rect 257 24825 291 24859
rect 257 24757 291 24791
rect 257 24689 291 24723
rect 257 24621 291 24655
rect 257 24553 291 24587
rect 257 24485 291 24519
rect 257 24417 291 24451
rect 257 24349 291 24383
rect 257 24281 291 24315
rect 257 24213 291 24247
rect 257 24145 291 24179
rect 257 24077 291 24111
rect 257 24009 291 24043
rect 257 23941 291 23975
rect 257 23873 291 23907
rect 257 23805 291 23839
rect 2145 27469 2179 27503
rect 2145 27401 2179 27435
rect 2145 27333 2179 27367
rect 2145 27265 2179 27299
rect 2145 27197 2179 27231
rect 2145 27129 2179 27163
rect 2145 27061 2179 27095
rect 2145 26993 2179 27027
rect 2145 26925 2179 26959
rect 2145 26857 2179 26891
rect 2145 26789 2179 26823
rect 2145 26721 2179 26755
rect 2145 26653 2179 26687
rect 2145 26585 2179 26619
rect 2145 26517 2179 26551
rect 2145 26449 2179 26483
rect 2145 26381 2179 26415
rect 2145 26313 2179 26347
rect 2145 26245 2179 26279
rect 2145 26177 2179 26211
rect 2145 26109 2179 26143
rect 2145 26041 2179 26075
rect 2145 25973 2179 26007
rect 2145 25905 2179 25939
rect 2145 25837 2179 25871
rect 2145 25769 2179 25803
rect 2145 25701 2179 25735
rect 2145 25633 2179 25667
rect 2145 25565 2179 25599
rect 2145 25497 2179 25531
rect 2145 25429 2179 25463
rect 2145 25361 2179 25395
rect 2145 25293 2179 25327
rect 2145 25225 2179 25259
rect 2145 25157 2179 25191
rect 2145 25089 2179 25123
rect 2145 25021 2179 25055
rect 2145 24953 2179 24987
rect 2145 24885 2179 24919
rect 2145 24817 2179 24851
rect 2145 24749 2179 24783
rect 2145 24681 2179 24715
rect 2145 24613 2179 24647
rect 2145 24545 2179 24579
rect 2145 24477 2179 24511
rect 2145 24409 2179 24443
rect 2145 24341 2179 24375
rect 2145 24273 2179 24307
rect 2145 24205 2179 24239
rect 2145 24137 2179 24171
rect 2145 24069 2179 24103
rect 2145 24001 2179 24035
rect 2145 23933 2179 23967
rect 2145 23865 2179 23899
rect 257 23737 291 23771
rect 2145 23797 2179 23831
rect 257 23669 291 23703
rect 2145 23729 2179 23763
rect 257 23601 291 23635
rect 2145 23661 2179 23695
rect 257 23533 291 23567
rect 257 23465 291 23499
rect 257 23397 291 23431
rect 257 23329 291 23363
rect 257 23261 291 23295
rect 257 23193 291 23227
rect 257 23125 291 23159
rect 257 23057 291 23091
rect 257 22989 291 23023
rect 257 22921 291 22955
rect 257 22853 291 22887
rect 257 22785 291 22819
rect 257 22717 291 22751
rect 257 22649 291 22683
rect 257 22581 291 22615
rect 257 22513 291 22547
rect 257 22445 291 22479
rect 257 22377 291 22411
rect 257 22309 291 22343
rect 2145 23593 2179 23627
rect 2145 23525 2179 23559
rect 2145 23457 2179 23491
rect 2145 23389 2179 23423
rect 2145 23321 2179 23355
rect 2145 23253 2179 23287
rect 2145 23185 2179 23219
rect 2145 23117 2179 23151
rect 2145 23049 2179 23083
rect 2145 22981 2179 23015
rect 2145 22913 2179 22947
rect 2145 22845 2179 22879
rect 2145 22777 2179 22811
rect 2145 22709 2179 22743
rect 2145 22641 2179 22675
rect 2145 22573 2179 22607
rect 2145 22505 2179 22539
rect 2145 22437 2179 22471
rect 2145 22369 2179 22403
rect 257 22241 291 22275
rect 257 22173 291 22207
rect 257 22105 291 22139
rect 257 22037 291 22071
rect 257 21969 291 22003
rect 257 21901 291 21935
rect 257 21833 291 21867
rect 257 21765 291 21799
rect 257 21697 291 21731
rect 257 21629 291 21663
rect 257 21561 291 21595
rect 257 21493 291 21527
rect 257 21425 291 21459
rect 257 21357 291 21391
rect 257 21289 291 21323
rect 257 21221 291 21255
rect 257 21153 291 21187
rect 257 21085 291 21119
rect 257 21017 291 21051
rect 257 20949 291 20983
rect 257 20881 291 20915
rect 257 20813 291 20847
rect 257 20745 291 20779
rect 257 20677 291 20711
rect 257 20609 291 20643
rect 257 20541 291 20575
rect 257 20473 291 20507
rect 257 20405 291 20439
rect 257 20337 291 20371
rect 257 20269 291 20303
rect 257 20201 291 20235
rect 257 20133 291 20167
rect 257 20065 291 20099
rect 257 19997 291 20031
rect 257 19929 291 19963
rect 257 19861 291 19895
rect 2145 22301 2179 22335
rect 2145 22233 2179 22267
rect 2145 22165 2179 22199
rect 2145 22097 2179 22131
rect 2145 22029 2179 22063
rect 2145 21961 2179 21995
rect 2145 21893 2179 21927
rect 2145 21825 2179 21859
rect 2145 21757 2179 21791
rect 2145 21689 2179 21723
rect 2145 21621 2179 21655
rect 2145 21553 2179 21587
rect 2145 21485 2179 21519
rect 2145 21417 2179 21451
rect 2145 21349 2179 21383
rect 2145 21281 2179 21315
rect 2145 21213 2179 21247
rect 2145 21145 2179 21179
rect 2145 21077 2179 21111
rect 2145 21009 2179 21043
rect 2145 20941 2179 20975
rect 2145 20873 2179 20907
rect 2145 20805 2179 20839
rect 2145 20737 2179 20771
rect 2145 20669 2179 20703
rect 2145 20601 2179 20635
rect 2145 20533 2179 20567
rect 2145 20465 2179 20499
rect 2145 20397 2179 20431
rect 2145 20329 2179 20363
rect 2145 20261 2179 20295
rect 2145 20193 2179 20227
rect 2145 20125 2179 20159
rect 2145 20057 2179 20091
rect 2145 19989 2179 20023
rect 2145 19921 2179 19955
rect 2145 19853 2179 19887
rect 257 19793 291 19827
rect 2145 19785 2179 19819
rect 257 19725 291 19759
rect 2145 19717 2179 19751
rect 257 19657 291 19691
rect 257 19589 291 19623
rect 257 19521 291 19555
rect 257 19453 291 19487
rect 257 19385 291 19419
rect 257 19317 291 19351
rect 257 19249 291 19283
rect 257 19181 291 19215
rect 257 19113 291 19147
rect 257 19045 291 19079
rect 257 18977 291 19011
rect 257 18909 291 18943
rect 257 18841 291 18875
rect 257 18773 291 18807
rect 257 18705 291 18739
rect 257 18637 291 18671
rect 257 18569 291 18603
rect 257 18501 291 18535
rect 257 18433 291 18467
rect 257 18365 291 18399
rect 257 18297 291 18331
rect 257 18229 291 18263
rect 257 18161 291 18195
rect 257 18093 291 18127
rect 257 18025 291 18059
rect 257 17957 291 17991
rect 257 17889 291 17923
rect 257 17821 291 17855
rect 257 17753 291 17787
rect 257 17685 291 17719
rect 257 17617 291 17651
rect 257 17549 291 17583
rect 257 17481 291 17515
rect 257 17413 291 17447
rect 257 17345 291 17379
rect 257 17277 291 17311
rect 257 17209 291 17243
rect 257 17141 291 17175
rect 257 17073 291 17107
rect 257 17005 291 17039
rect 257 16937 291 16971
rect 257 16869 291 16903
rect 257 16801 291 16835
rect 257 16733 291 16767
rect 257 16665 291 16699
rect 257 16597 291 16631
rect 257 16529 291 16563
rect 257 16461 291 16495
rect 257 16393 291 16427
rect 257 16325 291 16359
rect 257 16257 291 16291
rect 257 16189 291 16223
rect 257 16121 291 16155
rect 257 16053 291 16087
rect 257 15985 291 16019
rect 2145 19649 2179 19683
rect 2145 19581 2179 19615
rect 2145 19513 2179 19547
rect 2145 19445 2179 19479
rect 2145 19377 2179 19411
rect 2145 19309 2179 19343
rect 2145 19241 2179 19275
rect 2145 19173 2179 19207
rect 2145 19105 2179 19139
rect 2145 19037 2179 19071
rect 2145 18969 2179 19003
rect 2145 18901 2179 18935
rect 2145 18833 2179 18867
rect 2145 18765 2179 18799
rect 2145 18697 2179 18731
rect 2145 18629 2179 18663
rect 2145 18561 2179 18595
rect 2145 18493 2179 18527
rect 2145 18425 2179 18459
rect 2145 18357 2179 18391
rect 2145 18289 2179 18323
rect 2145 18221 2179 18255
rect 2145 18153 2179 18187
rect 2145 18085 2179 18119
rect 2145 18017 2179 18051
rect 2145 17949 2179 17983
rect 2145 17881 2179 17915
rect 2145 17813 2179 17847
rect 2145 17745 2179 17779
rect 2145 17677 2179 17711
rect 2145 17609 2179 17643
rect 2145 17541 2179 17575
rect 2145 17473 2179 17507
rect 2145 17405 2179 17439
rect 2145 17337 2179 17371
rect 2145 17269 2179 17303
rect 2145 17201 2179 17235
rect 2145 17133 2179 17167
rect 2145 17065 2179 17099
rect 2145 16997 2179 17031
rect 2145 16929 2179 16963
rect 2145 16861 2179 16895
rect 2145 16793 2179 16827
rect 2145 16725 2179 16759
rect 2145 16657 2179 16691
rect 2145 16589 2179 16623
rect 2145 16521 2179 16555
rect 2145 16453 2179 16487
rect 2145 16385 2179 16419
rect 2145 16317 2179 16351
rect 2145 16249 2179 16283
rect 2145 16181 2179 16215
rect 2145 16113 2179 16147
rect 2145 16045 2179 16079
rect 257 15917 291 15951
rect 2145 15977 2179 16011
rect 2145 15909 2179 15943
rect 257 15849 291 15883
rect 2145 15841 2179 15875
rect 257 15781 291 15815
rect 257 15713 291 15747
rect 257 15645 291 15679
rect 257 15577 291 15611
rect 257 15509 291 15543
rect 257 15441 291 15475
rect 257 15373 291 15407
rect 257 15305 291 15339
rect 257 15237 291 15271
rect 257 15169 291 15203
rect 257 15101 291 15135
rect 257 15033 291 15067
rect 257 14965 291 14999
rect 257 14897 291 14931
rect 257 14829 291 14863
rect 257 14761 291 14795
rect 257 14693 291 14727
rect 257 14625 291 14659
rect 257 14557 291 14591
rect 257 14489 291 14523
rect 257 14421 291 14455
rect 257 14353 291 14387
rect 257 14285 291 14319
rect 257 14217 291 14251
rect 257 14149 291 14183
rect 257 14081 291 14115
rect 257 14013 291 14047
rect 257 13945 291 13979
rect 257 13877 291 13911
rect 257 13809 291 13843
rect 257 13741 291 13775
rect 257 13673 291 13707
rect 257 13605 291 13639
rect 257 13537 291 13571
rect 257 13469 291 13503
rect 257 13401 291 13435
rect 257 13333 291 13367
rect 257 13265 291 13299
rect 257 13197 291 13231
rect 257 13129 291 13163
rect 257 13061 291 13095
rect 257 12993 291 13027
rect 257 12925 291 12959
rect 257 12857 291 12891
rect 257 12789 291 12823
rect 257 12721 291 12755
rect 257 12653 291 12687
rect 257 12585 291 12619
rect 257 12517 291 12551
rect 257 12449 291 12483
rect 257 12381 291 12415
rect 257 12313 291 12347
rect 257 12245 291 12279
rect 257 12177 291 12211
rect 257 12109 291 12143
rect 2145 15773 2179 15807
rect 2145 15705 2179 15739
rect 2145 15637 2179 15671
rect 2145 15569 2179 15603
rect 2145 15501 2179 15535
rect 2145 15433 2179 15467
rect 2145 15365 2179 15399
rect 2145 15297 2179 15331
rect 2145 15229 2179 15263
rect 2145 15161 2179 15195
rect 2145 15093 2179 15127
rect 2145 15025 2179 15059
rect 2145 14957 2179 14991
rect 2145 14889 2179 14923
rect 2145 14821 2179 14855
rect 2145 14753 2179 14787
rect 2145 14685 2179 14719
rect 2145 14617 2179 14651
rect 2145 14549 2179 14583
rect 2145 14481 2179 14515
rect 2145 14413 2179 14447
rect 2145 14345 2179 14379
rect 2145 14277 2179 14311
rect 2145 14209 2179 14243
rect 2145 14141 2179 14175
rect 2145 14073 2179 14107
rect 2145 14005 2179 14039
rect 2145 13937 2179 13971
rect 2145 13869 2179 13903
rect 2145 13801 2179 13835
rect 2145 13733 2179 13767
rect 2145 13665 2179 13699
rect 2145 13597 2179 13631
rect 2145 13529 2179 13563
rect 2145 13461 2179 13495
rect 2145 13393 2179 13427
rect 2145 13325 2179 13359
rect 2145 13257 2179 13291
rect 2145 13189 2179 13223
rect 2145 13121 2179 13155
rect 2145 13053 2179 13087
rect 2145 12985 2179 13019
rect 2145 12917 2179 12951
rect 2145 12849 2179 12883
rect 2145 12781 2179 12815
rect 2145 12713 2179 12747
rect 2145 12645 2179 12679
rect 2145 12577 2179 12611
rect 2145 12509 2179 12543
rect 2145 12441 2179 12475
rect 2145 12373 2179 12407
rect 2145 12305 2179 12339
rect 2145 12237 2179 12271
rect 2145 12169 2179 12203
rect 257 12041 291 12075
rect 2145 12101 2179 12135
rect 257 11973 291 12007
rect 2145 12033 2179 12067
rect 257 11905 291 11939
rect 2145 11965 2179 11999
rect 257 11837 291 11871
rect 257 11769 291 11803
rect 257 11701 291 11735
rect 257 11633 291 11667
rect 257 11565 291 11599
rect 257 11497 291 11531
rect 257 11429 291 11463
rect 257 11361 291 11395
rect 257 11293 291 11327
rect 257 11225 291 11259
rect 257 11157 291 11191
rect 257 11089 291 11123
rect 257 11021 291 11055
rect 257 10953 291 10987
rect 257 10885 291 10919
rect 257 10817 291 10851
rect 257 10749 291 10783
rect 257 10681 291 10715
rect 257 10613 291 10647
rect 257 10545 291 10579
rect 257 10477 291 10511
rect 257 10409 291 10443
rect 257 10341 291 10375
rect 257 10273 291 10307
rect 257 10205 291 10239
rect 257 10137 291 10171
rect 257 10069 291 10103
rect 257 10001 291 10035
rect 257 9933 291 9967
rect 257 9865 291 9899
rect 257 9797 291 9831
rect 257 9729 291 9763
rect 257 9661 291 9695
rect 257 9593 291 9627
rect 257 9525 291 9559
rect 257 9457 291 9491
rect 257 9389 291 9423
rect 257 9321 291 9355
rect 257 9253 291 9287
rect 257 9185 291 9219
rect 257 9117 291 9151
rect 257 9049 291 9083
rect 257 8981 291 9015
rect 257 8913 291 8947
rect 257 8845 291 8879
rect 257 8777 291 8811
rect 257 8709 291 8743
rect 257 8641 291 8675
rect 257 8573 291 8607
rect 257 8505 291 8539
rect 257 8437 291 8471
rect 257 8369 291 8403
rect 257 8301 291 8335
rect 257 8233 291 8267
rect 2145 11897 2179 11931
rect 2145 11829 2179 11863
rect 2145 11761 2179 11795
rect 2145 11693 2179 11727
rect 2145 11625 2179 11659
rect 2145 11557 2179 11591
rect 2145 11489 2179 11523
rect 2145 11421 2179 11455
rect 2145 11353 2179 11387
rect 2145 11285 2179 11319
rect 2145 11217 2179 11251
rect 2145 11149 2179 11183
rect 2145 11081 2179 11115
rect 2145 11013 2179 11047
rect 2145 10945 2179 10979
rect 2145 10877 2179 10911
rect 2145 10809 2179 10843
rect 2145 10741 2179 10775
rect 2145 10673 2179 10707
rect 2145 10605 2179 10639
rect 2145 10537 2179 10571
rect 2145 10469 2179 10503
rect 2145 10401 2179 10435
rect 2145 10333 2179 10367
rect 2145 10265 2179 10299
rect 2145 10197 2179 10231
rect 2145 10129 2179 10163
rect 2145 10061 2179 10095
rect 2145 9993 2179 10027
rect 2145 9925 2179 9959
rect 2145 9857 2179 9891
rect 2145 9789 2179 9823
rect 2145 9721 2179 9755
rect 2145 9653 2179 9687
rect 2145 9585 2179 9619
rect 2145 9517 2179 9551
rect 2145 9449 2179 9483
rect 2145 9381 2179 9415
rect 2145 9313 2179 9347
rect 2145 9245 2179 9279
rect 2145 9177 2179 9211
rect 2145 9109 2179 9143
rect 2145 9041 2179 9075
rect 2145 8973 2179 9007
rect 2145 8905 2179 8939
rect 2145 8837 2179 8871
rect 2145 8769 2179 8803
rect 2145 8701 2179 8735
rect 2145 8633 2179 8667
rect 2145 8565 2179 8599
rect 2145 8497 2179 8531
rect 2145 8429 2179 8463
rect 2145 8361 2179 8395
rect 2145 8293 2179 8327
rect 2145 8225 2179 8259
rect 257 8165 291 8199
rect 257 8097 291 8131
rect 257 8029 291 8063
rect 257 7961 291 7995
rect 257 7893 291 7927
rect 257 7825 291 7859
rect 257 7757 291 7791
rect 257 7689 291 7723
rect 257 7621 291 7655
rect 257 7553 291 7587
rect 257 7485 291 7519
rect 257 7417 291 7451
rect 257 7349 291 7383
rect 257 7281 291 7315
rect 257 7213 291 7247
rect 257 7145 291 7179
rect 257 7077 291 7111
rect 257 7009 291 7043
rect 257 6941 291 6975
rect 257 6873 291 6907
rect 231 6732 265 6766
rect 231 6660 265 6694
rect 231 6589 265 6623
rect 231 6518 265 6552
rect 231 6447 265 6481
rect 231 6376 265 6410
rect 231 6305 265 6339
rect 231 6234 265 6268
rect 231 6163 265 6197
rect 231 6092 265 6126
rect 231 6021 265 6055
rect 231 5950 265 5984
rect 231 5879 265 5913
rect 231 5808 265 5842
rect 253 5672 287 5706
rect 253 5604 287 5638
rect 253 5536 287 5570
rect 2145 8157 2179 8191
rect 2145 8089 2179 8123
rect 2145 8021 2179 8055
rect 2145 7953 2179 7987
rect 2145 7885 2179 7919
rect 2145 7817 2179 7851
rect 2145 7749 2179 7783
rect 2145 7681 2179 7715
rect 2145 7613 2179 7647
rect 2145 7545 2179 7579
rect 2145 7477 2179 7511
rect 2145 7409 2179 7443
rect 2145 7341 2179 7375
rect 2145 7273 2179 7307
rect 2145 7205 2179 7239
rect 2145 7137 2179 7171
rect 2145 7069 2179 7103
rect 2145 7001 2179 7035
rect 2145 6933 2179 6967
rect 2145 6865 2179 6899
rect 2145 6797 2179 6831
rect 2145 6729 2179 6763
rect 2145 6661 2179 6695
rect 2145 6593 2179 6627
rect 2145 6525 2179 6559
rect 2145 6457 2179 6491
rect 2145 6389 2179 6423
rect 2145 6321 2179 6355
rect 2145 6253 2179 6287
rect 2145 6185 2179 6219
rect 2145 6117 2179 6151
rect 2145 6049 2179 6083
rect 2743 10822 2777 10856
rect 2835 10855 2869 10889
rect 2903 10855 2937 10889
rect 2971 10855 3005 10889
rect 3039 10855 3073 10889
rect 3107 10855 3141 10889
rect 3175 10855 3209 10889
rect 3243 10855 3277 10889
rect 3311 10855 3345 10889
rect 3379 10855 3413 10889
rect 3447 10855 3481 10889
rect 3515 10855 3549 10889
rect 3583 10855 3617 10889
rect 3651 10855 3685 10889
rect 3719 10855 3753 10889
rect 3787 10855 3821 10889
rect 3855 10855 3889 10889
rect 3923 10855 3957 10889
rect 3991 10855 4025 10889
rect 4059 10855 4093 10889
rect 4127 10855 4161 10889
rect 4195 10855 4229 10889
rect 4263 10855 4297 10889
rect 4331 10855 4365 10889
rect 4399 10855 4433 10889
rect 4467 10855 4501 10889
rect 4535 10855 4569 10889
rect 4603 10855 4637 10889
rect 4671 10855 4705 10889
rect 4799 10855 4833 10889
rect 4867 10855 4901 10889
rect 4935 10855 4969 10889
rect 5003 10855 5037 10889
rect 5071 10855 5105 10889
rect 5139 10855 5173 10889
rect 5207 10855 5241 10889
rect 5275 10855 5309 10889
rect 5343 10855 5377 10889
rect 5411 10855 5445 10889
rect 5479 10855 5513 10889
rect 5547 10855 5581 10889
rect 5615 10855 5649 10889
rect 5683 10855 5717 10889
rect 5751 10855 5785 10889
rect 5819 10855 5853 10889
rect 5887 10855 5921 10889
rect 5955 10855 5989 10889
rect 6023 10855 6057 10889
rect 6091 10855 6125 10889
rect 6159 10855 6193 10889
rect 6227 10855 6261 10889
rect 6295 10855 6329 10889
rect 6363 10855 6397 10889
rect 6431 10855 6465 10889
rect 6499 10855 6533 10889
rect 6567 10855 6601 10889
rect 2743 10754 2777 10788
rect 6665 10822 6699 10856
rect 2743 10686 2777 10720
rect 2743 10618 2777 10652
rect 2743 10550 2777 10584
rect 2743 10482 2777 10516
rect 2743 10414 2777 10448
rect 2743 10346 2777 10380
rect 2743 10278 2777 10312
rect 2743 10210 2777 10244
rect 2743 10142 2777 10176
rect 2743 10074 2777 10108
rect 2743 10006 2777 10040
rect 2743 9938 2777 9972
rect 2743 9870 2777 9904
rect 2743 9802 2777 9836
rect 2743 9734 2777 9768
rect 2743 9666 2777 9700
rect 2743 9598 2777 9632
rect 2743 9530 2777 9564
rect 2743 9462 2777 9496
rect 2743 9394 2777 9428
rect 2743 9326 2777 9360
rect 2743 9258 2777 9292
rect 2743 9190 2777 9224
rect 2743 9122 2777 9156
rect 2743 9054 2777 9088
rect 2743 8986 2777 9020
rect 2743 8918 2777 8952
rect 2743 8850 2777 8884
rect 2743 8782 2777 8816
rect 2743 8714 2777 8748
rect 2743 8646 2777 8680
rect 2743 8578 2777 8612
rect 2743 8510 2777 8544
rect 2743 8442 2777 8476
rect 2743 8374 2777 8408
rect 2743 8306 2777 8340
rect 2743 8238 2777 8272
rect 2743 8170 2777 8204
rect 2743 8102 2777 8136
rect 2743 8034 2777 8068
rect 2743 7966 2777 8000
rect 2743 7898 2777 7932
rect 2743 7830 2777 7864
rect 2743 7762 2777 7796
rect 2743 7694 2777 7728
rect 2743 7626 2777 7660
rect 2743 7558 2777 7592
rect 2743 7490 2777 7524
rect 2743 7422 2777 7456
rect 2743 7354 2777 7388
rect 2743 7286 2777 7320
rect 2743 7218 2777 7252
rect 2743 7150 2777 7184
rect 2743 7082 2777 7116
rect 2743 7014 2777 7048
rect 2743 6946 2777 6980
rect 2743 6878 2777 6912
rect 2743 6810 2777 6844
rect 2743 6742 2777 6776
rect 2743 6674 2777 6708
rect 2743 6606 2777 6640
rect 2743 6538 2777 6572
rect 4704 10742 4738 10776
rect 6665 10754 6699 10788
rect 4704 10674 4738 10708
rect 4704 10606 4738 10640
rect 4704 10538 4738 10572
rect 4704 10470 4738 10504
rect 4704 10402 4738 10436
rect 4704 10334 4738 10368
rect 4704 10266 4738 10300
rect 4704 10198 4738 10232
rect 4704 10130 4738 10164
rect 4704 10062 4738 10096
rect 4704 9994 4738 10028
rect 4704 9926 4738 9960
rect 4704 9858 4738 9892
rect 4704 9790 4738 9824
rect 4704 9722 4738 9756
rect 4704 9654 4738 9688
rect 4704 9586 4738 9620
rect 4704 9518 4738 9552
rect 4704 9450 4738 9484
rect 4704 9382 4738 9416
rect 4704 9314 4738 9348
rect 4704 9246 4738 9280
rect 4704 9178 4738 9212
rect 4704 9110 4738 9144
rect 4704 9042 4738 9076
rect 4704 8974 4738 9008
rect 4704 8906 4738 8940
rect 4704 8838 4738 8872
rect 4704 8770 4738 8804
rect 4704 8702 4738 8736
rect 4704 8634 4738 8668
rect 4704 8566 4738 8600
rect 4704 8498 4738 8532
rect 4704 8430 4738 8464
rect 4704 8362 4738 8396
rect 4704 8294 4738 8328
rect 4704 8226 4738 8260
rect 4704 8158 4738 8192
rect 4704 8090 4738 8124
rect 4704 8022 4738 8056
rect 4704 7954 4738 7988
rect 4704 7886 4738 7920
rect 4704 7818 4738 7852
rect 4704 7750 4738 7784
rect 4704 7682 4738 7716
rect 4704 7614 4738 7648
rect 4704 7546 4738 7580
rect 4704 7478 4738 7512
rect 4704 7410 4738 7444
rect 4704 7342 4738 7376
rect 4704 7274 4738 7308
rect 4704 7206 4738 7240
rect 4704 7138 4738 7172
rect 4704 7070 4738 7104
rect 4704 7002 4738 7036
rect 4704 6934 4738 6968
rect 4704 6866 4738 6900
rect 4704 6798 4738 6832
rect 4704 6730 4738 6764
rect 4704 6662 4738 6696
rect 4704 6594 4738 6628
rect 6665 10686 6699 10720
rect 6665 10618 6699 10652
rect 6665 10550 6699 10584
rect 6665 10482 6699 10516
rect 6665 10414 6699 10448
rect 6665 10346 6699 10380
rect 6665 10278 6699 10312
rect 6665 10210 6699 10244
rect 6665 10142 6699 10176
rect 6665 10074 6699 10108
rect 6665 10006 6699 10040
rect 6665 9938 6699 9972
rect 6665 9870 6699 9904
rect 6665 9802 6699 9836
rect 6665 9734 6699 9768
rect 6665 9666 6699 9700
rect 6665 9598 6699 9632
rect 6665 9530 6699 9564
rect 6665 9462 6699 9496
rect 6665 9394 6699 9428
rect 6665 9326 6699 9360
rect 6665 9258 6699 9292
rect 6665 9190 6699 9224
rect 6665 9122 6699 9156
rect 6665 9054 6699 9088
rect 6665 8986 6699 9020
rect 6665 8918 6699 8952
rect 6665 8850 6699 8884
rect 6665 8782 6699 8816
rect 6665 8714 6699 8748
rect 6665 8646 6699 8680
rect 6665 8578 6699 8612
rect 6665 8510 6699 8544
rect 6665 8442 6699 8476
rect 6665 8374 6699 8408
rect 6665 8306 6699 8340
rect 6665 8238 6699 8272
rect 6665 8170 6699 8204
rect 6665 8102 6699 8136
rect 6665 8034 6699 8068
rect 6665 7966 6699 8000
rect 6665 7898 6699 7932
rect 6665 7830 6699 7864
rect 6665 7762 6699 7796
rect 6665 7694 6699 7728
rect 6665 7626 6699 7660
rect 6665 7558 6699 7592
rect 6665 7490 6699 7524
rect 6665 7422 6699 7456
rect 6665 7354 6699 7388
rect 6665 7286 6699 7320
rect 6665 7218 6699 7252
rect 6665 7150 6699 7184
rect 6665 7082 6699 7116
rect 6665 7014 6699 7048
rect 6665 6946 6699 6980
rect 6665 6878 6699 6912
rect 6665 6810 6699 6844
rect 6665 6742 6699 6776
rect 6665 6674 6699 6708
rect 6665 6606 6699 6640
rect 4704 6526 4738 6560
rect 2776 6425 2810 6459
rect 2844 6425 2878 6459
rect 2912 6425 2946 6459
rect 2980 6425 3014 6459
rect 3048 6425 3082 6459
rect 3116 6425 3150 6459
rect 3184 6425 3218 6459
rect 3252 6425 3286 6459
rect 3320 6425 3354 6459
rect 3388 6425 3422 6459
rect 3456 6425 3490 6459
rect 3524 6425 3558 6459
rect 3592 6425 3626 6459
rect 3660 6425 3694 6459
rect 3728 6425 3762 6459
rect 3796 6425 3830 6459
rect 3864 6425 3898 6459
rect 3932 6425 3966 6459
rect 4000 6425 4034 6459
rect 4068 6425 4102 6459
rect 4136 6425 4170 6459
rect 4204 6425 4238 6459
rect 4272 6425 4306 6459
rect 4340 6425 4374 6459
rect 4408 6425 4442 6459
rect 4476 6425 4510 6459
rect 4544 6425 4578 6459
rect 4612 6425 4646 6459
rect 4704 6458 4738 6492
rect 6665 6538 6699 6572
rect 4796 6425 4830 6459
rect 4864 6425 4898 6459
rect 4932 6425 4966 6459
rect 5000 6425 5034 6459
rect 5068 6425 5102 6459
rect 5136 6425 5170 6459
rect 5204 6425 5238 6459
rect 5272 6425 5306 6459
rect 5340 6425 5374 6459
rect 5408 6425 5442 6459
rect 5476 6425 5510 6459
rect 5544 6425 5578 6459
rect 5612 6425 5646 6459
rect 5680 6425 5714 6459
rect 5748 6425 5782 6459
rect 5816 6425 5850 6459
rect 5884 6425 5918 6459
rect 5952 6425 5986 6459
rect 6020 6425 6054 6459
rect 6088 6425 6122 6459
rect 6156 6425 6190 6459
rect 6224 6425 6258 6459
rect 6292 6425 6326 6459
rect 6360 6425 6394 6459
rect 6428 6425 6462 6459
rect 6496 6425 6530 6459
rect 6564 6425 6598 6459
rect 6632 6425 6666 6459
rect 2145 5981 2179 6015
rect 2145 5913 2179 5947
rect 2145 5845 2179 5879
rect 2145 5777 2179 5811
rect 2145 5709 2179 5743
rect 2145 5641 2179 5675
rect 2145 5573 2179 5607
rect 2280 5540 2314 5574
rect 2576 5540 2610 5574
rect 2644 5540 2678 5574
rect 2712 5540 2746 5574
rect 2780 5540 2814 5574
rect 2848 5540 2882 5574
rect 2916 5540 2950 5574
rect 2984 5540 3018 5574
rect 3052 5540 3086 5574
rect 3120 5540 3154 5574
rect 253 5468 287 5502
rect 231 5368 265 5402
rect 3153 5458 3187 5492
rect 231 5295 265 5329
rect 231 5222 265 5256
rect 231 5149 265 5183
rect 231 5076 265 5110
rect 231 5003 265 5037
rect 231 4931 265 4965
rect 231 4859 265 4893
rect 231 4787 265 4821
rect 231 4715 265 4749
rect 231 4643 265 4677
rect 231 4571 265 4605
rect 231 4499 265 4533
rect 231 4427 265 4461
rect 257 4319 291 4353
rect 3153 5390 3187 5424
rect 3153 5322 3187 5356
rect 3153 5254 3187 5288
rect 3153 5186 3187 5220
rect 3153 5118 3187 5152
rect 3153 5050 3187 5084
rect 3153 4982 3187 5016
rect 3153 4914 3187 4948
rect 3153 4846 3187 4880
rect 3153 4778 3187 4812
rect 3153 4710 3187 4744
rect 3153 4642 3187 4676
rect 3153 4574 3187 4608
rect 3153 4506 3187 4540
rect 3153 4438 3187 4472
rect 3153 4370 3187 4404
rect 257 4250 291 4284
rect 3153 4302 3187 4336
rect 3531 5508 3565 5542
rect 3651 5541 3685 5575
rect 3719 5541 3753 5575
rect 3787 5541 3821 5575
rect 3855 5541 3889 5575
rect 3923 5541 3957 5575
rect 3991 5541 4025 5575
rect 4059 5541 4093 5575
rect 4127 5541 4161 5575
rect 4195 5541 4229 5575
rect 4263 5541 4297 5575
rect 4331 5541 4365 5575
rect 4399 5541 4433 5575
rect 4467 5541 4501 5575
rect 4535 5541 4569 5575
rect 4603 5541 4637 5575
rect 4671 5541 4705 5575
rect 4739 5541 4773 5575
rect 4807 5541 4841 5575
rect 4875 5541 4909 5575
rect 4943 5541 4977 5575
rect 5011 5541 5045 5575
rect 5079 5541 5113 5575
rect 5147 5541 5181 5575
rect 5215 5541 5249 5575
rect 5283 5541 5317 5575
rect 5351 5541 5385 5575
rect 5588 5541 5622 5575
rect 3531 5440 3565 5474
rect 3531 5372 3565 5406
rect 3531 5304 3565 5338
rect 3531 5236 3565 5270
rect 3531 5168 3565 5202
rect 3531 5100 3565 5134
rect 3531 5032 3565 5066
rect 3531 4964 3565 4998
rect 3531 4896 3565 4930
rect 3531 4828 3565 4862
rect 3531 4760 3565 4794
rect 3531 4692 3565 4726
rect 3531 4624 3565 4658
rect 3531 4556 3565 4590
rect 3531 4488 3565 4522
rect 3531 4420 3565 4454
rect 5621 5422 5655 5456
rect 5621 5354 5655 5388
rect 5621 5286 5655 5320
rect 5621 5218 5655 5252
rect 5621 5150 5655 5184
rect 5621 5082 5655 5116
rect 5621 5014 5655 5048
rect 5621 4946 5655 4980
rect 5621 4878 5655 4912
rect 5621 4810 5655 4844
rect 5621 4742 5655 4776
rect 5621 4674 5655 4708
rect 5621 4606 5655 4640
rect 5621 4538 5655 4572
rect 5621 4470 5655 4504
rect 5621 4402 5655 4436
rect 3564 4301 3598 4335
rect 3632 4301 3666 4335
rect 3700 4301 3734 4335
rect 3768 4301 3802 4335
rect 3836 4301 3870 4335
rect 3904 4301 3938 4335
rect 3972 4301 4006 4335
rect 4040 4301 4074 4335
rect 4108 4301 4142 4335
rect 4176 4301 4210 4335
rect 4244 4301 4278 4335
rect 4312 4301 4346 4335
rect 4380 4301 4414 4335
rect 4448 4301 4482 4335
rect 4516 4301 4550 4335
rect 4584 4301 4618 4335
rect 4652 4301 4686 4335
rect 4720 4301 4754 4335
rect 4788 4301 4822 4335
rect 4856 4301 4890 4335
rect 4924 4301 4958 4335
rect 4992 4301 5026 4335
rect 5060 4301 5094 4335
rect 5128 4301 5162 4335
rect 5196 4301 5230 4335
rect 5264 4301 5298 4335
rect 5332 4301 5366 4335
rect 5400 4301 5434 4335
rect 5468 4301 5502 4335
rect 5536 4301 5570 4335
rect 5621 4334 5655 4368
rect 257 4181 291 4215
rect 3153 4234 3187 4268
rect 257 4112 291 4146
rect 3153 4166 3187 4200
rect 3153 4098 3187 4132
rect 257 4043 291 4077
rect 257 3974 291 4008
rect 257 3905 291 3939
rect 257 3836 291 3870
rect 257 3767 291 3801
rect 257 3698 291 3732
rect 257 3629 291 3663
rect 257 3560 291 3594
rect 257 3491 291 3525
rect 257 3422 291 3456
rect 257 3353 291 3387
rect 257 3284 291 3318
rect 257 3215 291 3249
rect 257 3146 291 3180
rect 257 3077 291 3111
rect 257 3008 291 3042
rect 257 2939 291 2973
rect 257 2870 291 2904
rect 257 2801 291 2835
rect 257 2732 291 2766
rect 257 2663 291 2697
rect 257 2594 291 2628
rect 257 2525 291 2559
rect 257 2456 291 2490
rect 257 2387 291 2421
rect 257 2318 291 2352
rect 257 2249 291 2283
rect 257 2180 291 2214
rect 257 2111 291 2145
rect 257 2042 291 2076
rect 257 1973 291 2007
rect 257 1904 291 1938
rect 257 1835 291 1869
rect 257 1766 291 1800
rect 257 1697 291 1731
rect 257 1628 291 1662
rect 257 1559 291 1593
rect 257 1490 291 1524
rect 257 1422 291 1456
rect 257 1354 291 1388
rect 257 1286 291 1320
rect 257 1218 291 1252
rect 257 1150 291 1184
rect 257 1082 291 1116
rect 257 1014 291 1048
rect 257 946 291 980
rect 257 878 291 912
rect 257 810 291 844
rect 257 742 291 776
rect 257 674 291 708
rect 257 606 291 640
rect 257 538 291 572
rect 257 470 291 504
rect 257 402 291 436
rect 3153 4030 3187 4064
rect 3153 3962 3187 3996
rect 3153 3894 3187 3928
rect 3153 3826 3187 3860
rect 3153 3758 3187 3792
rect 3153 3690 3187 3724
rect 3153 3622 3187 3656
rect 3153 3554 3187 3588
rect 3153 3486 3187 3520
rect 3153 3418 3187 3452
rect 3153 3350 3187 3384
rect 3153 3282 3187 3316
rect 3153 3214 3187 3248
rect 3153 3146 3187 3180
rect 3153 3078 3187 3112
rect 3153 3010 3187 3044
rect 3153 2942 3187 2976
rect 3153 2874 3187 2908
rect 3153 2806 3187 2840
rect 3153 2738 3187 2772
rect 3153 2670 3187 2704
rect 3153 2602 3187 2636
rect 3153 2534 3187 2568
rect 3153 2466 3187 2500
rect 3153 2398 3187 2432
rect 3153 2330 3187 2364
rect 3153 2262 3187 2296
rect 3153 2194 3187 2228
rect 3153 2126 3187 2160
rect 3153 2058 3187 2092
rect 3153 1990 3187 2024
rect 3153 1922 3187 1956
rect 3153 1854 3187 1888
rect 3153 1786 3187 1820
rect 3153 1718 3187 1752
rect 3153 1650 3187 1684
rect 3153 1582 3187 1616
rect 3153 1514 3187 1548
rect 3153 1446 3187 1480
rect 3153 1378 3187 1412
rect 3153 1310 3187 1344
rect 3153 1242 3187 1276
rect 3153 1174 3187 1208
rect 3153 1106 3187 1140
rect 3153 1038 3187 1072
rect 3153 970 3187 1004
rect 3153 902 3187 936
rect 3153 834 3187 868
rect 3153 766 3187 800
rect 3153 698 3187 732
rect 3153 630 3187 664
rect 3153 562 3187 596
rect 3153 494 3187 528
rect 3153 426 3187 460
rect 3153 358 3187 392
rect 290 257 324 291
rect 358 257 392 291
rect 426 257 460 291
rect 494 257 528 291
rect 562 257 596 291
rect 630 257 664 291
rect 698 257 732 291
rect 766 257 800 291
rect 834 257 868 291
rect 902 257 936 291
rect 970 257 1004 291
rect 1038 257 1072 291
rect 1106 257 1140 291
rect 1174 257 1208 291
rect 1242 257 1276 291
rect 1310 257 1344 291
rect 1378 257 1412 291
rect 1446 257 1480 291
rect 1514 257 1548 291
rect 1582 257 1616 291
rect 1650 257 1684 291
rect 1718 257 1752 291
rect 1786 257 1820 291
rect 1854 257 1888 291
rect 1922 257 1956 291
rect 1990 257 2024 291
rect 2058 257 2092 291
rect 2126 257 2160 291
rect 2194 257 2228 291
rect 2262 257 2296 291
rect 2330 257 2364 291
rect 2398 257 2432 291
rect 2466 257 2500 291
rect 2534 257 2568 291
rect 2602 257 2636 291
rect 2670 257 2704 291
rect 2738 257 2772 291
rect 2806 257 2840 291
rect 2874 257 2908 291
rect 2942 257 2976 291
rect 3010 257 3044 291
rect 3078 257 3112 291
rect 3153 290 3187 324
<< mvnsubdiffcont >>
rect 68 27802 102 27836
rect 165 27835 199 27869
rect 233 27835 267 27869
rect 301 27835 335 27869
rect 369 27835 403 27869
rect 437 27835 471 27869
rect 505 27835 539 27869
rect 573 27835 607 27869
rect 641 27835 675 27869
rect 709 27835 743 27869
rect 777 27835 811 27869
rect 845 27835 879 27869
rect 913 27835 947 27869
rect 981 27835 1015 27869
rect 1049 27835 1083 27869
rect 1117 27835 1151 27869
rect 1185 27835 1219 27869
rect 1253 27835 1287 27869
rect 1321 27835 1355 27869
rect 1389 27835 1423 27869
rect 1457 27835 1491 27869
rect 1525 27835 1559 27869
rect 1593 27835 1627 27869
rect 1661 27835 1695 27869
rect 1729 27835 1763 27869
rect 1797 27835 1831 27869
rect 1865 27835 1899 27869
rect 1998 27835 2032 27869
rect 2066 27835 2100 27869
rect 2134 27835 2168 27869
rect 2202 27835 2236 27869
rect 68 27734 102 27768
rect 68 27666 102 27700
rect 2334 27763 2368 27797
rect 2334 27695 2368 27729
rect 68 27598 102 27632
rect 68 27530 102 27564
rect 68 27462 102 27496
rect 68 27394 102 27428
rect 68 27326 102 27360
rect 68 27258 102 27292
rect 68 27190 102 27224
rect 68 27122 102 27156
rect 68 27054 102 27088
rect 68 26986 102 27020
rect 68 26918 102 26952
rect 68 26850 102 26884
rect 68 26782 102 26816
rect 68 26714 102 26748
rect 68 26646 102 26680
rect 68 26578 102 26612
rect 68 26510 102 26544
rect 68 26442 102 26476
rect 68 26374 102 26408
rect 68 26306 102 26340
rect 68 26238 102 26272
rect 68 26170 102 26204
rect 68 26102 102 26136
rect 68 26034 102 26068
rect 68 25966 102 26000
rect 68 25898 102 25932
rect 68 25830 102 25864
rect 68 25762 102 25796
rect 2334 27627 2368 27661
rect 2334 27559 2368 27593
rect 2334 27491 2368 27525
rect 2334 27423 2368 27457
rect 2334 27355 2368 27389
rect 2334 27287 2368 27321
rect 2334 27219 2368 27253
rect 2334 27151 2368 27185
rect 2334 27083 2368 27117
rect 2334 27015 2368 27049
rect 2334 26947 2368 26981
rect 2334 26879 2368 26913
rect 2334 26811 2368 26845
rect 2334 26743 2368 26777
rect 2334 26675 2368 26709
rect 2334 26607 2368 26641
rect 2334 26539 2368 26573
rect 2334 26471 2368 26505
rect 2334 26403 2368 26437
rect 2334 26335 2368 26369
rect 2334 26267 2368 26301
rect 2334 26199 2368 26233
rect 2334 26131 2368 26165
rect 2334 26063 2368 26097
rect 2334 25995 2368 26029
rect 2334 25927 2368 25961
rect 2334 25859 2368 25893
rect 2334 25791 2368 25825
rect 2334 25723 2368 25757
rect 2334 25655 2368 25689
rect 2334 25587 2368 25621
rect 2334 25519 2368 25553
rect 2334 25451 2368 25485
rect 2334 25383 2368 25417
rect 2334 25315 2368 25349
rect 2334 25247 2368 25281
rect 2334 25179 2368 25213
rect 2334 25111 2368 25145
rect 2334 25043 2368 25077
rect 2334 24975 2368 25009
rect 2334 24907 2368 24941
rect 2334 24839 2368 24873
rect 2334 24771 2368 24805
rect 2334 24703 2368 24737
rect 2334 24635 2368 24669
rect 2334 24567 2368 24601
rect 2334 24499 2368 24533
rect 2334 24431 2368 24465
rect 2334 24363 2368 24397
rect 2334 24295 2368 24329
rect 2334 24227 2368 24261
rect 2334 24159 2368 24193
rect 2334 24091 2368 24125
rect 2334 24023 2368 24057
rect 2334 23955 2368 23989
rect 2334 23887 2368 23921
rect 2334 23819 2368 23853
rect 2334 23751 2368 23785
rect 2334 23683 2368 23717
rect 2334 23615 2368 23649
rect 2334 23547 2368 23581
rect 2334 23479 2368 23513
rect 2334 23411 2368 23445
rect 2334 23343 2368 23377
rect 2334 23275 2368 23309
rect 2334 23207 2368 23241
rect 2334 23139 2368 23173
rect 2334 23071 2368 23105
rect 2334 23003 2368 23037
rect 2334 22935 2368 22969
rect 2334 22867 2368 22901
rect 2334 22799 2368 22833
rect 2334 22731 2368 22765
rect 2334 22663 2368 22697
rect 2334 22595 2368 22629
rect 2334 22527 2368 22561
rect 2334 22459 2368 22493
rect 2334 22391 2368 22425
rect 2334 22323 2368 22357
rect 2334 22255 2368 22289
rect 2334 22187 2368 22221
rect 2334 22119 2368 22153
rect 2334 22051 2368 22085
rect 2334 21983 2368 22017
rect 2334 21915 2368 21949
rect 2334 21847 2368 21881
rect 2334 21779 2368 21813
rect 2334 21711 2368 21745
rect 2334 21643 2368 21677
rect 2334 21575 2368 21609
rect 2334 21507 2368 21541
rect 2334 21439 2368 21473
rect 2334 21371 2368 21405
rect 2334 21303 2368 21337
rect 2334 21235 2368 21269
rect 2334 21167 2368 21201
rect 2334 21099 2368 21133
rect 2334 21031 2368 21065
rect 2334 20963 2368 20997
rect 2334 20895 2368 20929
rect 2334 20827 2368 20861
rect 2334 20759 2368 20793
rect 2334 20691 2368 20725
rect 2334 20623 2368 20657
rect 2334 20555 2368 20589
rect 2334 20487 2368 20521
rect 2334 20419 2368 20453
rect 2334 20351 2368 20385
rect 2334 20283 2368 20317
rect 2334 20215 2368 20249
rect 2334 20147 2368 20181
rect 2334 20079 2368 20113
rect 2334 20011 2368 20045
rect 2334 19943 2368 19977
rect 2334 19875 2368 19909
rect 2334 19807 2368 19841
rect 2334 19739 2368 19773
rect 2334 19671 2368 19705
rect 2334 19603 2368 19637
rect 2334 19535 2368 19569
rect 2334 19467 2368 19501
rect 2334 19399 2368 19433
rect 2334 19331 2368 19365
rect 2334 19263 2368 19297
rect 2334 19195 2368 19229
rect 2334 19127 2368 19161
rect 2334 19059 2368 19093
rect 2334 18991 2368 19025
rect 2334 18923 2368 18957
rect 2334 18855 2368 18889
rect 2334 18787 2368 18821
rect 2334 18719 2368 18753
rect 2334 18651 2368 18685
rect 2334 18583 2368 18617
rect 2334 18515 2368 18549
rect 2334 18447 2368 18481
rect 2334 18379 2368 18413
rect 2334 18311 2368 18345
rect 2334 18243 2368 18277
rect 2334 18175 2368 18209
rect 2334 18107 2368 18141
rect 2334 18039 2368 18073
rect 2334 17971 2368 18005
rect 2334 17903 2368 17937
rect 2334 17835 2368 17869
rect 2334 17767 2368 17801
rect 2334 17699 2368 17733
rect 2334 17631 2368 17665
rect 2334 17563 2368 17597
rect 2334 17495 2368 17529
rect 2334 17427 2368 17461
rect 2334 17359 2368 17393
rect 2334 17291 2368 17325
rect 2334 17223 2368 17257
rect 2334 17155 2368 17189
rect 2334 17087 2368 17121
rect 2334 17019 2368 17053
rect 2334 16951 2368 16985
rect 2334 16883 2368 16917
rect 2334 16815 2368 16849
rect 2334 16747 2368 16781
rect 2334 16679 2368 16713
rect 2334 16611 2368 16645
rect 2334 16543 2368 16577
rect 2334 16475 2368 16509
rect 2334 16407 2368 16441
rect 2334 16339 2368 16373
rect 2334 16271 2368 16305
rect 2334 16203 2368 16237
rect 2334 16135 2368 16169
rect 2334 16067 2368 16101
rect 2334 15999 2368 16033
rect 2334 15931 2368 15965
rect 2334 15863 2368 15897
rect 2334 15795 2368 15829
rect 2334 15727 2368 15761
rect 2334 15659 2368 15693
rect 2334 15591 2368 15625
rect 2334 15523 2368 15557
rect 2334 15455 2368 15489
rect 2334 15387 2368 15421
rect 2334 15319 2368 15353
rect 2334 15251 2368 15285
rect 2334 15183 2368 15217
rect 2334 15115 2368 15149
rect 2334 15047 2368 15081
rect 2334 14979 2368 15013
rect 2334 14911 2368 14945
rect 2334 14843 2368 14877
rect 2334 14775 2368 14809
rect 2334 14707 2368 14741
rect 2334 14639 2368 14673
rect 2334 14571 2368 14605
rect 2334 14503 2368 14537
rect 2334 14435 2368 14469
rect 2334 14367 2368 14401
rect 2334 14299 2368 14333
rect 2334 14231 2368 14265
rect 2334 14163 2368 14197
rect 2334 14095 2368 14129
rect 2334 14027 2368 14061
rect 2334 13959 2368 13993
rect 2334 13891 2368 13925
rect 2334 13823 2368 13857
rect 2334 13755 2368 13789
rect 2334 13687 2368 13721
rect 2334 13619 2368 13653
rect 2334 13551 2368 13585
rect 2334 13483 2368 13517
rect 2334 13415 2368 13449
rect 2334 13347 2368 13381
rect 2334 13279 2368 13313
rect 2334 13211 2368 13245
rect 2334 13143 2368 13177
rect 2334 13075 2368 13109
rect 2334 13007 2368 13041
rect 2334 12939 2368 12973
rect 2334 12871 2368 12905
rect 2334 12803 2368 12837
rect 2334 12735 2368 12769
rect 2334 12667 2368 12701
rect 2334 12599 2368 12633
rect 2334 12531 2368 12565
rect 2334 12463 2368 12497
rect 2334 12395 2368 12429
rect 2334 12327 2368 12361
rect 2334 12259 2368 12293
rect 2334 12191 2368 12225
rect 2334 12123 2368 12157
rect 2334 12055 2368 12089
rect 2334 11987 2368 12021
rect 2334 11919 2368 11953
rect 2334 11851 2368 11885
rect 2334 11783 2368 11817
rect 2334 11715 2368 11749
rect 2334 11647 2368 11681
rect 2334 11579 2368 11613
rect 2334 11511 2368 11545
rect 2334 11443 2368 11477
rect 2334 11375 2368 11409
rect 2334 11307 2368 11341
rect 2334 11239 2368 11273
rect 2334 11171 2368 11205
rect 2334 11103 2368 11137
rect 2334 11035 2368 11069
rect 2334 10967 2368 11001
rect 2334 10899 2368 10933
rect 2334 10831 2368 10865
rect 2334 10763 2368 10797
rect 2334 10695 2368 10729
rect 2334 10627 2368 10661
rect 2334 10559 2368 10593
rect 2334 10491 2368 10525
rect 2334 10423 2368 10457
rect 2334 10355 2368 10389
rect 2334 10287 2368 10321
rect 2334 10219 2368 10253
rect 2334 10151 2368 10185
rect 2334 10083 2368 10117
rect 2334 10015 2368 10049
rect 2334 9947 2368 9981
rect 2334 9879 2368 9913
rect 2334 9811 2368 9845
rect 2334 9743 2368 9777
rect 2334 9675 2368 9709
rect 2334 9607 2368 9641
rect 2334 9539 2368 9573
rect 2334 9471 2368 9505
rect 2334 9403 2368 9437
rect 2334 9335 2368 9369
rect 2334 9267 2368 9301
rect 2334 9199 2368 9233
rect 2334 9131 2368 9165
rect 2334 9063 2368 9097
rect 2334 8995 2368 9029
rect 2334 8927 2368 8961
rect 2334 8859 2368 8893
rect 2334 8791 2368 8825
rect 2334 8723 2368 8757
rect 2334 8655 2368 8689
rect 2334 8587 2368 8621
rect 2334 8519 2368 8553
rect 2334 8451 2368 8485
rect 2334 8383 2368 8417
rect 2334 8315 2368 8349
rect 2334 8247 2368 8281
rect 2334 8179 2368 8213
rect 2334 8111 2368 8145
rect 2334 8043 2368 8077
rect 2334 7975 2368 8009
rect 2334 7907 2368 7941
rect 2334 7839 2368 7873
rect 2334 7771 2368 7805
rect 2334 7703 2368 7737
rect 2334 7635 2368 7669
rect 2334 7567 2368 7601
rect 2334 7499 2368 7533
rect 2334 7431 2368 7465
rect 2334 7363 2368 7397
rect 2334 7295 2368 7329
rect 2334 7227 2368 7261
rect 2334 7159 2368 7193
rect 2334 7091 2368 7125
rect 2334 7023 2368 7057
rect 2334 6955 2368 6989
rect 2334 6887 2368 6921
rect 2334 6819 2368 6853
rect 2334 6751 2368 6785
rect 2334 6683 2368 6717
rect 2334 6615 2368 6649
rect 2334 6547 2368 6581
rect 2334 6479 2368 6513
rect 2334 6411 2368 6445
rect 2334 6343 2368 6377
rect 2334 6275 2368 6309
rect 2334 6207 2368 6241
rect 2554 10975 2588 11009
rect 2554 10907 2588 10941
rect 6854 10961 6888 10995
rect 6854 10893 6888 10927
rect 2554 10839 2588 10873
rect 2554 10771 2588 10805
rect 2554 10703 2588 10737
rect 2554 10635 2588 10669
rect 2554 10567 2588 10601
rect 2554 10499 2588 10533
rect 2554 10431 2588 10465
rect 2554 10363 2588 10397
rect 2554 10295 2588 10329
rect 2554 10227 2588 10261
rect 2554 10159 2588 10193
rect 2554 10091 2588 10125
rect 2554 10023 2588 10057
rect 2554 9955 2588 9989
rect 2554 9887 2588 9921
rect 2554 9819 2588 9853
rect 2554 9751 2588 9785
rect 2554 9683 2588 9717
rect 2554 9615 2588 9649
rect 2554 9547 2588 9581
rect 2554 9479 2588 9513
rect 2554 9411 2588 9445
rect 2554 9343 2588 9377
rect 2554 9275 2588 9309
rect 2554 9207 2588 9241
rect 2554 9139 2588 9173
rect 2554 9071 2588 9105
rect 2554 9003 2588 9037
rect 2554 8935 2588 8969
rect 2554 8867 2588 8901
rect 2554 8799 2588 8833
rect 2554 8731 2588 8765
rect 2554 8663 2588 8697
rect 2554 8595 2588 8629
rect 2554 8527 2588 8561
rect 2554 8459 2588 8493
rect 2554 8391 2588 8425
rect 2554 8323 2588 8357
rect 2554 8255 2588 8289
rect 2554 8187 2588 8221
rect 2554 8119 2588 8153
rect 2554 8051 2588 8085
rect 2554 7983 2588 8017
rect 2554 7915 2588 7949
rect 2554 7847 2588 7881
rect 2554 7779 2588 7813
rect 2554 7711 2588 7745
rect 2554 7643 2588 7677
rect 2554 7575 2588 7609
rect 2554 7507 2588 7541
rect 2554 7439 2588 7473
rect 2554 7371 2588 7405
rect 2554 7303 2588 7337
rect 2554 7235 2588 7269
rect 2554 7167 2588 7201
rect 2554 7099 2588 7133
rect 2554 7031 2588 7065
rect 2554 6963 2588 6997
rect 2554 6895 2588 6929
rect 2554 6827 2588 6861
rect 2554 6759 2588 6793
rect 2554 6691 2588 6725
rect 2554 6623 2588 6657
rect 2554 6555 2588 6589
rect 2554 6487 2588 6521
rect 2554 6419 2588 6453
rect 6854 10825 6888 10859
rect 6854 10757 6888 10791
rect 6854 10689 6888 10723
rect 6854 10621 6888 10655
rect 6854 10553 6888 10587
rect 6854 10485 6888 10519
rect 6854 10417 6888 10451
rect 6854 10349 6888 10383
rect 6854 10281 6888 10315
rect 6854 10213 6888 10247
rect 6854 10145 6888 10179
rect 6854 10077 6888 10111
rect 6854 10009 6888 10043
rect 6854 9941 6888 9975
rect 6854 9873 6888 9907
rect 6854 9805 6888 9839
rect 6854 9737 6888 9771
rect 6854 9669 6888 9703
rect 6854 9601 6888 9635
rect 6854 9533 6888 9567
rect 6854 9465 6888 9499
rect 6854 9397 6888 9431
rect 6854 9329 6888 9363
rect 6854 9261 6888 9295
rect 6854 9193 6888 9227
rect 6854 9125 6888 9159
rect 6854 9057 6888 9091
rect 6854 8989 6888 9023
rect 6854 8921 6888 8955
rect 6854 8853 6888 8887
rect 6854 8785 6888 8819
rect 6854 8717 6888 8751
rect 6854 8649 6888 8683
rect 6854 8581 6888 8615
rect 6854 8513 6888 8547
rect 6854 8445 6888 8479
rect 6854 8377 6888 8411
rect 6854 8309 6888 8343
rect 6854 8241 6888 8275
rect 6854 8173 6888 8207
rect 6854 8105 6888 8139
rect 6854 8037 6888 8071
rect 6854 7969 6888 8003
rect 6854 7901 6888 7935
rect 6854 7833 6888 7867
rect 6854 7765 6888 7799
rect 6854 7697 6888 7731
rect 6854 7629 6888 7663
rect 6854 7561 6888 7595
rect 6854 7493 6888 7527
rect 6854 7425 6888 7459
rect 6854 7357 6888 7391
rect 6854 7289 6888 7323
rect 6854 7221 6888 7255
rect 6854 7153 6888 7187
rect 6854 7085 6888 7119
rect 6854 7017 6888 7051
rect 6854 6949 6888 6983
rect 6854 6881 6888 6915
rect 6854 6813 6888 6847
rect 6854 6745 6888 6779
rect 6854 6677 6888 6711
rect 6854 6609 6888 6643
rect 6854 6541 6888 6575
rect 6854 6473 6888 6507
rect 2554 6351 2588 6385
rect 6854 6405 6888 6439
rect 6854 6337 6888 6371
rect 2587 6236 2621 6270
rect 2655 6236 2689 6270
rect 2723 6236 2757 6270
rect 2791 6236 2825 6270
rect 2859 6236 2893 6270
rect 2927 6236 2961 6270
rect 2995 6236 3029 6270
rect 3063 6236 3097 6270
rect 3131 6236 3165 6270
rect 3199 6236 3233 6270
rect 3267 6236 3301 6270
rect 3335 6236 3369 6270
rect 3403 6236 3437 6270
rect 3471 6236 3505 6270
rect 3539 6236 3573 6270
rect 3607 6236 3641 6270
rect 3675 6236 3709 6270
rect 3743 6236 3777 6270
rect 3811 6236 3845 6270
rect 3879 6236 3913 6270
rect 3947 6236 3981 6270
rect 4015 6236 4049 6270
rect 4083 6236 4117 6270
rect 4151 6236 4185 6270
rect 4219 6236 4253 6270
rect 4287 6236 4321 6270
rect 4355 6236 4389 6270
rect 4423 6236 4457 6270
rect 4491 6236 4525 6270
rect 4559 6236 4593 6270
rect 4627 6236 4661 6270
rect 4695 6236 4729 6270
rect 4763 6236 4797 6270
rect 4831 6236 4865 6270
rect 4899 6236 4933 6270
rect 4967 6236 5001 6270
rect 5035 6236 5069 6270
rect 5103 6236 5137 6270
rect 5171 6236 5205 6270
rect 5239 6236 5273 6270
rect 5307 6236 5341 6270
rect 5375 6236 5409 6270
rect 5443 6236 5477 6270
rect 5511 6236 5545 6270
rect 5579 6236 5613 6270
rect 5647 6236 5681 6270
rect 5715 6236 5749 6270
rect 5783 6236 5817 6270
rect 5851 6236 5885 6270
rect 5919 6236 5953 6270
rect 5987 6236 6021 6270
rect 6055 6236 6089 6270
rect 6123 6236 6157 6270
rect 6191 6236 6225 6270
rect 6259 6236 6293 6270
rect 6327 6236 6361 6270
rect 6395 6236 6429 6270
rect 6463 6236 6497 6270
rect 6531 6236 6565 6270
rect 6599 6236 6633 6270
rect 6667 6236 6701 6270
rect 6735 6236 6769 6270
rect 6854 6269 6888 6303
rect 2334 6139 2368 6173
rect 6854 6177 6888 6211
rect 6854 6105 6888 6139
rect 2357 6071 2391 6105
rect 2426 6071 2460 6105
rect 2495 6071 2529 6105
rect 2564 6071 2598 6105
rect 2633 6071 2667 6105
rect 2702 6071 2736 6105
rect 2771 6071 2805 6105
rect 2840 6071 2874 6105
rect 2909 6071 2943 6105
rect 2978 6071 3012 6105
rect 3047 6071 3081 6105
rect 3116 6071 3150 6105
rect 3185 6071 3219 6105
rect 3254 6071 3288 6105
rect 3323 6071 3357 6105
rect 3392 6071 3426 6105
rect 3461 6071 3495 6105
rect 3530 6071 3564 6105
rect 3599 6071 3633 6105
rect 3668 6071 3702 6105
rect 3737 6071 3771 6105
rect 3806 6071 3840 6105
rect 3875 6071 3909 6105
rect 3944 6071 3978 6105
rect 4013 6071 4047 6105
rect 4082 6071 4116 6105
rect 4151 6071 4185 6105
rect 4220 6071 4254 6105
rect 4289 6071 4323 6105
rect 4358 6071 4392 6105
rect 4427 6071 4461 6105
rect 4496 6071 4530 6105
rect 4565 6071 4599 6105
rect 4634 6071 4668 6105
rect 4703 6071 4737 6105
rect 4772 6071 4806 6105
rect 4841 6071 4875 6105
rect 4910 6071 4944 6105
rect 4979 6071 5013 6105
rect 5048 6071 5082 6105
rect 5117 6071 5151 6105
rect 5186 6071 5220 6105
rect 5255 6071 5289 6105
rect 5324 6071 5358 6105
rect 5392 6071 5426 6105
rect 5460 6071 5494 6105
rect 5528 6071 5562 6105
rect 5596 6071 5630 6105
rect 5664 6071 5698 6105
rect 5732 6071 5766 6105
rect 5800 6071 5834 6105
rect 5868 6071 5902 6105
rect 5936 6071 5970 6105
rect 6004 6071 6038 6105
rect 6072 6071 6106 6105
rect 6140 6071 6174 6105
rect 6208 6071 6242 6105
rect 6276 6071 6310 6105
rect 6344 6071 6378 6105
rect 6412 6071 6446 6105
rect 6480 6071 6514 6105
rect 6548 6071 6582 6105
rect 6616 6071 6650 6105
rect 6684 6071 6718 6105
rect 6752 6071 6786 6105
rect 3342 781 3376 815
rect 3342 713 3376 747
rect 3342 645 3376 679
rect 3342 577 3376 611
rect 3342 509 3376 543
rect 3342 441 3376 475
rect 3342 373 3376 407
rect 3342 305 3376 339
rect 3342 237 3376 271
rect 3342 169 3376 203
rect 743 35 777 69
rect 887 68 921 102
rect 955 68 989 102
rect 1023 68 1057 102
rect 1091 68 1125 102
rect 1159 68 1193 102
rect 1227 68 1261 102
rect 1295 68 1329 102
rect 1363 68 1397 102
rect 1431 68 1465 102
rect 1499 68 1533 102
rect 1567 68 1601 102
rect 1635 68 1669 102
rect 1703 68 1737 102
rect 1771 68 1805 102
rect 1839 68 1873 102
rect 1907 68 1941 102
rect 1975 68 2009 102
rect 2043 68 2077 102
rect 2111 68 2145 102
rect 2179 68 2213 102
rect 2247 68 2281 102
rect 2315 68 2349 102
rect 2383 68 2417 102
rect 2451 68 2485 102
rect 2519 68 2553 102
rect 2587 68 2621 102
rect 2655 68 2689 102
rect 2723 68 2757 102
rect 2791 68 2825 102
rect 2859 68 2893 102
rect 2927 68 2961 102
rect 2995 68 3029 102
rect 3063 68 3097 102
rect 3131 68 3165 102
rect 3199 68 3233 102
rect 3267 68 3301 102
rect 3342 101 3376 135
rect 743 -33 777 1
rect 743 -101 777 -67
rect 743 -169 777 -135
rect 743 -237 777 -203
rect 3605 -26 3639 8
rect 3605 -94 3639 -60
rect 3605 -162 3639 -128
rect 3605 -230 3639 -196
rect 743 -305 777 -271
rect 3605 -298 3639 -264
rect 743 -373 777 -339
rect 743 -441 777 -407
rect 743 -509 777 -475
rect 743 -577 777 -543
rect 1714 -399 1748 -365
rect 1861 -399 1895 -365
rect 1929 -399 1963 -365
rect 1997 -399 2031 -365
rect 2065 -399 2099 -365
rect 2133 -399 2167 -365
rect 2201 -399 2235 -365
rect 2269 -399 2303 -365
rect 2337 -399 2371 -365
rect 2405 -399 2439 -365
rect 2473 -399 2507 -365
rect 2541 -399 2575 -365
rect 2609 -399 2643 -365
rect 2677 -399 2711 -365
rect 2745 -399 2779 -365
rect 2813 -399 2847 -365
rect 2881 -399 2915 -365
rect 2949 -399 2983 -365
rect 3017 -399 3051 -365
rect 3085 -399 3119 -365
rect 3153 -399 3187 -365
rect 3221 -399 3255 -365
rect 3289 -399 3323 -365
rect 3357 -399 3391 -365
rect 3425 -399 3459 -365
rect 3493 -399 3527 -365
rect 3605 -366 3639 -332
rect 1681 -494 1715 -460
rect 1681 -562 1715 -528
rect 776 -663 810 -629
rect 844 -663 878 -629
rect 912 -663 946 -629
rect 980 -663 1014 -629
rect 1048 -663 1082 -629
rect 1116 -663 1150 -629
rect 1184 -663 1218 -629
rect 1252 -663 1286 -629
rect 1320 -663 1354 -629
rect 1388 -663 1422 -629
rect 1456 -663 1490 -629
rect 1524 -663 1558 -629
rect 1592 -663 1626 -629
rect 1681 -630 1715 -596
<< poly >>
rect 2905 10748 3705 10820
rect 3761 10748 4561 10820
rect 4881 10748 5681 10820
rect 5737 10748 6537 10820
rect 2905 6491 3705 6566
rect 3761 6491 4561 6566
rect 4881 6491 5681 6566
rect 5737 6491 6537 6566
rect 3693 5442 3712 5508
rect 4866 5442 4885 5508
rect 3693 5436 3793 5442
rect 3849 5436 3949 5442
rect 4005 5436 4105 5442
rect 4161 5436 4261 5442
rect 4317 5436 4417 5442
rect 4473 5436 4573 5442
rect 4629 5436 4729 5442
rect 4785 5436 4885 5442
rect 4941 5492 5237 5508
rect 4941 5458 4970 5492
rect 5004 5458 5038 5492
rect 5072 5458 5106 5492
rect 5140 5458 5174 5492
rect 5208 5458 5237 5492
rect 4941 5442 5237 5458
rect 4941 5436 5061 5442
rect 5117 5436 5237 5442
rect 5293 5492 5495 5508
rect 5293 5458 5309 5492
rect 5343 5458 5377 5492
rect 5411 5458 5445 5492
rect 5479 5458 5495 5492
rect 5293 5442 5495 5458
rect 5293 5436 5493 5442
rect 905 -280 2081 -256
rect 905 -314 943 -280
rect 977 -314 1011 -280
rect 1045 -314 1079 -280
rect 1113 -314 1147 -280
rect 1181 -314 1215 -280
rect 1249 -314 1283 -280
rect 1317 -314 1351 -280
rect 1385 -314 1419 -280
rect 1453 -314 1487 -280
rect 1521 -314 1555 -280
rect 1589 -314 1623 -280
rect 1657 -314 1691 -280
rect 1725 -314 1759 -280
rect 1793 -314 1827 -280
rect 1861 -314 1895 -280
rect 1929 -314 1963 -280
rect 1997 -314 2031 -280
rect 2065 -314 2081 -280
rect 905 -330 2081 -314
rect 2137 -280 2337 -256
rect 2137 -314 2153 -280
rect 2187 -314 2287 -280
rect 2321 -314 2337 -280
rect 2137 -330 2337 -314
rect 2503 -280 2903 -256
rect 2503 -314 2519 -280
rect 2553 -314 2603 -280
rect 2637 -314 2687 -280
rect 2721 -314 2770 -280
rect 2804 -314 2853 -280
rect 2887 -314 2903 -280
rect 2503 -330 2903 -314
rect 2959 -280 3359 -256
rect 2959 -314 2975 -280
rect 3009 -314 3059 -280
rect 3093 -314 3143 -280
rect 3177 -314 3226 -280
rect 3260 -314 3309 -280
rect 3343 -314 3359 -280
rect 2959 -330 3359 -314
rect 905 -338 1025 -330
rect 1081 -338 1201 -330
rect 1257 -338 1377 -330
rect 1433 -338 1553 -330
rect 2287 -639 2421 -623
rect 2287 -673 2303 -639
rect 2337 -673 2371 -639
rect 2405 -673 2421 -639
rect 2287 -689 2421 -673
rect 2527 -639 2687 -623
rect 2527 -673 2543 -639
rect 2577 -673 2637 -639
rect 2671 -673 2687 -639
rect 2311 -694 2471 -689
rect 2527 -694 2687 -673
rect 2743 -639 2903 -623
rect 2743 -673 2759 -639
rect 2793 -673 2853 -639
rect 2887 -673 2903 -639
rect 2743 -694 2903 -673
rect 2959 -639 3119 -623
rect 2959 -673 2975 -639
rect 3009 -673 3069 -639
rect 3103 -673 3119 -639
rect 2959 -694 3119 -673
rect 3175 -639 3335 -623
rect 3175 -673 3191 -639
rect 3225 -673 3285 -639
rect 3319 -673 3335 -639
rect 3175 -694 3335 -673
<< polycont >>
rect 4970 5458 5004 5492
rect 5038 5458 5072 5492
rect 5106 5458 5140 5492
rect 5174 5458 5208 5492
rect 5309 5458 5343 5492
rect 5377 5458 5411 5492
rect 5445 5458 5479 5492
rect 943 -314 977 -280
rect 1011 -314 1045 -280
rect 1079 -314 1113 -280
rect 1147 -314 1181 -280
rect 1215 -314 1249 -280
rect 1283 -314 1317 -280
rect 1351 -314 1385 -280
rect 1419 -314 1453 -280
rect 1487 -314 1521 -280
rect 1555 -314 1589 -280
rect 1623 -314 1657 -280
rect 1691 -314 1725 -280
rect 1759 -314 1793 -280
rect 1827 -314 1861 -280
rect 1895 -314 1929 -280
rect 1963 -314 1997 -280
rect 2031 -314 2065 -280
rect 2153 -314 2187 -280
rect 2287 -314 2321 -280
rect 2519 -314 2553 -280
rect 2603 -314 2637 -280
rect 2687 -314 2721 -280
rect 2770 -314 2804 -280
rect 2853 -314 2887 -280
rect 2975 -314 3009 -280
rect 3059 -314 3093 -280
rect 3143 -314 3177 -280
rect 3226 -314 3260 -280
rect 3309 -314 3343 -280
rect 2303 -673 2337 -639
rect 2371 -673 2405 -639
rect 2543 -673 2577 -639
rect 2637 -673 2671 -639
rect 2759 -673 2793 -639
rect 2853 -673 2887 -639
rect 2975 -673 3009 -639
rect 3069 -673 3103 -639
rect 3191 -673 3225 -639
rect 3285 -673 3319 -639
<< locali >>
rect 67 27869 2369 27870
rect 67 27836 165 27869
rect 67 27802 68 27836
rect 102 27835 165 27836
rect 206 27835 233 27869
rect 278 27835 301 27869
rect 335 27835 369 27869
rect 403 27835 437 27869
rect 471 27835 505 27869
rect 539 27835 573 27869
rect 607 27835 641 27869
rect 675 27835 709 27869
rect 743 27835 777 27869
rect 811 27835 845 27869
rect 879 27835 913 27869
rect 947 27835 981 27869
rect 1015 27835 1049 27869
rect 1083 27835 1117 27869
rect 1151 27835 1185 27869
rect 1219 27835 1253 27869
rect 1287 27835 1321 27869
rect 1355 27835 1389 27869
rect 1423 27835 1457 27869
rect 1491 27835 1525 27869
rect 1559 27835 1593 27869
rect 1627 27835 1661 27869
rect 1707 27835 1729 27869
rect 1779 27835 1797 27869
rect 1851 27835 1865 27869
rect 1923 27835 1998 27869
rect 2032 27835 2066 27869
rect 2100 27835 2134 27869
rect 2168 27835 2202 27869
rect 2236 27835 2369 27869
rect 102 27834 2369 27835
rect 102 27802 103 27834
rect 67 27785 103 27802
rect 67 27734 68 27785
rect 102 27734 103 27785
rect 67 27711 103 27734
rect 67 27666 68 27711
rect 102 27666 103 27711
rect 2333 27797 2369 27834
rect 2333 27763 2334 27797
rect 2368 27763 2369 27797
rect 2333 27729 2369 27763
rect 67 27637 103 27666
rect 67 27598 68 27637
rect 102 27598 103 27637
rect 67 27564 103 27598
rect 67 27529 68 27564
rect 102 27529 103 27564
rect 67 27496 103 27529
rect 67 27455 68 27496
rect 102 27455 103 27496
rect 67 27428 103 27455
rect 67 27381 68 27428
rect 102 27381 103 27428
rect 67 27360 103 27381
rect 67 27308 68 27360
rect 102 27308 103 27360
rect 67 27292 103 27308
rect 67 27235 68 27292
rect 102 27235 103 27292
rect 67 27224 103 27235
rect 67 27162 68 27224
rect 102 27162 103 27224
rect 67 27156 103 27162
rect 67 27089 68 27156
rect 102 27089 103 27156
rect 67 27088 103 27089
rect 67 27054 68 27088
rect 102 27054 103 27088
rect 67 27050 103 27054
rect 67 26986 68 27050
rect 102 26986 103 27050
rect 67 26977 103 26986
rect 67 26918 68 26977
rect 102 26918 103 26977
rect 67 26904 103 26918
rect 67 26850 68 26904
rect 102 26850 103 26904
rect 67 26831 103 26850
rect 67 26782 68 26831
rect 102 26782 103 26831
rect 67 26758 103 26782
rect 67 26714 68 26758
rect 102 26714 103 26758
rect 67 26685 103 26714
rect 67 26646 68 26685
rect 102 26646 103 26685
rect 67 26612 103 26646
rect 67 26578 68 26612
rect 102 26578 103 26612
rect 67 26544 103 26578
rect 67 26505 68 26544
rect 102 26505 103 26544
rect 67 26476 103 26505
rect 67 26432 68 26476
rect 102 26432 103 26476
rect 67 26408 103 26432
rect 67 26359 68 26408
rect 102 26359 103 26408
rect 67 26340 103 26359
rect 67 26286 68 26340
rect 102 26286 103 26340
rect 67 26272 103 26286
rect 67 26213 68 26272
rect 102 26213 103 26272
rect 67 26204 103 26213
rect 67 26140 68 26204
rect 102 26140 103 26204
rect 67 26136 103 26140
rect 67 26102 68 26136
rect 102 26102 103 26136
rect 67 26101 103 26102
rect 67 26034 68 26101
rect 102 26034 103 26101
rect 67 26028 103 26034
rect 67 25966 68 26028
rect 102 25966 103 26028
rect 67 25955 103 25966
rect 67 25898 68 25955
rect 102 25898 103 25955
rect 67 25882 103 25898
rect 67 25830 68 25882
rect 102 25830 103 25882
rect 67 25809 103 25830
rect 67 25762 68 25809
rect 102 25762 103 25809
rect 67 25736 103 25762
rect 67 25702 68 25736
rect 102 25702 103 25736
rect 67 25690 103 25702
rect 256 27680 2180 27707
rect 256 27647 344 27680
rect 256 27613 257 27647
rect 291 27646 344 27647
rect 378 27646 412 27680
rect 446 27646 480 27680
rect 514 27646 548 27680
rect 582 27646 616 27680
rect 650 27646 684 27680
rect 718 27646 752 27680
rect 786 27646 820 27680
rect 854 27646 888 27680
rect 922 27646 956 27680
rect 990 27646 1024 27680
rect 1058 27646 1092 27680
rect 1126 27646 1160 27680
rect 1194 27646 1228 27680
rect 1262 27646 1296 27680
rect 1330 27646 1364 27680
rect 1398 27646 1432 27680
rect 1466 27646 1500 27680
rect 1534 27646 1568 27680
rect 1602 27646 1636 27680
rect 1670 27646 1704 27680
rect 1738 27646 1772 27680
rect 1806 27646 1840 27680
rect 1874 27646 1908 27680
rect 1942 27646 1976 27680
rect 2010 27646 2044 27680
rect 2078 27646 2112 27680
rect 2146 27646 2180 27680
rect 291 27645 2180 27646
rect 291 27613 330 27645
rect 256 27579 330 27613
rect 256 27545 257 27579
rect 291 27545 330 27579
rect 2144 27571 2180 27645
rect 256 27511 330 27545
rect 256 27477 257 27511
rect 291 27477 330 27511
rect 366 27517 382 27563
rect 416 27517 432 27563
rect 366 27495 432 27517
rect 492 27517 508 27563
rect 542 27517 558 27563
rect 492 27495 558 27517
rect 618 27517 634 27563
rect 668 27517 684 27563
rect 618 27495 684 27517
rect 744 27517 760 27563
rect 794 27517 810 27563
rect 744 27495 810 27517
rect 870 27517 886 27563
rect 920 27517 936 27563
rect 870 27495 936 27517
rect 996 27517 1012 27563
rect 1046 27517 1062 27563
rect 996 27495 1062 27517
rect 1122 27517 1138 27563
rect 1172 27517 1188 27563
rect 1122 27495 1188 27517
rect 1248 27517 1264 27563
rect 1298 27517 1314 27563
rect 1248 27495 1314 27517
rect 1374 27517 1390 27563
rect 1424 27517 1440 27563
rect 1374 27495 1440 27517
rect 1500 27517 1516 27563
rect 1550 27517 1566 27563
rect 1500 27495 1566 27517
rect 1626 27517 1642 27563
rect 1676 27517 1692 27563
rect 1626 27495 1692 27517
rect 1752 27517 1768 27563
rect 1802 27517 1818 27563
rect 1752 27495 1818 27517
rect 1878 27517 1894 27563
rect 1928 27517 1944 27563
rect 1878 27495 1944 27517
rect 2004 27517 2020 27563
rect 2054 27517 2070 27563
rect 2004 27495 2070 27517
rect 2144 27537 2145 27571
rect 2179 27537 2180 27571
rect 2144 27503 2180 27537
rect 256 27443 330 27477
rect 382 27479 416 27495
rect 256 27409 257 27443
rect 291 27409 330 27443
rect 366 27445 382 27461
rect 508 27479 542 27495
rect 416 27445 432 27461
rect 366 27433 432 27445
rect 492 27445 508 27461
rect 634 27479 668 27495
rect 542 27445 558 27461
rect 492 27433 558 27445
rect 618 27445 634 27461
rect 760 27479 794 27495
rect 668 27445 684 27461
rect 618 27433 684 27445
rect 744 27445 760 27461
rect 886 27479 920 27495
rect 794 27445 810 27461
rect 744 27433 810 27445
rect 870 27445 886 27461
rect 1012 27479 1046 27495
rect 920 27445 936 27461
rect 870 27433 936 27445
rect 996 27445 1012 27461
rect 1138 27479 1172 27495
rect 1046 27445 1062 27461
rect 996 27433 1062 27445
rect 1122 27445 1138 27461
rect 1264 27479 1298 27495
rect 1172 27445 1188 27461
rect 1122 27433 1188 27445
rect 1248 27445 1264 27461
rect 1390 27479 1424 27495
rect 1298 27445 1314 27461
rect 1248 27433 1314 27445
rect 1374 27445 1390 27461
rect 1516 27479 1550 27495
rect 1424 27445 1440 27461
rect 1374 27433 1440 27445
rect 1500 27445 1516 27461
rect 1642 27479 1676 27495
rect 1550 27445 1566 27461
rect 1500 27433 1566 27445
rect 1626 27445 1642 27461
rect 1768 27479 1802 27495
rect 1676 27445 1692 27461
rect 1626 27433 1692 27445
rect 1752 27445 1768 27461
rect 1894 27479 1928 27495
rect 1802 27445 1818 27461
rect 1752 27433 1818 27445
rect 1878 27445 1894 27461
rect 2020 27479 2054 27495
rect 1928 27445 1944 27461
rect 1878 27433 1944 27445
rect 2004 27445 2020 27461
rect 2144 27469 2145 27503
rect 2179 27469 2180 27503
rect 2054 27445 2070 27461
rect 2004 27433 2070 27445
rect 2144 27435 2180 27469
rect 256 27375 330 27409
rect 256 27341 257 27375
rect 291 27341 330 27375
rect 256 27307 330 27341
rect 256 27273 257 27307
rect 291 27273 330 27307
rect 256 27239 330 27273
rect 256 27205 257 27239
rect 291 27205 330 27239
rect 256 27171 330 27205
rect 256 27137 257 27171
rect 291 27137 330 27171
rect 256 27103 330 27137
rect 256 27069 257 27103
rect 291 27069 330 27103
rect 256 27035 330 27069
rect 256 27001 257 27035
rect 291 27001 330 27035
rect 256 26967 330 27001
rect 256 26933 257 26967
rect 291 26933 330 26967
rect 256 26899 330 26933
rect 256 26865 257 26899
rect 291 26865 330 26899
rect 256 26831 330 26865
rect 256 26797 257 26831
rect 291 26797 330 26831
rect 256 26763 330 26797
rect 256 26729 257 26763
rect 291 26729 330 26763
rect 256 26695 330 26729
rect 256 26661 257 26695
rect 291 26661 330 26695
rect 256 26627 330 26661
rect 256 26593 257 26627
rect 291 26593 330 26627
rect 256 26559 330 26593
rect 256 26525 257 26559
rect 291 26525 330 26559
rect 256 26491 330 26525
rect 256 26457 257 26491
rect 291 26457 330 26491
rect 256 26423 330 26457
rect 256 26389 257 26423
rect 291 26389 330 26423
rect 256 26355 330 26389
rect 256 26321 257 26355
rect 291 26321 330 26355
rect 256 26287 330 26321
rect 256 26253 257 26287
rect 291 26253 330 26287
rect 256 26219 330 26253
rect 256 26185 257 26219
rect 291 26185 330 26219
rect 256 26151 330 26185
rect 256 26117 257 26151
rect 291 26117 330 26151
rect 256 26083 330 26117
rect 256 26049 257 26083
rect 291 26049 330 26083
rect 256 26015 330 26049
rect 256 25981 257 26015
rect 291 25981 330 26015
rect 256 25947 330 25981
rect 256 25913 257 25947
rect 291 25913 330 25947
rect 256 25879 330 25913
rect 256 25845 257 25879
rect 291 25845 330 25879
rect 256 25811 330 25845
rect 256 25777 257 25811
rect 291 25777 330 25811
rect 256 25743 330 25777
rect 256 25709 257 25743
rect 291 25709 330 25743
rect 256 25675 330 25709
rect 256 25641 257 25675
rect 291 25641 330 25675
rect 256 25607 330 25641
rect 256 25573 257 25607
rect 291 25573 330 25607
rect 256 25539 330 25573
rect 256 25505 257 25539
rect 291 25505 330 25539
rect 256 25471 330 25505
rect 256 25437 257 25471
rect 291 25437 330 25471
rect 256 25403 330 25437
rect 256 25369 257 25403
rect 291 25369 330 25403
rect 256 25335 330 25369
rect 256 25301 257 25335
rect 291 25301 330 25335
rect 256 25267 330 25301
rect 256 25233 257 25267
rect 291 25233 330 25267
rect 256 25199 330 25233
rect 256 25165 257 25199
rect 291 25165 330 25199
rect 256 25131 330 25165
rect 256 25097 257 25131
rect 291 25097 330 25131
rect 256 25063 330 25097
rect 256 25029 257 25063
rect 291 25029 330 25063
rect 256 24995 330 25029
rect 256 24961 257 24995
rect 291 24961 330 24995
rect 256 24927 330 24961
rect 256 24893 257 24927
rect 291 24893 330 24927
rect 256 24859 330 24893
rect 256 24825 257 24859
rect 291 24825 330 24859
rect 256 24791 330 24825
rect 256 24757 257 24791
rect 291 24757 330 24791
rect 256 24723 330 24757
rect 256 24689 257 24723
rect 291 24689 330 24723
rect 256 24655 330 24689
rect 256 24621 257 24655
rect 291 24621 330 24655
rect 256 24587 330 24621
rect 256 24553 257 24587
rect 291 24553 330 24587
rect 256 24519 330 24553
rect 256 24485 257 24519
rect 291 24485 330 24519
rect 256 24451 330 24485
rect 256 24417 257 24451
rect 291 24417 330 24451
rect 256 24383 330 24417
rect 256 24349 257 24383
rect 291 24349 330 24383
rect 256 24315 330 24349
rect 256 24281 257 24315
rect 291 24281 330 24315
rect 256 24247 330 24281
rect 256 24213 257 24247
rect 291 24213 330 24247
rect 256 24179 330 24213
rect 256 24145 257 24179
rect 291 24145 330 24179
rect 256 24111 330 24145
rect 256 24077 257 24111
rect 291 24077 330 24111
rect 256 24043 330 24077
rect 256 24009 257 24043
rect 291 24009 330 24043
rect 256 23975 330 24009
rect 256 23941 257 23975
rect 291 23941 330 23975
rect 256 23907 330 23941
rect 256 23873 257 23907
rect 291 23873 330 23907
rect 2144 27401 2145 27435
rect 2179 27401 2180 27435
rect 2144 27367 2180 27401
rect 2144 27333 2145 27367
rect 2179 27333 2180 27367
rect 2144 27299 2180 27333
rect 2144 27265 2145 27299
rect 2179 27265 2180 27299
rect 2144 27231 2180 27265
rect 2144 27197 2145 27231
rect 2179 27197 2180 27231
rect 2144 27163 2180 27197
rect 2144 27129 2145 27163
rect 2179 27129 2180 27163
rect 2144 27095 2180 27129
rect 2144 27061 2145 27095
rect 2179 27061 2180 27095
rect 2144 27027 2180 27061
rect 2144 26993 2145 27027
rect 2179 26993 2180 27027
rect 2144 26959 2180 26993
rect 2144 26925 2145 26959
rect 2179 26925 2180 26959
rect 2144 26891 2180 26925
rect 2144 26857 2145 26891
rect 2179 26857 2180 26891
rect 2144 26823 2180 26857
rect 2144 26789 2145 26823
rect 2179 26789 2180 26823
rect 2144 26755 2180 26789
rect 2144 26721 2145 26755
rect 2179 26721 2180 26755
rect 2144 26687 2180 26721
rect 2144 26653 2145 26687
rect 2179 26653 2180 26687
rect 2144 26619 2180 26653
rect 2144 26585 2145 26619
rect 2179 26585 2180 26619
rect 2144 26551 2180 26585
rect 2144 26517 2145 26551
rect 2179 26517 2180 26551
rect 2144 26483 2180 26517
rect 2144 26449 2145 26483
rect 2179 26449 2180 26483
rect 2144 26415 2180 26449
rect 2144 26381 2145 26415
rect 2179 26381 2180 26415
rect 2144 26347 2180 26381
rect 2144 26313 2145 26347
rect 2179 26313 2180 26347
rect 2144 26279 2180 26313
rect 2144 26245 2145 26279
rect 2179 26245 2180 26279
rect 2144 26211 2180 26245
rect 2144 26177 2145 26211
rect 2179 26177 2180 26211
rect 2144 26143 2180 26177
rect 2144 26109 2145 26143
rect 2179 26109 2180 26143
rect 2144 26075 2180 26109
rect 2144 26041 2145 26075
rect 2179 26041 2180 26075
rect 2144 26007 2180 26041
rect 2144 25973 2145 26007
rect 2179 25973 2180 26007
rect 2144 25939 2180 25973
rect 2144 25905 2145 25939
rect 2179 25905 2180 25939
rect 2144 25871 2180 25905
rect 2144 25837 2145 25871
rect 2179 25837 2180 25871
rect 2144 25803 2180 25837
rect 2144 25769 2145 25803
rect 2179 25769 2180 25803
rect 2144 25735 2180 25769
rect 2144 25701 2145 25735
rect 2179 25701 2180 25735
rect 2144 25667 2180 25701
rect 2144 25633 2145 25667
rect 2179 25633 2180 25667
rect 2144 25599 2180 25633
rect 2144 25565 2145 25599
rect 2179 25565 2180 25599
rect 2144 25531 2180 25565
rect 2144 25497 2145 25531
rect 2179 25497 2180 25531
rect 2144 25463 2180 25497
rect 2144 25429 2145 25463
rect 2179 25429 2180 25463
rect 2144 25395 2180 25429
rect 2144 25361 2145 25395
rect 2179 25361 2180 25395
rect 2144 25327 2180 25361
rect 2144 25293 2145 25327
rect 2179 25293 2180 25327
rect 2144 25259 2180 25293
rect 2144 25225 2145 25259
rect 2179 25225 2180 25259
rect 2144 25191 2180 25225
rect 2144 25157 2145 25191
rect 2179 25157 2180 25191
rect 2144 25123 2180 25157
rect 2144 25089 2145 25123
rect 2179 25089 2180 25123
rect 2144 25055 2180 25089
rect 2144 25021 2145 25055
rect 2179 25021 2180 25055
rect 2144 24987 2180 25021
rect 2144 24953 2145 24987
rect 2179 24953 2180 24987
rect 2144 24919 2180 24953
rect 2144 24885 2145 24919
rect 2179 24885 2180 24919
rect 2144 24851 2180 24885
rect 2144 24817 2145 24851
rect 2179 24817 2180 24851
rect 2144 24783 2180 24817
rect 2144 24749 2145 24783
rect 2179 24749 2180 24783
rect 2144 24715 2180 24749
rect 2144 24681 2145 24715
rect 2179 24681 2180 24715
rect 2144 24647 2180 24681
rect 2144 24613 2145 24647
rect 2179 24613 2180 24647
rect 2144 24579 2180 24613
rect 2144 24545 2145 24579
rect 2179 24545 2180 24579
rect 2144 24511 2180 24545
rect 2144 24477 2145 24511
rect 2179 24477 2180 24511
rect 2144 24443 2180 24477
rect 2144 24409 2145 24443
rect 2179 24409 2180 24443
rect 2144 24375 2180 24409
rect 2144 24341 2145 24375
rect 2179 24341 2180 24375
rect 2144 24307 2180 24341
rect 2144 24273 2145 24307
rect 2179 24273 2180 24307
rect 2144 24239 2180 24273
rect 2144 24205 2145 24239
rect 2179 24205 2180 24239
rect 2144 24171 2180 24205
rect 2144 24137 2145 24171
rect 2179 24137 2180 24171
rect 2144 24103 2180 24137
rect 2144 24069 2145 24103
rect 2179 24069 2180 24103
rect 2144 24035 2180 24069
rect 2144 24001 2145 24035
rect 2179 24001 2180 24035
rect 2144 23967 2180 24001
rect 2144 23933 2145 23967
rect 2179 23933 2180 23967
rect 2144 23899 2180 23933
rect 256 23839 330 23873
rect 366 23862 432 23874
rect 366 23846 382 23862
rect 256 23805 257 23839
rect 291 23805 330 23839
rect 416 23846 432 23862
rect 492 23862 558 23874
rect 492 23846 508 23862
rect 382 23812 416 23828
rect 542 23846 558 23862
rect 618 23862 684 23874
rect 618 23846 634 23862
rect 508 23812 542 23828
rect 668 23846 684 23862
rect 744 23862 810 23874
rect 744 23846 760 23862
rect 634 23812 668 23828
rect 794 23846 810 23862
rect 870 23862 936 23874
rect 870 23846 886 23862
rect 760 23812 794 23828
rect 920 23846 936 23862
rect 996 23862 1062 23874
rect 996 23846 1012 23862
rect 886 23812 920 23828
rect 1046 23846 1062 23862
rect 1122 23862 1188 23874
rect 1122 23846 1138 23862
rect 1012 23812 1046 23828
rect 1172 23846 1188 23862
rect 1248 23862 1314 23874
rect 1248 23846 1264 23862
rect 1138 23812 1172 23828
rect 1298 23846 1314 23862
rect 1374 23862 1440 23874
rect 1374 23846 1390 23862
rect 1264 23812 1298 23828
rect 1424 23846 1440 23862
rect 1500 23862 1566 23874
rect 1500 23846 1516 23862
rect 1390 23812 1424 23828
rect 1550 23846 1566 23862
rect 1626 23862 1692 23874
rect 1626 23846 1642 23862
rect 1516 23812 1550 23828
rect 1676 23846 1692 23862
rect 1752 23862 1818 23874
rect 1752 23846 1768 23862
rect 1642 23812 1676 23828
rect 1802 23846 1818 23862
rect 1878 23862 1944 23874
rect 1878 23846 1894 23862
rect 1768 23812 1802 23828
rect 1928 23846 1944 23862
rect 2004 23862 2070 23874
rect 2004 23846 2020 23862
rect 1894 23812 1928 23828
rect 2054 23846 2070 23862
rect 2144 23865 2145 23899
rect 2179 23865 2180 23899
rect 2020 23812 2054 23828
rect 2144 23831 2180 23865
rect 256 23771 330 23805
rect 256 23737 257 23771
rect 291 23737 330 23771
rect 366 23790 432 23812
rect 366 23744 382 23790
rect 416 23744 432 23790
rect 492 23790 558 23812
rect 492 23744 508 23790
rect 542 23744 558 23790
rect 618 23790 684 23812
rect 618 23744 634 23790
rect 668 23744 684 23790
rect 744 23790 810 23812
rect 744 23744 760 23790
rect 794 23744 810 23790
rect 870 23790 936 23812
rect 870 23744 886 23790
rect 920 23744 936 23790
rect 996 23790 1062 23812
rect 996 23744 1012 23790
rect 1046 23744 1062 23790
rect 1122 23790 1188 23812
rect 1122 23744 1138 23790
rect 1172 23744 1188 23790
rect 1248 23790 1314 23812
rect 1248 23744 1264 23790
rect 1298 23744 1314 23790
rect 1374 23790 1440 23812
rect 1374 23744 1390 23790
rect 1424 23744 1440 23790
rect 1500 23790 1566 23812
rect 1500 23744 1516 23790
rect 1550 23744 1566 23790
rect 1626 23790 1692 23812
rect 1626 23744 1642 23790
rect 1676 23744 1692 23790
rect 1752 23790 1818 23812
rect 1752 23744 1768 23790
rect 1802 23744 1818 23790
rect 1878 23790 1944 23812
rect 1878 23744 1894 23790
rect 1928 23744 1944 23790
rect 2004 23790 2070 23812
rect 2004 23744 2020 23790
rect 2054 23744 2070 23790
rect 2144 23797 2145 23831
rect 2179 23797 2180 23831
rect 2144 23763 2180 23797
rect 256 23703 330 23737
rect 256 23669 257 23703
rect 291 23669 330 23703
rect 256 23635 330 23669
rect 2144 23729 2145 23763
rect 2179 23729 2180 23763
rect 2144 23695 2180 23729
rect 256 23601 257 23635
rect 291 23601 330 23635
rect 256 23567 330 23601
rect 366 23622 382 23668
rect 416 23622 432 23668
rect 366 23600 432 23622
rect 492 23622 508 23668
rect 542 23622 558 23668
rect 492 23600 558 23622
rect 618 23622 634 23668
rect 668 23622 684 23668
rect 618 23600 684 23622
rect 744 23622 760 23668
rect 794 23622 810 23668
rect 744 23600 810 23622
rect 870 23622 886 23668
rect 920 23622 936 23668
rect 870 23600 936 23622
rect 996 23622 1012 23668
rect 1046 23622 1062 23668
rect 996 23600 1062 23622
rect 1122 23622 1138 23668
rect 1172 23622 1188 23668
rect 1122 23600 1188 23622
rect 1248 23622 1264 23668
rect 1298 23622 1314 23668
rect 1248 23600 1314 23622
rect 1374 23622 1390 23668
rect 1424 23622 1440 23668
rect 1374 23600 1440 23622
rect 1500 23622 1516 23668
rect 1550 23622 1566 23668
rect 1500 23600 1566 23622
rect 1626 23622 1642 23668
rect 1676 23622 1692 23668
rect 1626 23600 1692 23622
rect 1752 23622 1768 23668
rect 1802 23622 1818 23668
rect 1752 23600 1818 23622
rect 1878 23622 1894 23668
rect 1928 23622 1944 23668
rect 1878 23600 1944 23622
rect 2004 23622 2020 23668
rect 2054 23622 2070 23668
rect 2004 23600 2070 23622
rect 2144 23661 2145 23695
rect 2179 23661 2180 23695
rect 2144 23627 2180 23661
rect 256 23533 257 23567
rect 291 23533 330 23567
rect 382 23584 416 23600
rect 366 23550 382 23566
rect 508 23584 542 23600
rect 416 23550 432 23566
rect 366 23538 432 23550
rect 492 23550 508 23566
rect 634 23584 668 23600
rect 542 23550 558 23566
rect 492 23538 558 23550
rect 618 23550 634 23566
rect 760 23584 794 23600
rect 668 23550 684 23566
rect 618 23538 684 23550
rect 744 23550 760 23566
rect 886 23584 920 23600
rect 794 23550 810 23566
rect 744 23538 810 23550
rect 870 23550 886 23566
rect 1012 23584 1046 23600
rect 920 23550 936 23566
rect 870 23538 936 23550
rect 996 23550 1012 23566
rect 1138 23584 1172 23600
rect 1046 23550 1062 23566
rect 996 23538 1062 23550
rect 1122 23550 1138 23566
rect 1264 23584 1298 23600
rect 1172 23550 1188 23566
rect 1122 23538 1188 23550
rect 1248 23550 1264 23566
rect 1390 23584 1424 23600
rect 1298 23550 1314 23566
rect 1248 23538 1314 23550
rect 1374 23550 1390 23566
rect 1516 23584 1550 23600
rect 1424 23550 1440 23566
rect 1374 23538 1440 23550
rect 1500 23550 1516 23566
rect 1642 23584 1676 23600
rect 1550 23550 1566 23566
rect 1768 23584 1802 23600
rect 1752 23550 1768 23566
rect 1894 23584 1928 23600
rect 1802 23550 1818 23566
rect 1500 23538 1566 23550
rect 1752 23538 1818 23550
rect 1878 23550 1894 23566
rect 2020 23584 2054 23600
rect 1928 23550 1944 23566
rect 1878 23538 1944 23550
rect 2004 23550 2020 23566
rect 2144 23593 2145 23627
rect 2179 23593 2180 23627
rect 2054 23550 2070 23566
rect 2004 23538 2070 23550
rect 2144 23559 2180 23593
rect 256 23499 330 23533
rect 256 23465 257 23499
rect 291 23465 330 23499
rect 256 23431 330 23465
rect 256 23397 257 23431
rect 291 23397 330 23431
rect 256 23363 330 23397
rect 256 23329 257 23363
rect 291 23329 330 23363
rect 256 23295 330 23329
rect 256 23261 257 23295
rect 291 23261 330 23295
rect 256 23227 330 23261
rect 256 23193 257 23227
rect 291 23193 330 23227
rect 256 23159 330 23193
rect 256 23125 257 23159
rect 291 23125 330 23159
rect 256 23091 330 23125
rect 256 23057 257 23091
rect 291 23057 330 23091
rect 256 23023 330 23057
rect 256 22989 257 23023
rect 291 22989 330 23023
rect 256 22955 330 22989
rect 256 22921 257 22955
rect 291 22921 330 22955
rect 256 22887 330 22921
rect 256 22853 257 22887
rect 291 22853 330 22887
rect 256 22819 330 22853
rect 256 22785 257 22819
rect 291 22785 330 22819
rect 256 22751 330 22785
rect 256 22717 257 22751
rect 291 22717 330 22751
rect 256 22683 330 22717
rect 256 22649 257 22683
rect 291 22649 330 22683
rect 256 22615 330 22649
rect 256 22581 257 22615
rect 291 22581 330 22615
rect 256 22547 330 22581
rect 256 22513 257 22547
rect 291 22513 330 22547
rect 256 22479 330 22513
rect 256 22445 257 22479
rect 291 22445 330 22479
rect 256 22411 330 22445
rect 256 22377 257 22411
rect 291 22377 330 22411
rect 2144 23525 2145 23559
rect 2179 23525 2180 23559
rect 2144 23491 2180 23525
rect 2144 23457 2145 23491
rect 2179 23457 2180 23491
rect 2144 23423 2180 23457
rect 2144 23389 2145 23423
rect 2179 23389 2180 23423
rect 2144 23355 2180 23389
rect 2144 23321 2145 23355
rect 2179 23321 2180 23355
rect 2144 23287 2180 23321
rect 2144 23253 2145 23287
rect 2179 23253 2180 23287
rect 2144 23219 2180 23253
rect 2144 23185 2145 23219
rect 2179 23185 2180 23219
rect 2144 23151 2180 23185
rect 2144 23117 2145 23151
rect 2179 23117 2180 23151
rect 2144 23083 2180 23117
rect 2144 23049 2145 23083
rect 2179 23049 2180 23083
rect 2144 23015 2180 23049
rect 2144 22981 2145 23015
rect 2179 22981 2180 23015
rect 2144 22947 2180 22981
rect 2144 22913 2145 22947
rect 2179 22913 2180 22947
rect 2144 22879 2180 22913
rect 2144 22845 2145 22879
rect 2179 22845 2180 22879
rect 2144 22811 2180 22845
rect 2144 22777 2145 22811
rect 2179 22777 2180 22811
rect 2144 22743 2180 22777
rect 2144 22709 2145 22743
rect 2179 22709 2180 22743
rect 2144 22675 2180 22709
rect 2144 22641 2145 22675
rect 2179 22641 2180 22675
rect 2144 22607 2180 22641
rect 2144 22573 2145 22607
rect 2179 22573 2180 22607
rect 2144 22539 2180 22573
rect 2144 22505 2145 22539
rect 2179 22505 2180 22539
rect 2144 22471 2180 22505
rect 2144 22437 2145 22471
rect 2179 22437 2180 22471
rect 2144 22403 2180 22437
rect 256 22343 330 22377
rect 1374 22391 1440 22403
rect 1374 22375 1390 22391
rect 256 22309 257 22343
rect 291 22309 330 22343
rect 1424 22375 1440 22391
rect 1626 22391 1692 22403
rect 1626 22375 1642 22391
rect 1390 22341 1424 22357
rect 1676 22375 1692 22391
rect 1878 22391 1944 22403
rect 1878 22375 1894 22391
rect 1642 22341 1676 22357
rect 1928 22375 1944 22391
rect 1894 22341 1928 22357
rect 2144 22369 2145 22403
rect 2179 22369 2180 22403
rect 256 22275 330 22309
rect 256 22241 257 22275
rect 291 22241 330 22275
rect 1374 22319 1440 22341
rect 1374 22273 1390 22319
rect 1424 22273 1440 22319
rect 1626 22319 1692 22341
rect 1626 22273 1642 22319
rect 1676 22273 1692 22319
rect 1878 22319 1944 22341
rect 1878 22273 1894 22319
rect 1928 22273 1944 22319
rect 2144 22335 2180 22369
rect 2144 22301 2145 22335
rect 2179 22301 2180 22335
rect 256 22207 330 22241
rect 256 22173 257 22207
rect 291 22173 330 22207
rect 256 22139 330 22173
rect 256 22105 257 22139
rect 291 22105 330 22139
rect 256 22071 330 22105
rect 256 22037 257 22071
rect 291 22037 330 22071
rect 256 22003 330 22037
rect 256 21969 257 22003
rect 291 21969 330 22003
rect 256 21935 330 21969
rect 256 21901 257 21935
rect 291 21901 330 21935
rect 256 21867 330 21901
rect 256 21833 257 21867
rect 291 21833 330 21867
rect 256 21799 330 21833
rect 256 21765 257 21799
rect 291 21765 330 21799
rect 256 21731 330 21765
rect 256 21697 257 21731
rect 291 21697 330 21731
rect 256 21663 330 21697
rect 256 21629 257 21663
rect 291 21629 330 21663
rect 256 21595 330 21629
rect 256 21561 257 21595
rect 291 21561 330 21595
rect 256 21527 330 21561
rect 256 21493 257 21527
rect 291 21493 330 21527
rect 256 21459 330 21493
rect 256 21425 257 21459
rect 291 21425 330 21459
rect 256 21391 330 21425
rect 256 21357 257 21391
rect 291 21357 330 21391
rect 256 21323 330 21357
rect 256 21289 257 21323
rect 291 21289 330 21323
rect 256 21255 330 21289
rect 256 21221 257 21255
rect 291 21221 330 21255
rect 256 21187 330 21221
rect 256 21153 257 21187
rect 291 21153 330 21187
rect 256 21119 330 21153
rect 256 21085 257 21119
rect 291 21085 330 21119
rect 256 21051 330 21085
rect 256 21017 257 21051
rect 291 21017 330 21051
rect 256 20983 330 21017
rect 256 20949 257 20983
rect 291 20949 330 20983
rect 256 20915 330 20949
rect 256 20881 257 20915
rect 291 20881 330 20915
rect 256 20847 330 20881
rect 256 20813 257 20847
rect 291 20813 330 20847
rect 256 20779 330 20813
rect 256 20745 257 20779
rect 291 20745 330 20779
rect 256 20711 330 20745
rect 256 20677 257 20711
rect 291 20677 330 20711
rect 256 20643 330 20677
rect 256 20609 257 20643
rect 291 20609 330 20643
rect 256 20575 330 20609
rect 256 20541 257 20575
rect 291 20541 330 20575
rect 256 20507 330 20541
rect 256 20473 257 20507
rect 291 20473 330 20507
rect 256 20439 330 20473
rect 256 20405 257 20439
rect 291 20405 330 20439
rect 256 20371 330 20405
rect 256 20337 257 20371
rect 291 20337 330 20371
rect 256 20303 330 20337
rect 256 20269 257 20303
rect 291 20269 330 20303
rect 256 20235 330 20269
rect 256 20201 257 20235
rect 291 20201 330 20235
rect 256 20167 330 20201
rect 256 20133 257 20167
rect 291 20133 330 20167
rect 256 20099 330 20133
rect 256 20065 257 20099
rect 291 20065 330 20099
rect 256 20031 330 20065
rect 256 19997 257 20031
rect 291 19997 330 20031
rect 256 19963 330 19997
rect 2144 22267 2180 22301
rect 2144 22233 2145 22267
rect 2179 22233 2180 22267
rect 2144 22199 2180 22233
rect 2144 22165 2145 22199
rect 2179 22165 2180 22199
rect 2144 22131 2180 22165
rect 2144 22097 2145 22131
rect 2179 22097 2180 22131
rect 2144 22063 2180 22097
rect 2144 22029 2145 22063
rect 2179 22029 2180 22063
rect 2144 21995 2180 22029
rect 2144 21961 2145 21995
rect 2179 21961 2180 21995
rect 2144 21927 2180 21961
rect 2144 21893 2145 21927
rect 2179 21893 2180 21927
rect 2144 21859 2180 21893
rect 2144 21825 2145 21859
rect 2179 21825 2180 21859
rect 2144 21791 2180 21825
rect 2144 21757 2145 21791
rect 2179 21757 2180 21791
rect 2144 21723 2180 21757
rect 2144 21689 2145 21723
rect 2179 21689 2180 21723
rect 2144 21655 2180 21689
rect 2144 21621 2145 21655
rect 2179 21621 2180 21655
rect 2144 21587 2180 21621
rect 2144 21553 2145 21587
rect 2179 21553 2180 21587
rect 2144 21519 2180 21553
rect 2144 21485 2145 21519
rect 2179 21485 2180 21519
rect 2144 21451 2180 21485
rect 2144 21417 2145 21451
rect 2179 21417 2180 21451
rect 2144 21383 2180 21417
rect 2144 21349 2145 21383
rect 2179 21349 2180 21383
rect 2144 21315 2180 21349
rect 2144 21281 2145 21315
rect 2179 21281 2180 21315
rect 2144 21247 2180 21281
rect 2144 21213 2145 21247
rect 2179 21213 2180 21247
rect 2144 21179 2180 21213
rect 2144 21145 2145 21179
rect 2179 21145 2180 21179
rect 2144 21111 2180 21145
rect 2144 21077 2145 21111
rect 2179 21077 2180 21111
rect 2144 21043 2180 21077
rect 2144 21009 2145 21043
rect 2179 21009 2180 21043
rect 2144 20975 2180 21009
rect 2144 20941 2145 20975
rect 2179 20941 2180 20975
rect 2144 20907 2180 20941
rect 2144 20873 2145 20907
rect 2179 20873 2180 20907
rect 2144 20839 2180 20873
rect 2144 20805 2145 20839
rect 2179 20805 2180 20839
rect 2144 20771 2180 20805
rect 2144 20737 2145 20771
rect 2179 20737 2180 20771
rect 2144 20703 2180 20737
rect 2144 20669 2145 20703
rect 2179 20669 2180 20703
rect 2144 20635 2180 20669
rect 2144 20601 2145 20635
rect 2179 20601 2180 20635
rect 2144 20567 2180 20601
rect 2144 20533 2145 20567
rect 2179 20533 2180 20567
rect 2144 20499 2180 20533
rect 2144 20465 2145 20499
rect 2179 20465 2180 20499
rect 2144 20431 2180 20465
rect 2144 20397 2145 20431
rect 2179 20397 2180 20431
rect 2144 20363 2180 20397
rect 2144 20329 2145 20363
rect 2179 20329 2180 20363
rect 2144 20295 2180 20329
rect 2144 20261 2145 20295
rect 2179 20261 2180 20295
rect 2144 20227 2180 20261
rect 2144 20193 2145 20227
rect 2179 20193 2180 20227
rect 2144 20159 2180 20193
rect 2144 20125 2145 20159
rect 2179 20125 2180 20159
rect 2144 20091 2180 20125
rect 2144 20057 2145 20091
rect 2179 20057 2180 20091
rect 2144 20023 2180 20057
rect 2144 19989 2145 20023
rect 2179 19989 2180 20023
rect 256 19929 257 19963
rect 291 19929 330 19963
rect 366 19967 432 19979
rect 366 19951 382 19967
rect 256 19895 330 19929
rect 416 19951 432 19967
rect 492 19967 558 19979
rect 492 19951 508 19967
rect 382 19917 416 19933
rect 542 19951 558 19967
rect 618 19967 684 19979
rect 618 19951 634 19967
rect 508 19917 542 19933
rect 668 19951 684 19967
rect 744 19967 810 19979
rect 744 19951 760 19967
rect 634 19917 668 19933
rect 794 19951 810 19967
rect 870 19967 936 19979
rect 870 19951 886 19967
rect 760 19917 794 19933
rect 920 19951 936 19967
rect 996 19967 1062 19979
rect 996 19951 1012 19967
rect 886 19917 920 19933
rect 1046 19951 1062 19967
rect 1122 19967 1188 19979
rect 1122 19951 1138 19967
rect 1012 19917 1046 19933
rect 1172 19951 1188 19967
rect 1248 19967 1314 19979
rect 1248 19951 1264 19967
rect 1138 19917 1172 19933
rect 1298 19951 1314 19967
rect 1500 19967 1566 19979
rect 1500 19951 1516 19967
rect 1264 19917 1298 19933
rect 1550 19951 1566 19967
rect 1752 19967 1818 19979
rect 1752 19951 1768 19967
rect 1516 19917 1550 19933
rect 1802 19951 1818 19967
rect 2004 19967 2070 19979
rect 2004 19951 2020 19967
rect 1768 19917 1802 19933
rect 2054 19951 2070 19967
rect 2144 19955 2180 19989
rect 2020 19917 2054 19933
rect 2144 19921 2145 19955
rect 2179 19921 2180 19955
rect 256 19861 257 19895
rect 291 19861 330 19895
rect 256 19827 330 19861
rect 366 19895 432 19917
rect 366 19849 382 19895
rect 416 19849 432 19895
rect 492 19895 558 19917
rect 492 19849 508 19895
rect 542 19849 558 19895
rect 618 19895 684 19917
rect 618 19849 634 19895
rect 668 19849 684 19895
rect 744 19895 810 19917
rect 744 19849 760 19895
rect 794 19849 810 19895
rect 870 19895 936 19917
rect 870 19849 886 19895
rect 920 19849 936 19895
rect 996 19895 1062 19917
rect 996 19849 1012 19895
rect 1046 19849 1062 19895
rect 1122 19895 1188 19917
rect 1122 19849 1138 19895
rect 1172 19849 1188 19895
rect 1248 19895 1314 19917
rect 1248 19849 1264 19895
rect 1298 19849 1314 19895
rect 1500 19895 1566 19917
rect 1500 19849 1516 19895
rect 1550 19849 1566 19895
rect 1752 19895 1818 19917
rect 1752 19849 1768 19895
rect 1802 19849 1818 19895
rect 2004 19895 2070 19917
rect 2004 19849 2020 19895
rect 2054 19849 2070 19895
rect 2144 19887 2180 19921
rect 2144 19853 2145 19887
rect 2179 19853 2180 19887
rect 256 19793 257 19827
rect 291 19793 330 19827
rect 256 19759 330 19793
rect 2144 19819 2180 19853
rect 2144 19785 2145 19819
rect 2179 19785 2180 19819
rect 256 19725 257 19759
rect 291 19725 330 19759
rect 256 19691 330 19725
rect 366 19727 382 19773
rect 416 19727 432 19773
rect 366 19705 432 19727
rect 492 19727 508 19773
rect 542 19727 558 19773
rect 492 19705 558 19727
rect 618 19727 634 19773
rect 668 19727 684 19773
rect 618 19705 684 19727
rect 744 19727 760 19773
rect 794 19727 810 19773
rect 744 19705 810 19727
rect 870 19727 886 19773
rect 920 19727 936 19773
rect 870 19705 936 19727
rect 996 19727 1012 19773
rect 1046 19727 1062 19773
rect 996 19705 1062 19727
rect 1122 19727 1138 19773
rect 1172 19727 1188 19773
rect 1122 19705 1188 19727
rect 1248 19727 1264 19773
rect 1298 19727 1314 19773
rect 1248 19705 1314 19727
rect 1374 19727 1390 19773
rect 1424 19727 1440 19773
rect 1374 19705 1440 19727
rect 1500 19727 1516 19773
rect 1550 19727 1566 19773
rect 1500 19705 1566 19727
rect 1626 19727 1642 19773
rect 1676 19727 1692 19773
rect 1626 19705 1692 19727
rect 1752 19727 1768 19773
rect 1802 19727 1818 19773
rect 1752 19705 1818 19727
rect 1878 19727 1894 19773
rect 1928 19727 1944 19773
rect 1878 19705 1944 19727
rect 2004 19727 2020 19773
rect 2054 19727 2070 19773
rect 2004 19705 2070 19727
rect 2144 19751 2180 19785
rect 2144 19717 2145 19751
rect 2179 19717 2180 19751
rect 256 19657 257 19691
rect 291 19657 330 19691
rect 382 19689 416 19705
rect 256 19623 330 19657
rect 366 19655 382 19671
rect 508 19689 542 19705
rect 416 19655 432 19671
rect 366 19643 432 19655
rect 492 19655 508 19671
rect 634 19689 668 19705
rect 542 19655 558 19671
rect 492 19643 558 19655
rect 618 19655 634 19671
rect 760 19689 794 19705
rect 668 19655 684 19671
rect 618 19643 684 19655
rect 744 19655 760 19671
rect 886 19689 920 19705
rect 794 19655 810 19671
rect 744 19643 810 19655
rect 870 19655 886 19671
rect 1012 19689 1046 19705
rect 920 19655 936 19671
rect 870 19643 936 19655
rect 996 19655 1012 19671
rect 1138 19689 1172 19705
rect 1046 19655 1062 19671
rect 996 19643 1062 19655
rect 1122 19655 1138 19671
rect 1264 19689 1298 19705
rect 1172 19655 1188 19671
rect 1122 19643 1188 19655
rect 1248 19655 1264 19671
rect 1390 19689 1424 19705
rect 1298 19655 1314 19671
rect 1248 19643 1314 19655
rect 1374 19655 1390 19671
rect 1516 19689 1550 19705
rect 1424 19655 1440 19671
rect 1374 19643 1440 19655
rect 1500 19655 1516 19671
rect 1642 19689 1676 19705
rect 1550 19655 1566 19671
rect 1500 19643 1566 19655
rect 1626 19655 1642 19671
rect 1768 19689 1802 19705
rect 1676 19655 1692 19671
rect 1626 19643 1692 19655
rect 1752 19655 1768 19671
rect 1894 19689 1928 19705
rect 1802 19655 1818 19671
rect 1752 19643 1818 19655
rect 1878 19655 1894 19671
rect 2020 19689 2054 19705
rect 1928 19655 1944 19671
rect 1878 19643 1944 19655
rect 2004 19655 2020 19671
rect 2144 19683 2180 19717
rect 2054 19655 2070 19671
rect 2004 19643 2070 19655
rect 2144 19649 2145 19683
rect 2179 19649 2180 19683
rect 256 19589 257 19623
rect 291 19589 330 19623
rect 256 19555 330 19589
rect 256 19521 257 19555
rect 291 19521 330 19555
rect 256 19487 330 19521
rect 256 19453 257 19487
rect 291 19453 330 19487
rect 256 19419 330 19453
rect 256 19385 257 19419
rect 291 19385 330 19419
rect 256 19351 330 19385
rect 256 19317 257 19351
rect 291 19317 330 19351
rect 256 19283 330 19317
rect 256 19249 257 19283
rect 291 19249 330 19283
rect 256 19215 330 19249
rect 256 19181 257 19215
rect 291 19181 330 19215
rect 256 19147 330 19181
rect 256 19113 257 19147
rect 291 19113 330 19147
rect 256 19079 330 19113
rect 256 19045 257 19079
rect 291 19045 330 19079
rect 256 19011 330 19045
rect 256 18977 257 19011
rect 291 18977 330 19011
rect 256 18943 330 18977
rect 256 18909 257 18943
rect 291 18909 330 18943
rect 256 18875 330 18909
rect 256 18841 257 18875
rect 291 18841 330 18875
rect 256 18807 330 18841
rect 256 18773 257 18807
rect 291 18773 330 18807
rect 256 18739 330 18773
rect 256 18705 257 18739
rect 291 18705 330 18739
rect 256 18671 330 18705
rect 256 18637 257 18671
rect 291 18637 330 18671
rect 256 18603 330 18637
rect 256 18569 257 18603
rect 291 18569 330 18603
rect 256 18535 330 18569
rect 256 18501 257 18535
rect 291 18501 330 18535
rect 256 18467 330 18501
rect 256 18433 257 18467
rect 291 18433 330 18467
rect 256 18399 330 18433
rect 256 18365 257 18399
rect 291 18365 330 18399
rect 256 18331 330 18365
rect 256 18297 257 18331
rect 291 18297 330 18331
rect 256 18263 330 18297
rect 256 18229 257 18263
rect 291 18229 330 18263
rect 256 18195 330 18229
rect 256 18161 257 18195
rect 291 18161 330 18195
rect 256 18127 330 18161
rect 256 18093 257 18127
rect 291 18093 330 18127
rect 256 18059 330 18093
rect 256 18025 257 18059
rect 291 18025 330 18059
rect 256 17991 330 18025
rect 256 17957 257 17991
rect 291 17957 330 17991
rect 256 17923 330 17957
rect 256 17889 257 17923
rect 291 17889 330 17923
rect 256 17855 330 17889
rect 256 17821 257 17855
rect 291 17821 330 17855
rect 256 17787 330 17821
rect 256 17753 257 17787
rect 291 17753 330 17787
rect 256 17719 330 17753
rect 256 17685 257 17719
rect 291 17685 330 17719
rect 256 17651 330 17685
rect 256 17617 257 17651
rect 291 17617 330 17651
rect 256 17583 330 17617
rect 256 17549 257 17583
rect 291 17549 330 17583
rect 256 17515 330 17549
rect 256 17481 257 17515
rect 291 17481 330 17515
rect 256 17447 330 17481
rect 256 17413 257 17447
rect 291 17413 330 17447
rect 256 17379 330 17413
rect 256 17345 257 17379
rect 291 17345 330 17379
rect 256 17311 330 17345
rect 256 17277 257 17311
rect 291 17277 330 17311
rect 256 17243 330 17277
rect 256 17209 257 17243
rect 291 17209 330 17243
rect 256 17175 330 17209
rect 256 17141 257 17175
rect 291 17141 330 17175
rect 256 17107 330 17141
rect 256 17073 257 17107
rect 291 17073 330 17107
rect 256 17039 330 17073
rect 256 17005 257 17039
rect 291 17005 330 17039
rect 256 16971 330 17005
rect 256 16937 257 16971
rect 291 16937 330 16971
rect 256 16903 330 16937
rect 256 16869 257 16903
rect 291 16869 330 16903
rect 256 16835 330 16869
rect 256 16801 257 16835
rect 291 16801 330 16835
rect 256 16767 330 16801
rect 256 16733 257 16767
rect 291 16733 330 16767
rect 256 16699 330 16733
rect 256 16665 257 16699
rect 291 16665 330 16699
rect 256 16631 330 16665
rect 256 16597 257 16631
rect 291 16597 330 16631
rect 256 16563 330 16597
rect 256 16529 257 16563
rect 291 16529 330 16563
rect 256 16495 330 16529
rect 256 16461 257 16495
rect 291 16461 330 16495
rect 256 16427 330 16461
rect 256 16393 257 16427
rect 291 16393 330 16427
rect 256 16359 330 16393
rect 256 16325 257 16359
rect 291 16325 330 16359
rect 256 16291 330 16325
rect 256 16257 257 16291
rect 291 16257 330 16291
rect 256 16223 330 16257
rect 256 16189 257 16223
rect 291 16189 330 16223
rect 256 16155 330 16189
rect 256 16121 257 16155
rect 291 16121 330 16155
rect 256 16087 330 16121
rect 256 16053 257 16087
rect 291 16053 330 16087
rect 2144 19615 2180 19649
rect 2144 19581 2145 19615
rect 2179 19581 2180 19615
rect 2144 19547 2180 19581
rect 2144 19513 2145 19547
rect 2179 19513 2180 19547
rect 2144 19479 2180 19513
rect 2144 19445 2145 19479
rect 2179 19445 2180 19479
rect 2144 19411 2180 19445
rect 2144 19377 2145 19411
rect 2179 19377 2180 19411
rect 2144 19343 2180 19377
rect 2144 19309 2145 19343
rect 2179 19309 2180 19343
rect 2144 19275 2180 19309
rect 2144 19241 2145 19275
rect 2179 19241 2180 19275
rect 2144 19207 2180 19241
rect 2144 19173 2145 19207
rect 2179 19173 2180 19207
rect 2144 19139 2180 19173
rect 2144 19105 2145 19139
rect 2179 19105 2180 19139
rect 2144 19071 2180 19105
rect 2144 19037 2145 19071
rect 2179 19037 2180 19071
rect 2144 19003 2180 19037
rect 2144 18969 2145 19003
rect 2179 18969 2180 19003
rect 2144 18935 2180 18969
rect 2144 18901 2145 18935
rect 2179 18901 2180 18935
rect 2144 18867 2180 18901
rect 2144 18833 2145 18867
rect 2179 18833 2180 18867
rect 2144 18799 2180 18833
rect 2144 18765 2145 18799
rect 2179 18765 2180 18799
rect 2144 18731 2180 18765
rect 2144 18697 2145 18731
rect 2179 18697 2180 18731
rect 2144 18663 2180 18697
rect 2144 18629 2145 18663
rect 2179 18629 2180 18663
rect 2144 18595 2180 18629
rect 2144 18561 2145 18595
rect 2179 18561 2180 18595
rect 2144 18527 2180 18561
rect 2144 18493 2145 18527
rect 2179 18493 2180 18527
rect 2144 18459 2180 18493
rect 2144 18425 2145 18459
rect 2179 18425 2180 18459
rect 2144 18391 2180 18425
rect 2144 18357 2145 18391
rect 2179 18357 2180 18391
rect 2144 18323 2180 18357
rect 2144 18289 2145 18323
rect 2179 18289 2180 18323
rect 2144 18255 2180 18289
rect 2144 18221 2145 18255
rect 2179 18221 2180 18255
rect 2144 18187 2180 18221
rect 2144 18153 2145 18187
rect 2179 18153 2180 18187
rect 2144 18119 2180 18153
rect 2144 18085 2145 18119
rect 2179 18085 2180 18119
rect 2144 18051 2180 18085
rect 2144 18017 2145 18051
rect 2179 18017 2180 18051
rect 2144 17983 2180 18017
rect 2144 17949 2145 17983
rect 2179 17949 2180 17983
rect 2144 17915 2180 17949
rect 2144 17881 2145 17915
rect 2179 17881 2180 17915
rect 2144 17847 2180 17881
rect 2144 17813 2145 17847
rect 2179 17813 2180 17847
rect 2144 17779 2180 17813
rect 2144 17745 2145 17779
rect 2179 17745 2180 17779
rect 2144 17711 2180 17745
rect 2144 17677 2145 17711
rect 2179 17677 2180 17711
rect 2144 17643 2180 17677
rect 2144 17609 2145 17643
rect 2179 17609 2180 17643
rect 2144 17575 2180 17609
rect 2144 17541 2145 17575
rect 2179 17541 2180 17575
rect 2144 17507 2180 17541
rect 2144 17473 2145 17507
rect 2179 17473 2180 17507
rect 2144 17439 2180 17473
rect 2144 17405 2145 17439
rect 2179 17405 2180 17439
rect 2144 17371 2180 17405
rect 2144 17337 2145 17371
rect 2179 17337 2180 17371
rect 2144 17303 2180 17337
rect 2144 17269 2145 17303
rect 2179 17269 2180 17303
rect 2144 17235 2180 17269
rect 2144 17201 2145 17235
rect 2179 17201 2180 17235
rect 2144 17167 2180 17201
rect 2144 17133 2145 17167
rect 2179 17133 2180 17167
rect 2144 17099 2180 17133
rect 2144 17065 2145 17099
rect 2179 17065 2180 17099
rect 2144 17031 2180 17065
rect 2144 16997 2145 17031
rect 2179 16997 2180 17031
rect 2144 16963 2180 16997
rect 2144 16929 2145 16963
rect 2179 16929 2180 16963
rect 2144 16895 2180 16929
rect 2144 16861 2145 16895
rect 2179 16861 2180 16895
rect 2144 16827 2180 16861
rect 2144 16793 2145 16827
rect 2179 16793 2180 16827
rect 2144 16759 2180 16793
rect 2144 16725 2145 16759
rect 2179 16725 2180 16759
rect 2144 16691 2180 16725
rect 2144 16657 2145 16691
rect 2179 16657 2180 16691
rect 2144 16623 2180 16657
rect 2144 16589 2145 16623
rect 2179 16589 2180 16623
rect 2144 16555 2180 16589
rect 2144 16521 2145 16555
rect 2179 16521 2180 16555
rect 2144 16487 2180 16521
rect 2144 16453 2145 16487
rect 2179 16453 2180 16487
rect 2144 16419 2180 16453
rect 2144 16385 2145 16419
rect 2179 16385 2180 16419
rect 2144 16351 2180 16385
rect 2144 16317 2145 16351
rect 2179 16317 2180 16351
rect 2144 16283 2180 16317
rect 2144 16249 2145 16283
rect 2179 16249 2180 16283
rect 2144 16215 2180 16249
rect 2144 16181 2145 16215
rect 2179 16181 2180 16215
rect 2144 16147 2180 16181
rect 2144 16113 2145 16147
rect 2179 16113 2180 16147
rect 366 16072 432 16084
rect 366 16056 382 16072
rect 256 16019 330 16053
rect 416 16056 432 16072
rect 492 16072 558 16084
rect 492 16056 508 16072
rect 382 16022 416 16038
rect 542 16056 558 16072
rect 618 16072 684 16084
rect 618 16056 634 16072
rect 508 16022 542 16038
rect 668 16056 684 16072
rect 744 16072 810 16084
rect 744 16056 760 16072
rect 634 16022 668 16038
rect 794 16056 810 16072
rect 870 16072 936 16084
rect 870 16056 886 16072
rect 760 16022 794 16038
rect 920 16056 936 16072
rect 996 16072 1062 16084
rect 996 16056 1012 16072
rect 886 16022 920 16038
rect 1046 16056 1062 16072
rect 1122 16072 1188 16084
rect 1122 16056 1138 16072
rect 1012 16022 1046 16038
rect 1172 16056 1188 16072
rect 1248 16072 1314 16084
rect 1248 16056 1264 16072
rect 1138 16022 1172 16038
rect 1298 16056 1314 16072
rect 1374 16072 1440 16084
rect 1374 16056 1390 16072
rect 1264 16022 1298 16038
rect 1424 16056 1440 16072
rect 1500 16072 1566 16084
rect 1500 16056 1516 16072
rect 1390 16022 1424 16038
rect 1550 16056 1566 16072
rect 1626 16072 1692 16084
rect 1626 16056 1642 16072
rect 1516 16022 1550 16038
rect 1676 16056 1692 16072
rect 1752 16072 1818 16084
rect 1752 16056 1768 16072
rect 1642 16022 1676 16038
rect 1802 16056 1818 16072
rect 1878 16072 1944 16084
rect 1878 16056 1894 16072
rect 1768 16022 1802 16038
rect 1928 16056 1944 16072
rect 2004 16072 2070 16084
rect 2004 16056 2020 16072
rect 1894 16022 1928 16038
rect 2054 16056 2070 16072
rect 2144 16079 2180 16113
rect 2020 16022 2054 16038
rect 2144 16045 2145 16079
rect 2179 16045 2180 16079
rect 256 15985 257 16019
rect 291 15985 330 16019
rect 256 15951 330 15985
rect 366 16000 432 16022
rect 366 15954 382 16000
rect 416 15954 432 16000
rect 492 16000 558 16022
rect 492 15954 508 16000
rect 542 15954 558 16000
rect 618 16000 684 16022
rect 618 15954 634 16000
rect 668 15954 684 16000
rect 744 16000 810 16022
rect 744 15954 760 16000
rect 794 15954 810 16000
rect 870 16000 936 16022
rect 870 15954 886 16000
rect 920 15954 936 16000
rect 996 16000 1062 16022
rect 996 15954 1012 16000
rect 1046 15954 1062 16000
rect 1122 16000 1188 16022
rect 1122 15954 1138 16000
rect 1172 15954 1188 16000
rect 1248 16000 1314 16022
rect 1248 15954 1264 16000
rect 1298 15954 1314 16000
rect 1374 16000 1440 16022
rect 1374 15954 1390 16000
rect 1424 15954 1440 16000
rect 1500 16000 1566 16022
rect 1500 15954 1516 16000
rect 1550 15954 1566 16000
rect 1626 16000 1692 16022
rect 1626 15954 1642 16000
rect 1676 15954 1692 16000
rect 1752 16000 1818 16022
rect 1752 15954 1768 16000
rect 1802 15954 1818 16000
rect 1878 16000 1944 16022
rect 1878 15954 1894 16000
rect 1928 15954 1944 16000
rect 2004 16000 2070 16022
rect 2004 15954 2020 16000
rect 2054 15954 2070 16000
rect 2144 16011 2180 16045
rect 2144 15977 2145 16011
rect 2179 15977 2180 16011
rect 256 15917 257 15951
rect 291 15917 330 15951
rect 256 15883 330 15917
rect 256 15849 257 15883
rect 291 15849 330 15883
rect 2144 15943 2180 15977
rect 2144 15909 2145 15943
rect 2179 15909 2180 15943
rect 256 15815 330 15849
rect 256 15781 257 15815
rect 291 15781 330 15815
rect 366 15832 382 15878
rect 416 15832 432 15878
rect 366 15810 432 15832
rect 492 15832 508 15878
rect 542 15832 558 15878
rect 492 15810 558 15832
rect 618 15832 634 15878
rect 668 15832 684 15878
rect 618 15810 684 15832
rect 744 15832 760 15878
rect 794 15832 810 15878
rect 744 15810 810 15832
rect 870 15832 886 15878
rect 920 15832 936 15878
rect 870 15810 936 15832
rect 996 15832 1012 15878
rect 1046 15832 1062 15878
rect 996 15810 1062 15832
rect 1122 15832 1138 15878
rect 1172 15832 1188 15878
rect 1122 15810 1188 15832
rect 1248 15832 1264 15878
rect 1298 15832 1314 15878
rect 1248 15810 1314 15832
rect 1374 15832 1390 15878
rect 1424 15832 1440 15878
rect 1374 15810 1440 15832
rect 1500 15832 1516 15878
rect 1550 15832 1566 15878
rect 1500 15810 1566 15832
rect 1626 15832 1642 15878
rect 1676 15832 1692 15878
rect 1626 15810 1692 15832
rect 1752 15832 1768 15878
rect 1802 15832 1818 15878
rect 1752 15810 1818 15832
rect 1878 15832 1894 15878
rect 1928 15832 1944 15878
rect 1878 15810 1944 15832
rect 2004 15832 2020 15878
rect 2054 15832 2070 15878
rect 2004 15810 2070 15832
rect 2144 15875 2180 15909
rect 2144 15841 2145 15875
rect 2179 15841 2180 15875
rect 256 15747 330 15781
rect 382 15794 416 15810
rect 366 15760 382 15776
rect 508 15794 542 15810
rect 416 15760 432 15776
rect 366 15748 432 15760
rect 492 15760 508 15776
rect 634 15794 668 15810
rect 542 15760 558 15776
rect 492 15748 558 15760
rect 618 15760 634 15776
rect 760 15794 794 15810
rect 668 15760 684 15776
rect 618 15748 684 15760
rect 744 15760 760 15776
rect 886 15794 920 15810
rect 794 15760 810 15776
rect 744 15748 810 15760
rect 870 15760 886 15776
rect 1012 15794 1046 15810
rect 920 15760 936 15776
rect 870 15748 936 15760
rect 996 15760 1012 15776
rect 1138 15794 1172 15810
rect 1046 15760 1062 15776
rect 996 15748 1062 15760
rect 1122 15760 1138 15776
rect 1264 15794 1298 15810
rect 1172 15760 1188 15776
rect 1122 15748 1188 15760
rect 1248 15760 1264 15776
rect 1390 15794 1424 15810
rect 1298 15760 1314 15776
rect 1248 15748 1314 15760
rect 1374 15760 1390 15776
rect 1516 15794 1550 15810
rect 1424 15760 1440 15776
rect 1374 15748 1440 15760
rect 1500 15760 1516 15776
rect 1642 15794 1676 15810
rect 1550 15760 1566 15776
rect 1500 15748 1566 15760
rect 1626 15760 1642 15776
rect 1768 15794 1802 15810
rect 1676 15760 1692 15776
rect 1626 15748 1692 15760
rect 1752 15760 1768 15776
rect 1894 15794 1928 15810
rect 1802 15760 1818 15776
rect 1752 15748 1818 15760
rect 1878 15760 1894 15776
rect 2020 15794 2054 15810
rect 1928 15760 1944 15776
rect 1878 15748 1944 15760
rect 2004 15760 2020 15776
rect 2144 15807 2180 15841
rect 2054 15760 2070 15776
rect 2004 15748 2070 15760
rect 2144 15773 2145 15807
rect 2179 15773 2180 15807
rect 256 15713 257 15747
rect 291 15713 330 15747
rect 256 15679 330 15713
rect 256 15645 257 15679
rect 291 15645 330 15679
rect 256 15611 330 15645
rect 256 15577 257 15611
rect 291 15577 330 15611
rect 256 15543 330 15577
rect 256 15509 257 15543
rect 291 15509 330 15543
rect 256 15475 330 15509
rect 256 15441 257 15475
rect 291 15441 330 15475
rect 256 15407 330 15441
rect 256 15373 257 15407
rect 291 15373 330 15407
rect 256 15339 330 15373
rect 256 15305 257 15339
rect 291 15305 330 15339
rect 256 15271 330 15305
rect 256 15237 257 15271
rect 291 15237 330 15271
rect 256 15203 330 15237
rect 256 15169 257 15203
rect 291 15169 330 15203
rect 256 15135 330 15169
rect 256 15101 257 15135
rect 291 15101 330 15135
rect 256 15067 330 15101
rect 256 15033 257 15067
rect 291 15033 330 15067
rect 256 14999 330 15033
rect 256 14965 257 14999
rect 291 14965 330 14999
rect 256 14931 330 14965
rect 256 14897 257 14931
rect 291 14897 330 14931
rect 256 14863 330 14897
rect 256 14829 257 14863
rect 291 14829 330 14863
rect 256 14795 330 14829
rect 256 14761 257 14795
rect 291 14761 330 14795
rect 256 14727 330 14761
rect 256 14693 257 14727
rect 291 14693 330 14727
rect 256 14659 330 14693
rect 256 14625 257 14659
rect 291 14625 330 14659
rect 256 14591 330 14625
rect 256 14557 257 14591
rect 291 14557 330 14591
rect 256 14523 330 14557
rect 256 14489 257 14523
rect 291 14489 330 14523
rect 256 14455 330 14489
rect 256 14421 257 14455
rect 291 14421 330 14455
rect 256 14387 330 14421
rect 256 14353 257 14387
rect 291 14353 330 14387
rect 256 14319 330 14353
rect 256 14285 257 14319
rect 291 14285 330 14319
rect 256 14251 330 14285
rect 256 14217 257 14251
rect 291 14217 330 14251
rect 256 14183 330 14217
rect 256 14149 257 14183
rect 291 14149 330 14183
rect 256 14115 330 14149
rect 256 14081 257 14115
rect 291 14081 330 14115
rect 256 14047 330 14081
rect 256 14013 257 14047
rect 291 14013 330 14047
rect 256 13979 330 14013
rect 256 13945 257 13979
rect 291 13945 330 13979
rect 256 13911 330 13945
rect 256 13877 257 13911
rect 291 13877 330 13911
rect 256 13843 330 13877
rect 256 13809 257 13843
rect 291 13809 330 13843
rect 256 13775 330 13809
rect 256 13741 257 13775
rect 291 13741 330 13775
rect 256 13707 330 13741
rect 256 13673 257 13707
rect 291 13673 330 13707
rect 256 13639 330 13673
rect 256 13605 257 13639
rect 291 13605 330 13639
rect 256 13571 330 13605
rect 256 13537 257 13571
rect 291 13537 330 13571
rect 256 13503 330 13537
rect 256 13469 257 13503
rect 291 13469 330 13503
rect 256 13435 330 13469
rect 256 13401 257 13435
rect 291 13401 330 13435
rect 256 13367 330 13401
rect 256 13333 257 13367
rect 291 13333 330 13367
rect 256 13299 330 13333
rect 256 13265 257 13299
rect 291 13265 330 13299
rect 256 13231 330 13265
rect 256 13197 257 13231
rect 291 13197 330 13231
rect 256 13163 330 13197
rect 256 13129 257 13163
rect 291 13129 330 13163
rect 256 13095 330 13129
rect 256 13061 257 13095
rect 291 13061 330 13095
rect 256 13027 330 13061
rect 256 12993 257 13027
rect 291 12993 330 13027
rect 256 12959 330 12993
rect 256 12925 257 12959
rect 291 12925 330 12959
rect 256 12891 330 12925
rect 256 12857 257 12891
rect 291 12857 330 12891
rect 256 12823 330 12857
rect 256 12789 257 12823
rect 291 12789 330 12823
rect 256 12755 330 12789
rect 256 12721 257 12755
rect 291 12721 330 12755
rect 256 12687 330 12721
rect 256 12653 257 12687
rect 291 12653 330 12687
rect 256 12619 330 12653
rect 256 12585 257 12619
rect 291 12585 330 12619
rect 256 12551 330 12585
rect 256 12517 257 12551
rect 291 12517 330 12551
rect 256 12483 330 12517
rect 256 12449 257 12483
rect 291 12449 330 12483
rect 256 12415 330 12449
rect 256 12381 257 12415
rect 291 12381 330 12415
rect 256 12347 330 12381
rect 256 12313 257 12347
rect 291 12313 330 12347
rect 256 12279 330 12313
rect 256 12245 257 12279
rect 291 12245 330 12279
rect 256 12211 330 12245
rect 256 12177 257 12211
rect 291 12177 330 12211
rect 2144 15739 2180 15773
rect 2144 15705 2145 15739
rect 2179 15705 2180 15739
rect 2144 15671 2180 15705
rect 2144 15637 2145 15671
rect 2179 15637 2180 15671
rect 2144 15603 2180 15637
rect 2144 15569 2145 15603
rect 2179 15569 2180 15603
rect 2144 15535 2180 15569
rect 2144 15501 2145 15535
rect 2179 15501 2180 15535
rect 2144 15467 2180 15501
rect 2144 15433 2145 15467
rect 2179 15433 2180 15467
rect 2144 15399 2180 15433
rect 2144 15365 2145 15399
rect 2179 15365 2180 15399
rect 2144 15331 2180 15365
rect 2144 15297 2145 15331
rect 2179 15297 2180 15331
rect 2144 15263 2180 15297
rect 2144 15229 2145 15263
rect 2179 15229 2180 15263
rect 2144 15195 2180 15229
rect 2144 15161 2145 15195
rect 2179 15161 2180 15195
rect 2144 15127 2180 15161
rect 2144 15093 2145 15127
rect 2179 15093 2180 15127
rect 2144 15059 2180 15093
rect 2144 15025 2145 15059
rect 2179 15025 2180 15059
rect 2144 14991 2180 15025
rect 2144 14957 2145 14991
rect 2179 14957 2180 14991
rect 2144 14923 2180 14957
rect 2144 14889 2145 14923
rect 2179 14889 2180 14923
rect 2144 14855 2180 14889
rect 2144 14821 2145 14855
rect 2179 14821 2180 14855
rect 2144 14787 2180 14821
rect 2144 14753 2145 14787
rect 2179 14753 2180 14787
rect 2144 14719 2180 14753
rect 2144 14685 2145 14719
rect 2179 14685 2180 14719
rect 2144 14651 2180 14685
rect 2144 14617 2145 14651
rect 2179 14617 2180 14651
rect 2144 14583 2180 14617
rect 2144 14549 2145 14583
rect 2179 14549 2180 14583
rect 2144 14515 2180 14549
rect 2144 14481 2145 14515
rect 2179 14481 2180 14515
rect 2144 14447 2180 14481
rect 2144 14413 2145 14447
rect 2179 14413 2180 14447
rect 2144 14379 2180 14413
rect 2144 14345 2145 14379
rect 2179 14345 2180 14379
rect 2144 14311 2180 14345
rect 2144 14277 2145 14311
rect 2179 14277 2180 14311
rect 2144 14243 2180 14277
rect 2144 14209 2145 14243
rect 2179 14209 2180 14243
rect 2144 14175 2180 14209
rect 2144 14141 2145 14175
rect 2179 14141 2180 14175
rect 2144 14107 2180 14141
rect 2144 14073 2145 14107
rect 2179 14073 2180 14107
rect 2144 14039 2180 14073
rect 2144 14005 2145 14039
rect 2179 14005 2180 14039
rect 2144 13971 2180 14005
rect 2144 13937 2145 13971
rect 2179 13937 2180 13971
rect 2144 13903 2180 13937
rect 2144 13869 2145 13903
rect 2179 13869 2180 13903
rect 2144 13835 2180 13869
rect 2144 13801 2145 13835
rect 2179 13801 2180 13835
rect 2144 13767 2180 13801
rect 2144 13733 2145 13767
rect 2179 13733 2180 13767
rect 2144 13699 2180 13733
rect 2144 13665 2145 13699
rect 2179 13665 2180 13699
rect 2144 13631 2180 13665
rect 2144 13597 2145 13631
rect 2179 13597 2180 13631
rect 2144 13563 2180 13597
rect 2144 13529 2145 13563
rect 2179 13529 2180 13563
rect 2144 13495 2180 13529
rect 2144 13461 2145 13495
rect 2179 13461 2180 13495
rect 2144 13427 2180 13461
rect 2144 13393 2145 13427
rect 2179 13393 2180 13427
rect 2144 13359 2180 13393
rect 2144 13325 2145 13359
rect 2179 13325 2180 13359
rect 2144 13291 2180 13325
rect 2144 13257 2145 13291
rect 2179 13257 2180 13291
rect 2144 13223 2180 13257
rect 2144 13189 2145 13223
rect 2179 13189 2180 13223
rect 2144 13155 2180 13189
rect 2144 13121 2145 13155
rect 2179 13121 2180 13155
rect 2144 13087 2180 13121
rect 2144 13053 2145 13087
rect 2179 13053 2180 13087
rect 2144 13019 2180 13053
rect 2144 12985 2145 13019
rect 2179 12985 2180 13019
rect 2144 12951 2180 12985
rect 2144 12917 2145 12951
rect 2179 12917 2180 12951
rect 2144 12883 2180 12917
rect 2144 12849 2145 12883
rect 2179 12849 2180 12883
rect 2144 12815 2180 12849
rect 2144 12781 2145 12815
rect 2179 12781 2180 12815
rect 2144 12747 2180 12781
rect 2144 12713 2145 12747
rect 2179 12713 2180 12747
rect 2144 12679 2180 12713
rect 2144 12645 2145 12679
rect 2179 12645 2180 12679
rect 2144 12611 2180 12645
rect 2144 12577 2145 12611
rect 2179 12577 2180 12611
rect 2144 12543 2180 12577
rect 2144 12509 2145 12543
rect 2179 12509 2180 12543
rect 2144 12475 2180 12509
rect 2144 12441 2145 12475
rect 2179 12441 2180 12475
rect 2144 12407 2180 12441
rect 2144 12373 2145 12407
rect 2179 12373 2180 12407
rect 2144 12339 2180 12373
rect 2144 12305 2145 12339
rect 2179 12305 2180 12339
rect 2144 12271 2180 12305
rect 2144 12237 2145 12271
rect 2179 12237 2180 12271
rect 2144 12203 2180 12237
rect 256 12143 330 12177
rect 366 12177 432 12189
rect 366 12161 382 12177
rect 256 12109 257 12143
rect 291 12109 330 12143
rect 416 12161 432 12177
rect 492 12177 558 12189
rect 492 12161 508 12177
rect 382 12127 416 12143
rect 542 12161 558 12177
rect 618 12177 684 12189
rect 618 12161 634 12177
rect 508 12127 542 12143
rect 668 12161 684 12177
rect 744 12177 810 12189
rect 744 12161 760 12177
rect 634 12127 668 12143
rect 794 12161 810 12177
rect 870 12177 936 12189
rect 870 12161 886 12177
rect 760 12127 794 12143
rect 920 12161 936 12177
rect 996 12177 1062 12189
rect 996 12161 1012 12177
rect 886 12127 920 12143
rect 1046 12161 1062 12177
rect 1122 12177 1188 12189
rect 1122 12161 1138 12177
rect 1012 12127 1046 12143
rect 1172 12161 1188 12177
rect 1248 12177 1314 12189
rect 1248 12161 1264 12177
rect 1138 12127 1172 12143
rect 1298 12161 1314 12177
rect 1374 12177 1440 12189
rect 1374 12161 1390 12177
rect 1264 12127 1298 12143
rect 1424 12161 1440 12177
rect 1500 12177 1566 12189
rect 1500 12161 1516 12177
rect 1390 12127 1424 12143
rect 1550 12161 1566 12177
rect 1626 12177 1692 12189
rect 1626 12161 1642 12177
rect 1516 12127 1550 12143
rect 1676 12161 1692 12177
rect 1752 12177 1818 12189
rect 1752 12161 1768 12177
rect 1642 12127 1676 12143
rect 1802 12161 1818 12177
rect 1878 12177 1944 12189
rect 1878 12161 1894 12177
rect 1768 12127 1802 12143
rect 1928 12161 1944 12177
rect 2004 12177 2070 12189
rect 2004 12161 2020 12177
rect 1894 12127 1928 12143
rect 2054 12161 2070 12177
rect 2144 12169 2145 12203
rect 2179 12169 2180 12203
rect 2020 12127 2054 12143
rect 2144 12135 2180 12169
rect 256 12075 330 12109
rect 256 12041 257 12075
rect 291 12041 330 12075
rect 366 12105 432 12127
rect 366 12059 382 12105
rect 416 12059 432 12105
rect 492 12105 558 12127
rect 492 12059 508 12105
rect 542 12059 558 12105
rect 618 12105 684 12127
rect 618 12059 634 12105
rect 668 12059 684 12105
rect 744 12105 810 12127
rect 744 12059 760 12105
rect 794 12059 810 12105
rect 870 12105 936 12127
rect 870 12059 886 12105
rect 920 12059 936 12105
rect 996 12105 1062 12127
rect 996 12059 1012 12105
rect 1046 12059 1062 12105
rect 1122 12105 1188 12127
rect 1122 12059 1138 12105
rect 1172 12059 1188 12105
rect 1248 12105 1314 12127
rect 1248 12059 1264 12105
rect 1298 12059 1314 12105
rect 1374 12105 1440 12127
rect 1374 12059 1390 12105
rect 1424 12059 1440 12105
rect 1500 12105 1566 12127
rect 1500 12059 1516 12105
rect 1550 12059 1566 12105
rect 1626 12105 1692 12127
rect 1626 12059 1642 12105
rect 1676 12059 1692 12105
rect 1752 12105 1818 12127
rect 1752 12059 1768 12105
rect 1802 12059 1818 12105
rect 1878 12105 1944 12127
rect 1878 12059 1894 12105
rect 1928 12059 1944 12105
rect 2004 12105 2070 12127
rect 2004 12059 2020 12105
rect 2054 12059 2070 12105
rect 2144 12101 2145 12135
rect 2179 12101 2180 12135
rect 2144 12067 2180 12101
rect 256 12007 330 12041
rect 256 11973 257 12007
rect 291 11973 330 12007
rect 2144 12033 2145 12067
rect 2179 12033 2180 12067
rect 2144 11999 2180 12033
rect 256 11939 330 11973
rect 256 11905 257 11939
rect 291 11905 330 11939
rect 366 11937 382 11983
rect 416 11937 432 11983
rect 366 11915 432 11937
rect 492 11937 508 11983
rect 542 11937 558 11983
rect 492 11915 558 11937
rect 618 11937 634 11983
rect 668 11937 684 11983
rect 618 11915 684 11937
rect 744 11937 760 11983
rect 794 11937 810 11983
rect 744 11915 810 11937
rect 870 11937 886 11983
rect 920 11937 936 11983
rect 870 11915 936 11937
rect 996 11937 1012 11983
rect 1046 11937 1062 11983
rect 996 11915 1062 11937
rect 1122 11937 1138 11983
rect 1172 11937 1188 11983
rect 1122 11915 1188 11937
rect 1248 11937 1264 11983
rect 1298 11937 1314 11983
rect 1248 11915 1314 11937
rect 1374 11937 1390 11983
rect 1424 11937 1440 11983
rect 1374 11915 1440 11937
rect 1500 11937 1516 11983
rect 1550 11937 1566 11983
rect 1500 11915 1566 11937
rect 1626 11937 1642 11983
rect 1676 11937 1692 11983
rect 1626 11915 1692 11937
rect 1752 11937 1768 11983
rect 1802 11937 1818 11983
rect 1752 11915 1818 11937
rect 1878 11937 1894 11983
rect 1928 11937 1944 11983
rect 1878 11915 1944 11937
rect 2004 11937 2020 11983
rect 2054 11937 2070 11983
rect 2004 11915 2070 11937
rect 2144 11965 2145 11999
rect 2179 11965 2180 11999
rect 2144 11931 2180 11965
rect 256 11871 330 11905
rect 382 11899 416 11915
rect 256 11837 257 11871
rect 291 11837 330 11871
rect 366 11865 382 11881
rect 508 11899 542 11915
rect 416 11865 432 11881
rect 366 11853 432 11865
rect 492 11865 508 11881
rect 634 11899 668 11915
rect 542 11865 558 11881
rect 492 11853 558 11865
rect 618 11865 634 11881
rect 760 11899 794 11915
rect 668 11865 684 11881
rect 618 11853 684 11865
rect 744 11865 760 11881
rect 886 11899 920 11915
rect 794 11865 810 11881
rect 744 11853 810 11865
rect 870 11865 886 11881
rect 1012 11899 1046 11915
rect 920 11865 936 11881
rect 870 11853 936 11865
rect 996 11865 1012 11881
rect 1138 11899 1172 11915
rect 1046 11865 1062 11881
rect 996 11853 1062 11865
rect 1122 11865 1138 11881
rect 1264 11899 1298 11915
rect 1172 11865 1188 11881
rect 1122 11853 1188 11865
rect 1248 11865 1264 11881
rect 1390 11899 1424 11915
rect 1298 11865 1314 11881
rect 1248 11853 1314 11865
rect 1374 11865 1390 11881
rect 1516 11899 1550 11915
rect 1424 11865 1440 11881
rect 1374 11853 1440 11865
rect 1500 11865 1516 11881
rect 1642 11899 1676 11915
rect 1550 11865 1566 11881
rect 1500 11853 1566 11865
rect 1626 11865 1642 11881
rect 1768 11899 1802 11915
rect 1676 11865 1692 11881
rect 1626 11853 1692 11865
rect 1752 11865 1768 11881
rect 1894 11899 1928 11915
rect 1802 11865 1818 11881
rect 1752 11853 1818 11865
rect 1878 11865 1894 11881
rect 2020 11899 2054 11915
rect 1928 11865 1944 11881
rect 1878 11853 1944 11865
rect 2004 11865 2020 11881
rect 2144 11897 2145 11931
rect 2179 11897 2180 11931
rect 2054 11865 2070 11881
rect 2004 11853 2070 11865
rect 2144 11863 2180 11897
rect 256 11803 330 11837
rect 256 11769 257 11803
rect 291 11769 330 11803
rect 256 11735 330 11769
rect 256 11701 257 11735
rect 291 11701 330 11735
rect 256 11667 330 11701
rect 256 11633 257 11667
rect 291 11633 330 11667
rect 256 11599 330 11633
rect 256 11565 257 11599
rect 291 11565 330 11599
rect 256 11531 330 11565
rect 256 11497 257 11531
rect 291 11497 330 11531
rect 256 11463 330 11497
rect 256 11429 257 11463
rect 291 11429 330 11463
rect 256 11395 330 11429
rect 256 11361 257 11395
rect 291 11361 330 11395
rect 256 11327 330 11361
rect 256 11293 257 11327
rect 291 11293 330 11327
rect 256 11259 330 11293
rect 256 11225 257 11259
rect 291 11225 330 11259
rect 256 11191 330 11225
rect 256 11157 257 11191
rect 291 11157 330 11191
rect 256 11123 330 11157
rect 256 11089 257 11123
rect 291 11089 330 11123
rect 256 11055 330 11089
rect 256 11021 257 11055
rect 291 11021 330 11055
rect 256 10987 330 11021
rect 256 10953 257 10987
rect 291 10953 330 10987
rect 256 10919 330 10953
rect 256 10885 257 10919
rect 291 10885 330 10919
rect 256 10851 330 10885
rect 256 10817 257 10851
rect 291 10817 330 10851
rect 256 10783 330 10817
rect 256 10749 257 10783
rect 291 10749 330 10783
rect 256 10715 330 10749
rect 256 10681 257 10715
rect 291 10681 330 10715
rect 256 10647 330 10681
rect 256 10613 257 10647
rect 291 10613 330 10647
rect 256 10579 330 10613
rect 256 10545 257 10579
rect 291 10545 330 10579
rect 256 10511 330 10545
rect 256 10477 257 10511
rect 291 10477 330 10511
rect 256 10443 330 10477
rect 256 10409 257 10443
rect 291 10409 330 10443
rect 256 10375 330 10409
rect 256 10341 257 10375
rect 291 10341 330 10375
rect 256 10307 330 10341
rect 256 10273 257 10307
rect 291 10273 330 10307
rect 256 10239 330 10273
rect 256 10205 257 10239
rect 291 10205 330 10239
rect 256 10171 330 10205
rect 256 10137 257 10171
rect 291 10137 330 10171
rect 256 10103 330 10137
rect 256 10069 257 10103
rect 291 10069 330 10103
rect 256 10035 330 10069
rect 256 10001 257 10035
rect 291 10001 330 10035
rect 256 9967 330 10001
rect 256 9933 257 9967
rect 291 9933 330 9967
rect 256 9899 330 9933
rect 256 9865 257 9899
rect 291 9865 330 9899
rect 256 9831 330 9865
rect 256 9797 257 9831
rect 291 9797 330 9831
rect 256 9763 330 9797
rect 256 9729 257 9763
rect 291 9729 330 9763
rect 256 9695 330 9729
rect 256 9661 257 9695
rect 291 9661 330 9695
rect 256 9627 330 9661
rect 256 9593 257 9627
rect 291 9593 330 9627
rect 256 9559 330 9593
rect 256 9525 257 9559
rect 291 9525 330 9559
rect 256 9491 330 9525
rect 256 9457 257 9491
rect 291 9457 330 9491
rect 256 9423 330 9457
rect 256 9389 257 9423
rect 291 9389 330 9423
rect 256 9355 330 9389
rect 256 9321 257 9355
rect 291 9321 330 9355
rect 256 9287 330 9321
rect 256 9253 257 9287
rect 291 9253 330 9287
rect 256 9219 330 9253
rect 256 9185 257 9219
rect 291 9185 330 9219
rect 256 9151 330 9185
rect 256 9117 257 9151
rect 291 9117 330 9151
rect 256 9083 330 9117
rect 256 9049 257 9083
rect 291 9049 330 9083
rect 256 9015 330 9049
rect 256 8981 257 9015
rect 291 8981 330 9015
rect 256 8947 330 8981
rect 256 8913 257 8947
rect 291 8913 330 8947
rect 256 8879 330 8913
rect 256 8845 257 8879
rect 291 8845 330 8879
rect 256 8811 330 8845
rect 256 8777 257 8811
rect 291 8777 330 8811
rect 256 8743 330 8777
rect 256 8709 257 8743
rect 291 8709 330 8743
rect 256 8675 330 8709
rect 256 8641 257 8675
rect 291 8641 330 8675
rect 256 8607 330 8641
rect 256 8573 257 8607
rect 291 8573 330 8607
rect 256 8539 330 8573
rect 256 8505 257 8539
rect 291 8505 330 8539
rect 256 8471 330 8505
rect 256 8437 257 8471
rect 291 8437 330 8471
rect 256 8403 330 8437
rect 256 8369 257 8403
rect 291 8369 330 8403
rect 256 8335 330 8369
rect 256 8301 257 8335
rect 291 8301 330 8335
rect 256 8267 330 8301
rect 2144 11829 2145 11863
rect 2179 11829 2180 11863
rect 2144 11795 2180 11829
rect 2144 11761 2145 11795
rect 2179 11761 2180 11795
rect 2144 11727 2180 11761
rect 2144 11693 2145 11727
rect 2179 11693 2180 11727
rect 2144 11659 2180 11693
rect 2144 11625 2145 11659
rect 2179 11625 2180 11659
rect 2144 11591 2180 11625
rect 2144 11557 2145 11591
rect 2179 11557 2180 11591
rect 2144 11523 2180 11557
rect 2144 11489 2145 11523
rect 2179 11489 2180 11523
rect 2144 11455 2180 11489
rect 2144 11421 2145 11455
rect 2179 11421 2180 11455
rect 2144 11387 2180 11421
rect 2144 11353 2145 11387
rect 2179 11353 2180 11387
rect 2144 11319 2180 11353
rect 2144 11285 2145 11319
rect 2179 11285 2180 11319
rect 2144 11251 2180 11285
rect 2144 11217 2145 11251
rect 2179 11217 2180 11251
rect 2144 11183 2180 11217
rect 2144 11149 2145 11183
rect 2179 11149 2180 11183
rect 2144 11115 2180 11149
rect 2144 11081 2145 11115
rect 2179 11081 2180 11115
rect 2144 11047 2180 11081
rect 2144 11013 2145 11047
rect 2179 11013 2180 11047
rect 2144 10979 2180 11013
rect 2144 10945 2145 10979
rect 2179 10945 2180 10979
rect 2144 10911 2180 10945
rect 2144 10877 2145 10911
rect 2179 10877 2180 10911
rect 2144 10843 2180 10877
rect 2144 10809 2145 10843
rect 2179 10809 2180 10843
rect 2144 10775 2180 10809
rect 2144 10741 2145 10775
rect 2179 10741 2180 10775
rect 2144 10707 2180 10741
rect 2144 10673 2145 10707
rect 2179 10673 2180 10707
rect 2144 10639 2180 10673
rect 2144 10605 2145 10639
rect 2179 10605 2180 10639
rect 2144 10571 2180 10605
rect 2144 10537 2145 10571
rect 2179 10537 2180 10571
rect 2144 10503 2180 10537
rect 2144 10469 2145 10503
rect 2179 10469 2180 10503
rect 2144 10435 2180 10469
rect 2144 10401 2145 10435
rect 2179 10401 2180 10435
rect 2144 10367 2180 10401
rect 2144 10333 2145 10367
rect 2179 10333 2180 10367
rect 2144 10299 2180 10333
rect 2144 10265 2145 10299
rect 2179 10265 2180 10299
rect 2144 10231 2180 10265
rect 2144 10197 2145 10231
rect 2179 10197 2180 10231
rect 2144 10163 2180 10197
rect 2144 10129 2145 10163
rect 2179 10129 2180 10163
rect 2144 10095 2180 10129
rect 2144 10061 2145 10095
rect 2179 10061 2180 10095
rect 2144 10027 2180 10061
rect 2144 9993 2145 10027
rect 2179 9993 2180 10027
rect 2144 9959 2180 9993
rect 2144 9925 2145 9959
rect 2179 9925 2180 9959
rect 2144 9891 2180 9925
rect 2144 9857 2145 9891
rect 2179 9857 2180 9891
rect 2144 9823 2180 9857
rect 2144 9789 2145 9823
rect 2179 9789 2180 9823
rect 2144 9755 2180 9789
rect 2144 9721 2145 9755
rect 2179 9721 2180 9755
rect 2144 9687 2180 9721
rect 2144 9653 2145 9687
rect 2179 9653 2180 9687
rect 2144 9619 2180 9653
rect 2144 9585 2145 9619
rect 2179 9585 2180 9619
rect 2144 9551 2180 9585
rect 2144 9517 2145 9551
rect 2179 9517 2180 9551
rect 2144 9483 2180 9517
rect 2144 9449 2145 9483
rect 2179 9449 2180 9483
rect 2144 9415 2180 9449
rect 2144 9381 2145 9415
rect 2179 9381 2180 9415
rect 2144 9347 2180 9381
rect 2144 9313 2145 9347
rect 2179 9313 2180 9347
rect 2144 9279 2180 9313
rect 2144 9245 2145 9279
rect 2179 9245 2180 9279
rect 2144 9211 2180 9245
rect 2144 9177 2145 9211
rect 2179 9177 2180 9211
rect 2144 9143 2180 9177
rect 2144 9109 2145 9143
rect 2179 9109 2180 9143
rect 2144 9075 2180 9109
rect 2144 9041 2145 9075
rect 2179 9041 2180 9075
rect 2144 9007 2180 9041
rect 2144 8973 2145 9007
rect 2179 8973 2180 9007
rect 2144 8939 2180 8973
rect 2144 8905 2145 8939
rect 2179 8905 2180 8939
rect 2144 8871 2180 8905
rect 2144 8837 2145 8871
rect 2179 8837 2180 8871
rect 2144 8803 2180 8837
rect 2144 8769 2145 8803
rect 2179 8769 2180 8803
rect 2144 8735 2180 8769
rect 2144 8701 2145 8735
rect 2179 8701 2180 8735
rect 2144 8667 2180 8701
rect 2144 8633 2145 8667
rect 2179 8633 2180 8667
rect 2144 8599 2180 8633
rect 2144 8565 2145 8599
rect 2179 8565 2180 8599
rect 2144 8531 2180 8565
rect 2144 8497 2145 8531
rect 2179 8497 2180 8531
rect 2144 8463 2180 8497
rect 2144 8429 2145 8463
rect 2179 8429 2180 8463
rect 2144 8395 2180 8429
rect 2144 8361 2145 8395
rect 2179 8361 2180 8395
rect 2144 8327 2180 8361
rect 256 8233 257 8267
rect 291 8233 330 8267
rect 366 8282 432 8294
rect 366 8266 382 8282
rect 256 8199 330 8233
rect 416 8266 432 8282
rect 492 8282 558 8294
rect 492 8266 508 8282
rect 382 8232 416 8248
rect 542 8266 558 8282
rect 618 8282 684 8294
rect 618 8266 634 8282
rect 508 8232 542 8248
rect 668 8266 684 8282
rect 744 8282 810 8294
rect 744 8266 760 8282
rect 634 8232 668 8248
rect 794 8266 810 8282
rect 870 8282 936 8294
rect 870 8266 886 8282
rect 760 8232 794 8248
rect 920 8266 936 8282
rect 996 8282 1062 8294
rect 996 8266 1012 8282
rect 886 8232 920 8248
rect 1046 8266 1062 8282
rect 1122 8282 1188 8294
rect 1122 8266 1138 8282
rect 1012 8232 1046 8248
rect 1172 8266 1188 8282
rect 1248 8282 1314 8294
rect 1248 8266 1264 8282
rect 1138 8232 1172 8248
rect 1298 8266 1314 8282
rect 1374 8282 1440 8294
rect 1374 8266 1390 8282
rect 1264 8232 1298 8248
rect 1424 8266 1440 8282
rect 1500 8282 1566 8294
rect 1500 8266 1516 8282
rect 1390 8232 1424 8248
rect 1550 8266 1566 8282
rect 1626 8282 1692 8294
rect 1626 8266 1642 8282
rect 1516 8232 1550 8248
rect 1676 8266 1692 8282
rect 1752 8282 1818 8294
rect 1752 8266 1768 8282
rect 1642 8232 1676 8248
rect 1802 8266 1818 8282
rect 1878 8282 1944 8294
rect 1878 8266 1894 8282
rect 1768 8232 1802 8248
rect 1928 8266 1944 8282
rect 2004 8266 2070 8294
rect 2144 8293 2145 8327
rect 2179 8293 2180 8327
rect 1894 8232 1928 8248
rect 2144 8259 2180 8293
rect 256 8165 257 8199
rect 291 8165 330 8199
rect 256 8131 330 8165
rect 366 8210 432 8232
rect 366 8164 382 8210
rect 416 8164 432 8210
rect 492 8210 558 8232
rect 492 8164 508 8210
rect 542 8164 558 8210
rect 618 8210 684 8232
rect 618 8164 634 8210
rect 668 8164 684 8210
rect 744 8210 810 8232
rect 744 8164 760 8210
rect 794 8164 810 8210
rect 870 8210 936 8232
rect 870 8164 886 8210
rect 920 8164 936 8210
rect 996 8210 1062 8232
rect 996 8164 1012 8210
rect 1046 8164 1062 8210
rect 1122 8210 1188 8232
rect 1122 8164 1138 8210
rect 1172 8164 1188 8210
rect 1248 8210 1314 8232
rect 1248 8164 1264 8210
rect 1298 8164 1314 8210
rect 1374 8210 1440 8232
rect 1374 8164 1390 8210
rect 1424 8164 1440 8210
rect 1500 8210 1566 8232
rect 1500 8164 1516 8210
rect 1550 8164 1566 8210
rect 1626 8210 1692 8232
rect 1626 8164 1642 8210
rect 1676 8164 1692 8210
rect 1752 8210 1818 8232
rect 1752 8164 1768 8210
rect 1802 8164 1818 8210
rect 1878 8210 1944 8232
rect 1878 8164 1894 8210
rect 1928 8164 1944 8210
rect 2004 8198 2070 8232
rect 2004 8164 2020 8198
rect 2054 8164 2070 8198
rect 2144 8225 2145 8259
rect 2179 8225 2180 8259
rect 2144 8191 2180 8225
rect 256 8097 257 8131
rect 291 8097 330 8131
rect 256 8063 330 8097
rect 1752 8088 1818 8164
rect 2144 8157 2145 8191
rect 2179 8157 2180 8191
rect 2144 8123 2180 8157
rect 2144 8089 2145 8123
rect 2179 8089 2180 8123
rect 256 8029 257 8063
rect 291 8029 330 8063
rect 256 7995 330 8029
rect 366 8042 382 8088
rect 416 8042 432 8088
rect 366 8020 432 8042
rect 492 8042 508 8088
rect 542 8042 558 8088
rect 492 8020 558 8042
rect 618 8042 634 8088
rect 668 8042 684 8088
rect 618 8020 684 8042
rect 744 8042 760 8088
rect 794 8042 810 8088
rect 744 8020 810 8042
rect 870 8042 886 8088
rect 920 8042 936 8088
rect 870 8020 936 8042
rect 996 8042 1012 8088
rect 1046 8042 1062 8088
rect 996 8020 1062 8042
rect 1122 8042 1138 8088
rect 1172 8042 1188 8088
rect 1122 8020 1188 8042
rect 1248 8042 1264 8088
rect 1298 8042 1314 8088
rect 1248 8020 1314 8042
rect 1374 8042 1390 8088
rect 1424 8042 1440 8088
rect 1374 8020 1440 8042
rect 1500 8042 1516 8088
rect 1550 8042 1566 8088
rect 1500 8020 1566 8042
rect 1626 8042 1642 8088
rect 1676 8042 1692 8088
rect 1626 8020 1692 8042
rect 1752 8054 1768 8088
rect 1802 8054 1818 8088
rect 256 7961 257 7995
rect 291 7961 330 7995
rect 382 8004 416 8020
rect 256 7927 330 7961
rect 366 7970 382 7986
rect 508 8004 542 8020
rect 416 7970 432 7986
rect 366 7958 432 7970
rect 492 7970 508 7986
rect 634 8004 668 8020
rect 542 7970 558 7986
rect 492 7958 558 7970
rect 618 7970 634 7986
rect 760 8004 794 8020
rect 668 7970 684 7986
rect 618 7958 684 7970
rect 744 7970 760 7986
rect 886 8004 920 8020
rect 794 7970 810 7986
rect 744 7958 810 7970
rect 870 7970 886 7986
rect 1012 8004 1046 8020
rect 920 7970 936 7986
rect 870 7958 936 7970
rect 996 7970 1012 7986
rect 1138 8004 1172 8020
rect 1046 7970 1062 7986
rect 996 7958 1062 7970
rect 1122 7970 1138 7986
rect 1264 8004 1298 8020
rect 1172 7970 1188 7986
rect 1122 7958 1188 7970
rect 1248 7970 1264 7986
rect 1390 8004 1424 8020
rect 1298 7970 1314 7986
rect 1248 7958 1314 7970
rect 1374 7970 1390 7986
rect 1516 8004 1550 8020
rect 1424 7970 1440 7986
rect 1374 7958 1440 7970
rect 1500 7970 1516 7986
rect 1642 8004 1676 8020
rect 1550 7970 1566 7986
rect 1500 7958 1566 7970
rect 1626 7970 1642 7986
rect 1752 7986 1818 8054
rect 1878 8054 1894 8088
rect 1928 8054 1944 8088
rect 1878 7988 1944 8054
rect 1676 7970 1692 7986
rect 1626 7958 1692 7970
rect 256 7893 257 7927
rect 291 7893 330 7927
rect 256 7859 330 7893
rect 1878 7954 1894 7988
rect 1928 7954 1944 7988
rect 1878 7916 1944 7954
rect 1878 7882 1894 7916
rect 1928 7882 1944 7916
rect 1878 7876 1944 7882
rect 2144 8055 2180 8089
rect 2144 8021 2145 8055
rect 2179 8021 2180 8055
rect 2144 7987 2180 8021
rect 2144 7953 2145 7987
rect 2179 7953 2180 7987
rect 2144 7919 2180 7953
rect 2144 7885 2145 7919
rect 2179 7885 2180 7919
rect 256 7825 257 7859
rect 291 7825 330 7859
rect 256 7791 330 7825
rect 256 7757 257 7791
rect 291 7757 330 7791
rect 256 7723 330 7757
rect 256 7689 257 7723
rect 291 7689 330 7723
rect 256 7655 330 7689
rect 256 7621 257 7655
rect 291 7621 330 7655
rect 256 7587 330 7621
rect 256 7553 257 7587
rect 291 7553 330 7587
rect 256 7519 330 7553
rect 256 7485 257 7519
rect 291 7485 330 7519
rect 256 7451 330 7485
rect 256 7417 257 7451
rect 291 7417 330 7451
rect 256 7383 330 7417
rect 256 7349 257 7383
rect 291 7349 330 7383
rect 256 7315 330 7349
rect 256 7281 257 7315
rect 291 7281 330 7315
rect 256 7247 330 7281
rect 256 7213 257 7247
rect 291 7213 330 7247
rect 256 7179 330 7213
rect 256 7145 257 7179
rect 291 7145 330 7179
rect 256 7111 330 7145
rect 256 7077 257 7111
rect 291 7077 330 7111
rect 256 7043 330 7077
rect 256 7009 257 7043
rect 291 7009 330 7043
rect 256 6975 330 7009
rect 256 6941 257 6975
rect 291 6941 330 6975
rect 256 6907 330 6941
rect 256 6873 257 6907
rect 291 6873 330 6907
rect 256 6797 330 6873
rect 231 6766 330 6797
rect 265 6725 330 6766
rect 231 6694 330 6725
rect 265 6651 330 6694
rect 231 6623 330 6651
rect 265 6577 330 6623
rect 231 6552 330 6577
rect 265 6503 330 6552
rect 231 6481 330 6503
rect 265 6429 330 6481
rect 231 6410 330 6429
rect 265 6355 330 6410
rect 231 6339 330 6355
rect 265 6281 330 6339
rect 231 6268 330 6281
rect 265 6207 330 6268
rect 231 6197 330 6207
rect 265 6133 330 6197
rect 231 6126 330 6133
rect 265 6060 330 6126
rect 231 6055 330 6060
rect 265 5987 330 6055
rect 231 5984 330 5987
rect 265 5950 330 5984
rect 231 5948 330 5950
rect 265 5914 330 5948
rect 231 5913 330 5914
rect 265 5879 330 5913
rect 231 5875 330 5879
rect 265 5808 330 5875
rect 231 5802 330 5808
rect 265 5768 330 5802
rect 231 5729 330 5768
rect 265 5706 330 5729
rect 231 5672 253 5695
rect 287 5672 330 5706
rect 231 5656 330 5672
rect 265 5638 330 5656
rect 231 5604 253 5622
rect 287 5604 330 5638
rect 231 5583 330 5604
rect 265 5570 330 5583
rect 2144 7851 2180 7885
rect 2144 7817 2145 7851
rect 2179 7817 2180 7851
rect 2144 7783 2180 7817
rect 2144 7749 2145 7783
rect 2179 7749 2180 7783
rect 2144 7715 2180 7749
rect 2144 7681 2145 7715
rect 2179 7681 2180 7715
rect 2144 7647 2180 7681
rect 2144 7613 2145 7647
rect 2179 7613 2180 7647
rect 2144 7579 2180 7613
rect 2144 7545 2145 7579
rect 2179 7545 2180 7579
rect 2144 7511 2180 7545
rect 2144 7477 2145 7511
rect 2179 7477 2180 7511
rect 2144 7443 2180 7477
rect 2144 7409 2145 7443
rect 2179 7409 2180 7443
rect 2144 7375 2180 7409
rect 2144 7341 2145 7375
rect 2179 7341 2180 7375
rect 2144 7307 2180 7341
rect 2144 7273 2145 7307
rect 2179 7273 2180 7307
rect 2144 7239 2180 7273
rect 2144 7205 2145 7239
rect 2179 7205 2180 7239
rect 2144 7171 2180 7205
rect 2144 7137 2145 7171
rect 2179 7137 2180 7171
rect 2144 7103 2180 7137
rect 2144 7069 2145 7103
rect 2179 7069 2180 7103
rect 2144 7035 2180 7069
rect 2144 7001 2145 7035
rect 2179 7001 2180 7035
rect 2144 6967 2180 7001
rect 2144 6933 2145 6967
rect 2179 6933 2180 6967
rect 2144 6899 2180 6933
rect 2144 6865 2145 6899
rect 2179 6865 2180 6899
rect 2144 6831 2180 6865
rect 2144 6797 2145 6831
rect 2179 6797 2180 6831
rect 2144 6763 2180 6797
rect 2144 6729 2145 6763
rect 2179 6729 2180 6763
rect 2144 6695 2180 6729
rect 2144 6661 2145 6695
rect 2179 6661 2180 6695
rect 2144 6627 2180 6661
rect 2144 6593 2145 6627
rect 2179 6593 2180 6627
rect 2144 6559 2180 6593
rect 2144 6525 2145 6559
rect 2179 6525 2180 6559
rect 2144 6491 2180 6525
rect 2144 6457 2145 6491
rect 2179 6457 2180 6491
rect 2144 6423 2180 6457
rect 2144 6389 2145 6423
rect 2179 6389 2180 6423
rect 2144 6355 2180 6389
rect 2144 6321 2145 6355
rect 2179 6321 2180 6355
rect 2144 6287 2180 6321
rect 2144 6253 2145 6287
rect 2179 6253 2180 6287
rect 2144 6219 2180 6253
rect 2144 6185 2145 6219
rect 2179 6185 2180 6219
rect 2144 6151 2180 6185
rect 2144 6117 2145 6151
rect 2179 6117 2180 6151
rect 2144 6083 2180 6117
rect 2144 6049 2145 6083
rect 2179 6049 2180 6083
rect 2333 27695 2334 27729
rect 2368 27695 2369 27729
rect 2333 27661 2369 27695
rect 2333 27627 2334 27661
rect 2368 27627 2369 27661
rect 2333 27593 2369 27627
rect 2333 27559 2334 27593
rect 2368 27559 2369 27593
rect 2333 27525 2369 27559
rect 2333 27491 2334 27525
rect 2368 27491 2369 27525
rect 2333 27457 2369 27491
rect 2333 27423 2334 27457
rect 2368 27423 2369 27457
rect 2333 27389 2369 27423
rect 2333 27355 2334 27389
rect 2368 27355 2369 27389
rect 2333 27321 2369 27355
rect 2333 27287 2334 27321
rect 2368 27287 2369 27321
rect 2333 27253 2369 27287
rect 2333 27219 2334 27253
rect 2368 27219 2369 27253
rect 2333 27185 2369 27219
rect 2333 27151 2334 27185
rect 2368 27151 2369 27185
rect 2333 27117 2369 27151
rect 2333 27083 2334 27117
rect 2368 27083 2369 27117
rect 2333 27049 2369 27083
rect 2333 27015 2334 27049
rect 2368 27015 2369 27049
rect 2333 26981 2369 27015
rect 2333 26947 2334 26981
rect 2368 26947 2369 26981
rect 2333 26913 2369 26947
rect 2333 26879 2334 26913
rect 2368 26879 2369 26913
rect 2333 26845 2369 26879
rect 2333 26811 2334 26845
rect 2368 26811 2369 26845
rect 2333 26777 2369 26811
rect 2333 26743 2334 26777
rect 2368 26743 2369 26777
rect 2333 26709 2369 26743
rect 2333 26675 2334 26709
rect 2368 26675 2369 26709
rect 2333 26641 2369 26675
rect 2333 26607 2334 26641
rect 2368 26607 2369 26641
rect 2333 26573 2369 26607
rect 2333 26539 2334 26573
rect 2368 26539 2369 26573
rect 2333 26505 2369 26539
rect 2333 26471 2334 26505
rect 2368 26471 2369 26505
rect 2333 26437 2369 26471
rect 2333 26403 2334 26437
rect 2368 26403 2369 26437
rect 2333 26369 2369 26403
rect 2333 26335 2334 26369
rect 2368 26335 2369 26369
rect 2333 26301 2369 26335
rect 2333 26267 2334 26301
rect 2368 26267 2369 26301
rect 2333 26233 2369 26267
rect 2333 26199 2334 26233
rect 2368 26199 2369 26233
rect 2333 26165 2369 26199
rect 2333 26131 2334 26165
rect 2368 26131 2369 26165
rect 2333 26097 2369 26131
rect 2333 26063 2334 26097
rect 2368 26063 2369 26097
rect 2333 26029 2369 26063
rect 2333 25995 2334 26029
rect 2368 25995 2369 26029
rect 2333 25961 2369 25995
rect 2333 25927 2334 25961
rect 2368 25927 2369 25961
rect 2333 25893 2369 25927
rect 2333 25859 2334 25893
rect 2368 25859 2369 25893
rect 2333 25825 2369 25859
rect 2333 25791 2334 25825
rect 2368 25791 2369 25825
rect 2333 25757 2369 25791
rect 2333 25723 2334 25757
rect 2368 25723 2369 25757
rect 2333 25689 2369 25723
rect 2333 25655 2334 25689
rect 2368 25655 2369 25689
rect 2333 25621 2369 25655
rect 2333 25587 2334 25621
rect 2368 25587 2369 25621
rect 2333 25553 2369 25587
rect 2333 25519 2334 25553
rect 2368 25519 2369 25553
rect 2333 25485 2369 25519
rect 2333 25451 2334 25485
rect 2368 25451 2369 25485
rect 2333 25417 2369 25451
rect 2333 25383 2334 25417
rect 2368 25383 2369 25417
rect 2333 25349 2369 25383
rect 2333 25315 2334 25349
rect 2368 25315 2369 25349
rect 2333 25281 2369 25315
rect 2333 25247 2334 25281
rect 2368 25247 2369 25281
rect 2333 25213 2369 25247
rect 2333 25179 2334 25213
rect 2368 25179 2369 25213
rect 2333 25145 2369 25179
rect 2333 25111 2334 25145
rect 2368 25111 2369 25145
rect 2333 25077 2369 25111
rect 2333 25043 2334 25077
rect 2368 25043 2369 25077
rect 2333 25009 2369 25043
rect 2333 24975 2334 25009
rect 2368 24975 2369 25009
rect 2333 24941 2369 24975
rect 2333 24907 2334 24941
rect 2368 24907 2369 24941
rect 2333 24873 2369 24907
rect 2333 24839 2334 24873
rect 2368 24839 2369 24873
rect 2333 24805 2369 24839
rect 2333 24771 2334 24805
rect 2368 24771 2369 24805
rect 2333 24737 2369 24771
rect 2333 24703 2334 24737
rect 2368 24703 2369 24737
rect 2333 24669 2369 24703
rect 2333 24635 2334 24669
rect 2368 24635 2369 24669
rect 2333 24601 2369 24635
rect 2333 24567 2334 24601
rect 2368 24567 2369 24601
rect 2333 24533 2369 24567
rect 2333 24499 2334 24533
rect 2368 24499 2369 24533
rect 2333 24465 2369 24499
rect 2333 24431 2334 24465
rect 2368 24431 2369 24465
rect 2333 24397 2369 24431
rect 2333 24363 2334 24397
rect 2368 24363 2369 24397
rect 2333 24329 2369 24363
rect 2333 24295 2334 24329
rect 2368 24295 2369 24329
rect 2333 24261 2369 24295
rect 2333 24227 2334 24261
rect 2368 24227 2369 24261
rect 2333 24193 2369 24227
rect 2333 24159 2334 24193
rect 2368 24159 2369 24193
rect 2333 24125 2369 24159
rect 2333 24091 2334 24125
rect 2368 24091 2369 24125
rect 2333 24057 2369 24091
rect 2333 24023 2334 24057
rect 2368 24023 2369 24057
rect 2333 23989 2369 24023
rect 2333 23955 2334 23989
rect 2368 23955 2369 23989
rect 2333 23921 2369 23955
rect 2333 23887 2334 23921
rect 2368 23887 2369 23921
rect 2333 23853 2369 23887
rect 2333 23819 2334 23853
rect 2368 23819 2369 23853
rect 2333 23785 2369 23819
rect 2333 23751 2334 23785
rect 2368 23751 2369 23785
rect 2333 23717 2369 23751
rect 2333 23683 2334 23717
rect 2368 23683 2369 23717
rect 2333 23649 2369 23683
rect 2333 23615 2334 23649
rect 2368 23615 2369 23649
rect 2333 23581 2369 23615
rect 2333 23547 2334 23581
rect 2368 23547 2369 23581
rect 2333 23513 2369 23547
rect 2333 23479 2334 23513
rect 2368 23479 2369 23513
rect 2333 23445 2369 23479
rect 2333 23411 2334 23445
rect 2368 23411 2369 23445
rect 2333 23377 2369 23411
rect 2333 23343 2334 23377
rect 2368 23343 2369 23377
rect 2333 23309 2369 23343
rect 2333 23275 2334 23309
rect 2368 23275 2369 23309
rect 2333 23241 2369 23275
rect 2333 23207 2334 23241
rect 2368 23207 2369 23241
rect 2333 23173 2369 23207
rect 2333 23139 2334 23173
rect 2368 23139 2369 23173
rect 2333 23105 2369 23139
rect 2333 23071 2334 23105
rect 2368 23071 2369 23105
rect 2333 23037 2369 23071
rect 2333 23003 2334 23037
rect 2368 23003 2369 23037
rect 2333 22969 2369 23003
rect 2333 22935 2334 22969
rect 2368 22935 2369 22969
rect 2333 22901 2369 22935
rect 2333 22867 2334 22901
rect 2368 22867 2369 22901
rect 2333 22833 2369 22867
rect 2333 22799 2334 22833
rect 2368 22799 2369 22833
rect 2333 22765 2369 22799
rect 2333 22731 2334 22765
rect 2368 22731 2369 22765
rect 2333 22697 2369 22731
rect 2333 22663 2334 22697
rect 2368 22663 2369 22697
rect 2333 22629 2369 22663
rect 2333 22595 2334 22629
rect 2368 22595 2369 22629
rect 2333 22561 2369 22595
rect 2333 22527 2334 22561
rect 2368 22527 2369 22561
rect 2333 22493 2369 22527
rect 2333 22459 2334 22493
rect 2368 22459 2369 22493
rect 2333 22425 2369 22459
rect 2333 22391 2334 22425
rect 2368 22391 2369 22425
rect 2333 22357 2369 22391
rect 2333 22323 2334 22357
rect 2368 22323 2369 22357
rect 2333 22289 2369 22323
rect 2333 22255 2334 22289
rect 2368 22255 2369 22289
rect 2333 22221 2369 22255
rect 2333 22187 2334 22221
rect 2368 22187 2369 22221
rect 2333 22153 2369 22187
rect 2333 22119 2334 22153
rect 2368 22119 2369 22153
rect 2333 22085 2369 22119
rect 2333 22051 2334 22085
rect 2368 22051 2369 22085
rect 2333 22017 2369 22051
rect 2333 21983 2334 22017
rect 2368 21983 2369 22017
rect 2333 21949 2369 21983
rect 2333 21915 2334 21949
rect 2368 21915 2369 21949
rect 2333 21881 2369 21915
rect 2333 21847 2334 21881
rect 2368 21847 2369 21881
rect 2333 21813 2369 21847
rect 2333 21779 2334 21813
rect 2368 21779 2369 21813
rect 2333 21745 2369 21779
rect 2333 21711 2334 21745
rect 2368 21711 2369 21745
rect 2333 21677 2369 21711
rect 2333 21643 2334 21677
rect 2368 21643 2369 21677
rect 2333 21609 2369 21643
rect 2333 21575 2334 21609
rect 2368 21575 2369 21609
rect 2333 21541 2369 21575
rect 2333 21507 2334 21541
rect 2368 21507 2369 21541
rect 2333 21473 2369 21507
rect 2333 21439 2334 21473
rect 2368 21439 2369 21473
rect 2333 21405 2369 21439
rect 2333 21371 2334 21405
rect 2368 21371 2369 21405
rect 2333 21337 2369 21371
rect 2333 21303 2334 21337
rect 2368 21303 2369 21337
rect 2333 21269 2369 21303
rect 2333 21235 2334 21269
rect 2368 21235 2369 21269
rect 2333 21201 2369 21235
rect 2333 21167 2334 21201
rect 2368 21167 2369 21201
rect 2333 21133 2369 21167
rect 2333 21099 2334 21133
rect 2368 21099 2369 21133
rect 2333 21065 2369 21099
rect 2333 21031 2334 21065
rect 2368 21031 2369 21065
rect 2333 20997 2369 21031
rect 2333 20963 2334 20997
rect 2368 20963 2369 20997
rect 2333 20929 2369 20963
rect 2333 20895 2334 20929
rect 2368 20895 2369 20929
rect 2333 20861 2369 20895
rect 2333 20827 2334 20861
rect 2368 20827 2369 20861
rect 2333 20793 2369 20827
rect 2333 20759 2334 20793
rect 2368 20759 2369 20793
rect 2333 20725 2369 20759
rect 2333 20691 2334 20725
rect 2368 20691 2369 20725
rect 2333 20657 2369 20691
rect 2333 20623 2334 20657
rect 2368 20623 2369 20657
rect 2333 20589 2369 20623
rect 2333 20555 2334 20589
rect 2368 20555 2369 20589
rect 2333 20521 2369 20555
rect 2333 20487 2334 20521
rect 2368 20487 2369 20521
rect 2333 20453 2369 20487
rect 2333 20419 2334 20453
rect 2368 20419 2369 20453
rect 2333 20385 2369 20419
rect 2333 20351 2334 20385
rect 2368 20351 2369 20385
rect 2333 20317 2369 20351
rect 2333 20283 2334 20317
rect 2368 20283 2369 20317
rect 2333 20249 2369 20283
rect 2333 20215 2334 20249
rect 2368 20215 2369 20249
rect 2333 20181 2369 20215
rect 2333 20147 2334 20181
rect 2368 20147 2369 20181
rect 2333 20113 2369 20147
rect 2333 20079 2334 20113
rect 2368 20079 2369 20113
rect 2333 20045 2369 20079
rect 2333 20011 2334 20045
rect 2368 20011 2369 20045
rect 2333 19977 2369 20011
rect 2333 19943 2334 19977
rect 2368 19943 2369 19977
rect 2333 19909 2369 19943
rect 2333 19875 2334 19909
rect 2368 19875 2369 19909
rect 2333 19841 2369 19875
rect 2333 19807 2334 19841
rect 2368 19807 2369 19841
rect 2333 19773 2369 19807
rect 2333 19739 2334 19773
rect 2368 19739 2369 19773
rect 2333 19705 2369 19739
rect 2333 19671 2334 19705
rect 2368 19671 2369 19705
rect 2333 19637 2369 19671
rect 2333 19603 2334 19637
rect 2368 19603 2369 19637
rect 2333 19569 2369 19603
rect 2333 19535 2334 19569
rect 2368 19535 2369 19569
rect 2333 19501 2369 19535
rect 2333 19467 2334 19501
rect 2368 19467 2369 19501
rect 2333 19433 2369 19467
rect 2333 19399 2334 19433
rect 2368 19399 2369 19433
rect 2333 19365 2369 19399
rect 2333 19331 2334 19365
rect 2368 19331 2369 19365
rect 2333 19297 2369 19331
rect 2333 19263 2334 19297
rect 2368 19263 2369 19297
rect 2333 19229 2369 19263
rect 2333 19195 2334 19229
rect 2368 19195 2369 19229
rect 2333 19161 2369 19195
rect 2333 19127 2334 19161
rect 2368 19127 2369 19161
rect 2333 19093 2369 19127
rect 2333 19059 2334 19093
rect 2368 19059 2369 19093
rect 2333 19025 2369 19059
rect 2333 18991 2334 19025
rect 2368 18991 2369 19025
rect 2333 18957 2369 18991
rect 2333 18923 2334 18957
rect 2368 18923 2369 18957
rect 2333 18889 2369 18923
rect 2333 18855 2334 18889
rect 2368 18855 2369 18889
rect 2333 18821 2369 18855
rect 2333 18787 2334 18821
rect 2368 18787 2369 18821
rect 2333 18753 2369 18787
rect 2333 18719 2334 18753
rect 2368 18719 2369 18753
rect 2333 18685 2369 18719
rect 2333 18651 2334 18685
rect 2368 18651 2369 18685
rect 2333 18617 2369 18651
rect 2333 18583 2334 18617
rect 2368 18583 2369 18617
rect 2333 18549 2369 18583
rect 2333 18515 2334 18549
rect 2368 18515 2369 18549
rect 2333 18481 2369 18515
rect 2333 18447 2334 18481
rect 2368 18447 2369 18481
rect 2333 18413 2369 18447
rect 2333 18379 2334 18413
rect 2368 18379 2369 18413
rect 2333 18345 2369 18379
rect 2333 18311 2334 18345
rect 2368 18311 2369 18345
rect 2333 18277 2369 18311
rect 2333 18243 2334 18277
rect 2368 18243 2369 18277
rect 2333 18209 2369 18243
rect 2333 18175 2334 18209
rect 2368 18175 2369 18209
rect 2333 18141 2369 18175
rect 2333 18107 2334 18141
rect 2368 18107 2369 18141
rect 2333 18073 2369 18107
rect 2333 18039 2334 18073
rect 2368 18039 2369 18073
rect 2333 18005 2369 18039
rect 2333 17971 2334 18005
rect 2368 17971 2369 18005
rect 2333 17937 2369 17971
rect 2333 17903 2334 17937
rect 2368 17903 2369 17937
rect 2333 17869 2369 17903
rect 2333 17835 2334 17869
rect 2368 17835 2369 17869
rect 2333 17801 2369 17835
rect 2333 17767 2334 17801
rect 2368 17767 2369 17801
rect 2333 17733 2369 17767
rect 2333 17699 2334 17733
rect 2368 17699 2369 17733
rect 2333 17665 2369 17699
rect 2333 17631 2334 17665
rect 2368 17631 2369 17665
rect 2333 17597 2369 17631
rect 2333 17563 2334 17597
rect 2368 17563 2369 17597
rect 2333 17529 2369 17563
rect 2333 17495 2334 17529
rect 2368 17495 2369 17529
rect 2333 17461 2369 17495
rect 2333 17427 2334 17461
rect 2368 17427 2369 17461
rect 2333 17393 2369 17427
rect 2333 17359 2334 17393
rect 2368 17359 2369 17393
rect 2333 17325 2369 17359
rect 2333 17291 2334 17325
rect 2368 17291 2369 17325
rect 2333 17257 2369 17291
rect 2333 17223 2334 17257
rect 2368 17223 2369 17257
rect 2333 17189 2369 17223
rect 2333 17155 2334 17189
rect 2368 17155 2369 17189
rect 2333 17121 2369 17155
rect 2333 17087 2334 17121
rect 2368 17087 2369 17121
rect 2333 17053 2369 17087
rect 2333 17019 2334 17053
rect 2368 17019 2369 17053
rect 2333 16985 2369 17019
rect 2333 16951 2334 16985
rect 2368 16951 2369 16985
rect 2333 16917 2369 16951
rect 2333 16883 2334 16917
rect 2368 16883 2369 16917
rect 2333 16849 2369 16883
rect 2333 16815 2334 16849
rect 2368 16815 2369 16849
rect 2333 16781 2369 16815
rect 2333 16747 2334 16781
rect 2368 16747 2369 16781
rect 2333 16713 2369 16747
rect 2333 16679 2334 16713
rect 2368 16679 2369 16713
rect 2333 16645 2369 16679
rect 2333 16611 2334 16645
rect 2368 16611 2369 16645
rect 2333 16577 2369 16611
rect 2333 16543 2334 16577
rect 2368 16543 2369 16577
rect 2333 16509 2369 16543
rect 2333 16475 2334 16509
rect 2368 16475 2369 16509
rect 2333 16441 2369 16475
rect 2333 16407 2334 16441
rect 2368 16407 2369 16441
rect 2333 16373 2369 16407
rect 2333 16339 2334 16373
rect 2368 16339 2369 16373
rect 2333 16305 2369 16339
rect 2333 16271 2334 16305
rect 2368 16271 2369 16305
rect 2333 16237 2369 16271
rect 2333 16203 2334 16237
rect 2368 16203 2369 16237
rect 2333 16169 2369 16203
rect 2333 16135 2334 16169
rect 2368 16135 2369 16169
rect 2333 16101 2369 16135
rect 2333 16067 2334 16101
rect 2368 16067 2369 16101
rect 2333 16033 2369 16067
rect 2333 15999 2334 16033
rect 2368 15999 2369 16033
rect 2333 15965 2369 15999
rect 2333 15931 2334 15965
rect 2368 15931 2369 15965
rect 2333 15897 2369 15931
rect 2333 15863 2334 15897
rect 2368 15863 2369 15897
rect 2333 15829 2369 15863
rect 2333 15795 2334 15829
rect 2368 15795 2369 15829
rect 2333 15761 2369 15795
rect 2333 15727 2334 15761
rect 2368 15727 2369 15761
rect 2333 15693 2369 15727
rect 2333 15659 2334 15693
rect 2368 15659 2369 15693
rect 2333 15625 2369 15659
rect 2333 15591 2334 15625
rect 2368 15591 2369 15625
rect 2333 15557 2369 15591
rect 2333 15523 2334 15557
rect 2368 15523 2369 15557
rect 2333 15489 2369 15523
rect 2333 15455 2334 15489
rect 2368 15455 2369 15489
rect 2333 15421 2369 15455
rect 2333 15387 2334 15421
rect 2368 15387 2369 15421
rect 2333 15353 2369 15387
rect 2333 15319 2334 15353
rect 2368 15319 2369 15353
rect 2333 15285 2369 15319
rect 2333 15251 2334 15285
rect 2368 15251 2369 15285
rect 2333 15217 2369 15251
rect 2333 15183 2334 15217
rect 2368 15183 2369 15217
rect 2333 15149 2369 15183
rect 2333 15115 2334 15149
rect 2368 15115 2369 15149
rect 2333 15081 2369 15115
rect 2333 15047 2334 15081
rect 2368 15047 2369 15081
rect 2333 15013 2369 15047
rect 2333 14979 2334 15013
rect 2368 14979 2369 15013
rect 2333 14945 2369 14979
rect 2333 14911 2334 14945
rect 2368 14911 2369 14945
rect 2333 14877 2369 14911
rect 2333 14843 2334 14877
rect 2368 14843 2369 14877
rect 2333 14809 2369 14843
rect 2333 14775 2334 14809
rect 2368 14775 2369 14809
rect 2333 14741 2369 14775
rect 2333 14707 2334 14741
rect 2368 14707 2369 14741
rect 2333 14673 2369 14707
rect 2333 14639 2334 14673
rect 2368 14639 2369 14673
rect 2333 14605 2369 14639
rect 2333 14571 2334 14605
rect 2368 14571 2369 14605
rect 2333 14537 2369 14571
rect 2333 14503 2334 14537
rect 2368 14503 2369 14537
rect 2333 14469 2369 14503
rect 2333 14435 2334 14469
rect 2368 14435 2369 14469
rect 2333 14401 2369 14435
rect 2333 14367 2334 14401
rect 2368 14367 2369 14401
rect 2333 14333 2369 14367
rect 2333 14299 2334 14333
rect 2368 14299 2369 14333
rect 2333 14265 2369 14299
rect 2333 14231 2334 14265
rect 2368 14231 2369 14265
rect 2333 14197 2369 14231
rect 2333 14163 2334 14197
rect 2368 14163 2369 14197
rect 2333 14129 2369 14163
rect 2333 14095 2334 14129
rect 2368 14095 2369 14129
rect 2333 14061 2369 14095
rect 2333 14027 2334 14061
rect 2368 14027 2369 14061
rect 2333 13993 2369 14027
rect 2333 13959 2334 13993
rect 2368 13959 2369 13993
rect 2333 13925 2369 13959
rect 2333 13891 2334 13925
rect 2368 13891 2369 13925
rect 2333 13857 2369 13891
rect 2333 13823 2334 13857
rect 2368 13823 2369 13857
rect 2333 13789 2369 13823
rect 2333 13755 2334 13789
rect 2368 13755 2369 13789
rect 2333 13721 2369 13755
rect 2333 13687 2334 13721
rect 2368 13687 2369 13721
rect 2333 13653 2369 13687
rect 2333 13619 2334 13653
rect 2368 13619 2369 13653
rect 2333 13585 2369 13619
rect 2333 13551 2334 13585
rect 2368 13551 2369 13585
rect 2333 13517 2369 13551
rect 2333 13483 2334 13517
rect 2368 13483 2369 13517
rect 2333 13449 2369 13483
rect 2333 13415 2334 13449
rect 2368 13415 2369 13449
rect 2333 13381 2369 13415
rect 2333 13347 2334 13381
rect 2368 13347 2369 13381
rect 2333 13313 2369 13347
rect 2333 13279 2334 13313
rect 2368 13279 2369 13313
rect 2333 13245 2369 13279
rect 2333 13211 2334 13245
rect 2368 13211 2369 13245
rect 2333 13177 2369 13211
rect 2333 13143 2334 13177
rect 2368 13143 2369 13177
rect 2333 13109 2369 13143
rect 2333 13075 2334 13109
rect 2368 13075 2369 13109
rect 2333 13041 2369 13075
rect 2333 13007 2334 13041
rect 2368 13007 2369 13041
rect 2333 12973 2369 13007
rect 2333 12939 2334 12973
rect 2368 12939 2369 12973
rect 2333 12905 2369 12939
rect 2333 12871 2334 12905
rect 2368 12871 2369 12905
rect 2333 12837 2369 12871
rect 2333 12803 2334 12837
rect 2368 12803 2369 12837
rect 2333 12769 2369 12803
rect 2333 12735 2334 12769
rect 2368 12735 2369 12769
rect 2333 12701 2369 12735
rect 2333 12667 2334 12701
rect 2368 12667 2369 12701
rect 2333 12633 2369 12667
rect 2333 12599 2334 12633
rect 2368 12599 2369 12633
rect 2333 12565 2369 12599
rect 2333 12531 2334 12565
rect 2368 12531 2369 12565
rect 2333 12497 2369 12531
rect 2333 12463 2334 12497
rect 2368 12463 2369 12497
rect 2333 12429 2369 12463
rect 2333 12395 2334 12429
rect 2368 12395 2369 12429
rect 2333 12361 2369 12395
rect 2333 12327 2334 12361
rect 2368 12327 2369 12361
rect 2333 12293 2369 12327
rect 2333 12259 2334 12293
rect 2368 12259 2369 12293
rect 2333 12225 2369 12259
rect 2333 12191 2334 12225
rect 2368 12191 2369 12225
rect 2333 12157 2369 12191
rect 2333 12123 2334 12157
rect 2368 12123 2369 12157
rect 2333 12089 2369 12123
rect 2333 12055 2334 12089
rect 2368 12055 2369 12089
rect 2333 12021 2369 12055
rect 2333 11987 2334 12021
rect 2368 11987 2369 12021
rect 2333 11953 2369 11987
rect 2333 11919 2334 11953
rect 2368 11919 2369 11953
rect 2333 11885 2369 11919
rect 2333 11851 2334 11885
rect 2368 11851 2369 11885
rect 2333 11817 2369 11851
rect 2333 11783 2334 11817
rect 2368 11783 2369 11817
rect 2333 11749 2369 11783
rect 2333 11715 2334 11749
rect 2368 11715 2369 11749
rect 2333 11681 2369 11715
rect 2333 11647 2334 11681
rect 2368 11647 2369 11681
rect 2333 11613 2369 11647
rect 2333 11579 2334 11613
rect 2368 11579 2369 11613
rect 2333 11545 2369 11579
rect 2333 11511 2334 11545
rect 2368 11511 2369 11545
rect 2333 11477 2369 11511
rect 2333 11443 2334 11477
rect 2368 11443 2369 11477
rect 2333 11409 2369 11443
rect 2333 11375 2334 11409
rect 2368 11375 2369 11409
rect 2333 11341 2369 11375
rect 2333 11307 2334 11341
rect 2368 11307 2369 11341
rect 2333 11273 2369 11307
rect 2333 11239 2334 11273
rect 2368 11239 2369 11273
rect 2333 11205 2369 11239
rect 2333 11171 2334 11205
rect 2368 11171 2369 11205
rect 2333 11137 2369 11171
rect 2333 11103 2334 11137
rect 2368 11103 2369 11137
rect 2333 11069 2369 11103
rect 2333 11035 2334 11069
rect 2368 11035 2369 11069
rect 2333 11001 2369 11035
rect 2333 10967 2334 11001
rect 2368 10967 2369 11001
rect 2333 10933 2369 10967
rect 2333 10899 2334 10933
rect 2368 10899 2369 10933
rect 2333 10865 2369 10899
rect 2333 10831 2334 10865
rect 2368 10831 2369 10865
rect 2333 10797 2369 10831
rect 2333 10763 2334 10797
rect 2368 10763 2369 10797
rect 2333 10729 2369 10763
rect 2333 10695 2334 10729
rect 2368 10695 2369 10729
rect 2333 10661 2369 10695
rect 2333 10627 2334 10661
rect 2368 10627 2369 10661
rect 2333 10593 2369 10627
rect 2333 10559 2334 10593
rect 2368 10559 2369 10593
rect 2333 10525 2369 10559
rect 2333 10491 2334 10525
rect 2368 10491 2369 10525
rect 2333 10457 2369 10491
rect 2333 10423 2334 10457
rect 2368 10423 2369 10457
rect 2333 10389 2369 10423
rect 2333 10355 2334 10389
rect 2368 10355 2369 10389
rect 2333 10321 2369 10355
rect 2333 10287 2334 10321
rect 2368 10287 2369 10321
rect 2333 10253 2369 10287
rect 2333 10219 2334 10253
rect 2368 10219 2369 10253
rect 2333 10185 2369 10219
rect 2333 10151 2334 10185
rect 2368 10151 2369 10185
rect 2333 10117 2369 10151
rect 2333 10083 2334 10117
rect 2368 10083 2369 10117
rect 2333 10049 2369 10083
rect 2333 10015 2334 10049
rect 2368 10015 2369 10049
rect 2333 9981 2369 10015
rect 2333 9947 2334 9981
rect 2368 9947 2369 9981
rect 2333 9913 2369 9947
rect 2333 9879 2334 9913
rect 2368 9879 2369 9913
rect 2333 9845 2369 9879
rect 2333 9811 2334 9845
rect 2368 9811 2369 9845
rect 2333 9777 2369 9811
rect 2333 9743 2334 9777
rect 2368 9743 2369 9777
rect 2333 9709 2369 9743
rect 2333 9675 2334 9709
rect 2368 9675 2369 9709
rect 2333 9641 2369 9675
rect 2333 9607 2334 9641
rect 2368 9607 2369 9641
rect 2333 9573 2369 9607
rect 2333 9539 2334 9573
rect 2368 9539 2369 9573
rect 2333 9505 2369 9539
rect 2333 9471 2334 9505
rect 2368 9471 2369 9505
rect 2333 9437 2369 9471
rect 2333 9403 2334 9437
rect 2368 9403 2369 9437
rect 2333 9369 2369 9403
rect 2333 9335 2334 9369
rect 2368 9335 2369 9369
rect 2333 9301 2369 9335
rect 2333 9267 2334 9301
rect 2368 9267 2369 9301
rect 2333 9233 2369 9267
rect 2333 9199 2334 9233
rect 2368 9199 2369 9233
rect 2333 9165 2369 9199
rect 2333 9131 2334 9165
rect 2368 9131 2369 9165
rect 2333 9097 2369 9131
rect 2333 9063 2334 9097
rect 2368 9063 2369 9097
rect 2333 9029 2369 9063
rect 2333 8995 2334 9029
rect 2368 8995 2369 9029
rect 2333 8961 2369 8995
rect 2333 8927 2334 8961
rect 2368 8927 2369 8961
rect 2333 8893 2369 8927
rect 2333 8859 2334 8893
rect 2368 8859 2369 8893
rect 2333 8825 2369 8859
rect 2333 8791 2334 8825
rect 2368 8791 2369 8825
rect 2333 8757 2369 8791
rect 2333 8723 2334 8757
rect 2368 8723 2369 8757
rect 2333 8689 2369 8723
rect 2333 8655 2334 8689
rect 2368 8655 2369 8689
rect 2333 8621 2369 8655
rect 2333 8587 2334 8621
rect 2368 8587 2369 8621
rect 2333 8553 2369 8587
rect 2333 8519 2334 8553
rect 2368 8519 2369 8553
rect 2333 8485 2369 8519
rect 2333 8451 2334 8485
rect 2368 8451 2369 8485
rect 2333 8417 2369 8451
rect 2333 8383 2334 8417
rect 2368 8383 2369 8417
rect 2333 8349 2369 8383
rect 2333 8315 2334 8349
rect 2368 8315 2369 8349
rect 2333 8281 2369 8315
rect 2333 8247 2334 8281
rect 2368 8247 2369 8281
rect 2333 8213 2369 8247
rect 2333 8179 2334 8213
rect 2368 8179 2369 8213
rect 2333 8145 2369 8179
rect 2333 8111 2334 8145
rect 2368 8111 2369 8145
rect 2333 8077 2369 8111
rect 2333 8043 2334 8077
rect 2368 8043 2369 8077
rect 2333 8009 2369 8043
rect 2333 7975 2334 8009
rect 2368 7975 2369 8009
rect 2333 7941 2369 7975
rect 2333 7907 2334 7941
rect 2368 7907 2369 7941
rect 2333 7873 2369 7907
rect 2333 7839 2334 7873
rect 2368 7839 2369 7873
rect 2333 7805 2369 7839
rect 2333 7771 2334 7805
rect 2368 7771 2369 7805
rect 2333 7737 2369 7771
rect 2333 7703 2334 7737
rect 2368 7703 2369 7737
rect 2333 7669 2369 7703
rect 2333 7635 2334 7669
rect 2368 7635 2369 7669
rect 2333 7601 2369 7635
rect 2333 7567 2334 7601
rect 2368 7567 2369 7601
rect 2333 7533 2369 7567
rect 2333 7499 2334 7533
rect 2368 7499 2369 7533
rect 2333 7465 2369 7499
rect 2333 7431 2334 7465
rect 2368 7431 2369 7465
rect 2333 7397 2369 7431
rect 2333 7363 2334 7397
rect 2368 7363 2369 7397
rect 2333 7329 2369 7363
rect 2333 7295 2334 7329
rect 2368 7295 2369 7329
rect 2333 7261 2369 7295
rect 2333 7227 2334 7261
rect 2368 7227 2369 7261
rect 2333 7193 2369 7227
rect 2333 7159 2334 7193
rect 2368 7159 2369 7193
rect 2333 7125 2369 7159
rect 2333 7091 2334 7125
rect 2368 7091 2369 7125
rect 2333 7057 2369 7091
rect 2333 7023 2334 7057
rect 2368 7023 2369 7057
rect 2333 6989 2369 7023
rect 2333 6955 2334 6989
rect 2368 6955 2369 6989
rect 2333 6921 2369 6955
rect 2333 6887 2334 6921
rect 2368 6887 2369 6921
rect 2333 6853 2369 6887
rect 2333 6819 2334 6853
rect 2368 6819 2369 6853
rect 2333 6785 2369 6819
rect 2333 6751 2334 6785
rect 2368 6751 2369 6785
rect 2333 6717 2369 6751
rect 2333 6683 2334 6717
rect 2368 6683 2369 6717
rect 2333 6649 2369 6683
rect 2333 6615 2334 6649
rect 2368 6615 2369 6649
rect 2333 6581 2369 6615
rect 2333 6547 2334 6581
rect 2368 6547 2369 6581
rect 2333 6513 2369 6547
rect 2333 6479 2334 6513
rect 2368 6479 2369 6513
rect 2333 6445 2369 6479
rect 2333 6411 2334 6445
rect 2368 6411 2369 6445
rect 2333 6377 2369 6411
rect 2333 6343 2334 6377
rect 2368 6343 2369 6377
rect 2333 6309 2369 6343
rect 2333 6275 2334 6309
rect 2368 6275 2369 6309
rect 2333 6264 2369 6275
rect 2333 6207 2334 6264
rect 2368 6207 2369 6264
rect 2553 11009 2589 11043
rect 2553 10975 2554 11009
rect 2588 10975 2589 11009
rect 2553 10941 2589 10975
rect 2553 10907 2554 10941
rect 2588 10907 2589 10941
rect 2553 10873 2589 10907
rect 6853 10995 6889 11043
rect 6853 10961 6854 10995
rect 6888 10961 6889 10995
rect 6853 10927 6889 10961
rect 6853 10893 6854 10927
rect 6888 10893 6889 10927
rect 2553 10839 2554 10873
rect 2588 10839 2589 10873
rect 2553 10805 2589 10839
rect 2553 10771 2554 10805
rect 2588 10771 2589 10805
rect 2553 10737 2589 10771
rect 2553 10703 2554 10737
rect 2588 10703 2589 10737
rect 2553 10669 2589 10703
rect 2553 10635 2554 10669
rect 2588 10635 2589 10669
rect 2553 10601 2589 10635
rect 2553 10567 2554 10601
rect 2588 10567 2589 10601
rect 2553 10533 2589 10567
rect 2553 10499 2554 10533
rect 2588 10499 2589 10533
rect 2553 10465 2589 10499
rect 2553 10431 2554 10465
rect 2588 10431 2589 10465
rect 2553 10397 2589 10431
rect 2553 10363 2554 10397
rect 2588 10363 2589 10397
rect 2553 10329 2589 10363
rect 2553 10295 2554 10329
rect 2588 10295 2589 10329
rect 2553 10261 2589 10295
rect 2553 10227 2554 10261
rect 2588 10227 2589 10261
rect 2553 10193 2589 10227
rect 2553 10159 2554 10193
rect 2588 10159 2589 10193
rect 2553 10125 2589 10159
rect 2553 10091 2554 10125
rect 2588 10091 2589 10125
rect 2553 10057 2589 10091
rect 2553 10023 2554 10057
rect 2588 10023 2589 10057
rect 2553 9989 2589 10023
rect 2553 9955 2554 9989
rect 2588 9955 2589 9989
rect 2553 9921 2589 9955
rect 2553 9887 2554 9921
rect 2588 9887 2589 9921
rect 2553 9853 2589 9887
rect 2553 9819 2554 9853
rect 2588 9819 2589 9853
rect 2553 9785 2589 9819
rect 2553 9751 2554 9785
rect 2588 9751 2589 9785
rect 2553 9717 2589 9751
rect 2553 9683 2554 9717
rect 2588 9683 2589 9717
rect 2553 9649 2589 9683
rect 2553 9615 2554 9649
rect 2588 9615 2589 9649
rect 2553 9581 2589 9615
rect 2553 9547 2554 9581
rect 2588 9547 2589 9581
rect 2553 9513 2589 9547
rect 2553 9479 2554 9513
rect 2588 9479 2589 9513
rect 2553 9445 2589 9479
rect 2553 9411 2554 9445
rect 2588 9411 2589 9445
rect 2553 9377 2589 9411
rect 2553 9343 2554 9377
rect 2588 9343 2589 9377
rect 2553 9309 2589 9343
rect 2553 9275 2554 9309
rect 2588 9275 2589 9309
rect 2553 9241 2589 9275
rect 2553 9207 2554 9241
rect 2588 9207 2589 9241
rect 2553 9173 2589 9207
rect 2553 9139 2554 9173
rect 2588 9139 2589 9173
rect 2553 9105 2589 9139
rect 2553 9071 2554 9105
rect 2588 9071 2589 9105
rect 2553 9037 2589 9071
rect 2553 9003 2554 9037
rect 2588 9003 2589 9037
rect 2553 8969 2589 9003
rect 2553 8935 2554 8969
rect 2588 8935 2589 8969
rect 2553 8901 2589 8935
rect 2553 8867 2554 8901
rect 2588 8867 2589 8901
rect 2553 8833 2589 8867
rect 2553 8799 2554 8833
rect 2588 8799 2589 8833
rect 2553 8765 2589 8799
rect 2553 8731 2554 8765
rect 2588 8731 2589 8765
rect 2553 8697 2589 8731
rect 2553 8663 2554 8697
rect 2588 8663 2589 8697
rect 2553 8629 2589 8663
rect 2553 8595 2554 8629
rect 2588 8595 2589 8629
rect 2553 8561 2589 8595
rect 2553 8527 2554 8561
rect 2588 8527 2589 8561
rect 2553 8493 2589 8527
rect 2553 8459 2554 8493
rect 2588 8459 2589 8493
rect 2553 8425 2589 8459
rect 2553 8391 2554 8425
rect 2588 8391 2589 8425
rect 2553 8357 2589 8391
rect 2553 8323 2554 8357
rect 2588 8323 2589 8357
rect 2553 8289 2589 8323
rect 2553 8255 2554 8289
rect 2588 8255 2589 8289
rect 2553 8221 2589 8255
rect 2553 8187 2554 8221
rect 2588 8187 2589 8221
rect 2553 8153 2589 8187
rect 2553 8119 2554 8153
rect 2588 8119 2589 8153
rect 2553 8085 2589 8119
rect 2553 8051 2554 8085
rect 2588 8051 2589 8085
rect 2553 8017 2589 8051
rect 2553 7983 2554 8017
rect 2588 7983 2589 8017
rect 2553 7949 2589 7983
rect 2553 7915 2554 7949
rect 2588 7915 2589 7949
rect 2553 7881 2589 7915
rect 2553 7847 2554 7881
rect 2588 7847 2589 7881
rect 2553 7813 2589 7847
rect 2553 7779 2554 7813
rect 2588 7779 2589 7813
rect 2553 7745 2589 7779
rect 2553 7711 2554 7745
rect 2588 7711 2589 7745
rect 2553 7677 2589 7711
rect 2553 7643 2554 7677
rect 2588 7643 2589 7677
rect 2553 7609 2589 7643
rect 2553 7575 2554 7609
rect 2588 7575 2589 7609
rect 2553 7541 2589 7575
rect 2553 7507 2554 7541
rect 2588 7507 2589 7541
rect 2553 7473 2589 7507
rect 2553 7439 2554 7473
rect 2588 7439 2589 7473
rect 2553 7405 2589 7439
rect 2553 7371 2554 7405
rect 2588 7371 2589 7405
rect 2553 7337 2589 7371
rect 2553 7303 2554 7337
rect 2588 7303 2589 7337
rect 2553 7269 2589 7303
rect 2553 7235 2554 7269
rect 2588 7235 2589 7269
rect 2553 7201 2589 7235
rect 2553 7167 2554 7201
rect 2588 7167 2589 7201
rect 2553 7133 2589 7167
rect 2553 7099 2554 7133
rect 2588 7099 2589 7133
rect 2553 7065 2589 7099
rect 2553 7031 2554 7065
rect 2588 7031 2589 7065
rect 2553 6997 2589 7031
rect 2553 6963 2554 6997
rect 2588 6963 2589 6997
rect 2553 6929 2589 6963
rect 2553 6895 2554 6929
rect 2588 6895 2589 6929
rect 2553 6861 2589 6895
rect 2553 6827 2554 6861
rect 2588 6827 2589 6861
rect 2553 6793 2589 6827
rect 2553 6759 2554 6793
rect 2588 6759 2589 6793
rect 2553 6725 2589 6759
rect 2553 6691 2554 6725
rect 2588 6691 2589 6725
rect 2553 6657 2589 6691
rect 2553 6623 2554 6657
rect 2588 6623 2589 6657
rect 2553 6589 2589 6623
rect 2553 6555 2554 6589
rect 2588 6555 2589 6589
rect 2553 6521 2589 6555
rect 2553 6487 2554 6521
rect 2588 6487 2589 6521
rect 2553 6453 2589 6487
rect 2553 6419 2554 6453
rect 2588 6419 2589 6453
rect 2742 10889 6700 10890
rect 2742 10856 2835 10889
rect 2742 10822 2743 10856
rect 2777 10855 2835 10856
rect 2869 10855 2903 10889
rect 2937 10855 2971 10889
rect 3005 10855 3039 10889
rect 3073 10855 3107 10889
rect 3141 10855 3175 10889
rect 3209 10855 3243 10889
rect 3277 10855 3311 10889
rect 3345 10855 3379 10889
rect 3413 10855 3447 10889
rect 3481 10855 3515 10889
rect 3549 10855 3583 10889
rect 3617 10855 3651 10889
rect 3685 10855 3719 10889
rect 3753 10855 3787 10889
rect 3821 10855 3855 10889
rect 3889 10855 3923 10889
rect 3957 10855 3991 10889
rect 4025 10855 4059 10889
rect 4093 10855 4127 10889
rect 4161 10855 4195 10889
rect 4229 10855 4263 10889
rect 4297 10855 4331 10889
rect 4365 10855 4399 10889
rect 4433 10855 4467 10889
rect 4501 10855 4535 10889
rect 4569 10855 4603 10889
rect 4637 10855 4671 10889
rect 4705 10855 4799 10889
rect 4833 10855 4867 10889
rect 4901 10855 4935 10889
rect 4969 10855 5003 10889
rect 5037 10855 5071 10889
rect 5105 10855 5139 10889
rect 5173 10855 5207 10889
rect 5241 10855 5275 10889
rect 5309 10855 5343 10889
rect 5377 10855 5411 10889
rect 5445 10855 5479 10889
rect 5513 10855 5547 10889
rect 5581 10855 5615 10889
rect 5649 10855 5683 10889
rect 5717 10855 5751 10889
rect 5785 10855 5819 10889
rect 5853 10855 5887 10889
rect 5921 10855 5955 10889
rect 5989 10855 6023 10889
rect 6057 10855 6091 10889
rect 6125 10855 6159 10889
rect 6193 10855 6227 10889
rect 6261 10855 6295 10889
rect 6329 10855 6363 10889
rect 6397 10855 6431 10889
rect 6465 10855 6499 10889
rect 6533 10855 6567 10889
rect 6601 10856 6700 10889
rect 6601 10855 6665 10856
rect 2777 10854 6665 10855
rect 2777 10822 2778 10854
rect 2742 10788 2778 10822
rect 2742 10754 2743 10788
rect 2777 10754 2778 10788
rect 2742 10720 2778 10754
rect 2932 10723 4534 10804
rect 4703 10776 4739 10854
rect 6664 10822 6665 10854
rect 6699 10822 6700 10856
rect 4703 10742 4704 10776
rect 4738 10742 4739 10776
rect 2742 10686 2743 10720
rect 2777 10686 2778 10720
rect 2742 10652 2778 10686
rect 2742 10618 2743 10652
rect 2777 10618 2778 10652
rect 2742 10584 2778 10618
rect 2742 10550 2743 10584
rect 2777 10550 2778 10584
rect 2742 10516 2778 10550
rect 2742 10482 2743 10516
rect 2777 10482 2778 10516
rect 2742 10448 2778 10482
rect 2742 10414 2743 10448
rect 2777 10414 2778 10448
rect 2742 10380 2778 10414
rect 2742 10346 2743 10380
rect 2777 10346 2778 10380
rect 2742 10312 2778 10346
rect 2742 10278 2743 10312
rect 2777 10278 2778 10312
rect 2742 10244 2778 10278
rect 2742 10210 2743 10244
rect 2777 10210 2778 10244
rect 2742 10176 2778 10210
rect 2742 10142 2743 10176
rect 2777 10142 2778 10176
rect 2742 10108 2778 10142
rect 2742 10074 2743 10108
rect 2777 10074 2778 10108
rect 2742 10040 2778 10074
rect 2742 10006 2743 10040
rect 2777 10006 2778 10040
rect 2742 9972 2778 10006
rect 2742 9938 2743 9972
rect 2777 9938 2778 9972
rect 2742 9904 2778 9938
rect 2742 9870 2743 9904
rect 2777 9870 2778 9904
rect 2742 9836 2778 9870
rect 2742 9802 2743 9836
rect 2777 9802 2778 9836
rect 2742 9768 2778 9802
rect 2742 9734 2743 9768
rect 2777 9734 2778 9768
rect 2742 9700 2778 9734
rect 2742 9666 2743 9700
rect 2777 9666 2778 9700
rect 2742 9632 2778 9666
rect 2742 9598 2743 9632
rect 2777 9598 2778 9632
rect 2742 9564 2778 9598
rect 2742 9530 2743 9564
rect 2777 9530 2778 9564
rect 2742 9496 2778 9530
rect 2742 9462 2743 9496
rect 2777 9462 2778 9496
rect 2742 9428 2778 9462
rect 2742 9394 2743 9428
rect 2777 9394 2778 9428
rect 2742 9360 2778 9394
rect 2742 9326 2743 9360
rect 2777 9326 2778 9360
rect 2742 9292 2778 9326
rect 2742 9258 2743 9292
rect 2777 9258 2778 9292
rect 2742 9224 2778 9258
rect 2742 9190 2743 9224
rect 2777 9190 2778 9224
rect 2742 9156 2778 9190
rect 2742 9122 2743 9156
rect 2777 9122 2778 9156
rect 2742 9088 2778 9122
rect 2742 9054 2743 9088
rect 2777 9054 2778 9088
rect 2742 9020 2778 9054
rect 2742 8986 2743 9020
rect 2777 8986 2778 9020
rect 2742 8952 2778 8986
rect 2742 8918 2743 8952
rect 2777 8918 2778 8952
rect 2742 8884 2778 8918
rect 2742 8850 2743 8884
rect 2777 8850 2778 8884
rect 2742 8816 2778 8850
rect 2742 8782 2743 8816
rect 2777 8782 2778 8816
rect 2742 8748 2778 8782
rect 2742 8714 2743 8748
rect 2777 8714 2778 8748
rect 2742 8680 2778 8714
rect 2742 8646 2743 8680
rect 2777 8646 2778 8680
rect 2742 8612 2778 8646
rect 2742 8578 2743 8612
rect 2777 8578 2778 8612
rect 2742 8544 2778 8578
rect 2742 8510 2743 8544
rect 2777 8510 2778 8544
rect 2742 8476 2778 8510
rect 2742 8442 2743 8476
rect 2777 8442 2778 8476
rect 2742 8408 2778 8442
rect 2742 8374 2743 8408
rect 2777 8374 2778 8408
rect 2742 8340 2778 8374
rect 2742 8306 2743 8340
rect 2777 8306 2778 8340
rect 2742 8272 2778 8306
rect 2742 8238 2743 8272
rect 2777 8238 2778 8272
rect 2742 8204 2778 8238
rect 2742 8170 2743 8204
rect 2777 8170 2778 8204
rect 2742 8136 2778 8170
rect 2742 8102 2743 8136
rect 2777 8102 2778 8136
rect 2742 8068 2778 8102
rect 2742 8034 2743 8068
rect 2777 8034 2778 8068
rect 2742 8000 2778 8034
rect 2742 7966 2743 8000
rect 2777 7966 2778 8000
rect 2742 7932 2778 7966
rect 2742 7898 2743 7932
rect 2777 7898 2778 7932
rect 2742 7864 2778 7898
rect 2742 7830 2743 7864
rect 2777 7830 2778 7864
rect 2742 7796 2778 7830
rect 2742 7762 2743 7796
rect 2777 7762 2778 7796
rect 2742 7728 2778 7762
rect 2742 7694 2743 7728
rect 2777 7694 2778 7728
rect 2742 7660 2778 7694
rect 2742 7626 2743 7660
rect 2777 7626 2778 7660
rect 2742 7592 2778 7626
rect 2742 7558 2743 7592
rect 2777 7558 2778 7592
rect 2742 7524 2778 7558
rect 2742 7490 2743 7524
rect 2777 7490 2778 7524
rect 2742 7456 2778 7490
rect 2742 7422 2743 7456
rect 2777 7422 2778 7456
rect 2742 7388 2778 7422
rect 2742 7354 2743 7388
rect 2777 7354 2778 7388
rect 2742 7320 2778 7354
rect 2742 7286 2743 7320
rect 2777 7286 2778 7320
rect 2742 7252 2778 7286
rect 2742 7218 2743 7252
rect 2777 7218 2778 7252
rect 2742 7184 2778 7218
rect 2742 7150 2743 7184
rect 2777 7150 2778 7184
rect 2742 7116 2778 7150
rect 2742 7082 2743 7116
rect 2777 7082 2778 7116
rect 2742 7048 2778 7082
rect 2742 7014 2743 7048
rect 2777 7014 2778 7048
rect 2742 6980 2778 7014
rect 2742 6946 2743 6980
rect 2777 6946 2778 6980
rect 2742 6912 2778 6946
rect 2742 6878 2743 6912
rect 2777 6878 2778 6912
rect 2742 6844 2778 6878
rect 2742 6810 2743 6844
rect 2777 6810 2778 6844
rect 2742 6776 2778 6810
rect 2742 6742 2743 6776
rect 2777 6742 2778 6776
rect 2742 6708 2778 6742
rect 2742 6674 2743 6708
rect 2777 6674 2778 6708
rect 2742 6640 2778 6674
rect 2742 6606 2743 6640
rect 2777 6606 2778 6640
rect 2742 6572 2778 6606
rect 4703 10708 4739 10742
rect 4908 10723 6510 10804
rect 6664 10788 6700 10822
rect 6664 10754 6665 10788
rect 6699 10754 6700 10788
rect 4703 10674 4704 10708
rect 4738 10674 4739 10708
rect 4703 10640 4739 10674
rect 4703 10606 4704 10640
rect 4738 10606 4739 10640
rect 4703 10572 4739 10606
rect 4703 10538 4704 10572
rect 4738 10538 4739 10572
rect 4703 10504 4739 10538
rect 4703 10470 4704 10504
rect 4738 10470 4739 10504
rect 4703 10436 4739 10470
rect 4703 10402 4704 10436
rect 4738 10402 4739 10436
rect 4703 10368 4739 10402
rect 4703 10334 4704 10368
rect 4738 10334 4739 10368
rect 4703 10300 4739 10334
rect 4703 10266 4704 10300
rect 4738 10266 4739 10300
rect 4703 10232 4739 10266
rect 4703 10198 4704 10232
rect 4738 10198 4739 10232
rect 4703 10164 4739 10198
rect 4703 10130 4704 10164
rect 4738 10130 4739 10164
rect 4703 10096 4739 10130
rect 4703 10062 4704 10096
rect 4738 10062 4739 10096
rect 4703 10028 4739 10062
rect 4703 9994 4704 10028
rect 4738 9994 4739 10028
rect 4703 9960 4739 9994
rect 4703 9926 4704 9960
rect 4738 9926 4739 9960
rect 4703 9892 4739 9926
rect 4703 9858 4704 9892
rect 4738 9858 4739 9892
rect 4703 9824 4739 9858
rect 4703 9790 4704 9824
rect 4738 9790 4739 9824
rect 4703 9756 4739 9790
rect 4703 9722 4704 9756
rect 4738 9722 4739 9756
rect 4703 9688 4739 9722
rect 4703 9654 4704 9688
rect 4738 9654 4739 9688
rect 4703 9620 4739 9654
rect 4703 9586 4704 9620
rect 4738 9586 4739 9620
rect 4703 9552 4739 9586
rect 4703 9518 4704 9552
rect 4738 9518 4739 9552
rect 4703 9484 4739 9518
rect 4703 9450 4704 9484
rect 4738 9450 4739 9484
rect 4703 9416 4739 9450
rect 4703 9382 4704 9416
rect 4738 9382 4739 9416
rect 4703 9348 4739 9382
rect 4703 9314 4704 9348
rect 4738 9314 4739 9348
rect 4703 9280 4739 9314
rect 4703 9246 4704 9280
rect 4738 9246 4739 9280
rect 4703 9212 4739 9246
rect 4703 9178 4704 9212
rect 4738 9178 4739 9212
rect 4703 9144 4739 9178
rect 4703 9110 4704 9144
rect 4738 9110 4739 9144
rect 4703 9076 4739 9110
rect 4703 9042 4704 9076
rect 4738 9042 4739 9076
rect 4703 9008 4739 9042
rect 4703 8974 4704 9008
rect 4738 8974 4739 9008
rect 4703 8940 4739 8974
rect 4703 8906 4704 8940
rect 4738 8906 4739 8940
rect 4703 8872 4739 8906
rect 4703 8838 4704 8872
rect 4738 8838 4739 8872
rect 4703 8804 4739 8838
rect 4703 8770 4704 8804
rect 4738 8770 4739 8804
rect 4703 8736 4739 8770
rect 4703 8702 4704 8736
rect 4738 8702 4739 8736
rect 4703 8668 4739 8702
rect 4703 8634 4704 8668
rect 4738 8634 4739 8668
rect 4703 8600 4739 8634
rect 4703 8566 4704 8600
rect 4738 8566 4739 8600
rect 4703 8532 4739 8566
rect 4703 8498 4704 8532
rect 4738 8498 4739 8532
rect 4703 8464 4739 8498
rect 4703 8430 4704 8464
rect 4738 8430 4739 8464
rect 4703 8396 4739 8430
rect 4703 8362 4704 8396
rect 4738 8362 4739 8396
rect 4703 8328 4739 8362
rect 4703 8294 4704 8328
rect 4738 8294 4739 8328
rect 4703 8260 4739 8294
rect 4703 8226 4704 8260
rect 4738 8226 4739 8260
rect 4703 8192 4739 8226
rect 4703 8158 4704 8192
rect 4738 8158 4739 8192
rect 4703 8124 4739 8158
rect 4703 8090 4704 8124
rect 4738 8090 4739 8124
rect 4703 8056 4739 8090
rect 4703 8022 4704 8056
rect 4738 8022 4739 8056
rect 4703 7988 4739 8022
rect 4703 7954 4704 7988
rect 4738 7954 4739 7988
rect 4703 7920 4739 7954
rect 4703 7886 4704 7920
rect 4738 7886 4739 7920
rect 4703 7852 4739 7886
rect 4703 7818 4704 7852
rect 4738 7818 4739 7852
rect 4703 7784 4739 7818
rect 4703 7750 4704 7784
rect 4738 7750 4739 7784
rect 4703 7716 4739 7750
rect 4703 7682 4704 7716
rect 4738 7682 4739 7716
rect 4703 7648 4739 7682
rect 4703 7614 4704 7648
rect 4738 7614 4739 7648
rect 4703 7580 4739 7614
rect 4703 7546 4704 7580
rect 4738 7546 4739 7580
rect 4703 7512 4739 7546
rect 4703 7478 4704 7512
rect 4738 7478 4739 7512
rect 4703 7444 4739 7478
rect 4703 7410 4704 7444
rect 4738 7410 4739 7444
rect 4703 7376 4739 7410
rect 4703 7342 4704 7376
rect 4738 7342 4739 7376
rect 4703 7308 4739 7342
rect 4703 7274 4704 7308
rect 4738 7274 4739 7308
rect 4703 7240 4739 7274
rect 4703 7206 4704 7240
rect 4738 7206 4739 7240
rect 4703 7172 4739 7206
rect 4703 7138 4704 7172
rect 4738 7138 4739 7172
rect 4703 7104 4739 7138
rect 4703 7070 4704 7104
rect 4738 7070 4739 7104
rect 4703 7036 4739 7070
rect 4703 7002 4704 7036
rect 4738 7002 4739 7036
rect 4703 6968 4739 7002
rect 4703 6934 4704 6968
rect 4738 6934 4739 6968
rect 4703 6900 4739 6934
rect 4703 6866 4704 6900
rect 4738 6866 4739 6900
rect 4703 6832 4739 6866
rect 4703 6798 4704 6832
rect 4738 6798 4739 6832
rect 4703 6764 4739 6798
rect 4703 6730 4704 6764
rect 4738 6730 4739 6764
rect 4703 6696 4739 6730
rect 4703 6662 4704 6696
rect 4738 6662 4739 6696
rect 4703 6628 4739 6662
rect 4703 6594 4704 6628
rect 4738 6594 4739 6628
rect 2742 6538 2743 6572
rect 2777 6538 2778 6572
rect 2742 6460 2778 6538
rect 2932 6510 4534 6591
rect 4703 6560 4739 6594
rect 6664 10720 6700 10754
rect 6664 10686 6665 10720
rect 6699 10686 6700 10720
rect 6664 10652 6700 10686
rect 6664 10618 6665 10652
rect 6699 10618 6700 10652
rect 6664 10584 6700 10618
rect 6664 10550 6665 10584
rect 6699 10550 6700 10584
rect 6664 10516 6700 10550
rect 6664 10482 6665 10516
rect 6699 10482 6700 10516
rect 6664 10448 6700 10482
rect 6664 10414 6665 10448
rect 6699 10414 6700 10448
rect 6664 10380 6700 10414
rect 6664 10346 6665 10380
rect 6699 10346 6700 10380
rect 6664 10312 6700 10346
rect 6664 10278 6665 10312
rect 6699 10278 6700 10312
rect 6664 10244 6700 10278
rect 6664 10210 6665 10244
rect 6699 10210 6700 10244
rect 6664 10176 6700 10210
rect 6664 10142 6665 10176
rect 6699 10142 6700 10176
rect 6664 10108 6700 10142
rect 6664 10074 6665 10108
rect 6699 10074 6700 10108
rect 6664 10040 6700 10074
rect 6664 10006 6665 10040
rect 6699 10006 6700 10040
rect 6664 9972 6700 10006
rect 6664 9938 6665 9972
rect 6699 9938 6700 9972
rect 6664 9904 6700 9938
rect 6664 9870 6665 9904
rect 6699 9870 6700 9904
rect 6664 9836 6700 9870
rect 6664 9802 6665 9836
rect 6699 9802 6700 9836
rect 6664 9768 6700 9802
rect 6664 9734 6665 9768
rect 6699 9734 6700 9768
rect 6664 9700 6700 9734
rect 6664 9666 6665 9700
rect 6699 9666 6700 9700
rect 6664 9632 6700 9666
rect 6664 9598 6665 9632
rect 6699 9598 6700 9632
rect 6664 9564 6700 9598
rect 6664 9530 6665 9564
rect 6699 9530 6700 9564
rect 6664 9496 6700 9530
rect 6664 9462 6665 9496
rect 6699 9462 6700 9496
rect 6664 9428 6700 9462
rect 6664 9394 6665 9428
rect 6699 9394 6700 9428
rect 6664 9360 6700 9394
rect 6664 9326 6665 9360
rect 6699 9326 6700 9360
rect 6664 9292 6700 9326
rect 6664 9258 6665 9292
rect 6699 9258 6700 9292
rect 6664 9224 6700 9258
rect 6664 9190 6665 9224
rect 6699 9190 6700 9224
rect 6664 9156 6700 9190
rect 6664 9122 6665 9156
rect 6699 9122 6700 9156
rect 6664 9088 6700 9122
rect 6664 9054 6665 9088
rect 6699 9054 6700 9088
rect 6664 9020 6700 9054
rect 6664 8986 6665 9020
rect 6699 8986 6700 9020
rect 6664 8952 6700 8986
rect 6664 8918 6665 8952
rect 6699 8918 6700 8952
rect 6664 8884 6700 8918
rect 6664 8850 6665 8884
rect 6699 8850 6700 8884
rect 6664 8816 6700 8850
rect 6664 8782 6665 8816
rect 6699 8782 6700 8816
rect 6664 8748 6700 8782
rect 6664 8714 6665 8748
rect 6699 8714 6700 8748
rect 6664 8680 6700 8714
rect 6664 8646 6665 8680
rect 6699 8646 6700 8680
rect 6664 8612 6700 8646
rect 6664 8578 6665 8612
rect 6699 8578 6700 8612
rect 6664 8544 6700 8578
rect 6664 8510 6665 8544
rect 6699 8510 6700 8544
rect 6664 8476 6700 8510
rect 6664 8442 6665 8476
rect 6699 8442 6700 8476
rect 6664 8408 6700 8442
rect 6664 8374 6665 8408
rect 6699 8374 6700 8408
rect 6664 8340 6700 8374
rect 6664 8306 6665 8340
rect 6699 8306 6700 8340
rect 6664 8272 6700 8306
rect 6664 8238 6665 8272
rect 6699 8238 6700 8272
rect 6664 8204 6700 8238
rect 6664 8170 6665 8204
rect 6699 8170 6700 8204
rect 6664 8136 6700 8170
rect 6664 8102 6665 8136
rect 6699 8102 6700 8136
rect 6664 8068 6700 8102
rect 6664 8034 6665 8068
rect 6699 8034 6700 8068
rect 6664 8000 6700 8034
rect 6664 7966 6665 8000
rect 6699 7966 6700 8000
rect 6664 7932 6700 7966
rect 6664 7898 6665 7932
rect 6699 7898 6700 7932
rect 6664 7864 6700 7898
rect 6664 7830 6665 7864
rect 6699 7830 6700 7864
rect 6664 7796 6700 7830
rect 6664 7762 6665 7796
rect 6699 7762 6700 7796
rect 6664 7728 6700 7762
rect 6664 7694 6665 7728
rect 6699 7694 6700 7728
rect 6664 7660 6700 7694
rect 6664 7626 6665 7660
rect 6699 7626 6700 7660
rect 6664 7592 6700 7626
rect 6664 7558 6665 7592
rect 6699 7558 6700 7592
rect 6664 7524 6700 7558
rect 6664 7490 6665 7524
rect 6699 7490 6700 7524
rect 6664 7456 6700 7490
rect 6664 7422 6665 7456
rect 6699 7422 6700 7456
rect 6664 7388 6700 7422
rect 6664 7354 6665 7388
rect 6699 7354 6700 7388
rect 6664 7320 6700 7354
rect 6664 7286 6665 7320
rect 6699 7286 6700 7320
rect 6664 7252 6700 7286
rect 6664 7218 6665 7252
rect 6699 7218 6700 7252
rect 6664 7184 6700 7218
rect 6664 7150 6665 7184
rect 6699 7150 6700 7184
rect 6664 7116 6700 7150
rect 6664 7082 6665 7116
rect 6699 7082 6700 7116
rect 6664 7048 6700 7082
rect 6664 7014 6665 7048
rect 6699 7014 6700 7048
rect 6664 6980 6700 7014
rect 6664 6946 6665 6980
rect 6699 6946 6700 6980
rect 6664 6912 6700 6946
rect 6664 6878 6665 6912
rect 6699 6878 6700 6912
rect 6664 6844 6700 6878
rect 6664 6810 6665 6844
rect 6699 6810 6700 6844
rect 6664 6776 6700 6810
rect 6664 6742 6665 6776
rect 6699 6742 6700 6776
rect 6664 6708 6700 6742
rect 6664 6674 6665 6708
rect 6699 6674 6700 6708
rect 6664 6640 6700 6674
rect 6664 6606 6665 6640
rect 6699 6606 6700 6640
rect 4703 6526 4704 6560
rect 4738 6526 4739 6560
rect 4703 6492 4739 6526
rect 4908 6510 6510 6591
rect 6664 6572 6700 6606
rect 6664 6538 6665 6572
rect 6699 6538 6700 6572
rect 4703 6460 4704 6492
rect 2742 6459 4704 6460
rect 2742 6425 2776 6459
rect 2810 6425 2844 6459
rect 2878 6425 2912 6459
rect 2946 6425 2980 6459
rect 3014 6425 3048 6459
rect 3082 6425 3116 6459
rect 3150 6425 3184 6459
rect 3218 6425 3252 6459
rect 3286 6425 3320 6459
rect 3354 6425 3388 6459
rect 3422 6425 3456 6459
rect 3490 6425 3524 6459
rect 3558 6425 3592 6459
rect 3626 6425 3660 6459
rect 3694 6425 3728 6459
rect 3762 6425 3796 6459
rect 3830 6425 3864 6459
rect 3898 6425 3932 6459
rect 3966 6425 4000 6459
rect 4034 6425 4068 6459
rect 4102 6425 4136 6459
rect 4170 6425 4204 6459
rect 4238 6425 4272 6459
rect 4306 6425 4340 6459
rect 4374 6425 4408 6459
rect 4442 6425 4476 6459
rect 4510 6425 4544 6459
rect 4578 6425 4612 6459
rect 4646 6458 4704 6459
rect 4738 6460 4739 6492
rect 6664 6460 6700 6538
rect 4738 6459 6700 6460
rect 4738 6458 4796 6459
rect 4646 6425 4796 6458
rect 4830 6425 4864 6459
rect 4898 6425 4932 6459
rect 4966 6425 5000 6459
rect 5034 6425 5068 6459
rect 5102 6425 5136 6459
rect 5170 6425 5204 6459
rect 5238 6425 5272 6459
rect 5306 6425 5340 6459
rect 5374 6425 5408 6459
rect 5442 6425 5476 6459
rect 5510 6425 5544 6459
rect 5578 6425 5612 6459
rect 5646 6425 5680 6459
rect 5714 6425 5748 6459
rect 5782 6425 5816 6459
rect 5850 6425 5884 6459
rect 5918 6425 5952 6459
rect 5986 6425 6020 6459
rect 6054 6425 6088 6459
rect 6122 6425 6156 6459
rect 6190 6425 6224 6459
rect 6258 6425 6292 6459
rect 6326 6425 6360 6459
rect 6394 6425 6428 6459
rect 6462 6425 6496 6459
rect 6530 6425 6564 6459
rect 6598 6425 6632 6459
rect 6666 6425 6700 6459
rect 2742 6424 6700 6425
rect 6853 10859 6889 10893
rect 6853 10825 6854 10859
rect 6888 10825 6889 10859
rect 6853 10791 6889 10825
rect 6853 10757 6854 10791
rect 6888 10757 6889 10791
rect 6853 10723 6889 10757
rect 6853 10689 6854 10723
rect 6888 10689 6889 10723
rect 6853 10655 6889 10689
rect 6853 10621 6854 10655
rect 6888 10621 6889 10655
rect 6853 10587 6889 10621
rect 6853 10553 6854 10587
rect 6888 10553 6889 10587
rect 6853 10519 6889 10553
rect 6853 10485 6854 10519
rect 6888 10485 6889 10519
rect 6853 10451 6889 10485
rect 6853 10417 6854 10451
rect 6888 10417 6889 10451
rect 6853 10383 6889 10417
rect 6853 10349 6854 10383
rect 6888 10349 6889 10383
rect 6853 10315 6889 10349
rect 6853 10281 6854 10315
rect 6888 10281 6889 10315
rect 6853 10247 6889 10281
rect 6853 10213 6854 10247
rect 6888 10213 6889 10247
rect 6853 10179 6889 10213
rect 6853 10145 6854 10179
rect 6888 10145 6889 10179
rect 6853 10111 6889 10145
rect 6853 10077 6854 10111
rect 6888 10077 6889 10111
rect 6853 10043 6889 10077
rect 6853 10009 6854 10043
rect 6888 10009 6889 10043
rect 6853 9975 6889 10009
rect 6853 9941 6854 9975
rect 6888 9941 6889 9975
rect 6853 9907 6889 9941
rect 6853 9873 6854 9907
rect 6888 9873 6889 9907
rect 6853 9839 6889 9873
rect 6853 9805 6854 9839
rect 6888 9805 6889 9839
rect 6853 9771 6889 9805
rect 6853 9737 6854 9771
rect 6888 9737 6889 9771
rect 6853 9703 6889 9737
rect 6853 9669 6854 9703
rect 6888 9669 6889 9703
rect 6853 9635 6889 9669
rect 6853 9601 6854 9635
rect 6888 9601 6889 9635
rect 6853 9567 6889 9601
rect 6853 9533 6854 9567
rect 6888 9533 6889 9567
rect 6853 9499 6889 9533
rect 6853 9465 6854 9499
rect 6888 9465 6889 9499
rect 6853 9431 6889 9465
rect 6853 9397 6854 9431
rect 6888 9397 6889 9431
rect 6853 9363 6889 9397
rect 6853 9329 6854 9363
rect 6888 9329 6889 9363
rect 6853 9295 6889 9329
rect 6853 9261 6854 9295
rect 6888 9261 6889 9295
rect 6853 9227 6889 9261
rect 6853 9193 6854 9227
rect 6888 9193 6889 9227
rect 6853 9159 6889 9193
rect 6853 9125 6854 9159
rect 6888 9125 6889 9159
rect 6853 9091 6889 9125
rect 6853 9057 6854 9091
rect 6888 9057 6889 9091
rect 6853 9023 6889 9057
rect 6853 8989 6854 9023
rect 6888 8989 6889 9023
rect 6853 8955 6889 8989
rect 6853 8921 6854 8955
rect 6888 8921 6889 8955
rect 6853 8887 6889 8921
rect 6853 8853 6854 8887
rect 6888 8853 6889 8887
rect 6853 8819 6889 8853
rect 6853 8785 6854 8819
rect 6888 8785 6889 8819
rect 6853 8751 6889 8785
rect 6853 8717 6854 8751
rect 6888 8717 6889 8751
rect 6853 8683 6889 8717
rect 6853 8649 6854 8683
rect 6888 8649 6889 8683
rect 6853 8615 6889 8649
rect 6853 8581 6854 8615
rect 6888 8581 6889 8615
rect 6853 8547 6889 8581
rect 6853 8513 6854 8547
rect 6888 8513 6889 8547
rect 6853 8479 6889 8513
rect 6853 8445 6854 8479
rect 6888 8445 6889 8479
rect 6853 8411 6889 8445
rect 6853 8377 6854 8411
rect 6888 8377 6889 8411
rect 6853 8343 6889 8377
rect 6853 8309 6854 8343
rect 6888 8309 6889 8343
rect 6853 8275 6889 8309
rect 6853 8241 6854 8275
rect 6888 8241 6889 8275
rect 6853 8207 6889 8241
rect 6853 8173 6854 8207
rect 6888 8173 6889 8207
rect 6853 8139 6889 8173
rect 6853 8105 6854 8139
rect 6888 8105 6889 8139
rect 6853 8071 6889 8105
rect 6853 8037 6854 8071
rect 6888 8037 6889 8071
rect 6853 8003 6889 8037
rect 6853 7969 6854 8003
rect 6888 7969 6889 8003
rect 6853 7935 6889 7969
rect 6853 7901 6854 7935
rect 6888 7901 6889 7935
rect 6853 7867 6889 7901
rect 6853 7833 6854 7867
rect 6888 7833 6889 7867
rect 6853 7799 6889 7833
rect 6853 7765 6854 7799
rect 6888 7765 6889 7799
rect 6853 7731 6889 7765
rect 6853 7697 6854 7731
rect 6888 7697 6889 7731
rect 6853 7663 6889 7697
rect 6853 7629 6854 7663
rect 6888 7629 6889 7663
rect 6853 7595 6889 7629
rect 6853 7561 6854 7595
rect 6888 7561 6889 7595
rect 6853 7527 6889 7561
rect 6853 7493 6854 7527
rect 6888 7493 6889 7527
rect 6853 7459 6889 7493
rect 6853 7425 6854 7459
rect 6888 7425 6889 7459
rect 6853 7391 6889 7425
rect 6853 7357 6854 7391
rect 6888 7357 6889 7391
rect 6853 7323 6889 7357
rect 6853 7289 6854 7323
rect 6888 7289 6889 7323
rect 6853 7255 6889 7289
rect 6853 7221 6854 7255
rect 6888 7221 6889 7255
rect 6853 7187 6889 7221
rect 6853 7153 6854 7187
rect 6888 7153 6889 7187
rect 6853 7119 6889 7153
rect 6853 7085 6854 7119
rect 6888 7085 6889 7119
rect 6853 7051 6889 7085
rect 6853 7017 6854 7051
rect 6888 7017 6889 7051
rect 6853 6983 6889 7017
rect 6853 6949 6854 6983
rect 6888 6949 6889 6983
rect 6853 6915 6889 6949
rect 6853 6881 6854 6915
rect 6888 6881 6889 6915
rect 6853 6847 6889 6881
rect 6853 6813 6854 6847
rect 6888 6813 6889 6847
rect 6853 6779 6889 6813
rect 6853 6745 6854 6779
rect 6888 6745 6889 6779
rect 6853 6711 6889 6745
rect 6853 6677 6854 6711
rect 6888 6677 6889 6711
rect 6853 6643 6889 6677
rect 6853 6609 6854 6643
rect 6888 6609 6889 6643
rect 6853 6575 6889 6609
rect 6853 6541 6854 6575
rect 6888 6541 6889 6575
rect 6853 6507 6889 6541
rect 6853 6473 6854 6507
rect 6888 6473 6889 6507
rect 6853 6439 6889 6473
rect 2553 6385 2589 6419
rect 2553 6351 2554 6385
rect 2588 6351 2589 6385
rect 2553 6271 2589 6351
rect 6853 6405 6854 6439
rect 6888 6405 6889 6439
rect 6853 6371 6889 6405
rect 6853 6337 6854 6371
rect 6888 6337 6889 6371
rect 6853 6303 6889 6337
rect 6853 6271 6854 6303
rect 2553 6270 6854 6271
rect 2553 6236 2587 6270
rect 2621 6236 2655 6270
rect 2689 6236 2723 6270
rect 2757 6236 2791 6270
rect 2825 6236 2859 6270
rect 2893 6236 2927 6270
rect 2961 6236 2995 6270
rect 3029 6236 3063 6270
rect 3097 6236 3131 6270
rect 3165 6236 3199 6270
rect 3233 6236 3267 6270
rect 3301 6236 3335 6270
rect 3369 6236 3403 6270
rect 3437 6236 3471 6270
rect 3505 6236 3539 6270
rect 3573 6236 3607 6270
rect 3641 6236 3675 6270
rect 3709 6236 3743 6270
rect 3777 6236 3811 6270
rect 3845 6236 3879 6270
rect 3913 6236 3947 6270
rect 3981 6236 4015 6270
rect 4049 6236 4083 6270
rect 4117 6236 4151 6270
rect 4185 6236 4219 6270
rect 4253 6236 4287 6270
rect 4321 6236 4355 6270
rect 4389 6236 4423 6270
rect 4457 6236 4491 6270
rect 4525 6236 4559 6270
rect 4593 6236 4627 6270
rect 4661 6236 4695 6270
rect 4729 6236 4763 6270
rect 4797 6236 4831 6270
rect 4865 6236 4899 6270
rect 4933 6236 4967 6270
rect 5001 6236 5035 6270
rect 5069 6236 5103 6270
rect 5137 6236 5171 6270
rect 5205 6236 5239 6270
rect 5273 6236 5307 6270
rect 5341 6236 5375 6270
rect 5409 6236 5443 6270
rect 5477 6236 5511 6270
rect 5545 6236 5579 6270
rect 5613 6236 5647 6270
rect 5681 6236 5715 6270
rect 5749 6236 5783 6270
rect 5817 6236 5851 6270
rect 5885 6236 5919 6270
rect 5953 6236 5987 6270
rect 6021 6236 6055 6270
rect 6089 6236 6123 6270
rect 6157 6236 6191 6270
rect 6225 6236 6259 6270
rect 6293 6236 6327 6270
rect 6361 6236 6395 6270
rect 6429 6236 6463 6270
rect 6497 6236 6531 6270
rect 6565 6236 6599 6270
rect 6633 6236 6667 6270
rect 6701 6236 6735 6270
rect 6769 6269 6854 6270
rect 6888 6269 6889 6303
rect 6769 6236 6889 6269
rect 2553 6235 6889 6236
rect 2333 6192 2369 6207
rect 2333 6139 2334 6192
rect 2368 6139 2369 6192
rect 2333 6135 2369 6139
rect 6854 6211 6888 6235
rect 6854 6139 6888 6177
rect 2333 6105 6854 6135
rect 2333 6071 2357 6105
rect 2391 6071 2426 6105
rect 2460 6071 2495 6105
rect 2529 6071 2564 6105
rect 2598 6071 2633 6105
rect 2667 6071 2702 6105
rect 2736 6071 2771 6105
rect 2805 6071 2840 6105
rect 2874 6071 2909 6105
rect 2943 6071 2978 6105
rect 3012 6071 3047 6105
rect 3081 6071 3116 6105
rect 3150 6071 3185 6105
rect 3219 6071 3254 6105
rect 3288 6071 3323 6105
rect 3357 6071 3392 6105
rect 3426 6071 3461 6105
rect 3495 6071 3530 6105
rect 3564 6071 3599 6105
rect 3633 6071 3668 6105
rect 3702 6071 3737 6105
rect 3771 6071 3806 6105
rect 3840 6071 3875 6105
rect 3909 6071 3944 6105
rect 3978 6071 4013 6105
rect 4047 6071 4082 6105
rect 4116 6071 4151 6105
rect 4185 6071 4220 6105
rect 4254 6071 4289 6105
rect 4323 6071 4358 6105
rect 4392 6071 4427 6105
rect 4461 6071 4496 6105
rect 4530 6071 4565 6105
rect 4599 6071 4634 6105
rect 4668 6071 4703 6105
rect 4737 6071 4772 6105
rect 4806 6071 4841 6105
rect 4875 6071 4910 6105
rect 4944 6071 4979 6105
rect 5013 6071 5048 6105
rect 5082 6071 5117 6105
rect 5151 6071 5186 6105
rect 5220 6071 5255 6105
rect 5289 6071 5324 6105
rect 5358 6071 5392 6105
rect 5426 6071 5460 6105
rect 5494 6071 5528 6105
rect 5562 6071 5596 6105
rect 5630 6071 5664 6105
rect 5698 6071 5732 6105
rect 5766 6071 5800 6105
rect 5834 6071 5868 6105
rect 5902 6071 5936 6105
rect 5970 6071 6004 6105
rect 6038 6071 6072 6105
rect 6106 6071 6140 6105
rect 6174 6071 6208 6105
rect 6242 6071 6276 6105
rect 6310 6071 6344 6105
rect 6378 6071 6412 6105
rect 6446 6071 6480 6105
rect 6514 6071 6548 6105
rect 6582 6071 6616 6105
rect 6650 6071 6684 6105
rect 6718 6071 6752 6105
rect 6786 6071 6888 6105
rect 2144 6015 2180 6049
rect 2144 5981 2145 6015
rect 2179 5981 2180 6015
rect 2144 5947 2180 5981
rect 2144 5913 2145 5947
rect 2179 5913 2180 5947
rect 2144 5879 2180 5913
rect 2144 5845 2145 5879
rect 2179 5845 2180 5879
rect 2144 5811 2180 5845
rect 2144 5777 2145 5811
rect 2179 5777 2180 5811
rect 2144 5743 2180 5777
rect 2144 5709 2145 5743
rect 2179 5709 2180 5743
rect 2144 5675 2180 5709
rect 2144 5641 2145 5675
rect 2179 5641 2180 5675
rect 5453 5959 5465 5993
rect 5499 5959 5537 5993
rect 2144 5607 2180 5641
rect 2144 5573 2145 5607
rect 2179 5575 2180 5607
rect 2382 5620 2388 5654
rect 2422 5620 2460 5654
rect 2179 5574 2348 5575
rect 2179 5573 2230 5574
rect 231 5536 253 5549
rect 287 5536 330 5570
rect 231 5510 330 5536
rect 265 5502 330 5510
rect 231 5468 253 5476
rect 287 5468 330 5502
rect 231 5437 330 5468
rect 265 5403 330 5437
rect 231 5402 330 5403
rect 265 5368 330 5402
rect 231 5364 330 5368
rect 265 5330 330 5364
rect 231 5329 330 5330
rect 265 5295 330 5329
rect 231 5291 330 5295
rect 265 5257 330 5291
rect 231 5256 330 5257
rect 265 5222 330 5256
rect 231 5218 330 5222
rect 265 5184 330 5218
rect 231 5183 330 5184
rect 265 5149 330 5183
rect 1878 5564 1944 5570
rect 1878 5530 1894 5564
rect 1928 5530 1944 5564
rect 1878 5492 1944 5530
rect 1878 5458 1894 5492
rect 1928 5458 1944 5492
rect 1878 5270 1944 5458
rect 2004 5564 2070 5570
rect 2004 5530 2020 5564
rect 2054 5530 2070 5564
rect 2144 5540 2230 5573
rect 2264 5540 2280 5574
rect 2336 5540 2348 5574
rect 2144 5539 2348 5540
rect 2004 5492 2070 5530
rect 2004 5458 2020 5492
rect 2054 5458 2070 5492
rect 2004 5457 2070 5458
rect 2382 5457 2448 5620
rect 3530 5575 5419 5576
rect 2482 5574 3188 5575
rect 2482 5540 2576 5574
rect 2610 5540 2644 5574
rect 2678 5540 2712 5574
rect 2746 5540 2780 5574
rect 2814 5540 2848 5574
rect 2882 5540 2916 5574
rect 2950 5540 2984 5574
rect 3018 5540 3052 5574
rect 3086 5540 3120 5574
rect 3154 5540 3188 5574
rect 2482 5539 3188 5540
rect 3152 5498 3188 5539
rect 3152 5458 3153 5498
rect 3187 5458 3188 5498
rect 2004 5423 2020 5457
rect 2054 5423 2070 5457
rect 2004 5389 2070 5423
rect 2130 5423 2146 5457
rect 2180 5423 2196 5457
rect 2130 5389 2196 5423
rect 2256 5423 2272 5457
rect 2306 5423 2322 5457
rect 2256 5389 2322 5423
rect 2382 5423 2398 5457
rect 2432 5423 2448 5457
rect 1878 5236 1894 5270
rect 1928 5236 1944 5270
rect 1878 5198 1944 5236
rect 1878 5164 1894 5198
rect 1928 5164 1944 5198
rect 1878 5158 1944 5164
rect 2004 5270 2070 5355
rect 2004 5236 2020 5270
rect 2054 5236 2070 5270
rect 2004 5198 2070 5236
rect 2004 5164 2020 5198
rect 2054 5164 2070 5198
rect 2004 5158 2070 5164
rect 2130 5270 2196 5355
rect 2130 5236 2146 5270
rect 2180 5236 2196 5270
rect 2130 5198 2196 5236
rect 2130 5164 2146 5198
rect 2180 5164 2196 5198
rect 2130 5158 2196 5164
rect 2256 5270 2322 5355
rect 2256 5236 2272 5270
rect 2306 5236 2322 5270
rect 2256 5198 2322 5236
rect 2256 5164 2272 5198
rect 2306 5164 2322 5198
rect 2256 5158 2322 5164
rect 2382 5270 2448 5423
rect 2508 5423 2524 5457
rect 2558 5423 2574 5457
rect 2508 5389 2574 5423
rect 2634 5423 2650 5457
rect 2684 5423 2700 5457
rect 2634 5389 2700 5423
rect 2760 5423 2776 5457
rect 2810 5423 2826 5457
rect 2760 5389 2826 5423
rect 2886 5423 2902 5457
rect 2936 5423 2952 5457
rect 2886 5389 2952 5423
rect 3012 5423 3028 5457
rect 3062 5423 3078 5457
rect 3012 5389 3078 5423
rect 3152 5424 3188 5458
rect 3152 5390 3153 5424
rect 3187 5390 3188 5424
rect 3152 5356 3188 5390
rect 2382 5236 2398 5270
rect 2432 5236 2448 5270
rect 2382 5198 2448 5236
rect 2382 5164 2398 5198
rect 2432 5164 2448 5198
rect 2382 5158 2448 5164
rect 2508 5270 2574 5355
rect 2508 5236 2524 5270
rect 2558 5236 2574 5270
rect 2508 5198 2574 5236
rect 2508 5164 2524 5198
rect 2558 5164 2574 5198
rect 2508 5158 2574 5164
rect 2634 5270 2700 5355
rect 2634 5236 2650 5270
rect 2684 5236 2700 5270
rect 2634 5198 2700 5236
rect 2634 5164 2650 5198
rect 2684 5164 2700 5198
rect 2634 5158 2700 5164
rect 2760 5270 2826 5355
rect 2760 5236 2776 5270
rect 2810 5236 2826 5270
rect 2760 5198 2826 5236
rect 2760 5164 2776 5198
rect 2810 5164 2826 5198
rect 2760 5158 2826 5164
rect 2886 5270 2952 5355
rect 2886 5236 2902 5270
rect 2936 5236 2952 5270
rect 2886 5198 2952 5236
rect 2886 5164 2902 5198
rect 2936 5164 2952 5198
rect 2886 5158 2952 5164
rect 3012 5270 3078 5355
rect 3012 5236 3028 5270
rect 3062 5236 3078 5270
rect 3012 5198 3078 5236
rect 3012 5164 3028 5198
rect 3062 5164 3078 5198
rect 3012 5158 3078 5164
rect 3152 5322 3153 5356
rect 3187 5322 3188 5356
rect 3152 5288 3188 5322
rect 3152 5254 3153 5288
rect 3187 5254 3188 5288
rect 3152 5220 3188 5254
rect 3152 5186 3153 5220
rect 3187 5186 3188 5220
rect 231 5145 330 5149
rect 265 5111 330 5145
rect 231 5110 330 5111
rect 265 5076 330 5110
rect 231 5072 330 5076
rect 265 5038 330 5072
rect 231 5037 330 5038
rect 265 5003 330 5037
rect 231 4999 330 5003
rect 265 4931 330 4999
rect 231 4926 330 4931
rect 265 4859 330 4926
rect 231 4853 330 4859
rect 265 4787 330 4853
rect 231 4780 330 4787
rect 265 4715 330 4780
rect 231 4707 330 4715
rect 265 4643 330 4707
rect 3152 5152 3188 5186
rect 3152 5118 3153 5152
rect 3187 5118 3188 5152
rect 3152 5084 3188 5118
rect 3152 5050 3153 5084
rect 3187 5050 3188 5084
rect 3152 5016 3188 5050
rect 3152 4982 3153 5016
rect 3187 4982 3188 5016
rect 3152 4948 3188 4982
rect 3152 4914 3153 4948
rect 3187 4914 3188 4948
rect 3152 4880 3188 4914
rect 3152 4846 3153 4880
rect 3187 4846 3188 4880
rect 3152 4812 3188 4846
rect 3152 4778 3153 4812
rect 3187 4778 3188 4812
rect 3152 4744 3188 4778
rect 3152 4710 3153 4744
rect 3187 4710 3188 4744
rect 3152 4676 3188 4710
rect 231 4634 330 4643
rect 265 4571 330 4634
rect 231 4561 330 4571
rect 265 4499 330 4561
rect 231 4488 330 4499
rect 265 4427 330 4488
rect 231 4415 330 4427
rect 265 4381 330 4415
rect 1248 4644 1314 4656
rect 1248 4610 1264 4644
rect 1298 4610 1314 4644
rect 1248 4572 1314 4610
rect 1248 4538 1264 4572
rect 1298 4538 1314 4572
rect 231 4353 330 4381
rect 231 4333 257 4353
rect 291 4319 330 4353
rect 265 4299 330 4319
rect 231 4284 330 4299
rect 231 4257 257 4284
rect 256 4250 257 4257
rect 291 4250 330 4284
rect 256 4215 330 4250
rect 256 4181 257 4215
rect 291 4181 330 4215
rect 256 4146 330 4181
rect 256 4112 257 4146
rect 291 4112 330 4146
rect 256 4077 330 4112
rect 256 4043 257 4077
rect 291 4043 330 4077
rect 256 4008 330 4043
rect 256 3974 257 4008
rect 291 3974 330 4008
rect 366 4387 432 4399
rect 366 4353 382 4387
rect 416 4353 432 4387
rect 366 4315 432 4353
rect 366 4269 382 4315
rect 416 4269 432 4315
rect 366 4193 432 4269
rect 366 4159 382 4193
rect 416 4159 432 4193
rect 366 4107 432 4159
rect 366 4073 382 4107
rect 416 4073 432 4107
rect 366 4035 432 4073
rect 366 4001 382 4035
rect 416 4001 432 4035
rect 366 3989 432 4001
rect 492 4387 558 4399
rect 492 4353 508 4387
rect 542 4353 558 4387
rect 492 4315 558 4353
rect 492 4269 508 4315
rect 542 4269 558 4315
rect 492 4193 558 4269
rect 492 4159 508 4193
rect 542 4159 558 4193
rect 492 4107 558 4159
rect 492 4073 508 4107
rect 542 4073 558 4107
rect 492 4035 558 4073
rect 492 4001 508 4035
rect 542 4001 558 4035
rect 492 3989 558 4001
rect 618 4387 684 4399
rect 618 4353 634 4387
rect 668 4353 684 4387
rect 618 4315 684 4353
rect 618 4269 634 4315
rect 668 4269 684 4315
rect 618 4193 684 4269
rect 618 4159 634 4193
rect 668 4159 684 4193
rect 618 4107 684 4159
rect 618 4073 634 4107
rect 668 4073 684 4107
rect 618 4035 684 4073
rect 618 4001 634 4035
rect 668 4001 684 4035
rect 618 3989 684 4001
rect 744 4387 810 4399
rect 744 4353 760 4387
rect 794 4353 810 4387
rect 744 4315 810 4353
rect 744 4269 760 4315
rect 794 4269 810 4315
rect 744 4193 810 4269
rect 744 4159 760 4193
rect 794 4159 810 4193
rect 744 4107 810 4159
rect 744 4073 760 4107
rect 794 4073 810 4107
rect 744 4035 810 4073
rect 744 4001 760 4035
rect 794 4001 810 4035
rect 744 3989 810 4001
rect 870 4387 936 4399
rect 870 4353 886 4387
rect 920 4353 936 4387
rect 870 4315 936 4353
rect 870 4269 886 4315
rect 920 4269 936 4315
rect 870 4193 936 4269
rect 870 4159 886 4193
rect 920 4159 936 4193
rect 870 4107 936 4159
rect 870 4073 886 4107
rect 920 4073 936 4107
rect 870 4035 936 4073
rect 870 4001 886 4035
rect 920 4001 936 4035
rect 870 3989 936 4001
rect 996 4387 1062 4399
rect 996 4353 1012 4387
rect 1046 4353 1062 4387
rect 996 4315 1062 4353
rect 996 4269 1012 4315
rect 1046 4269 1062 4315
rect 996 4193 1062 4269
rect 996 4159 1012 4193
rect 1046 4159 1062 4193
rect 996 4107 1062 4159
rect 996 4073 1012 4107
rect 1046 4073 1062 4107
rect 996 4035 1062 4073
rect 996 4001 1012 4035
rect 1046 4001 1062 4035
rect 996 3989 1062 4001
rect 1122 4387 1188 4399
rect 1122 4353 1138 4387
rect 1172 4353 1188 4387
rect 1122 4315 1188 4353
rect 1122 4269 1138 4315
rect 1172 4269 1188 4315
rect 1122 4193 1188 4269
rect 1122 4159 1138 4193
rect 1172 4159 1188 4193
rect 1122 4107 1188 4159
rect 1122 4073 1138 4107
rect 1172 4073 1188 4107
rect 1122 4035 1188 4073
rect 1122 4001 1138 4035
rect 1172 4001 1188 4035
rect 1122 3989 1188 4001
rect 1248 4303 1314 4538
rect 3152 4642 3153 4676
rect 3187 4642 3188 4676
rect 3152 4608 3188 4642
rect 3152 4574 3153 4608
rect 3187 4574 3188 4608
rect 3152 4540 3188 4574
rect 3152 4506 3153 4540
rect 3187 4506 3188 4540
rect 3152 4472 3188 4506
rect 3152 4438 3153 4472
rect 3187 4438 3188 4472
rect 1248 4269 1264 4303
rect 1298 4269 1314 4303
rect 1248 4193 1314 4269
rect 1248 4159 1264 4193
rect 1298 4159 1314 4193
rect 1248 4107 1314 4159
rect 1248 4073 1264 4107
rect 1298 4073 1314 4107
rect 1248 4035 1314 4073
rect 1248 4001 1264 4035
rect 1298 4001 1314 4035
rect 1248 3989 1314 4001
rect 1374 4407 1440 4419
rect 1374 4373 1390 4407
rect 1424 4373 1440 4407
rect 1374 4335 1440 4373
rect 1374 4269 1390 4335
rect 1424 4269 1440 4335
rect 1374 4193 1440 4269
rect 1374 4159 1390 4193
rect 1424 4159 1440 4193
rect 1374 4107 1440 4159
rect 1374 4073 1390 4107
rect 1424 4073 1440 4107
rect 1374 4035 1440 4073
rect 1374 4001 1390 4035
rect 1424 4001 1440 4035
rect 1374 3989 1440 4001
rect 1500 4407 1566 4419
rect 1500 4373 1516 4407
rect 1550 4373 1566 4407
rect 1500 4335 1566 4373
rect 1500 4269 1516 4335
rect 1550 4269 1566 4335
rect 1500 4193 1566 4269
rect 1500 4159 1516 4193
rect 1550 4159 1566 4193
rect 1500 4107 1566 4159
rect 1500 4073 1516 4107
rect 1550 4073 1566 4107
rect 1500 4035 1566 4073
rect 1500 4001 1516 4035
rect 1550 4001 1566 4035
rect 1500 3989 1566 4001
rect 1626 4407 1692 4419
rect 1626 4373 1642 4407
rect 1676 4373 1692 4407
rect 1626 4335 1692 4373
rect 1626 4269 1642 4335
rect 1676 4269 1692 4335
rect 1626 4193 1692 4269
rect 1626 4159 1642 4193
rect 1676 4159 1692 4193
rect 1626 4107 1692 4159
rect 1626 4073 1642 4107
rect 1676 4073 1692 4107
rect 1626 4035 1692 4073
rect 1626 4001 1642 4035
rect 1676 4001 1692 4035
rect 1626 3989 1692 4001
rect 1752 4407 1818 4419
rect 1752 4373 1768 4407
rect 1802 4373 1818 4407
rect 1752 4335 1818 4373
rect 1752 4269 1768 4335
rect 1802 4269 1818 4335
rect 1752 4193 1818 4269
rect 1752 4159 1768 4193
rect 1802 4159 1818 4193
rect 1752 4107 1818 4159
rect 1752 4073 1768 4107
rect 1802 4073 1818 4107
rect 1752 4035 1818 4073
rect 1752 4001 1768 4035
rect 1802 4001 1818 4035
rect 1752 3989 1818 4001
rect 1878 4407 1944 4419
rect 1878 4373 1894 4407
rect 1928 4373 1944 4407
rect 1878 4335 1944 4373
rect 1878 4269 1894 4335
rect 1928 4269 1944 4335
rect 1878 4193 1944 4269
rect 1878 4159 1894 4193
rect 1928 4159 1944 4193
rect 1878 4072 1944 4159
rect 1878 4038 1894 4072
rect 1928 4038 1944 4072
rect 1878 4000 1944 4038
rect 256 3939 330 3974
rect 1878 3966 1894 4000
rect 1928 3966 1944 4000
rect 2004 4407 2070 4413
rect 2004 4373 2020 4407
rect 2054 4373 2070 4407
rect 2004 4335 2070 4373
rect 2004 4301 2020 4335
rect 2054 4301 2070 4335
rect 2004 4107 2070 4301
rect 2004 4073 2020 4107
rect 2054 4073 2070 4107
rect 2004 4035 2070 4073
rect 2004 4001 2020 4035
rect 2054 4001 2070 4035
rect 2004 3989 2070 4001
rect 2130 4407 2196 4413
rect 2130 4373 2146 4407
rect 2180 4373 2196 4407
rect 2130 4335 2196 4373
rect 2130 4301 2146 4335
rect 2180 4301 2196 4335
rect 2130 4072 2196 4301
rect 2130 4038 2146 4072
rect 2180 4038 2196 4072
rect 2130 4000 2196 4038
rect 1878 3954 1944 3966
rect 2130 3966 2146 4000
rect 2180 3966 2196 4000
rect 2256 4407 2322 4413
rect 2256 4373 2272 4407
rect 2306 4373 2322 4407
rect 2256 4335 2322 4373
rect 2256 4301 2272 4335
rect 2306 4301 2322 4335
rect 2256 4107 2322 4301
rect 2256 4073 2272 4107
rect 2306 4073 2322 4107
rect 2256 4035 2322 4073
rect 2256 4001 2272 4035
rect 2306 4001 2322 4035
rect 2256 3989 2322 4001
rect 2382 4407 2448 4413
rect 2382 4373 2398 4407
rect 2432 4373 2448 4407
rect 2382 4335 2448 4373
rect 2382 4301 2398 4335
rect 2432 4301 2448 4335
rect 2382 4072 2448 4301
rect 2382 4038 2398 4072
rect 2432 4038 2448 4072
rect 2382 4000 2448 4038
rect 2130 3954 2196 3966
rect 2382 3966 2398 4000
rect 2432 3966 2448 4000
rect 2508 4407 2574 4413
rect 2508 4373 2524 4407
rect 2558 4373 2574 4407
rect 2508 4335 2574 4373
rect 2508 4301 2524 4335
rect 2558 4301 2574 4335
rect 2508 4107 2574 4301
rect 2508 4073 2524 4107
rect 2558 4073 2574 4107
rect 2508 4035 2574 4073
rect 2508 4001 2524 4035
rect 2558 4001 2574 4035
rect 2508 3989 2574 4001
rect 2634 4407 2700 4413
rect 2634 4373 2650 4407
rect 2684 4373 2700 4407
rect 2634 4335 2700 4373
rect 2634 4301 2650 4335
rect 2684 4301 2700 4335
rect 2634 4072 2700 4301
rect 2634 4038 2650 4072
rect 2684 4038 2700 4072
rect 2634 4000 2700 4038
rect 2382 3954 2448 3966
rect 2634 3966 2650 4000
rect 2684 3966 2700 4000
rect 2760 4407 2826 4413
rect 2760 4373 2776 4407
rect 2810 4373 2826 4407
rect 2760 4335 2826 4373
rect 2760 4301 2776 4335
rect 2810 4301 2826 4335
rect 2760 4107 2826 4301
rect 2760 4073 2776 4107
rect 2810 4073 2826 4107
rect 2760 4035 2826 4073
rect 2760 4001 2776 4035
rect 2810 4001 2826 4035
rect 2760 3989 2826 4001
rect 2886 4407 2952 4413
rect 2886 4373 2902 4407
rect 2936 4373 2952 4407
rect 2886 4335 2952 4373
rect 2886 4301 2902 4335
rect 2936 4301 2952 4335
rect 2886 4019 2952 4301
rect 2634 3954 2700 3966
rect 2886 3985 2902 4019
rect 2936 3985 2952 4019
rect 3012 4407 3078 4413
rect 3012 4373 3028 4407
rect 3062 4373 3078 4407
rect 3012 4335 3078 4373
rect 3012 4301 3028 4335
rect 3062 4301 3078 4335
rect 3012 4107 3078 4301
rect 3012 4073 3028 4107
rect 3062 4073 3078 4107
rect 3012 4035 3078 4073
rect 3012 4001 3028 4035
rect 3062 4001 3078 4035
rect 3012 3989 3078 4001
rect 3152 4404 3188 4438
rect 3152 4370 3153 4404
rect 3187 4370 3188 4404
rect 3152 4336 3188 4370
rect 3152 4302 3153 4336
rect 3187 4302 3188 4336
rect 3152 4268 3188 4302
rect 3530 5542 3651 5575
rect 3530 5508 3531 5542
rect 3565 5541 3651 5542
rect 3685 5541 3719 5575
rect 3753 5541 3787 5575
rect 3821 5541 3855 5575
rect 3889 5541 3923 5575
rect 3957 5541 3991 5575
rect 4025 5541 4059 5575
rect 4093 5541 4127 5575
rect 4161 5541 4195 5575
rect 4229 5541 4263 5575
rect 4297 5541 4331 5575
rect 4365 5541 4399 5575
rect 4433 5541 4467 5575
rect 4501 5541 4535 5575
rect 4569 5541 4603 5575
rect 4637 5541 4671 5575
rect 4705 5541 4739 5575
rect 4773 5541 4807 5575
rect 4841 5541 4875 5575
rect 4909 5541 4943 5575
rect 4977 5541 5011 5575
rect 5045 5541 5079 5575
rect 5113 5541 5147 5575
rect 5181 5541 5215 5575
rect 5249 5541 5283 5575
rect 5317 5541 5351 5575
rect 5385 5541 5419 5575
rect 3565 5540 5419 5541
rect 3565 5508 3566 5540
rect 3530 5498 3566 5508
rect 3530 5440 3531 5498
rect 3565 5440 3566 5498
rect 5453 5492 5495 5959
rect 5529 5575 5656 5576
rect 5529 5541 5588 5575
rect 5622 5541 5656 5575
rect 5529 5540 5656 5541
rect 4954 5458 4962 5492
rect 5004 5458 5034 5492
rect 5072 5458 5106 5492
rect 5140 5458 5174 5492
rect 5212 5458 5224 5492
rect 5293 5458 5309 5492
rect 5343 5458 5377 5492
rect 5411 5458 5445 5492
rect 5479 5458 5495 5492
rect 3530 5406 3566 5440
rect 3530 5372 3531 5406
rect 3565 5372 3566 5406
rect 3530 5338 3566 5372
rect 3530 5304 3531 5338
rect 3565 5304 3566 5338
rect 3530 5270 3566 5304
rect 3530 5236 3531 5270
rect 3565 5236 3566 5270
rect 5620 5456 5656 5540
rect 5620 5422 5621 5456
rect 5655 5422 5656 5456
rect 5620 5388 5656 5422
rect 5620 5354 5621 5388
rect 5655 5354 5656 5388
rect 5620 5320 5656 5354
rect 5620 5286 5621 5320
rect 5655 5286 5656 5320
rect 5620 5252 5656 5286
rect 3530 5202 3566 5236
rect 3530 5168 3531 5202
rect 3565 5168 3566 5202
rect 3530 5134 3566 5168
rect 3530 5100 3531 5134
rect 3565 5100 3566 5134
rect 3530 5066 3566 5100
rect 3530 5032 3531 5066
rect 3565 5032 3566 5066
rect 3530 4998 3566 5032
rect 3530 4964 3531 4998
rect 3565 4964 3566 4998
rect 3530 4930 3566 4964
rect 3530 4896 3531 4930
rect 3565 4896 3566 4930
rect 3530 4862 3566 4896
rect 3530 4828 3531 4862
rect 3565 4828 3566 4862
rect 3530 4794 3566 4828
rect 3530 4760 3531 4794
rect 3565 4760 3566 4794
rect 3530 4726 3566 4760
rect 3530 4692 3531 4726
rect 3565 4692 3566 4726
rect 5504 5166 5538 5214
rect 5504 5084 5538 5132
rect 5504 5002 5538 5050
rect 5504 4920 5538 4968
rect 5504 4838 5538 4886
rect 5504 4755 5538 4804
rect 5620 5218 5621 5252
rect 5655 5218 5656 5252
rect 5620 5184 5656 5218
rect 5620 5150 5621 5184
rect 5655 5150 5656 5184
rect 5620 5116 5656 5150
rect 5620 5082 5621 5116
rect 5655 5082 5656 5116
rect 5620 5048 5656 5082
rect 5620 5014 5621 5048
rect 5655 5014 5656 5048
rect 5620 4980 5656 5014
rect 5620 4946 5621 4980
rect 5655 4946 5656 4980
rect 5620 4912 5656 4946
rect 5620 4878 5621 4912
rect 5655 4878 5656 4912
rect 5620 4844 5656 4878
rect 5620 4810 5621 4844
rect 5655 4810 5656 4844
rect 5620 4776 5656 4810
rect 5620 4742 5621 4776
rect 5655 4742 5656 4776
rect 3530 4658 3566 4692
rect 3530 4624 3531 4658
rect 3565 4624 3566 4658
rect 3530 4590 3566 4624
rect 3530 4556 3531 4590
rect 3565 4556 3566 4590
rect 3530 4522 3566 4556
rect 3530 4488 3531 4522
rect 3565 4488 3566 4522
rect 3530 4454 3566 4488
rect 3530 4420 3531 4454
rect 3565 4420 3566 4454
rect 3530 4336 3566 4420
rect 5620 4708 5656 4742
rect 5620 4674 5621 4708
rect 5655 4674 5656 4708
rect 5620 4640 5656 4674
rect 5620 4606 5621 4640
rect 5655 4606 5656 4640
rect 5620 4572 5656 4606
rect 5620 4538 5621 4572
rect 5655 4538 5656 4572
rect 5620 4504 5656 4538
rect 5620 4470 5621 4504
rect 5655 4470 5656 4504
rect 5620 4436 5656 4470
rect 5620 4402 5621 4436
rect 5655 4402 5656 4436
rect 5620 4368 5656 4402
rect 5620 4336 5621 4368
rect 3530 4335 5621 4336
rect 3530 4301 3564 4335
rect 3598 4301 3632 4335
rect 3666 4301 3700 4335
rect 3734 4301 3768 4335
rect 3802 4301 3836 4335
rect 3870 4301 3904 4335
rect 3938 4301 3972 4335
rect 4006 4301 4040 4335
rect 4074 4301 4108 4335
rect 4142 4301 4176 4335
rect 4210 4301 4244 4335
rect 4278 4301 4312 4335
rect 4346 4301 4380 4335
rect 4414 4301 4448 4335
rect 4482 4301 4516 4335
rect 4550 4301 4584 4335
rect 4618 4301 4652 4335
rect 4686 4301 4720 4335
rect 4754 4301 4788 4335
rect 4822 4301 4856 4335
rect 4890 4301 4924 4335
rect 4958 4301 4992 4335
rect 5026 4301 5060 4335
rect 5094 4301 5128 4335
rect 5162 4301 5196 4335
rect 5230 4301 5264 4335
rect 5298 4301 5332 4335
rect 5366 4301 5400 4335
rect 5434 4301 5468 4335
rect 5502 4301 5536 4335
rect 5570 4334 5621 4335
rect 5655 4334 5656 4368
rect 5570 4301 5656 4334
rect 3530 4300 5656 4301
rect 3152 4234 3153 4268
rect 3187 4234 3188 4268
rect 3152 4200 3188 4234
rect 3152 4166 3153 4200
rect 3187 4166 3188 4200
rect 3152 4132 3188 4166
rect 3152 4098 3153 4132
rect 3187 4098 3188 4132
rect 3152 4064 3188 4098
rect 3152 4030 3153 4064
rect 3187 4030 3188 4064
rect 3152 3996 3188 4030
rect 256 3905 257 3939
rect 291 3905 330 3939
rect 256 3870 330 3905
rect 2886 3947 2952 3985
rect 2886 3913 2902 3947
rect 2936 3913 2952 3947
rect 2886 3901 2952 3913
rect 3152 3962 3153 3996
rect 3187 3962 3188 3996
rect 3152 3928 3188 3962
rect 256 3836 257 3870
rect 291 3836 330 3870
rect 256 3801 330 3836
rect 256 3767 257 3801
rect 291 3767 330 3801
rect 256 3732 330 3767
rect 256 3698 257 3732
rect 291 3698 330 3732
rect 256 3663 330 3698
rect 256 3629 257 3663
rect 291 3629 330 3663
rect 256 3594 330 3629
rect 256 3560 257 3594
rect 291 3560 330 3594
rect 256 3525 330 3560
rect 256 3491 257 3525
rect 291 3491 330 3525
rect 256 3456 330 3491
rect 256 3422 257 3456
rect 291 3422 330 3456
rect 256 3387 330 3422
rect 256 3353 257 3387
rect 291 3353 330 3387
rect 256 3318 330 3353
rect 256 3284 257 3318
rect 291 3284 330 3318
rect 256 3249 330 3284
rect 256 3215 257 3249
rect 291 3215 330 3249
rect 256 3180 330 3215
rect 256 3146 257 3180
rect 291 3146 330 3180
rect 256 3111 330 3146
rect 256 3077 257 3111
rect 291 3077 330 3111
rect 256 3042 330 3077
rect 256 3008 257 3042
rect 291 3008 330 3042
rect 256 2973 330 3008
rect 256 2939 257 2973
rect 291 2939 330 2973
rect 256 2904 330 2939
rect 256 2870 257 2904
rect 291 2870 330 2904
rect 256 2835 330 2870
rect 256 2801 257 2835
rect 291 2801 330 2835
rect 256 2766 330 2801
rect 256 2732 257 2766
rect 291 2732 330 2766
rect 256 2697 330 2732
rect 256 2663 257 2697
rect 291 2663 330 2697
rect 256 2628 330 2663
rect 256 2594 257 2628
rect 291 2594 330 2628
rect 256 2559 330 2594
rect 256 2525 257 2559
rect 291 2525 330 2559
rect 256 2490 330 2525
rect 256 2456 257 2490
rect 291 2456 330 2490
rect 256 2421 330 2456
rect 256 2387 257 2421
rect 291 2387 330 2421
rect 256 2352 330 2387
rect 256 2318 257 2352
rect 291 2318 330 2352
rect 256 2283 330 2318
rect 256 2249 257 2283
rect 291 2249 330 2283
rect 256 2214 330 2249
rect 256 2180 257 2214
rect 291 2180 330 2214
rect 256 2145 330 2180
rect 256 2111 257 2145
rect 291 2111 330 2145
rect 256 2076 330 2111
rect 256 2042 257 2076
rect 291 2042 330 2076
rect 256 2007 330 2042
rect 256 1973 257 2007
rect 291 1973 330 2007
rect 256 1938 330 1973
rect 256 1904 257 1938
rect 291 1904 330 1938
rect 256 1869 330 1904
rect 256 1835 257 1869
rect 291 1835 330 1869
rect 256 1800 330 1835
rect 256 1766 257 1800
rect 291 1766 330 1800
rect 256 1731 330 1766
rect 256 1697 257 1731
rect 291 1697 330 1731
rect 256 1662 330 1697
rect 256 1628 257 1662
rect 291 1628 330 1662
rect 256 1593 330 1628
rect 256 1559 257 1593
rect 291 1559 330 1593
rect 256 1524 330 1559
rect 256 1490 257 1524
rect 291 1490 330 1524
rect 256 1456 330 1490
rect 256 1422 257 1456
rect 291 1422 330 1456
rect 256 1388 330 1422
rect 256 1354 257 1388
rect 291 1354 330 1388
rect 256 1320 330 1354
rect 256 1286 257 1320
rect 291 1286 330 1320
rect 256 1252 330 1286
rect 256 1218 257 1252
rect 291 1218 330 1252
rect 256 1184 330 1218
rect 256 1150 257 1184
rect 291 1150 330 1184
rect 256 1116 330 1150
rect 256 1082 257 1116
rect 291 1082 330 1116
rect 256 1048 330 1082
rect 256 1014 257 1048
rect 291 1014 330 1048
rect 256 980 330 1014
rect 256 946 257 980
rect 291 946 330 980
rect 256 912 330 946
rect 256 878 257 912
rect 291 878 330 912
rect 256 844 330 878
rect 256 810 257 844
rect 291 810 330 844
rect 256 776 330 810
rect 256 742 257 776
rect 291 742 330 776
rect 256 708 330 742
rect 256 674 257 708
rect 291 674 330 708
rect 256 640 330 674
rect 256 606 257 640
rect 291 606 330 640
rect 256 572 330 606
rect 3152 3894 3153 3928
rect 3187 3894 3188 3928
rect 3152 3860 3188 3894
rect 3152 3826 3153 3860
rect 3187 3826 3188 3860
rect 3152 3792 3188 3826
rect 3152 3758 3153 3792
rect 3187 3758 3188 3792
rect 3152 3724 3188 3758
rect 3152 3690 3153 3724
rect 3187 3690 3188 3724
rect 3152 3656 3188 3690
rect 3152 3622 3153 3656
rect 3187 3622 3188 3656
rect 3152 3588 3188 3622
rect 3152 3554 3153 3588
rect 3187 3554 3188 3588
rect 3152 3520 3188 3554
rect 3152 3486 3153 3520
rect 3187 3486 3188 3520
rect 3152 3452 3188 3486
rect 3152 3418 3153 3452
rect 3187 3418 3188 3452
rect 3152 3384 3188 3418
rect 3152 3350 3153 3384
rect 3187 3350 3188 3384
rect 3152 3316 3188 3350
rect 3152 3282 3153 3316
rect 3187 3282 3188 3316
rect 3152 3248 3188 3282
rect 3152 3214 3153 3248
rect 3187 3214 3188 3248
rect 3152 3180 3188 3214
rect 3152 3146 3153 3180
rect 3187 3146 3188 3180
rect 3152 3112 3188 3146
rect 3152 3078 3153 3112
rect 3187 3078 3188 3112
rect 3152 3044 3188 3078
rect 3152 3010 3153 3044
rect 3187 3010 3188 3044
rect 3152 2976 3188 3010
rect 3152 2942 3153 2976
rect 3187 2942 3188 2976
rect 3152 2908 3188 2942
rect 3152 2874 3153 2908
rect 3187 2874 3188 2908
rect 3152 2840 3188 2874
rect 3152 2806 3153 2840
rect 3187 2806 3188 2840
rect 3152 2772 3188 2806
rect 3152 2738 3153 2772
rect 3187 2738 3188 2772
rect 3152 2704 3188 2738
rect 3152 2670 3153 2704
rect 3187 2670 3188 2704
rect 3152 2636 3188 2670
rect 3152 2602 3153 2636
rect 3187 2602 3188 2636
rect 3152 2568 3188 2602
rect 3152 2534 3153 2568
rect 3187 2534 3188 2568
rect 3152 2500 3188 2534
rect 3152 2466 3153 2500
rect 3187 2466 3188 2500
rect 3152 2432 3188 2466
rect 3152 2398 3153 2432
rect 3187 2398 3188 2432
rect 3152 2364 3188 2398
rect 3152 2330 3153 2364
rect 3187 2330 3188 2364
rect 3152 2296 3188 2330
rect 3152 2262 3153 2296
rect 3187 2262 3188 2296
rect 3152 2228 3188 2262
rect 3152 2194 3153 2228
rect 3187 2194 3188 2228
rect 3152 2160 3188 2194
rect 3152 2126 3153 2160
rect 3187 2126 3188 2160
rect 3152 2092 3188 2126
rect 3152 2058 3153 2092
rect 3187 2058 3188 2092
rect 3152 2024 3188 2058
rect 3152 1990 3153 2024
rect 3187 1990 3188 2024
rect 3152 1956 3188 1990
rect 3152 1922 3153 1956
rect 3187 1922 3188 1956
rect 3152 1888 3188 1922
rect 3152 1854 3153 1888
rect 3187 1854 3188 1888
rect 3152 1820 3188 1854
rect 3152 1786 3153 1820
rect 3187 1786 3188 1820
rect 3152 1752 3188 1786
rect 3152 1718 3153 1752
rect 3187 1718 3188 1752
rect 3152 1684 3188 1718
rect 3152 1650 3153 1684
rect 3187 1650 3188 1684
rect 3152 1616 3188 1650
rect 3152 1582 3153 1616
rect 3187 1582 3188 1616
rect 3152 1548 3188 1582
rect 3152 1514 3153 1548
rect 3187 1514 3188 1548
rect 3152 1480 3188 1514
rect 3152 1446 3153 1480
rect 3187 1446 3188 1480
rect 3152 1412 3188 1446
rect 3152 1378 3153 1412
rect 3187 1378 3188 1412
rect 3152 1344 3188 1378
rect 3152 1310 3153 1344
rect 3187 1310 3188 1344
rect 3152 1276 3188 1310
rect 3152 1242 3153 1276
rect 3187 1242 3188 1276
rect 3152 1208 3188 1242
rect 3152 1174 3153 1208
rect 3187 1174 3188 1208
rect 3152 1140 3188 1174
rect 3152 1106 3153 1140
rect 3187 1106 3188 1140
rect 3152 1072 3188 1106
rect 3152 1038 3153 1072
rect 3187 1038 3188 1072
rect 3152 1004 3188 1038
rect 3152 970 3153 1004
rect 3187 970 3188 1004
rect 3152 936 3188 970
rect 3152 902 3153 936
rect 3187 902 3188 936
rect 3152 868 3188 902
rect 3152 834 3153 868
rect 3187 834 3188 868
rect 3152 800 3188 834
rect 3152 766 3153 800
rect 3187 766 3188 800
rect 3152 732 3188 766
rect 3152 698 3153 732
rect 3187 698 3188 732
rect 3152 664 3188 698
rect 3152 630 3153 664
rect 3187 630 3188 664
rect 3152 596 3188 630
rect 256 538 257 572
rect 291 538 330 572
rect 256 504 330 538
rect 2004 572 2070 578
rect 2004 538 2020 572
rect 2054 538 2070 572
rect 256 470 257 504
rect 291 470 330 504
rect 366 492 432 504
rect 366 476 382 492
rect 256 436 330 470
rect 416 476 432 492
rect 492 492 558 504
rect 492 476 508 492
rect 382 442 416 458
rect 542 476 558 492
rect 618 492 684 504
rect 618 476 634 492
rect 508 442 542 458
rect 668 476 684 492
rect 744 492 810 504
rect 744 476 760 492
rect 634 442 668 458
rect 794 476 810 492
rect 870 492 936 504
rect 870 476 886 492
rect 760 442 794 458
rect 920 476 936 492
rect 996 492 1062 504
rect 996 476 1012 492
rect 886 442 920 458
rect 1046 476 1062 492
rect 1122 492 1188 504
rect 1122 476 1138 492
rect 1012 442 1046 458
rect 1172 476 1188 492
rect 1248 492 1314 504
rect 1248 476 1264 492
rect 1138 442 1172 458
rect 1298 476 1314 492
rect 1374 492 1440 504
rect 1374 476 1390 492
rect 1264 442 1298 458
rect 1424 476 1440 492
rect 1500 492 1566 504
rect 1500 476 1516 492
rect 1390 442 1424 458
rect 1550 476 1566 492
rect 1626 492 1692 504
rect 1626 476 1642 492
rect 1516 442 1550 458
rect 1676 476 1692 492
rect 1752 492 1818 504
rect 1752 476 1768 492
rect 1642 442 1676 458
rect 1802 476 1818 492
rect 1878 492 1944 504
rect 1878 476 1894 492
rect 1768 442 1802 458
rect 1928 476 1944 492
rect 2004 500 2070 538
rect 2004 476 2020 500
rect 2054 476 2070 500
rect 2130 572 2196 578
rect 2130 538 2146 572
rect 2180 538 2196 572
rect 2130 500 2196 538
rect 2130 476 2146 500
rect 2180 476 2196 500
rect 2256 572 2322 578
rect 2256 538 2272 572
rect 2306 538 2322 572
rect 2256 500 2322 538
rect 2256 476 2272 500
rect 2306 476 2322 500
rect 2382 572 2448 578
rect 2382 538 2398 572
rect 2432 538 2448 572
rect 2382 500 2448 538
rect 3152 562 3153 596
rect 3187 562 3188 596
rect 3152 528 3188 562
rect 2382 476 2398 500
rect 2432 476 2448 500
rect 2508 492 2574 498
rect 1894 442 1928 458
rect 2508 458 2524 492
rect 2558 458 2574 492
rect 256 402 257 436
rect 291 402 330 436
rect 256 292 330 402
rect 366 420 432 442
rect 366 374 382 420
rect 416 374 432 420
rect 492 420 558 442
rect 492 374 508 420
rect 542 374 558 420
rect 618 420 684 442
rect 618 374 634 420
rect 668 374 684 420
rect 744 420 810 442
rect 744 374 760 420
rect 794 374 810 420
rect 870 420 936 442
rect 870 374 886 420
rect 920 374 936 420
rect 996 420 1062 442
rect 996 374 1012 420
rect 1046 374 1062 420
rect 1122 420 1188 442
rect 1122 374 1138 420
rect 1172 374 1188 420
rect 1248 420 1314 442
rect 1248 374 1264 420
rect 1298 374 1314 420
rect 1374 420 1440 442
rect 1374 374 1390 420
rect 1424 374 1440 420
rect 1500 420 1566 442
rect 1500 374 1516 420
rect 1550 374 1566 420
rect 1626 420 1692 442
rect 1626 374 1642 420
rect 1676 374 1692 420
rect 1752 420 1818 442
rect 1752 374 1768 420
rect 1802 374 1818 420
rect 1878 420 1944 442
rect 1878 374 1894 420
rect 1928 374 1944 420
rect 2004 408 2070 442
rect 2004 374 2020 408
rect 2054 374 2070 408
rect 2130 408 2196 442
rect 2130 374 2146 408
rect 2180 374 2196 408
rect 2256 408 2322 442
rect 2256 374 2272 408
rect 2306 374 2322 408
rect 2382 408 2448 442
rect 2382 374 2398 408
rect 2432 374 2448 408
rect 2508 420 2574 458
rect 2508 374 2524 420
rect 2558 374 2574 420
rect 2634 492 2700 498
rect 2634 458 2650 492
rect 2684 458 2700 492
rect 2634 420 2700 458
rect 2634 374 2650 420
rect 2684 374 2700 420
rect 2760 492 2826 498
rect 2760 458 2776 492
rect 2810 458 2826 492
rect 2886 492 2952 504
rect 2886 476 2902 492
rect 2760 420 2826 458
rect 2936 476 2952 492
rect 3012 492 3078 504
rect 3012 476 3028 492
rect 2902 442 2936 458
rect 3062 476 3078 492
rect 3152 494 3153 528
rect 3187 494 3188 528
rect 3028 442 3062 458
rect 3152 460 3188 494
rect 2760 374 2776 420
rect 2810 374 2826 420
rect 2886 420 2952 442
rect 2886 374 2902 420
rect 2936 374 2952 420
rect 3012 420 3078 442
rect 3012 374 3028 420
rect 3062 374 3078 420
rect 3152 426 3153 460
rect 3187 426 3188 460
rect 3152 392 3188 426
rect 3152 358 3153 392
rect 3187 358 3188 392
rect 3152 324 3188 358
rect 3152 292 3153 324
rect 256 291 3153 292
rect 256 257 290 291
rect 324 257 358 291
rect 392 257 426 291
rect 460 257 494 291
rect 528 257 562 291
rect 596 257 630 291
rect 664 257 698 291
rect 732 257 766 291
rect 800 257 834 291
rect 868 257 902 291
rect 936 257 970 291
rect 1004 257 1038 291
rect 1072 257 1106 291
rect 1140 257 1174 291
rect 1208 257 1242 291
rect 1276 257 1310 291
rect 1344 257 1378 291
rect 1412 257 1446 291
rect 1480 257 1514 291
rect 1548 257 1582 291
rect 1616 257 1650 291
rect 1684 257 1718 291
rect 1752 257 1786 291
rect 1820 257 1854 291
rect 1888 257 1922 291
rect 1956 257 1990 291
rect 2024 257 2058 291
rect 2092 257 2126 291
rect 2160 257 2194 291
rect 2228 257 2262 291
rect 2296 257 2330 291
rect 2364 257 2398 291
rect 2432 257 2466 291
rect 2500 257 2534 291
rect 2568 257 2602 291
rect 2636 257 2670 291
rect 2704 257 2738 291
rect 2772 257 2806 291
rect 2840 257 2874 291
rect 2908 257 2942 291
rect 2976 257 3010 291
rect 3044 257 3078 291
rect 3112 290 3153 291
rect 3187 290 3188 324
rect 3112 257 3188 290
rect 256 142 3188 257
rect 3341 862 3377 899
rect 3341 828 3342 862
rect 3376 828 3377 862
rect 3341 815 3377 828
rect 3341 752 3342 815
rect 3376 752 3377 815
rect 3341 747 3377 752
rect 3341 713 3342 747
rect 3376 713 3377 747
rect 3341 710 3377 713
rect 3341 645 3342 710
rect 3376 645 3377 710
rect 3341 634 3377 645
rect 3341 577 3342 634
rect 3376 577 3377 634
rect 3341 558 3377 577
rect 3341 509 3342 558
rect 3376 509 3377 558
rect 3341 482 3377 509
rect 3341 441 3342 482
rect 3376 441 3377 482
rect 3341 407 3377 441
rect 3341 372 3342 407
rect 3376 372 3377 407
rect 3341 339 3377 372
rect 3341 296 3342 339
rect 3376 296 3377 339
rect 3341 271 3377 296
rect 3341 220 3342 271
rect 3376 220 3377 271
rect 3341 203 3377 220
rect 3341 144 3342 203
rect 3376 144 3377 203
rect 3341 135 3377 144
rect 3341 103 3342 135
rect 742 102 3342 103
rect 742 70 887 102
rect 776 69 887 70
rect 777 68 887 69
rect 921 68 955 102
rect 989 68 1023 102
rect 1057 68 1091 102
rect 1125 68 1159 102
rect 1193 68 1227 102
rect 1261 68 1295 102
rect 1329 68 1363 102
rect 1397 68 1431 102
rect 1465 68 1499 102
rect 1533 68 1567 102
rect 1601 68 1635 102
rect 1669 68 1703 102
rect 1737 68 1771 102
rect 1805 68 1839 102
rect 1873 68 1907 102
rect 1941 68 1975 102
rect 2009 68 2043 102
rect 2077 68 2111 102
rect 2145 68 2179 102
rect 2213 68 2247 102
rect 2281 68 2315 102
rect 2349 68 2383 102
rect 2417 68 2451 102
rect 2485 68 2519 102
rect 2553 68 2587 102
rect 2621 68 2655 102
rect 2689 68 2723 102
rect 2757 68 2791 102
rect 2825 68 2859 102
rect 2893 68 2927 102
rect 2961 68 2995 102
rect 3029 68 3063 102
rect 3097 68 3131 102
rect 3165 68 3199 102
rect 3233 68 3267 102
rect 3301 68 3342 102
rect 3376 78 3377 135
rect 3376 68 3640 78
rect 777 67 3640 68
rect 742 35 743 36
rect 777 35 778 67
rect 3341 44 3640 67
rect 742 1 778 35
rect 742 -18 743 1
rect 777 -33 778 1
rect 776 -52 778 -33
rect 3604 8 3640 44
rect 3604 -28 3605 8
rect 3639 -28 3640 8
rect 742 -67 778 -52
rect 742 -101 743 -67
rect 777 -101 778 -67
rect 742 -107 778 -101
rect 776 -135 778 -107
rect 742 -169 743 -141
rect 777 -169 778 -135
rect 742 -196 778 -169
rect 776 -203 778 -196
rect 742 -237 743 -230
rect 777 -237 778 -203
rect 2458 -128 2492 -90
rect 2914 -116 2948 -78
rect 3370 -128 3404 -90
rect 2458 -200 2492 -162
rect 3370 -200 3404 -162
rect 742 -271 778 -237
rect 742 -305 743 -271
rect 777 -305 778 -271
rect 2526 -240 2547 -206
rect 2581 -240 2619 -206
rect 2653 -240 2691 -206
rect 2725 -240 2763 -206
rect 2797 -240 2835 -206
rect 2869 -240 2880 -206
rect 3604 -60 3640 -28
rect 3604 -101 3605 -60
rect 3639 -101 3640 -60
rect 3604 -128 3640 -101
rect 3604 -174 3605 -128
rect 3639 -174 3640 -128
rect 3604 -196 3640 -174
rect 2526 -280 2880 -240
rect 3604 -247 3605 -196
rect 3639 -247 3640 -196
rect 3604 -264 3640 -247
rect 742 -339 778 -305
rect 905 -314 943 -280
rect 977 -314 1011 -280
rect 1045 -314 1079 -280
rect 1113 -314 1147 -280
rect 1181 -314 1215 -280
rect 1249 -314 1283 -280
rect 1317 -314 1351 -280
rect 1385 -314 1419 -280
rect 1453 -314 1487 -280
rect 1521 -314 1555 -280
rect 1589 -314 1623 -280
rect 1657 -314 1691 -280
rect 1725 -314 1759 -280
rect 1793 -314 1827 -280
rect 1861 -314 1895 -280
rect 1929 -314 1963 -280
rect 2065 -314 2069 -280
rect 2137 -314 2153 -280
rect 2187 -314 2287 -280
rect 2321 -314 2337 -280
rect 2371 -314 2409 -280
rect 2503 -314 2519 -280
rect 2553 -314 2603 -280
rect 2637 -314 2687 -280
rect 2721 -314 2770 -280
rect 2804 -314 2853 -280
rect 2887 -314 2903 -280
rect 2959 -314 2975 -280
rect 3032 -314 3059 -280
rect 3104 -314 3142 -280
rect 3177 -314 3214 -280
rect 3260 -314 3309 -280
rect 3343 -314 3359 -280
rect 742 -373 743 -339
rect 777 -373 778 -339
rect 3604 -320 3605 -264
rect 3639 -320 3640 -264
rect 3604 -332 3640 -320
rect 3604 -364 3605 -332
rect 742 -381 778 -373
rect 776 -407 778 -381
rect 742 -441 743 -415
rect 777 -441 778 -407
rect 742 -462 778 -441
rect 776 -475 778 -462
rect 742 -509 743 -496
rect 777 -509 778 -475
rect 742 -543 778 -509
rect 777 -577 778 -543
rect 742 -623 778 -577
rect 776 -628 778 -623
rect 1680 -365 3605 -364
rect 1680 -371 1714 -365
rect 1680 -405 1681 -371
rect 1748 -399 1756 -365
rect 1790 -399 1830 -365
rect 1895 -399 1904 -365
rect 1963 -399 1978 -365
rect 2031 -399 2052 -365
rect 2099 -399 2126 -365
rect 2167 -399 2200 -365
rect 2235 -399 2269 -365
rect 2308 -399 2337 -365
rect 2382 -399 2405 -365
rect 2456 -399 2473 -365
rect 2530 -399 2541 -365
rect 2604 -399 2609 -365
rect 2643 -399 2644 -365
rect 2711 -399 2718 -365
rect 2779 -399 2792 -365
rect 2847 -399 2866 -365
rect 2915 -399 2940 -365
rect 2983 -399 3014 -365
rect 3051 -399 3085 -365
rect 3122 -399 3153 -365
rect 3196 -399 3221 -365
rect 3270 -399 3289 -365
rect 3344 -399 3357 -365
rect 3418 -399 3425 -365
rect 3492 -399 3493 -365
rect 3527 -399 3533 -365
rect 3567 -393 3605 -365
rect 3639 -393 3640 -332
rect 3567 -399 3640 -393
rect 1715 -400 3640 -399
rect 1715 -405 1716 -400
rect 1680 -460 1716 -405
rect 1680 -498 1681 -460
rect 1715 -498 1716 -460
rect 1680 -528 1716 -498
rect 1680 -591 1681 -528
rect 1715 -591 1716 -528
rect 1680 -596 1716 -591
rect 1680 -628 1681 -596
rect 776 -629 1681 -628
rect 742 -663 776 -657
rect 810 -663 844 -629
rect 878 -663 912 -629
rect 946 -663 980 -629
rect 1014 -663 1048 -629
rect 1082 -663 1116 -629
rect 1150 -663 1184 -629
rect 1218 -663 1252 -629
rect 1286 -663 1320 -629
rect 1354 -663 1388 -629
rect 1422 -663 1456 -629
rect 1490 -663 1524 -629
rect 1558 -663 1592 -629
rect 1626 -630 1681 -629
rect 1715 -630 1716 -596
rect 1626 -663 1716 -630
rect 742 -664 1716 -663
rect 2148 -554 3498 -553
rect 2148 -560 2221 -554
rect 2148 -621 2149 -560
rect 2183 -588 2221 -560
rect 2255 -588 2274 -554
rect 2328 -588 2342 -554
rect 2401 -588 2410 -554
rect 2474 -588 2478 -554
rect 2512 -588 2513 -554
rect 2580 -588 2586 -554
rect 2648 -588 2659 -554
rect 2716 -588 2732 -554
rect 2784 -588 2805 -554
rect 2852 -588 2878 -554
rect 2920 -588 2951 -554
rect 2988 -588 3022 -554
rect 3058 -588 3090 -554
rect 3131 -588 3158 -554
rect 3204 -588 3226 -554
rect 3277 -588 3294 -554
rect 3351 -588 3362 -554
rect 3425 -588 3430 -554
rect 3464 -560 3498 -554
rect 2183 -589 3463 -588
rect 2183 -621 2184 -589
rect 2148 -645 2184 -621
rect 3462 -594 3463 -589
rect 3497 -594 3498 -560
rect 3462 -622 3498 -594
rect 2148 -689 2149 -645
rect 2183 -689 2184 -645
rect 2337 -673 2357 -639
rect 2405 -673 2421 -639
rect 2489 -673 2527 -639
rect 2577 -673 2637 -639
rect 2671 -673 2759 -639
rect 2793 -673 2853 -639
rect 2887 -673 2903 -639
rect 2959 -673 2975 -639
rect 3009 -673 3047 -639
rect 3103 -673 3191 -639
rect 3225 -673 3285 -639
rect 3319 -673 3335 -639
rect 2148 -723 2184 -689
rect 2148 -765 2149 -723
rect 2183 -765 2184 -723
rect 2148 -791 2184 -765
rect 2148 -851 2149 -791
rect 2183 -851 2184 -791
rect 2266 -791 2300 -753
rect 2698 -791 2732 -753
rect 2148 -859 2184 -851
rect 2148 -893 2149 -859
rect 2183 -893 2184 -859
rect 2148 -903 2184 -893
rect 2148 -937 2149 -903
rect 2183 -937 2184 -903
rect 3130 -791 3164 -753
rect 2482 -890 2516 -852
rect 3232 -837 3278 -673
rect 3462 -680 3463 -622
rect 3497 -680 3498 -622
rect 3462 -690 3498 -680
rect 3462 -724 3463 -690
rect 3497 -724 3498 -690
rect 3462 -732 3498 -724
rect 3462 -792 3463 -732
rect 3497 -792 3498 -732
rect 2914 -890 2948 -852
rect 3346 -890 3380 -852
rect 3462 -826 3498 -792
rect 3462 -860 3463 -826
rect 3497 -860 3498 -826
rect 3462 -894 3498 -860
rect 2148 -989 2184 -937
rect 2148 -1023 2149 -989
rect 2183 -994 2184 -989
rect 3462 -928 3463 -894
rect 3497 -928 3498 -894
rect 3462 -962 3498 -928
rect 3462 -994 3463 -962
rect 2183 -995 3463 -994
rect 2148 -1029 2182 -1023
rect 2216 -1029 2221 -995
rect 2284 -1029 2294 -995
rect 2352 -1029 2367 -995
rect 2420 -1029 2440 -995
rect 2488 -1029 2513 -995
rect 2556 -1029 2586 -995
rect 2624 -1029 2658 -995
rect 2693 -1029 2726 -995
rect 2766 -1029 2794 -995
rect 2839 -1029 2862 -995
rect 2912 -1029 2930 -995
rect 2985 -1029 2998 -995
rect 3058 -1029 3066 -995
rect 3131 -1029 3134 -995
rect 3168 -1029 3170 -995
rect 3236 -1029 3243 -995
rect 3304 -1029 3317 -995
rect 3372 -1029 3391 -995
rect 3425 -996 3463 -995
rect 3497 -996 3498 -962
rect 3425 -1029 3498 -996
rect 2148 -1030 3498 -1029
<< viali >>
rect 172 27835 199 27869
rect 199 27835 206 27869
rect 244 27835 267 27869
rect 267 27835 278 27869
rect 1673 27835 1695 27869
rect 1695 27835 1707 27869
rect 1745 27835 1763 27869
rect 1763 27835 1779 27869
rect 1817 27835 1831 27869
rect 1831 27835 1851 27869
rect 1889 27835 1899 27869
rect 1899 27835 1923 27869
rect 68 27768 102 27785
rect 68 27751 102 27768
rect 68 27700 102 27711
rect 68 27677 102 27700
rect 68 27632 102 27637
rect 68 27603 102 27632
rect 68 27530 102 27563
rect 68 27529 102 27530
rect 68 27462 102 27489
rect 68 27455 102 27462
rect 68 27394 102 27415
rect 68 27381 102 27394
rect 68 27326 102 27342
rect 68 27308 102 27326
rect 68 27258 102 27269
rect 68 27235 102 27258
rect 68 27190 102 27196
rect 68 27162 102 27190
rect 68 27122 102 27123
rect 68 27089 102 27122
rect 68 27020 102 27050
rect 68 27016 102 27020
rect 68 26952 102 26977
rect 68 26943 102 26952
rect 68 26884 102 26904
rect 68 26870 102 26884
rect 68 26816 102 26831
rect 68 26797 102 26816
rect 68 26748 102 26758
rect 68 26724 102 26748
rect 68 26680 102 26685
rect 68 26651 102 26680
rect 68 26578 102 26612
rect 68 26510 102 26539
rect 68 26505 102 26510
rect 68 26442 102 26466
rect 68 26432 102 26442
rect 68 26374 102 26393
rect 68 26359 102 26374
rect 68 26306 102 26320
rect 68 26286 102 26306
rect 68 26238 102 26247
rect 68 26213 102 26238
rect 68 26170 102 26174
rect 68 26140 102 26170
rect 68 26068 102 26101
rect 68 26067 102 26068
rect 68 26000 102 26028
rect 68 25994 102 26000
rect 68 25932 102 25955
rect 68 25921 102 25932
rect 68 25864 102 25882
rect 68 25848 102 25864
rect 68 25796 102 25809
rect 68 25775 102 25796
rect 68 25702 102 25736
rect 382 27529 416 27551
rect 382 27517 416 27529
rect 508 27529 542 27551
rect 508 27517 542 27529
rect 634 27529 668 27551
rect 634 27517 668 27529
rect 760 27529 794 27551
rect 760 27517 794 27529
rect 886 27529 920 27551
rect 886 27517 920 27529
rect 1012 27529 1046 27551
rect 1012 27517 1046 27529
rect 1138 27529 1172 27551
rect 1138 27517 1172 27529
rect 1264 27529 1298 27551
rect 1264 27517 1298 27529
rect 1390 27529 1424 27551
rect 1390 27517 1424 27529
rect 1516 27529 1550 27551
rect 1516 27517 1550 27529
rect 1642 27529 1676 27551
rect 1642 27517 1676 27529
rect 1768 27529 1802 27551
rect 1768 27517 1802 27529
rect 1894 27529 1928 27551
rect 1894 27517 1928 27529
rect 2020 27529 2054 27551
rect 2020 27517 2054 27529
rect 382 27445 416 27479
rect 508 27445 542 27479
rect 634 27445 668 27479
rect 760 27445 794 27479
rect 886 27445 920 27479
rect 1012 27445 1046 27479
rect 1138 27445 1172 27479
rect 1264 27445 1298 27479
rect 1390 27445 1424 27479
rect 1516 27445 1550 27479
rect 1642 27445 1676 27479
rect 1768 27445 1802 27479
rect 1894 27445 1928 27479
rect 2020 27445 2054 27479
rect 382 23828 416 23862
rect 508 23828 542 23862
rect 634 23828 668 23862
rect 760 23828 794 23862
rect 886 23828 920 23862
rect 1012 23828 1046 23862
rect 1138 23828 1172 23862
rect 1264 23828 1298 23862
rect 1390 23828 1424 23862
rect 1516 23828 1550 23862
rect 1642 23828 1676 23862
rect 1768 23828 1802 23862
rect 1894 23828 1928 23862
rect 2020 23828 2054 23862
rect 382 23778 416 23790
rect 382 23756 416 23778
rect 508 23778 542 23790
rect 508 23756 542 23778
rect 634 23778 668 23790
rect 634 23756 668 23778
rect 760 23778 794 23790
rect 760 23756 794 23778
rect 886 23778 920 23790
rect 886 23756 920 23778
rect 1012 23778 1046 23790
rect 1012 23756 1046 23778
rect 1138 23778 1172 23790
rect 1138 23756 1172 23778
rect 1264 23778 1298 23790
rect 1264 23756 1298 23778
rect 1390 23778 1424 23790
rect 1390 23756 1424 23778
rect 1516 23778 1550 23790
rect 1516 23756 1550 23778
rect 1642 23778 1676 23790
rect 1642 23756 1676 23778
rect 1768 23778 1802 23790
rect 1768 23756 1802 23778
rect 1894 23778 1928 23790
rect 1894 23756 1928 23778
rect 2020 23778 2054 23790
rect 2020 23756 2054 23778
rect 382 23634 416 23656
rect 382 23622 416 23634
rect 508 23634 542 23656
rect 508 23622 542 23634
rect 634 23634 668 23656
rect 634 23622 668 23634
rect 760 23634 794 23656
rect 760 23622 794 23634
rect 886 23634 920 23656
rect 886 23622 920 23634
rect 1012 23634 1046 23656
rect 1012 23622 1046 23634
rect 1138 23634 1172 23656
rect 1138 23622 1172 23634
rect 1264 23634 1298 23656
rect 1264 23622 1298 23634
rect 1390 23634 1424 23656
rect 1390 23622 1424 23634
rect 1516 23634 1550 23656
rect 1516 23622 1550 23634
rect 1642 23634 1676 23656
rect 1642 23622 1676 23634
rect 1768 23634 1802 23656
rect 1768 23622 1802 23634
rect 1894 23634 1928 23656
rect 1894 23622 1928 23634
rect 2020 23634 2054 23656
rect 2020 23622 2054 23634
rect 382 23550 416 23584
rect 508 23550 542 23584
rect 634 23550 668 23584
rect 760 23550 794 23584
rect 886 23550 920 23584
rect 1012 23550 1046 23584
rect 1138 23550 1172 23584
rect 1264 23550 1298 23584
rect 1390 23550 1424 23584
rect 1516 23550 1550 23584
rect 1642 23550 1676 23584
rect 1768 23550 1802 23584
rect 1894 23550 1928 23584
rect 2020 23550 2054 23584
rect 1390 22357 1424 22391
rect 1642 22357 1676 22391
rect 1894 22357 1928 22391
rect 1390 22307 1424 22319
rect 1390 22285 1424 22307
rect 1642 22307 1676 22319
rect 1642 22285 1676 22307
rect 1894 22307 1928 22319
rect 1894 22285 1928 22307
rect 382 19933 416 19967
rect 508 19933 542 19967
rect 634 19933 668 19967
rect 760 19933 794 19967
rect 886 19933 920 19967
rect 1012 19933 1046 19967
rect 1138 19933 1172 19967
rect 1264 19933 1298 19967
rect 1516 19933 1550 19967
rect 1768 19933 1802 19967
rect 2020 19933 2054 19967
rect 382 19883 416 19895
rect 382 19861 416 19883
rect 508 19883 542 19895
rect 508 19861 542 19883
rect 634 19883 668 19895
rect 634 19861 668 19883
rect 760 19883 794 19895
rect 760 19861 794 19883
rect 886 19883 920 19895
rect 886 19861 920 19883
rect 1012 19883 1046 19895
rect 1012 19861 1046 19883
rect 1138 19883 1172 19895
rect 1138 19861 1172 19883
rect 1264 19883 1298 19895
rect 1264 19861 1298 19883
rect 1516 19883 1550 19895
rect 1516 19861 1550 19883
rect 1768 19883 1802 19895
rect 1768 19861 1802 19883
rect 2020 19883 2054 19895
rect 2020 19861 2054 19883
rect 382 19739 416 19761
rect 382 19727 416 19739
rect 508 19739 542 19761
rect 508 19727 542 19739
rect 634 19739 668 19761
rect 634 19727 668 19739
rect 760 19739 794 19761
rect 760 19727 794 19739
rect 886 19739 920 19761
rect 886 19727 920 19739
rect 1012 19739 1046 19761
rect 1012 19727 1046 19739
rect 1138 19739 1172 19761
rect 1138 19727 1172 19739
rect 1264 19739 1298 19761
rect 1264 19727 1298 19739
rect 1390 19739 1424 19761
rect 1390 19727 1424 19739
rect 1516 19739 1550 19761
rect 1516 19727 1550 19739
rect 1642 19739 1676 19761
rect 1642 19727 1676 19739
rect 1768 19739 1802 19761
rect 1768 19727 1802 19739
rect 1894 19739 1928 19761
rect 1894 19727 1928 19739
rect 2020 19739 2054 19761
rect 2020 19727 2054 19739
rect 382 19655 416 19689
rect 508 19655 542 19689
rect 634 19655 668 19689
rect 760 19655 794 19689
rect 886 19655 920 19689
rect 1012 19655 1046 19689
rect 1138 19655 1172 19689
rect 1264 19655 1298 19689
rect 1390 19655 1424 19689
rect 1516 19655 1550 19689
rect 1642 19655 1676 19689
rect 1768 19655 1802 19689
rect 1894 19655 1928 19689
rect 2020 19655 2054 19689
rect 382 16038 416 16072
rect 508 16038 542 16072
rect 634 16038 668 16072
rect 760 16038 794 16072
rect 886 16038 920 16072
rect 1012 16038 1046 16072
rect 1138 16038 1172 16072
rect 1264 16038 1298 16072
rect 1390 16038 1424 16072
rect 1516 16038 1550 16072
rect 1642 16038 1676 16072
rect 1768 16038 1802 16072
rect 1894 16038 1928 16072
rect 2020 16038 2054 16072
rect 382 15988 416 16000
rect 382 15966 416 15988
rect 508 15988 542 16000
rect 508 15966 542 15988
rect 634 15988 668 16000
rect 634 15966 668 15988
rect 760 15988 794 16000
rect 760 15966 794 15988
rect 886 15988 920 16000
rect 886 15966 920 15988
rect 1012 15988 1046 16000
rect 1012 15966 1046 15988
rect 1138 15988 1172 16000
rect 1138 15966 1172 15988
rect 1264 15988 1298 16000
rect 1264 15966 1298 15988
rect 1390 15988 1424 16000
rect 1390 15966 1424 15988
rect 1516 15988 1550 16000
rect 1516 15966 1550 15988
rect 1642 15988 1676 16000
rect 1642 15966 1676 15988
rect 1768 15988 1802 16000
rect 1768 15966 1802 15988
rect 1894 15988 1928 16000
rect 1894 15966 1928 15988
rect 2020 15988 2054 16000
rect 2020 15966 2054 15988
rect 382 15844 416 15866
rect 382 15832 416 15844
rect 508 15844 542 15866
rect 508 15832 542 15844
rect 634 15844 668 15866
rect 634 15832 668 15844
rect 760 15844 794 15866
rect 760 15832 794 15844
rect 886 15844 920 15866
rect 886 15832 920 15844
rect 1012 15844 1046 15866
rect 1012 15832 1046 15844
rect 1138 15844 1172 15866
rect 1138 15832 1172 15844
rect 1264 15844 1298 15866
rect 1264 15832 1298 15844
rect 1390 15844 1424 15866
rect 1390 15832 1424 15844
rect 1516 15844 1550 15866
rect 1516 15832 1550 15844
rect 1642 15844 1676 15866
rect 1642 15832 1676 15844
rect 1768 15844 1802 15866
rect 1768 15832 1802 15844
rect 1894 15844 1928 15866
rect 1894 15832 1928 15844
rect 2020 15844 2054 15866
rect 2020 15832 2054 15844
rect 382 15760 416 15794
rect 508 15760 542 15794
rect 634 15760 668 15794
rect 760 15760 794 15794
rect 886 15760 920 15794
rect 1012 15760 1046 15794
rect 1138 15760 1172 15794
rect 1264 15760 1298 15794
rect 1390 15760 1424 15794
rect 1516 15760 1550 15794
rect 1642 15760 1676 15794
rect 1768 15760 1802 15794
rect 1894 15760 1928 15794
rect 2020 15760 2054 15794
rect 382 12143 416 12177
rect 508 12143 542 12177
rect 634 12143 668 12177
rect 760 12143 794 12177
rect 886 12143 920 12177
rect 1012 12143 1046 12177
rect 1138 12143 1172 12177
rect 1264 12143 1298 12177
rect 1390 12143 1424 12177
rect 1516 12143 1550 12177
rect 1642 12143 1676 12177
rect 1768 12143 1802 12177
rect 1894 12143 1928 12177
rect 2020 12143 2054 12177
rect 382 12093 416 12105
rect 382 12071 416 12093
rect 508 12093 542 12105
rect 508 12071 542 12093
rect 634 12093 668 12105
rect 634 12071 668 12093
rect 760 12093 794 12105
rect 760 12071 794 12093
rect 886 12093 920 12105
rect 886 12071 920 12093
rect 1012 12093 1046 12105
rect 1012 12071 1046 12093
rect 1138 12093 1172 12105
rect 1138 12071 1172 12093
rect 1264 12093 1298 12105
rect 1264 12071 1298 12093
rect 1390 12093 1424 12105
rect 1390 12071 1424 12093
rect 1516 12093 1550 12105
rect 1516 12071 1550 12093
rect 1642 12093 1676 12105
rect 1642 12071 1676 12093
rect 1768 12093 1802 12105
rect 1768 12071 1802 12093
rect 1894 12093 1928 12105
rect 1894 12071 1928 12093
rect 2020 12093 2054 12105
rect 2020 12071 2054 12093
rect 382 11949 416 11971
rect 382 11937 416 11949
rect 508 11949 542 11971
rect 508 11937 542 11949
rect 634 11949 668 11971
rect 634 11937 668 11949
rect 760 11949 794 11971
rect 760 11937 794 11949
rect 886 11949 920 11971
rect 886 11937 920 11949
rect 1012 11949 1046 11971
rect 1012 11937 1046 11949
rect 1138 11949 1172 11971
rect 1138 11937 1172 11949
rect 1264 11949 1298 11971
rect 1264 11937 1298 11949
rect 1390 11949 1424 11971
rect 1390 11937 1424 11949
rect 1516 11949 1550 11971
rect 1516 11937 1550 11949
rect 1642 11949 1676 11971
rect 1642 11937 1676 11949
rect 1768 11949 1802 11971
rect 1768 11937 1802 11949
rect 1894 11949 1928 11971
rect 1894 11937 1928 11949
rect 2020 11949 2054 11971
rect 2020 11937 2054 11949
rect 382 11865 416 11899
rect 508 11865 542 11899
rect 634 11865 668 11899
rect 760 11865 794 11899
rect 886 11865 920 11899
rect 1012 11865 1046 11899
rect 1138 11865 1172 11899
rect 1264 11865 1298 11899
rect 1390 11865 1424 11899
rect 1516 11865 1550 11899
rect 1642 11865 1676 11899
rect 1768 11865 1802 11899
rect 1894 11865 1928 11899
rect 2020 11865 2054 11899
rect 382 8248 416 8282
rect 508 8248 542 8282
rect 634 8248 668 8282
rect 760 8248 794 8282
rect 886 8248 920 8282
rect 1012 8248 1046 8282
rect 1138 8248 1172 8282
rect 1264 8248 1298 8282
rect 1390 8248 1424 8282
rect 1516 8248 1550 8282
rect 1642 8248 1676 8282
rect 1768 8248 1802 8282
rect 1894 8248 1928 8282
rect 382 8198 416 8210
rect 382 8176 416 8198
rect 508 8198 542 8210
rect 508 8176 542 8198
rect 634 8198 668 8210
rect 634 8176 668 8198
rect 760 8198 794 8210
rect 760 8176 794 8198
rect 886 8198 920 8210
rect 886 8176 920 8198
rect 1012 8198 1046 8210
rect 1012 8176 1046 8198
rect 1138 8198 1172 8210
rect 1138 8176 1172 8198
rect 1264 8198 1298 8210
rect 1264 8176 1298 8198
rect 1390 8198 1424 8210
rect 1390 8176 1424 8198
rect 1516 8198 1550 8210
rect 1516 8176 1550 8198
rect 1642 8198 1676 8210
rect 1642 8176 1676 8198
rect 1768 8198 1802 8210
rect 1768 8176 1802 8198
rect 1894 8198 1928 8210
rect 1894 8176 1928 8198
rect 382 8054 416 8076
rect 382 8042 416 8054
rect 508 8054 542 8076
rect 508 8042 542 8054
rect 634 8054 668 8076
rect 634 8042 668 8054
rect 760 8054 794 8076
rect 760 8042 794 8054
rect 886 8054 920 8076
rect 886 8042 920 8054
rect 1012 8054 1046 8076
rect 1012 8042 1046 8054
rect 1138 8054 1172 8076
rect 1138 8042 1172 8054
rect 1264 8054 1298 8076
rect 1264 8042 1298 8054
rect 1390 8054 1424 8076
rect 1390 8042 1424 8054
rect 1516 8054 1550 8076
rect 1516 8042 1550 8054
rect 1642 8054 1676 8076
rect 1642 8042 1676 8054
rect 382 7970 416 8004
rect 508 7970 542 8004
rect 634 7970 668 8004
rect 760 7970 794 8004
rect 886 7970 920 8004
rect 1012 7970 1046 8004
rect 1138 7970 1172 8004
rect 1264 7970 1298 8004
rect 1390 7970 1424 8004
rect 1516 7970 1550 8004
rect 1642 7970 1676 8004
rect 1894 7954 1928 7988
rect 1894 7882 1928 7916
rect 231 6732 265 6759
rect 231 6725 265 6732
rect 231 6660 265 6685
rect 231 6651 265 6660
rect 231 6589 265 6611
rect 231 6577 265 6589
rect 231 6518 265 6537
rect 231 6503 265 6518
rect 231 6447 265 6463
rect 231 6429 265 6447
rect 231 6376 265 6389
rect 231 6355 265 6376
rect 231 6305 265 6315
rect 231 6281 265 6305
rect 231 6234 265 6241
rect 231 6207 265 6234
rect 231 6163 265 6167
rect 231 6133 265 6163
rect 231 6092 265 6094
rect 231 6060 265 6092
rect 231 5987 265 6021
rect 231 5914 265 5948
rect 231 5842 265 5875
rect 231 5841 265 5842
rect 231 5768 265 5802
rect 231 5706 265 5729
rect 231 5695 253 5706
rect 253 5695 265 5706
rect 231 5638 265 5656
rect 231 5622 253 5638
rect 253 5622 265 5638
rect 231 5570 265 5583
rect 2334 6241 2368 6264
rect 2334 6230 2368 6241
rect 2334 6173 2368 6192
rect 2334 6158 2368 6173
rect 5465 5959 5499 5993
rect 5537 5959 5571 5993
rect 2388 5620 2422 5654
rect 2460 5620 2494 5654
rect 231 5549 253 5570
rect 253 5549 265 5570
rect 231 5502 265 5510
rect 231 5476 253 5502
rect 253 5476 265 5502
rect 231 5403 265 5437
rect 231 5330 265 5364
rect 231 5257 265 5291
rect 231 5184 265 5218
rect 1894 5530 1928 5564
rect 1894 5458 1928 5492
rect 2020 5530 2054 5564
rect 2230 5540 2264 5574
rect 2302 5540 2314 5574
rect 2314 5540 2336 5574
rect 2020 5458 2054 5492
rect 3153 5492 3187 5498
rect 3153 5464 3187 5492
rect 1894 5236 1928 5270
rect 1894 5164 1928 5198
rect 2020 5236 2054 5270
rect 2020 5164 2054 5198
rect 2146 5236 2180 5270
rect 2146 5164 2180 5198
rect 2272 5236 2306 5270
rect 2272 5164 2306 5198
rect 2398 5236 2432 5270
rect 2398 5164 2432 5198
rect 2524 5236 2558 5270
rect 2524 5164 2558 5198
rect 2650 5236 2684 5270
rect 2650 5164 2684 5198
rect 2776 5236 2810 5270
rect 2776 5164 2810 5198
rect 2902 5236 2936 5270
rect 2902 5164 2936 5198
rect 3028 5236 3062 5270
rect 3028 5164 3062 5198
rect 231 5111 265 5145
rect 231 5038 265 5072
rect 231 4965 265 4999
rect 231 4893 265 4926
rect 231 4892 265 4893
rect 231 4821 265 4853
rect 231 4819 265 4821
rect 231 4749 265 4780
rect 231 4746 265 4749
rect 231 4677 265 4707
rect 231 4673 265 4677
rect 231 4605 265 4634
rect 231 4600 265 4605
rect 231 4533 265 4561
rect 231 4527 265 4533
rect 231 4461 265 4488
rect 231 4454 265 4461
rect 231 4381 265 4415
rect 1264 4610 1298 4644
rect 1264 4538 1298 4572
rect 231 4319 257 4333
rect 257 4319 265 4333
rect 231 4299 265 4319
rect 382 4353 416 4387
rect 382 4303 416 4315
rect 382 4281 416 4303
rect 382 4073 416 4107
rect 382 4001 416 4035
rect 508 4353 542 4387
rect 508 4303 542 4315
rect 508 4281 542 4303
rect 508 4073 542 4107
rect 508 4001 542 4035
rect 634 4353 668 4387
rect 634 4303 668 4315
rect 634 4281 668 4303
rect 634 4073 668 4107
rect 634 4001 668 4035
rect 760 4353 794 4387
rect 760 4303 794 4315
rect 760 4281 794 4303
rect 760 4073 794 4107
rect 760 4001 794 4035
rect 886 4353 920 4387
rect 886 4303 920 4315
rect 886 4281 920 4303
rect 886 4073 920 4107
rect 886 4001 920 4035
rect 1012 4353 1046 4387
rect 1012 4303 1046 4315
rect 1012 4281 1046 4303
rect 1012 4073 1046 4107
rect 1012 4001 1046 4035
rect 1138 4353 1172 4387
rect 1138 4303 1172 4315
rect 1138 4281 1172 4303
rect 1138 4073 1172 4107
rect 1138 4001 1172 4035
rect 1264 4073 1298 4107
rect 1264 4001 1298 4035
rect 1390 4373 1424 4407
rect 1390 4303 1424 4335
rect 1390 4301 1424 4303
rect 1390 4073 1424 4107
rect 1390 4001 1424 4035
rect 1516 4373 1550 4407
rect 1516 4303 1550 4335
rect 1516 4301 1550 4303
rect 1516 4073 1550 4107
rect 1516 4001 1550 4035
rect 1642 4373 1676 4407
rect 1642 4303 1676 4335
rect 1642 4301 1676 4303
rect 1642 4073 1676 4107
rect 1642 4001 1676 4035
rect 1768 4373 1802 4407
rect 1768 4303 1802 4335
rect 1768 4301 1802 4303
rect 1768 4073 1802 4107
rect 1768 4001 1802 4035
rect 1894 4373 1928 4407
rect 1894 4303 1928 4335
rect 1894 4301 1928 4303
rect 1894 4038 1928 4072
rect 1894 3966 1928 4000
rect 2020 4373 2054 4407
rect 2020 4301 2054 4335
rect 2020 4073 2054 4107
rect 2020 4001 2054 4035
rect 2146 4373 2180 4407
rect 2146 4301 2180 4335
rect 2146 4038 2180 4072
rect 2146 3966 2180 4000
rect 2272 4373 2306 4407
rect 2272 4301 2306 4335
rect 2272 4073 2306 4107
rect 2272 4001 2306 4035
rect 2398 4373 2432 4407
rect 2398 4301 2432 4335
rect 2398 4038 2432 4072
rect 2398 3966 2432 4000
rect 2524 4373 2558 4407
rect 2524 4301 2558 4335
rect 2524 4073 2558 4107
rect 2524 4001 2558 4035
rect 2650 4373 2684 4407
rect 2650 4301 2684 4335
rect 2650 4038 2684 4072
rect 2650 3966 2684 4000
rect 2776 4373 2810 4407
rect 2776 4301 2810 4335
rect 2776 4073 2810 4107
rect 2776 4001 2810 4035
rect 2902 4373 2936 4407
rect 2902 4301 2936 4335
rect 2902 3985 2936 4019
rect 3028 4373 3062 4407
rect 3028 4301 3062 4335
rect 3028 4073 3062 4107
rect 3028 4001 3062 4035
rect 3531 5474 3565 5498
rect 3531 5464 3565 5474
rect 4962 5458 4970 5492
rect 4970 5458 4996 5492
rect 5034 5458 5038 5492
rect 5038 5458 5068 5492
rect 5106 5458 5140 5492
rect 5178 5458 5208 5492
rect 5208 5458 5212 5492
rect 5504 5214 5538 5248
rect 5504 5132 5538 5166
rect 5504 5050 5538 5084
rect 5504 4968 5538 5002
rect 5504 4886 5538 4920
rect 5504 4804 5538 4838
rect 5504 4721 5538 4755
rect 2902 3913 2936 3947
rect 2020 538 2054 572
rect 382 458 416 492
rect 508 458 542 492
rect 634 458 668 492
rect 760 458 794 492
rect 886 458 920 492
rect 1012 458 1046 492
rect 1138 458 1172 492
rect 1264 458 1298 492
rect 1390 458 1424 492
rect 1516 458 1550 492
rect 1642 458 1676 492
rect 1768 458 1802 492
rect 1894 458 1928 492
rect 2020 466 2054 500
rect 2146 538 2180 572
rect 2146 466 2180 500
rect 2272 538 2306 572
rect 2272 466 2306 500
rect 2398 538 2432 572
rect 2398 466 2432 500
rect 2524 458 2558 492
rect 382 408 416 420
rect 382 386 416 408
rect 508 408 542 420
rect 508 386 542 408
rect 634 408 668 420
rect 634 386 668 408
rect 760 408 794 420
rect 760 386 794 408
rect 886 408 920 420
rect 886 386 920 408
rect 1012 408 1046 420
rect 1012 386 1046 408
rect 1138 408 1172 420
rect 1138 386 1172 408
rect 1264 408 1298 420
rect 1264 386 1298 408
rect 1390 408 1424 420
rect 1390 386 1424 408
rect 1516 408 1550 420
rect 1516 386 1550 408
rect 1642 408 1676 420
rect 1642 386 1676 408
rect 1768 408 1802 420
rect 1768 386 1802 408
rect 1894 408 1928 420
rect 1894 386 1928 408
rect 2524 408 2558 420
rect 2524 386 2558 408
rect 2650 458 2684 492
rect 2650 408 2684 420
rect 2650 386 2684 408
rect 2776 458 2810 492
rect 2902 458 2936 492
rect 3028 458 3062 492
rect 2776 408 2810 420
rect 2776 386 2810 408
rect 2902 408 2936 420
rect 2902 386 2936 408
rect 3028 408 3062 420
rect 3028 386 3062 408
rect 3342 828 3376 862
rect 3342 781 3376 786
rect 3342 752 3376 781
rect 3342 679 3376 710
rect 3342 676 3376 679
rect 3342 611 3376 634
rect 3342 600 3376 611
rect 3342 543 3376 558
rect 3342 524 3376 543
rect 3342 475 3376 482
rect 3342 448 3376 475
rect 3342 373 3376 406
rect 3342 372 3376 373
rect 3342 305 3376 330
rect 3342 296 3376 305
rect 3342 237 3376 254
rect 3342 220 3376 237
rect 3342 169 3376 178
rect 3342 144 3376 169
rect 742 69 776 70
rect 742 36 743 69
rect 743 36 776 69
rect 3342 101 3376 102
rect 3342 68 3376 101
rect 742 -33 743 -18
rect 743 -33 776 -18
rect 742 -52 776 -33
rect 3605 -26 3639 6
rect 3605 -28 3639 -26
rect 742 -135 776 -107
rect 742 -141 743 -135
rect 743 -141 776 -135
rect 742 -203 776 -196
rect 742 -230 743 -203
rect 743 -230 776 -203
rect 2458 -90 2492 -56
rect 2458 -162 2492 -128
rect 2914 -78 2948 -44
rect 2914 -150 2948 -116
rect 3370 -90 3404 -56
rect 2458 -234 2492 -200
rect 3370 -162 3404 -128
rect 2547 -240 2581 -206
rect 2619 -240 2653 -206
rect 2691 -240 2725 -206
rect 2763 -240 2797 -206
rect 2835 -240 2869 -206
rect 3370 -234 3404 -200
rect 3605 -94 3639 -67
rect 3605 -101 3639 -94
rect 3605 -162 3639 -140
rect 3605 -174 3639 -162
rect 3605 -230 3639 -213
rect 3605 -247 3639 -230
rect 1997 -314 2031 -280
rect 2069 -314 2103 -280
rect 2337 -314 2371 -280
rect 2409 -314 2443 -280
rect 2998 -314 3009 -280
rect 3009 -314 3032 -280
rect 3070 -314 3093 -280
rect 3093 -314 3104 -280
rect 3142 -314 3143 -280
rect 3143 -314 3176 -280
rect 3214 -314 3226 -280
rect 3226 -314 3248 -280
rect 3605 -298 3639 -286
rect 3605 -320 3639 -298
rect 742 -407 776 -381
rect 742 -415 743 -407
rect 743 -415 776 -407
rect 742 -475 776 -462
rect 742 -496 743 -475
rect 743 -496 776 -475
rect 742 -577 743 -543
rect 743 -577 776 -543
rect 742 -657 776 -623
rect 1681 -399 1714 -371
rect 1714 -399 1715 -371
rect 1756 -399 1790 -365
rect 1830 -399 1861 -365
rect 1861 -399 1864 -365
rect 1904 -399 1929 -365
rect 1929 -399 1938 -365
rect 1978 -399 1997 -365
rect 1997 -399 2012 -365
rect 2052 -399 2065 -365
rect 2065 -399 2086 -365
rect 2126 -399 2133 -365
rect 2133 -399 2160 -365
rect 2200 -399 2201 -365
rect 2201 -399 2234 -365
rect 2274 -399 2303 -365
rect 2303 -399 2308 -365
rect 2348 -399 2371 -365
rect 2371 -399 2382 -365
rect 2422 -399 2439 -365
rect 2439 -399 2456 -365
rect 2496 -399 2507 -365
rect 2507 -399 2530 -365
rect 2570 -399 2575 -365
rect 2575 -399 2604 -365
rect 2644 -399 2677 -365
rect 2677 -399 2678 -365
rect 2718 -399 2745 -365
rect 2745 -399 2752 -365
rect 2792 -399 2813 -365
rect 2813 -399 2826 -365
rect 2866 -399 2881 -365
rect 2881 -399 2900 -365
rect 2940 -399 2949 -365
rect 2949 -399 2974 -365
rect 3014 -399 3017 -365
rect 3017 -399 3048 -365
rect 3088 -399 3119 -365
rect 3119 -399 3122 -365
rect 3162 -399 3187 -365
rect 3187 -399 3196 -365
rect 3236 -399 3255 -365
rect 3255 -399 3270 -365
rect 3310 -399 3323 -365
rect 3323 -399 3344 -365
rect 3384 -399 3391 -365
rect 3391 -399 3418 -365
rect 3458 -399 3459 -365
rect 3459 -399 3492 -365
rect 3533 -399 3567 -365
rect 3605 -366 3639 -359
rect 3605 -393 3639 -366
rect 1681 -405 1715 -399
rect 1681 -494 1715 -464
rect 1681 -498 1715 -494
rect 1681 -562 1715 -557
rect 1681 -591 1715 -562
rect 2149 -587 2183 -560
rect 2149 -594 2183 -587
rect 2221 -588 2255 -554
rect 2294 -588 2308 -554
rect 2308 -588 2328 -554
rect 2367 -588 2376 -554
rect 2376 -588 2401 -554
rect 2440 -588 2444 -554
rect 2444 -588 2474 -554
rect 2513 -588 2546 -554
rect 2546 -588 2547 -554
rect 2586 -588 2614 -554
rect 2614 -588 2620 -554
rect 2659 -588 2682 -554
rect 2682 -588 2693 -554
rect 2732 -588 2750 -554
rect 2750 -588 2766 -554
rect 2805 -588 2818 -554
rect 2818 -588 2839 -554
rect 2878 -588 2886 -554
rect 2886 -588 2912 -554
rect 2951 -588 2954 -554
rect 2954 -588 2985 -554
rect 3024 -588 3056 -554
rect 3056 -588 3058 -554
rect 3097 -588 3124 -554
rect 3124 -588 3131 -554
rect 3170 -588 3192 -554
rect 3192 -588 3204 -554
rect 3243 -588 3260 -554
rect 3260 -588 3277 -554
rect 3317 -588 3328 -554
rect 3328 -588 3351 -554
rect 3391 -588 3396 -554
rect 3396 -588 3425 -554
rect 3463 -588 3464 -560
rect 3464 -588 3497 -560
rect 3463 -594 3497 -588
rect 2149 -655 2183 -645
rect 2149 -679 2183 -655
rect 2285 -673 2303 -639
rect 2303 -673 2319 -639
rect 2357 -673 2371 -639
rect 2371 -673 2391 -639
rect 2455 -673 2489 -639
rect 2527 -673 2543 -639
rect 2543 -673 2561 -639
rect 2975 -673 3009 -639
rect 3047 -673 3069 -639
rect 3069 -673 3081 -639
rect 2149 -757 2183 -731
rect 2149 -765 2183 -757
rect 2149 -825 2183 -817
rect 2149 -851 2183 -825
rect 2266 -753 2300 -719
rect 2266 -825 2300 -791
rect 2698 -753 2732 -719
rect 2149 -937 2183 -903
rect 2482 -852 2516 -818
rect 2698 -825 2732 -791
rect 3130 -753 3164 -719
rect 2482 -924 2516 -890
rect 2914 -852 2948 -818
rect 3130 -825 3164 -791
rect 3463 -656 3497 -646
rect 3463 -680 3497 -656
rect 3463 -758 3497 -732
rect 3463 -766 3497 -758
rect 2914 -924 2948 -890
rect 3346 -852 3380 -818
rect 3346 -924 3380 -890
rect 2149 -995 2183 -989
rect 2149 -1023 2182 -995
rect 2182 -1023 2183 -995
rect 2221 -1029 2250 -995
rect 2250 -1029 2255 -995
rect 2294 -1029 2318 -995
rect 2318 -1029 2328 -995
rect 2367 -1029 2386 -995
rect 2386 -1029 2401 -995
rect 2440 -1029 2454 -995
rect 2454 -1029 2474 -995
rect 2513 -1029 2522 -995
rect 2522 -1029 2547 -995
rect 2586 -1029 2590 -995
rect 2590 -1029 2620 -995
rect 2659 -1029 2692 -995
rect 2692 -1029 2693 -995
rect 2732 -1029 2760 -995
rect 2760 -1029 2766 -995
rect 2805 -1029 2828 -995
rect 2828 -1029 2839 -995
rect 2878 -1029 2896 -995
rect 2896 -1029 2912 -995
rect 2951 -1029 2964 -995
rect 2964 -1029 2985 -995
rect 3024 -1029 3032 -995
rect 3032 -1029 3058 -995
rect 3097 -1029 3100 -995
rect 3100 -1029 3131 -995
rect 3170 -1029 3202 -995
rect 3202 -1029 3204 -995
rect 3243 -1029 3270 -995
rect 3270 -1029 3277 -995
rect 3317 -1029 3338 -995
rect 3338 -1029 3351 -995
rect 3391 -1029 3425 -995
<< metal1 >>
tri 1604 27912 1606 27914 se
rect 1606 27912 1652 27914
tri 310 27878 344 27912 se
rect 344 27878 394 27912
tri 394 27878 428 27912 sw
tri 1570 27878 1604 27912 se
rect 1604 27878 1652 27912
tri 1652 27878 1688 27914 sw
tri 99 27869 108 27878 se
rect 108 27869 138 27878
rect 190 27869 202 27878
rect 254 27869 266 27878
rect 318 27877 1936 27878
tri 1936 27877 1937 27878 sw
rect 318 27875 1937 27877
tri 1937 27875 1939 27877 sw
tri 2118 27875 2120 27877 se
rect 2120 27875 2373 27877
rect 318 27871 1939 27875
tri 1939 27871 1943 27875 sw
tri 2114 27871 2118 27875 se
rect 2118 27871 2373 27875
rect 318 27869 2373 27871
tri 65 27835 99 27869 se
rect 99 27835 138 27869
rect 318 27835 1673 27869
rect 1707 27835 1745 27869
rect 1779 27835 1817 27869
rect 1851 27835 1889 27869
rect 1923 27835 2373 27869
tri 62 27832 65 27835 se
rect 65 27832 138 27835
rect 62 27826 138 27832
rect 190 27826 202 27835
rect 254 27826 266 27835
rect 318 27826 2373 27835
rect 62 27785 108 27826
tri 108 27798 136 27826 nw
tri 2097 27798 2125 27826 ne
rect 2125 27798 2373 27826
rect 62 27751 68 27785
rect 102 27751 108 27785
rect 62 27711 108 27751
rect 62 27677 68 27711
rect 102 27677 108 27711
tri 273 27699 357 27783 se
rect 357 27713 540 27783
tri 357 27699 371 27713 nw
rect 62 27637 108 27677
rect 62 27603 68 27637
rect 102 27603 108 27637
rect 62 27563 108 27603
rect 62 27529 68 27563
rect 102 27529 108 27563
rect 62 27489 108 27529
rect 62 27455 68 27489
rect 102 27455 108 27489
tri 248 27674 273 27699 se
rect 273 27674 332 27699
tri 332 27674 357 27699 nw
rect 248 27667 325 27674
tri 325 27667 332 27674 nw
rect 534 27667 540 27713
rect 656 27731 724 27783
rect 776 27731 796 27783
rect 848 27731 868 27783
rect 920 27731 940 27783
rect 992 27731 1011 27783
rect 1063 27731 1082 27783
rect 1134 27731 1153 27783
rect 1205 27731 1224 27783
rect 1276 27731 1344 27783
rect 656 27719 1344 27731
rect 656 27713 724 27719
rect 656 27667 662 27713
rect 718 27667 724 27713
rect 776 27667 796 27719
rect 848 27667 868 27719
rect 920 27667 940 27719
rect 992 27667 1011 27719
rect 1063 27667 1082 27719
rect 1134 27667 1153 27719
rect 1205 27667 1224 27719
rect 1276 27713 1344 27719
rect 1276 27667 1282 27713
rect 1338 27667 1344 27713
rect 1460 27746 1569 27783
tri 1569 27746 1606 27783 sw
rect 1685 27746 1691 27798
rect 1743 27746 1755 27798
rect 1807 27746 1819 27798
rect 1871 27782 2063 27798
tri 2063 27782 2079 27798 sw
tri 2125 27782 2141 27798 ne
rect 2141 27782 2373 27798
rect 1871 27764 2079 27782
tri 2079 27764 2097 27782 sw
tri 2141 27764 2159 27782 ne
rect 2159 27764 2373 27782
rect 1871 27746 2097 27764
tri 2097 27746 2115 27764 sw
tri 2159 27746 2177 27764 ne
rect 2177 27746 2373 27764
rect 1460 27718 1606 27746
tri 1606 27718 1634 27746 sw
tri 2047 27718 2075 27746 ne
rect 2075 27718 2115 27746
tri 2115 27718 2143 27746 sw
tri 2177 27718 2205 27746 ne
rect 2205 27718 2373 27746
rect 1460 27713 1634 27718
tri 1634 27713 1639 27718 sw
tri 1785 27713 1790 27718 se
rect 1790 27713 1802 27718
rect 1460 27667 1466 27713
rect 1796 27667 1802 27713
rect 248 27666 324 27667
tri 324 27666 325 27667 nw
tri 1787 27666 1788 27667 ne
rect 1788 27666 1802 27667
rect 1854 27666 1866 27718
rect 1918 27666 1930 27718
rect 1982 27713 2004 27718
tri 2004 27713 2009 27718 sw
tri 2075 27714 2079 27718 ne
rect 2079 27714 2143 27718
tri 2143 27714 2147 27718 sw
tri 2205 27714 2209 27718 ne
rect 2209 27714 2373 27718
tri 2079 27713 2080 27714 ne
rect 2080 27713 2147 27714
tri 2147 27713 2148 27714 sw
tri 2209 27713 2210 27714 ne
rect 2210 27713 2373 27714
rect 1982 27667 1988 27713
tri 2080 27696 2097 27713 ne
rect 2097 27696 2148 27713
tri 2097 27667 2126 27696 ne
rect 2126 27667 2148 27696
rect 1982 27666 2039 27667
tri 2126 27666 2127 27667 ne
rect 2127 27666 2148 27667
tri 2148 27666 2195 27713 sw
tri 2210 27666 2257 27713 ne
rect 2257 27666 2373 27713
rect 248 27465 300 27666
tri 300 27642 324 27666 nw
tri 2127 27646 2147 27666 ne
rect 2147 27646 2195 27666
tri 2195 27646 2215 27666 sw
tri 2257 27646 2277 27666 ne
rect 2277 27646 2373 27666
tri 2147 27642 2151 27646 ne
rect 2151 27642 2215 27646
tri 2215 27642 2219 27646 sw
tri 2277 27642 2281 27646 ne
rect 2281 27642 2373 27646
tri 2151 27637 2156 27642 ne
rect 2156 27637 2219 27642
tri 2219 27637 2224 27642 sw
tri 2281 27637 2286 27642 ne
rect 2286 27637 2373 27642
rect 1010 27585 1016 27637
rect 1068 27585 1080 27637
rect 1132 27585 1144 27637
rect 1196 27585 1208 27637
rect 1260 27585 1344 27637
rect 1396 27585 1408 27637
rect 1460 27585 1802 27637
rect 1854 27585 1866 27637
rect 1918 27585 1930 27637
rect 1982 27595 2015 27637
tri 2015 27595 2057 27637 sw
tri 2156 27595 2198 27637 ne
rect 2198 27595 2224 27637
tri 2224 27595 2266 27637 sw
tri 2286 27595 2328 27637 ne
rect 1982 27586 2057 27595
tri 2057 27586 2066 27595 sw
rect 1982 27585 2066 27586
tri 2198 27585 2208 27595 ne
rect 2208 27585 2266 27595
tri 2266 27585 2276 27595 sw
tri 1983 27578 1990 27585 ne
rect 1990 27578 2066 27585
tri 2208 27578 2215 27585 ne
rect 2215 27578 2276 27585
tri 2276 27578 2283 27585 sw
tri 1990 27562 2006 27578 ne
rect 2006 27562 2066 27578
tri 2215 27562 2231 27578 ne
tri 2006 27560 2008 27562 ne
rect 370 27551 428 27557
rect 370 27517 382 27551
rect 416 27517 428 27551
rect 370 27479 428 27517
rect 62 27415 108 27455
rect 62 27381 68 27415
rect 102 27381 108 27415
rect 62 27342 108 27381
rect 62 27308 68 27342
rect 102 27308 108 27342
rect 62 27269 108 27308
rect 62 27235 68 27269
rect 102 27235 108 27269
rect 62 27196 108 27235
rect 62 27162 68 27196
rect 102 27162 108 27196
rect 62 27123 108 27162
rect 62 27089 68 27123
rect 102 27089 108 27123
rect 62 27050 108 27089
rect 62 27016 68 27050
rect 102 27016 108 27050
rect 62 26977 108 27016
rect 62 26943 68 26977
rect 102 26943 108 26977
rect 62 26904 108 26943
rect 62 26870 68 26904
rect 102 26870 108 26904
rect 62 26831 108 26870
rect 62 26797 68 26831
rect 102 26797 108 26831
rect 62 26758 108 26797
rect 62 26724 68 26758
rect 102 26724 108 26758
rect 62 26685 108 26724
rect 62 26651 68 26685
rect 102 26651 108 26685
rect 62 26612 108 26651
rect 62 26578 68 26612
rect 102 26578 108 26612
rect 62 26539 108 26578
rect 62 26505 68 26539
rect 102 26505 108 26539
rect 62 26466 108 26505
rect 62 26432 68 26466
rect 102 26432 108 26466
rect 62 26393 108 26432
rect 62 26359 68 26393
rect 102 26359 108 26393
rect 62 26320 108 26359
rect 62 26286 68 26320
rect 102 26286 108 26320
rect 62 26247 108 26286
rect 62 26213 68 26247
rect 102 26213 108 26247
rect 62 26174 108 26213
rect 62 26140 68 26174
rect 102 26140 108 26174
rect 62 26101 108 26140
rect 62 26067 68 26101
rect 102 26067 108 26101
rect 62 26028 108 26067
rect 62 25994 68 26028
rect 102 25994 108 26028
rect 62 25955 108 25994
rect 62 25921 68 25955
rect 102 25921 108 25955
rect 62 25882 108 25921
rect 62 25848 68 25882
rect 102 25848 108 25882
rect 62 25809 108 25848
rect 62 25775 68 25809
rect 102 25775 108 25809
rect 62 25736 108 25775
rect 62 25702 68 25736
rect 102 25702 108 25736
rect 62 25690 108 25702
rect 370 27445 382 27479
rect 416 27445 428 27479
rect 370 23862 428 27445
rect 496 27551 680 27557
rect 496 27517 508 27551
rect 542 27517 634 27551
rect 668 27517 680 27551
rect 496 27479 680 27517
rect 496 27445 508 27479
rect 542 27445 634 27479
rect 668 27445 680 27479
rect 496 27439 680 27445
rect 748 27551 932 27557
rect 748 27517 760 27551
rect 794 27517 886 27551
rect 920 27517 932 27551
rect 748 27479 932 27517
rect 748 27445 760 27479
rect 794 27445 886 27479
rect 920 27445 932 27479
rect 748 27439 932 27445
rect 496 27387 538 27439
tri 538 27414 563 27439 nw
tri 597 27414 622 27439 ne
rect 497 27385 537 27386
rect 370 23828 382 23862
rect 416 23828 428 23862
rect 370 23790 428 23828
rect 370 23756 382 23790
rect 416 23756 428 23790
rect 370 23656 428 23756
rect 370 23622 382 23656
rect 416 23622 428 23656
rect 370 23584 428 23622
rect 370 23550 382 23584
rect 416 23550 428 23584
rect 370 19967 428 23550
rect 497 27348 537 27349
rect 496 27295 538 27347
tri 538 27295 554 27311 sw
rect 496 23862 554 27295
rect 622 23960 680 27439
tri 849 27414 874 27439 ne
rect 623 23958 679 23959
rect 874 23960 932 27439
rect 1000 27551 1184 27557
rect 1000 27517 1012 27551
rect 1046 27517 1138 27551
rect 1172 27517 1184 27551
rect 1000 27479 1184 27517
rect 1000 27445 1012 27479
rect 1046 27445 1138 27479
rect 1172 27445 1184 27479
rect 1000 27439 1184 27445
rect 1252 27551 1436 27557
rect 1252 27517 1264 27551
rect 1298 27517 1390 27551
rect 1424 27517 1436 27551
rect 1252 27479 1436 27517
rect 1252 27445 1264 27479
rect 1298 27445 1390 27479
rect 1424 27445 1436 27479
rect 1252 27439 1436 27445
rect 1504 27551 1688 27557
rect 1504 27517 1516 27551
rect 1550 27517 1642 27551
rect 1676 27517 1688 27551
rect 1504 27479 1688 27517
rect 1504 27445 1516 27479
rect 1550 27445 1642 27479
rect 1676 27445 1688 27479
rect 1504 27439 1688 27445
rect 1756 27551 1940 27557
rect 1756 27517 1768 27551
rect 1802 27517 1894 27551
rect 1928 27517 1940 27551
rect 1756 27479 1940 27517
rect 1756 27445 1768 27479
rect 1802 27445 1894 27479
rect 1928 27445 1940 27479
rect 1756 27439 1940 27445
rect 2008 27551 2066 27562
rect 2008 27517 2020 27551
rect 2054 27517 2066 27551
rect 2008 27479 2066 27517
rect 2008 27445 2020 27479
rect 2054 27445 2066 27479
rect 2008 27439 2066 27445
rect 1000 27387 1048 27439
tri 1048 27414 1073 27439 nw
tri 2124 27387 2139 27402 se
tri 2123 27386 2124 27387 se
rect 2124 27386 2139 27387
rect 1001 27385 1047 27386
tri 2122 27385 2123 27386 se
rect 2123 27385 2139 27386
tri 2114 27377 2122 27385 se
rect 2122 27377 2139 27385
rect 875 23958 931 23959
rect 1001 27348 1047 27349
rect 1000 27295 1048 27347
tri 1048 27295 1058 27305 sw
rect 496 23828 508 23862
rect 542 23828 554 23862
rect 496 23790 554 23828
rect 496 23756 508 23790
rect 542 23756 554 23790
rect 496 23656 554 23756
rect 496 23622 508 23656
rect 542 23622 554 23656
rect 496 23584 554 23622
rect 496 23550 508 23584
rect 542 23550 554 23584
rect 496 23492 554 23550
rect 497 23490 553 23491
rect 623 23921 679 23922
rect 622 23862 680 23920
rect 875 23921 931 23922
rect 622 23828 634 23862
rect 668 23828 680 23862
rect 622 23790 680 23828
rect 622 23756 634 23790
rect 668 23756 680 23790
rect 622 23656 680 23756
rect 622 23622 634 23656
rect 668 23622 680 23656
rect 622 23584 680 23622
rect 622 23550 634 23584
rect 668 23550 680 23584
rect 370 19933 382 19967
rect 416 19933 428 19967
rect 370 19895 428 19933
rect 370 19861 382 19895
rect 416 19861 428 19895
rect 370 19761 428 19861
rect 370 19727 382 19761
rect 416 19727 428 19761
rect 370 19689 428 19727
rect 370 19655 382 19689
rect 416 19655 428 19689
rect 370 16072 428 19655
rect 497 23453 553 23454
rect 496 19967 554 23452
rect 622 20065 680 23550
rect 748 23862 806 23868
rect 748 23828 760 23862
rect 794 23828 806 23862
rect 748 23790 806 23828
rect 748 23756 760 23790
rect 794 23756 806 23790
rect 748 23656 806 23756
rect 748 23622 760 23656
rect 794 23622 806 23656
rect 748 23584 806 23622
rect 748 23550 760 23584
rect 794 23550 806 23584
rect 748 23544 806 23550
rect 874 23862 932 23920
rect 874 23828 886 23862
rect 920 23828 932 23862
rect 874 23790 932 23828
rect 874 23756 886 23790
rect 920 23756 932 23790
rect 874 23656 932 23756
rect 874 23622 886 23656
rect 920 23622 932 23656
rect 874 23584 932 23622
rect 874 23550 886 23584
rect 920 23550 932 23584
rect 623 20063 679 20064
rect 874 20065 932 23550
rect 1000 23862 1058 27295
rect 2017 23921 2185 27377
tri 2114 23896 2139 23921 ne
rect 2139 23896 2185 23921
rect 1000 23828 1012 23862
rect 1046 23828 1058 23862
rect 1000 23790 1058 23828
rect 1000 23756 1012 23790
rect 1046 23756 1058 23790
rect 1000 23656 1058 23756
rect 1000 23622 1012 23656
rect 1046 23622 1058 23656
rect 1000 23584 1058 23622
rect 1000 23550 1012 23584
rect 1046 23550 1058 23584
rect 1000 23492 1058 23550
rect 1126 23862 1184 23868
rect 1126 23828 1138 23862
rect 1172 23828 1184 23862
rect 1126 23790 1184 23828
rect 1126 23756 1138 23790
rect 1172 23756 1184 23790
rect 1126 23656 1184 23756
rect 1126 23622 1138 23656
rect 1172 23622 1184 23656
rect 1126 23584 1184 23622
rect 1126 23550 1138 23584
rect 1172 23550 1184 23584
rect 1126 23544 1184 23550
rect 1252 23862 1310 23868
rect 1252 23828 1264 23862
rect 1298 23828 1310 23862
rect 1252 23790 1310 23828
rect 1252 23756 1264 23790
rect 1298 23756 1310 23790
rect 1252 23656 1310 23756
rect 1252 23622 1264 23656
rect 1298 23622 1310 23656
rect 1252 23584 1310 23622
rect 1252 23550 1264 23584
rect 1298 23550 1310 23584
rect 1252 23544 1310 23550
rect 1378 23862 1436 23868
rect 1378 23828 1390 23862
rect 1424 23828 1436 23862
rect 1378 23790 1436 23828
rect 1378 23756 1390 23790
rect 1424 23756 1436 23790
rect 1378 23656 1436 23756
rect 1378 23622 1390 23656
rect 1424 23622 1436 23656
rect 1378 23584 1436 23622
rect 1378 23550 1390 23584
rect 1424 23550 1436 23584
rect 1378 23544 1436 23550
rect 1504 23862 1562 23868
rect 1504 23828 1516 23862
rect 1550 23828 1562 23862
rect 1504 23790 1562 23828
rect 1504 23756 1516 23790
rect 1550 23756 1562 23790
rect 1504 23656 1562 23756
rect 1504 23622 1516 23656
rect 1550 23622 1562 23656
rect 1504 23584 1562 23622
rect 1504 23550 1516 23584
rect 1550 23550 1562 23584
rect 1504 23544 1562 23550
rect 1630 23862 1688 23868
rect 1630 23828 1642 23862
rect 1676 23828 1688 23862
rect 1630 23790 1688 23828
rect 1630 23756 1642 23790
rect 1676 23756 1688 23790
rect 1630 23656 1688 23756
rect 1630 23622 1642 23656
rect 1676 23622 1688 23656
rect 1630 23584 1688 23622
rect 1630 23550 1642 23584
rect 1676 23550 1688 23584
rect 1630 23544 1688 23550
rect 1756 23862 1814 23868
rect 1756 23828 1768 23862
rect 1802 23828 1814 23862
rect 1756 23790 1814 23828
rect 1756 23756 1768 23790
rect 1802 23756 1814 23790
rect 1756 23656 1814 23756
rect 1756 23622 1768 23656
rect 1802 23622 1814 23656
rect 1756 23584 1814 23622
rect 1756 23550 1768 23584
rect 1802 23550 1814 23584
rect 1756 23544 1814 23550
rect 1882 23862 1940 23868
rect 1882 23828 1894 23862
rect 1928 23828 1940 23862
rect 1882 23790 1940 23828
rect 1882 23756 1894 23790
rect 1928 23756 1940 23790
rect 1882 23656 1940 23756
rect 1882 23622 1894 23656
rect 1928 23622 1940 23656
rect 1882 23584 1940 23622
rect 1882 23550 1894 23584
rect 1928 23550 1940 23584
rect 1882 23544 1940 23550
rect 2008 23862 2066 23868
rect 2008 23828 2020 23862
rect 2054 23828 2066 23862
rect 2008 23790 2066 23828
rect 2008 23756 2020 23790
rect 2054 23756 2066 23790
rect 2008 23656 2066 23756
rect 2008 23622 2020 23656
rect 2054 23622 2066 23656
rect 2008 23584 2066 23622
rect 2008 23550 2020 23584
rect 2054 23550 2066 23584
rect 2008 23544 2066 23550
tri 2114 23503 2139 23528 se
rect 2139 23503 2185 23528
rect 1001 23490 1057 23491
rect 875 20063 931 20064
rect 1001 23453 1057 23454
rect 496 19933 508 19967
rect 542 19933 554 19967
rect 496 19895 554 19933
rect 496 19861 508 19895
rect 542 19861 554 19895
rect 496 19761 554 19861
rect 496 19727 508 19761
rect 542 19727 554 19761
rect 496 19689 554 19727
rect 496 19655 508 19689
rect 542 19655 554 19689
rect 496 19649 554 19655
rect 623 20026 679 20027
rect 622 19967 680 20025
rect 875 20026 931 20027
rect 622 19933 634 19967
rect 668 19933 680 19967
rect 622 19895 680 19933
rect 622 19861 634 19895
rect 668 19861 680 19895
rect 622 19761 680 19861
rect 622 19727 634 19761
rect 668 19727 680 19761
rect 622 19689 680 19727
rect 622 19655 634 19689
rect 668 19655 680 19689
rect 622 16170 680 19655
rect 748 19967 806 19973
rect 748 19933 760 19967
rect 794 19933 806 19967
rect 748 19895 806 19933
rect 748 19861 760 19895
rect 794 19861 806 19895
rect 748 19761 806 19861
rect 748 19727 760 19761
rect 794 19727 806 19761
rect 748 19689 806 19727
rect 748 19655 760 19689
rect 794 19655 806 19689
rect 748 19597 806 19655
rect 749 19595 805 19596
rect 874 19967 932 20025
rect 874 19933 886 19967
rect 920 19933 932 19967
rect 874 19895 932 19933
rect 874 19861 886 19895
rect 920 19861 932 19895
rect 874 19761 932 19861
rect 874 19727 886 19761
rect 920 19727 932 19761
rect 874 19689 932 19727
rect 874 19655 886 19689
rect 920 19655 932 19689
rect 623 16168 679 16169
rect 749 19558 805 19559
rect 623 16131 679 16132
rect 370 16038 382 16072
rect 416 16038 428 16072
rect 370 16000 428 16038
rect 370 15966 382 16000
rect 416 15966 428 16000
rect 370 15866 428 15966
rect 370 15832 382 15866
rect 416 15832 428 15866
rect 370 15794 428 15832
rect 370 15760 382 15794
rect 416 15760 428 15794
rect 370 12177 428 15760
rect 496 16072 554 16078
rect 496 16038 508 16072
rect 542 16038 554 16072
rect 496 16000 554 16038
rect 496 15966 508 16000
rect 542 15966 554 16000
rect 496 15866 554 15966
rect 496 15832 508 15866
rect 542 15832 554 15866
rect 496 15794 554 15832
rect 496 15760 508 15794
rect 542 15760 554 15794
rect 496 15754 554 15760
rect 622 16072 680 16130
rect 622 16038 634 16072
rect 668 16038 680 16072
rect 622 16000 680 16038
rect 622 15966 634 16000
rect 668 15966 680 16000
rect 622 15866 680 15966
rect 622 15832 634 15866
rect 668 15832 680 15866
rect 622 15794 680 15832
rect 622 15760 634 15794
rect 668 15760 680 15794
rect 622 12275 680 15760
rect 748 16072 806 19557
rect 874 16170 932 19655
rect 1000 19967 1058 23452
tri 1965 22427 2017 22479 ne
rect 1378 22391 1436 22397
rect 1378 22357 1390 22391
rect 1424 22357 1436 22391
rect 1378 22319 1436 22357
rect 1378 22285 1390 22319
rect 1424 22285 1436 22319
rect 1000 19933 1012 19967
rect 1046 19933 1058 19967
rect 1000 19895 1058 19933
rect 1000 19861 1012 19895
rect 1046 19861 1058 19895
rect 1000 19761 1058 19861
rect 1000 19727 1012 19761
rect 1046 19727 1058 19761
rect 1000 19689 1058 19727
rect 1000 19655 1012 19689
rect 1046 19655 1058 19689
rect 1000 19597 1058 19655
rect 1001 19595 1057 19596
rect 1126 19967 1184 19973
rect 1126 19933 1138 19967
rect 1172 19933 1184 19967
rect 1126 19895 1184 19933
rect 1126 19861 1138 19895
rect 1172 19861 1184 19895
rect 1126 19761 1184 19861
rect 1126 19727 1138 19761
rect 1172 19727 1184 19761
rect 1126 19689 1184 19727
rect 1126 19655 1138 19689
rect 1172 19655 1184 19689
rect 875 16168 931 16169
rect 1001 19558 1057 19559
rect 748 16038 760 16072
rect 794 16038 806 16072
rect 748 16000 806 16038
rect 748 15966 760 16000
rect 794 15966 806 16000
rect 748 15866 806 15966
rect 748 15832 760 15866
rect 794 15832 806 15866
rect 748 15794 806 15832
rect 748 15760 760 15794
rect 794 15760 806 15794
rect 748 15702 806 15760
rect 749 15700 805 15701
rect 875 16131 931 16132
rect 874 16072 932 16130
rect 874 16038 886 16072
rect 920 16038 932 16072
rect 874 16000 932 16038
rect 874 15966 886 16000
rect 920 15966 932 16000
rect 874 15866 932 15966
rect 874 15832 886 15866
rect 920 15832 932 15866
rect 874 15794 932 15832
rect 874 15760 886 15794
rect 920 15760 932 15794
rect 623 12273 679 12274
rect 749 15663 805 15664
rect 623 12236 679 12237
rect 370 12143 382 12177
rect 416 12143 428 12177
rect 370 12105 428 12143
rect 370 12071 382 12105
rect 416 12071 428 12105
rect 370 11971 428 12071
rect 370 11937 382 11971
rect 416 11937 428 11971
rect 370 11899 428 11937
rect 370 11865 382 11899
rect 416 11865 428 11899
rect 370 8282 428 11865
rect 496 12177 554 12183
rect 496 12143 508 12177
rect 542 12143 554 12177
rect 496 12105 554 12143
rect 496 12071 508 12105
rect 542 12071 554 12105
rect 496 11971 554 12071
rect 496 11937 508 11971
rect 542 11937 554 11971
rect 496 11899 554 11937
rect 496 11865 508 11899
rect 542 11865 554 11899
rect 496 11807 554 11865
rect 622 12177 680 12235
rect 622 12143 634 12177
rect 668 12143 680 12177
rect 622 12105 680 12143
rect 622 12071 634 12105
rect 668 12071 680 12105
rect 622 11971 680 12071
rect 622 11937 634 11971
rect 668 11937 680 11971
rect 622 11899 680 11937
rect 622 11865 634 11899
rect 668 11865 680 11899
rect 622 11859 680 11865
rect 748 12177 806 15662
rect 874 12275 932 15760
rect 1000 16072 1058 19557
rect 1126 16170 1184 19655
rect 1252 19967 1310 19973
rect 1252 19933 1264 19967
rect 1298 19933 1310 19967
rect 1252 19895 1310 19933
rect 1252 19861 1264 19895
rect 1298 19861 1310 19895
rect 1252 19761 1310 19861
rect 1252 19727 1264 19761
rect 1298 19727 1310 19761
rect 1252 19689 1310 19727
rect 1252 19655 1264 19689
rect 1298 19655 1310 19689
rect 1252 19649 1310 19655
rect 1378 19761 1436 22285
rect 1630 22391 1688 22397
rect 1630 22357 1642 22391
rect 1676 22357 1688 22391
rect 1630 22319 1688 22357
rect 1630 22285 1642 22319
rect 1676 22285 1688 22319
rect 1378 19727 1390 19761
rect 1424 19727 1436 19761
rect 1378 19689 1436 19727
rect 1378 19655 1390 19689
rect 1424 19655 1436 19689
rect 1127 16168 1183 16169
rect 1378 16170 1436 19655
rect 1504 19967 1562 19973
rect 1504 19933 1516 19967
rect 1550 19933 1562 19967
rect 1504 19895 1562 19933
rect 1504 19861 1516 19895
rect 1550 19861 1562 19895
rect 1504 19761 1562 19861
rect 1504 19727 1516 19761
rect 1550 19727 1562 19761
rect 1504 19689 1562 19727
rect 1504 19655 1516 19689
rect 1550 19655 1562 19689
rect 1504 19649 1562 19655
rect 1630 19761 1688 22285
rect 1882 22391 1940 22397
rect 1882 22357 1894 22391
rect 1928 22357 1940 22391
rect 1882 22319 1940 22357
rect 1882 22285 1894 22319
rect 1928 22285 1940 22319
rect 1882 22279 1940 22285
rect 1630 19727 1642 19761
rect 1676 19727 1688 19761
rect 1630 19689 1688 19727
rect 1630 19655 1642 19689
rect 1676 19655 1688 19689
rect 1379 16168 1435 16169
rect 1630 16170 1688 19655
rect 1756 19967 1814 19973
rect 1756 19933 1768 19967
rect 1802 19933 1814 19967
rect 1756 19895 1814 19933
rect 1756 19861 1768 19895
rect 1802 19861 1814 19895
rect 1756 19761 1814 19861
rect 1756 19727 1768 19761
rect 1802 19727 1814 19761
rect 1756 19689 1814 19727
rect 1756 19655 1768 19689
rect 1802 19655 1814 19689
rect 1756 19649 1814 19655
rect 1882 19767 1937 22279
tri 1937 22276 1940 22279 nw
tri 1965 22223 2017 22275 se
rect 2017 20047 2185 23503
tri 2114 20022 2139 20047 ne
rect 2139 20022 2185 20047
rect 2008 19967 2066 19973
rect 2008 19933 2020 19967
rect 2054 19933 2066 19967
rect 2008 19895 2066 19933
rect 2008 19861 2020 19895
rect 2054 19861 2066 19895
tri 1937 19767 1940 19770 sw
rect 1882 19761 1940 19767
rect 1882 19727 1894 19761
rect 1928 19727 1940 19761
rect 1882 19689 1940 19727
rect 1882 19655 1894 19689
rect 1928 19655 1940 19689
rect 1882 19649 1940 19655
rect 2008 19761 2066 19861
rect 2008 19727 2020 19761
rect 2054 19727 2066 19761
rect 2008 19689 2066 19727
rect 2008 19655 2020 19689
rect 2054 19655 2066 19689
rect 2008 19649 2066 19655
rect 1631 16168 1687 16169
rect 1882 16170 1937 19649
tri 1937 19646 1940 19649 nw
tri 2114 19608 2139 19633 se
rect 2139 19608 2185 19633
rect 1883 16168 1936 16169
rect 2017 16152 2185 19608
tri 2114 16132 2134 16152 ne
rect 2134 16132 2185 16152
rect 1000 16038 1012 16072
rect 1046 16038 1058 16072
rect 1000 16000 1058 16038
rect 1000 15966 1012 16000
rect 1046 15966 1058 16000
rect 1000 15866 1058 15966
rect 1000 15832 1012 15866
rect 1046 15832 1058 15866
rect 1000 15794 1058 15832
rect 1000 15760 1012 15794
rect 1046 15760 1058 15794
rect 1000 15702 1058 15760
rect 1001 15700 1057 15701
rect 1127 16131 1183 16132
rect 1126 16072 1184 16130
rect 1379 16131 1435 16132
rect 1126 16038 1138 16072
rect 1172 16038 1184 16072
rect 1126 16000 1184 16038
rect 1126 15966 1138 16000
rect 1172 15966 1184 16000
rect 1126 15866 1184 15966
rect 1126 15832 1138 15866
rect 1172 15832 1184 15866
rect 1126 15794 1184 15832
rect 1126 15760 1138 15794
rect 1172 15760 1184 15794
rect 875 12273 931 12274
rect 1001 15663 1057 15664
rect 748 12143 760 12177
rect 794 12143 806 12177
rect 748 12105 806 12143
rect 748 12071 760 12105
rect 794 12071 806 12105
rect 748 11971 806 12071
rect 748 11937 760 11971
rect 794 11937 806 11971
rect 748 11899 806 11937
rect 748 11865 760 11899
rect 794 11865 806 11899
rect 497 11805 553 11806
rect 748 11807 806 11865
rect 749 11805 805 11806
rect 875 12236 931 12237
rect 874 12177 932 12235
rect 874 12143 886 12177
rect 920 12143 932 12177
rect 874 12105 932 12143
rect 874 12071 886 12105
rect 920 12071 932 12105
rect 874 11971 932 12071
rect 874 11937 886 11971
rect 920 11937 932 11971
rect 874 11899 932 11937
rect 874 11865 886 11899
rect 920 11865 932 11899
rect 370 8248 382 8282
rect 416 8248 428 8282
rect 370 8210 428 8248
rect 370 8176 382 8210
rect 416 8176 428 8210
rect 370 8076 428 8176
rect 370 8042 382 8076
rect 416 8042 428 8076
rect 370 8004 428 8042
rect 370 7970 382 8004
rect 416 7970 428 8004
tri 225 6834 248 6857 se
rect 248 6834 300 6857
rect 225 6759 300 6834
rect 225 6725 231 6759
rect 265 6725 300 6759
rect 225 6685 300 6725
rect 225 6651 231 6685
rect 265 6651 300 6685
rect 225 6611 300 6651
rect 225 6577 231 6611
rect 265 6577 300 6611
rect 225 6537 300 6577
rect 225 6503 231 6537
rect 265 6503 300 6537
rect 225 6463 300 6503
rect 225 6429 231 6463
rect 265 6429 300 6463
rect 225 6389 300 6429
rect 225 6355 231 6389
rect 265 6355 300 6389
rect 225 6315 300 6355
rect 225 6281 231 6315
rect 265 6281 300 6315
rect 225 6241 300 6281
rect 225 6207 231 6241
rect 265 6207 300 6241
rect 225 6167 300 6207
rect 225 6133 231 6167
rect 265 6133 300 6167
rect 225 6094 300 6133
rect 225 6060 231 6094
rect 265 6060 300 6094
rect 225 6021 300 6060
rect 225 5987 231 6021
rect 265 5987 300 6021
rect 225 5948 300 5987
rect 225 5914 231 5948
rect 265 5914 300 5948
rect 225 5875 300 5914
rect 225 5841 231 5875
rect 265 5841 300 5875
rect 225 5802 300 5841
rect 225 5768 231 5802
rect 265 5768 300 5802
rect 225 5729 300 5768
rect 225 5695 231 5729
rect 265 5695 300 5729
rect 225 5656 300 5695
rect 225 5622 231 5656
rect 265 5622 300 5656
rect 225 5583 300 5622
rect 225 5549 231 5583
rect 265 5549 300 5583
rect 225 5510 300 5549
rect 225 5476 231 5510
rect 265 5476 300 5510
rect 225 5437 300 5476
rect 225 5403 231 5437
rect 265 5403 300 5437
rect 225 5364 300 5403
rect 225 5330 231 5364
rect 265 5330 300 5364
rect 225 5291 300 5330
rect 225 5257 231 5291
rect 265 5257 300 5291
rect 225 5218 300 5257
rect 225 5184 231 5218
rect 265 5184 300 5218
rect 225 5145 300 5184
rect 225 5111 231 5145
rect 265 5111 300 5145
rect 225 5072 300 5111
rect 225 5038 231 5072
rect 265 5038 300 5072
rect 225 4999 300 5038
rect 225 4965 231 4999
rect 265 4965 300 4999
rect 225 4926 300 4965
rect 225 4892 231 4926
rect 265 4892 300 4926
rect 225 4853 300 4892
rect 225 4819 231 4853
rect 265 4819 300 4853
rect 225 4780 300 4819
rect 225 4746 231 4780
rect 265 4746 300 4780
rect 225 4707 300 4746
rect 225 4673 231 4707
rect 265 4673 300 4707
rect 225 4634 300 4673
rect 225 4600 231 4634
rect 265 4600 300 4634
rect 225 4561 300 4600
rect 225 4527 231 4561
rect 265 4527 300 4561
rect 225 4488 300 4527
rect 225 4454 231 4488
rect 265 4454 300 4488
rect 225 4415 300 4454
rect 225 4381 231 4415
rect 265 4381 300 4415
rect 225 4333 300 4381
rect 225 4299 231 4333
rect 265 4299 300 4333
rect 225 4221 300 4299
rect 370 4387 428 7970
rect 497 11768 553 11769
rect 496 8282 554 11767
rect 749 11768 805 11769
rect 496 8248 508 8282
rect 542 8248 554 8282
rect 496 8210 554 8248
rect 496 8176 508 8210
rect 542 8176 554 8210
rect 496 8076 554 8176
rect 496 8042 508 8076
rect 542 8042 554 8076
rect 496 8004 554 8042
rect 496 7970 508 8004
rect 542 7970 554 8004
rect 496 7912 554 7970
rect 622 8282 680 8288
rect 622 8248 634 8282
rect 668 8248 680 8282
rect 622 8210 680 8248
rect 622 8176 634 8210
rect 668 8176 680 8210
rect 622 8076 680 8176
rect 622 8042 634 8076
rect 668 8042 680 8076
rect 622 8004 680 8042
rect 622 7970 634 8004
rect 668 7970 680 8004
rect 622 7964 680 7970
rect 748 8282 806 11767
rect 874 8380 932 11865
rect 1000 12177 1058 15662
rect 1126 12275 1184 15760
rect 1252 16072 1310 16078
rect 1252 16038 1264 16072
rect 1298 16038 1310 16072
rect 1252 16000 1310 16038
rect 1252 15966 1264 16000
rect 1298 15966 1310 16000
rect 1252 15866 1310 15966
rect 1252 15832 1264 15866
rect 1298 15832 1310 15866
rect 1252 15794 1310 15832
rect 1252 15760 1264 15794
rect 1298 15760 1310 15794
rect 1252 15754 1310 15760
rect 1378 16072 1436 16130
rect 1631 16131 1687 16132
rect 1378 16038 1390 16072
rect 1424 16038 1436 16072
rect 1378 16000 1436 16038
rect 1378 15966 1390 16000
rect 1424 15966 1436 16000
rect 1378 15866 1436 15966
rect 1378 15832 1390 15866
rect 1424 15832 1436 15866
rect 1378 15794 1436 15832
rect 1378 15760 1390 15794
rect 1424 15760 1436 15794
rect 1127 12273 1183 12274
rect 1378 12275 1436 15760
rect 1504 16072 1562 16078
rect 1504 16038 1516 16072
rect 1550 16038 1562 16072
rect 1504 16000 1562 16038
rect 1504 15966 1516 16000
rect 1550 15966 1562 16000
rect 1504 15866 1562 15966
rect 1504 15832 1516 15866
rect 1550 15832 1562 15866
rect 1504 15794 1562 15832
rect 1504 15760 1516 15794
rect 1550 15760 1562 15794
rect 1504 15754 1562 15760
rect 1630 16072 1688 16130
rect 1883 16131 1936 16132
tri 2134 16131 2135 16132 ne
rect 2135 16131 2185 16132
tri 2135 16130 2136 16131 ne
rect 2136 16130 2185 16131
rect 1882 16078 1937 16130
tri 2136 16127 2139 16130 ne
rect 2139 16127 2185 16130
tri 1937 16078 1940 16081 sw
rect 1630 16038 1642 16072
rect 1676 16038 1688 16072
rect 1630 16000 1688 16038
rect 1630 15966 1642 16000
rect 1676 15966 1688 16000
rect 1630 15866 1688 15966
rect 1630 15832 1642 15866
rect 1676 15832 1688 15866
rect 1630 15794 1688 15832
rect 1630 15760 1642 15794
rect 1676 15760 1688 15794
rect 1379 12273 1435 12274
rect 1630 12275 1688 15760
rect 1756 16072 1814 16078
rect 1756 16038 1768 16072
rect 1802 16038 1814 16072
rect 1756 16000 1814 16038
rect 1756 15966 1768 16000
rect 1802 15966 1814 16000
rect 1756 15866 1814 15966
rect 1756 15832 1768 15866
rect 1802 15832 1814 15866
rect 1756 15794 1814 15832
rect 1756 15760 1768 15794
rect 1802 15760 1814 15794
rect 1756 15754 1814 15760
rect 1882 16072 1940 16078
rect 1882 16038 1894 16072
rect 1928 16038 1940 16072
rect 1882 16000 1940 16038
rect 1882 15966 1894 16000
rect 1928 15966 1940 16000
rect 1882 15866 1940 15966
rect 1882 15832 1894 15866
rect 1928 15832 1940 15866
rect 1882 15794 1940 15832
rect 1882 15760 1894 15794
rect 1928 15760 1940 15794
rect 1882 15754 1940 15760
rect 2008 16072 2066 16078
rect 2008 16038 2020 16072
rect 2054 16038 2066 16072
rect 2008 16000 2066 16038
rect 2008 15966 2020 16000
rect 2054 15966 2066 16000
rect 2008 15866 2066 15966
rect 2008 15832 2020 15866
rect 2054 15832 2066 15866
rect 2008 15794 2066 15832
rect 2008 15760 2020 15794
rect 2054 15760 2066 15794
rect 2008 15754 2066 15760
rect 1631 12273 1687 12274
rect 1882 12275 1937 15754
tri 1937 15751 1940 15754 nw
tri 2114 15680 2139 15705 se
rect 2139 15680 2185 15705
rect 1883 12273 1936 12274
rect 1000 12143 1012 12177
rect 1046 12143 1058 12177
rect 1000 12105 1058 12143
rect 1000 12071 1012 12105
rect 1046 12071 1058 12105
rect 1000 11971 1058 12071
rect 1000 11937 1012 11971
rect 1046 11937 1058 11971
rect 1000 11899 1058 11937
rect 1000 11865 1012 11899
rect 1046 11865 1058 11899
rect 1000 11807 1058 11865
rect 1001 11805 1057 11806
rect 1127 12236 1183 12237
rect 1126 12177 1184 12235
rect 1379 12236 1435 12237
rect 1126 12143 1138 12177
rect 1172 12143 1184 12177
rect 1126 12105 1184 12143
rect 1126 12071 1138 12105
rect 1172 12071 1184 12105
rect 1126 11971 1184 12071
rect 1126 11937 1138 11971
rect 1172 11937 1184 11971
rect 1126 11899 1184 11937
rect 1126 11865 1138 11899
rect 1172 11865 1184 11899
rect 875 8378 931 8379
rect 1001 11768 1057 11769
rect 748 8248 760 8282
rect 794 8248 806 8282
rect 748 8210 806 8248
rect 748 8176 760 8210
rect 794 8176 806 8210
rect 748 8076 806 8176
rect 748 8042 760 8076
rect 794 8042 806 8076
rect 748 8004 806 8042
rect 748 7970 760 8004
rect 794 7970 806 8004
rect 497 7910 553 7911
rect 748 7912 806 7970
rect 749 7910 805 7911
rect 875 8341 931 8342
rect 874 8282 932 8340
rect 874 8248 886 8282
rect 920 8248 932 8282
rect 874 8210 932 8248
rect 874 8176 886 8210
rect 920 8176 932 8210
rect 874 8076 932 8176
rect 874 8042 886 8076
rect 920 8042 932 8076
rect 874 8004 932 8042
rect 874 7970 886 8004
rect 920 7970 932 8004
rect 370 4353 382 4387
rect 416 4353 428 4387
rect 370 4315 428 4353
rect 370 4281 382 4315
rect 416 4281 428 4315
rect 370 4275 428 4281
rect 497 7873 553 7874
rect 496 4387 554 7872
rect 749 7873 805 7874
rect 496 4353 508 4387
rect 542 4353 554 4387
rect 496 4315 554 4353
rect 496 4281 508 4315
rect 542 4281 554 4315
rect 496 4275 554 4281
rect 622 4387 680 4393
rect 622 4353 634 4387
rect 668 4353 680 4387
rect 622 4315 680 4353
rect 622 4281 634 4315
rect 668 4281 680 4315
rect 622 4275 680 4281
rect 748 4387 806 7872
rect 874 4485 932 7970
rect 1000 8282 1058 11767
rect 1126 8380 1184 11865
rect 1252 12177 1310 12183
rect 1252 12143 1264 12177
rect 1298 12143 1310 12177
rect 1252 12105 1310 12143
rect 1252 12071 1264 12105
rect 1298 12071 1310 12105
rect 1252 11971 1310 12071
rect 1252 11937 1264 11971
rect 1298 11937 1310 11971
rect 1252 11899 1310 11937
rect 1252 11865 1264 11899
rect 1298 11865 1310 11899
rect 1252 11859 1310 11865
rect 1378 12177 1436 12235
rect 1631 12236 1687 12237
rect 1378 12143 1390 12177
rect 1424 12143 1436 12177
rect 1378 12105 1436 12143
rect 1378 12071 1390 12105
rect 1424 12071 1436 12105
rect 1378 11971 1436 12071
rect 1378 11937 1390 11971
rect 1424 11937 1436 11971
rect 1378 11899 1436 11937
rect 1378 11865 1390 11899
rect 1424 11865 1436 11899
rect 1127 8378 1183 8379
rect 1378 8380 1436 11865
rect 1504 12177 1562 12183
rect 1504 12143 1516 12177
rect 1550 12143 1562 12177
rect 1504 12105 1562 12143
rect 1504 12071 1516 12105
rect 1550 12071 1562 12105
rect 1504 11971 1562 12071
rect 1504 11937 1516 11971
rect 1550 11937 1562 11971
rect 1504 11899 1562 11937
rect 1504 11865 1516 11899
rect 1550 11865 1562 11899
rect 1504 11859 1562 11865
rect 1630 12177 1688 12235
rect 1883 12236 1936 12237
rect 1882 12183 1937 12235
rect 2017 12224 2185 15680
tri 2114 12199 2139 12224 ne
rect 2139 12199 2185 12224
tri 1937 12183 1940 12186 sw
rect 1630 12143 1642 12177
rect 1676 12143 1688 12177
rect 1630 12105 1688 12143
rect 1630 12071 1642 12105
rect 1676 12071 1688 12105
rect 1630 11971 1688 12071
rect 1630 11937 1642 11971
rect 1676 11937 1688 11971
rect 1630 11899 1688 11937
rect 1630 11865 1642 11899
rect 1676 11865 1688 11899
rect 1379 8378 1435 8379
rect 1630 8380 1688 11865
rect 1756 12177 1814 12183
rect 1756 12143 1768 12177
rect 1802 12143 1814 12177
rect 1756 12105 1814 12143
rect 1756 12071 1768 12105
rect 1802 12071 1814 12105
rect 1756 11971 1814 12071
rect 1756 11937 1768 11971
rect 1802 11937 1814 11971
rect 1756 11899 1814 11937
rect 1756 11865 1768 11899
rect 1802 11865 1814 11899
rect 1756 11859 1814 11865
rect 1882 12177 1940 12183
rect 1882 12143 1894 12177
rect 1928 12143 1940 12177
rect 1882 12105 1940 12143
rect 1882 12071 1894 12105
rect 1928 12071 1940 12105
rect 1882 11971 1940 12071
rect 1882 11937 1894 11971
rect 1928 11937 1940 11971
rect 1882 11899 1940 11937
rect 1882 11865 1894 11899
rect 1928 11865 1940 11899
rect 1882 11859 1940 11865
rect 2008 12177 2066 12183
rect 2008 12143 2020 12177
rect 2054 12143 2066 12177
rect 2008 12105 2066 12143
rect 2008 12071 2020 12105
rect 2054 12071 2066 12105
rect 2008 11971 2066 12071
rect 2008 11937 2020 11971
rect 2054 11937 2066 11971
rect 2008 11899 2066 11937
rect 2008 11865 2020 11899
rect 2054 11865 2066 11899
rect 2008 11859 2066 11865
rect 1631 8378 1687 8379
rect 1882 8380 1937 11859
tri 1937 11856 1940 11859 nw
tri 2017 11721 2139 11843 se
rect 2139 11721 2185 11843
tri 1992 10410 2017 10435 se
rect 1883 8378 1936 8379
rect 2017 8362 2185 11721
rect 2231 10992 2283 27578
rect 2328 27550 2373 27637
rect 2325 11038 2377 22742
tri 2283 10992 2308 11017 sw
rect 2231 10941 6806 10992
tri 6729 10913 6757 10941 ne
rect 6757 10913 6806 10941
rect 2734 10907 6706 10913
rect 2734 10895 3015 10907
rect 1000 8248 1012 8282
rect 1046 8248 1058 8282
rect 1000 8210 1058 8248
rect 1000 8176 1012 8210
rect 1046 8176 1058 8210
rect 1000 8076 1058 8176
rect 1000 8042 1012 8076
rect 1046 8042 1058 8076
rect 1000 8004 1058 8042
rect 1000 7970 1012 8004
rect 1046 7970 1058 8004
rect 1000 7912 1058 7970
rect 1001 7910 1057 7911
rect 1127 8341 1183 8342
rect 1126 8282 1184 8340
rect 1379 8341 1435 8342
rect 1126 8248 1138 8282
rect 1172 8248 1184 8282
rect 1126 8210 1184 8248
rect 1126 8176 1138 8210
rect 1172 8176 1184 8210
rect 1126 8076 1184 8176
rect 1126 8042 1138 8076
rect 1172 8042 1184 8076
rect 1126 8004 1184 8042
rect 1126 7970 1138 8004
rect 1172 7970 1184 8004
rect 875 4483 931 4484
rect 1001 7873 1057 7874
rect 748 4353 760 4387
rect 794 4353 806 4387
rect 748 4315 806 4353
rect 748 4281 760 4315
rect 794 4281 806 4315
rect 748 4275 806 4281
rect 875 4446 931 4447
rect 874 4387 932 4445
rect 874 4353 886 4387
rect 920 4353 932 4387
rect 874 4315 932 4353
rect 874 4281 886 4315
rect 920 4281 932 4315
rect 874 4275 932 4281
rect 1000 4387 1058 7872
rect 1126 4504 1184 7970
rect 1252 8282 1310 8288
rect 1252 8248 1264 8282
rect 1298 8248 1310 8282
rect 1252 8210 1310 8248
rect 1252 8176 1264 8210
rect 1298 8176 1310 8210
rect 1252 8076 1310 8176
rect 1252 8042 1264 8076
rect 1298 8042 1310 8076
rect 1252 8004 1310 8042
rect 1252 7970 1264 8004
rect 1298 7970 1310 8004
rect 1252 7964 1310 7970
rect 1378 8282 1436 8340
rect 1631 8341 1687 8342
rect 1378 8248 1390 8282
rect 1424 8248 1436 8282
rect 1378 8210 1436 8248
rect 1378 8176 1390 8210
rect 1424 8176 1436 8210
rect 1378 8076 1436 8176
rect 1378 8042 1390 8076
rect 1424 8042 1436 8076
rect 1378 8004 1436 8042
rect 1378 7970 1390 8004
rect 1424 7970 1436 8004
rect 1252 4644 1310 4650
rect 1252 4610 1264 4644
rect 1298 4610 1310 4644
rect 1252 4572 1310 4610
rect 1252 4538 1264 4572
rect 1298 4538 1310 4572
rect 1252 4532 1310 4538
tri 1184 4504 1209 4529 sw
rect 1378 4505 1436 7970
rect 1504 8282 1562 8288
rect 1504 8248 1516 8282
rect 1550 8248 1562 8282
rect 1504 8210 1562 8248
rect 1504 8176 1516 8210
rect 1550 8176 1562 8210
rect 1504 8076 1562 8176
rect 1504 8042 1516 8076
rect 1550 8042 1562 8076
rect 1504 8004 1562 8042
rect 1504 7970 1516 8004
rect 1550 7970 1562 8004
rect 1504 7964 1562 7970
rect 1630 8282 1688 8340
rect 1883 8341 1936 8342
rect 1882 8288 1937 8340
rect 2045 8328 2279 8334
tri 1937 8288 1940 8291 sw
rect 1630 8248 1642 8282
rect 1676 8248 1688 8282
rect 1630 8210 1688 8248
rect 1630 8176 1642 8210
rect 1676 8176 1688 8210
rect 1630 8076 1688 8176
rect 1756 8282 1814 8288
rect 1756 8248 1768 8282
rect 1802 8248 1814 8282
rect 1756 8210 1814 8248
rect 1756 8176 1768 8210
rect 1802 8176 1814 8210
rect 1756 8170 1814 8176
rect 1882 8282 1940 8288
rect 1882 8248 1894 8282
rect 1928 8248 1940 8282
rect 1882 8210 1940 8248
rect 1882 8176 1894 8210
rect 1928 8176 1940 8210
rect 2097 8276 2279 8328
rect 2045 8264 2279 8276
rect 2097 8212 2279 8264
rect 2045 8206 2279 8212
rect 1882 8170 1940 8176
tri 1874 8150 1882 8158 se
rect 1882 8150 1937 8170
tri 1937 8167 1940 8170 nw
tri 2180 8167 2219 8206 ne
rect 2219 8167 2279 8206
tri 2219 8155 2231 8167 ne
tri 1853 8129 1874 8150 se
rect 1874 8129 1937 8150
tri 1814 8090 1853 8129 se
rect 1853 8090 1898 8129
tri 1898 8090 1937 8129 nw
rect 1965 8144 2139 8150
rect 2017 8092 2139 8144
tri 1806 8082 1814 8090 se
rect 1814 8082 1890 8090
tri 1890 8082 1898 8090 nw
rect 1630 8042 1642 8076
rect 1676 8042 1688 8076
rect 1630 8004 1688 8042
rect 1630 7970 1642 8004
rect 1676 7970 1688 8004
rect 1126 4503 1257 4504
tri 1257 4503 1258 4504 sw
rect 1379 4503 1435 4504
rect 1630 5350 1688 7970
tri 1756 8032 1806 8082 se
rect 1806 8032 1830 8082
rect 1756 8022 1830 8032
tri 1830 8022 1890 8082 nw
rect 1965 8080 2139 8092
rect 2017 8028 2029 8080
rect 2081 8028 2139 8080
rect 1965 8022 2139 8028
rect 1756 5424 1814 8022
tri 1814 8006 1830 8022 nw
tri 2100 8006 2116 8022 ne
rect 2116 8006 2139 8022
tri 2116 7994 2128 8006 ne
rect 2128 7994 2139 8006
rect 1882 7988 2066 7994
rect 1882 7954 1894 7988
rect 1928 7954 2066 7988
tri 2128 7983 2139 7994 ne
rect 1882 7916 2066 7954
rect 1882 7882 1894 7916
rect 1928 7882 2066 7916
rect 1882 7876 2066 7882
tri 1983 7851 2008 7876 ne
tri 1998 5588 2008 5598 se
rect 2008 5588 2066 7876
rect 2231 6373 2279 8167
rect 2325 6409 2594 10889
rect 2734 10849 2820 10895
rect 2961 10855 3015 10878
rect 3067 10855 3079 10907
rect 3131 10855 3143 10907
rect 3195 10855 3207 10907
rect 3259 10895 3429 10907
rect 3259 10855 3429 10878
rect 3481 10855 3493 10907
rect 3545 10855 3557 10907
rect 3609 10855 3621 10907
rect 3673 10855 3685 10907
rect 3737 10855 3749 10907
rect 3801 10895 3973 10907
rect 3801 10855 3973 10878
rect 4025 10855 4037 10907
rect 4089 10855 4101 10907
rect 4153 10855 4165 10907
rect 4217 10855 4229 10907
rect 4281 10855 4293 10907
rect 4345 10855 4357 10907
rect 4409 10895 5109 10907
rect 2961 10849 4409 10855
rect 5081 10855 5109 10878
rect 5161 10855 5173 10907
rect 5225 10855 5237 10907
rect 5289 10855 5301 10907
rect 5353 10855 5365 10907
rect 5417 10855 5429 10907
rect 5481 10895 5637 10907
rect 5481 10855 5637 10878
rect 5689 10855 5701 10907
rect 5753 10855 5765 10907
rect 5817 10855 5829 10907
rect 5881 10855 5893 10907
rect 5945 10855 5957 10907
rect 6009 10855 6021 10907
rect 6073 10895 6269 10907
rect 6073 10855 6269 10878
rect 6321 10855 6333 10907
rect 6385 10855 6397 10907
rect 6449 10855 6461 10907
rect 6513 10855 6525 10907
rect 6577 10855 6589 10907
rect 6641 10855 6653 10907
rect 6705 10905 6706 10907
tri 6706 10905 6714 10913 sw
tri 6757 10905 6765 10913 ne
rect 6705 10882 6714 10905
tri 6714 10882 6737 10905 sw
rect 6705 10855 6737 10882
rect 5081 10849 6737 10855
rect 2734 10846 2826 10849
rect 2737 6597 2826 10846
tri 2826 10824 2851 10849 nw
tri 2936 10824 2961 10849 ne
rect 2961 10826 4363 10849
tri 4363 10826 4386 10849 nw
tri 4615 10826 4638 10849 ne
rect 4638 10826 4802 10849
rect 4361 10825 4362 10826
tri 4362 10825 4363 10826 nw
tri 4638 10825 4639 10826 ne
rect 4639 10825 4802 10826
rect 2962 10824 4360 10825
tri 4361 10824 4362 10825 nw
tri 4639 10824 4640 10825 ne
tri 2936 10763 2961 10788 se
rect 2962 10787 4360 10788
tri 4361 10787 4362 10788 sw
tri 4467 10787 4468 10788 se
rect 4468 10787 4474 10788
rect 4361 10786 4362 10787
tri 4362 10786 4363 10787 sw
tri 4466 10786 4467 10787 se
rect 4467 10786 4474 10787
rect 2961 10763 4363 10786
tri 4363 10763 4386 10786 sw
tri 4443 10763 4466 10786 se
rect 4466 10763 4474 10786
rect 2961 10717 4394 10763
rect 4396 10762 4432 10763
rect 2936 10711 4394 10717
rect 4395 10712 4433 10762
rect 4396 10711 4432 10712
rect 4434 10711 4474 10763
tri 2936 10686 2961 10711 ne
rect 2961 10688 4363 10711
tri 4363 10688 4386 10711 nw
tri 4443 10688 4466 10711 ne
rect 4466 10688 4474 10711
rect 4361 10687 4362 10688
tri 4362 10687 4363 10688 nw
tri 4466 10687 4467 10688 ne
rect 4467 10687 4474 10688
rect 2962 10686 4360 10687
tri 4361 10686 4362 10687 nw
tri 4467 10686 4468 10687 ne
rect 4468 10672 4474 10687
rect 4590 10672 4596 10788
tri 2936 10625 2961 10650 se
rect 2962 10649 4360 10650
tri 4361 10649 4362 10650 sw
rect 4361 10648 4362 10649
tri 4362 10648 4363 10649 sw
rect 2961 10625 4363 10648
tri 4363 10625 4386 10648 sw
rect 2734 6419 2826 6597
rect 2854 10425 4612 10625
rect 2854 8920 3041 10425
tri 3041 10283 3183 10425 nw
tri 3436 10283 3578 10425 ne
tri 3041 8920 3183 9062 sw
tri 3436 8920 3578 9062 se
rect 3578 8920 3892 10425
tri 3892 10283 4034 10425 nw
tri 4287 10283 4429 10425 ne
tri 3892 8920 4034 9062 sw
tri 4287 8920 4429 9062 se
rect 4429 8920 4612 10425
rect 2854 8677 4612 8920
rect 2855 8675 4611 8676
rect 2854 8639 4612 8675
rect 2855 8638 4611 8639
rect 2854 8394 4612 8637
rect 2854 8378 3167 8394
tri 3167 8378 3183 8394 nw
tri 3436 8378 3452 8394 ne
rect 3452 8378 4018 8394
tri 4018 8378 4034 8394 nw
tri 4287 8378 4303 8394 ne
rect 4303 8378 4612 8394
rect 2854 8342 3131 8378
tri 3131 8342 3167 8378 nw
tri 3452 8342 3488 8378 ne
rect 3488 8342 3982 8378
tri 3982 8342 4018 8378 nw
tri 4303 8342 4339 8378 ne
rect 4339 8342 4612 8378
rect 2854 8334 3123 8342
tri 3123 8334 3131 8342 nw
tri 3488 8334 3496 8342 ne
rect 3496 8334 3974 8342
tri 3974 8334 3982 8342 nw
tri 4339 8334 4347 8342 ne
rect 4347 8334 4612 8342
rect 2854 6889 3041 8334
tri 3041 8252 3123 8334 nw
tri 3496 8252 3578 8334 ne
tri 3041 6889 3183 7031 sw
tri 3436 6889 3578 7031 se
rect 3578 6889 3892 8334
tri 3892 8252 3974 8334 nw
tri 4347 8252 4429 8334 ne
tri 3892 6889 4034 7031 sw
tri 4287 6889 4429 7031 se
rect 4429 6889 4612 8334
rect 2854 6689 4612 6889
rect 2854 6666 3023 6689
tri 3023 6666 3046 6689 nw
tri 3080 6666 3103 6689 ne
rect 3103 6666 4363 6689
tri 4363 6666 4386 6689 nw
rect 3021 6665 3022 6666
tri 3022 6665 3023 6666 nw
tri 3103 6665 3104 6666 ne
rect 3104 6665 3105 6666
rect 4361 6665 4362 6666
tri 4362 6665 4363 6666 nw
rect 2855 6664 3020 6665
tri 3021 6664 3022 6665 nw
tri 3104 6664 3105 6665 ne
rect 3106 6664 4360 6665
tri 4361 6664 4362 6665 nw
rect 2854 6628 3021 6664
rect 2855 6627 3020 6628
tri 3104 6627 3105 6628 se
rect 3106 6627 4360 6628
tri 4361 6627 4362 6628 sw
tri 4467 6627 4468 6628 se
rect 4468 6627 4474 6642
tri 3103 6626 3104 6627 se
rect 3104 6626 3105 6627
rect 4361 6626 4362 6627
tri 4362 6626 4363 6627 sw
tri 4466 6626 4467 6627 se
rect 4467 6626 4474 6627
rect 2854 6548 3021 6626
tri 3080 6603 3103 6626 se
rect 3103 6603 4363 6626
tri 4363 6603 4386 6626 sw
tri 4443 6603 4466 6626 se
rect 4466 6603 4474 6626
rect 3080 6597 4394 6603
rect 4396 6602 4432 6603
rect 3105 6551 4394 6597
rect 4395 6552 4433 6602
rect 4396 6551 4432 6552
rect 4434 6551 4474 6603
tri 3080 6548 3083 6551 ne
rect 3083 6548 4363 6551
rect 2854 6496 2906 6548
rect 2958 6496 3021 6548
tri 3083 6526 3105 6548 ne
rect 3105 6528 4363 6548
tri 4363 6528 4386 6551 nw
tri 4443 6528 4466 6551 ne
rect 4466 6528 4474 6551
rect 4361 6527 4362 6528
tri 4362 6527 4363 6528 nw
tri 4466 6527 4467 6528 ne
rect 4467 6527 4474 6528
rect 3106 6526 4360 6527
tri 4361 6526 4362 6527 nw
tri 4467 6526 4468 6527 ne
rect 4468 6526 4474 6527
rect 4590 6526 4596 6642
rect 2854 6484 3021 6496
rect 2854 6432 2906 6484
rect 2958 6432 3021 6484
tri 3080 6465 3105 6490 se
rect 3106 6489 4360 6490
tri 4361 6489 4362 6490 sw
tri 4639 6489 4640 6490 se
rect 4640 6489 4802 10825
tri 4802 10824 4827 10849 nw
tri 5056 10824 5081 10849 ne
rect 5081 10826 6483 10849
tri 6483 10826 6506 10849 nw
tri 6591 10826 6614 10849 ne
rect 6614 10826 6737 10849
rect 6481 10825 6482 10826
tri 6482 10825 6483 10826 nw
tri 6614 10825 6615 10826 ne
rect 6615 10825 6737 10826
rect 5082 10824 6480 10825
tri 6481 10824 6482 10825 nw
tri 6615 10824 6616 10825 ne
rect 4840 10672 4846 10788
rect 4962 10763 4968 10788
tri 4968 10763 4993 10788 sw
tri 5056 10763 5081 10788 se
rect 5082 10787 6480 10788
tri 6481 10787 6482 10788 sw
rect 6481 10786 6482 10787
tri 6482 10786 6483 10787 sw
rect 5081 10763 6483 10786
tri 6483 10763 6506 10786 sw
rect 4962 10711 5008 10763
rect 5010 10762 5046 10763
rect 5009 10712 5047 10762
rect 5048 10717 6481 10763
rect 5010 10711 5046 10712
rect 5048 10711 6506 10717
rect 4962 10672 4968 10711
tri 4968 10686 4993 10711 nw
tri 5056 10686 5081 10711 ne
rect 5081 10688 6483 10711
tri 6483 10688 6506 10711 nw
rect 6481 10687 6482 10688
tri 6482 10687 6483 10688 nw
rect 5082 10686 6480 10687
tri 6481 10686 6482 10687 nw
tri 5056 10625 5081 10650 se
rect 5082 10649 6480 10650
tri 6481 10649 6482 10650 sw
rect 6481 10648 6482 10649
tri 6482 10648 6483 10649 sw
rect 5081 10625 6483 10648
tri 6483 10625 6506 10648 sw
rect 4830 10425 6588 10625
rect 4830 8920 5013 10425
tri 5013 10283 5155 10425 nw
tri 5408 10283 5550 10425 ne
tri 5013 8920 5155 9062 sw
tri 5408 8920 5550 9062 se
rect 5550 8920 5864 10425
tri 5864 10283 6006 10425 nw
tri 6259 10283 6401 10425 ne
tri 5864 8920 6006 9062 sw
tri 6259 8920 6401 9062 se
rect 6401 8920 6588 10425
rect 4830 8677 6588 8920
rect 4831 8675 6587 8676
rect 4830 8639 6588 8675
rect 4831 8638 6587 8639
rect 4830 8394 6588 8637
rect 4830 6889 5013 8394
tri 5013 8252 5155 8394 nw
tri 5408 8252 5550 8394 ne
tri 5013 6889 5155 7031 sw
tri 5408 6889 5550 7031 se
rect 5550 6889 5864 8394
tri 5864 8252 6006 8394 nw
tri 6259 8252 6401 8394 ne
tri 5864 6889 6006 7031 sw
tri 6259 6889 6401 7031 se
rect 6401 6889 6588 8394
rect 4830 6689 6588 6889
tri 5056 6664 5081 6689 ne
rect 5081 6666 6339 6689
tri 6339 6666 6362 6689 nw
tri 6396 6666 6419 6689 ne
rect 6419 6666 6588 6689
rect 6337 6665 6338 6666
tri 6338 6665 6339 6666 nw
tri 6419 6665 6420 6666 ne
rect 6420 6665 6421 6666
rect 5082 6664 6336 6665
tri 6337 6664 6338 6665 nw
tri 6420 6664 6421 6665 ne
rect 6422 6664 6587 6665
rect 4840 6526 4846 6642
rect 4962 6603 4968 6642
rect 6421 6628 6588 6664
tri 4968 6603 4993 6628 sw
tri 5056 6603 5081 6628 se
rect 5082 6627 6336 6628
tri 6337 6627 6338 6628 sw
rect 6422 6627 6587 6628
rect 6337 6626 6338 6627
tri 6338 6626 6339 6627 sw
rect 5081 6603 6339 6626
tri 6339 6603 6362 6626 sw
rect 4962 6551 5008 6603
rect 5010 6602 5046 6603
rect 5009 6552 5047 6602
rect 5048 6597 6362 6603
rect 5010 6551 5046 6552
rect 5048 6551 6337 6597
rect 4962 6526 4968 6551
tri 4968 6526 4993 6551 nw
tri 5056 6526 5081 6551 ne
rect 5081 6528 6339 6551
tri 6339 6528 6362 6551 nw
rect 6337 6527 6338 6528
tri 6338 6527 6339 6528 nw
rect 5082 6526 6336 6527
tri 6337 6526 6338 6527 nw
rect 4361 6488 4362 6489
tri 4362 6488 4363 6489 sw
tri 4638 6488 4639 6489 se
rect 4639 6488 4802 6489
rect 3105 6465 4363 6488
tri 4363 6465 4386 6488 sw
tri 4615 6465 4638 6488 se
rect 4638 6465 4802 6488
tri 4802 6465 4827 6490 sw
tri 5056 6465 5081 6490 se
rect 5082 6489 6336 6490
tri 6337 6489 6338 6490 sw
rect 6337 6488 6338 6489
tri 6338 6488 6339 6489 sw
rect 5081 6465 6339 6488
tri 6339 6465 6362 6488 sw
rect 3105 6459 4409 6465
rect 3105 6436 3143 6459
rect 3063 6407 3143 6419
rect 3195 6407 3207 6459
rect 3259 6436 3424 6459
rect 3259 6407 3424 6419
rect 3476 6407 3488 6459
rect 3540 6407 3552 6459
rect 3604 6407 3616 6459
rect 3668 6436 3973 6459
rect 3668 6407 3973 6419
rect 4025 6407 4037 6459
rect 4089 6407 4101 6459
rect 4153 6407 4165 6459
rect 4217 6407 4229 6459
rect 4281 6407 4293 6459
rect 4345 6407 4357 6459
rect 5081 6459 6337 6465
rect 5081 6436 5109 6459
rect 4409 6407 5109 6419
rect 5161 6407 5173 6459
rect 5225 6407 5237 6459
rect 5289 6407 5301 6459
rect 5353 6436 5777 6459
rect 5353 6419 5403 6436
rect 5353 6407 5777 6419
rect 5829 6407 5841 6459
rect 5893 6407 5905 6459
rect 5957 6407 5969 6459
rect 6021 6407 6033 6459
rect 6085 6436 6337 6459
tri 6408 6419 6421 6432 se
rect 6421 6419 6588 6626
rect 6616 6588 6737 10825
rect 6765 10709 6806 10913
tri 6806 10709 6831 10734 sw
rect 6765 10658 7306 10709
rect 6848 8206 7083 10630
tri 7083 8206 7186 8309 sw
rect 6848 8167 7186 8206
tri 7186 8167 7225 8206 sw
rect 6848 7952 7306 8167
rect 6848 7876 7149 7952
tri 7149 7876 7225 7952 nw
rect 6848 7424 7083 7876
tri 7083 7810 7149 7876 nw
tri 7083 7424 7225 7566 sw
rect 6848 7148 7306 7424
rect 6848 6662 7083 7148
tri 7083 7006 7225 7148 nw
rect 6085 6407 6350 6419
rect 3063 6401 6350 6407
tri 6350 6401 6368 6419 nw
tri 6390 6401 6408 6419 se
rect 6408 6401 6588 6419
tri 6371 6382 6390 6401 se
rect 6390 6382 6588 6401
tri 2279 6373 2288 6382 sw
tri 6362 6373 6371 6382 se
rect 6371 6373 6588 6382
rect 2231 6357 2288 6373
tri 2288 6357 2304 6373 sw
rect 2231 6341 5506 6357
tri 5506 6341 5522 6357 sw
rect 2231 6321 5522 6341
tri 5522 6321 5542 6341 sw
rect 5594 6321 5600 6373
rect 5652 6321 5664 6373
rect 5716 6321 6588 6373
tri 6737 6321 6773 6357 se
rect 6773 6321 7306 6357
rect 2231 6309 5542 6321
tri 5483 6276 5516 6309 ne
rect 5516 6286 5542 6309
tri 5542 6286 5577 6321 sw
tri 5594 6298 5617 6321 ne
rect 5617 6298 6588 6321
tri 6714 6298 6737 6321 se
rect 6737 6309 7306 6321
rect 6737 6298 6773 6309
tri 6702 6286 6714 6298 se
rect 6714 6286 6773 6298
tri 6773 6286 6796 6309 nw
rect 5516 6276 5577 6286
tri 5577 6276 5587 6286 sw
tri 6692 6276 6702 6286 se
rect 6702 6276 6757 6286
rect 2325 6264 4393 6276
tri 5516 6270 5522 6276 ne
rect 5522 6270 5587 6276
tri 5587 6270 5593 6276 sw
tri 6686 6270 6692 6276 se
rect 6692 6270 6757 6276
tri 6757 6270 6773 6286 nw
rect 2325 6230 2334 6264
rect 2368 6230 4393 6264
tri 5522 6230 5562 6270 ne
rect 5562 6230 6709 6270
rect 2325 6229 2445 6230
rect 2377 6177 2445 6229
rect 2325 6165 2334 6177
rect 2368 6165 2445 6177
rect 2377 6159 2445 6165
tri 2445 6159 2516 6230 nw
tri 5562 6222 5570 6230 ne
rect 5570 6222 6709 6230
tri 6709 6222 6757 6270 nw
rect 2377 6113 2393 6159
rect 2325 6107 2393 6113
tri 2393 6107 2445 6159 nw
rect 2507 6107 2513 6159
rect 2565 6107 2577 6159
rect 2629 6107 6259 6159
rect 6311 6107 6323 6159
rect 6375 6107 7306 6159
rect 4996 6069 5048 6075
tri 4971 5999 4996 6024 se
rect 5321 6027 5327 6079
rect 5379 6027 5391 6079
rect 5443 6027 7306 6079
rect 4996 6005 5048 6017
rect 2488 5947 2494 5999
rect 2546 5953 4996 5999
tri 5048 5999 5073 6024 sw
rect 5048 5993 6000 5999
rect 5048 5959 5465 5993
rect 5499 5959 5537 5993
rect 5571 5959 6000 5993
rect 5048 5953 6000 5959
rect 2546 5947 6000 5953
rect 6052 5947 6064 5999
rect 6116 5947 7306 5999
rect 2488 5935 2552 5947
rect 2488 5883 2494 5935
rect 2546 5883 2552 5935
tri 2552 5922 2577 5947 nw
rect 3023 5861 3029 5913
rect 3081 5867 3087 5913
tri 3087 5867 3090 5870 sw
rect 5000 5867 5006 5919
rect 5058 5867 5070 5919
rect 5122 5873 7306 5919
rect 5122 5867 5128 5873
tri 5128 5867 5134 5873 nw
rect 3081 5861 3090 5867
rect 3023 5849 3090 5861
rect 3023 5797 3029 5849
rect 3081 5845 3090 5849
tri 3090 5845 3112 5867 sw
rect 3081 5839 4982 5845
tri 4982 5839 4988 5845 sw
tri 5140 5839 5146 5845 se
rect 5146 5839 5614 5845
rect 3081 5797 5614 5839
tri 5604 5793 5608 5797 ne
rect 5608 5793 5614 5797
rect 5666 5793 5678 5845
rect 5730 5793 5736 5845
rect 3240 5682 3246 5734
rect 3298 5682 3310 5734
rect 3362 5682 5682 5734
rect 2382 5654 2500 5666
tri 2500 5654 2512 5666 sw
rect 2382 5620 2388 5654
rect 2422 5620 2460 5654
rect 2494 5620 5682 5654
rect 2382 5608 5682 5620
tri 2185 5588 2202 5605 sw
tri 1984 5574 1998 5588 se
rect 1998 5574 2066 5588
tri 1980 5570 1984 5574 se
rect 1984 5570 2066 5574
rect 1882 5564 1940 5570
rect 1882 5530 1894 5564
rect 1928 5530 1940 5564
rect 1882 5492 1940 5530
rect 1882 5458 1894 5492
rect 1928 5458 1940 5492
rect 1882 5452 1940 5458
rect 1941 5453 1942 5569
rect 1978 5453 1979 5569
rect 1980 5564 2066 5570
rect 1980 5530 2020 5564
rect 2054 5530 2066 5564
rect 2139 5580 2202 5588
tri 2202 5580 2210 5588 sw
rect 2139 5574 2500 5580
rect 2139 5540 2230 5574
rect 2264 5540 2302 5574
rect 2336 5540 2500 5574
rect 2139 5534 2500 5540
rect 3134 5574 3596 5580
rect 3134 5534 3144 5574
rect 1980 5492 2066 5530
tri 3117 5507 3144 5534 ne
rect 1980 5458 2020 5492
rect 2054 5458 2066 5492
rect 1980 5452 2066 5458
rect 3260 5534 3596 5574
rect 3260 5510 3572 5534
tri 3572 5510 3596 5534 nw
rect 5608 5574 5685 5580
rect 5660 5534 5685 5574
rect 5608 5510 5660 5522
rect 3260 5498 3571 5510
tri 3571 5509 3572 5510 nw
rect 3260 5464 3531 5498
rect 3565 5464 3571 5498
rect 3260 5458 3571 5464
rect 3144 5452 3571 5458
rect 4950 5492 5224 5498
rect 4950 5458 4962 5492
rect 4996 5458 5034 5492
rect 5068 5458 5106 5492
rect 5140 5458 5178 5492
rect 5212 5458 5224 5492
rect 4950 5452 5224 5458
tri 5660 5509 5685 5534 nw
rect 5608 5452 5660 5458
tri 4800 5449 4803 5452 ne
rect 4803 5449 4866 5452
tri 4866 5449 4869 5452 sw
tri 5158 5449 5161 5452 ne
rect 5161 5449 5224 5452
tri 5224 5449 5227 5452 sw
tri 1814 5424 1839 5449 sw
tri 4803 5424 4828 5449 ne
rect 4828 5424 4869 5449
tri 4869 5424 4894 5449 sw
tri 5161 5424 5186 5449 ne
rect 5186 5424 5227 5449
tri 5227 5424 5252 5449 sw
rect 1756 5408 4776 5424
tri 4776 5408 4792 5424 sw
tri 4828 5416 4836 5424 ne
rect 4836 5416 4894 5424
tri 4894 5416 4902 5424 sw
tri 5186 5416 5194 5424 ne
rect 5194 5416 5682 5424
tri 4836 5408 4844 5416 ne
rect 4844 5408 4902 5416
tri 4902 5408 4910 5416 sw
tri 5194 5408 5202 5416 ne
rect 5202 5408 5682 5416
rect 1756 5400 4792 5408
tri 4792 5400 4800 5408 sw
tri 4844 5400 4852 5408 ne
rect 4852 5400 4910 5408
rect 1756 5386 4800 5400
tri 4800 5386 4814 5400 sw
tri 4852 5386 4866 5400 ne
rect 4866 5386 4910 5400
rect 1756 5378 4814 5386
tri 4756 5375 4759 5378 ne
rect 4759 5375 4814 5378
tri 1688 5350 1713 5375 sw
tri 4759 5350 4784 5375 ne
rect 4784 5350 4814 5375
rect 1630 5342 4729 5350
tri 4729 5342 4737 5350 sw
tri 4784 5342 4792 5350 ne
rect 4792 5342 4814 5350
tri 4814 5342 4858 5386 sw
tri 4866 5350 4902 5386 ne
rect 4902 5350 4910 5386
tri 4910 5350 4968 5408 sw
tri 5202 5386 5224 5408 ne
rect 5224 5386 5682 5408
tri 5224 5378 5232 5386 ne
rect 5232 5378 5682 5386
tri 4902 5342 4910 5350 ne
rect 4910 5342 5682 5350
rect 1630 5304 4737 5342
rect 1630 5299 1708 5304
tri 1708 5299 1713 5304 nw
tri 3773 5299 3778 5304 ne
rect 3778 5299 3864 5304
tri 3864 5299 3869 5304 nw
tri 4085 5299 4090 5304 ne
rect 4090 5299 4176 5304
tri 4176 5299 4181 5304 nw
tri 4397 5299 4402 5304 ne
rect 4402 5299 4488 5304
tri 4488 5299 4493 5304 nw
tri 4709 5299 4714 5304 ne
rect 4714 5299 4737 5304
tri 4737 5299 4780 5342 sw
rect 1630 4505 1688 5299
tri 1688 5279 1708 5299 nw
tri 3778 5279 3798 5299 ne
rect 1631 4503 1687 4504
rect 1882 5270 1940 5276
rect 1882 5236 1894 5270
rect 1928 5236 1940 5270
rect 1882 5198 1940 5236
rect 1882 5164 1894 5198
rect 1928 5164 1940 5198
rect 1126 4485 1258 4503
tri 1258 4485 1276 4503 sw
rect 1126 4467 1276 4485
tri 1276 4467 1294 4485 sw
rect 1126 4458 1294 4467
rect 1126 4453 1204 4458
tri 1204 4453 1209 4458 nw
tri 1237 4453 1242 4458 ne
rect 1242 4453 1294 4458
tri 1294 4453 1308 4467 sw
rect 1126 4433 1184 4453
tri 1184 4433 1204 4453 nw
tri 1242 4438 1257 4453 ne
rect 1257 4438 1308 4453
tri 1257 4433 1262 4438 ne
rect 1127 4431 1183 4432
rect 1000 4353 1012 4387
rect 1046 4353 1058 4387
rect 1000 4315 1058 4353
rect 1000 4281 1012 4315
rect 1046 4281 1058 4315
rect 1000 4275 1058 4281
rect 1127 4394 1183 4395
rect 1126 4387 1184 4393
rect 1126 4353 1138 4387
rect 1172 4353 1184 4387
rect 1126 4315 1184 4353
rect 1126 4281 1138 4315
rect 1172 4281 1184 4315
rect 1126 4221 1184 4281
rect 1262 4275 1308 4438
rect 1379 4466 1435 4467
rect 1378 4407 1436 4465
rect 1631 4466 1687 4467
rect 1378 4373 1390 4407
rect 1424 4373 1436 4407
rect 1378 4335 1436 4373
rect 1378 4301 1390 4335
rect 1424 4301 1436 4335
rect 1378 4295 1436 4301
rect 1504 4407 1562 4413
rect 1504 4373 1516 4407
rect 1550 4373 1562 4407
rect 1504 4335 1562 4373
rect 1504 4301 1516 4335
rect 1550 4301 1562 4335
rect 1504 4295 1562 4301
rect 1630 4407 1688 4465
rect 1630 4373 1642 4407
rect 1676 4373 1688 4407
rect 1630 4335 1688 4373
rect 1630 4301 1642 4335
rect 1676 4301 1688 4335
rect 1630 4295 1688 4301
rect 1756 4407 1814 4413
rect 1756 4373 1768 4407
rect 1802 4373 1814 4407
rect 1756 4335 1814 4373
rect 1756 4301 1768 4335
rect 1802 4301 1814 4335
rect 1756 4295 1814 4301
rect 1882 4407 1940 5164
rect 1882 4373 1894 4407
rect 1928 4373 1940 4407
rect 1882 4335 1940 4373
rect 1882 4301 1894 4335
rect 1928 4301 1940 4335
rect 1882 4295 1940 4301
rect 2008 5270 2066 5276
rect 2008 5236 2020 5270
rect 2054 5236 2066 5270
rect 2008 5198 2066 5236
rect 2008 5164 2020 5198
rect 2054 5164 2066 5198
rect 2008 4407 2066 5164
rect 2134 5270 2318 5276
rect 2134 5236 2146 5270
rect 2180 5236 2272 5270
rect 2306 5236 2318 5270
rect 2134 5198 2318 5236
rect 2134 5164 2146 5198
rect 2180 5164 2272 5198
rect 2306 5164 2318 5198
rect 2134 5158 2318 5164
rect 2134 5091 2184 5158
tri 2184 5133 2209 5158 nw
tri 2243 5133 2268 5158 ne
tri 2184 5091 2192 5099 sw
rect 2134 4505 2192 5091
rect 2135 4503 2191 4504
tri 2260 5091 2268 5099 se
rect 2268 5091 2318 5158
rect 2008 4373 2020 4407
rect 2054 4373 2066 4407
rect 2008 4335 2066 4373
rect 2008 4301 2020 4335
rect 2054 4301 2066 4335
rect 2008 4295 2066 4301
rect 2135 4466 2191 4467
rect 2134 4407 2192 4465
rect 2134 4373 2146 4407
rect 2180 4373 2192 4407
rect 2134 4335 2192 4373
rect 2134 4301 2146 4335
rect 2180 4301 2192 4335
rect 2134 4295 2192 4301
rect 2260 4407 2318 5091
rect 2386 5270 2444 5276
rect 2386 5236 2398 5270
rect 2432 5236 2444 5270
rect 2386 5198 2444 5236
rect 2386 5164 2398 5198
rect 2432 5164 2444 5198
rect 2386 4505 2444 5164
rect 2387 4503 2443 4504
rect 2512 5270 2696 5276
rect 2512 5236 2524 5270
rect 2558 5236 2650 5270
rect 2684 5236 2696 5270
rect 2512 5198 2696 5236
rect 2512 5164 2524 5198
rect 2558 5164 2650 5198
rect 2684 5164 2696 5198
rect 2512 5158 2696 5164
rect 2512 5091 2562 5158
tri 2562 5133 2587 5158 nw
tri 2621 5133 2646 5158 ne
tri 2562 5091 2570 5099 sw
rect 2260 4373 2272 4407
rect 2306 4373 2318 4407
rect 2260 4335 2318 4373
rect 2260 4301 2272 4335
rect 2306 4301 2318 4335
rect 2260 4295 2318 4301
rect 2387 4466 2443 4467
rect 2386 4407 2444 4465
rect 2386 4373 2398 4407
rect 2432 4373 2444 4407
rect 2386 4335 2444 4373
rect 2386 4301 2398 4335
rect 2432 4301 2444 4335
rect 2386 4295 2444 4301
rect 2512 4407 2570 5091
rect 2512 4373 2524 4407
rect 2558 4373 2570 4407
rect 2512 4335 2570 4373
rect 2512 4301 2524 4335
rect 2558 4301 2570 4335
rect 2512 4295 2570 4301
tri 2638 5091 2646 5099 se
rect 2646 5091 2696 5158
rect 2638 4407 2696 5091
rect 2638 4373 2650 4407
rect 2684 4373 2696 4407
rect 2638 4335 2696 4373
rect 2638 4301 2650 4335
rect 2684 4301 2696 4335
rect 2638 4295 2696 4301
rect 2764 5270 2948 5276
rect 2764 5236 2776 5270
rect 2810 5236 2902 5270
rect 2936 5236 2948 5270
rect 2764 5198 2948 5236
rect 2764 5164 2776 5198
rect 2810 5164 2902 5198
rect 2936 5164 2948 5198
rect 2764 5158 2948 5164
rect 2764 5091 2814 5158
tri 2814 5133 2839 5158 nw
tri 2873 5133 2898 5158 ne
tri 2814 5091 2822 5099 sw
rect 2764 4407 2822 5091
rect 2764 4373 2776 4407
rect 2810 4373 2822 4407
rect 2764 4335 2822 4373
rect 2764 4301 2776 4335
rect 2810 4301 2822 4335
rect 2764 4295 2822 4301
tri 2890 5091 2898 5099 se
rect 2898 5091 2948 5158
rect 2890 4407 2948 5091
rect 2890 4373 2902 4407
rect 2936 4373 2948 4407
rect 2890 4335 2948 4373
rect 2890 4301 2902 4335
rect 2936 4301 2948 4335
rect 2890 4295 2948 4301
rect 3016 5270 3074 5276
rect 3016 5236 3028 5270
rect 3062 5236 3074 5270
rect 3798 5260 3844 5299
tri 3844 5279 3864 5299 nw
tri 4090 5279 4110 5299 ne
rect 4110 5260 4156 5299
tri 4156 5279 4176 5299 nw
tri 4402 5279 4422 5299 ne
rect 4422 5260 4468 5299
tri 4468 5279 4488 5299 nw
tri 4714 5284 4729 5299 ne
rect 4729 5284 4780 5299
tri 4729 5279 4734 5284 ne
rect 4734 5260 4780 5284
tri 4792 5276 4858 5342 ne
tri 4858 5304 4896 5342 sw
tri 4910 5304 4948 5342 ne
rect 4948 5304 5682 5342
rect 4858 5276 4896 5304
tri 4896 5276 4924 5304 sw
tri 4858 5260 4874 5276 ne
rect 4874 5260 5066 5276
rect 3016 5198 3074 5236
rect 3016 5164 3028 5198
rect 3062 5164 3074 5198
rect 3016 4407 3074 5164
rect 3016 4373 3028 4407
rect 3062 4373 3074 4407
rect 3016 4335 3074 4373
rect 3016 4301 3028 4335
rect 3062 4301 3074 4335
rect 3016 4295 3074 4301
rect 3144 4341 3525 5260
tri 4874 5248 4886 5260 ne
rect 4886 5248 5066 5260
tri 4886 5230 4904 5248 ne
rect 4904 5230 5066 5248
tri 5041 5214 5057 5230 ne
rect 5057 5214 5066 5230
tri 5057 5205 5066 5214 ne
rect 5498 5248 5580 5260
rect 5498 5214 5504 5248
rect 5538 5214 5580 5248
rect 5498 5166 5580 5214
rect 5498 5132 5504 5166
rect 5538 5132 5580 5166
rect 5498 5084 5580 5132
rect 5498 5050 5504 5084
rect 5538 5050 5580 5084
rect 5498 5002 5580 5050
rect 5498 4968 5504 5002
rect 5538 4968 5580 5002
rect 5498 4920 5580 4968
rect 5498 4886 5504 4920
rect 5538 4886 5580 4920
rect 5498 4838 5580 4886
rect 5498 4804 5504 4838
rect 5538 4804 5580 4838
rect 5498 4755 5580 4804
rect 5498 4721 5504 4755
rect 5538 4721 5580 4755
rect 5498 4708 5580 4721
tri 5498 4678 5528 4708 ne
tri 3688 4602 3713 4627 sw
tri 3929 4602 3954 4627 se
tri 4000 4602 4025 4627 sw
tri 4241 4602 4266 4627 se
tri 4312 4602 4337 4627 sw
tri 4553 4602 4578 4627 se
tri 4624 4602 4649 4627 sw
tri 4865 4602 4890 4627 se
tri 4936 4602 4961 4627 sw
tri 5217 4602 5242 4627 se
rect 5528 4603 5580 4708
rect 3642 4596 5288 4602
rect 5529 4601 5579 4602
tri 5661 4601 5662 4602 sw
rect 3758 4416 5172 4596
rect 5661 4577 5662 4601
tri 5662 4577 5686 4601 sw
rect 3642 4410 5288 4416
rect 5529 4564 5579 4565
rect 5528 4505 5580 4563
rect 5661 4531 5686 4577
tri 5661 4506 5686 4531 nw
rect 5528 4441 5580 4453
rect 5528 4383 5580 4389
tri 3571 4341 3596 4366 sw
tri 5590 4341 5615 4366 se
rect 3144 4295 3592 4341
rect 5594 4295 5661 4341
tri 1308 4275 1325 4292 sw
rect 1262 4272 1325 4275
tri 1262 4267 1267 4272 ne
rect 1267 4267 1325 4272
tri 1325 4267 1333 4275 sw
tri 1267 4226 1308 4267 ne
rect 1308 4226 5682 4267
tri 1308 4221 1313 4226 ne
rect 1313 4221 5682 4226
rect 59 4187 5534 4193
rect 59 4141 2896 4187
tri 1857 4116 1882 4141 ne
rect 1882 4118 1942 4141
tri 1942 4118 1965 4141 nw
tri 2109 4118 2132 4141 ne
rect 2132 4118 2192 4141
tri 2192 4118 2215 4141 nw
tri 2361 4118 2384 4141 ne
rect 2384 4118 2444 4141
tri 2444 4118 2467 4141 nw
tri 2613 4118 2636 4141 ne
rect 2636 4118 2696 4141
tri 2696 4118 2719 4141 nw
tri 2865 4118 2888 4141 ne
rect 2888 4135 2896 4141
rect 2948 4141 5534 4187
rect 5586 4141 5598 4193
rect 5650 4141 5682 4193
rect 2888 4123 2948 4135
rect 2888 4118 2896 4123
rect 1940 4117 1941 4118
tri 1941 4117 1942 4118 nw
tri 2132 4117 2133 4118 ne
rect 2133 4117 2134 4118
tri 2384 4117 2385 4118 ne
rect 2385 4117 2386 4118
tri 2636 4117 2637 4118 ne
rect 2637 4117 2638 4118
tri 2888 4117 2889 4118 ne
rect 2889 4117 2896 4118
rect 1883 4116 1939 4117
tri 1940 4116 1941 4117 nw
tri 2133 4116 2134 4117 ne
rect 2135 4116 2191 4117
tri 2385 4116 2386 4117 ne
rect 2387 4116 2443 4117
tri 2637 4116 2638 4117 ne
rect 2639 4116 2695 4117
tri 2889 4116 2890 4117 ne
rect 248 3468 300 4108
rect 370 4107 428 4113
rect 370 4073 382 4107
rect 416 4073 428 4107
rect 370 4035 428 4073
rect 370 4001 382 4035
rect 416 4001 428 4035
rect 370 493 428 4001
rect 496 4107 554 4113
rect 496 4073 508 4107
rect 542 4073 554 4107
rect 496 4035 554 4073
rect 496 4001 508 4035
rect 542 4001 554 4035
rect 496 3943 554 4001
rect 497 3941 553 3942
rect 622 4107 680 4113
rect 622 4073 634 4107
rect 668 4073 680 4107
rect 622 4035 680 4073
rect 622 4001 634 4035
rect 668 4001 680 4035
rect 370 441 373 493
rect 425 441 428 493
rect 370 429 428 441
rect 370 377 373 429
rect 425 377 428 429
rect 370 371 428 377
rect 497 3904 553 3905
rect 496 493 554 3903
rect 622 642 680 4001
rect 748 4107 806 4113
rect 748 4073 760 4107
rect 794 4073 806 4107
rect 748 4035 806 4073
rect 748 4001 760 4035
rect 794 4001 806 4035
rect 748 3943 806 4001
rect 874 4107 932 4113
rect 874 4073 886 4107
rect 920 4073 932 4107
rect 874 4035 932 4073
rect 874 4001 886 4035
rect 920 4001 932 4035
rect 874 3995 932 4001
rect 1000 4107 1058 4113
rect 1000 4073 1012 4107
rect 1046 4073 1058 4107
rect 1000 4035 1058 4073
rect 1000 4001 1012 4035
rect 1046 4001 1058 4035
rect 1000 3995 1058 4001
rect 1126 4107 1184 4113
rect 1126 4073 1138 4107
rect 1172 4073 1184 4107
rect 1126 4035 1184 4073
rect 1126 4001 1138 4035
rect 1172 4001 1184 4035
rect 749 3941 805 3942
rect 622 634 672 642
tri 672 634 680 642 nw
rect 749 3904 805 3905
rect 622 590 664 634
tri 664 626 672 634 nw
rect 623 588 663 589
rect 496 441 499 493
rect 551 441 554 493
rect 496 429 554 441
rect 496 377 499 429
rect 551 377 554 429
rect 623 551 663 552
rect 622 500 664 550
tri 664 500 687 523 sw
tri 725 500 748 523 se
rect 748 500 806 3903
rect 1126 642 1184 4001
rect 1252 4107 1310 4113
rect 1252 4073 1264 4107
rect 1298 4073 1310 4107
rect 1252 4035 1310 4073
rect 1252 4001 1264 4035
rect 1298 4001 1310 4035
rect 1252 3943 1310 4001
rect 1253 3941 1309 3942
rect 1378 4107 1436 4113
rect 1378 4073 1390 4107
rect 1424 4073 1436 4107
rect 1378 4035 1436 4073
rect 1378 4001 1390 4035
rect 1424 4001 1436 4035
rect 1126 634 1176 642
tri 1176 634 1184 642 nw
rect 1253 3904 1309 3905
rect 1126 590 1168 634
tri 1168 626 1176 634 nw
rect 1127 588 1167 589
rect 622 498 687 500
tri 687 498 689 500 sw
tri 723 498 725 500 se
rect 725 498 806 500
rect 1127 551 1167 552
rect 1126 500 1168 550
tri 1168 500 1191 523 sw
tri 1229 500 1252 523 se
rect 1252 500 1310 3903
rect 1378 642 1436 4001
rect 1504 4107 1562 4113
rect 1504 4073 1516 4107
rect 1550 4073 1562 4107
rect 1504 4035 1562 4073
rect 1504 4001 1516 4035
rect 1550 4001 1562 4035
rect 1504 3943 1562 4001
rect 1505 3941 1561 3942
rect 1630 4107 1688 4113
rect 1630 4073 1642 4107
rect 1676 4073 1688 4107
rect 1630 4035 1688 4073
rect 1630 4001 1642 4035
rect 1676 4001 1688 4035
rect 1378 634 1428 642
tri 1428 634 1436 642 nw
rect 1505 3904 1561 3905
rect 1378 590 1420 634
tri 1420 626 1428 634 nw
rect 1379 588 1419 589
rect 1126 498 1191 500
tri 1191 498 1193 500 sw
tri 1227 498 1229 500 se
rect 1229 498 1310 500
rect 622 492 806 498
rect 622 458 634 492
rect 668 458 760 492
rect 794 458 806 492
rect 622 420 806 458
rect 622 386 634 420
rect 668 386 760 420
rect 794 386 806 420
rect 622 380 806 386
rect 874 492 1058 498
rect 874 458 886 492
rect 920 458 1012 492
rect 1046 458 1058 492
rect 874 420 1058 458
rect 874 386 886 420
rect 920 386 1012 420
rect 1046 386 1058 420
rect 874 380 1058 386
rect 1126 492 1310 498
rect 1126 458 1138 492
rect 1172 458 1264 492
rect 1298 458 1310 492
rect 1126 420 1310 458
rect 1126 386 1138 420
rect 1172 386 1264 420
rect 1298 386 1310 420
rect 1126 380 1310 386
rect 1379 551 1419 552
rect 1378 500 1420 550
tri 1420 500 1443 523 sw
tri 1481 500 1504 523 se
rect 1504 500 1562 3903
rect 1630 642 1688 4001
rect 1756 4107 1814 4113
rect 1756 4073 1768 4107
rect 1802 4073 1814 4107
rect 1756 4035 1814 4073
rect 1756 4001 1768 4035
rect 1802 4001 1814 4035
rect 1756 3943 1814 4001
rect 1757 3941 1813 3942
rect 1882 4080 1940 4116
rect 1883 4079 1939 4080
rect 1882 4072 1940 4078
rect 1882 4038 1894 4072
rect 1928 4038 1940 4072
rect 1882 4000 1940 4038
rect 1882 3966 1894 4000
rect 1928 3966 1940 4000
rect 1882 3943 1940 3966
rect 1883 3941 1939 3942
rect 2008 4107 2066 4113
rect 2008 4073 2020 4107
rect 2054 4073 2066 4107
rect 2260 4107 2318 4113
rect 2008 4035 2066 4073
rect 2008 4001 2020 4035
rect 2054 4001 2066 4035
rect 2008 3943 2066 4001
rect 2009 3941 2065 3942
rect 2135 4079 2191 4080
rect 2134 4072 2192 4078
rect 2134 4038 2146 4072
rect 2180 4038 2192 4072
rect 2134 4000 2192 4038
rect 2134 3966 2146 4000
rect 2180 3966 2192 4000
rect 1630 634 1680 642
tri 1680 634 1688 642 nw
rect 1757 3904 1813 3905
rect 1630 590 1672 634
tri 1672 626 1680 634 nw
rect 1631 588 1671 589
rect 1378 498 1443 500
tri 1443 498 1445 500 sw
tri 1479 498 1481 500 se
rect 1481 498 1562 500
rect 1378 492 1562 498
rect 1378 458 1390 492
rect 1424 458 1516 492
rect 1550 458 1562 492
rect 1378 420 1562 458
rect 1378 386 1390 420
rect 1424 386 1516 420
rect 1550 386 1562 420
rect 1378 380 1562 386
rect 1631 551 1671 552
rect 1630 500 1672 550
tri 1672 500 1695 523 sw
tri 1733 500 1756 523 se
rect 1756 500 1814 3903
rect 1630 498 1695 500
tri 1695 498 1697 500 sw
tri 1731 498 1733 500 se
rect 1733 498 1814 500
rect 1630 492 1814 498
rect 1630 458 1642 492
rect 1676 458 1768 492
rect 1802 458 1814 492
rect 1630 420 1814 458
rect 1630 386 1642 420
rect 1676 386 1768 420
rect 1802 386 1814 420
rect 1630 380 1814 386
rect 1883 3904 1939 3905
rect 1882 492 1940 3903
rect 1882 458 1894 492
rect 1928 458 1940 492
rect 2009 3904 2065 3905
rect 2008 645 2066 3903
rect 2008 642 2063 645
tri 2063 642 2066 645 nw
rect 2134 645 2192 3966
rect 2260 4073 2272 4107
rect 2306 4073 2318 4107
rect 2512 4107 2570 4113
rect 2260 4035 2318 4073
rect 2260 4001 2272 4035
rect 2306 4001 2318 4035
rect 2260 3943 2318 4001
rect 2261 3941 2317 3942
rect 2387 4079 2443 4080
rect 2386 4072 2444 4078
rect 2386 4038 2398 4072
rect 2432 4038 2444 4072
rect 2386 4000 2444 4038
rect 2386 3966 2398 4000
rect 2432 3966 2444 4000
tri 2134 642 2137 645 ne
rect 2137 642 2192 645
rect 2008 600 2058 642
tri 2058 637 2063 642 nw
tri 2137 637 2142 642 ne
tri 2058 600 2061 603 sw
tri 2139 600 2142 603 se
rect 2142 600 2192 642
rect 2008 588 2061 600
tri 2061 588 2073 600 sw
tri 2127 588 2139 600 se
rect 2139 588 2192 600
rect 2008 578 2073 588
tri 2073 578 2083 588 sw
tri 2117 578 2127 588 se
rect 2127 578 2192 588
rect 2008 572 2192 578
rect 2008 538 2020 572
rect 2054 538 2146 572
rect 2180 538 2192 572
rect 2008 500 2192 538
rect 2008 466 2020 500
rect 2054 466 2146 500
rect 2180 466 2192 500
rect 2008 460 2192 466
rect 2261 3904 2317 3905
rect 2260 645 2318 3903
rect 2260 642 2315 645
tri 2315 642 2318 645 nw
rect 2386 645 2444 3966
rect 2512 4073 2524 4107
rect 2558 4073 2570 4107
rect 2764 4107 2822 4113
rect 2512 4035 2570 4073
rect 2512 4001 2524 4035
rect 2558 4001 2570 4035
rect 2512 3943 2570 4001
rect 2513 3941 2569 3942
rect 2639 4079 2695 4080
rect 2638 4072 2696 4078
rect 2638 4038 2650 4072
rect 2684 4038 2696 4072
rect 2638 4000 2696 4038
rect 2638 3966 2650 4000
rect 2684 3966 2696 4000
rect 2638 3943 2696 3966
rect 2639 3941 2695 3942
rect 2764 4073 2776 4107
rect 2810 4073 2822 4107
rect 2764 4035 2822 4073
rect 2890 4071 2896 4117
tri 2948 4116 2973 4141 nw
rect 2890 4065 2948 4071
rect 2891 4063 2947 4064
rect 3014 4107 3078 4113
rect 3014 4073 3028 4107
rect 3062 4073 3078 4107
rect 2764 4001 2776 4035
rect 2810 4001 2822 4035
rect 3014 4035 3078 4073
rect 3144 4061 5682 4113
tri 3260 4036 3285 4061 nw
rect 2764 3943 2822 4001
rect 2765 3941 2821 3942
rect 2891 4026 2947 4027
rect 2890 4019 2948 4025
rect 2890 3985 2902 4019
rect 2936 3985 2948 4019
rect 2890 3947 2948 3985
rect 2890 3913 2902 3947
rect 2936 3913 2948 3947
tri 2386 642 2389 645 ne
rect 2389 642 2444 645
rect 2260 600 2310 642
tri 2310 637 2315 642 nw
tri 2389 637 2394 642 ne
tri 2310 600 2313 603 sw
tri 2391 600 2394 603 se
rect 2394 600 2444 642
rect 2260 588 2313 600
tri 2313 588 2325 600 sw
tri 2379 588 2391 600 se
rect 2391 588 2444 600
rect 2260 578 2325 588
tri 2325 578 2335 588 sw
tri 2369 578 2379 588 se
rect 2379 578 2444 588
rect 2260 572 2444 578
rect 2260 538 2272 572
rect 2306 538 2398 572
rect 2432 538 2444 572
rect 2260 500 2444 538
rect 2260 466 2272 500
rect 2306 466 2398 500
rect 2432 466 2444 500
rect 2260 460 2444 466
rect 2513 3904 2569 3905
rect 2512 492 2570 3903
rect 1882 448 1940 458
rect 2512 458 2524 492
rect 2558 458 2570 492
tri 1940 448 1949 457 sw
tri 2503 448 2512 457 se
rect 2512 448 2570 458
rect 1882 432 1949 448
tri 1949 432 1965 448 sw
tri 2487 432 2503 448 se
rect 2503 432 2570 448
rect 1882 420 2570 432
rect 1882 386 1894 420
rect 1928 386 2524 420
rect 2558 386 2570 420
rect 1882 380 2570 386
rect 2639 3904 2695 3905
rect 2638 565 2696 3903
rect 2638 558 2689 565
tri 2689 558 2696 565 nw
rect 2765 3904 2821 3905
rect 2764 565 2822 3903
rect 2890 3890 2948 3913
rect 2891 3888 2947 3889
rect 3014 4001 3028 4035
rect 3062 4001 3078 4035
tri 2764 558 2771 565 ne
rect 2771 558 2822 565
rect 2638 498 2688 558
tri 2688 557 2689 558 nw
tri 2771 557 2772 558 ne
tri 2688 498 2713 523 sw
tri 2747 498 2772 523 se
rect 2772 498 2822 558
rect 2638 492 2822 498
rect 2638 458 2650 492
rect 2684 458 2776 492
rect 2810 458 2822 492
rect 2638 420 2822 458
rect 2638 386 2650 420
rect 2684 386 2776 420
rect 2810 386 2822 420
rect 2638 380 2822 386
rect 2891 3851 2947 3852
rect 2890 492 2948 3850
rect 2890 458 2902 492
rect 2936 458 2948 492
rect 2890 420 2948 458
rect 2890 386 2902 420
rect 2936 386 2948 420
rect 2890 380 2948 386
rect 3014 496 3078 4001
tri 3260 3719 3285 3744 sw
rect 3260 3589 3621 3719
tri 3260 3564 3285 3589 nw
tri 3260 3150 3285 3175 sw
rect 3260 3098 3573 3150
tri 3260 3073 3285 3098 nw
tri 3260 2880 3285 2905 sw
rect 3260 2828 3573 2880
tri 3260 2803 3285 2828 nw
tri 3260 1619 3285 1644 sw
rect 3260 1567 3604 1619
tri 3260 1542 3285 1567 nw
tri 3260 1110 3285 1135 sw
rect 3260 1064 3592 1110
tri 3260 1039 3285 1064 nw
rect 3014 444 3020 496
rect 3072 444 3078 496
rect 3014 432 3078 444
rect 3014 380 3020 432
rect 3072 380 3078 432
rect 3336 862 3382 874
rect 3336 828 3342 862
rect 3376 828 3382 862
rect 3336 786 3382 828
rect 3336 752 3342 786
rect 3376 752 3382 786
rect 3336 710 3382 752
rect 3336 676 3342 710
rect 3376 676 3382 710
rect 3336 634 3382 676
rect 3336 600 3342 634
rect 3376 600 3382 634
rect 3336 558 3382 600
rect 3336 524 3342 558
rect 3376 524 3382 558
rect 3336 482 3382 524
rect 3336 448 3342 482
rect 3376 448 3382 482
rect 3336 406 3382 448
rect 496 371 554 377
rect 3336 372 3342 406
rect 3376 372 3382 406
rect 3336 330 3382 372
rect 248 182 300 306
rect 729 210 735 262
rect 787 210 799 262
rect 851 210 863 262
rect 915 210 921 262
rect 1005 210 1011 262
rect 1063 210 1075 262
rect 1127 210 1139 262
rect 1191 210 1197 262
tri 1306 220 1338 252 se
rect 1338 220 1344 252
tri 1296 210 1306 220 se
rect 1306 210 1344 220
tri 1293 207 1296 210 se
rect 1296 207 1344 210
tri 300 182 325 207 sw
tri 1268 182 1293 207 se
rect 1293 182 1344 207
rect 248 175 326 182
tri 248 144 279 175 ne
rect 279 144 326 175
tri 279 136 287 144 ne
rect 287 136 326 144
rect 1338 136 1344 182
rect 1460 241 2049 252
tri 2049 241 2060 252 sw
rect 1460 220 2060 241
tri 2060 220 2081 241 sw
tri 3123 220 3144 241 se
rect 3144 220 3193 306
rect 1460 196 2081 220
tri 2081 196 2105 220 sw
tri 3099 196 3123 220 se
rect 3123 196 3193 220
rect 1460 182 3193 196
rect 1460 136 1466 182
rect 3120 171 3193 182
rect 3120 144 3166 171
tri 3166 144 3193 171 nw
rect 3336 296 3342 330
rect 3376 296 3382 330
rect 3336 254 3382 296
rect 3336 220 3342 254
rect 3376 220 3382 254
rect 3336 178 3382 220
rect 3336 144 3342 178
rect 3376 144 3382 178
rect 3120 136 3158 144
tri 3158 136 3166 144 nw
tri 3328 136 3336 144 se
rect 3336 136 3382 144
tri 3300 108 3328 136 se
rect 3328 108 3382 136
rect 326 102 3382 108
rect 326 70 3342 102
rect 326 38 742 70
rect 409 36 742 38
rect 776 68 3342 70
rect 3376 84 3382 102
tri 3382 84 3442 144 sw
rect 3376 68 3670 84
rect 776 38 3670 68
rect 776 36 3650 38
rect 409 18 3650 36
tri 3650 18 3670 38 nw
rect 409 6 3645 18
tri 3645 13 3650 18 nw
rect 409 -16 3605 6
rect 229 -18 475 -16
tri 475 -18 477 -16 nw
tri 711 -18 713 -16 ne
rect 713 -18 795 -16
rect 229 -32 461 -18
tri 461 -32 475 -18 nw
tri 713 -32 727 -18 ne
rect 727 -32 742 -18
rect 229 -44 449 -32
tri 449 -44 461 -32 nw
tri 727 -41 736 -32 ne
rect 229 -52 441 -44
tri 441 -52 449 -44 nw
rect 736 -52 742 -32
rect 776 -28 795 -18
tri 795 -28 807 -16 nw
tri 1005 -28 1017 -16 ne
rect 1017 -28 1089 -16
tri 1089 -28 1101 -16 nw
tri 1357 -28 1369 -16 ne
rect 1369 -28 1441 -16
tri 1441 -28 1453 -16 nw
tri 1709 -28 1721 -16 ne
rect 1721 -28 1793 -16
tri 1793 -28 1805 -16 nw
tri 2061 -28 2073 -16 ne
rect 2073 -28 2145 -16
tri 2145 -28 2157 -16 nw
tri 2883 -28 2895 -16 ne
rect 2895 -28 2967 -16
tri 2967 -28 2979 -16 nw
tri 3574 -28 3586 -16 ne
rect 3586 -28 3605 -16
rect 3639 -28 3645 6
rect 776 -32 791 -28
tri 791 -32 795 -28 nw
tri 1017 -32 1021 -28 ne
rect 1021 -32 1085 -28
tri 1085 -32 1089 -28 nw
tri 1369 -32 1373 -28 ne
rect 1373 -32 1437 -28
tri 1437 -32 1441 -28 nw
tri 1721 -32 1725 -28 ne
rect 1725 -32 1789 -28
tri 1789 -32 1793 -28 nw
tri 2073 -32 2077 -28 ne
rect 2077 -32 2141 -28
tri 2141 -32 2145 -28 nw
tri 2895 -32 2899 -28 ne
rect 2899 -32 2963 -28
tri 2963 -32 2967 -28 nw
tri 3586 -32 3590 -28 ne
rect 3590 -32 3645 -28
rect 776 -52 782 -32
tri 782 -41 791 -32 nw
tri 1021 -41 1030 -32 ne
rect 1030 -44 1076 -32
tri 1076 -41 1085 -32 nw
tri 1373 -41 1382 -32 ne
rect 1382 -44 1428 -32
tri 1428 -41 1437 -32 nw
tri 1725 -41 1734 -32 ne
rect 1734 -44 1780 -32
tri 1780 -41 1789 -32 nw
tri 2077 -41 2086 -32 ne
rect 2086 -44 2132 -32
tri 2132 -41 2141 -32 nw
tri 2899 -41 2908 -32 ne
rect 2908 -44 2954 -32
tri 2954 -41 2963 -32 nw
tri 3590 -41 3599 -32 ne
rect 229 -56 437 -52
tri 437 -56 441 -52 nw
rect 229 -320 409 -56
tri 409 -84 437 -56 nw
rect 736 -107 782 -52
rect 499 -143 551 -137
rect 499 -207 551 -195
rect 736 -141 742 -107
rect 776 -141 782 -107
rect 736 -196 782 -141
rect 2452 -56 2498 -44
rect 2452 -90 2458 -56
rect 2492 -90 2498 -56
rect 2452 -128 2498 -90
rect 2452 -162 2458 -128
rect 2492 -162 2498 -128
rect 2908 -78 2914 -44
rect 2948 -78 2954 -44
rect 2908 -116 2954 -78
rect 2908 -150 2914 -116
rect 2948 -150 2954 -116
rect 3364 -56 3410 -44
rect 3364 -90 3370 -56
rect 3404 -90 3410 -56
rect 2908 -162 2954 -150
rect 3054 -124 3106 -118
tri 2337 -174 2342 -169 se
tri 2317 -194 2337 -174 se
rect 2337 -194 2342 -174
rect 736 -230 742 -196
rect 776 -230 782 -196
rect 736 -242 782 -230
rect 2241 -246 2266 -194
rect 2318 -246 2330 -194
rect 2382 -246 2388 -194
rect 2452 -200 2498 -162
tri 3029 -200 3054 -175 se
rect 3364 -128 3410 -90
rect 3364 -162 3370 -128
rect 3404 -162 3410 -128
rect 3054 -188 3106 -176
rect 2452 -234 2458 -200
rect 2492 -234 2498 -200
tri 551 -257 553 -255 sw
rect 551 -259 553 -257
rect 499 -271 553 -259
tri 409 -320 413 -316 sw
rect 229 -329 413 -320
tri 413 -329 422 -320 sw
rect 551 -280 553 -271
tri 553 -280 576 -257 sw
tri 831 -280 854 -257 se
rect 854 -280 900 -246
tri 900 -280 923 -257 sw
tri 1183 -280 1206 -257 se
rect 1206 -280 1252 -246
tri 1252 -280 1275 -257 sw
tri 1535 -280 1558 -257 se
rect 1558 -274 1604 -246
tri 1604 -274 1621 -257 sw
tri 1893 -274 1910 -257 se
rect 1910 -274 1956 -246
rect 2241 -247 2312 -246
tri 2312 -247 2313 -246 nw
rect 2241 -248 2311 -247
tri 2311 -248 2312 -247 nw
tri 2240 -249 2241 -248 se
rect 2241 -249 2310 -248
tri 2310 -249 2311 -248 nw
tri 2215 -274 2240 -249 se
rect 2240 -274 2285 -249
tri 2285 -274 2310 -249 nw
tri 2427 -274 2452 -249 se
rect 2452 -274 2498 -234
rect 2535 -206 3054 -200
rect 2535 -240 2547 -206
rect 2581 -240 2619 -206
rect 2653 -240 2691 -206
rect 2725 -240 2763 -206
rect 2797 -240 2835 -206
rect 2869 -240 3054 -206
tri 3106 -200 3131 -175 sw
tri 3339 -200 3364 -175 se
rect 3364 -200 3410 -162
rect 3106 -234 3370 -200
rect 3404 -234 3410 -200
rect 3106 -240 3410 -234
rect 2535 -246 3410 -240
rect 3599 -67 3645 -32
rect 3599 -101 3605 -67
rect 3639 -101 3645 -67
rect 3599 -140 3645 -101
rect 3599 -174 3605 -140
rect 3639 -174 3645 -140
rect 3599 -213 3645 -174
rect 3599 -247 3605 -213
rect 3639 -247 3645 -213
tri 2498 -274 2523 -249 sw
rect 1558 -280 1621 -274
tri 1621 -280 1627 -274 sw
tri 1887 -280 1893 -274 se
rect 1893 -280 1956 -274
rect 551 -282 576 -280
tri 576 -282 578 -280 sw
tri 829 -282 831 -280 se
rect 831 -282 923 -280
tri 923 -282 925 -280 sw
tri 1181 -282 1183 -280 se
rect 1183 -282 1275 -280
tri 1275 -282 1277 -280 sw
tri 1533 -282 1535 -280 se
rect 1535 -282 1627 -280
tri 1627 -282 1629 -280 sw
tri 1885 -282 1887 -280 se
rect 1887 -282 1956 -280
rect 551 -285 1956 -282
rect 551 -314 1927 -285
tri 1927 -314 1956 -285 nw
rect 1985 -280 2279 -274
tri 2279 -280 2285 -274 nw
rect 2325 -280 2696 -274
rect 1985 -314 1997 -280
rect 2031 -314 2069 -280
rect 2103 -314 2245 -280
tri 2245 -314 2279 -280 nw
rect 2325 -314 2337 -280
rect 2371 -314 2409 -280
rect 2443 -314 2696 -280
rect 551 -320 1921 -314
tri 1921 -320 1927 -314 nw
rect 1985 -320 2239 -314
tri 2239 -320 2245 -314 nw
rect 2325 -320 2696 -314
rect 551 -323 1915 -320
rect 499 -326 1915 -323
tri 1915 -326 1921 -320 nw
tri 2684 -326 2690 -320 ne
rect 2690 -326 2696 -320
rect 2748 -326 2760 -274
rect 2812 -280 3260 -274
rect 2812 -314 2998 -280
rect 3032 -314 3070 -280
rect 3104 -314 3142 -280
rect 3176 -314 3214 -280
rect 3248 -314 3260 -280
rect 2812 -320 3260 -314
rect 3599 -286 3645 -247
rect 3599 -320 3605 -286
rect 3639 -320 3645 -286
rect 2812 -326 2818 -320
tri 2818 -326 2824 -320 nw
rect 499 -329 1912 -326
tri 1912 -329 1915 -326 nw
rect 229 -359 422 -329
tri 422 -359 452 -329 sw
tri 829 -334 834 -329 ne
rect 834 -334 920 -329
tri 920 -334 925 -329 nw
tri 1181 -334 1186 -329 ne
rect 1186 -334 1272 -329
tri 1272 -334 1277 -329 nw
tri 1533 -334 1538 -329 ne
rect 1538 -334 1624 -329
tri 1624 -334 1629 -329 nw
tri 834 -354 854 -334 ne
rect 229 -365 452 -359
tri 452 -365 458 -359 sw
rect 229 -369 458 -365
tri 458 -369 462 -365 sw
rect 229 -381 782 -369
rect 854 -378 900 -334
tri 900 -354 920 -334 nw
tri 1186 -354 1206 -334 ne
rect 1206 -378 1252 -334
tri 1252 -354 1272 -334 nw
tri 1538 -354 1558 -334 ne
rect 1558 -378 1604 -334
tri 1604 -354 1624 -334 nw
tri 3579 -354 3599 -334 se
rect 3599 -354 3645 -320
tri 3574 -359 3579 -354 se
rect 3579 -359 3645 -354
rect 1675 -365 3605 -359
rect 1675 -371 1756 -365
rect 229 -415 742 -381
rect 776 -415 782 -381
rect 229 -462 782 -415
rect 229 -496 742 -462
rect 776 -496 782 -462
rect 229 -543 782 -496
rect 229 -577 742 -543
rect 776 -577 782 -543
rect 229 -580 782 -577
rect 1675 -405 1681 -371
rect 1715 -399 1756 -371
rect 1790 -399 1830 -365
rect 1864 -399 1904 -365
rect 1938 -399 1978 -365
rect 2012 -399 2052 -365
rect 2086 -399 2126 -365
rect 2160 -399 2200 -365
rect 2234 -399 2274 -365
rect 2308 -399 2348 -365
rect 2382 -399 2422 -365
rect 2456 -399 2496 -365
rect 2530 -399 2570 -365
rect 2604 -399 2644 -365
rect 2678 -399 2718 -365
rect 2752 -399 2792 -365
rect 2826 -399 2866 -365
rect 2900 -399 2940 -365
rect 2974 -399 3014 -365
rect 3048 -399 3088 -365
rect 3122 -399 3162 -365
rect 3196 -399 3236 -365
rect 3270 -399 3310 -365
rect 3344 -399 3384 -365
rect 3418 -399 3458 -365
rect 3492 -399 3533 -365
rect 3567 -393 3605 -365
rect 3639 -393 3645 -359
rect 3567 -399 3645 -393
rect 1715 -405 3645 -399
rect 1675 -464 1724 -405
tri 1724 -430 1749 -405 nw
rect 1675 -498 1681 -464
rect 1715 -498 1724 -464
rect 1675 -557 1724 -498
tri 229 -591 240 -580 ne
rect 240 -591 782 -580
tri 1028 -591 1030 -589 se
rect 1030 -591 1076 -580
tri 1076 -591 1078 -589 sw
tri 1380 -591 1382 -589 se
rect 1382 -591 1428 -580
tri 1428 -591 1430 -589 sw
rect 1675 -591 1681 -557
rect 1715 -591 1724 -557
tri 240 -594 243 -591 ne
rect 243 -594 782 -591
tri 1025 -594 1028 -591 se
rect 1028 -594 1078 -591
tri 1078 -594 1081 -591 sw
tri 1377 -594 1380 -591 se
rect 1380 -594 1430 -591
tri 1430 -594 1433 -591 sw
tri 243 -603 252 -594 ne
rect 252 -603 782 -594
tri 1021 -598 1025 -594 se
rect 1025 -598 1081 -594
tri 252 -623 272 -603 ne
rect 272 -623 782 -603
tri 782 -623 807 -598 sw
tri 996 -623 1021 -598 se
rect 1021 -623 1081 -598
tri 1081 -623 1110 -594 sw
tri 1348 -623 1377 -594 se
rect 1377 -598 1433 -594
tri 1433 -598 1437 -594 sw
rect 1377 -603 1437 -598
tri 1437 -603 1442 -598 sw
tri 1670 -603 1675 -598 se
rect 1675 -603 1724 -591
rect 1976 -536 3503 -530
rect 2028 -588 2040 -536
rect 2092 -588 2104 -536
rect 2156 -560 2168 -536
rect 2220 -554 3139 -536
rect 3191 -554 3203 -536
rect 3255 -554 3503 -536
rect 2220 -588 2221 -554
rect 2255 -588 2294 -554
rect 2328 -588 2367 -554
rect 2401 -588 2440 -554
rect 2474 -588 2513 -554
rect 2547 -588 2586 -554
rect 2620 -588 2659 -554
rect 2693 -588 2732 -554
rect 2766 -588 2805 -554
rect 2839 -588 2878 -554
rect 2912 -588 2951 -554
rect 2985 -588 3024 -554
rect 3058 -588 3097 -554
rect 3131 -588 3139 -554
rect 3277 -588 3317 -554
rect 3351 -588 3391 -554
rect 3425 -560 3503 -554
rect 3425 -588 3463 -560
rect 1976 -594 2149 -588
rect 2183 -594 3463 -588
rect 3497 -594 3503 -560
rect 1377 -623 1442 -603
tri 1442 -623 1462 -603 sw
tri 1650 -623 1670 -603 se
rect 1670 -623 1724 -603
tri 2118 -619 2143 -594 ne
tri 272 -657 306 -623 ne
rect 306 -657 742 -623
rect 776 -657 1724 -623
tri 306 -679 328 -657 ne
rect 328 -679 1724 -657
tri 328 -680 329 -679 ne
rect 329 -680 1724 -679
tri 329 -719 368 -680 ne
rect 368 -719 1724 -680
tri 368 -731 380 -719 ne
rect 380 -731 1724 -719
rect 2143 -645 2189 -594
tri 2189 -619 2214 -594 nw
tri 3432 -619 3457 -594 ne
rect 2143 -679 2149 -645
rect 2183 -679 2189 -645
rect 2273 -639 2403 -633
rect 2273 -673 2285 -639
rect 2319 -673 2357 -639
rect 2391 -673 2403 -639
rect 2273 -679 2403 -673
rect 2443 -679 2451 -627
rect 2503 -679 2515 -627
rect 2567 -679 2573 -627
rect 2601 -679 2607 -627
rect 2659 -679 2671 -627
rect 2723 -639 3093 -627
rect 2723 -673 2975 -639
rect 3009 -673 3047 -639
rect 3081 -673 3093 -639
rect 2723 -679 3093 -673
rect 3457 -646 3503 -594
rect 2143 -731 2189 -679
tri 2333 -680 2334 -679 ne
rect 2334 -680 2403 -679
tri 2403 -680 2404 -679 sw
rect 3457 -680 3463 -646
rect 3497 -680 3503 -646
tri 2334 -707 2361 -680 ne
rect 2361 -707 2404 -680
tri 2404 -707 2431 -680 sw
rect 2143 -765 2149 -731
rect 2183 -765 2189 -731
rect 2143 -817 2189 -765
rect 2143 -851 2149 -817
rect 2183 -851 2189 -817
rect 2260 -713 2312 -707
tri 2361 -719 2373 -707 ne
rect 2373 -719 2696 -707
tri 2373 -749 2403 -719 ne
rect 2403 -749 2696 -719
tri 2403 -753 2407 -749 ne
rect 2407 -753 2696 -749
tri 2667 -759 2673 -753 ne
rect 2673 -759 2696 -753
rect 2748 -759 2760 -707
rect 2812 -759 2818 -707
rect 3054 -713 3170 -707
rect 2260 -777 2312 -765
tri 2673 -766 2680 -759 ne
rect 2680 -766 2756 -759
tri 2756 -766 2763 -759 nw
rect 3106 -719 3170 -713
rect 3106 -753 3130 -719
rect 3164 -753 3170 -719
rect 3106 -765 3170 -753
tri 2680 -778 2692 -766 ne
rect 2692 -791 2738 -766
tri 2738 -784 2756 -766 nw
rect 3054 -777 3170 -765
rect 2260 -837 2312 -829
rect 2476 -818 2522 -806
rect 2143 -903 2189 -851
rect 2143 -937 2149 -903
rect 2183 -937 2189 -903
tri 2118 -971 2143 -946 se
rect 2143 -971 2189 -937
rect 2476 -852 2482 -818
rect 2516 -852 2522 -818
rect 2692 -825 2698 -791
rect 2732 -825 2738 -791
rect 2692 -837 2738 -825
rect 2837 -814 3017 -806
tri 2522 -852 2534 -840 sw
tri 2825 -852 2837 -840 se
rect 3106 -791 3170 -777
rect 3457 -732 3503 -680
rect 3457 -766 3463 -732
rect 3497 -766 3503 -732
rect 3457 -778 3503 -766
rect 3106 -825 3130 -791
rect 3164 -825 3170 -791
rect 3106 -829 3170 -825
rect 3054 -837 3170 -829
rect 3340 -814 3604 -806
rect 3340 -818 3424 -814
tri 3017 -852 3029 -840 sw
tri 3328 -852 3340 -840 se
rect 3340 -852 3346 -818
rect 3380 -852 3424 -818
rect 2476 -865 2534 -852
tri 2534 -865 2547 -852 sw
tri 2812 -865 2825 -852 se
rect 2825 -865 2837 -852
rect 2476 -890 2837 -865
rect 3017 -865 3029 -852
tri 3029 -865 3042 -852 sw
tri 3315 -865 3328 -852 se
rect 3328 -865 3424 -852
rect 3017 -890 3424 -865
rect 2476 -924 2482 -890
rect 2516 -924 2837 -890
rect 3017 -924 3346 -890
rect 3380 -924 3424 -890
rect 2476 -930 2837 -924
rect 3017 -930 3424 -924
rect 2476 -943 3604 -930
tri 2189 -971 2214 -946 sw
rect 1976 -977 3457 -971
rect 2028 -1029 2040 -977
rect 2092 -1029 2104 -977
rect 2156 -989 2168 -977
rect 2220 -995 3139 -977
rect 3191 -995 3203 -977
rect 3255 -995 3457 -977
rect 2156 -1029 2168 -1023
rect 2220 -1029 2221 -995
rect 2255 -1029 2294 -995
rect 2328 -1029 2367 -995
rect 2401 -1029 2440 -995
rect 2474 -1029 2513 -995
rect 2547 -1029 2586 -995
rect 2620 -1029 2659 -995
rect 2693 -1029 2732 -995
rect 2766 -1029 2805 -995
rect 2839 -1029 2878 -995
rect 2912 -1029 2951 -995
rect 2985 -1029 3024 -995
rect 3058 -1029 3097 -995
rect 3131 -1029 3139 -995
rect 3277 -1029 3317 -995
rect 3351 -1029 3391 -995
rect 3425 -1029 3457 -995
rect 1976 -1035 3457 -1029
<< rmetal1 >>
rect 496 27386 538 27387
rect 496 27385 497 27386
rect 537 27385 538 27386
rect 496 27348 497 27349
rect 537 27348 538 27349
rect 496 27347 538 27348
rect 622 23959 680 23960
rect 622 23958 623 23959
rect 679 23958 680 23959
rect 1000 27386 1048 27387
rect 1000 27385 1001 27386
rect 1047 27385 1048 27386
rect 874 23959 932 23960
rect 874 23958 875 23959
rect 931 23958 932 23959
rect 1000 27348 1001 27349
rect 1047 27348 1048 27349
rect 1000 27347 1048 27348
rect 496 23491 554 23492
rect 496 23490 497 23491
rect 553 23490 554 23491
rect 622 23921 623 23922
rect 679 23921 680 23922
rect 622 23920 680 23921
rect 874 23921 875 23922
rect 931 23921 932 23922
rect 874 23920 932 23921
rect 496 23453 497 23454
rect 553 23453 554 23454
rect 496 23452 554 23453
rect 622 20064 680 20065
rect 622 20063 623 20064
rect 679 20063 680 20064
rect 1000 23491 1058 23492
rect 1000 23490 1001 23491
rect 1057 23490 1058 23491
rect 874 20064 932 20065
rect 874 20063 875 20064
rect 931 20063 932 20064
rect 1000 23453 1001 23454
rect 1057 23453 1058 23454
rect 1000 23452 1058 23453
rect 622 20026 623 20027
rect 679 20026 680 20027
rect 622 20025 680 20026
rect 874 20026 875 20027
rect 931 20026 932 20027
rect 874 20025 932 20026
rect 748 19596 806 19597
rect 748 19595 749 19596
rect 805 19595 806 19596
rect 622 16169 680 16170
rect 622 16168 623 16169
rect 679 16168 680 16169
rect 748 19558 749 19559
rect 805 19558 806 19559
rect 748 19557 806 19558
rect 622 16131 623 16132
rect 679 16131 680 16132
rect 622 16130 680 16131
rect 1000 19596 1058 19597
rect 1000 19595 1001 19596
rect 1057 19595 1058 19596
rect 874 16169 932 16170
rect 874 16168 875 16169
rect 931 16168 932 16169
rect 1000 19558 1001 19559
rect 1057 19558 1058 19559
rect 1000 19557 1058 19558
rect 748 15701 806 15702
rect 748 15700 749 15701
rect 805 15700 806 15701
rect 874 16131 875 16132
rect 931 16131 932 16132
rect 874 16130 932 16131
rect 622 12274 680 12275
rect 622 12273 623 12274
rect 679 12273 680 12274
rect 748 15663 749 15664
rect 805 15663 806 15664
rect 748 15662 806 15663
rect 622 12236 623 12237
rect 679 12236 680 12237
rect 622 12235 680 12236
rect 1126 16169 1184 16170
rect 1126 16168 1127 16169
rect 1183 16168 1184 16169
rect 1378 16169 1436 16170
rect 1378 16168 1379 16169
rect 1435 16168 1436 16169
rect 1630 16169 1688 16170
rect 1630 16168 1631 16169
rect 1687 16168 1688 16169
rect 1882 16169 1937 16170
rect 1882 16168 1883 16169
rect 1936 16168 1937 16169
rect 1000 15701 1058 15702
rect 1000 15700 1001 15701
rect 1057 15700 1058 15701
rect 1126 16131 1127 16132
rect 1183 16131 1184 16132
rect 1126 16130 1184 16131
rect 1378 16131 1379 16132
rect 1435 16131 1436 16132
rect 1378 16130 1436 16131
rect 874 12274 932 12275
rect 874 12273 875 12274
rect 931 12273 932 12274
rect 1000 15663 1001 15664
rect 1057 15663 1058 15664
rect 1000 15662 1058 15663
rect 496 11806 554 11807
rect 496 11805 497 11806
rect 553 11805 554 11806
rect 748 11806 806 11807
rect 748 11805 749 11806
rect 805 11805 806 11806
rect 874 12236 875 12237
rect 931 12236 932 12237
rect 874 12235 932 12236
rect 496 11768 497 11769
rect 553 11768 554 11769
rect 496 11767 554 11768
rect 748 11768 749 11769
rect 805 11768 806 11769
rect 748 11767 806 11768
rect 1630 16131 1631 16132
rect 1687 16131 1688 16132
rect 1630 16130 1688 16131
rect 1126 12274 1184 12275
rect 1126 12273 1127 12274
rect 1183 12273 1184 12274
rect 1882 16131 1883 16132
rect 1936 16131 1937 16132
rect 1882 16130 1937 16131
rect 1378 12274 1436 12275
rect 1378 12273 1379 12274
rect 1435 12273 1436 12274
rect 1630 12274 1688 12275
rect 1630 12273 1631 12274
rect 1687 12273 1688 12274
rect 1882 12274 1937 12275
rect 1882 12273 1883 12274
rect 1936 12273 1937 12274
rect 1000 11806 1058 11807
rect 1000 11805 1001 11806
rect 1057 11805 1058 11806
rect 1126 12236 1127 12237
rect 1183 12236 1184 12237
rect 1126 12235 1184 12236
rect 1378 12236 1379 12237
rect 1435 12236 1436 12237
rect 1378 12235 1436 12236
rect 874 8379 932 8380
rect 874 8378 875 8379
rect 931 8378 932 8379
rect 1000 11768 1001 11769
rect 1057 11768 1058 11769
rect 1000 11767 1058 11768
rect 496 7911 554 7912
rect 496 7910 497 7911
rect 553 7910 554 7911
rect 748 7911 806 7912
rect 748 7910 749 7911
rect 805 7910 806 7911
rect 874 8341 875 8342
rect 931 8341 932 8342
rect 874 8340 932 8341
rect 496 7873 497 7874
rect 553 7873 554 7874
rect 496 7872 554 7873
rect 748 7873 749 7874
rect 805 7873 806 7874
rect 748 7872 806 7873
rect 1630 12236 1631 12237
rect 1687 12236 1688 12237
rect 1630 12235 1688 12236
rect 1126 8379 1184 8380
rect 1126 8378 1127 8379
rect 1183 8378 1184 8379
rect 1882 12236 1883 12237
rect 1936 12236 1937 12237
rect 1882 12235 1937 12236
rect 1378 8379 1436 8380
rect 1378 8378 1379 8379
rect 1435 8378 1436 8379
rect 1630 8379 1688 8380
rect 1630 8378 1631 8379
rect 1687 8378 1688 8379
rect 1882 8379 1937 8380
rect 1882 8378 1883 8379
rect 1936 8378 1937 8379
rect 1000 7911 1058 7912
rect 1000 7910 1001 7911
rect 1057 7910 1058 7911
rect 1126 8341 1127 8342
rect 1183 8341 1184 8342
rect 1126 8340 1184 8341
rect 1378 8341 1379 8342
rect 1435 8341 1436 8342
rect 1378 8340 1436 8341
rect 874 4484 932 4485
rect 874 4483 875 4484
rect 931 4483 932 4484
rect 1000 7873 1001 7874
rect 1057 7873 1058 7874
rect 1000 7872 1058 7873
rect 874 4446 875 4447
rect 931 4446 932 4447
rect 874 4445 932 4446
rect 1630 8341 1631 8342
rect 1687 8341 1688 8342
rect 1630 8340 1688 8341
rect 1882 8341 1883 8342
rect 1936 8341 1937 8342
rect 1882 8340 1937 8341
rect 1378 4504 1436 4505
rect 1378 4503 1379 4504
rect 1435 4503 1436 4504
rect 2961 10825 4361 10826
rect 2961 10824 2962 10825
rect 4360 10824 4361 10825
rect 2961 10787 2962 10788
rect 4360 10787 4361 10788
rect 2961 10786 4361 10787
rect 4394 10762 4396 10763
rect 4432 10762 4434 10763
rect 4394 10712 4395 10762
rect 4433 10712 4434 10762
rect 4394 10711 4396 10712
rect 4432 10711 4434 10712
rect 2961 10687 4361 10688
rect 2961 10686 2962 10687
rect 4360 10686 4361 10687
rect 2961 10649 2962 10650
rect 4360 10649 4361 10650
rect 2961 10648 4361 10649
rect 2854 8676 4612 8677
rect 2854 8675 2855 8676
rect 4611 8675 4612 8676
rect 2854 8638 2855 8639
rect 4611 8638 4612 8639
rect 2854 8637 4612 8638
rect 2854 6665 3021 6666
rect 3105 6665 4361 6666
rect 2854 6664 2855 6665
rect 3020 6664 3021 6665
rect 3105 6664 3106 6665
rect 4360 6664 4361 6665
rect 2854 6627 2855 6628
rect 3020 6627 3021 6628
rect 3105 6627 3106 6628
rect 4360 6627 4361 6628
rect 2854 6626 3021 6627
rect 3105 6626 4361 6627
rect 4394 6602 4396 6603
rect 4432 6602 4434 6603
rect 4394 6552 4395 6602
rect 4433 6552 4434 6602
rect 4394 6551 4396 6552
rect 4432 6551 4434 6552
rect 3105 6527 4361 6528
rect 3105 6526 3106 6527
rect 4360 6526 4361 6527
rect 3105 6489 3106 6490
rect 4360 6489 4361 6490
rect 5081 10825 6481 10826
rect 5081 10824 5082 10825
rect 6480 10824 6481 10825
rect 5081 10787 5082 10788
rect 6480 10787 6481 10788
rect 5081 10786 6481 10787
rect 5008 10762 5010 10763
rect 5046 10762 5048 10763
rect 5008 10712 5009 10762
rect 5047 10712 5048 10762
rect 5008 10711 5010 10712
rect 5046 10711 5048 10712
rect 5081 10687 6481 10688
rect 5081 10686 5082 10687
rect 6480 10686 6481 10687
rect 5081 10649 5082 10650
rect 6480 10649 6481 10650
rect 5081 10648 6481 10649
rect 4830 8676 6588 8677
rect 4830 8675 4831 8676
rect 6587 8675 6588 8676
rect 4830 8638 4831 8639
rect 6587 8638 6588 8639
rect 4830 8637 6588 8638
rect 5081 6665 6337 6666
rect 6421 6665 6588 6666
rect 5081 6664 5082 6665
rect 6336 6664 6337 6665
rect 6421 6664 6422 6665
rect 6587 6664 6588 6665
rect 5081 6627 5082 6628
rect 6336 6627 6337 6628
rect 6421 6627 6422 6628
rect 6587 6627 6588 6628
rect 5081 6626 6337 6627
rect 6421 6626 6588 6627
rect 5008 6602 5010 6603
rect 5046 6602 5048 6603
rect 5008 6552 5009 6602
rect 5047 6552 5048 6602
rect 5008 6551 5010 6552
rect 5046 6551 5048 6552
rect 5081 6527 6337 6528
rect 5081 6526 5082 6527
rect 6336 6526 6337 6527
rect 3105 6488 4361 6489
rect 5081 6489 5082 6490
rect 6336 6489 6337 6490
rect 5081 6488 6337 6489
rect 1940 5569 1942 5570
rect 1940 5453 1941 5569
rect 1940 5452 1942 5453
rect 1978 5569 1980 5570
rect 1979 5453 1980 5569
rect 1978 5452 1980 5453
rect 1630 4504 1688 4505
rect 1630 4503 1631 4504
rect 1687 4503 1688 4504
rect 1126 4432 1184 4433
rect 1126 4431 1127 4432
rect 1183 4431 1184 4432
rect 1126 4394 1127 4395
rect 1183 4394 1184 4395
rect 1126 4393 1184 4394
rect 1378 4466 1379 4467
rect 1435 4466 1436 4467
rect 1378 4465 1436 4466
rect 1630 4466 1631 4467
rect 1687 4466 1688 4467
rect 1630 4465 1688 4466
rect 2134 4504 2192 4505
rect 2134 4503 2135 4504
rect 2191 4503 2192 4504
rect 2134 4466 2135 4467
rect 2191 4466 2192 4467
rect 2134 4465 2192 4466
rect 2386 4504 2444 4505
rect 2386 4503 2387 4504
rect 2443 4503 2444 4504
rect 2386 4466 2387 4467
rect 2443 4466 2444 4467
rect 2386 4465 2444 4466
rect 5528 4602 5580 4603
rect 5528 4601 5529 4602
rect 5579 4601 5580 4602
rect 5528 4564 5529 4565
rect 5579 4564 5580 4565
rect 5528 4563 5580 4564
rect 1882 4117 1940 4118
rect 2134 4117 2192 4118
rect 2386 4117 2444 4118
rect 2638 4117 2696 4118
rect 1882 4116 1883 4117
rect 1939 4116 1940 4117
rect 2134 4116 2135 4117
rect 2191 4116 2192 4117
rect 2386 4116 2387 4117
rect 2443 4116 2444 4117
rect 2638 4116 2639 4117
rect 2695 4116 2696 4117
rect 496 3942 554 3943
rect 496 3941 497 3942
rect 553 3941 554 3942
rect 496 3904 497 3905
rect 553 3904 554 3905
rect 496 3903 554 3904
rect 748 3942 806 3943
rect 748 3941 749 3942
rect 805 3941 806 3942
rect 748 3904 749 3905
rect 805 3904 806 3905
rect 748 3903 806 3904
rect 622 589 664 590
rect 622 588 623 589
rect 663 588 664 589
rect 622 551 623 552
rect 663 551 664 552
rect 622 550 664 551
rect 1252 3942 1310 3943
rect 1252 3941 1253 3942
rect 1309 3941 1310 3942
rect 1252 3904 1253 3905
rect 1309 3904 1310 3905
rect 1252 3903 1310 3904
rect 1126 589 1168 590
rect 1126 588 1127 589
rect 1167 588 1168 589
rect 1126 551 1127 552
rect 1167 551 1168 552
rect 1126 550 1168 551
rect 1504 3942 1562 3943
rect 1504 3941 1505 3942
rect 1561 3941 1562 3942
rect 1504 3904 1505 3905
rect 1561 3904 1562 3905
rect 1504 3903 1562 3904
rect 1378 589 1420 590
rect 1378 588 1379 589
rect 1419 588 1420 589
rect 1378 551 1379 552
rect 1419 551 1420 552
rect 1378 550 1420 551
rect 1756 3942 1814 3943
rect 1756 3941 1757 3942
rect 1813 3941 1814 3942
rect 1882 4079 1883 4080
rect 1939 4079 1940 4080
rect 1882 4078 1940 4079
rect 1882 3942 1940 3943
rect 1882 3941 1883 3942
rect 1939 3941 1940 3942
rect 2008 3942 2066 3943
rect 2008 3941 2009 3942
rect 2065 3941 2066 3942
rect 2134 4079 2135 4080
rect 2191 4079 2192 4080
rect 2134 4078 2192 4079
rect 1756 3904 1757 3905
rect 1813 3904 1814 3905
rect 1756 3903 1814 3904
rect 1630 589 1672 590
rect 1630 588 1631 589
rect 1671 588 1672 589
rect 1630 551 1631 552
rect 1671 551 1672 552
rect 1630 550 1672 551
rect 1882 3904 1883 3905
rect 1939 3904 1940 3905
rect 1882 3903 1940 3904
rect 2008 3904 2009 3905
rect 2065 3904 2066 3905
rect 2008 3903 2066 3904
rect 2260 3942 2318 3943
rect 2260 3941 2261 3942
rect 2317 3941 2318 3942
rect 2386 4079 2387 4080
rect 2443 4079 2444 4080
rect 2386 4078 2444 4079
rect 2260 3904 2261 3905
rect 2317 3904 2318 3905
rect 2260 3903 2318 3904
rect 2512 3942 2570 3943
rect 2512 3941 2513 3942
rect 2569 3941 2570 3942
rect 2638 4079 2639 4080
rect 2695 4079 2696 4080
rect 2638 4078 2696 4079
rect 2638 3942 2696 3943
rect 2638 3941 2639 3942
rect 2695 3941 2696 3942
rect 2890 4064 2948 4065
rect 2890 4063 2891 4064
rect 2947 4063 2948 4064
rect 2764 3942 2822 3943
rect 2764 3941 2765 3942
rect 2821 3941 2822 3942
rect 2890 4026 2891 4027
rect 2947 4026 2948 4027
rect 2890 4025 2948 4026
rect 2512 3904 2513 3905
rect 2569 3904 2570 3905
rect 2512 3903 2570 3904
rect 2638 3904 2639 3905
rect 2695 3904 2696 3905
rect 2638 3903 2696 3904
rect 2764 3904 2765 3905
rect 2821 3904 2822 3905
rect 2764 3903 2822 3904
rect 2890 3889 2948 3890
rect 2890 3888 2891 3889
rect 2947 3888 2948 3889
rect 2890 3851 2891 3852
rect 2947 3851 2948 3852
rect 2890 3850 2948 3851
<< via1 >>
rect 138 27869 190 27878
rect 202 27869 254 27878
rect 266 27869 318 27878
rect 138 27835 172 27869
rect 172 27835 190 27869
rect 202 27835 206 27869
rect 206 27835 244 27869
rect 244 27835 254 27869
rect 266 27835 278 27869
rect 278 27835 318 27869
rect 138 27826 190 27835
rect 202 27826 254 27835
rect 266 27826 318 27835
rect 540 27667 656 27783
rect 724 27731 776 27783
rect 796 27731 848 27783
rect 868 27731 920 27783
rect 940 27731 992 27783
rect 1011 27731 1063 27783
rect 1082 27731 1134 27783
rect 1153 27731 1205 27783
rect 1224 27731 1276 27783
rect 724 27667 776 27719
rect 796 27667 848 27719
rect 868 27667 920 27719
rect 940 27667 992 27719
rect 1011 27667 1063 27719
rect 1082 27667 1134 27719
rect 1153 27667 1205 27719
rect 1224 27667 1276 27719
rect 1344 27667 1460 27783
rect 1691 27746 1743 27798
rect 1755 27746 1807 27798
rect 1819 27746 1871 27798
rect 1802 27666 1854 27718
rect 1866 27666 1918 27718
rect 1930 27666 1982 27718
rect 1016 27585 1068 27637
rect 1080 27585 1132 27637
rect 1144 27585 1196 27637
rect 1208 27585 1260 27637
rect 1344 27585 1396 27637
rect 1408 27585 1460 27637
rect 1802 27585 1854 27637
rect 1866 27585 1918 27637
rect 1930 27585 1982 27637
rect 2045 8276 2097 8328
rect 2045 8212 2097 8264
rect 1965 8092 2017 8144
rect 1965 8028 2017 8080
rect 2029 8028 2081 8080
rect 3015 10855 3067 10907
rect 3079 10855 3131 10907
rect 3143 10855 3195 10907
rect 3207 10855 3259 10907
rect 3429 10855 3481 10907
rect 3493 10855 3545 10907
rect 3557 10855 3609 10907
rect 3621 10855 3673 10907
rect 3685 10855 3737 10907
rect 3749 10855 3801 10907
rect 3973 10855 4025 10907
rect 4037 10855 4089 10907
rect 4101 10855 4153 10907
rect 4165 10855 4217 10907
rect 4229 10855 4281 10907
rect 4293 10855 4345 10907
rect 4357 10855 4409 10907
rect 5109 10855 5161 10907
rect 5173 10855 5225 10907
rect 5237 10855 5289 10907
rect 5301 10855 5353 10907
rect 5365 10855 5417 10907
rect 5429 10855 5481 10907
rect 5637 10855 5689 10907
rect 5701 10855 5753 10907
rect 5765 10855 5817 10907
rect 5829 10855 5881 10907
rect 5893 10855 5945 10907
rect 5957 10855 6009 10907
rect 6021 10855 6073 10907
rect 6269 10855 6321 10907
rect 6333 10855 6385 10907
rect 6397 10855 6449 10907
rect 6461 10855 6513 10907
rect 6525 10855 6577 10907
rect 6589 10855 6641 10907
rect 6653 10855 6705 10907
rect 4474 10672 4590 10788
rect 2906 6496 2958 6548
rect 4474 6526 4590 6642
rect 2906 6432 2958 6484
rect 4846 10672 4962 10788
rect 4846 6526 4962 6642
rect 3143 6407 3195 6459
rect 3207 6407 3259 6459
rect 3424 6407 3476 6459
rect 3488 6407 3540 6459
rect 3552 6407 3604 6459
rect 3616 6407 3668 6459
rect 3973 6407 4025 6459
rect 4037 6407 4089 6459
rect 4101 6407 4153 6459
rect 4165 6407 4217 6459
rect 4229 6407 4281 6459
rect 4293 6407 4345 6459
rect 4357 6407 4409 6459
rect 5109 6407 5161 6459
rect 5173 6407 5225 6459
rect 5237 6407 5289 6459
rect 5301 6407 5353 6459
rect 5777 6407 5829 6459
rect 5841 6407 5893 6459
rect 5905 6407 5957 6459
rect 5969 6407 6021 6459
rect 6033 6407 6085 6459
rect 5600 6321 5652 6373
rect 5664 6321 5716 6373
rect 2325 6192 2377 6229
rect 2325 6177 2334 6192
rect 2334 6177 2368 6192
rect 2368 6177 2377 6192
rect 2325 6158 2334 6165
rect 2334 6158 2368 6165
rect 2368 6158 2377 6165
rect 2325 6113 2377 6158
rect 2513 6107 2565 6159
rect 2577 6107 2629 6159
rect 6259 6107 6311 6159
rect 6323 6107 6375 6159
rect 4996 6017 5048 6069
rect 5327 6027 5379 6079
rect 5391 6027 5443 6079
rect 2494 5947 2546 5999
rect 4996 5953 5048 6005
rect 6000 5947 6052 5999
rect 6064 5947 6116 5999
rect 2494 5883 2546 5935
rect 3029 5861 3081 5913
rect 5006 5867 5058 5919
rect 5070 5867 5122 5919
rect 3029 5797 3081 5849
rect 5614 5793 5666 5845
rect 5678 5793 5730 5845
rect 3246 5682 3298 5734
rect 3310 5682 3362 5734
rect 3144 5498 3260 5574
rect 5608 5522 5660 5574
rect 3144 5464 3153 5498
rect 3153 5464 3187 5498
rect 3187 5464 3260 5498
rect 3144 5458 3260 5464
rect 5608 5458 5660 5510
rect 3642 4416 3758 4596
rect 5172 4416 5288 4596
rect 5528 4453 5580 4505
rect 5528 4389 5580 4441
rect 2896 4135 2948 4187
rect 5534 4141 5586 4193
rect 5598 4141 5650 4193
rect 373 492 425 493
rect 373 458 382 492
rect 382 458 416 492
rect 416 458 425 492
rect 373 441 425 458
rect 373 420 425 429
rect 373 386 382 420
rect 382 386 416 420
rect 416 386 425 420
rect 373 377 425 386
rect 499 492 551 493
rect 499 458 508 492
rect 508 458 542 492
rect 542 458 551 492
rect 499 441 551 458
rect 499 420 551 429
rect 499 386 508 420
rect 508 386 542 420
rect 542 386 551 420
rect 499 377 551 386
rect 2896 4071 2948 4123
rect 3020 492 3072 496
rect 3020 458 3028 492
rect 3028 458 3062 492
rect 3062 458 3072 492
rect 3020 444 3072 458
rect 3020 420 3072 432
rect 3020 386 3028 420
rect 3028 386 3062 420
rect 3062 386 3072 420
rect 3020 380 3072 386
rect 735 210 787 262
rect 799 210 851 262
rect 863 210 915 262
rect 1011 210 1063 262
rect 1075 210 1127 262
rect 1139 210 1191 262
rect 1344 136 1460 252
rect 499 -195 551 -143
rect 499 -259 551 -207
rect 2266 -246 2318 -194
rect 2330 -246 2382 -194
rect 3054 -176 3106 -124
rect 499 -323 551 -271
rect 3054 -240 3106 -188
rect 2696 -326 2748 -274
rect 2760 -326 2812 -274
rect 1976 -588 2028 -536
rect 2040 -588 2092 -536
rect 2104 -560 2156 -536
rect 2168 -560 2220 -536
rect 3139 -554 3191 -536
rect 3203 -554 3255 -536
rect 2104 -588 2149 -560
rect 2149 -588 2156 -560
rect 2168 -588 2183 -560
rect 2183 -588 2220 -560
rect 3139 -588 3170 -554
rect 3170 -588 3191 -554
rect 3203 -588 3204 -554
rect 3204 -588 3243 -554
rect 3243 -588 3255 -554
rect 2451 -639 2503 -627
rect 2451 -673 2455 -639
rect 2455 -673 2489 -639
rect 2489 -673 2503 -639
rect 2451 -679 2503 -673
rect 2515 -639 2567 -627
rect 2515 -673 2527 -639
rect 2527 -673 2561 -639
rect 2561 -673 2567 -639
rect 2515 -679 2567 -673
rect 2607 -679 2659 -627
rect 2671 -679 2723 -627
rect 2260 -719 2312 -713
rect 2696 -719 2748 -707
rect 2260 -753 2266 -719
rect 2266 -753 2300 -719
rect 2300 -753 2312 -719
rect 2696 -753 2698 -719
rect 2698 -753 2732 -719
rect 2732 -753 2748 -719
rect 2260 -765 2312 -753
rect 2696 -759 2748 -753
rect 2760 -759 2812 -707
rect 3054 -765 3106 -713
rect 2260 -791 2312 -777
rect 2260 -825 2266 -791
rect 2266 -825 2300 -791
rect 2300 -825 2312 -791
rect 2260 -829 2312 -825
rect 2837 -818 3017 -814
rect 2837 -852 2914 -818
rect 2914 -852 2948 -818
rect 2948 -852 3017 -818
rect 3054 -829 3106 -777
rect 2837 -890 3017 -852
rect 2837 -924 2914 -890
rect 2914 -924 2948 -890
rect 2948 -924 3017 -890
rect 2837 -930 3017 -924
rect 3424 -930 3604 -814
rect 1976 -1029 2028 -977
rect 2040 -1029 2092 -977
rect 2104 -989 2156 -977
rect 2168 -989 2220 -977
rect 2104 -1023 2149 -989
rect 2149 -1023 2156 -989
rect 2168 -1023 2183 -989
rect 2183 -1023 2220 -989
rect 3139 -995 3191 -977
rect 3203 -995 3255 -977
rect 2104 -1029 2156 -1023
rect 2168 -1029 2220 -1023
rect 3139 -1029 3170 -995
rect 3170 -1029 3191 -995
rect 3203 -1029 3204 -995
rect 3204 -1029 3243 -995
rect 3243 -1029 3255 -995
<< metal2 >>
tri 108 27878 126 27896 se
rect 126 27878 478 27896
tri 59 27829 108 27878 se
rect 108 27829 138 27878
rect 59 27826 138 27829
rect 190 27826 202 27878
rect 254 27826 266 27878
rect 318 27826 478 27878
rect 59 27784 478 27826
rect 534 27783 662 27784
tri 441 27667 534 27760 se
rect 534 27667 540 27783
rect 656 27667 662 27783
tri 440 27666 441 27667 se
rect 441 27666 662 27667
tri 411 27637 440 27666 se
rect 440 27644 662 27666
rect 440 27637 655 27644
tri 655 27637 662 27644 nw
rect 718 27783 1282 27784
rect 718 27731 724 27783
rect 776 27731 796 27783
rect 848 27731 868 27783
rect 920 27731 940 27783
rect 992 27731 1011 27783
rect 1063 27731 1082 27783
rect 1134 27731 1153 27783
rect 1205 27731 1224 27783
rect 1276 27731 1282 27783
rect 718 27719 1282 27731
rect 718 27667 724 27719
rect 776 27667 796 27719
rect 848 27667 868 27719
rect 920 27667 940 27719
rect 992 27667 1011 27719
rect 1063 27667 1082 27719
rect 1134 27667 1153 27719
rect 1205 27667 1224 27719
rect 1276 27667 1282 27719
rect 718 27637 1282 27667
tri 359 27585 411 27637 se
rect 411 27585 603 27637
tri 603 27585 655 27637 nw
rect 718 27585 1016 27637
rect 1068 27585 1080 27637
rect 1132 27585 1144 27637
rect 1196 27585 1208 27637
rect 1260 27585 1282 27637
tri 344 27570 359 27585 se
rect 359 27570 588 27585
tri 588 27570 603 27585 nw
tri 290 27516 344 27570 se
rect 344 27516 534 27570
tri 534 27516 588 27570 nw
tri 664 27516 718 27570 se
rect 718 27516 1282 27585
tri 59 27285 290 27516 se
rect 290 27386 404 27516
tri 404 27386 534 27516 nw
tri 534 27386 664 27516 se
rect 664 27386 1282 27516
rect 290 27285 381 27386
tri 381 27363 404 27386 nw
tri 511 27363 534 27386 se
rect 534 27363 1282 27386
rect 59 4916 381 27285
tri 59 4620 355 4916 ne
rect 355 4703 381 4916
tri 459 27311 511 27363 se
rect 511 27311 1282 27363
rect 459 27224 1282 27311
rect 459 26634 658 27224
tri 658 27097 785 27224 nw
tri 985 27126 1083 27224 ne
tri 1054 26897 1083 26926 se
rect 1083 26897 1282 27224
tri 658 26634 921 26897 sw
rect 459 4785 921 26634
tri 1010 26853 1054 26897 se
rect 1054 26853 1282 26897
tri 966 5953 1010 5997 se
rect 1010 5953 1282 26853
rect 966 5143 1282 5953
tri 966 5104 1005 5143 ne
tri 459 4783 461 4785 ne
rect 461 4783 921 4785
tri 381 4703 461 4783 sw
tri 461 4703 541 4783 ne
rect 541 4703 921 4783
rect 355 4676 461 4703
tri 461 4676 488 4703 sw
tri 541 4676 568 4703 ne
rect 568 4676 921 4703
rect 355 4620 488 4676
tri 488 4620 544 4676 sw
tri 568 4620 624 4676 ne
tri 355 4596 379 4620 ne
rect 379 4596 544 4620
tri 544 4596 568 4620 sw
tri 379 4594 381 4596 ne
rect 381 4594 568 4596
tri 381 4540 435 4594 ne
rect 59 3706 379 4516
rect 59 3682 355 3706
tri 355 3682 379 3706 nw
rect 59 3602 275 3682
tri 275 3602 355 3682 nw
tri 355 3602 435 3682 se
rect 435 3626 568 4594
rect 435 3602 544 3626
tri 544 3602 568 3626 nw
rect 59 3575 248 3602
tri 248 3575 275 3602 nw
tri 328 3575 355 3602 se
rect 355 3575 488 3602
rect 59 150 192 3575
tri 192 3519 248 3575 nw
tri 272 3519 328 3575 se
rect 328 3546 488 3575
tri 488 3546 544 3602 nw
tri 568 3546 624 3602 se
rect 624 3546 921 4676
rect 328 3519 461 3546
tri 461 3519 488 3546 nw
tri 541 3519 568 3546 se
rect 568 3519 921 3546
tri 248 3495 272 3519 se
rect 272 3495 437 3519
tri 437 3495 461 3519 nw
tri 517 3495 541 3519 se
rect 541 3495 921 3519
rect 248 584 381 3495
tri 381 3439 437 3495 nw
tri 461 3439 517 3495 se
rect 517 3439 921 3495
rect 248 514 311 584
tri 311 514 381 584 nw
tri 459 3437 461 3439 se
rect 461 3437 921 3439
rect 459 671 921 3437
tri 966 3158 1005 3197 se
rect 1005 3158 1282 5143
rect 966 2348 1282 3158
tri 966 2309 1005 2348 ne
tri 459 514 616 671 ne
rect 248 268 300 514
tri 300 503 311 514 nw
rect 370 493 428 499
rect 370 441 373 493
rect 425 441 428 493
rect 370 429 428 441
rect 370 377 373 429
rect 425 377 428 429
tri 192 150 217 175 sw
tri 345 150 370 175 se
rect 370 150 428 377
rect 59 86 428 150
tri 59 -84 229 86 ne
rect 229 -65 428 86
rect 229 -84 409 -65
tri 409 -84 428 -65 nw
rect 499 493 551 499
rect 499 429 551 441
rect 499 -143 551 377
rect 616 262 921 671
rect 616 210 735 262
rect 787 210 799 262
rect 851 210 863 262
rect 915 210 921 262
rect 616 62 921 210
rect 1005 262 1282 2348
rect 1005 210 1011 262
rect 1063 210 1075 262
rect 1127 210 1139 262
rect 1191 210 1282 262
rect 1005 62 1282 210
rect 1338 27783 1477 27784
rect 1338 27667 1344 27783
rect 1460 27667 1477 27783
rect 1685 27746 1691 27798
rect 1743 27746 1755 27798
rect 1807 27746 1819 27798
rect 1871 27746 1877 27798
rect 1338 27637 1477 27667
rect 1338 27585 1344 27637
rect 1396 27585 1408 27637
rect 1460 27585 1477 27637
rect 1338 11385 1477 27585
rect 1793 27666 1802 27718
rect 1854 27666 1866 27718
rect 1918 27666 1930 27718
rect 1982 27666 2017 27718
rect 1793 27637 2017 27666
rect 1793 27585 1802 27637
rect 1854 27585 1866 27637
rect 1918 27585 1930 27637
rect 1982 27585 2017 27637
rect 1793 11533 2017 27585
tri 1477 11385 1535 11443 sw
tri 1735 11385 1793 11443 se
rect 1793 11385 1934 11533
tri 1934 11450 2017 11533 nw
rect 1338 10575 1934 11385
rect 1338 3745 1477 10575
tri 1477 10517 1535 10575 nw
tri 1735 10517 1793 10575 ne
rect 1793 10517 1934 10575
tri 1793 10512 1798 10517 ne
rect 1798 10512 1934 10517
tri 1934 10512 2017 10595 sw
tri 1798 10492 1818 10512 ne
rect 1818 8150 2017 10512
rect 2045 8328 2097 11017
rect 2045 8264 2097 8276
rect 2045 8206 2097 8212
tri 2017 8150 2042 8175 sw
rect 1818 8144 2042 8150
rect 1818 8092 1965 8144
rect 2017 8111 2042 8144
tri 2042 8111 2081 8150 sw
rect 2017 8092 2081 8111
rect 1818 8080 2081 8092
rect 1818 8028 1965 8080
rect 2017 8028 2029 8080
tri 1749 3791 1818 3860 se
rect 1818 3791 2081 8028
tri 2121 7311 2125 7315 se
rect 2125 7311 2432 11017
tri 2432 7311 2437 7316 sw
rect 2121 6501 2437 7311
tri 2121 6497 2125 6501 ne
rect 2125 6497 2433 6501
tri 2433 6497 2437 6501 nw
rect 2125 6229 2432 6497
tri 2432 6496 2433 6497 nw
rect 2488 6386 2850 11017
rect 2906 6648 2958 11017
rect 3014 10907 3260 11017
rect 3014 10855 3015 10907
rect 3067 10855 3079 10907
rect 3131 10855 3143 10907
rect 3195 10855 3207 10907
rect 3259 10855 3260 10907
rect 3014 6719 3260 10855
tri 3014 6678 3055 6719 ne
rect 3055 6678 3260 6719
tri 2906 6642 2912 6648 ne
rect 2912 6642 2958 6648
tri 2958 6642 2994 6678 sw
tri 3055 6642 3091 6678 ne
rect 3091 6642 3260 6678
tri 2912 6631 2923 6642 ne
rect 2923 6631 2994 6642
tri 2994 6631 3005 6642 sw
tri 3091 6631 3102 6642 ne
rect 3102 6631 3260 6642
tri 2923 6596 2958 6631 ne
rect 2958 6622 3005 6631
tri 3005 6622 3014 6631 sw
tri 3102 6622 3111 6631 ne
rect 3111 6622 3260 6631
rect 2958 6596 3014 6622
tri 2958 6549 3005 6596 ne
rect 3005 6590 3014 6596
tri 3014 6590 3046 6622 sw
tri 3111 6590 3143 6622 ne
rect 3005 6549 3046 6590
tri 3046 6549 3087 6590 sw
tri 3005 6548 3006 6549 ne
rect 3006 6548 3087 6549
tri 2488 6373 2501 6386 ne
rect 2501 6373 2850 6386
tri 2501 6321 2553 6373 ne
rect 2553 6321 2850 6373
rect 2125 6177 2325 6229
rect 2377 6177 2432 6229
tri 2553 6183 2691 6321 ne
rect 2125 6165 2432 6177
rect 2125 6113 2325 6165
rect 2377 6113 2432 6165
rect 2125 4774 2432 6113
rect 2507 6107 2513 6159
rect 2565 6107 2577 6159
rect 2629 6107 2635 6159
tri 2507 6079 2535 6107 ne
rect 2535 6079 2635 6107
tri 2535 6069 2545 6079 ne
rect 2545 6069 2635 6079
tri 2545 6034 2580 6069 ne
rect 2488 5947 2494 5999
rect 2546 5947 2552 5999
rect 2488 5935 2552 5947
rect 2488 5883 2494 5935
rect 2546 5883 2552 5935
tri 1724 3766 1749 3791 se
rect 1749 3766 2081 3791
tri 1703 3745 1724 3766 se
rect 1724 3745 2081 3766
rect 1338 252 1466 3745
tri 1466 3734 1477 3745 nw
tri 1692 3734 1703 3745 se
rect 1703 3734 2081 3745
rect 1338 136 1344 252
rect 1460 136 1466 252
rect 1338 62 1466 136
tri 1577 3619 1692 3734 se
rect 1692 3619 2081 3734
tri 2121 4517 2125 4521 se
rect 2125 4517 2432 4521
rect 2121 4516 2432 4517
tri 2432 4516 2437 4521 sw
rect 2121 3706 2437 4516
rect 2121 3705 2432 3706
tri 2121 3701 2125 3705 ne
rect 1577 62 2081 3619
tri 1577 -55 1694 62 ne
rect 1694 -55 2081 62
rect 2125 -16 2432 3705
tri 2432 3701 2437 3706 nw
tri 2432 100 2445 113 sw
tri 1694 -124 1763 -55 ne
rect 1763 -118 2081 -55
tri 2081 -118 2144 -55 sw
rect 1763 -124 2144 -118
tri 2144 -124 2150 -118 sw
tri 1763 -176 1815 -124 ne
rect 1815 -176 2150 -124
tri 2150 -176 2202 -124 sw
tri 1815 -188 1827 -176 ne
rect 1827 -188 2202 -176
tri 2202 -188 2214 -176 sw
tri 1827 -194 1833 -188 ne
rect 1833 -194 2214 -188
tri 2214 -194 2220 -188 sw
rect 499 -207 551 -195
tri 1833 -246 1885 -194 ne
rect 1885 -246 2220 -194
rect 499 -271 551 -259
tri 1885 -274 1913 -246 ne
rect 1913 -274 2220 -246
rect 499 -329 551 -323
tri 1913 -326 1965 -274 ne
rect 1965 -326 2220 -274
tri 1965 -329 1968 -326 ne
rect 1968 -329 2220 -326
tri 1968 -337 1976 -329 ne
rect 1976 -536 2220 -329
rect 2028 -588 2040 -536
rect 2092 -588 2104 -536
rect 2156 -588 2168 -536
rect 1976 -977 2220 -588
rect 2260 -246 2266 -194
rect 2318 -246 2330 -194
rect 2382 -246 2388 -194
rect 2260 -713 2312 -246
tri 2312 -271 2337 -246 nw
tri 2484 -588 2488 -584 se
rect 2488 -588 2543 5883
tri 2543 5874 2552 5883 nw
tri 2475 -597 2484 -588 se
rect 2484 -597 2543 -588
rect 2580 -588 2635 6069
rect 2691 3327 2850 6321
rect 2900 6496 2906 6548
rect 2958 6496 2964 6548
tri 3006 6531 3023 6548 ne
rect 2900 6484 2964 6496
rect 2900 6432 2906 6484
rect 2958 6432 2964 6484
tri 2896 4193 2900 4197 se
rect 2900 4193 2964 6432
rect 3023 5913 3087 6548
rect 3143 6459 3260 6622
rect 3195 6407 3207 6459
rect 3259 6407 3260 6459
rect 3143 6401 3260 6407
tri 3143 6373 3171 6401 ne
rect 3171 6373 3260 6401
tri 3171 6348 3196 6373 ne
rect 3023 5861 3029 5913
rect 3081 5861 3087 5913
rect 3023 5849 3087 5861
rect 3023 5797 3029 5849
rect 3081 5797 3087 5849
tri 3184 5810 3196 5822 se
rect 3196 5810 3260 6373
tri 3171 5797 3184 5810 se
rect 3184 5797 3260 5810
tri 3303 5797 3316 5810 se
rect 3316 5797 3368 11017
tri 3167 5793 3171 5797 se
rect 3171 5794 3260 5797
tri 3300 5794 3303 5797 se
rect 3303 5794 3368 5797
rect 3171 5793 3259 5794
tri 3259 5793 3260 5794 nw
tri 3299 5793 3300 5794 se
rect 3300 5793 3368 5794
tri 3108 5734 3167 5793 se
rect 3167 5754 3220 5793
tri 3220 5754 3259 5793 nw
tri 3260 5754 3299 5793 se
rect 3299 5754 3368 5793
rect 3167 5734 3200 5754
tri 3200 5734 3220 5754 nw
tri 3240 5734 3260 5754 se
rect 3260 5734 3368 5754
tri 3104 5730 3108 5734 se
rect 3108 5730 3196 5734
tri 3196 5730 3200 5734 nw
tri 3056 5682 3104 5730 se
rect 3104 5682 3148 5730
tri 3148 5682 3196 5730 nw
rect 3240 5682 3246 5734
rect 3298 5682 3310 5734
rect 3362 5682 3368 5734
rect 3424 10907 3806 11017
rect 3424 10855 3429 10907
rect 3481 10855 3493 10907
rect 3545 10855 3557 10907
rect 3609 10855 3621 10907
rect 3673 10855 3685 10907
rect 3737 10855 3749 10907
rect 3801 10855 3806 10907
rect 3424 6459 3806 10855
rect 3476 6407 3488 6459
rect 3540 6407 3552 6459
rect 3604 6407 3616 6459
rect 3668 6407 3806 6459
rect 2896 4187 2964 4193
rect 2948 4135 2964 4187
rect 2896 4123 2964 4135
rect 2948 4071 2964 4123
rect 2896 4065 2964 4071
tri 3014 5640 3056 5682 se
rect 3056 5640 3106 5682
tri 3106 5640 3148 5682 nw
tri 2850 3327 2881 3358 sw
tri 2983 3327 3014 3358 se
rect 3014 3327 3078 5640
tri 3078 5612 3106 5640 nw
rect 2691 496 3078 3327
rect 2691 444 3020 496
rect 3072 444 3078 496
rect 2691 432 3078 444
rect 2691 380 3020 432
rect 3072 380 3078 432
rect 2691 153 3026 380
tri 3026 328 3078 380 nw
rect 3134 5574 3260 5580
rect 3134 5458 3144 5574
tri 2704 11 2846 153 ne
rect 2690 -326 2696 -274
rect 2748 -326 2760 -274
rect 2812 -326 2818 -274
tri 2741 -351 2766 -326 ne
tri 2635 -588 2652 -571 sw
rect 2580 -594 2652 -588
tri 2580 -597 2583 -594 ne
rect 2583 -597 2652 -594
tri 2445 -627 2475 -597 se
rect 2475 -615 2543 -597
tri 2543 -615 2561 -597 sw
tri 2583 -615 2601 -597 ne
rect 2475 -627 2561 -615
tri 2561 -627 2573 -615 sw
rect 2445 -679 2451 -627
rect 2503 -679 2515 -627
rect 2567 -679 2573 -627
rect 2601 -627 2652 -597
tri 2652 -627 2691 -588 sw
rect 2601 -679 2607 -627
rect 2659 -679 2671 -627
rect 2723 -679 2729 -627
tri 2741 -707 2766 -682 se
rect 2766 -707 2818 -326
rect 2690 -759 2696 -707
rect 2748 -759 2760 -707
rect 2812 -759 2818 -707
rect 2260 -777 2312 -765
rect 2260 -835 2312 -829
tri 2837 -808 2846 -799 se
rect 2846 -808 3026 153
rect 2837 -814 3026 -808
rect 3017 -930 3026 -814
rect 3054 -124 3106 -118
rect 3054 -188 3106 -176
rect 3054 -713 3106 -240
rect 3054 -777 3106 -765
rect 3054 -835 3106 -829
rect 3134 -536 3260 5458
rect 3424 4596 3806 6407
rect 3424 4416 3642 4596
rect 3758 4416 3806 4596
rect 3424 4274 3806 4416
rect 3862 10907 4412 11017
rect 3862 10855 3973 10907
rect 4025 10855 4037 10907
rect 4089 10855 4101 10907
rect 4153 10855 4165 10907
rect 4217 10855 4229 10907
rect 4281 10855 4293 10907
rect 4345 10855 4357 10907
rect 4409 10855 4412 10907
rect 3862 6459 4412 10855
rect 3862 6407 3973 6459
rect 4025 6407 4037 6459
rect 4089 6407 4101 6459
rect 4153 6407 4165 6459
rect 4217 6407 4229 6459
rect 4281 6407 4293 6459
rect 4345 6407 4357 6459
rect 4409 6407 4412 6459
rect 3862 4274 4412 6407
rect 4468 10788 4968 11017
rect 4468 10672 4474 10788
rect 4590 10672 4846 10788
rect 4962 10672 4968 10788
rect 4468 6642 4968 10672
rect 4468 6526 4474 6642
rect 4590 6526 4846 6642
rect 4962 6526 4968 6642
rect 4468 4917 4968 6526
rect 4996 6069 5048 11017
rect 5104 10907 5486 11017
rect 5104 10855 5109 10907
rect 5161 10855 5173 10907
rect 5225 10855 5237 10907
rect 5289 10855 5301 10907
rect 5353 10855 5365 10907
rect 5417 10855 5429 10907
rect 5481 10855 5486 10907
rect 5104 6551 5486 10855
rect 5622 10907 6085 11017
rect 5622 10855 5637 10907
rect 5689 10855 5701 10907
rect 5753 10855 5765 10907
rect 5817 10855 5829 10907
rect 5881 10855 5893 10907
rect 5945 10855 5957 10907
rect 6009 10855 6021 10907
rect 6073 10855 6085 10907
rect 5622 6789 6085 10855
tri 5622 6647 5764 6789 ne
rect 5104 6526 5461 6551
tri 5461 6526 5486 6551 nw
rect 5104 6465 5400 6526
tri 5400 6465 5461 6526 nw
rect 5104 6459 5394 6465
tri 5394 6459 5400 6465 nw
rect 5764 6459 6085 6789
rect 5104 6407 5109 6459
rect 5161 6407 5173 6459
rect 5225 6407 5237 6459
rect 5289 6407 5301 6459
rect 5353 6407 5391 6459
tri 5391 6456 5394 6459 nw
rect 5104 6203 5391 6407
rect 5764 6407 5777 6459
rect 5829 6407 5841 6459
rect 5893 6407 5905 6459
rect 5957 6407 5969 6459
rect 6021 6407 6033 6459
rect 5104 6159 5347 6203
tri 5347 6159 5391 6203 nw
rect 5528 6321 5600 6373
rect 5652 6321 5664 6373
rect 5716 6321 5722 6373
rect 5104 6157 5345 6159
tri 5345 6157 5347 6159 nw
tri 5104 6107 5154 6157 ne
rect 5154 6107 5295 6157
tri 5295 6107 5345 6157 nw
tri 5154 6105 5156 6107 ne
rect 4996 6005 5048 6017
rect 4996 5947 5048 5953
rect 5000 5867 5006 5919
rect 5058 5867 5070 5919
rect 5122 5867 5128 5919
tri 5000 5845 5022 5867 ne
rect 5022 5845 5128 5867
tri 5022 5797 5070 5845 ne
rect 5070 5797 5128 5845
tri 5070 5793 5074 5797 ne
rect 5074 5793 5128 5797
tri 5074 5791 5076 5793 ne
rect 4468 4602 4653 4917
tri 4653 4602 4968 4917 nw
rect 4468 4596 4647 4602
tri 4647 4596 4653 4602 nw
rect 4468 4274 4600 4596
tri 4600 4549 4647 4596 nw
tri 5065 4194 5076 4205 se
rect 5076 4194 5128 5793
rect 5156 4596 5293 6107
tri 5293 6105 5295 6107 nw
rect 5156 4416 5172 4596
rect 5288 4416 5293 4596
rect 5156 4274 5293 4416
rect 5321 6027 5327 6079
rect 5379 6027 5391 6079
rect 5443 6027 5449 6079
rect 5321 5999 5421 6027
tri 5421 5999 5449 6027 nw
rect 5065 4180 5128 4194
rect 5065 4133 5117 4180
tri 5117 4169 5128 4180 nw
rect 5321 4133 5373 5999
tri 5373 5951 5421 5999 nw
rect 5528 4505 5580 6321
tri 5580 6179 5722 6321 nw
rect 5764 6326 6085 6407
rect 5764 6321 6080 6326
tri 6080 6321 6085 6326 nw
rect 5764 6235 5994 6321
tri 5994 6235 6080 6321 nw
rect 5608 5793 5614 5845
rect 5666 5793 5678 5845
rect 5730 5793 5736 5845
rect 5608 5750 5693 5793
tri 5693 5750 5736 5793 nw
rect 5764 5750 5966 6235
tri 5966 6207 5994 6235 nw
rect 6141 6108 6193 11017
rect 6249 10907 6911 11017
rect 6249 10855 6269 10907
rect 6321 10855 6333 10907
rect 6385 10855 6397 10907
rect 6449 10855 6461 10907
rect 6513 10855 6525 10907
rect 6577 10855 6589 10907
rect 6641 10855 6653 10907
rect 6705 10855 6911 10907
rect 6249 10447 6911 10855
tri 6249 10075 6621 10447 ne
rect 6249 6766 6565 10051
rect 6621 7461 6911 10447
rect 6621 7421 6871 7461
tri 6871 7421 6911 7461 nw
tri 6911 7421 6967 7477 se
rect 6967 7421 7117 11017
rect 6621 7391 6841 7421
tri 6841 7391 6871 7421 nw
tri 6881 7391 6911 7421 se
rect 6911 7391 7117 7421
rect 6621 7351 6801 7391
tri 6801 7351 6841 7391 nw
tri 6841 7351 6881 7391 se
rect 6881 7351 7117 7391
rect 6621 6830 6773 7351
tri 6773 7323 6801 7351 nw
tri 6813 7323 6841 7351 se
rect 6841 7323 7117 7351
tri 6621 6806 6645 6830 ne
rect 6645 6806 6773 6830
tri 6565 6766 6605 6806 sw
tri 6645 6766 6685 6806 ne
rect 6685 6766 6773 6806
tri 6801 7311 6813 7323 se
rect 6813 7311 7117 7323
rect 6249 6734 6605 6766
tri 6605 6734 6637 6766 sw
rect 6801 6734 7117 7311
rect 6249 6570 6637 6734
tri 6637 6570 6801 6734 sw
tri 6801 6570 6965 6734 ne
rect 6965 6570 7117 6734
rect 6249 6568 6801 6570
tri 6801 6568 6803 6570 sw
tri 6965 6568 6967 6570 ne
rect 6249 6460 6803 6568
tri 6803 6460 6911 6568 sw
rect 6249 6372 6911 6460
tri 6249 6210 6411 6372 ne
tri 6193 6108 6202 6117 sw
rect 6141 6095 6202 6108
tri 6141 6086 6150 6095 ne
rect 5994 5947 6000 5999
rect 6052 5947 6064 5999
rect 6116 5947 6122 5999
rect 5994 5750 6046 5947
tri 6046 5922 6071 5947 nw
tri 6141 5893 6150 5902 se
rect 6150 5893 6202 6095
rect 6141 5880 6202 5893
rect 6141 5750 6193 5880
tri 6193 5871 6202 5880 nw
rect 6253 6107 6259 6159
rect 6311 6107 6323 6159
rect 6375 6107 6381 6159
rect 6253 5750 6305 6107
tri 6305 6031 6381 6107 nw
rect 6411 5750 6911 6372
rect 6967 5750 7117 6570
rect 7176 10575 7492 11017
rect 7176 5750 7306 10575
tri 7306 10389 7492 10575 nw
rect 5608 5574 5660 5750
tri 5660 5717 5693 5750 nw
rect 5608 5510 5660 5522
rect 5608 5452 5660 5458
rect 5528 4441 5580 4453
rect 5528 4193 5580 4389
tri 5580 4193 5608 4221 sw
rect 5528 4141 5534 4193
rect 5586 4141 5598 4193
rect 5650 4141 5656 4193
rect 3134 -588 3139 -536
rect 3191 -588 3203 -536
rect 3255 -588 3260 -536
rect 2837 -936 3026 -930
rect 2028 -1029 2040 -977
rect 2092 -1029 2104 -977
rect 2156 -1029 2168 -977
rect 1976 -1035 2220 -1029
rect 3134 -977 3260 -588
rect 3424 -814 3652 62
rect 3604 -930 3652 -814
rect 3424 -936 3652 -930
rect 3134 -1029 3139 -977
rect 3191 -1029 3203 -977
rect 3255 -1029 3260 -977
rect 3134 -1035 3260 -1029
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_0
timestamp 1707688321
transform 0 -1 680 -1 0 27571
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_1
timestamp 1707688321
transform 0 -1 680 -1 0 23676
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_2
timestamp 1707688321
transform 0 -1 680 -1 0 19781
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_3
timestamp 1707688321
transform 0 -1 680 -1 0 15886
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_4
timestamp 1707688321
transform 0 -1 680 -1 0 11991
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_5
timestamp 1707688321
transform 0 -1 680 -1 0 4201
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_6
timestamp 1707688321
transform 0 -1 680 -1 0 8096
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_7
timestamp 1707688321
transform 0 -1 806 -1 0 4201
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_8
timestamp 1707688321
transform 0 -1 806 -1 0 8096
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_9
timestamp 1707688321
transform 0 -1 806 -1 0 11991
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_10
timestamp 1707688321
transform 0 -1 806 -1 0 15886
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_11
timestamp 1707688321
transform 0 -1 806 -1 0 19781
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_12
timestamp 1707688321
transform 0 -1 806 -1 0 23676
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_13
timestamp 1707688321
transform 0 -1 806 -1 0 27571
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_14
timestamp 1707688321
transform 0 -1 932 -1 0 4201
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_15
timestamp 1707688321
transform 0 -1 932 -1 0 8096
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_16
timestamp 1707688321
transform 0 -1 932 -1 0 11991
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_17
timestamp 1707688321
transform 0 -1 932 -1 0 15886
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_18
timestamp 1707688321
transform 0 -1 932 -1 0 19781
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_19
timestamp 1707688321
transform 0 -1 932 -1 0 23676
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_20
timestamp 1707688321
transform 0 -1 932 -1 0 27571
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_21
timestamp 1707688321
transform 0 -1 1184 -1 0 4201
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_22
timestamp 1707688321
transform 0 -1 1184 -1 0 8096
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_23
timestamp 1707688321
transform 0 -1 1184 -1 0 11991
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_24
timestamp 1707688321
transform 0 -1 1184 -1 0 15886
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_25
timestamp 1707688321
transform 0 -1 1184 -1 0 19781
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_26
timestamp 1707688321
transform 0 -1 1184 -1 0 23676
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_27
timestamp 1707688321
transform 0 -1 1184 -1 0 27571
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_28
timestamp 1707688321
transform 0 -1 1058 -1 0 27571
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_29
timestamp 1707688321
transform 0 -1 1058 -1 0 23676
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_30
timestamp 1707688321
transform 0 -1 1058 -1 0 19781
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_31
timestamp 1707688321
transform 0 -1 1058 -1 0 15886
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_32
timestamp 1707688321
transform 0 -1 1058 -1 0 11991
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_33
timestamp 1707688321
transform 0 -1 1058 -1 0 8096
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_34
timestamp 1707688321
transform 0 -1 1058 -1 0 4201
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_35
timestamp 1707688321
transform 0 -1 1688 -1 0 4201
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_36
timestamp 1707688321
transform 0 -1 1688 -1 0 8096
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_37
timestamp 1707688321
transform 0 -1 1688 -1 0 23676
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_38
timestamp 1707688321
transform 0 -1 1688 -1 0 11991
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_39
timestamp 1707688321
transform 0 -1 1688 -1 0 15886
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_40
timestamp 1707688321
transform 0 -1 1688 -1 0 19781
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_41
timestamp 1707688321
transform 0 -1 1688 -1 0 27571
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_42
timestamp 1707688321
transform 0 -1 1562 -1 0 27571
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_43
timestamp 1707688321
transform 0 -1 1562 -1 0 23676
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_44
timestamp 1707688321
transform 0 -1 1562 -1 0 19781
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_45
timestamp 1707688321
transform 0 -1 1562 -1 0 15886
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_46
timestamp 1707688321
transform 0 -1 1562 -1 0 11991
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_47
timestamp 1707688321
transform 0 -1 1562 -1 0 8096
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_48
timestamp 1707688321
transform 0 -1 1562 -1 0 4201
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_49
timestamp 1707688321
transform 0 -1 1436 -1 0 27571
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_50
timestamp 1707688321
transform 0 -1 1436 -1 0 23676
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_51
timestamp 1707688321
transform 0 -1 1436 -1 0 19781
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_52
timestamp 1707688321
transform 0 -1 1436 -1 0 15886
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_53
timestamp 1707688321
transform 0 -1 1436 -1 0 11991
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_54
timestamp 1707688321
transform 0 -1 1436 -1 0 8096
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_55
timestamp 1707688321
transform 0 -1 1436 -1 0 4201
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_56
timestamp 1707688321
transform 0 -1 1310 -1 0 27571
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_57
timestamp 1707688321
transform 0 -1 1310 -1 0 23676
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_58
timestamp 1707688321
transform 0 -1 1310 -1 0 19781
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_59
timestamp 1707688321
transform 0 -1 1310 -1 0 15886
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_60
timestamp 1707688321
transform 0 -1 1310 -1 0 11991
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_61
timestamp 1707688321
transform 0 -1 1310 -1 0 8096
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_62
timestamp 1707688321
transform 0 -1 1310 -1 0 4201
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_63
timestamp 1707688321
transform 0 -1 2066 -1 0 5465
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_64
timestamp 1707688321
transform 0 -1 2066 -1 0 11991
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_65
timestamp 1707688321
transform 0 -1 2066 -1 0 15886
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_66
timestamp 1707688321
transform 0 -1 2066 -1 0 19781
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_67
timestamp 1707688321
transform 0 -1 2066 -1 0 23676
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_68
timestamp 1707688321
transform 0 -1 2066 -1 0 27571
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_69
timestamp 1707688321
transform 0 -1 1940 -1 0 27571
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_70
timestamp 1707688321
transform 0 -1 1940 -1 0 23676
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_71
timestamp 1707688321
transform 0 -1 1940 -1 0 19781
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_72
timestamp 1707688321
transform 0 -1 1940 -1 0 15886
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_73
timestamp 1707688321
transform 0 -1 1940 -1 0 11991
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_74
timestamp 1707688321
transform 0 -1 1940 -1 0 8096
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_75
timestamp 1707688321
transform 0 -1 1940 -1 0 4201
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_76
timestamp 1707688321
transform 0 -1 1814 -1 0 27571
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_77
timestamp 1707688321
transform 0 -1 1814 -1 0 23676
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_78
timestamp 1707688321
transform 0 -1 1814 -1 0 19781
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_79
timestamp 1707688321
transform 0 -1 1814 -1 0 15886
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_80
timestamp 1707688321
transform 0 -1 1814 -1 0 11991
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_81
timestamp 1707688321
transform 0 -1 1814 -1 0 8096
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_82
timestamp 1707688321
transform 0 -1 1814 -1 0 4201
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_83
timestamp 1707688321
transform 0 -1 428 -1 0 27571
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_84
timestamp 1707688321
transform 0 -1 428 -1 0 23676
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_85
timestamp 1707688321
transform 0 -1 428 -1 0 19781
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_86
timestamp 1707688321
transform 0 -1 428 -1 0 15886
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_87
timestamp 1707688321
transform 0 -1 428 -1 0 11991
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_88
timestamp 1707688321
transform 0 -1 554 -1 0 8096
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_89
timestamp 1707688321
transform 0 -1 554 -1 0 4201
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_90
timestamp 1707688321
transform 0 -1 554 -1 0 11991
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_91
timestamp 1707688321
transform 0 -1 554 -1 0 15886
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_92
timestamp 1707688321
transform 0 -1 554 -1 0 19781
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_93
timestamp 1707688321
transform 0 -1 554 -1 0 23676
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_94
timestamp 1707688321
transform 0 -1 554 -1 0 27571
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_95
timestamp 1707688321
transform 0 -1 428 -1 0 4201
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_96
timestamp 1707688321
transform 0 -1 428 -1 0 8096
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_97
timestamp 1707688321
transform 0 -1 2192 -1 0 5465
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_98
timestamp 1707688321
transform 0 -1 2318 -1 0 5465
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_99
timestamp 1707688321
transform 0 -1 2444 -1 0 5465
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_100
timestamp 1707688321
transform 0 -1 2570 -1 0 5465
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_101
timestamp 1707688321
transform 0 -1 2696 -1 0 5465
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_102
timestamp 1707688321
transform 0 -1 2822 -1 0 5465
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_103
timestamp 1707688321
transform 0 -1 2948 -1 0 5465
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_104
timestamp 1707688321
transform 0 -1 3074 -1 0 5465
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_105
timestamp 1707688321
transform 0 -1 680 1 0 23736
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_106
timestamp 1707688321
transform 0 -1 680 1 0 19841
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_107
timestamp 1707688321
transform 0 -1 680 1 0 15946
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_108
timestamp 1707688321
transform 0 -1 680 1 0 12051
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_109
timestamp 1707688321
transform 0 -1 680 1 0 8156
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_110
timestamp 1707688321
transform 0 -1 680 1 0 366
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_111
timestamp 1707688321
transform 0 -1 680 1 0 4261
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_112
timestamp 1707688321
transform 0 -1 806 1 0 366
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_113
timestamp 1707688321
transform 0 -1 806 1 0 4261
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_114
timestamp 1707688321
transform 0 -1 806 1 0 8156
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_115
timestamp 1707688321
transform 0 -1 806 1 0 12051
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_116
timestamp 1707688321
transform 0 -1 806 1 0 15946
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_117
timestamp 1707688321
transform 0 -1 806 1 0 19841
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_118
timestamp 1707688321
transform 0 -1 806 1 0 23736
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_119
timestamp 1707688321
transform 0 -1 932 1 0 366
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_120
timestamp 1707688321
transform 0 -1 932 1 0 4261
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_121
timestamp 1707688321
transform 0 -1 932 1 0 8156
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_122
timestamp 1707688321
transform 0 -1 932 1 0 12051
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_123
timestamp 1707688321
transform 0 -1 932 1 0 15946
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_124
timestamp 1707688321
transform 0 -1 932 1 0 19841
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_125
timestamp 1707688321
transform 0 -1 932 1 0 23736
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_126
timestamp 1707688321
transform 0 -1 1184 1 0 366
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_127
timestamp 1707688321
transform 0 -1 1184 1 0 4261
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_128
timestamp 1707688321
transform 0 -1 1184 1 0 8156
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_129
timestamp 1707688321
transform 0 -1 1184 1 0 12051
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_130
timestamp 1707688321
transform 0 -1 1184 1 0 15946
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_131
timestamp 1707688321
transform 0 -1 1184 1 0 19841
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_132
timestamp 1707688321
transform 0 -1 1184 1 0 23736
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_133
timestamp 1707688321
transform 0 -1 1058 1 0 23736
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_134
timestamp 1707688321
transform 0 -1 1058 1 0 19841
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_135
timestamp 1707688321
transform 0 -1 1058 1 0 15946
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_136
timestamp 1707688321
transform 0 -1 1058 1 0 12051
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_137
timestamp 1707688321
transform 0 -1 1058 1 0 8156
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_138
timestamp 1707688321
transform 0 -1 1058 1 0 4261
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_139
timestamp 1707688321
transform 0 -1 1058 1 0 366
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_140
timestamp 1707688321
transform 0 -1 1688 1 0 366
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_141
timestamp 1707688321
transform 0 -1 1688 1 0 4261
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_142
timestamp 1707688321
transform 0 -1 1688 1 0 22265
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_143
timestamp 1707688321
transform 0 -1 1688 1 0 8156
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_144
timestamp 1707688321
transform 0 -1 1688 1 0 12051
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_145
timestamp 1707688321
transform 0 -1 1688 1 0 15946
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_146
timestamp 1707688321
transform 0 -1 1688 1 0 23736
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_147
timestamp 1707688321
transform 0 -1 1562 1 0 23736
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_148
timestamp 1707688321
transform 0 -1 1562 1 0 19841
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_149
timestamp 1707688321
transform 0 -1 1562 1 0 15946
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_150
timestamp 1707688321
transform 0 -1 1562 1 0 12051
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_151
timestamp 1707688321
transform 0 -1 1562 1 0 8156
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_152
timestamp 1707688321
transform 0 -1 1562 1 0 4261
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_153
timestamp 1707688321
transform 0 -1 1562 1 0 366
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_154
timestamp 1707688321
transform 0 -1 1436 1 0 23736
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_155
timestamp 1707688321
transform 0 -1 1436 1 0 22265
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_156
timestamp 1707688321
transform 0 -1 1436 1 0 15946
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_157
timestamp 1707688321
transform 0 -1 1436 1 0 12051
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_158
timestamp 1707688321
transform 0 -1 1436 1 0 8156
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_159
timestamp 1707688321
transform 0 -1 1436 1 0 4261
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_160
timestamp 1707688321
transform 0 -1 1436 1 0 366
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_161
timestamp 1707688321
transform 0 -1 1310 1 0 23736
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_162
timestamp 1707688321
transform 0 -1 1310 1 0 19841
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_163
timestamp 1707688321
transform 0 -1 1310 1 0 15946
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_164
timestamp 1707688321
transform 0 -1 1310 1 0 12051
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_165
timestamp 1707688321
transform 0 -1 1310 1 0 8156
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_166
timestamp 1707688321
transform 0 -1 1310 1 0 4261
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_167
timestamp 1707688321
transform 0 -1 1310 1 0 366
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_168
timestamp 1707688321
transform 0 -1 2066 1 0 366
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_169
timestamp 1707688321
transform 0 -1 2066 1 0 8156
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_170
timestamp 1707688321
transform 0 -1 2066 1 0 12051
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_171
timestamp 1707688321
transform 0 -1 2066 1 0 15946
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_172
timestamp 1707688321
transform 0 -1 2066 1 0 19841
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_173
timestamp 1707688321
transform 0 -1 2066 1 0 23736
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_174
timestamp 1707688321
transform 0 -1 1940 1 0 23736
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_175
timestamp 1707688321
transform 0 -1 1940 1 0 15946
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_176
timestamp 1707688321
transform 0 -1 1940 1 0 12051
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_177
timestamp 1707688321
transform 0 -1 1940 1 0 8156
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_178
timestamp 1707688321
transform 0 -1 1940 1 0 4261
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_179
timestamp 1707688321
transform 0 -1 1940 1 0 366
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_180
timestamp 1707688321
transform 0 -1 1814 1 0 23736
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_181
timestamp 1707688321
transform 0 -1 1814 1 0 19841
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_182
timestamp 1707688321
transform 0 -1 1814 1 0 15946
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_183
timestamp 1707688321
transform 0 -1 1814 1 0 12051
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_184
timestamp 1707688321
transform 0 -1 1814 1 0 8156
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_185
timestamp 1707688321
transform 0 -1 1814 1 0 4261
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_186
timestamp 1707688321
transform 0 -1 1814 1 0 366
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_187
timestamp 1707688321
transform 0 -1 428 1 0 23736
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_188
timestamp 1707688321
transform 0 -1 428 1 0 19841
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_189
timestamp 1707688321
transform 0 -1 428 1 0 15946
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_190
timestamp 1707688321
transform 0 -1 428 1 0 12051
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_191
timestamp 1707688321
transform 0 -1 428 1 0 8156
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_192
timestamp 1707688321
transform 0 -1 554 1 0 4261
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_193
timestamp 1707688321
transform 0 -1 554 1 0 366
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_194
timestamp 1707688321
transform 0 -1 554 1 0 8156
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_195
timestamp 1707688321
transform 0 -1 554 1 0 12051
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_196
timestamp 1707688321
transform 0 -1 554 1 0 15946
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_197
timestamp 1707688321
transform 0 -1 554 1 0 19841
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_198
timestamp 1707688321
transform 0 -1 554 1 0 23736
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_199
timestamp 1707688321
transform 0 -1 428 1 0 366
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_200
timestamp 1707688321
transform 0 -1 428 1 0 4261
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_201
timestamp 1707688321
transform 0 -1 1940 1 0 22265
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_202
timestamp 1707688321
transform 0 -1 2192 1 0 366
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_203
timestamp 1707688321
transform 0 -1 2318 1 0 366
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_204
timestamp 1707688321
transform 0 -1 2444 1 0 366
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_205
timestamp 1707688321
transform 0 -1 2570 1 0 366
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_206
timestamp 1707688321
transform 0 -1 2696 1 0 366
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_207
timestamp 1707688321
transform 0 -1 2822 1 0 366
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_208
timestamp 1707688321
transform 0 -1 2948 1 0 366
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_209
timestamp 1707688321
transform 0 -1 3074 1 0 366
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1707688321
transform 0 -1 2494 -1 0 5654
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_1
timestamp 1707688321
transform -1 0 668 0 1 27445
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_2
timestamp 1707688321
transform -1 0 668 0 1 23550
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_3
timestamp 1707688321
transform -1 0 668 0 1 19655
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_4
timestamp 1707688321
transform -1 0 668 0 1 15760
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_5
timestamp 1707688321
transform -1 0 668 0 1 11865
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_6
timestamp 1707688321
transform -1 0 668 0 1 4001
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_7
timestamp 1707688321
transform -1 0 668 0 1 7970
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_8
timestamp 1707688321
transform -1 0 794 0 1 4001
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_9
timestamp 1707688321
transform -1 0 794 0 1 7970
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_10
timestamp 1707688321
transform -1 0 794 0 1 11865
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_11
timestamp 1707688321
transform -1 0 794 0 1 15760
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_12
timestamp 1707688321
transform -1 0 794 0 1 19655
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_13
timestamp 1707688321
transform -1 0 794 0 1 23550
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_14
timestamp 1707688321
transform -1 0 794 0 1 27445
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_15
timestamp 1707688321
transform -1 0 920 0 1 4001
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_16
timestamp 1707688321
transform -1 0 920 0 1 7970
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_17
timestamp 1707688321
transform -1 0 920 0 1 11865
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_18
timestamp 1707688321
transform -1 0 920 0 1 15760
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_19
timestamp 1707688321
transform -1 0 920 0 1 19655
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_20
timestamp 1707688321
transform -1 0 920 0 1 23550
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_21
timestamp 1707688321
transform -1 0 920 0 1 27445
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_22
timestamp 1707688321
transform -1 0 1172 0 1 4001
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_23
timestamp 1707688321
transform -1 0 1172 0 1 7970
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_24
timestamp 1707688321
transform -1 0 1172 0 1 11865
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_25
timestamp 1707688321
transform -1 0 1172 0 1 15760
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_26
timestamp 1707688321
transform -1 0 1172 0 1 19655
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_27
timestamp 1707688321
transform -1 0 1172 0 1 23550
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_28
timestamp 1707688321
transform -1 0 1172 0 1 27445
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_29
timestamp 1707688321
transform -1 0 1046 0 1 27445
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_30
timestamp 1707688321
transform -1 0 1046 0 1 23550
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_31
timestamp 1707688321
transform -1 0 1046 0 1 19655
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_32
timestamp 1707688321
transform -1 0 1046 0 1 15760
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_33
timestamp 1707688321
transform -1 0 1046 0 1 11865
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_34
timestamp 1707688321
transform -1 0 1046 0 1 7970
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_35
timestamp 1707688321
transform -1 0 1046 0 1 4001
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_36
timestamp 1707688321
transform -1 0 1676 0 1 4001
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_37
timestamp 1707688321
transform -1 0 1676 0 1 7970
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_38
timestamp 1707688321
transform -1 0 1676 0 1 23550
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_39
timestamp 1707688321
transform -1 0 1676 0 1 11865
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_40
timestamp 1707688321
transform -1 0 1676 0 1 15760
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_41
timestamp 1707688321
transform -1 0 1676 0 1 19655
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_42
timestamp 1707688321
transform -1 0 1676 0 1 27445
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_43
timestamp 1707688321
transform -1 0 1550 0 1 27445
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_44
timestamp 1707688321
transform -1 0 1550 0 1 23550
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_45
timestamp 1707688321
transform -1 0 1550 0 1 19655
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_46
timestamp 1707688321
transform -1 0 1550 0 1 15760
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_47
timestamp 1707688321
transform -1 0 1550 0 1 11865
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_48
timestamp 1707688321
transform -1 0 1550 0 1 7970
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_49
timestamp 1707688321
transform -1 0 1550 0 1 4001
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_50
timestamp 1707688321
transform -1 0 1424 0 1 27445
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_51
timestamp 1707688321
transform -1 0 1424 0 1 23550
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_52
timestamp 1707688321
transform -1 0 1424 0 1 19655
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_53
timestamp 1707688321
transform -1 0 1424 0 1 15760
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_54
timestamp 1707688321
transform -1 0 1424 0 1 11865
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_55
timestamp 1707688321
transform -1 0 1424 0 1 7970
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_56
timestamp 1707688321
transform -1 0 1424 0 1 4001
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_57
timestamp 1707688321
transform -1 0 1298 0 1 27445
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_58
timestamp 1707688321
transform -1 0 1298 0 1 23550
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_59
timestamp 1707688321
transform -1 0 1298 0 1 19655
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_60
timestamp 1707688321
transform -1 0 1298 0 1 15760
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_61
timestamp 1707688321
transform -1 0 1298 0 1 11865
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_62
timestamp 1707688321
transform -1 0 1298 0 1 7970
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_63
timestamp 1707688321
transform -1 0 1298 0 1 4001
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_64
timestamp 1707688321
transform -1 0 2054 0 1 5458
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_65
timestamp 1707688321
transform -1 0 2054 0 1 11865
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_66
timestamp 1707688321
transform -1 0 2054 0 1 15760
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_67
timestamp 1707688321
transform -1 0 2054 0 1 19655
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_68
timestamp 1707688321
transform -1 0 2054 0 1 23550
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_69
timestamp 1707688321
transform -1 0 2054 0 1 27445
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_70
timestamp 1707688321
transform -1 0 1928 0 1 27445
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_71
timestamp 1707688321
transform -1 0 1928 0 1 23550
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_72
timestamp 1707688321
transform -1 0 1928 0 1 19655
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_73
timestamp 1707688321
transform -1 0 1928 0 1 15760
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_74
timestamp 1707688321
transform -1 0 1928 0 1 11865
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_75
timestamp 1707688321
transform -1 0 1928 0 1 3966
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_76
timestamp 1707688321
transform -1 0 1802 0 1 27445
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_77
timestamp 1707688321
transform -1 0 1802 0 1 23550
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_78
timestamp 1707688321
transform -1 0 1802 0 1 19655
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_79
timestamp 1707688321
transform -1 0 1802 0 1 15760
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_80
timestamp 1707688321
transform -1 0 1802 0 1 11865
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_81
timestamp 1707688321
transform -1 0 1928 0 1 7882
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_82
timestamp 1707688321
transform -1 0 1802 0 1 4001
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_83
timestamp 1707688321
transform -1 0 416 0 1 7970
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_84
timestamp 1707688321
transform -1 0 416 0 1 4001
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_85
timestamp 1707688321
transform -1 0 416 0 1 11865
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_86
timestamp 1707688321
transform -1 0 416 0 1 15760
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_87
timestamp 1707688321
transform -1 0 416 0 1 19655
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_88
timestamp 1707688321
transform -1 0 416 0 1 23550
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_89
timestamp 1707688321
transform -1 0 416 0 1 27445
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_90
timestamp 1707688321
transform -1 0 542 0 1 7970
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_91
timestamp 1707688321
transform -1 0 542 0 1 4001
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_92
timestamp 1707688321
transform -1 0 542 0 1 11865
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_93
timestamp 1707688321
transform -1 0 542 0 1 15760
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_94
timestamp 1707688321
transform -1 0 542 0 1 19655
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_95
timestamp 1707688321
transform -1 0 542 0 1 23550
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_96
timestamp 1707688321
transform -1 0 542 0 1 27445
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_97
timestamp 1707688321
transform -1 0 2180 0 1 5164
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_98
timestamp 1707688321
transform -1 0 2306 0 1 5164
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_99
timestamp 1707688321
transform -1 0 2432 0 1 5164
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_100
timestamp 1707688321
transform -1 0 2558 0 1 5164
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_101
timestamp 1707688321
transform -1 0 2684 0 1 5164
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_102
timestamp 1707688321
transform -1 0 2810 0 1 5164
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_103
timestamp 1707688321
transform -1 0 2936 0 1 5164
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_104
timestamp 1707688321
transform -1 0 3062 0 1 5164
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_105
timestamp 1707688321
transform -1 0 3062 0 1 4001
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_106
timestamp 1707688321
transform -1 0 2054 0 1 4001
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_107
timestamp 1707688321
transform -1 0 2180 0 1 3966
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_108
timestamp 1707688321
transform -1 0 2306 0 1 4001
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_109
timestamp 1707688321
transform -1 0 2432 0 1 3966
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_110
timestamp 1707688321
transform -1 0 2558 0 1 4001
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_111
timestamp 1707688321
transform -1 0 2684 0 1 3966
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_112
timestamp 1707688321
transform -1 0 2810 0 1 4001
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_113
timestamp 1707688321
transform -1 0 2054 0 1 5164
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_114
timestamp 1707688321
transform -1 0 2936 0 1 3913
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_115
timestamp 1707688321
transform -1 0 1928 0 1 5164
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_116
timestamp 1707688321
transform -1 0 1928 0 1 5458
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_117
timestamp 1707688321
transform -1 0 668 0 -1 23862
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_118
timestamp 1707688321
transform -1 0 668 0 -1 19967
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_119
timestamp 1707688321
transform -1 0 668 0 -1 16072
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_120
timestamp 1707688321
transform -1 0 668 0 -1 12177
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_121
timestamp 1707688321
transform -1 0 668 0 -1 8282
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_122
timestamp 1707688321
transform -1 0 668 0 -1 492
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_123
timestamp 1707688321
transform -1 0 668 0 -1 4387
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_124
timestamp 1707688321
transform -1 0 794 0 -1 492
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_125
timestamp 1707688321
transform -1 0 794 0 -1 4387
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_126
timestamp 1707688321
transform -1 0 794 0 -1 8282
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_127
timestamp 1707688321
transform -1 0 794 0 -1 12177
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_128
timestamp 1707688321
transform -1 0 794 0 -1 16072
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_129
timestamp 1707688321
transform -1 0 794 0 -1 19967
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_130
timestamp 1707688321
transform -1 0 794 0 -1 23862
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_131
timestamp 1707688321
transform -1 0 920 0 -1 492
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_132
timestamp 1707688321
transform -1 0 920 0 -1 4387
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_133
timestamp 1707688321
transform -1 0 920 0 -1 8282
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_134
timestamp 1707688321
transform -1 0 920 0 -1 12177
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_135
timestamp 1707688321
transform -1 0 920 0 -1 16072
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_136
timestamp 1707688321
transform -1 0 920 0 -1 19967
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_137
timestamp 1707688321
transform -1 0 920 0 -1 23862
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_138
timestamp 1707688321
transform -1 0 1172 0 -1 492
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_139
timestamp 1707688321
transform -1 0 1172 0 -1 4387
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_140
timestamp 1707688321
transform -1 0 1172 0 -1 8282
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_141
timestamp 1707688321
transform -1 0 1172 0 -1 12177
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_142
timestamp 1707688321
transform -1 0 1172 0 -1 16072
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_143
timestamp 1707688321
transform -1 0 1172 0 -1 19967
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_144
timestamp 1707688321
transform -1 0 1172 0 -1 23862
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_145
timestamp 1707688321
transform -1 0 1046 0 -1 23862
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_146
timestamp 1707688321
transform -1 0 1046 0 -1 19967
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_147
timestamp 1707688321
transform -1 0 1046 0 -1 16072
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_148
timestamp 1707688321
transform -1 0 1046 0 -1 12177
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_149
timestamp 1707688321
transform -1 0 1046 0 -1 8282
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_150
timestamp 1707688321
transform -1 0 1046 0 -1 4387
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_151
timestamp 1707688321
transform -1 0 1046 0 -1 492
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_152
timestamp 1707688321
transform -1 0 1676 0 -1 492
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_153
timestamp 1707688321
transform -1 0 1676 0 -1 8282
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_154
timestamp 1707688321
transform -1 0 1676 0 -1 12177
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_155
timestamp 1707688321
transform -1 0 1676 0 -1 16072
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_156
timestamp 1707688321
transform -1 0 1676 0 -1 22391
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_157
timestamp 1707688321
transform -1 0 1676 0 -1 23862
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_158
timestamp 1707688321
transform -1 0 1550 0 -1 23862
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_159
timestamp 1707688321
transform -1 0 1550 0 -1 19967
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_160
timestamp 1707688321
transform -1 0 1550 0 -1 16072
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_161
timestamp 1707688321
transform -1 0 1550 0 -1 12177
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_162
timestamp 1707688321
transform -1 0 1550 0 -1 8282
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_163
timestamp 1707688321
transform -1 0 1550 0 -1 4407
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_164
timestamp 1707688321
transform -1 0 1550 0 -1 492
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_165
timestamp 1707688321
transform -1 0 1424 0 -1 23862
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_166
timestamp 1707688321
transform -1 0 1424 0 -1 22391
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_167
timestamp 1707688321
transform -1 0 1424 0 -1 16072
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_168
timestamp 1707688321
transform -1 0 1424 0 -1 12177
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_169
timestamp 1707688321
transform -1 0 1424 0 -1 8282
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_170
timestamp 1707688321
transform -1 0 1424 0 -1 492
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_171
timestamp 1707688321
transform -1 0 1298 0 -1 23862
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_172
timestamp 1707688321
transform -1 0 1298 0 -1 19967
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_173
timestamp 1707688321
transform -1 0 1298 0 -1 16072
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_174
timestamp 1707688321
transform -1 0 1298 0 -1 12177
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_175
timestamp 1707688321
transform -1 0 1298 0 -1 8282
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_176
timestamp 1707688321
transform -1 0 1298 0 -1 4644
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_177
timestamp 1707688321
transform -1 0 1298 0 -1 492
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_178
timestamp 1707688321
transform -1 0 2054 0 -1 12177
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_179
timestamp 1707688321
transform -1 0 2054 0 -1 16072
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_180
timestamp 1707688321
transform -1 0 2054 0 -1 19967
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_181
timestamp 1707688321
transform -1 0 2054 0 -1 23862
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_182
timestamp 1707688321
transform -1 0 1928 0 -1 23862
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_183
timestamp 1707688321
transform -1 0 1928 0 -1 16072
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_184
timestamp 1707688321
transform -1 0 1928 0 -1 12177
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_185
timestamp 1707688321
transform -1 0 1928 0 -1 8282
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_186
timestamp 1707688321
transform -1 0 1928 0 -1 4407
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_187
timestamp 1707688321
transform -1 0 1928 0 -1 492
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_188
timestamp 1707688321
transform -1 0 1802 0 -1 23862
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_189
timestamp 1707688321
transform -1 0 1802 0 -1 19967
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_190
timestamp 1707688321
transform -1 0 1802 0 -1 16072
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_191
timestamp 1707688321
transform -1 0 1802 0 -1 12177
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_192
timestamp 1707688321
transform -1 0 1802 0 -1 8282
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_193
timestamp 1707688321
transform -1 0 1802 0 -1 4407
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_194
timestamp 1707688321
transform -1 0 1802 0 -1 492
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_195
timestamp 1707688321
transform -1 0 416 0 -1 4387
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_196
timestamp 1707688321
transform -1 0 416 0 -1 492
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_197
timestamp 1707688321
transform -1 0 416 0 -1 8282
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_198
timestamp 1707688321
transform -1 0 416 0 -1 12177
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_199
timestamp 1707688321
transform -1 0 416 0 -1 16072
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_200
timestamp 1707688321
transform -1 0 416 0 -1 19967
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_201
timestamp 1707688321
transform -1 0 416 0 -1 23862
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_202
timestamp 1707688321
transform -1 0 542 0 -1 4387
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_203
timestamp 1707688321
transform -1 0 542 0 -1 492
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_204
timestamp 1707688321
transform -1 0 542 0 -1 8282
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_205
timestamp 1707688321
transform -1 0 542 0 -1 12177
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_206
timestamp 1707688321
transform -1 0 542 0 -1 16072
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_207
timestamp 1707688321
transform -1 0 542 0 -1 19967
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_208
timestamp 1707688321
transform -1 0 542 0 -1 23862
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_209
timestamp 1707688321
transform -1 0 1928 0 -1 22391
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_210
timestamp 1707688321
transform -1 0 2180 0 -1 572
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_211
timestamp 1707688321
transform -1 0 2306 0 -1 572
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_212
timestamp 1707688321
transform -1 0 2432 0 -1 572
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_213
timestamp 1707688321
transform -1 0 2558 0 -1 492
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_214
timestamp 1707688321
transform -1 0 2684 0 -1 492
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_215
timestamp 1707688321
transform -1 0 2810 0 -1 492
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_216
timestamp 1707688321
transform -1 0 2936 0 -1 492
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_217
timestamp 1707688321
transform -1 0 3062 0 -1 492
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_218
timestamp 1707688321
transform -1 0 3062 0 -1 4407
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_219
timestamp 1707688321
transform -1 0 2936 0 -1 4407
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_220
timestamp 1707688321
transform -1 0 2054 0 -1 572
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_221
timestamp 1707688321
transform -1 0 2054 0 -1 4407
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_222
timestamp 1707688321
transform -1 0 2180 0 -1 4407
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_223
timestamp 1707688321
transform -1 0 2306 0 -1 4407
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_224
timestamp 1707688321
transform -1 0 2432 0 -1 4407
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_225
timestamp 1707688321
transform -1 0 2558 0 -1 4407
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_226
timestamp 1707688321
transform -1 0 2684 0 -1 4407
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_227
timestamp 1707688321
transform -1 0 2810 0 -1 4407
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_228
timestamp 1707688321
transform -1 0 1424 0 -1 4407
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_229
timestamp 1707688321
transform -1 0 1676 0 -1 4407
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1707688321
transform 0 -1 2948 -1 0 -44
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1707688321
transform 0 1 2334 -1 0 6264
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1707688321
transform -1 0 2391 0 1 -673
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1707688321
transform -1 0 2103 0 -1 -280
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1707688321
transform -1 0 2443 0 -1 -280
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1707688321
transform -1 0 3081 0 -1 -639
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1707688321
transform 0 1 2266 1 0 -825
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1707688321
transform 0 1 2698 1 0 -825
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1707688321
transform 0 -1 3164 1 0 -825
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_9
timestamp 1707688321
transform 0 -1 2516 1 0 -924
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_10
timestamp 1707688321
transform 0 -1 2948 1 0 -924
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_11
timestamp 1707688321
transform 0 -1 3380 1 0 -924
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_12
timestamp 1707688321
transform 1 0 172 0 -1 27869
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_13
timestamp 1707688321
transform 1 0 5465 0 1 5959
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_14
timestamp 1707688321
transform 1 0 2230 0 1 5540
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_15
timestamp 1707688321
transform 1 0 2455 0 1 -673
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1707688321
transform 0 -1 2492 1 0 -234
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1707688321
transform 0 -1 3404 1 0 -234
box 0 0 1 1
use L1M1_CDNS_52468879185191  L1M1_CDNS_52468879185191_0
timestamp 1707688321
transform 0 -1 3682 -1 0 5248
box -12 -6 838 40
use L1M1_CDNS_52468879185191  L1M1_CDNS_52468879185191_1
timestamp 1707688321
transform 0 -1 3994 -1 0 5248
box -12 -6 838 40
use L1M1_CDNS_52468879185191  L1M1_CDNS_52468879185191_2
timestamp 1707688321
transform 0 -1 4306 -1 0 5248
box -12 -6 838 40
use L1M1_CDNS_52468879185191  L1M1_CDNS_52468879185191_3
timestamp 1707688321
transform 0 -1 4618 -1 0 5248
box -12 -6 838 40
use L1M1_CDNS_52468879185191  L1M1_CDNS_52468879185191_4
timestamp 1707688321
transform 0 -1 5282 -1 0 5248
box -12 -6 838 40
use L1M1_CDNS_52468879185193  L1M1_CDNS_52468879185193_0
timestamp 1707688321
transform -1 0 2869 0 1 -240
box 0 0 1 1
use L1M1_CDNS_52468879185194  L1M1_CDNS_52468879185194_0
timestamp 1707688321
transform 0 -1 4930 1 0 4422
box -12 -6 766 40
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_0
timestamp 1707688321
transform -1 0 5212 0 1 5458
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_1
timestamp 1707688321
transform 1 0 1673 0 -1 27869
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_2
timestamp 1707688321
transform 1 0 2998 0 1 -314
box 0 0 1 1
use L1M1_CDNS_52468879185307  L1M1_CDNS_52468879185307_0
timestamp 1707688321
transform -1 0 6494 0 1 10723
box -12 -6 1414 40
use L1M1_CDNS_52468879185307  L1M1_CDNS_52468879185307_1
timestamp 1707688321
transform 1 0 2948 0 1 10723
box -12 -6 1414 40
use L1M1_CDNS_52468879185316  L1M1_CDNS_52468879185316_0
timestamp 1707688321
transform -1 0 3122 0 1 5540
box -12 -6 622 40
use L1M1_CDNS_52468879185316  L1M1_CDNS_52468879185316_1
timestamp 1707688321
transform 0 -1 4774 1 0 4656
box -12 -6 622 40
use L1M1_CDNS_52468879185316  L1M1_CDNS_52468879185316_2
timestamp 1707688321
transform 0 -1 5106 1 0 4654
box -12 -6 622 40
use L1M1_CDNS_52468879185326  L1M1_CDNS_52468879185326_0
timestamp 1707688321
transform 0 -1 3838 1 0 4656
box -12 -6 694 40
use L1M1_CDNS_52468879185326  L1M1_CDNS_52468879185326_1
timestamp 1707688321
transform 0 -1 4150 1 0 4656
box -12 -6 694 40
use L1M1_CDNS_52468879185326  L1M1_CDNS_52468879185326_2
timestamp 1707688321
transform 0 -1 4462 1 0 4656
box -12 -6 694 40
use L1M1_CDNS_52468879185335  L1M1_CDNS_52468879185335_0
timestamp 1707688321
transform -1 0 4854 0 1 5458
box -12 -6 1126 40
use L1M1_CDNS_52468879185381  L1M1_CDNS_52468879185381_0
timestamp 1707688321
transform 0 -1 5655 -1 0 5248
box -12 -6 910 40
use L1M1_CDNS_52468879185381  L1M1_CDNS_52468879185381_1
timestamp 1707688321
transform 0 -1 3565 -1 0 5248
box -12 -6 910 40
use L1M1_CDNS_52468879185381  L1M1_CDNS_52468879185381_2
timestamp 1707688321
transform 0 -1 3187 -1 0 5248
box -12 -6 910 40
use L1M1_CDNS_52468879185381  L1M1_CDNS_52468879185381_3
timestamp 1707688321
transform 1 0 814 0 -1 -629
box -12 -6 910 40
use L1M1_CDNS_52468879185448  L1M1_CDNS_52468879185448_0
timestamp 1707688321
transform -1 0 4350 0 -1 6591
box -12 -6 1270 40
use L1M1_CDNS_52468879185448  L1M1_CDNS_52468879185448_1
timestamp 1707688321
transform 1 0 5092 0 -1 6591
box -12 -6 1270 40
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_0
timestamp 1707688321
transform 0 -1 3187 1 0 5464
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_1
timestamp 1707688321
transform 0 -1 3565 1 0 5464
box 0 0 1 1
use L1M1_CDNS_52468879185939  L1M1_CDNS_52468879185939_0
timestamp 1707688321
transform 0 -1 291 -1 0 27594
box -12 -6 20710 40
use L1M1_CDNS_52468879185940  L1M1_CDNS_52468879185940_0
timestamp 1707688321
transform 1 0 338 0 -1 176
box -12 -6 2782 40
use L1M1_CDNS_52468879185941  L1M1_CDNS_52468879185941_0
timestamp 1707688321
transform 1 0 3604 0 -1 4335
box -12 -6 1990 40
use L1M1_CDNS_52468879185942  L1M1_CDNS_52468879185942_0
timestamp 1707688321
transform 0 1 2743 1 0 6480
box -12 -6 4366 40
use L1M1_CDNS_52468879185943  L1M1_CDNS_52468879185943_0
timestamp 1707688321
transform 0 1 6665 -1 0 10834
box -12 -6 4222 40
use L1M1_CDNS_52468879185944  L1M1_CDNS_52468879185944_0
timestamp 1707688321
transform 0 1 3153 1 0 318
box -12 -6 3790 40
use L1M1_CDNS_52468879185944  L1M1_CDNS_52468879185944_1
timestamp 1707688321
transform 0 1 257 1 0 318
box -12 -6 3790 40
use L1M1_CDNS_52468879185944  L1M1_CDNS_52468879185944_2
timestamp 1707688321
transform 1 0 2832 0 -1 10889
box -12 -6 3790 40
use L1M1_CDNS_52468879185945  L1M1_CDNS_52468879185945_0
timestamp 1707688321
transform 0 -1 5726 -1 0 8582
box -12 -6 1846 40
use L1M1_CDNS_52468879185945  L1M1_CDNS_52468879185945_1
timestamp 1707688321
transform 0 -1 6582 -1 0 8582
box -12 -6 1846 40
use L1M1_CDNS_52468879185945  L1M1_CDNS_52468879185945_2
timestamp 1707688321
transform 0 -1 4870 -1 0 8582
box -12 -6 1846 40
use L1M1_CDNS_52468879185945  L1M1_CDNS_52468879185945_3
timestamp 1707688321
transform 0 1 4572 -1 0 8582
box -12 -6 1846 40
use L1M1_CDNS_52468879185945  L1M1_CDNS_52468879185945_4
timestamp 1707688321
transform 0 1 3716 -1 0 8582
box -12 -6 1846 40
use L1M1_CDNS_52468879185945  L1M1_CDNS_52468879185945_5
timestamp 1707688321
transform 0 1 2860 -1 0 8582
box -12 -6 1846 40
use L1M1_CDNS_52468879185945  L1M1_CDNS_52468879185945_6
timestamp 1707688321
transform 0 1 4572 1 0 8732
box -12 -6 1846 40
use L1M1_CDNS_52468879185945  L1M1_CDNS_52468879185945_7
timestamp 1707688321
transform 0 1 2860 1 0 8732
box -12 -6 1846 40
use L1M1_CDNS_52468879185945  L1M1_CDNS_52468879185945_8
timestamp 1707688321
transform 0 1 3716 1 0 8732
box -12 -6 1846 40
use L1M1_CDNS_52468879185945  L1M1_CDNS_52468879185945_9
timestamp 1707688321
transform 0 -1 6582 1 0 8732
box -12 -6 1846 40
use L1M1_CDNS_52468879185945  L1M1_CDNS_52468879185945_10
timestamp 1707688321
transform 0 -1 5726 1 0 8732
box -12 -6 1846 40
use L1M1_CDNS_52468879185945  L1M1_CDNS_52468879185945_11
timestamp 1707688321
transform 0 -1 4870 1 0 8732
box -12 -6 1846 40
use L1M1_CDNS_52468879185945  L1M1_CDNS_52468879185945_12
timestamp 1707688321
transform 1 0 3573 0 1 5540
box -12 -6 1846 40
use L1M1_CDNS_52468879185946  L1M1_CDNS_52468879185946_0
timestamp 1707688321
transform 0 1 4704 1 0 6612
box -12 -6 4150 40
use L1M1_CDNS_52468879185947  L1M1_CDNS_52468879185947_0
timestamp 1707688321
transform 0 1 2145 1 0 5584
box -12 -6 2566 40
use L1M1_CDNS_52468879185948  L1M1_CDNS_52468879185948_0
timestamp 1707688321
transform 1 0 337 0 -1 27707
box -12 -6 1702 40
use L1M1_CDNS_52468879185949  L1M1_CDNS_52468879185949_0
timestamp 1707688321
transform 0 1 2145 1 0 8396
box -12 -6 19126 40
use L1M1_CDNS_52468879185950  L1M1_CDNS_52468879185950_0
timestamp 1707688321
transform 0 1 2334 -1 0 22730
box -12 -6 11638 40
use L1M1_CDNS_52468879185951  L1M1_CDNS_52468879185951_0
timestamp 1707688321
transform 0 1 2334 -1 0 10877
box -12 -6 4438 40
use L1M1_CDNS_52468879185951  L1M1_CDNS_52468879185951_1
timestamp 1707688321
transform 0 1 2554 1 0 6451
box -12 -6 4438 40
use L1M1_CDNS_52468879185952  L1M1_CDNS_52468879185952_0
timestamp 1707688321
transform 0 -1 6888 1 0 6696
box -12 -6 3934 40
use L1M1_CDNS_52468879185953  L1M1_CDNS_52468879185953_0
timestamp 1707688321
transform -1 0 5341 0 -1 6459
box -12 -6 2278 40
use L1M1_CDNS_52468879185954  L1M1_CDNS_52468879185954_0
timestamp 1707688321
transform 1 0 2616 0 -1 6270
box -12 -6 2854 40
use L1M1_CDNS_52468879185955  L1M1_CDNS_52468879185955_0
timestamp 1707688321
transform 1 0 5386 0 -1 6459
box -12 -6 982 40
use L1M1_CDNS_52468879185956  L1M1_CDNS_52468879185956_0
timestamp 1707688321
transform -1 0 3299 0 -1 102
box -12 -6 2494 40
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1707688321
transform 0 -1 5580 -1 0 4511
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1707688321
transform 0 -1 5660 -1 0 5580
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1707688321
transform 0 1 373 -1 0 499
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1707688321
transform 0 1 2325 -1 0 6235
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1707688321
transform 0 1 2260 -1 0 -707
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_5
timestamp 1707688321
transform 0 1 499 -1 0 499
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_6
timestamp 1707688321
transform -1 0 5656 0 1 4141
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_7
timestamp 1707688321
transform -1 0 5722 0 1 6321
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_8
timestamp 1707688321
transform -1 0 3368 0 1 5682
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_9
timestamp 1707688321
transform -1 0 2635 0 1 6107
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_10
timestamp 1707688321
transform -1 0 5128 0 1 5867
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_11
timestamp 1707688321
transform -1 0 5449 0 1 6027
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_12
timestamp 1707688321
transform -1 0 6381 0 1 6107
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_13
timestamp 1707688321
transform -1 0 6122 0 1 5947
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_14
timestamp 1707688321
transform -1 0 2729 0 1 -679
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_15
timestamp 1707688321
transform -1 0 2573 0 1 -679
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_16
timestamp 1707688321
transform -1 0 2388 0 -1 -194
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_17
timestamp 1707688321
transform -1 0 2818 0 -1 -707
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_18
timestamp 1707688321
transform 0 1 2045 1 0 8206
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_19
timestamp 1707688321
transform 0 1 4996 1 0 5947
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_20
timestamp 1707688321
transform 0 1 1965 1 0 8022
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_21
timestamp 1707688321
transform 0 1 3054 1 0 -835
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_22
timestamp 1707688321
transform 0 -1 2948 1 0 4065
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_23
timestamp 1707688321
transform 0 -1 3106 1 0 -246
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_24
timestamp 1707688321
transform 1 0 5608 0 -1 5845
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_25
timestamp 1707688321
transform 1 0 1338 0 -1 27637
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_26
timestamp 1707688321
transform 1 0 2690 0 1 -326
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_0
timestamp 1707688321
transform 0 1 3642 1 0 4410
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_1
timestamp 1707688321
transform 0 -1 5288 1 0 4410
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_0
timestamp 1707688321
transform 0 1 3144 -1 0 5580
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_1
timestamp 1707688321
transform -1 0 4968 0 1 6526
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_2
timestamp 1707688321
transform -1 0 4968 0 -1 10788
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_3
timestamp 1707688321
transform 1 0 4468 0 -1 10788
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_4
timestamp 1707688321
transform 1 0 4468 0 1 6526
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_5
timestamp 1707688321
transform 1 0 1338 0 1 27667
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_6
timestamp 1707688321
transform 1 0 534 0 1 27667
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_7
timestamp 1707688321
transform 1 0 1338 0 1 136
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_0
timestamp 1707688321
transform 0 1 3424 -1 0 -808
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_1
timestamp 1707688321
transform 0 1 2837 -1 0 -808
box 0 0 1 1
use M1M2_CDNS_52468879185201  M1M2_CDNS_52468879185201_0
timestamp 1707688321
transform 1 0 2125 0 1 -16
box 0 0 320 116
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_0
timestamp 1707688321
transform -1 0 1877 0 1 27746
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_1
timestamp 1707688321
transform 0 1 499 1 0 -329
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_2
timestamp 1707688321
transform 1 0 729 0 -1 262
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_3
timestamp 1707688321
transform 1 0 132 0 -1 27878
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_4
timestamp 1707688321
transform 1 0 1005 0 -1 262
box 0 0 1 1
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_0
timestamp 1707688321
transform 1 0 1010 0 -1 27637
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_0
timestamp 1707688321
transform -1 0 3087 0 1 5797
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_1
timestamp 1707688321
transform -1 0 2964 0 1 6432
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_2
timestamp 1707688321
transform -1 0 3078 0 1 380
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_3
timestamp 1707688321
transform -1 0 2552 0 -1 5999
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_4
timestamp 1707688321
transform 0 -1 3255 1 0 -1035
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_5
timestamp 1707688321
transform 0 -1 3255 1 0 -594
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_6
timestamp 1707688321
transform 0 -1 3259 1 0 6401
box 0 0 1 1
use M1M2_CDNS_52468879185957  M1M2_CDNS_52468879185957_0
timestamp 1707688321
transform 0 -1 300 -1 0 27465
box 0 0 20608 52
use M1M2_CDNS_52468879185958  M1M2_CDNS_52468879185958_0
timestamp 1707688321
transform 0 1 3973 1 0 4410
box 0 0 192 436
use M1M2_CDNS_52468879185959  M1M2_CDNS_52468879185959_0
timestamp 1707688321
transform 0 1 5109 1 0 10849
box 0 0 1 1
use M1M2_CDNS_52468879185959  M1M2_CDNS_52468879185959_1
timestamp 1707688321
transform 0 1 3429 1 0 10849
box 0 0 1 1
use M1M2_CDNS_52468879185960  M1M2_CDNS_52468879185960_0
timestamp 1707688321
transform 0 1 3973 1 0 10849
box 0 0 1 1
use M1M2_CDNS_52468879185960  M1M2_CDNS_52468879185960_1
timestamp 1707688321
transform 0 1 3973 1 0 6401
box 0 0 1 1
use M1M2_CDNS_52468879185960  M1M2_CDNS_52468879185960_2
timestamp 1707688321
transform 0 1 5637 1 0 10849
box 0 0 1 1
use M1M2_CDNS_52468879185960  M1M2_CDNS_52468879185960_3
timestamp 1707688321
transform 0 1 6269 1 0 10849
box 0 0 1 1
use M1M2_CDNS_52468879185961  M1M2_CDNS_52468879185961_0
timestamp 1707688321
transform 0 1 5109 1 0 6401
box 0 0 1 1
use M1M2_CDNS_52468879185961  M1M2_CDNS_52468879185961_1
timestamp 1707688321
transform 0 1 3424 1 0 6401
box 0 0 1 1
use M1M2_CDNS_52468879185961  M1M2_CDNS_52468879185961_2
timestamp 1707688321
transform 0 1 3015 1 0 10849
box 0 0 1 1
use M1M2_CDNS_52468879185961  M1M2_CDNS_52468879185961_3
timestamp 1707688321
transform 0 -1 2220 1 0 -1035
box 0 0 1 1
use M1M2_CDNS_52468879185961  M1M2_CDNS_52468879185961_4
timestamp 1707688321
transform 0 -1 2220 1 0 -594
box 0 0 1 1
use M1M2_CDNS_52468879185962  M1M2_CDNS_52468879185962_0
timestamp 1707688321
transform 0 1 1965 -1 0 27377
box 0 0 3456 52
use M1M2_CDNS_52468879185962  M1M2_CDNS_52468879185962_1
timestamp 1707688321
transform 0 1 1965 -1 0 19608
box 0 0 3456 52
use M1M2_CDNS_52468879185962  M1M2_CDNS_52468879185962_2
timestamp 1707688321
transform 0 1 1965 1 0 12224
box 0 0 3456 52
use M1M2_CDNS_52468879185963  M1M2_CDNS_52468879185963_0
timestamp 1707688321
transform 0 1 3144 -1 0 5255
box 0 0 960 116
use M1M2_CDNS_52468879185964  M1M2_CDNS_52468879185964_0
timestamp 1707688321
transform 0 1 3144 1 0 136
box 0 0 3968 116
use M1M2_CDNS_52468879185964  M1M2_CDNS_52468879185964_1
timestamp 1707688321
transform 0 -1 7083 1 0 6662
box 0 0 3968 116
use M1M2_CDNS_52468879185965  M1M2_CDNS_52468879185965_0
timestamp 1707688321
transform 0 1 1965 1 0 20047
box 0 0 2176 52
use M1M2_CDNS_52468879185966  M1M2_CDNS_52468879185966_0
timestamp 1707688321
transform 0 1 1965 1 0 22479
box 0 0 1024 52
use M1M2_CDNS_52468879185967  M1M2_CDNS_52468879185967_0
timestamp 1707688321
transform 1 0 1601 0 1 136
box 0 0 448 116
use M1M2_CDNS_52468879185968  M1M2_CDNS_52468879185968_0
timestamp 1707688321
transform 0 1 2325 1 0 6409
box 0 0 4480 52
use M1M2_CDNS_52468879185969  M1M2_CDNS_52468879185969_0
timestamp 1707688321
transform 0 1 1965 1 0 8362
box 0 0 2048 52
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_0
timestamp 1707688321
transform 0 1 2029 1 0 8022
box 0 0 1 1
use M1M2_CDNS_52468879185971  M1M2_CDNS_52468879185971_0
timestamp 1707688321
transform 0 -1 300 1 0 268
box 0 0 3200 52
use M1M2_CDNS_52468879185972  M1M2_CDNS_52468879185972_0
timestamp 1707688321
transform 0 -1 6085 1 0 6401
box 0 0 1 1
use M1M2_CDNS_52468879185973  M1M2_CDNS_52468879185973_0
timestamp 1707688321
transform 0 1 2734 -1 0 10885
box 0 0 4288 52
use M1M2_CDNS_52468879185974  M1M2_CDNS_52468879185974_0
timestamp 1707688321
transform 0 -1 6737 -1 0 10798
box 0 0 4032 52
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_0
timestamp 1707688321
transform 0 1 229 1 0 -84
box 0 0 192 180
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_0
timestamp 1707688321
transform 0 -1 684 -1 0 27461
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_1
timestamp 1707688321
transform 0 -1 684 -1 0 23566
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_2
timestamp 1707688321
transform 0 -1 684 -1 0 19671
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_3
timestamp 1707688321
transform 0 -1 684 -1 0 15776
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_4
timestamp 1707688321
transform 0 -1 684 -1 0 11881
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_5
timestamp 1707688321
transform 0 -1 684 -1 0 7986
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_6
timestamp 1707688321
transform 0 -1 684 -1 0 4091
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_7
timestamp 1707688321
transform 0 -1 810 -1 0 7986
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_8
timestamp 1707688321
transform 0 -1 810 -1 0 4091
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_9
timestamp 1707688321
transform 0 -1 810 -1 0 11881
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_10
timestamp 1707688321
transform 0 -1 810 -1 0 15776
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_11
timestamp 1707688321
transform 0 -1 810 -1 0 19671
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_12
timestamp 1707688321
transform 0 -1 810 -1 0 23566
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_13
timestamp 1707688321
transform 0 -1 810 -1 0 27461
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_14
timestamp 1707688321
transform 0 -1 936 -1 0 7986
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_15
timestamp 1707688321
transform 0 -1 936 -1 0 4091
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_16
timestamp 1707688321
transform 0 -1 936 -1 0 11881
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_17
timestamp 1707688321
transform 0 -1 936 -1 0 15776
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_18
timestamp 1707688321
transform 0 -1 936 -1 0 19671
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_19
timestamp 1707688321
transform 0 -1 936 -1 0 23566
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_20
timestamp 1707688321
transform 0 -1 936 -1 0 27461
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_21
timestamp 1707688321
transform 0 -1 1188 -1 0 7986
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_22
timestamp 1707688321
transform 0 -1 1188 -1 0 4091
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_23
timestamp 1707688321
transform 0 -1 1188 -1 0 11881
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_24
timestamp 1707688321
transform 0 -1 1188 -1 0 15776
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_25
timestamp 1707688321
transform 0 -1 1188 -1 0 19671
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_26
timestamp 1707688321
transform 0 -1 1188 -1 0 23566
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_27
timestamp 1707688321
transform 0 -1 1188 -1 0 27461
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_28
timestamp 1707688321
transform 0 -1 1062 -1 0 27461
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_29
timestamp 1707688321
transform 0 -1 1062 -1 0 23566
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_30
timestamp 1707688321
transform 0 -1 1062 -1 0 19671
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_31
timestamp 1707688321
transform 0 -1 1062 -1 0 15776
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_32
timestamp 1707688321
transform 0 -1 1062 -1 0 11881
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_33
timestamp 1707688321
transform 0 -1 1062 -1 0 4091
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_34
timestamp 1707688321
transform 0 -1 1062 -1 0 7986
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_35
timestamp 1707688321
transform 0 -1 1692 -1 0 7986
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_36
timestamp 1707688321
transform 0 -1 1692 -1 0 4091
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_37
timestamp 1707688321
transform 0 -1 1692 -1 0 11881
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_38
timestamp 1707688321
transform 0 -1 1692 -1 0 15776
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_39
timestamp 1707688321
transform 0 -1 1692 -1 0 19671
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_40
timestamp 1707688321
transform 0 -1 1692 -1 0 27461
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_41
timestamp 1707688321
transform 0 -1 1566 -1 0 27461
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_42
timestamp 1707688321
transform 0 -1 1566 -1 0 23566
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_43
timestamp 1707688321
transform 0 -1 1566 -1 0 19671
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_44
timestamp 1707688321
transform 0 -1 1566 -1 0 15776
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_45
timestamp 1707688321
transform 0 -1 1566 -1 0 11881
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_46
timestamp 1707688321
transform 0 -1 1566 -1 0 4091
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_47
timestamp 1707688321
transform 0 -1 1566 -1 0 7986
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_48
timestamp 1707688321
transform 0 -1 1440 -1 0 27461
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_49
timestamp 1707688321
transform 0 -1 1440 -1 0 19671
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_50
timestamp 1707688321
transform 0 -1 1440 -1 0 15776
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_51
timestamp 1707688321
transform 0 -1 1440 -1 0 11881
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_52
timestamp 1707688321
transform 0 -1 1440 -1 0 4091
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_53
timestamp 1707688321
transform 0 -1 1440 -1 0 7986
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_54
timestamp 1707688321
transform 0 -1 1314 -1 0 27461
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_55
timestamp 1707688321
transform 0 -1 1314 -1 0 23566
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_56
timestamp 1707688321
transform 0 -1 1314 -1 0 19671
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_57
timestamp 1707688321
transform 0 -1 1314 -1 0 15776
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_58
timestamp 1707688321
transform 0 -1 1314 -1 0 11881
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_59
timestamp 1707688321
transform 0 -1 1314 -1 0 4091
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_60
timestamp 1707688321
transform 0 -1 1314 -1 0 7986
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_61
timestamp 1707688321
transform 0 -1 2070 -1 0 11881
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_62
timestamp 1707688321
transform 0 -1 2070 -1 0 15776
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_63
timestamp 1707688321
transform 0 -1 2070 -1 0 19671
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_64
timestamp 1707688321
transform 0 -1 2070 -1 0 23566
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_65
timestamp 1707688321
transform 0 -1 2070 -1 0 27461
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_66
timestamp 1707688321
transform 0 -1 1944 -1 0 27461
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_67
timestamp 1707688321
transform 0 -1 1944 -1 0 19671
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_68
timestamp 1707688321
transform 0 -1 1944 -1 0 15776
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_69
timestamp 1707688321
transform 0 -1 1944 -1 0 11881
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_70
timestamp 1707688321
transform 0 -1 1944 -1 0 4091
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_71
timestamp 1707688321
transform 0 -1 1944 -1 0 7986
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_72
timestamp 1707688321
transform 0 -1 1818 -1 0 27461
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_73
timestamp 1707688321
transform 0 -1 1818 -1 0 23566
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_74
timestamp 1707688321
transform 0 -1 1818 -1 0 19671
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_75
timestamp 1707688321
transform 0 -1 1818 -1 0 15776
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_76
timestamp 1707688321
transform 0 -1 1818 -1 0 11881
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_77
timestamp 1707688321
transform 0 -1 1818 -1 0 4091
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_78
timestamp 1707688321
transform 0 -1 1818 -1 0 7986
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_79
timestamp 1707688321
transform 0 -1 558 -1 0 4091
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_80
timestamp 1707688321
transform 0 -1 558 -1 0 7986
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_81
timestamp 1707688321
transform 0 -1 558 -1 0 11881
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_82
timestamp 1707688321
transform 0 -1 558 -1 0 15776
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_83
timestamp 1707688321
transform 0 -1 558 -1 0 19671
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_84
timestamp 1707688321
transform 0 -1 558 -1 0 23566
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_85
timestamp 1707688321
transform 0 -1 558 -1 0 27461
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_86
timestamp 1707688321
transform 0 -1 432 -1 0 27461
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_87
timestamp 1707688321
transform 0 -1 432 -1 0 23566
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_88
timestamp 1707688321
transform 0 -1 432 -1 0 19671
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_89
timestamp 1707688321
transform 0 -1 432 -1 0 15776
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_90
timestamp 1707688321
transform 0 -1 432 -1 0 11881
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_91
timestamp 1707688321
transform 0 -1 432 -1 0 7986
box -68 -26 3683 92
use nDFres_CDNS_52468879185986  nDFres_CDNS_52468879185986_92
timestamp 1707688321
transform 0 -1 432 -1 0 4091
box -68 -26 3683 92
use nDFres_CDNS_52468879185987  nDFres_CDNS_52468879185987_0
timestamp 1707688321
transform 0 -1 1692 -1 0 23566
box -68 -26 1259 92
use nDFres_CDNS_52468879185987  nDFres_CDNS_52468879185987_1
timestamp 1707688321
transform 0 -1 1440 -1 0 23566
box -68 -26 1259 92
use nDFres_CDNS_52468879185987  nDFres_CDNS_52468879185987_2
timestamp 1707688321
transform 0 -1 1944 -1 0 23566
box -68 -26 1259 92
use nDFres_CDNS_52468879185988  nDFres_CDNS_52468879185988_0
timestamp 1707688321
transform 0 -1 2070 -1 0 5355
box -68 -26 4947 92
use nDFres_CDNS_52468879185988  nDFres_CDNS_52468879185988_1
timestamp 1707688321
transform 0 -1 2196 -1 0 5355
box -68 -26 4947 92
use nDFres_CDNS_52468879185988  nDFres_CDNS_52468879185988_2
timestamp 1707688321
transform 0 -1 2322 -1 0 5355
box -68 -26 4947 92
use nDFres_CDNS_52468879185988  nDFres_CDNS_52468879185988_3
timestamp 1707688321
transform 0 -1 2448 -1 0 5355
box -68 -26 4947 92
use nDFres_CDNS_52468879185988  nDFres_CDNS_52468879185988_4
timestamp 1707688321
transform 0 -1 2574 -1 0 5355
box -68 -26 4947 92
use nDFres_CDNS_52468879185988  nDFres_CDNS_52468879185988_5
timestamp 1707688321
transform 0 -1 2700 -1 0 5355
box -68 -26 4947 92
use nDFres_CDNS_52468879185988  nDFres_CDNS_52468879185988_6
timestamp 1707688321
transform 0 -1 2826 -1 0 5355
box -68 -26 4947 92
use nDFres_CDNS_52468879185988  nDFres_CDNS_52468879185988_7
timestamp 1707688321
transform 0 -1 2952 -1 0 5355
box -68 -26 4947 92
use nDFres_CDNS_52468879185988  nDFres_CDNS_52468879185988_8
timestamp 1707688321
transform 0 -1 3078 -1 0 5355
box -68 -26 4947 92
use nfet_CDNS_52468879185989  nfet_CDNS_52468879185989_0
timestamp 1707688321
transform -1 0 4561 0 1 8722
box -79 -26 1735 2026
use nfet_CDNS_52468879185989  nfet_CDNS_52468879185989_1
timestamp 1707688321
transform -1 0 4561 0 -1 8592
box -79 -26 1735 2026
use nfet_CDNS_52468879185989  nfet_CDNS_52468879185989_2
timestamp 1707688321
transform 1 0 4881 0 -1 8592
box -79 -26 1735 2026
use nfet_CDNS_52468879185989  nfet_CDNS_52468879185989_3
timestamp 1707688321
transform 1 0 4881 0 1 8722
box -79 -26 1735 2026
use nfet_CDNS_52468879185992  nfet_CDNS_52468879185992_0
timestamp 1707688321
transform 1 0 3693 0 1 4410
box -79 -26 1271 1026
use nfet_CDNS_52468879185993  nfet_CDNS_52468879185993_0
timestamp 1707688321
transform 1 0 4941 0 1 4410
box -79 -26 375 1026
use nfet_CDNS_52468879185994  nfet_CDNS_52468879185994_0
timestamp 1707688321
transform 1 0 5293 0 1 4410
box -79 -26 279 1026
use nfet_CDNS_52468879185995  nfet_CDNS_52468879185995_0
timestamp 1707688321
transform 1 0 2959 0 1 -920
box -79 -26 455 226
use nfet_CDNS_52468879185996  nfet_CDNS_52468879185996_0
timestamp 1707688321
transform 1 0 2527 0 1 -920
box -79 -26 455 226
use nfet_CDNS_52468879185997  nfet_CDNS_52468879185997_0
timestamp 1707688321
transform -1 0 2471 0 1 -920
box -79 -26 239 226
use pfet_CDNS_52468879185998  pfet_CDNS_52468879185998_0
timestamp 1707688321
transform 1 0 2137 0 1 -230
box -119 -66 319 266
use pfet_CDNS_52468879185999  pfet_CDNS_52468879185999_0
timestamp 1707688321
transform -1 0 3359 0 1 -230
box -119 -66 519 266
use pfet_CDNS_524688791851000  pfet_CDNS_524688791851000_0
timestamp 1707688321
transform 1 0 2503 0 1 -230
box -119 -66 519 266
use pfet_CDNS_524688791851001  pfet_CDNS_524688791851001_0
timestamp 1707688321
transform 1 0 905 0 1 -230
box -119 -66 1119 266
use pfet_CDNS_524688791851002  pfet_CDNS_524688791851002_0
timestamp 1707688321
transform 1 0 905 0 1 -564
box -119 -66 767 266
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_0
timestamp 1707688321
transform 0 1 5293 -1 0 5508
box 0 0 1 1
use PYL1_CDNS_52468879185309  PYL1_CDNS_52468879185309_0
timestamp 1707688321
transform 0 -1 5224 -1 0 5508
box 0 0 1 1
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_0
timestamp 1707688321
transform 0 1 5764 -1 0 6558
box 0 0 66 746
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_1
timestamp 1707688321
transform 0 1 4908 -1 0 6558
box 0 0 66 746
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_2
timestamp 1707688321
transform 0 1 3788 -1 0 6558
box 0 0 66 746
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_3
timestamp 1707688321
transform 0 1 2932 -1 0 6558
box 0 0 66 746
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_4
timestamp 1707688321
transform 0 1 3788 1 0 10754
box 0 0 66 746
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_5
timestamp 1707688321
transform 0 1 2932 1 0 10754
box 0 0 66 746
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_6
timestamp 1707688321
transform 0 1 5764 1 0 10754
box 0 0 66 746
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_7
timestamp 1707688321
transform 0 1 4908 1 0 10754
box 0 0 66 746
use PYL1_CDNS_52468879185331  PYL1_CDNS_52468879185331_0
timestamp 1707688321
transform 0 -1 4866 1 0 5442
box 0 0 66 1154
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_0
timestamp 1707688321
transform 0 -1 5580 1 0 4511
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185979  sky130_fd_io__tk_em1o_CDNS_52468879185979_0
timestamp 1707688321
transform 0 -1 6337 -1 0 6580
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185979  sky130_fd_io__tk_em1o_CDNS_52468879185979_1
timestamp 1707688321
transform 0 1 3105 -1 0 6580
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185979  sky130_fd_io__tk_em1o_CDNS_52468879185979_2
timestamp 1707688321
transform 0 1 3105 1 0 6574
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185979  sky130_fd_io__tk_em1o_CDNS_52468879185979_3
timestamp 1707688321
transform 0 -1 6337 1 0 6574
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185980  sky130_fd_io__tk_em1o_CDNS_52468879185980_0
timestamp 1707688321
transform 0 -1 6481 -1 0 10740
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185980  sky130_fd_io__tk_em1o_CDNS_52468879185980_1
timestamp 1707688321
transform 0 1 2961 -1 0 10740
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185980  sky130_fd_io__tk_em1o_CDNS_52468879185980_2
timestamp 1707688321
transform 0 1 2961 1 0 10734
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185980  sky130_fd_io__tk_em1o_CDNS_52468879185980_3
timestamp 1707688321
transform 0 -1 6481 1 0 10734
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185981  sky130_fd_io__tk_em1o_CDNS_52468879185981_0
timestamp 1707688321
transform 0 -1 538 -1 0 27439
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185981  sky130_fd_io__tk_em1o_CDNS_52468879185981_1
timestamp 1707688321
transform 0 -1 664 1 0 498
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185981  sky130_fd_io__tk_em1o_CDNS_52468879185981_2
timestamp 1707688321
transform 0 -1 1168 1 0 498
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185981  sky130_fd_io__tk_em1o_CDNS_52468879185981_3
timestamp 1707688321
transform 0 -1 1420 1 0 498
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185981  sky130_fd_io__tk_em1o_CDNS_52468879185981_4
timestamp 1707688321
transform 0 -1 1672 1 0 498
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185982  sky130_fd_io__tk_em1o_CDNS_52468879185982_0
timestamp 1707688321
transform 0 -1 1937 1 0 16078
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185982  sky130_fd_io__tk_em1o_CDNS_52468879185982_1
timestamp 1707688321
transform 0 -1 1937 1 0 12183
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185982  sky130_fd_io__tk_em1o_CDNS_52468879185982_2
timestamp 1707688321
transform 0 -1 1937 1 0 8288
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185983  sky130_fd_io__tk_em1o_CDNS_52468879185983_0
timestamp 1707688321
transform 1 0 1888 0 -1 5570
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185984  sky130_fd_io__tk_em1o_CDNS_52468879185984_0
timestamp 1707688321
transform 0 -1 1048 -1 0 27439
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_0
timestamp 1707688321
transform 0 -1 554 -1 0 23544
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_1
timestamp 1707688321
transform 0 -1 554 -1 0 7964
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_2
timestamp 1707688321
transform 0 -1 554 -1 0 11859
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_3
timestamp 1707688321
transform 0 -1 554 -1 0 3995
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_4
timestamp 1707688321
transform 0 -1 806 -1 0 3995
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_5
timestamp 1707688321
transform 0 -1 806 -1 0 7964
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_6
timestamp 1707688321
transform 0 -1 806 -1 0 11859
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_7
timestamp 1707688321
transform 0 -1 806 -1 0 15754
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_8
timestamp 1707688321
transform 0 -1 806 -1 0 19649
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_9
timestamp 1707688321
transform 0 -1 1058 -1 0 7964
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_10
timestamp 1707688321
transform 0 -1 1058 -1 0 11859
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_11
timestamp 1707688321
transform 0 -1 1058 -1 0 15754
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_12
timestamp 1707688321
transform 0 -1 1058 -1 0 19649
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_13
timestamp 1707688321
transform 0 -1 1058 -1 0 23544
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_14
timestamp 1707688321
transform 0 -1 1310 -1 0 3995
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_15
timestamp 1707688321
transform 0 -1 1562 -1 0 3995
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_16
timestamp 1707688321
transform 0 -1 1814 -1 0 3995
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_17
timestamp 1707688321
transform 0 -1 2822 -1 0 3995
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_18
timestamp 1707688321
transform 0 -1 2570 -1 0 3995
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_19
timestamp 1707688321
transform 0 -1 2066 -1 0 3995
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_20
timestamp 1707688321
transform 0 -1 2318 -1 0 3995
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_21
timestamp 1707688321
transform 0 -1 1940 1 0 3851
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_22
timestamp 1707688321
transform 0 -1 2948 1 0 3798
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_23
timestamp 1707688321
transform 0 -1 680 1 0 23868
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_24
timestamp 1707688321
transform 0 -1 680 1 0 12183
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_25
timestamp 1707688321
transform 0 -1 680 1 0 16078
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_26
timestamp 1707688321
transform 0 -1 680 1 0 19973
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_27
timestamp 1707688321
transform 0 -1 932 1 0 23868
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_28
timestamp 1707688321
transform 0 -1 932 1 0 19973
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_29
timestamp 1707688321
transform 0 -1 932 1 0 16078
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_30
timestamp 1707688321
transform 0 -1 932 1 0 4393
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_31
timestamp 1707688321
transform 0 -1 932 1 0 12183
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_32
timestamp 1707688321
transform 0 -1 932 1 0 8288
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_33
timestamp 1707688321
transform 0 -1 1184 1 0 16078
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_34
timestamp 1707688321
transform 0 -1 1184 1 0 12183
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_35
timestamp 1707688321
transform 0 -1 1184 1 0 8288
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_36
timestamp 1707688321
transform 0 -1 1184 1 0 4341
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_37
timestamp 1707688321
transform 0 -1 1436 1 0 16078
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_38
timestamp 1707688321
transform 0 -1 1436 1 0 12183
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_39
timestamp 1707688321
transform 0 -1 1436 1 0 8288
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_40
timestamp 1707688321
transform 0 -1 1436 1 0 4413
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_41
timestamp 1707688321
transform 0 -1 1688 1 0 16078
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_42
timestamp 1707688321
transform 0 -1 1688 1 0 12183
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_43
timestamp 1707688321
transform 0 -1 1688 1 0 8288
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_44
timestamp 1707688321
transform 0 -1 1688 1 0 4413
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_45
timestamp 1707688321
transform 0 -1 2444 1 0 4026
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_46
timestamp 1707688321
transform 0 -1 2192 1 0 4026
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_47
timestamp 1707688321
transform 0 -1 2696 1 0 4026
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_48
timestamp 1707688321
transform 0 -1 2948 1 0 3973
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_49
timestamp 1707688321
transform 0 -1 2696 1 0 3851
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_50
timestamp 1707688321
transform 0 -1 2192 1 0 4413
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_51
timestamp 1707688321
transform 0 -1 2444 1 0 4413
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_0
timestamp 1707688321
transform -1 0 5100 0 1 10711
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_1
timestamp 1707688321
transform -1 0 5100 0 -1 6603
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_2
timestamp 1707688321
transform 1 0 4342 0 -1 6603
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_3
timestamp 1707688321
transform 1 0 4342 0 1 10711
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185976  sky130_fd_io__tk_em1s_CDNS_52468879185976_0
timestamp 1707688321
transform 0 1 2854 1 0 6574
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185976  sky130_fd_io__tk_em1s_CDNS_52468879185976_1
timestamp 1707688321
transform 0 -1 6588 1 0 6574
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185977  sky130_fd_io__tk_em1s_CDNS_52468879185977_0
timestamp 1707688321
transform 0 -1 6588 -1 0 8729
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185977  sky130_fd_io__tk_em1s_CDNS_52468879185977_1
timestamp 1707688321
transform 0 1 2854 -1 0 8729
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185978  sky130_fd_io__tk_em1s_CDNS_52468879185978_0
timestamp 1707688321
transform 0 -1 1940 1 0 4026
box 0 0 1 1
<< labels >>
flabel comment s 3179 10782 3179 10782 0 FreeSans 1000 0 0 0 condiode
flabel comment s 399 4334 399 4334 0 FreeSans 100 90 0 0 li_jumper_ok
flabel comment s 3042 4359 3042 4359 0 FreeSans 100 90 0 0 li_jumper_ok
flabel comment s 2029 8229 2029 8229 0 FreeSans 100 90 0 0 resistive_li1_ok
flabel comment s 2418 4485 2418 4485 0 FreeSans 400 0 0 0 I16
flabel comment s 2291 3920 2291 3920 0 FreeSans 400 0 0 0 I17
flabel comment s 2167 4487 2167 4487 0 FreeSans 400 0 0 0 I18
flabel comment s 2042 3922 2042 3922 0 FreeSans 400 0 0 0 I19
flabel comment s 1954 5499 1954 5499 0 FreeSans 400 0 0 0 I20
flabel comment s 1922 3925 1922 3925 0 FreeSans 400 0 0 0 I21
flabel comment s 2540 3923 2540 3923 0 FreeSans 400 0 0 0 I22
flabel comment s 2667 3923 2667 3923 0 FreeSans 400 0 0 0 I23
flabel comment s 2809 3925 2809 3925 0 FreeSans 400 0 0 0 I24
flabel comment s 2915 3871 2915 3871 0 FreeSans 400 0 0 0 I25
flabel comment s 1914 4099 1914 4099 0 FreeSans 400 0 0 0 I44
flabel comment s 2670 4097 2670 4097 0 FreeSans 400 0 0 0 I45
flabel comment s 2923 4049 2923 4049 0 FreeSans 400 0 0 0 I46
flabel comment s 2166 4095 2166 4095 0 FreeSans 400 0 0 0 I43
flabel comment s 2416 4097 2416 4097 0 FreeSans 400 0 0 0 I42
flabel comment s 7285 10678 7285 10678 3 FreeSans 200 180 0 0 en_inpop_h
flabel comment s 2067 11011 2067 11011 3 FreeSans 200 270 0 0 en_outop_h
flabel comment s 7299 6135 7299 6135 3 FreeSans 200 180 0 0 ibuf_sel_h
flabel comment s 7299 6054 7299 6054 3 FreeSans 200 180 0 0 vtrip_sel_h_n
flabel comment s 7299 5902 7299 5902 3 FreeSans 200 180 0 0 vtrip_sel_h
flabel comment s 7299 6335 7299 6335 3 FreeSans 200 180 0 0 en_outop_h
flabel comment s 1714 27774 1714 27774 3 FreeSans 200 0 0 0 en_inpop_h
flabel comment s 6664 5788 6664 5788 3 FreeSans 200 90 0 0 vpwr
flabel comment s 1910 11828 1910 11828 3 FreeSans 200 270 0 0 R<7>
flabel comment s 1913 23513 1913 23513 3 FreeSans 200 270 0 0 R<7>
flabel comment s 1913 27408 1913 27408 3 FreeSans 200 270 0 0 R<7>
flabel comment s 1784 23899 1784 23899 3 FreeSans 200 90 0 0 R<7>
flabel comment s 1784 20004 1784 20004 3 FreeSans 200 90 0 0 R<7>
flabel comment s 1784 16109 1784 16109 3 FreeSans 200 90 0 0 R<7>
flabel comment s 1784 12214 1784 12214 3 FreeSans 200 90 0 0 R<7>
flabel comment s 1784 8319 1784 8319 3 FreeSans 200 90 0 0 R<7>
flabel comment s 1784 4187 1784 4187 3 FreeSans 200 90 0 0 R<7>
flabel comment s 1784 529 1784 529 3 FreeSans 200 90 0 0 R<7>
flabel comment s 1658 4032 1658 4032 3 FreeSans 200 270 0 0 R<7>
flabel comment s 1658 7933 1658 7933 3 FreeSans 200 270 0 0 R<7>
flabel comment s 1659 23513 1659 23513 3 FreeSans 200 270 0 0 R<5>
flabel comment s 1660 23513 1660 23513 3 FreeSans 200 270 0 0 R<6>
flabel comment s 1660 27408 1660 27408 3 FreeSans 200 270 0 0 R<6>
flabel comment s 1532 23899 1532 23899 3 FreeSans 200 90 0 0 R<6>
flabel comment s 1532 20004 1532 20004 3 FreeSans 200 90 0 0 R<6>
flabel comment s 1532 16109 1532 16109 3 FreeSans 200 90 0 0 R<6>
flabel comment s 1532 12214 1532 12214 3 FreeSans 200 90 0 0 R<6>
flabel comment s 1532 8319 1532 8319 3 FreeSans 200 90 0 0 R<6>
flabel comment s 1532 4187 1532 4187 3 FreeSans 200 90 0 0 R<6>
flabel comment s 1658 11828 1658 11828 3 FreeSans 200 270 0 0 R<6>
flabel comment s 1658 15723 1658 15723 3 FreeSans 200 270 0 0 R<6>
flabel comment s 1658 19618 1658 19618 3 FreeSans 200 270 0 0 R<6>
flabel comment s 1532 529 1532 529 3 FreeSans 200 90 0 0 R<6>
flabel comment s 1406 4032 1406 4032 3 FreeSans 200 270 0 0 R<6>
flabel comment s 1406 7933 1406 7933 3 FreeSans 200 270 0 0 R<6>
flabel comment s 1407 23513 1407 23513 3 FreeSans 200 270 0 0 R<5>
flabel comment s 1407 27408 1407 27408 3 FreeSans 200 270 0 0 R<5>
flabel comment s 1280 23899 1280 23899 3 FreeSans 200 90 0 0 R<5>
flabel comment s 1280 20004 1280 20004 3 FreeSans 200 90 0 0 R<5>
flabel comment s 1280 16109 1280 16109 3 FreeSans 200 90 0 0 R<5>
flabel comment s 1280 12214 1280 12214 3 FreeSans 200 90 0 0 R<5>
flabel comment s 1280 8319 1280 8319 3 FreeSans 200 90 0 0 R<5>
flabel comment s 1280 4424 1280 4424 3 FreeSans 200 90 0 0 R<5>
flabel comment s 1406 11828 1406 11828 3 FreeSans 200 270 0 0 R<5>
flabel comment s 1406 15723 1406 15723 3 FreeSans 200 270 0 0 R<5>
flabel comment s 1406 19618 1406 19618 3 FreeSans 200 270 0 0 R<5>
flabel comment s 1280 529 1280 529 3 FreeSans 200 90 0 0 R<5>
flabel comment s 1154 4032 1154 4032 3 FreeSans 200 270 0 0 R<5>
flabel comment s 1154 7933 1154 7933 3 FreeSans 200 270 0 0 R<5>
flabel comment s 1154 27408 1154 27408 3 FreeSans 200 270 0 0 R<4>
flabel comment s 1154 23513 1154 23513 3 FreeSans 200 270 0 0 R<4>
flabel comment s 1154 11828 1154 11828 3 FreeSans 200 270 0 0 R<4>
flabel comment s 1154 15723 1154 15723 3 FreeSans 200 270 0 0 R<4>
flabel comment s 1154 19618 1154 19618 3 FreeSans 200 270 0 0 R<4>
flabel comment s 1028 23899 1028 23899 3 FreeSans 200 90 0 0 R<4>
flabel comment s 1028 20004 1028 20004 3 FreeSans 200 90 0 0 R<4>
flabel comment s 1028 16109 1028 16109 3 FreeSans 200 90 0 0 R<4>
flabel comment s 1028 12214 1028 12214 3 FreeSans 200 90 0 0 R<3>
flabel comment s 1028 8319 1028 8319 3 FreeSans 200 90 0 0 R<3>
flabel comment s 1028 4424 1028 4424 3 FreeSans 200 90 0 0 R<3>
flabel comment s 899 7939 899 7939 3 FreeSans 200 270 0 0 R<3>
flabel comment s 899 11834 899 11834 3 FreeSans 200 270 0 0 R<3>
flabel comment s 899 15723 899 15723 3 FreeSans 200 270 0 0 R<3>
flabel comment s 899 19618 899 19618 3 FreeSans 200 270 0 0 R<2>
flabel comment s 899 23513 899 23513 3 FreeSans 200 270 0 0 R<2>
flabel comment s 899 27408 899 27408 3 FreeSans 200 270 0 0 R<2>
flabel comment s 772 23899 772 23899 3 FreeSans 200 90 0 0 R<2>
flabel comment s 772 19998 772 19998 3 FreeSans 200 90 0 0 R<2>
flabel comment s 772 16109 772 16109 3 FreeSans 200 90 0 0 R<2>
flabel comment s 772 12214 772 12214 3 FreeSans 200 90 0 0 R<2>
flabel comment s 772 8319 772 8319 3 FreeSans 200 90 0 0 R<2>
flabel comment s 772 4430 772 4430 3 FreeSans 200 90 0 0 R<1>
flabel comment s 772 535 772 535 3 FreeSans 200 90 0 0 R<1>
flabel comment s 649 4026 649 4026 3 FreeSans 200 270 0 0 R<1>
flabel comment s 649 7927 649 7927 3 FreeSans 200 270 0 0 R<1>
flabel comment s 649 11822 649 11822 3 FreeSans 200 270 0 0 R<1>
flabel comment s 649 15717 649 15717 3 FreeSans 200 270 0 0 R<1>
flabel comment s 649 19612 649 19612 3 FreeSans 200 270 0 0 R<1>
flabel comment s 649 23513 649 23513 3 FreeSans 200 270 0 0 R<1>
flabel comment s 649 27408 649 27408 3 FreeSans 200 270 0 0 R<0>
flabel comment s 524 23899 524 23899 3 FreeSans 200 90 0 0 R<0>
flabel comment s 524 20004 524 20004 3 FreeSans 200 90 0 0 R<0>
flabel comment s 524 16109 524 16109 3 FreeSans 200 90 0 0 R<0>
flabel comment s 524 12214 524 12214 3 FreeSans 200 90 0 0 R<0>
flabel comment s 524 8319 524 8319 3 FreeSans 200 90 0 0 R<0>
flabel comment s 524 4424 524 4424 3 FreeSans 200 90 0 0 R<0>
flabel comment s 524 523 524 523 3 FreeSans 200 90 0 0 R<0>
flabel comment s 899 4038 899 4038 3 FreeSans 200 270 0 0 R<3>
flabel comment s 1028 523 1028 523 3 FreeSans 200 90 0 0 R<3>
flabel comment s 1910 19618 1910 19618 3 FreeSans 200 270 0 0 R<7>
flabel comment s 1910 15723 1910 15723 3 FreeSans 200 270 0 0 R<7>
flabel metal1 s 59 4141 85 4193 3 FreeSans 200 0 0 0 vinref
port 3 nsew
flabel metal1 s 5661 4221 5682 4267 3 FreeSans 200 180 0 0 vcc_io_0p5
port 4 nsew
flabel metal1 s 5656 5304 5682 5350 3 FreeSans 200 180 0 0 sel_vcc_io_0p4
port 5 nsew
flabel metal1 s 5656 5378 5682 5424 3 FreeSans 200 180 0 0 sel_vcc_io
port 6 nsew
flabel metal1 s 5662 5608 5682 5654 3 FreeSans 200 180 0 0 in_lpf
port 7 nsew
flabel metal1 s 5661 4141 5682 4193 3 FreeSans 200 180 0 0 vinref
port 3 nsew
flabel metal1 s 7269 5947 7306 5999 3 FreeSans 200 180 0 0 ibuf_sel_h_n
port 2 nsew
flabel metal1 s 7273 7148 7306 7424 7 FreeSans 200 0 0 0 vcc_a
port 8 nsew
flabel metal2 s 7176 10797 7306 10838 3 FreeSans 200 270 0 0 vgnd
port 9 nsew
flabel metal2 s 1338 27767 1477 27784 3 FreeSans 200 270 0 0 vgnd
port 9 nsew
flabel metal2 s 5994 5750 6046 5771 3 FreeSans 200 90 0 0 ibuf_sel_h_n
port 2 nsew
flabel metal2 s 7176 10976 7306 11017 3 FreeSans 200 270 0 0 vgnd
port 9 nsew
flabel metal2 s 7176 5750 7306 5791 3 FreeSans 200 90 0 0 vgnd
port 9 nsew
flabel metal2 s 3424 4274 3806 4295 3 FreeSans 200 90 0 0 vgnd
port 9 nsew
flabel metal2 s 3862 4274 4412 4295 3 FreeSans 200 90 0 0 vgnd
port 9 nsew
flabel metal2 s 5156 4274 5293 4295 3 FreeSans 200 90 0 0 vgnd
port 9 nsew
flabel metal2 s 5622 10976 6085 11017 3 FreeSans 200 270 0 0 vgnd
port 9 nsew
flabel metal2 s 5764 5750 5966 5771 3 FreeSans 200 90 0 0 vgnd
port 9 nsew
flabel metal2 s 3862 10976 4412 11017 3 FreeSans 200 270 0 0 vgnd
port 9 nsew
flabel metal2 s 3424 10976 3806 11017 3 FreeSans 200 270 0 0 vgnd
port 9 nsew
flabel metal2 s 2488 10976 2850 11017 3 FreeSans 200 270 0 0 vgnd
port 9 nsew
flabel metal2 s 3014 10976 3260 11017 3 FreeSans 200 270 0 0 vgnd
port 9 nsew
flabel metal2 s 718 27767 1282 27784 3 FreeSans 200 270 0 0 vgnd
port 9 nsew
flabel metal2 s 5104 10976 5486 11017 3 FreeSans 200 270 0 0 vgnd
port 9 nsew
flabel metal2 s 6249 10976 6911 11017 3 FreeSans 200 270 0 0 vgnd
port 9 nsew
flabel metal2 s 2125 10976 2432 11017 7 FreeSans 200 90 0 0 vcc_a
port 8 nsew
flabel metal2 s 6967 10976 7117 11017 7 FreeSans 200 90 0 0 vcc_a
port 8 nsew
flabel metal2 s 4468 10976 4968 11017 7 FreeSans 200 90 0 0 vcc_a
port 8 nsew
flabel metal2 s 6967 5750 7117 5771 3 FreeSans 200 90 0 0 vcc_a
port 8 nsew
flabel metal2 s 6253 5750 6305 5771 3 FreeSans 200 90 0 0 ibuf_sel_h
port 10 nsew
flabel metal2 s 4468 4274 4600 4295 3 FreeSans 200 90 0 0 vcc_a
port 8 nsew
flabel metal2 s 59 4456 379 4516 0 FreeSans 200 0 0 0 vcc_io
port 11 nsew
flabel metal2 s 2121 4343 2437 4412 0 FreeSans 200 0 0 0 vcc_io
port 11 nsew
<< properties >>
string GDS_END 78907590
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 78610534
string path 44.900 692.300 49.700 692.300 
<< end >>
