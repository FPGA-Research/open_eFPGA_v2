magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -66 377 2562 897
<< pwell >>
rect 2032 225 2492 301
rect 1598 217 2492 225
rect 4 43 2492 217
rect -26 -43 2522 43
<< mvnmos >>
rect 83 107 183 191
rect 239 107 339 191
rect 381 107 481 191
rect 537 107 637 191
rect 679 107 779 191
rect 883 107 983 191
rect 1025 107 1125 191
rect 1181 107 1281 191
rect 1323 107 1423 191
rect 1681 115 1781 199
rect 1837 115 1937 199
rect 2115 191 2215 275
rect 2313 125 2413 275
<< mvpmos >>
rect 83 627 183 711
rect 239 627 339 711
rect 381 627 481 711
rect 537 627 637 711
rect 699 627 799 711
rect 855 627 955 711
rect 997 627 1097 711
rect 1153 627 1253 711
rect 1295 627 1395 711
rect 1569 615 1669 699
rect 1725 615 1825 699
rect 2115 443 2215 527
rect 2313 443 2413 743
<< mvndiff >>
rect 2058 250 2115 275
rect 2058 216 2070 250
rect 2104 216 2115 250
rect 30 166 83 191
rect 30 132 38 166
rect 72 132 83 166
rect 30 107 83 132
rect 183 166 239 191
rect 183 132 194 166
rect 228 132 239 166
rect 183 107 239 132
rect 339 107 381 191
rect 481 166 537 191
rect 481 132 492 166
rect 526 132 537 166
rect 481 107 537 132
rect 637 107 679 191
rect 779 166 883 191
rect 779 132 790 166
rect 824 132 883 166
rect 779 107 883 132
rect 983 107 1025 191
rect 1125 170 1181 191
rect 1125 136 1136 170
rect 1170 136 1181 170
rect 1125 107 1181 136
rect 1281 107 1323 191
rect 1423 166 1480 191
rect 1423 132 1434 166
rect 1468 132 1480 166
rect 1423 107 1480 132
rect 1624 182 1681 199
rect 1624 148 1636 182
rect 1670 148 1681 182
rect 1624 115 1681 148
rect 1781 157 1837 199
rect 1781 123 1792 157
rect 1826 123 1837 157
rect 1781 115 1837 123
rect 1937 174 1994 199
rect 2058 191 2115 216
rect 2215 267 2313 275
rect 2215 233 2268 267
rect 2302 233 2313 267
rect 2215 191 2313 233
rect 1937 140 1948 174
rect 1982 140 1994 174
rect 2256 167 2313 191
rect 1937 115 1994 140
rect 2256 133 2268 167
rect 2302 133 2313 167
rect 2256 125 2313 133
rect 2413 263 2466 275
rect 2413 229 2424 263
rect 2458 229 2466 263
rect 2413 171 2466 229
rect 2413 137 2424 171
rect 2458 137 2466 171
rect 2413 125 2466 137
<< mvpdiff >>
rect 2237 735 2313 743
rect 30 686 83 711
rect 30 652 38 686
rect 72 652 83 686
rect 30 627 83 652
rect 183 686 239 711
rect 183 652 194 686
rect 228 652 239 686
rect 183 627 239 652
rect 339 627 381 711
rect 481 680 537 711
rect 481 646 492 680
rect 526 646 537 680
rect 481 627 537 646
rect 637 627 699 711
rect 799 686 855 711
rect 799 652 810 686
rect 844 652 855 686
rect 799 627 855 652
rect 955 627 997 711
rect 1097 686 1153 711
rect 1097 652 1108 686
rect 1142 652 1153 686
rect 1097 627 1153 652
rect 1253 627 1295 711
rect 1395 686 1452 711
rect 2237 701 2249 735
rect 2283 701 2313 735
rect 1395 652 1406 686
rect 1440 652 1452 686
rect 1395 627 1452 652
rect 1512 674 1569 699
rect 1512 640 1524 674
rect 1558 640 1569 674
rect 1512 615 1569 640
rect 1669 686 1725 699
rect 1669 652 1680 686
rect 1714 652 1725 686
rect 1669 615 1725 652
rect 1825 674 1956 699
rect 1825 640 1910 674
rect 1944 640 1956 674
rect 1825 615 1956 640
rect 2237 652 2313 701
rect 2237 618 2249 652
rect 2283 618 2313 652
rect 2237 568 2313 618
rect 2237 534 2249 568
rect 2283 534 2313 568
rect 2237 527 2313 534
rect 2062 502 2115 527
rect 2062 468 2070 502
rect 2104 468 2115 502
rect 2062 443 2115 468
rect 2215 485 2313 527
rect 2215 451 2249 485
rect 2283 451 2313 485
rect 2215 443 2313 451
rect 2413 731 2466 743
rect 2413 697 2424 731
rect 2458 697 2466 731
rect 2413 651 2466 697
rect 2413 617 2424 651
rect 2458 617 2466 651
rect 2413 569 2466 617
rect 2413 535 2424 569
rect 2458 535 2466 569
rect 2413 489 2466 535
rect 2413 455 2424 489
rect 2458 455 2466 489
rect 2413 443 2466 455
<< mvndiffc >>
rect 2070 216 2104 250
rect 38 132 72 166
rect 194 132 228 166
rect 492 132 526 166
rect 790 132 824 166
rect 1136 136 1170 170
rect 1434 132 1468 166
rect 1636 148 1670 182
rect 1792 123 1826 157
rect 2268 233 2302 267
rect 1948 140 1982 174
rect 2268 133 2302 167
rect 2424 229 2458 263
rect 2424 137 2458 171
<< mvpdiffc >>
rect 38 652 72 686
rect 194 652 228 686
rect 492 646 526 680
rect 810 652 844 686
rect 1108 652 1142 686
rect 2249 701 2283 735
rect 1406 652 1440 686
rect 1524 640 1558 674
rect 1680 652 1714 686
rect 1910 640 1944 674
rect 2249 618 2283 652
rect 2249 534 2283 568
rect 2070 468 2104 502
rect 2249 451 2283 485
rect 2424 697 2458 731
rect 2424 617 2458 651
rect 2424 535 2458 569
rect 2424 455 2458 489
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2496 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2496 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
<< poly >>
rect 2313 743 2413 769
rect 83 711 183 737
rect 239 711 339 737
rect 381 711 481 737
rect 537 711 637 737
rect 699 711 799 737
rect 855 711 955 737
rect 997 711 1097 737
rect 1153 711 1253 737
rect 1295 711 1395 737
rect 1569 699 1669 725
rect 1725 699 1825 725
rect 83 575 183 627
rect 239 601 339 627
rect 83 541 129 575
rect 163 541 183 575
rect 83 507 183 541
rect 83 473 129 507
rect 163 473 183 507
rect 83 191 183 473
rect 233 418 339 601
rect 381 579 481 627
rect 381 545 397 579
rect 431 545 481 579
rect 381 516 481 545
rect 537 528 637 627
rect 699 601 799 627
rect 699 572 805 601
rect 699 538 719 572
rect 753 538 805 572
rect 381 511 447 516
rect 381 477 397 511
rect 431 477 447 511
rect 381 461 447 477
rect 537 508 657 528
rect 537 474 607 508
rect 641 474 657 508
rect 489 440 657 474
rect 699 504 805 538
rect 699 470 719 504
rect 753 470 805 504
rect 699 450 805 470
rect 489 419 607 440
rect 233 384 253 418
rect 287 384 339 418
rect 233 350 339 384
rect 233 316 253 350
rect 287 316 339 350
rect 233 296 339 316
rect 239 191 339 296
rect 381 406 607 419
rect 641 406 657 440
rect 381 391 657 406
rect 381 357 397 391
rect 431 381 657 391
rect 431 357 499 381
rect 381 323 499 357
rect 381 289 397 323
rect 431 311 499 323
rect 541 323 637 339
rect 431 289 481 311
rect 381 191 481 289
rect 541 289 557 323
rect 591 289 637 323
rect 705 317 805 450
rect 541 217 637 289
rect 537 191 637 217
rect 679 217 805 317
rect 855 579 955 627
rect 855 545 896 579
rect 930 545 955 579
rect 855 511 955 545
rect 855 477 896 511
rect 930 477 955 511
rect 855 317 955 477
rect 997 601 1097 627
rect 997 579 1067 601
rect 997 545 1017 579
rect 1051 545 1067 579
rect 1153 559 1253 627
rect 997 511 1067 545
rect 997 477 1017 511
rect 1051 477 1067 511
rect 997 461 1067 477
rect 1109 419 1253 559
rect 1025 389 1253 419
rect 1295 495 1395 627
rect 1569 589 1669 615
rect 1563 567 1669 589
rect 1563 533 1589 567
rect 1623 533 1669 567
rect 1563 499 1669 533
rect 1295 475 1429 495
rect 1295 441 1370 475
rect 1404 441 1429 475
rect 1563 465 1589 499
rect 1623 465 1669 499
rect 1563 445 1669 465
rect 1725 589 1825 615
rect 1725 567 2034 589
rect 1725 533 1980 567
rect 2014 533 2034 567
rect 1725 499 2034 533
rect 2115 527 2215 553
rect 1725 465 1980 499
rect 2014 465 2034 499
rect 1725 445 2034 465
rect 1295 407 1429 441
rect 1295 395 1370 407
rect 1025 338 1139 389
rect 1323 373 1370 395
rect 1404 373 1429 407
rect 855 217 983 317
rect 679 191 779 217
rect 883 191 983 217
rect 1025 304 1045 338
rect 1079 304 1139 338
rect 1025 270 1139 304
rect 1025 236 1045 270
rect 1079 236 1139 270
rect 1025 216 1139 236
rect 1181 331 1281 347
rect 1181 297 1198 331
rect 1232 297 1281 331
rect 1181 263 1281 297
rect 1181 229 1198 263
rect 1232 229 1281 263
rect 1025 191 1125 216
rect 1181 191 1281 229
rect 1323 217 1429 373
rect 1725 225 1781 445
rect 1823 397 1923 401
rect 2115 397 2215 443
rect 1823 381 2215 397
rect 1823 347 1840 381
rect 1874 347 2215 381
rect 1823 313 2215 347
rect 1823 279 1840 313
rect 1874 297 2215 313
rect 1874 279 1937 297
rect 1823 259 1937 279
rect 2115 275 2215 297
rect 2313 369 2413 443
rect 2313 335 2333 369
rect 2367 335 2413 369
rect 2313 275 2413 335
rect 1323 191 1423 217
rect 1681 199 1781 225
rect 1837 199 1937 259
rect 2115 165 2215 191
rect 83 81 183 107
rect 239 81 339 107
rect 381 81 481 107
rect 537 81 637 107
rect 679 81 779 107
rect 883 81 983 107
rect 1025 81 1125 107
rect 1181 81 1281 107
rect 1323 81 1423 107
rect 1681 89 1781 115
rect 1837 89 1937 115
rect 2313 99 2413 125
<< polycont >>
rect 129 541 163 575
rect 129 473 163 507
rect 397 545 431 579
rect 719 538 753 572
rect 397 477 431 511
rect 607 474 641 508
rect 719 470 753 504
rect 253 384 287 418
rect 253 316 287 350
rect 607 406 641 440
rect 397 357 431 391
rect 397 289 431 323
rect 557 289 591 323
rect 896 545 930 579
rect 896 477 930 511
rect 1017 545 1051 579
rect 1017 477 1051 511
rect 1589 533 1623 567
rect 1370 441 1404 475
rect 1589 465 1623 499
rect 1980 533 2014 567
rect 1980 465 2014 499
rect 1370 373 1404 407
rect 1045 304 1079 338
rect 1045 236 1079 270
rect 1198 297 1232 331
rect 1198 229 1232 263
rect 1840 347 1874 381
rect 1840 279 1874 313
rect 2333 335 2367 369
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2496 831
rect 124 735 314 741
rect 22 686 88 715
rect 22 652 38 686
rect 72 652 88 686
rect 22 623 88 652
rect 124 701 130 735
rect 164 701 202 735
rect 236 701 274 735
rect 308 701 314 735
rect 124 686 314 701
rect 124 652 194 686
rect 228 652 314 686
rect 22 269 56 623
rect 124 619 314 652
rect 381 727 612 761
rect 113 575 179 583
rect 113 541 129 575
rect 163 541 179 575
rect 113 507 179 541
rect 113 473 129 507
rect 163 500 179 507
rect 381 579 431 727
rect 381 545 397 579
rect 381 511 431 545
rect 381 500 397 511
rect 163 477 397 500
rect 163 473 431 477
rect 113 466 431 473
rect 381 461 431 466
rect 467 680 542 691
rect 467 646 492 680
rect 526 646 542 680
rect 467 635 542 646
rect 217 418 303 430
rect 217 384 253 418
rect 287 384 303 418
rect 217 350 303 384
rect 217 316 253 350
rect 287 316 303 350
rect 217 305 303 316
rect 381 391 431 407
rect 381 357 397 391
rect 381 323 431 357
rect 381 289 397 323
rect 381 269 431 289
rect 22 235 431 269
rect 467 253 501 635
rect 578 594 612 727
rect 654 735 844 741
rect 654 701 660 735
rect 694 701 732 735
rect 766 701 804 735
rect 838 701 844 735
rect 1266 735 1456 741
rect 654 686 844 701
rect 654 652 810 686
rect 1092 686 1158 719
rect 1092 652 1108 686
rect 1142 652 1158 686
rect 654 619 844 652
rect 537 560 612 594
rect 697 572 769 583
rect 537 354 571 560
rect 697 538 719 572
rect 753 538 769 572
rect 607 508 657 524
rect 641 474 657 508
rect 607 440 657 474
rect 697 504 769 538
rect 697 470 719 504
rect 753 470 769 504
rect 697 460 769 470
rect 880 579 946 652
rect 1092 619 1158 652
rect 1266 701 1272 735
rect 1306 701 1344 735
rect 1378 701 1416 735
rect 1450 701 1456 735
rect 1664 727 2174 761
rect 1266 686 1456 701
rect 1266 652 1406 686
rect 1440 652 1456 686
rect 1266 619 1456 652
rect 1492 674 1574 707
rect 1492 640 1524 674
rect 1558 640 1574 674
rect 1664 686 1730 727
rect 1664 652 1680 686
rect 1714 652 1730 686
rect 1664 647 1730 652
rect 1894 674 1960 691
rect 1492 623 1574 640
rect 1894 640 1910 674
rect 1944 640 1960 674
rect 1894 623 1960 640
rect 1124 583 1158 619
rect 1492 583 1526 623
rect 1610 583 1858 611
rect 880 545 896 579
rect 930 545 946 579
rect 880 511 946 545
rect 880 477 896 511
rect 930 477 946 511
rect 880 460 946 477
rect 1001 579 1067 583
rect 1001 545 1017 579
rect 1051 545 1067 579
rect 1124 549 1526 583
rect 1001 511 1067 545
rect 1001 477 1017 511
rect 1051 477 1067 511
rect 641 424 657 440
rect 1001 424 1067 477
rect 641 406 1248 424
rect 607 390 1248 406
rect 537 338 1084 354
rect 537 323 1045 338
rect 537 289 557 323
rect 591 304 1045 323
rect 1079 304 1084 338
rect 591 289 1084 304
rect 985 270 1084 289
rect 22 166 88 235
rect 467 219 910 253
rect 22 132 38 166
rect 72 132 88 166
rect 22 103 88 132
rect 124 166 314 199
rect 124 132 194 166
rect 228 132 314 166
rect 124 113 314 132
rect 124 79 130 113
rect 164 79 202 113
rect 236 79 274 113
rect 308 79 314 113
rect 467 166 542 219
rect 467 132 492 166
rect 526 132 542 166
rect 467 99 542 132
rect 650 166 840 183
rect 650 132 790 166
rect 824 132 840 166
rect 650 113 840 132
rect 124 73 314 79
rect 650 79 656 113
rect 690 79 728 113
rect 762 79 800 113
rect 834 79 840 113
rect 650 73 840 79
rect 876 87 910 219
rect 985 236 1045 270
rect 1079 236 1084 270
rect 985 162 1084 236
rect 1182 331 1248 390
rect 1182 297 1198 331
rect 1232 297 1248 331
rect 1182 263 1248 297
rect 1182 229 1198 263
rect 1232 229 1248 263
rect 1182 219 1248 229
rect 1284 183 1318 549
rect 1354 475 1420 504
rect 1354 441 1370 475
rect 1404 441 1420 475
rect 1354 407 1420 441
rect 1354 373 1370 407
rect 1404 373 1420 407
rect 1354 310 1420 373
rect 1492 348 1526 549
rect 1562 577 1858 583
rect 1562 567 1644 577
rect 1562 533 1589 567
rect 1623 533 1644 567
rect 1562 499 1644 533
rect 1562 465 1589 499
rect 1623 465 1644 499
rect 1562 384 1644 465
rect 1824 397 1858 577
rect 1824 381 1874 397
rect 1492 314 1670 348
rect 1120 170 1318 183
rect 1120 136 1136 170
rect 1170 136 1318 170
rect 1120 123 1318 136
rect 1354 235 1600 269
rect 1354 87 1388 235
rect 876 53 1388 87
rect 1424 166 1530 199
rect 1424 132 1434 166
rect 1468 132 1530 166
rect 1424 113 1530 132
rect 1458 79 1496 113
rect 1424 73 1530 79
rect 1566 87 1600 235
rect 1636 182 1670 314
rect 1824 347 1840 381
rect 1824 313 1874 347
rect 1824 279 1840 313
rect 1824 263 1874 279
rect 1910 227 1944 623
rect 1980 567 2030 583
rect 2014 533 2030 567
rect 1980 531 2030 533
rect 1980 502 2104 531
rect 1980 499 2070 502
rect 2014 468 2070 499
rect 2014 465 2104 468
rect 1980 423 2104 465
rect 1636 123 1670 148
rect 1706 207 1944 227
rect 2054 250 2104 423
rect 2054 216 2070 250
rect 1706 193 1998 207
rect 1706 87 1740 193
rect 1910 174 1998 193
rect 2054 183 2104 216
rect 2140 385 2174 727
rect 2210 735 2388 751
rect 2244 701 2249 735
rect 2316 701 2354 735
rect 2210 652 2388 701
rect 2210 618 2249 652
rect 2283 618 2388 652
rect 2210 568 2388 618
rect 2210 534 2249 568
rect 2283 534 2388 568
rect 2210 485 2388 534
rect 2210 451 2249 485
rect 2283 451 2388 485
rect 2210 435 2388 451
rect 2424 731 2474 747
rect 2458 697 2474 731
rect 2424 651 2474 697
rect 2458 617 2474 651
rect 2424 569 2474 617
rect 2458 535 2474 569
rect 2424 489 2474 535
rect 2458 455 2474 489
rect 2140 369 2383 385
rect 2140 335 2333 369
rect 2367 335 2383 369
rect 2140 319 2383 335
rect 1566 53 1740 87
rect 1776 123 1792 157
rect 1826 123 1842 157
rect 1910 140 1948 174
rect 1982 140 1998 174
rect 1910 123 1998 140
rect 1776 87 1842 123
rect 2140 87 2174 319
rect 1776 53 2174 87
rect 2210 267 2388 283
rect 2210 233 2268 267
rect 2302 233 2388 267
rect 2210 167 2388 233
rect 2210 133 2268 167
rect 2302 133 2388 167
rect 2210 113 2388 133
rect 2424 263 2474 455
rect 2458 229 2474 263
rect 2424 171 2474 229
rect 2458 137 2474 171
rect 2424 121 2474 137
rect 2244 79 2282 113
rect 2316 79 2354 113
rect 2210 73 2388 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2496 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 130 701 164 735
rect 202 701 236 735
rect 274 701 308 735
rect 660 701 694 735
rect 732 701 766 735
rect 804 701 838 735
rect 1272 701 1306 735
rect 1344 701 1378 735
rect 1416 701 1450 735
rect 130 79 164 113
rect 202 79 236 113
rect 274 79 308 113
rect 656 79 690 113
rect 728 79 762 113
rect 800 79 834 113
rect 1424 79 1458 113
rect 1496 79 1530 113
rect 2210 701 2244 735
rect 2282 701 2283 735
rect 2283 701 2316 735
rect 2354 701 2388 735
rect 2210 79 2244 113
rect 2282 79 2316 113
rect 2354 79 2388 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
<< metal1 >>
rect 0 831 2496 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2496 831
rect 0 791 2496 797
rect 0 735 2496 763
rect 0 701 130 735
rect 164 701 202 735
rect 236 701 274 735
rect 308 701 660 735
rect 694 701 732 735
rect 766 701 804 735
rect 838 701 1272 735
rect 1306 701 1344 735
rect 1378 701 1416 735
rect 1450 701 2210 735
rect 2244 701 2282 735
rect 2316 701 2354 735
rect 2388 701 2496 735
rect 0 689 2496 701
rect 0 113 2496 125
rect 0 79 130 113
rect 164 79 202 113
rect 236 79 274 113
rect 308 79 656 113
rect 690 79 728 113
rect 762 79 800 113
rect 834 79 1424 113
rect 1458 79 1496 113
rect 1530 79 2210 113
rect 2244 79 2282 113
rect 2316 79 2354 113
rect 2388 79 2496 113
rect 0 51 2496 79
rect 0 17 2496 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2496 17
rect 0 -23 2496 -17
<< labels >>
flabel comment s 523 410 523 410 0 FreeSans 200 0 0 0 no_jumper_check
rlabel comment s 0 0 0 0 4 mux4_1
flabel metal1 s 0 51 2496 125 0 FreeSans 340 0 0 0 VGND
port 7 nsew ground bidirectional
flabel metal1 s 0 0 2496 23 0 FreeSans 340 0 0 0 VNB
port 8 nsew ground bidirectional
flabel metal1 s 0 689 2496 763 0 FreeSans 340 0 0 0 VPWR
port 10 nsew power bidirectional
flabel metal1 s 0 791 2496 814 0 FreeSans 340 0 0 0 VPB
port 9 nsew power bidirectional
flabel locali s 1375 316 1409 350 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
flabel locali s 1375 390 1409 424 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
flabel locali s 1375 464 1409 498 0 FreeSans 340 0 0 0 A0
port 1 nsew signal input
flabel locali s 991 168 1025 202 0 FreeSans 340 0 0 0 S0
port 5 nsew signal input
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 S0
port 5 nsew signal input
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 S0
port 5 nsew signal input
flabel locali s 895 464 929 498 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 895 538 929 572 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 895 612 929 646 0 FreeSans 340 0 0 0 A1
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A2
port 3 nsew signal input
flabel locali s 223 390 257 424 0 FreeSans 340 0 0 0 A2
port 3 nsew signal input
flabel locali s 703 464 737 498 0 FreeSans 340 0 0 0 A3
port 4 nsew signal input
flabel locali s 703 538 737 572 0 FreeSans 340 0 0 0 A3
port 4 nsew signal input
flabel locali s 2431 168 2465 202 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 2431 242 2465 276 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 2431 316 2465 350 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 2431 390 2465 424 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 2431 464 2465 498 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 2431 538 2465 572 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 2431 612 2465 646 0 FreeSans 340 0 0 0 X
port 11 nsew signal output
flabel locali s 1567 390 1601 424 0 FreeSans 340 0 0 0 S1
port 6 nsew signal input
flabel locali s 1567 464 1601 498 0 FreeSans 340 0 0 0 S1
port 6 nsew signal input
flabel locali s 1567 538 1601 572 0 FreeSans 340 0 0 0 S1
port 6 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 2496 814
string GDS_END 236664
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 211614
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
