magic
tech sky130B
magscale 1 2
timestamp 1707688321
use sky130_fd_io__gnd2gnd_strap  sky130_fd_io__gnd2gnd_strap_0
timestamp 1707688321
transform 1 0 0 0 1 0
box 61 139 62 140
<< properties >>
string GDS_END 30713020
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 30712836
<< end >>
