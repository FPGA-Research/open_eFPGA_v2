magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -91 498 247 593
rect 651 66 817 798
rect 3093 1232 3211 1904
rect 2585 1138 3211 1232
rect 3093 466 3211 1138
<< pwell >>
rect 227 1451 313 2050
rect 2477 82 2563 2195
<< psubdiff >>
rect 2503 2145 2537 2169
rect 2503 2076 2537 2111
rect 253 2000 287 2024
rect 2503 2007 2537 2042
rect 253 1923 287 1966
rect 253 1846 287 1889
rect 253 1769 287 1812
rect 253 1691 287 1735
rect 253 1613 287 1657
rect 253 1535 287 1579
rect 253 1477 287 1501
rect 2503 1938 2537 1973
rect 2503 1869 2537 1904
rect 2503 1800 2537 1835
rect 2503 1731 2537 1766
rect 2503 1662 2537 1697
rect 2503 1594 2537 1628
rect 2503 1526 2537 1560
rect 2503 1458 2537 1492
rect 2503 1390 2537 1424
rect 2503 1322 2537 1356
rect 2503 1254 2537 1288
rect 2503 1186 2537 1220
rect 2503 1118 2537 1152
rect 2503 1050 2537 1084
rect 2503 982 2537 1016
rect 2503 914 2537 948
rect 2503 846 2537 880
rect 2503 778 2537 812
rect 2503 710 2537 744
rect 2503 642 2537 676
rect 2503 574 2537 608
rect 2503 506 2537 540
rect 2503 438 2537 472
rect 2503 370 2537 404
rect 2503 302 2537 336
rect 2503 234 2537 268
rect 2503 166 2537 200
rect 2503 108 2537 132
<< nsubdiff >>
rect 3130 1819 3166 1865
rect 3130 1785 3131 1819
rect 3165 1785 3166 1819
rect 3130 1751 3166 1785
rect 3130 1717 3131 1751
rect 3165 1717 3166 1751
rect 3130 1683 3166 1717
rect 3130 1649 3131 1683
rect 3165 1649 3166 1683
rect 3130 1615 3166 1649
rect 3130 1581 3131 1615
rect 3165 1581 3166 1615
rect 3130 1547 3166 1581
rect 3130 1513 3131 1547
rect 3165 1513 3166 1547
rect 3130 1472 3166 1513
rect 3130 1438 3131 1472
rect 3165 1438 3166 1472
rect 3130 1404 3166 1438
rect 3130 1370 3131 1404
rect 3165 1370 3166 1404
rect 3130 1336 3166 1370
rect 3130 1302 3131 1336
rect 3165 1302 3166 1336
rect 3130 1268 3166 1302
rect 3130 1234 3131 1268
rect 3165 1234 3166 1268
rect 3130 1200 3166 1234
rect 3130 1166 3131 1200
rect 3165 1166 3166 1200
rect 3130 1132 3166 1166
rect 3130 1098 3131 1132
rect 3165 1098 3166 1132
rect 3130 1064 3166 1098
rect 3130 1030 3131 1064
rect 3165 1030 3166 1064
rect 3130 996 3166 1030
rect 3130 962 3131 996
rect 3165 962 3166 996
rect 3130 921 3166 962
rect 3130 887 3131 921
rect 3165 887 3166 921
rect 3130 853 3166 887
rect 3130 819 3131 853
rect 3165 819 3166 853
rect 3130 785 3166 819
rect 3130 751 3131 785
rect 3165 751 3166 785
rect 3130 717 3166 751
rect 3130 683 3131 717
rect 3165 683 3166 717
rect 3130 649 3166 683
rect 3130 615 3131 649
rect 3165 615 3166 649
rect 3130 581 3166 615
rect 3130 547 3131 581
rect 3165 547 3166 581
rect 3130 511 3166 547
<< mvnsubdiff >>
rect 717 708 751 732
rect 717 634 751 674
rect 717 560 751 600
rect 717 486 751 526
rect 717 412 751 452
rect 717 338 751 378
rect 717 264 751 304
rect 717 190 751 230
rect 717 132 751 156
<< psubdiffcont >>
rect 2503 2111 2537 2145
rect 2503 2042 2537 2076
rect 253 1966 287 2000
rect 253 1889 287 1923
rect 253 1812 287 1846
rect 253 1735 287 1769
rect 253 1657 287 1691
rect 253 1579 287 1613
rect 253 1501 287 1535
rect 2503 1973 2537 2007
rect 2503 1904 2537 1938
rect 2503 1835 2537 1869
rect 2503 1766 2537 1800
rect 2503 1697 2537 1731
rect 2503 1628 2537 1662
rect 2503 1560 2537 1594
rect 2503 1492 2537 1526
rect 2503 1424 2537 1458
rect 2503 1356 2537 1390
rect 2503 1288 2537 1322
rect 2503 1220 2537 1254
rect 2503 1152 2537 1186
rect 2503 1084 2537 1118
rect 2503 1016 2537 1050
rect 2503 948 2537 982
rect 2503 880 2537 914
rect 2503 812 2537 846
rect 2503 744 2537 778
rect 2503 676 2537 710
rect 2503 608 2537 642
rect 2503 540 2537 574
rect 2503 472 2537 506
rect 2503 404 2537 438
rect 2503 336 2537 370
rect 2503 268 2537 302
rect 2503 200 2537 234
rect 2503 132 2537 166
<< nsubdiffcont >>
rect 3131 1785 3165 1819
rect 3131 1717 3165 1751
rect 3131 1649 3165 1683
rect 3131 1581 3165 1615
rect 3131 1513 3165 1547
rect 3131 1438 3165 1472
rect 3131 1370 3165 1404
rect 3131 1302 3165 1336
rect 3131 1234 3165 1268
rect 3131 1166 3165 1200
rect 3131 1098 3165 1132
rect 3131 1030 3165 1064
rect 3131 962 3165 996
rect 3131 887 3165 921
rect 3131 819 3165 853
rect 3131 751 3165 785
rect 3131 683 3165 717
rect 3131 615 3165 649
rect 3131 547 3165 581
<< mvnsubdiffcont >>
rect 717 674 751 708
rect 717 600 751 634
rect 717 526 751 560
rect 717 452 751 486
rect 717 378 751 412
rect 717 304 751 338
rect 717 230 751 264
rect 717 156 751 190
<< poly >>
rect 1311 2278 1720 2294
rect 1311 2244 1329 2278
rect 1363 2244 1397 2278
rect 1431 2244 1465 2278
rect 1499 2244 1533 2278
rect 1567 2244 1601 2278
rect 1635 2244 1669 2278
rect 1703 2244 1720 2278
rect 1311 2228 1720 2244
rect 1900 2278 2080 2294
rect 1900 2244 1939 2278
rect 1973 2244 2007 2278
rect 2041 2244 2080 2278
rect 1900 2228 2080 2244
rect 2251 2278 2385 2294
rect 2251 2244 2267 2278
rect 2301 2244 2335 2278
rect 2369 2244 2385 2278
rect 2251 2228 2385 2244
rect 420 2158 554 2174
rect 420 2124 436 2158
rect 470 2124 504 2158
rect 538 2124 554 2158
rect 420 2050 554 2124
rect 812 2106 946 2122
rect 812 2072 828 2106
rect 862 2072 896 2106
rect 930 2072 946 2106
rect 812 2050 946 2072
rect 1002 2106 1136 2122
rect 1002 2072 1018 2106
rect 1052 2072 1086 2106
rect 1120 2072 1136 2106
rect 1002 2050 1136 2072
rect 610 1794 646 1798
rect 610 1778 676 1794
rect 610 1744 626 1778
rect 660 1744 676 1778
rect 323 1710 554 1726
rect 323 1676 339 1710
rect 373 1676 407 1710
rect 441 1676 554 1710
rect 323 1660 554 1676
rect 518 1650 554 1660
rect 610 1710 676 1744
rect 610 1676 626 1710
rect 660 1676 676 1710
rect 610 1660 676 1676
rect 610 1650 646 1660
rect 1900 1182 2080 1976
rect 2260 1402 2290 1976
rect 2346 1402 2376 1976
rect 2590 1950 2724 1966
rect 2590 1916 2606 1950
rect 2640 1916 2674 1950
rect 2708 1916 2724 1950
rect 2590 1900 2724 1916
rect 2766 1950 3022 1966
rect 2766 1916 2782 1950
rect 2816 1916 2850 1950
rect 2884 1916 3022 1950
rect 2590 1894 2710 1900
rect 2766 1894 3022 1916
rect 1900 1148 1939 1182
rect 1973 1148 2007 1182
rect 2041 1148 2080 1182
rect 28 1030 206 1056
rect 28 928 67 1030
rect 169 928 206 1030
rect 28 885 206 928
rect 262 1034 414 1056
rect 262 932 278 1034
rect 380 932 414 1034
rect 262 758 414 932
rect 826 1040 946 1056
rect 826 1006 869 1040
rect 903 1006 946 1040
rect 826 972 946 1006
rect 826 938 869 972
rect 903 938 946 972
rect 826 922 946 938
rect 1002 1040 1122 1056
rect 1002 1006 1018 1040
rect 1052 1006 1122 1040
rect 1002 972 1122 1006
rect 1002 938 1018 972
rect 1052 938 1122 972
rect 1002 922 1122 938
rect 1304 353 1484 882
rect 1540 353 1720 882
rect 28 106 128 206
rect 28 14 414 106
rect 470 80 603 106
rect 1900 102 2080 1148
rect 2569 1184 2710 1200
rect 2569 1150 2585 1184
rect 2619 1150 2653 1184
rect 2687 1150 2710 1184
rect 2569 1128 2710 1150
rect 2766 1128 3022 1242
rect 2260 274 2290 882
rect 2346 274 2376 882
rect 2766 454 3036 476
rect 2766 420 2782 454
rect 2816 420 2850 454
rect 2884 420 2918 454
rect 2952 420 2986 454
rect 3020 420 3036 454
rect 2766 404 3036 420
rect 470 64 604 80
rect 470 30 486 64
rect 520 30 554 64
rect 588 30 604 64
rect 1304 36 2080 102
rect 2251 86 2385 102
rect 2251 52 2267 86
rect 2301 52 2335 86
rect 2369 52 2385 86
rect 2251 36 2385 52
rect 470 14 604 30
<< polycont >>
rect 1329 2244 1363 2278
rect 1397 2244 1431 2278
rect 1465 2244 1499 2278
rect 1533 2244 1567 2278
rect 1601 2244 1635 2278
rect 1669 2244 1703 2278
rect 1939 2244 1973 2278
rect 2007 2244 2041 2278
rect 2267 2244 2301 2278
rect 2335 2244 2369 2278
rect 436 2124 470 2158
rect 504 2124 538 2158
rect 828 2072 862 2106
rect 896 2072 930 2106
rect 1018 2072 1052 2106
rect 1086 2072 1120 2106
rect 626 1744 660 1778
rect 339 1676 373 1710
rect 407 1676 441 1710
rect 626 1676 660 1710
rect 2606 1916 2640 1950
rect 2674 1916 2708 1950
rect 2782 1916 2816 1950
rect 2850 1916 2884 1950
rect 1939 1148 1973 1182
rect 2007 1148 2041 1182
rect 67 928 169 1030
rect 278 932 380 1034
rect 869 1006 903 1040
rect 869 938 903 972
rect 1018 1006 1052 1040
rect 1018 938 1052 972
rect 2585 1150 2619 1184
rect 2653 1150 2687 1184
rect 2782 420 2816 454
rect 2850 420 2884 454
rect 2918 420 2952 454
rect 2986 420 3020 454
rect 486 30 520 64
rect 554 30 588 64
rect 2267 52 2301 86
rect 2335 52 2369 86
<< locali >>
rect 420 2280 432 2314
rect 466 2280 504 2314
rect 538 2280 554 2314
rect 420 2158 554 2280
rect 420 2124 436 2158
rect 470 2124 504 2158
rect 538 2124 554 2158
rect 812 2106 946 2379
rect 1096 2362 1136 2379
rect 381 2056 599 2090
rect 812 2072 828 2106
rect 862 2072 896 2106
rect 930 2072 946 2106
rect 1002 2106 1136 2362
rect 2251 2354 2279 2388
rect 2313 2354 2351 2388
rect 2251 2278 2385 2354
rect 1313 2244 1329 2278
rect 1363 2244 1397 2278
rect 1431 2244 1465 2278
rect 1499 2244 1533 2278
rect 1567 2244 1601 2278
rect 1635 2244 1669 2278
rect 1703 2244 1719 2278
rect 1923 2244 1939 2278
rect 1973 2244 2007 2278
rect 2041 2244 2057 2278
rect 2251 2244 2267 2278
rect 2301 2244 2335 2278
rect 2369 2244 2385 2278
rect 1002 2072 1018 2106
rect 1052 2072 1086 2106
rect 1120 2072 1136 2106
rect 253 2000 287 2024
rect 253 1923 287 1966
rect 253 1849 287 1889
rect 253 1777 287 1812
rect 253 1705 287 1735
rect 381 1735 415 2056
rect 339 1710 381 1726
rect 475 1849 515 2022
rect 565 2018 599 2056
rect 684 1849 747 2022
rect 475 1815 481 1849
rect 675 1815 713 1849
rect 475 1777 515 1815
rect 475 1743 481 1777
rect 610 1751 626 1778
rect 660 1751 676 1778
rect 415 1710 441 1726
rect 373 1701 381 1710
rect 373 1676 407 1701
rect 339 1663 441 1676
rect 339 1660 381 1663
rect 253 1633 287 1657
rect 415 1660 441 1663
rect 253 1561 287 1579
rect 253 1443 287 1501
rect 475 1444 515 1743
rect 604 1744 626 1751
rect 604 1717 642 1744
rect 610 1710 676 1717
rect 610 1676 626 1710
rect 660 1676 676 1710
rect 710 1642 747 1815
rect 565 1523 599 1561
rect 473 1410 515 1444
rect 657 1443 747 1642
rect 815 1489 853 1523
rect 323 1403 515 1410
rect 323 1369 409 1403
rect 443 1369 481 1403
rect 515 1369 641 1386
rect 323 1331 641 1369
rect 323 1320 494 1331
rect 482 1297 494 1320
rect 528 1297 566 1331
rect 600 1297 641 1331
rect 217 1259 251 1265
rect 414 1151 448 1286
rect 482 1265 641 1297
rect 781 1212 815 1486
rect 957 1443 991 1486
rect 957 1371 991 1409
rect 957 1299 991 1337
rect 957 1154 991 1265
rect 1133 1256 1300 2028
rect 1553 1489 1591 1523
rect 1133 1212 1167 1256
rect 1422 1180 1456 1266
rect 1731 1256 1889 2206
rect 217 1103 251 1146
rect 413 1105 448 1151
rect 1259 1140 1765 1180
rect 75 1064 113 1098
rect 278 1034 380 1050
rect 51 928 67 1030
rect 169 1018 185 1030
rect 169 928 185 984
rect -17 436 17 661
rect 51 436 105 928
rect 308 910 346 932
rect 274 894 380 910
rect 139 857 380 894
rect 139 829 173 857
rect 414 823 448 1105
rect 269 789 448 823
rect 516 1058 554 1092
rect 482 796 588 1058
rect 781 944 815 1116
rect 1259 1106 1293 1140
rect 1731 1106 1765 1140
rect 743 910 781 944
rect 853 1018 869 1040
rect 903 1018 919 1040
rect 903 1006 925 1018
rect 887 984 925 1006
rect 1002 1006 1018 1040
rect 1052 1006 1068 1040
rect 1133 1018 1167 1092
rect 853 972 919 984
rect 853 938 869 972
rect 903 938 919 972
rect 1002 972 1068 1006
rect 1137 984 1175 1018
rect 1002 944 1018 972
rect 1052 944 1068 972
rect 1495 950 1529 988
rect 1052 938 1074 944
rect 1036 910 1074 938
rect 269 736 303 789
rect 482 762 615 796
rect 581 736 615 762
rect 717 708 751 732
rect 717 634 751 674
rect 717 560 751 600
rect 717 486 751 526
rect -17 222 17 260
rect -17 150 17 188
rect 51 64 173 436
rect 717 412 751 452
rect 717 338 751 378
rect 1259 306 1293 904
rect 717 294 751 304
rect 1495 296 1529 904
rect 425 222 459 260
rect 425 150 459 188
rect 1731 286 1765 904
rect 1855 260 1889 1256
rect 1923 2090 2057 2244
rect 1923 1912 1937 2090
rect 2043 1912 2057 2090
rect 2503 2145 2537 2169
rect 2503 2076 2537 2111
rect 2503 2007 2537 2042
rect 1923 1182 2057 1912
rect 1923 1148 1939 1182
rect 1973 1148 2007 1182
rect 2041 1148 2057 1182
rect 717 222 751 230
rect 717 150 751 156
rect 1923 90 2057 1148
rect 2091 1595 2125 1998
rect 2091 1523 2125 1561
rect 2091 283 2125 1489
rect 2215 1443 2249 1998
rect 2215 1371 2249 1409
rect 2215 1299 2249 1337
rect 2301 1595 2335 1998
rect 2301 1523 2335 1561
rect 2301 1317 2335 1489
rect 2387 1443 2421 1998
rect 2387 1371 2421 1409
rect 2387 1299 2421 1337
rect 2503 1938 2537 1973
rect 2934 2022 2968 2060
rect 2934 1950 2968 1988
rect 2503 1869 2537 1904
rect 2590 1916 2606 1950
rect 2640 1916 2674 1950
rect 2708 1916 2724 1950
rect 2766 1916 2782 1950
rect 2816 1916 2850 1950
rect 2884 1916 2900 1950
rect 2590 1874 2724 1916
rect 2590 1840 2618 1874
rect 2652 1840 2690 1874
rect 2503 1800 2537 1835
rect 2503 1731 2537 1766
rect 2503 1662 2537 1697
rect 2585 1671 2663 1806
rect 2789 1755 2843 1916
rect 2934 1844 2968 1916
rect 2877 1810 2968 1844
rect 3131 1819 3165 1864
rect 2877 1806 2911 1810
rect 2789 1721 2799 1755
rect 2833 1721 2843 1755
rect 2789 1683 2843 1721
rect 2615 1637 2653 1671
rect 2789 1649 2799 1683
rect 2833 1649 2843 1683
rect 2503 1594 2537 1628
rect 2503 1526 2537 1560
rect 2503 1458 2537 1492
rect 2503 1390 2537 1409
rect 2503 1322 2537 1337
rect 2503 1254 2537 1265
rect 2215 1106 2249 1247
rect 2387 1106 2421 1237
rect 2503 1186 2537 1220
rect 2503 1118 2537 1152
rect 2585 1200 2663 1637
rect 2721 1523 2755 1561
rect 2585 1184 2687 1200
rect 2619 1150 2653 1184
rect 2585 1134 2687 1150
rect 2503 1050 2537 1084
rect 2301 950 2335 988
rect 2721 1040 2755 1264
rect 2503 982 2537 1016
rect 2503 914 2537 948
rect 2721 950 2755 988
rect 2215 276 2249 904
rect 2301 276 2335 904
rect 2387 276 2421 904
rect 2503 846 2537 880
rect 2629 864 2663 902
rect 2503 778 2537 812
rect 2503 710 2537 744
rect 2503 642 2537 676
rect 2503 574 2537 608
rect 2503 506 2537 540
rect 2503 452 2537 472
rect 2503 380 2537 404
rect 2503 302 2537 336
rect 2503 234 2537 268
rect 2503 166 2537 200
rect 2503 108 2537 132
rect 51 30 486 64
rect 520 30 554 64
rect 588 30 604 64
rect 1312 26 2058 90
rect 2251 52 2267 86
rect 2301 52 2335 86
rect 2369 74 2385 86
rect 2629 74 2663 565
rect 2789 454 2843 1649
rect 2945 1721 2956 1755
rect 2990 1721 2999 1755
rect 2945 1683 2999 1721
rect 2945 1649 2956 1683
rect 2990 1649 2999 1683
rect 2877 1039 2911 1264
rect 2877 873 2911 911
rect 2945 454 2999 1649
rect 3131 1751 3165 1785
rect 3131 1683 3165 1717
rect 3131 1615 3165 1649
rect 3033 1523 3067 1561
rect 3131 1547 3165 1561
rect 3131 1472 3165 1489
rect 3131 1404 3165 1438
rect 3131 1336 3165 1370
rect 3131 1268 3165 1302
rect 3033 1039 3067 1264
rect 3131 1200 3165 1234
rect 3131 1132 3165 1166
rect 3131 1083 3165 1098
rect 3033 950 3067 988
rect 3131 1011 3165 1030
rect 3131 939 3165 962
rect 3131 867 3165 887
rect 3131 785 3165 819
rect 3131 717 3165 751
rect 3131 649 3165 683
rect 3131 581 3165 615
rect 3131 512 3165 547
rect 2766 420 2782 454
rect 2816 420 2850 454
rect 2884 420 2918 454
rect 2952 420 2986 454
rect 3020 420 3036 454
rect 2369 52 2663 74
rect 2251 40 2663 52
<< viali >>
rect 432 2280 466 2314
rect 504 2280 538 2314
rect 2279 2354 2313 2388
rect 2351 2354 2385 2388
rect 253 1846 287 1849
rect 253 1815 287 1846
rect 253 1769 287 1777
rect 253 1743 287 1769
rect 253 1691 287 1705
rect 253 1671 287 1691
rect 381 1710 415 1735
rect 481 1815 515 1849
rect 641 1815 675 1849
rect 713 1815 747 1849
rect 481 1743 515 1777
rect 381 1701 407 1710
rect 407 1701 415 1710
rect 253 1613 287 1633
rect 381 1629 415 1663
rect 253 1599 287 1613
rect 253 1535 287 1561
rect 253 1527 287 1535
rect 570 1717 604 1751
rect 642 1744 660 1751
rect 660 1744 676 1751
rect 642 1717 676 1744
rect 565 1561 599 1595
rect 565 1489 599 1523
rect 217 1265 323 1443
rect 781 1489 815 1523
rect 853 1489 887 1523
rect 409 1369 443 1403
rect 481 1369 515 1403
rect 494 1297 528 1331
rect 566 1297 600 1331
rect 641 1265 747 1443
rect 957 1409 991 1443
rect 957 1337 991 1371
rect 957 1265 991 1299
rect 1519 1489 1553 1523
rect 1591 1489 1625 1523
rect 41 1064 75 1098
rect 113 1064 147 1098
rect 88 984 122 1018
rect 160 984 169 1018
rect 169 984 194 1018
rect 274 932 278 944
rect 278 932 308 944
rect 346 932 380 944
rect 274 910 308 932
rect 346 910 380 932
rect 482 1058 516 1092
rect 554 1058 588 1092
rect 709 910 743 944
rect 781 910 815 944
rect 853 1006 869 1018
rect 869 1006 887 1018
rect 853 984 887 1006
rect 925 984 959 1018
rect 1103 984 1137 1018
rect 1175 984 1209 1018
rect 1495 988 1529 1022
rect 1002 938 1018 944
rect 1018 938 1036 944
rect 1002 910 1036 938
rect 1074 910 1108 944
rect 1495 916 1529 950
rect -17 260 17 294
rect -17 188 17 222
rect -17 116 17 150
rect 959 346 1137 452
rect 425 260 459 294
rect 425 188 459 222
rect 425 116 459 150
rect 717 264 751 294
rect 717 260 751 264
rect 1937 1912 2043 2090
rect 717 190 751 222
rect 717 188 751 190
rect 717 116 751 150
rect 2091 1561 2125 1595
rect 2091 1489 2125 1523
rect 2215 1409 2249 1443
rect 2215 1337 2249 1371
rect 2301 1561 2335 1595
rect 2301 1489 2335 1523
rect 2387 1409 2421 1443
rect 2387 1337 2421 1371
rect 2215 1265 2249 1299
rect 2387 1265 2421 1299
rect 2934 2060 2968 2094
rect 2934 1988 2968 2022
rect 2934 1916 2968 1950
rect 2618 1840 2652 1874
rect 2690 1840 2724 1874
rect 2799 1721 2833 1755
rect 2581 1637 2615 1671
rect 2653 1637 2687 1671
rect 2799 1649 2833 1683
rect 2503 1424 2537 1443
rect 2503 1409 2537 1424
rect 2503 1356 2537 1371
rect 2503 1337 2537 1356
rect 2503 1288 2537 1299
rect 2503 1265 2537 1288
rect 2721 1561 2755 1595
rect 2721 1489 2755 1523
rect 2301 988 2335 1022
rect 2301 916 2335 950
rect 2721 988 2755 1022
rect 2629 902 2663 936
rect 2721 916 2755 950
rect 2629 830 2663 864
rect 2503 438 2537 452
rect 2503 418 2537 438
rect 2503 370 2537 380
rect 2503 346 2537 370
rect 2956 1721 2990 1755
rect 2956 1649 2990 1683
rect 2877 911 2911 945
rect 2877 839 2911 873
rect 3033 1561 3067 1595
rect 3033 1489 3067 1523
rect 3131 1581 3165 1595
rect 3131 1561 3165 1581
rect 3131 1513 3165 1523
rect 3131 1489 3165 1513
rect 3131 1064 3165 1083
rect 3131 1049 3165 1064
rect 3033 988 3067 1022
rect 3033 916 3067 950
rect 3131 996 3165 1011
rect 3131 977 3165 996
rect 3131 921 3165 939
rect 3131 905 3165 921
rect 3131 853 3165 867
rect 3131 833 3165 853
<< metal1 >>
rect 2267 2388 2424 2400
rect 2267 2354 2279 2388
rect 2313 2354 2351 2388
rect 2385 2354 2424 2388
rect 2267 2348 2424 2354
rect 2476 2348 2488 2400
rect 2540 2348 2546 2400
tri 2627 2320 2652 2345 se
rect 2652 2320 2658 2390
rect 420 2314 2658 2320
rect 420 2280 432 2314
rect 466 2280 504 2314
rect 538 2280 2658 2314
rect 420 2274 2658 2280
rect 2774 2274 2780 2390
rect 10 2194 3122 2246
rect 3174 2194 3312 2246
rect 10 2182 3312 2194
rect 10 2130 3122 2182
rect 3174 2130 3312 2182
rect 10 2118 3312 2130
rect 10 2094 3122 2118
rect 10 2090 2934 2094
rect 10 1912 1937 2090
rect 2043 2060 2934 2090
rect 2968 2066 3122 2094
rect 3174 2066 3312 2118
rect 2968 2060 3312 2066
rect 2043 2054 3312 2060
rect 2043 2022 3122 2054
rect 2043 1988 2934 2022
rect 2968 2002 3122 2022
rect 3174 2002 3312 2054
rect 2968 1990 3312 2002
rect 2968 1988 3122 1990
rect 2043 1950 3122 1988
rect 2043 1923 2934 1950
rect 2043 1916 2543 1923
tri 2543 1916 2550 1923 nw
tri 2780 1916 2787 1923 ne
rect 2787 1916 2934 1923
rect 2968 1938 3122 1950
rect 3174 1938 3312 1990
rect 2968 1916 3312 1938
rect 2043 1912 2537 1916
rect 10 1910 2537 1912
tri 2537 1910 2543 1916 nw
tri 2787 1910 2793 1916 ne
rect 2793 1910 3312 1916
rect 10 1906 2533 1910
tri 2533 1906 2537 1910 nw
tri 2793 1906 2797 1910 ne
rect 2797 1906 3312 1910
rect 10 1898 2525 1906
tri 2525 1898 2533 1906 nw
tri 2797 1898 2805 1906 ne
rect 2805 1898 3312 1906
rect 2606 1874 2658 1880
rect 2710 1874 2722 1880
rect 247 1849 293 1861
rect 247 1815 253 1849
rect 287 1815 293 1849
rect 247 1777 293 1815
rect 247 1743 253 1777
rect 287 1743 293 1777
rect 247 1705 293 1743
rect 475 1849 753 1861
rect 475 1815 481 1849
rect 515 1815 641 1849
rect 675 1815 713 1849
rect 747 1815 753 1849
rect 2606 1840 2618 1874
rect 2652 1840 2658 1874
rect 2606 1828 2658 1840
rect 2710 1828 2722 1840
rect 2774 1828 2780 1880
rect 475 1803 753 1815
rect 475 1777 521 1803
tri 521 1778 546 1803 nw
rect 475 1743 481 1777
rect 515 1743 521 1777
rect 247 1671 253 1705
rect 287 1671 293 1705
rect 247 1633 293 1671
rect 247 1599 253 1633
rect 287 1599 293 1633
rect 369 1735 427 1741
rect 369 1701 381 1735
rect 415 1701 427 1735
rect 475 1731 521 1743
rect 564 1755 3002 1763
rect 564 1751 2799 1755
rect 564 1717 570 1751
rect 604 1717 642 1751
rect 676 1721 2799 1751
rect 2833 1721 2956 1755
rect 2990 1721 3002 1755
rect 676 1717 3002 1721
rect 564 1705 3002 1717
tri 2762 1702 2765 1705 ne
rect 2765 1702 2848 1705
rect 369 1683 427 1701
tri 427 1683 446 1702 sw
tri 2765 1683 2784 1702 ne
rect 2784 1683 2848 1702
tri 2848 1683 2870 1705 nw
tri 2919 1683 2941 1705 ne
rect 2941 1683 3002 1705
rect 369 1677 446 1683
tri 446 1677 452 1683 sw
tri 2784 1680 2787 1683 ne
rect 369 1671 2699 1677
rect 369 1663 2395 1671
rect 369 1629 381 1663
rect 415 1630 2395 1663
rect 415 1629 427 1630
rect 369 1623 427 1629
tri 427 1623 434 1630 nw
tri 2378 1623 2385 1630 ne
rect 2385 1623 2395 1630
tri 2385 1613 2395 1623 ne
rect 2447 1619 2459 1671
rect 2511 1637 2581 1671
rect 2615 1637 2653 1671
rect 2687 1637 2699 1671
rect 2787 1649 2799 1683
rect 2833 1649 2845 1683
tri 2845 1680 2848 1683 nw
tri 2941 1680 2944 1683 ne
rect 2787 1643 2845 1649
rect 2944 1649 2956 1683
rect 2990 1649 3002 1683
rect 2944 1643 3002 1649
rect 2511 1630 2699 1637
rect 2395 1613 2511 1619
tri 2511 1613 2528 1630 nw
rect 247 1561 293 1599
rect 553 1600 698 1601
rect 553 1595 640 1600
tri 293 1561 316 1584 sw
rect 553 1561 565 1595
rect 599 1561 640 1595
rect 247 1527 253 1561
rect 287 1527 316 1561
rect 247 1523 316 1527
tri 316 1523 354 1561 sw
rect 553 1548 640 1561
rect 692 1548 698 1600
rect 553 1536 698 1548
rect 553 1523 640 1536
rect 247 1515 354 1523
tri 354 1515 362 1523 sw
rect 247 1489 362 1515
tri 362 1489 388 1515 sw
rect 553 1489 565 1523
rect 599 1489 640 1523
rect 247 1483 388 1489
tri 388 1483 394 1489 sw
rect 553 1484 640 1489
rect 692 1484 698 1536
rect 2079 1595 2347 1601
rect 2079 1561 2091 1595
rect 2125 1561 2301 1595
rect 2335 1561 2347 1595
rect 553 1483 698 1484
rect 769 1523 1637 1529
rect 769 1489 781 1523
rect 815 1489 853 1523
rect 887 1489 1519 1523
rect 1553 1489 1591 1523
rect 1625 1489 1637 1523
rect 769 1483 1637 1489
rect 2079 1523 2347 1561
rect 2079 1489 2091 1523
rect 2125 1489 2301 1523
rect 2335 1489 2347 1523
rect 2079 1483 2347 1489
rect 2709 1595 3079 1601
rect 2709 1561 2721 1595
rect 2755 1561 3033 1595
rect 3067 1561 3079 1595
rect 2709 1523 3079 1561
rect 2709 1489 2721 1523
rect 2755 1489 3033 1523
rect 3067 1489 3079 1523
rect 2709 1483 3079 1489
rect 3116 1549 3122 1601
rect 3174 1549 3180 1601
rect 3116 1537 3180 1549
rect 3116 1485 3122 1537
rect 3174 1485 3180 1537
rect 3116 1483 3180 1485
rect 247 1455 394 1483
tri 394 1455 422 1483 sw
rect -96 1443 3312 1455
rect -96 1265 217 1443
rect 323 1403 641 1443
rect 323 1369 409 1403
rect 443 1369 481 1403
rect 515 1369 641 1403
rect 323 1331 641 1369
rect 323 1297 494 1331
rect 528 1297 566 1331
rect 600 1297 641 1331
rect 323 1265 641 1297
rect 747 1409 957 1443
rect 991 1409 2215 1443
rect 2249 1409 2387 1443
rect 2421 1409 2503 1443
rect 2537 1409 3312 1443
rect 747 1371 3312 1409
rect 747 1337 957 1371
rect 991 1337 2215 1371
rect 2249 1337 2387 1371
rect 2421 1337 2503 1371
rect 2537 1337 3312 1371
rect 747 1299 3312 1337
rect 747 1265 957 1299
rect 991 1265 2215 1299
rect 2249 1265 2387 1299
rect 2421 1265 2503 1299
rect 2537 1265 3312 1299
rect -96 1253 3312 1265
rect 29 1098 600 1104
rect 29 1064 41 1098
rect 75 1064 113 1098
rect 147 1092 600 1098
rect 147 1064 482 1092
rect 29 1058 482 1064
rect 516 1058 554 1092
rect 588 1058 600 1092
rect 29 1052 600 1058
rect 3119 1083 3177 1089
rect 3119 1077 3131 1083
rect 3165 1077 3177 1083
rect 76 1018 1221 1024
rect 76 984 88 1018
rect 122 984 160 1018
rect 194 984 853 1018
rect 887 984 925 1018
rect 959 984 1103 1018
rect 1137 984 1175 1018
rect 1209 984 1221 1018
rect 76 978 1221 984
rect 1489 1022 2347 1034
rect 1489 988 1495 1022
rect 1529 988 2301 1022
rect 2335 988 2347 1022
rect 1489 950 2347 988
rect 262 944 1120 950
rect 262 910 274 944
rect 308 910 346 944
rect 380 910 709 944
rect 743 910 781 944
rect 815 910 1002 944
rect 1036 910 1074 944
rect 1108 910 1120 944
rect 262 904 1120 910
rect 1489 916 1495 950
rect 1529 916 2301 950
rect 2335 916 2347 950
rect 2715 1022 3073 1034
rect 2715 988 2721 1022
rect 2755 988 3033 1022
rect 3067 988 3073 1022
rect 2715 977 2775 988
tri 2775 977 2786 988 nw
tri 3002 977 3013 988 ne
rect 3013 977 3073 988
rect 2715 950 2761 977
tri 2761 963 2775 977 nw
tri 3013 963 3027 977 ne
rect 1489 904 2347 916
rect 2617 936 2675 942
rect 2617 902 2629 936
rect 2663 902 2675 936
rect 2715 916 2721 950
rect 2755 916 2761 950
rect 2715 904 2761 916
rect 2871 945 2917 957
rect 2871 911 2877 945
rect 2911 911 2917 945
rect 2871 904 2917 911
rect 3027 950 3073 977
rect 3027 916 3033 950
rect 3067 916 3073 950
tri 2917 904 2918 905 sw
rect 3027 904 3073 916
rect 3119 1025 3122 1077
rect 3174 1025 3177 1077
rect 3119 1013 3177 1025
rect 3119 961 3122 1013
rect 3174 961 3177 1013
rect 3119 949 3177 961
tri 3118 904 3119 905 se
rect 3119 904 3122 949
tri 2592 876 2617 901 se
rect 2617 876 2675 902
rect 570 824 576 876
rect 628 824 640 876
rect 692 864 2675 876
rect 692 830 2629 864
rect 2663 830 2675 864
rect 692 824 2675 830
rect 2871 873 2918 904
rect 2871 839 2877 873
rect 2911 871 2918 873
tri 2918 871 2951 904 sw
tri 3085 871 3118 904 se
rect 3118 897 3122 904
rect 3174 897 3177 949
rect 3118 885 3177 897
rect 3118 871 3122 885
rect 2911 839 3122 871
rect 2871 833 3122 839
rect 3174 833 3177 885
rect 2871 827 3177 833
rect -179 452 3312 464
rect -179 346 959 452
rect 1137 418 2503 452
rect 2537 418 3312 452
rect 1137 380 3312 418
rect 1137 346 2503 380
rect 2537 346 3312 380
rect -179 334 3312 346
rect -179 294 3312 306
rect -179 260 -17 294
rect 17 260 425 294
rect 459 260 717 294
rect 751 260 3312 294
rect -179 222 3312 260
rect -179 188 -17 222
rect 17 188 425 222
rect 459 188 717 222
rect 751 188 3312 222
rect -179 150 3312 188
rect -179 116 -17 150
rect 17 116 425 150
rect 459 116 717 150
rect 751 116 3312 150
rect -179 104 3312 116
<< via1 >>
rect 2424 2348 2476 2400
rect 2488 2348 2540 2400
rect 2658 2274 2774 2390
rect 3122 2194 3174 2246
rect 3122 2130 3174 2182
rect 3122 2066 3174 2118
rect 3122 2002 3174 2054
rect 3122 1938 3174 1990
rect 2658 1874 2710 1880
rect 2722 1874 2774 1880
rect 2658 1840 2690 1874
rect 2690 1840 2710 1874
rect 2722 1840 2724 1874
rect 2724 1840 2774 1874
rect 2658 1828 2710 1840
rect 2722 1828 2774 1840
rect 2395 1619 2447 1671
rect 2459 1619 2511 1671
rect 640 1548 692 1600
rect 640 1484 692 1536
rect 3122 1595 3174 1601
rect 3122 1561 3131 1595
rect 3131 1561 3165 1595
rect 3165 1561 3174 1595
rect 3122 1549 3174 1561
rect 3122 1523 3174 1537
rect 3122 1489 3131 1523
rect 3131 1489 3165 1523
rect 3165 1489 3174 1523
rect 3122 1485 3174 1489
rect 3122 1049 3131 1077
rect 3131 1049 3165 1077
rect 3165 1049 3174 1077
rect 3122 1025 3174 1049
rect 3122 1011 3174 1013
rect 3122 977 3131 1011
rect 3131 977 3165 1011
rect 3165 977 3174 1011
rect 3122 961 3174 977
rect 3122 939 3174 949
rect 3122 905 3131 939
rect 3131 905 3165 939
rect 3165 905 3174 939
rect 576 824 628 876
rect 640 824 692 876
rect 3122 897 3174 905
rect 3122 867 3174 885
rect 3122 833 3131 867
rect 3131 833 3165 867
rect 3165 833 3174 867
<< metal2 >>
rect 2418 2348 2424 2400
rect 2476 2348 2488 2400
rect 2540 2348 2546 2400
rect 2418 1700 2482 2348
tri 2482 2323 2507 2348 nw
rect 2652 2274 2658 2390
rect 2774 2274 2780 2390
rect 2652 1880 2780 2274
rect 2652 1828 2658 1880
rect 2710 1828 2722 1880
rect 2774 1828 2780 1880
rect 3116 2194 3122 2246
rect 3174 2194 3180 2246
rect 3116 2182 3180 2194
rect 3116 2130 3122 2182
rect 3174 2130 3180 2182
rect 3116 2118 3180 2130
rect 3116 2066 3122 2118
rect 3174 2066 3180 2118
rect 3116 2054 3180 2066
rect 3116 2002 3122 2054
rect 3174 2002 3180 2054
rect 3116 1990 3180 2002
rect 3116 1938 3122 1990
rect 3174 1938 3180 1990
tri 2482 1700 2488 1706 sw
tri 2395 1677 2418 1700 se
rect 2418 1677 2488 1700
tri 2488 1677 2511 1700 sw
rect 2395 1671 2511 1677
rect 2447 1619 2459 1671
rect 2395 1613 2511 1619
rect 3116 1601 3180 1938
rect 634 1600 698 1601
rect 634 1548 640 1600
rect 692 1548 698 1600
rect 634 1536 698 1548
rect 634 1484 640 1536
rect 692 1484 698 1536
tri 630 897 634 901 se
rect 634 897 698 1484
tri 618 885 630 897 se
rect 630 885 698 897
tri 609 876 618 885 se
rect 618 876 698 885
rect 570 824 576 876
rect 628 824 640 876
rect 692 824 698 876
rect 3116 1549 3122 1601
rect 3174 1549 3180 1601
rect 3116 1537 3180 1549
rect 3116 1485 3122 1537
rect 3174 1485 3180 1537
rect 3116 1077 3180 1485
rect 3116 1025 3122 1077
rect 3174 1025 3180 1077
rect 3116 1013 3180 1025
rect 3116 961 3122 1013
rect 3174 961 3180 1013
rect 3116 949 3180 961
rect 3116 897 3122 949
rect 3174 897 3180 949
rect 3116 885 3180 897
rect 3116 833 3122 885
rect 3174 833 3180 885
rect 3116 827 3180 833
<< comment >>
rect 2251 2333 2488 2420
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1707688321
transform -1 0 415 0 -1 1735
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_1
timestamp 1707688321
transform 0 1 641 1 0 1815
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_2
timestamp 1707688321
transform 0 1 570 1 0 1717
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_3
timestamp 1707688321
transform 1 0 3131 0 -1 1595
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_4
timestamp 1707688321
transform 1 0 2956 0 -1 1755
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_5
timestamp 1707688321
transform 1 0 2799 0 -1 1755
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_6
timestamp 1707688321
transform 1 0 2301 0 -1 1595
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_7
timestamp 1707688321
transform 1 0 2091 0 -1 1595
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_8
timestamp 1707688321
transform 1 0 2629 0 -1 936
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_9
timestamp 1707688321
transform 1 0 565 0 1 1489
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_10
timestamp 1707688321
transform 1 0 2721 0 1 1489
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_11
timestamp 1707688321
transform 1 0 3033 0 1 1489
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1707688321
transform 0 -1 2537 -1 0 452
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1707688321
transform 0 -1 1529 -1 0 1022
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1707688321
transform 0 -1 2335 -1 0 1022
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1707688321
transform 0 1 481 -1 0 1849
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1707688321
transform 0 1 2503 -1 0 452
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1707688321
transform -1 0 194 0 1 984
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1707688321
transform -1 0 380 0 1 910
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1707688321
transform -1 0 600 0 1 1297
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1707688321
transform -1 0 959 0 1 984
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_9
timestamp 1707688321
transform -1 0 1108 0 1 910
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_10
timestamp 1707688321
transform -1 0 815 0 1 910
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_11
timestamp 1707688321
transform -1 0 147 0 -1 1098
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_12
timestamp 1707688321
transform -1 0 515 0 -1 1403
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_13
timestamp 1707688321
transform 0 -1 2911 1 0 839
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_14
timestamp 1707688321
transform 0 -1 2755 1 0 916
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_15
timestamp 1707688321
transform 0 -1 3067 1 0 916
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_16
timestamp 1707688321
transform 1 0 2279 0 1 2354
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_17
timestamp 1707688321
transform 1 0 781 0 1 1489
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_18
timestamp 1707688321
transform 1 0 1519 0 1 1489
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_19
timestamp 1707688321
transform 1 0 2618 0 1 1840
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_20
timestamp 1707688321
transform 1 0 432 0 1 2280
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_21
timestamp 1707688321
transform 1 0 2581 0 1 1637
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_22
timestamp 1707688321
transform 1 0 482 0 1 1058
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_23
timestamp 1707688321
transform 1 0 1103 0 1 984
box 0 0 1 1
use L1M1_CDNS_5246887918558  L1M1_CDNS_5246887918558_0
timestamp 1707688321
transform 0 1 959 -1 0 452
box 0 0 1 1
use L1M1_CDNS_5246887918558  L1M1_CDNS_5246887918558_1
timestamp 1707688321
transform -1 0 2043 0 -1 2090
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1707688321
transform 0 -1 991 -1 0 1443
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1707688321
transform 0 -1 2421 -1 0 1443
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_2
timestamp 1707688321
transform 0 -1 2249 -1 0 1443
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_3
timestamp 1707688321
transform 0 1 2503 -1 0 1443
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_4
timestamp 1707688321
transform 0 -1 459 1 0 116
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_5
timestamp 1707688321
transform 0 -1 17 1 0 116
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_6
timestamp 1707688321
transform 0 -1 751 1 0 116
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_0
timestamp 1707688321
transform -1 0 2968 0 -1 2094
box 0 0 1 1
use L1M1_CDNS_52468879185193  L1M1_CDNS_52468879185193_0
timestamp 1707688321
transform 0 1 253 -1 0 1849
box 0 0 1 1
use L1M1_CDNS_52468879185334  L1M1_CDNS_52468879185334_0
timestamp 1707688321
transform 0 -1 747 -1 0 1443
box 0 0 1 1
use L1M1_CDNS_52468879185334  L1M1_CDNS_52468879185334_1
timestamp 1707688321
transform 0 1 217 -1 0 1443
box 0 0 1 1
use L1M1_CDNS_524688791851057  L1M1_CDNS_524688791851057_0
timestamp 1707688321
transform 1 0 3131 0 -1 1083
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1707688321
transform 1 0 570 0 -1 876
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1707688321
transform 1 0 2418 0 1 2348
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1707688321
transform 1 0 2652 0 1 1828
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_0
timestamp 1707688321
transform 1 0 2652 0 1 2274
box 0 0 1 1
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_0
timestamp 1707688321
transform 0 -1 3174 -1 0 1083
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_0
timestamp 1707688321
transform 0 1 2395 -1 0 1677
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_1
timestamp 1707688321
transform 1 0 3116 0 -1 1601
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_2
timestamp 1707688321
transform 1 0 634 0 1 1484
box 0 0 1 1
use M1M2_CDNS_52468879185972  M1M2_CDNS_52468879185972_0
timestamp 1707688321
transform 1 0 3116 0 -1 2246
box 0 0 1 1
use nfet_CDNS_52468879185411  nfet_CDNS_52468879185411_0
timestamp 1707688321
transform -1 0 206 0 -1 1282
box -79 -26 202 226
use nfet_CDNS_52468879185412  nfet_CDNS_52468879185412_0
timestamp 1707688321
transform 1 0 262 0 -1 1282
box -82 -26 202 226
use nfet_CDNS_52468879185413  nfet_CDNS_52468879185413_0
timestamp 1707688321
transform 1 0 1002 0 -1 2024
box -82 -26 199 626
use nfet_CDNS_52468879185414  nfet_CDNS_52468879185414_0
timestamp 1707688321
transform -1 0 946 0 -1 2024
box -82 -26 199 626
use nfet_CDNS_52468879185432  nfet_CDNS_52468879185432_0
timestamp 1707688321
transform 1 0 1620 0 -1 2202
box -79 -26 179 1026
use nfet_CDNS_52468879185433  nfet_CDNS_52468879185433_0
timestamp 1707688321
transform -1 0 1411 0 -1 2202
box -82 -26 179 1026
use nfet_CDNS_52468879185434  nfet_CDNS_52468879185434_0
timestamp 1707688321
transform -1 0 946 0 -1 1222
box -79 -26 199 166
use nfet_CDNS_52468879185435  nfet_CDNS_52468879185435_0
timestamp 1707688321
transform 1 0 1002 0 -1 1222
box -82 -26 199 166
use nfet_CDNS_52468879185436  nfet_CDNS_52468879185436_0
timestamp 1707688321
transform 1 0 1304 0 1 908
box -79 -26 495 226
use nfet_CDNS_52468879185436  nfet_CDNS_52468879185436_1
timestamp 1707688321
transform 1 0 1304 0 1 388
box -79 -26 495 226
use nfet_CDNS_52468879185436  nfet_CDNS_52468879185436_2
timestamp 1707688321
transform 1 0 1304 0 1 128
box -79 -26 495 226
use nfet_CDNS_52468879185436  nfet_CDNS_52468879185436_3
timestamp 1707688321
transform 1 0 1304 0 1 648
box -79 -26 495 226
use nfet_CDNS_52468879185437  nfet_CDNS_52468879185437_0
timestamp 1707688321
transform 1 0 1900 0 1 908
box -79 -26 259 226
use nfet_CDNS_52468879185437  nfet_CDNS_52468879185437_1
timestamp 1707688321
transform 1 0 1900 0 1 648
box -79 -26 259 226
use nfet_CDNS_52468879185437  nfet_CDNS_52468879185437_2
timestamp 1707688321
transform 1 0 1900 0 1 128
box -79 -26 259 226
use nfet_CDNS_52468879185437  nfet_CDNS_52468879185437_3
timestamp 1707688321
transform 1 0 1900 0 1 1482
box -79 -26 259 226
use nfet_CDNS_52468879185437  nfet_CDNS_52468879185437_4
timestamp 1707688321
transform 1 0 1900 0 1 388
box -79 -26 259 226
use nfet_CDNS_52468879185437  nfet_CDNS_52468879185437_5
timestamp 1707688321
transform 1 0 1900 0 1 1742
box -79 -26 259 226
use nfet_CDNS_52468879185437  nfet_CDNS_52468879185437_6
timestamp 1707688321
transform 1 0 1900 0 1 1222
box -79 -26 259 226
use nfet_CDNS_52468879185437  nfet_CDNS_52468879185437_7
timestamp 1707688321
transform 1 0 1900 0 1 2002
box -79 -26 259 226
use nfet_CDNS_52468879185438  nfet_CDNS_52468879185438_0
timestamp 1707688321
transform 1 0 2260 0 1 388
box -79 -26 195 226
use nfet_CDNS_52468879185438  nfet_CDNS_52468879185438_1
timestamp 1707688321
transform 1 0 2260 0 1 128
box -79 -26 195 226
use nfet_CDNS_52468879185438  nfet_CDNS_52468879185438_2
timestamp 1707688321
transform 1 0 2260 0 1 1742
box -79 -26 195 226
use nfet_CDNS_52468879185438  nfet_CDNS_52468879185438_3
timestamp 1707688321
transform 1 0 2260 0 1 2002
box -79 -26 195 226
use nfet_CDNS_52468879185438  nfet_CDNS_52468879185438_4
timestamp 1707688321
transform 1 0 2260 0 1 1222
box -79 -26 195 226
use nfet_CDNS_52468879185438  nfet_CDNS_52468879185438_5
timestamp 1707688321
transform 1 0 2260 0 1 1482
box -79 -26 195 226
use nfet_CDNS_52468879185438  nfet_CDNS_52468879185438_6
timestamp 1707688321
transform 1 0 2260 0 1 648
box -79 -26 195 226
use nfet_CDNS_52468879185438  nfet_CDNS_52468879185438_7
timestamp 1707688321
transform 1 0 2260 0 1 908
box -79 -26 195 226
use nfet_CDNS_524688791851425  nfet_CDNS_524688791851425_0
timestamp 1707688321
transform -1 0 646 0 1 1424
box -79 -26 115 226
use nfet_CDNS_524688791851425  nfet_CDNS_524688791851425_1
timestamp 1707688321
transform -1 0 646 0 1 1824
box -79 -26 115 226
use nfet_CDNS_524688791851425  nfet_CDNS_524688791851425_2
timestamp 1707688321
transform 1 0 518 0 1 1424
box -79 -26 115 226
use nfet_CDNS_524688791851425  nfet_CDNS_524688791851425_3
timestamp 1707688321
transform 1 0 518 0 1 1824
box -79 -26 115 226
use pfet_CDNS_52468879185440  pfet_CDNS_52468879185440_0
timestamp 1707688321
transform 1 0 28 0 -1 432
box -119 -66 219 266
use pfet_CDNS_52468879185441  pfet_CDNS_52468879185441_0
timestamp 1707688321
transform 1 0 28 0 -1 859
box -119 -66 219 266
use pfet_CDNS_52468879185442  pfet_CDNS_52468879185442_0
timestamp 1707688321
transform 1 0 470 0 -1 732
box -119 -66 219 666
use pfet_CDNS_52468879185443  pfet_CDNS_52468879185443_0
timestamp 1707688321
transform -1 0 414 0 -1 732
box -119 -66 219 666
use pfet_CDNS_524688791851426  pfet_CDNS_524688791851426_0
timestamp 1707688321
transform -1 0 3022 0 1 502
box -89 -36 345 636
use pfet_CDNS_524688791851426  pfet_CDNS_524688791851426_1
timestamp 1707688321
transform 1 0 2766 0 1 1268
box -89 -36 345 636
use pfet_CDNS_524688791851427  pfet_CDNS_524688791851427_0
timestamp 1707688321
transform -1 0 2710 0 1 502
box -89 -36 125 636
use pfet_CDNS_524688791851427  pfet_CDNS_524688791851427_1
timestamp 1707688321
transform -1 0 2710 0 1 1268
box -89 -36 125 636
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_0
timestamp 1707688321
transform -1 0 457 0 1 1660
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_1
timestamp 1707688321
transform -1 0 2703 0 -1 1200
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_2
timestamp 1707688321
transform 0 1 853 1 0 922
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_3
timestamp 1707688321
transform 0 1 1002 1 0 922
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_4
timestamp 1707688321
transform 0 -1 676 1 0 1660
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1707688321
transform 0 -1 2724 -1 0 1966
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_1
timestamp 1707688321
transform 0 1 420 -1 0 2174
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_2
timestamp 1707688321
transform 0 1 812 -1 0 2122
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_3
timestamp 1707688321
transform 0 1 1002 -1 0 2122
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_4
timestamp 1707688321
transform 0 1 1923 1 0 1132
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_5
timestamp 1707688321
transform 0 1 2766 1 0 1900
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_6
timestamp 1707688321
transform 0 1 470 1 0 14
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_7
timestamp 1707688321
transform 0 1 2251 1 0 2228
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_8
timestamp 1707688321
transform 0 1 2251 1 0 36
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_9
timestamp 1707688321
transform 0 1 1923 1 0 2228
box 0 0 1 1
use PYL1_CDNS_52468879185309  PYL1_CDNS_52468879185309_0
timestamp 1707688321
transform 0 1 2766 1 0 404
box 0 0 1 1
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_0
timestamp 1707688321
transform 0 1 1312 1 0 36
box 0 0 66 746
use PYL1_CDNS_52468879185327  PYL1_CDNS_52468879185327_0
timestamp 1707688321
transform 0 -1 1719 -1 0 2294
box 0 0 1 1
use PYL1_CDNS_52468879185429  PYL1_CDNS_52468879185429_0
timestamp 1707688321
transform 0 1 51 -1 0 1046
box 0 0 1 1
use PYL1_CDNS_52468879185429  PYL1_CDNS_52468879185429_1
timestamp 1707688321
transform 1 0 262 0 -1 1050
box 0 0 1 1
use TPL1_CDNS_52468879185430  TPL1_CDNS_52468879185430_0
timestamp 1707688321
transform -1 0 1161 0 1 92
box -26 -26 244 788
<< labels >>
flabel comment s 1213 1832 1213 1832 0 FreeSans 300 180 0 0 fbk_n
flabel comment s 2578 63 2578 63 0 FreeSans 400 0 0 0 in_i
flabel comment s 1197 1497 1197 1497 0 FreeSans 300 180 0 0 fbk
flabel comment s 2887 1546 2887 1546 0 FreeSans 300 0 0 0 virt_pwr
flabel comment s 388 727 388 727 0 FreeSans 200 0 0 0 out_h_n
flabel comment s 812 1318 812 1318 0 FreeSans 300 270 0 0 fbk
flabel comment s 1142 1338 1142 1338 0 FreeSans 300 90 0 0 fbk_n
flabel comment s 1512 1295 1512 1295 0 FreeSans 200 0 0 0 to hvnatives
flabel comment s 1405 1655 1405 1655 0 FreeSans 300 0 0 0 in_i_n
flabel comment s 1516 2251 1516 2251 0 FreeSans 200 180 0 0 hld_h_n
flabel comment s 2618 1197 2618 1197 0 FreeSans 400 180 0 0 in_i_n
flabel comment s 491 2167 491 2167 0 FreeSans 300 180 0 0 in
flabel comment s 579 1745 579 1745 0 FreeSans 300 180 0 0 in_dis
flabel comment s 572 2028 572 2028 0 FreeSans 400 180 0 0 in_i_n
flabel comment s 766 836 766 836 0 FreeSans 300 180 0 0 in_i
flabel comment s 1065 1048 1065 1048 0 FreeSans 300 0 0 0 fbk
flabel comment s 870 1048 870 1048 0 FreeSans 300 0 0 0 fbk_n
flabel metal1 s -96 1253 -56 1455 3 FreeSans 300 180 0 0 vgnd
port 2 nsew
flabel metal1 s 2607 1834 2657 1864 3 FreeSans 300 180 0 0 in
port 4 nsew
flabel metal1 s 10 1898 45 2246 3 FreeSans 300 180 0 0 vpwr_ka
port 5 nsew
flabel metal1 s 3277 1898 3312 2246 7 FreeSans 300 0 0 0 vpwr_ka
port 5 nsew
flabel metal1 s 3277 1253 3312 1455 7 FreeSans 300 180 0 0 vgnd
port 2 nsew
flabel metal1 s 543 1052 578 1104 7 FreeSans 400 180 0 0 out_h
port 1 nsew
flabel metal1 s 3277 334 3312 464 7 FreeSans 300 180 0 0 vgnd
port 2 nsew
flabel metal1 s -179 104 -144 306 3 FreeSans 300 180 0 0 vcc_io
port 3 nsew
flabel metal1 s -179 334 -144 464 3 FreeSans 300 180 0 0 vgnd
port 2 nsew
flabel metal1 s 3277 104 3312 306 7 FreeSans 300 180 0 0 vcc_io
port 3 nsew
flabel locali s 1496 2245 1536 2277 0 FreeSans 200 0 0 0 hld_h_n
port 7 nsew
flabel locali s 2986 420 3036 454 7 FreeSans 300 180 0 0 in_dis
port 8 nsew
flabel locali s 1096 2333 1136 2379 7 FreeSans 300 180 0 0 set_h
port 9 nsew
flabel locali s 812 2333 852 2379 3 FreeSans 300 180 0 0 rst_h
port 10 nsew
flabel locali s 413 1105 448 1151 7 FreeSans 300 180 0 0 out_h_n
port 11 nsew
<< properties >>
string GDS_END 87559834
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87534720
string path 18.350 2.650 18.350 18.950 
<< end >>
