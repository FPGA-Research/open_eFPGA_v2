magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect 0 2274 1022 2440
rect 0 166 166 2274
rect 856 166 1022 2274
rect 0 0 1022 166
<< mvnsubdiff >>
rect 66 2350 156 2374
rect 100 2340 156 2350
rect 190 2340 230 2374
rect 264 2340 304 2374
rect 338 2340 378 2374
rect 412 2340 452 2374
rect 486 2340 526 2374
rect 560 2340 600 2374
rect 634 2340 674 2374
rect 708 2340 747 2374
rect 781 2340 820 2374
rect 854 2350 956 2374
rect 854 2340 922 2350
rect 66 2279 100 2316
rect 922 2280 956 2316
rect 66 2208 100 2245
rect 66 2137 100 2174
rect 66 2066 100 2103
rect 66 1995 100 2032
rect 66 1924 100 1961
rect 66 1853 100 1890
rect 66 1782 100 1819
rect 66 1711 100 1748
rect 66 1640 100 1677
rect 66 1569 100 1606
rect 66 1498 100 1535
rect 66 1427 100 1464
rect 66 1356 100 1393
rect 66 1286 100 1322
rect 66 1216 100 1252
rect 66 1146 100 1182
rect 66 1076 100 1112
rect 66 1006 100 1042
rect 66 936 100 972
rect 66 866 100 902
rect 66 796 100 832
rect 66 590 100 762
rect 66 513 100 556
rect 66 436 100 479
rect 66 358 100 402
rect 66 280 100 324
rect 66 202 100 246
rect 922 2210 956 2246
rect 922 2140 956 2176
rect 922 2070 956 2106
rect 922 2000 956 2036
rect 922 1930 956 1966
rect 922 1860 956 1896
rect 922 1790 956 1826
rect 922 1720 956 1756
rect 922 1650 956 1686
rect 922 1580 956 1616
rect 922 1510 956 1546
rect 922 1440 956 1476
rect 922 1370 956 1406
rect 922 1300 956 1336
rect 922 1230 956 1266
rect 922 1160 956 1196
rect 922 1091 956 1126
rect 922 1022 956 1057
rect 922 953 956 988
rect 922 884 956 919
rect 922 815 956 850
rect 922 746 956 781
rect 922 677 956 712
rect 922 608 956 643
rect 922 539 956 574
rect 922 470 956 505
rect 922 401 956 436
rect 922 332 956 367
rect 922 263 956 298
rect 922 194 956 229
rect 66 124 100 168
rect 922 100 956 160
rect 100 90 168 100
rect 66 66 168 90
rect 202 66 241 100
rect 275 66 314 100
rect 348 66 387 100
rect 421 66 460 100
rect 494 66 533 100
rect 567 66 606 100
rect 640 66 679 100
rect 713 66 752 100
rect 786 66 825 100
rect 859 66 898 100
rect 932 66 956 100
<< mvnsubdiffcont >>
rect 66 2316 100 2350
rect 156 2340 190 2374
rect 230 2340 264 2374
rect 304 2340 338 2374
rect 378 2340 412 2374
rect 452 2340 486 2374
rect 526 2340 560 2374
rect 600 2340 634 2374
rect 674 2340 708 2374
rect 747 2340 781 2374
rect 820 2340 854 2374
rect 66 2245 100 2279
rect 922 2316 956 2350
rect 922 2246 956 2280
rect 66 2174 100 2208
rect 66 2103 100 2137
rect 66 2032 100 2066
rect 66 1961 100 1995
rect 66 1890 100 1924
rect 66 1819 100 1853
rect 66 1748 100 1782
rect 66 1677 100 1711
rect 66 1606 100 1640
rect 66 1535 100 1569
rect 66 1464 100 1498
rect 66 1393 100 1427
rect 66 1322 100 1356
rect 66 1252 100 1286
rect 66 1182 100 1216
rect 66 1112 100 1146
rect 66 1042 100 1076
rect 66 972 100 1006
rect 66 902 100 936
rect 66 832 100 866
rect 66 762 100 796
rect 66 556 100 590
rect 66 479 100 513
rect 66 402 100 436
rect 66 324 100 358
rect 66 246 100 280
rect 66 168 100 202
rect 922 2176 956 2210
rect 922 2106 956 2140
rect 922 2036 956 2070
rect 922 1966 956 2000
rect 922 1896 956 1930
rect 922 1826 956 1860
rect 922 1756 956 1790
rect 922 1686 956 1720
rect 922 1616 956 1650
rect 922 1546 956 1580
rect 922 1476 956 1510
rect 922 1406 956 1440
rect 922 1336 956 1370
rect 922 1266 956 1300
rect 922 1196 956 1230
rect 922 1126 956 1160
rect 922 1057 956 1091
rect 922 988 956 1022
rect 922 919 956 953
rect 922 850 956 884
rect 922 781 956 815
rect 922 712 956 746
rect 922 643 956 677
rect 922 574 956 608
rect 922 505 956 539
rect 922 436 956 470
rect 922 367 956 401
rect 922 298 956 332
rect 922 229 956 263
rect 66 90 100 124
rect 922 160 956 194
rect 168 66 202 100
rect 241 66 275 100
rect 314 66 348 100
rect 387 66 421 100
rect 460 66 494 100
rect 533 66 567 100
rect 606 66 640 100
rect 679 66 713 100
rect 752 66 786 100
rect 825 66 859 100
rect 898 66 932 100
<< poly >>
rect 227 2246 327 2318
rect 383 2246 483 2318
rect 539 2246 639 2318
rect 695 2246 795 2318
rect 227 122 327 194
rect 383 122 483 194
rect 539 122 639 194
rect 695 122 795 194
<< locali >>
rect 66 2350 156 2374
rect 100 2340 156 2350
rect 190 2340 230 2374
rect 264 2340 304 2374
rect 338 2340 378 2374
rect 412 2340 452 2374
rect 486 2340 526 2374
rect 560 2340 600 2374
rect 634 2340 674 2374
rect 708 2340 747 2374
rect 781 2340 820 2374
rect 854 2350 956 2374
rect 854 2340 922 2350
rect 66 2279 100 2316
rect 250 2300 304 2302
rect 406 2300 460 2302
rect 562 2300 616 2302
rect 718 2300 772 2302
rect 274 2266 312 2300
rect 346 2266 384 2300
rect 418 2266 456 2300
rect 490 2266 529 2300
rect 563 2266 602 2300
rect 636 2266 675 2300
rect 709 2266 748 2300
rect 922 2280 956 2316
rect 66 2208 100 2245
rect 66 2137 100 2174
rect 66 2066 100 2103
rect 66 1995 100 2032
rect 66 1924 100 1961
rect 66 1853 100 1890
rect 66 1782 100 1819
rect 66 1711 100 1748
rect 66 1640 100 1677
rect 66 1569 100 1606
rect 66 1498 100 1535
rect 66 1427 100 1464
rect 66 1356 100 1393
rect 66 1286 100 1322
rect 66 1216 100 1252
rect 66 1146 100 1182
rect 66 1076 100 1112
rect 66 1006 100 1042
rect 66 936 100 972
rect 66 866 100 902
rect 66 796 100 832
rect 66 590 100 762
rect 66 513 100 556
rect 66 436 100 479
rect 66 358 100 402
rect 66 280 100 324
rect 182 2112 216 2151
rect 182 2039 216 2078
rect 182 1966 216 2005
rect 182 1893 216 1932
rect 182 1820 216 1859
rect 182 1747 216 1786
rect 182 1674 216 1713
rect 182 1601 216 1640
rect 182 1528 216 1567
rect 182 1455 216 1494
rect 182 1382 216 1421
rect 182 1309 216 1348
rect 182 1236 216 1275
rect 182 1163 216 1202
rect 182 1090 216 1129
rect 182 1017 216 1056
rect 182 944 216 983
rect 182 871 216 910
rect 182 798 216 837
rect 182 725 216 764
rect 182 652 216 691
rect 182 579 216 618
rect 182 506 216 545
rect 182 433 216 472
rect 182 361 216 399
rect 182 289 216 327
rect 66 202 100 246
rect 250 174 304 2266
rect 338 2110 372 2151
rect 338 2035 372 2076
rect 338 1960 372 2001
rect 338 1885 372 1926
rect 338 1810 372 1851
rect 338 1735 372 1776
rect 338 1660 372 1701
rect 338 1585 372 1626
rect 338 1510 372 1551
rect 338 1435 372 1476
rect 338 1360 372 1401
rect 338 1285 372 1326
rect 338 1210 372 1251
rect 338 1135 372 1176
rect 338 1060 372 1101
rect 338 986 372 1026
rect 338 912 372 952
rect 338 838 372 878
rect 338 764 372 804
rect 338 690 372 730
rect 338 616 372 656
rect 406 174 460 2266
rect 494 1762 528 1802
rect 494 1688 528 1728
rect 494 1614 528 1654
rect 494 1540 528 1580
rect 494 1466 528 1506
rect 494 1392 528 1432
rect 494 1318 528 1358
rect 494 1244 528 1284
rect 494 1170 528 1210
rect 494 1096 528 1136
rect 494 1022 528 1062
rect 494 948 528 988
rect 494 874 528 914
rect 494 800 528 840
rect 494 727 528 766
rect 494 654 528 693
rect 494 581 528 620
rect 494 508 528 547
rect 494 435 528 474
rect 494 362 528 401
rect 494 289 528 328
rect 562 174 616 2266
rect 650 2110 684 2151
rect 650 2035 684 2076
rect 650 1960 684 2001
rect 650 1885 684 1926
rect 650 1810 684 1851
rect 650 1735 684 1776
rect 650 1660 684 1701
rect 650 1585 684 1626
rect 650 1510 684 1551
rect 650 1435 684 1476
rect 650 1360 684 1401
rect 650 1285 684 1326
rect 650 1210 684 1251
rect 650 1135 684 1176
rect 650 1060 684 1101
rect 650 986 684 1026
rect 650 912 684 952
rect 650 838 684 878
rect 650 764 684 804
rect 650 690 684 730
rect 650 616 684 656
rect 718 174 772 2266
rect 922 2210 956 2246
rect 806 2112 840 2151
rect 806 2039 840 2078
rect 806 1966 840 2005
rect 806 1893 840 1932
rect 806 1820 840 1859
rect 806 1747 840 1786
rect 806 1674 840 1713
rect 806 1601 840 1640
rect 806 1528 840 1567
rect 806 1455 840 1494
rect 806 1382 840 1421
rect 806 1309 840 1348
rect 806 1236 840 1275
rect 806 1163 840 1202
rect 806 1090 840 1129
rect 806 1017 840 1056
rect 806 944 840 983
rect 806 871 840 910
rect 806 798 840 837
rect 806 725 840 764
rect 806 652 840 691
rect 806 579 840 618
rect 806 506 840 545
rect 806 433 840 472
rect 806 361 840 399
rect 806 289 840 327
rect 922 2140 956 2176
rect 922 2070 956 2106
rect 922 2000 956 2036
rect 922 1930 956 1966
rect 922 1860 956 1896
rect 922 1790 956 1826
rect 922 1720 956 1756
rect 922 1650 956 1686
rect 922 1580 956 1616
rect 922 1510 956 1546
rect 922 1440 956 1476
rect 922 1370 956 1406
rect 922 1300 956 1336
rect 922 1230 956 1266
rect 922 1160 956 1196
rect 922 1091 956 1126
rect 922 1022 956 1057
rect 922 953 956 988
rect 922 884 956 919
rect 922 815 956 850
rect 922 746 956 781
rect 922 677 956 712
rect 922 608 956 643
rect 922 539 956 574
rect 922 470 956 505
rect 922 401 956 436
rect 922 332 956 367
rect 922 263 956 298
rect 922 194 956 229
rect 66 124 100 168
rect 274 140 312 174
rect 346 140 384 174
rect 418 140 456 174
rect 490 140 529 174
rect 563 140 602 174
rect 636 140 675 174
rect 709 140 748 174
rect 250 138 304 140
rect 406 138 460 140
rect 562 138 616 140
rect 718 138 772 140
rect 922 100 956 160
rect 100 90 168 100
rect 66 66 168 90
rect 202 66 241 100
rect 275 66 314 100
rect 348 66 387 100
rect 421 66 460 100
rect 494 66 533 100
rect 567 66 606 100
rect 640 66 679 100
rect 713 66 752 100
rect 786 66 825 100
rect 859 66 898 100
rect 932 66 956 100
<< viali >>
rect 240 2266 274 2300
rect 312 2266 346 2300
rect 384 2266 418 2300
rect 456 2266 490 2300
rect 529 2266 563 2300
rect 602 2266 636 2300
rect 675 2266 709 2300
rect 748 2266 782 2300
rect 182 2151 216 2185
rect 182 2078 216 2112
rect 182 2005 216 2039
rect 182 1932 216 1966
rect 182 1859 216 1893
rect 182 1786 216 1820
rect 182 1713 216 1747
rect 182 1640 216 1674
rect 182 1567 216 1601
rect 182 1494 216 1528
rect 182 1421 216 1455
rect 182 1348 216 1382
rect 182 1275 216 1309
rect 182 1202 216 1236
rect 182 1129 216 1163
rect 182 1056 216 1090
rect 182 983 216 1017
rect 182 910 216 944
rect 182 837 216 871
rect 182 764 216 798
rect 182 691 216 725
rect 182 618 216 652
rect 182 545 216 579
rect 182 472 216 506
rect 182 399 216 433
rect 182 327 216 361
rect 182 255 216 289
rect 338 2151 372 2185
rect 338 2076 372 2110
rect 338 2001 372 2035
rect 338 1926 372 1960
rect 338 1851 372 1885
rect 338 1776 372 1810
rect 338 1701 372 1735
rect 338 1626 372 1660
rect 338 1551 372 1585
rect 338 1476 372 1510
rect 338 1401 372 1435
rect 338 1326 372 1360
rect 338 1251 372 1285
rect 338 1176 372 1210
rect 338 1101 372 1135
rect 338 1026 372 1060
rect 338 952 372 986
rect 338 878 372 912
rect 338 804 372 838
rect 338 730 372 764
rect 338 656 372 690
rect 338 582 372 616
rect 494 1802 528 1836
rect 494 1728 528 1762
rect 494 1654 528 1688
rect 494 1580 528 1614
rect 494 1506 528 1540
rect 494 1432 528 1466
rect 494 1358 528 1392
rect 494 1284 528 1318
rect 494 1210 528 1244
rect 494 1136 528 1170
rect 494 1062 528 1096
rect 494 988 528 1022
rect 494 914 528 948
rect 494 840 528 874
rect 494 766 528 800
rect 494 693 528 727
rect 494 620 528 654
rect 494 547 528 581
rect 494 474 528 508
rect 494 401 528 435
rect 494 328 528 362
rect 494 255 528 289
rect 650 2151 684 2185
rect 650 2076 684 2110
rect 650 2001 684 2035
rect 650 1926 684 1960
rect 650 1851 684 1885
rect 650 1776 684 1810
rect 650 1701 684 1735
rect 650 1626 684 1660
rect 650 1551 684 1585
rect 650 1476 684 1510
rect 650 1401 684 1435
rect 650 1326 684 1360
rect 650 1251 684 1285
rect 650 1176 684 1210
rect 650 1101 684 1135
rect 650 1026 684 1060
rect 650 952 684 986
rect 650 878 684 912
rect 650 804 684 838
rect 650 730 684 764
rect 650 656 684 690
rect 650 582 684 616
rect 806 2151 840 2185
rect 806 2078 840 2112
rect 806 2005 840 2039
rect 806 1932 840 1966
rect 806 1859 840 1893
rect 806 1786 840 1820
rect 806 1713 840 1747
rect 806 1640 840 1674
rect 806 1567 840 1601
rect 806 1494 840 1528
rect 806 1421 840 1455
rect 806 1348 840 1382
rect 806 1275 840 1309
rect 806 1202 840 1236
rect 806 1129 840 1163
rect 806 1056 840 1090
rect 806 983 840 1017
rect 806 910 840 944
rect 806 837 840 871
rect 806 764 840 798
rect 806 691 840 725
rect 806 618 840 652
rect 806 545 840 579
rect 806 472 840 506
rect 806 399 840 433
rect 806 327 840 361
rect 806 255 840 289
rect 240 140 274 174
rect 312 140 346 174
rect 384 140 418 174
rect 456 140 490 174
rect 529 140 563 174
rect 602 140 636 174
rect 675 140 709 174
rect 748 140 782 174
<< metal1 >>
rect 228 2300 794 2306
rect 228 2266 240 2300
rect 274 2266 312 2300
rect 346 2266 384 2300
rect 418 2266 456 2300
rect 490 2266 529 2300
rect 563 2266 602 2300
rect 636 2266 675 2300
rect 709 2266 748 2300
rect 782 2266 794 2300
rect 228 2254 794 2266
rect 176 2185 222 2197
rect 176 2151 182 2185
rect 216 2151 222 2185
rect 176 2112 222 2151
rect 176 2078 182 2112
rect 216 2078 222 2112
rect 176 2039 222 2078
rect 176 2005 182 2039
rect 216 2005 222 2039
rect 176 1966 222 2005
rect 176 1932 182 1966
rect 216 1932 222 1966
rect 176 1893 222 1932
rect 176 1859 182 1893
rect 216 1859 222 1893
rect 176 1820 222 1859
rect 176 1786 182 1820
rect 216 1786 222 1820
rect 176 1747 222 1786
rect 176 1713 182 1747
rect 216 1713 222 1747
rect 176 1674 222 1713
rect 176 1640 182 1674
rect 216 1640 222 1674
rect 176 1601 222 1640
rect 176 1567 182 1601
rect 216 1567 222 1601
rect 176 1528 222 1567
rect 176 1494 182 1528
rect 216 1494 222 1528
rect 176 1455 222 1494
rect 176 1421 182 1455
rect 216 1421 222 1455
rect 176 1382 222 1421
rect 176 1348 182 1382
rect 216 1348 222 1382
rect 176 1309 222 1348
rect 176 1275 182 1309
rect 216 1275 222 1309
rect 176 1236 222 1275
rect 176 1202 182 1236
rect 216 1202 222 1236
rect 176 1163 222 1202
rect 176 1129 182 1163
rect 216 1129 222 1163
rect 176 1090 222 1129
rect 176 1056 182 1090
rect 216 1056 222 1090
rect 176 1017 222 1056
rect 176 983 182 1017
rect 216 983 222 1017
rect 176 944 222 983
rect 176 910 182 944
rect 216 910 222 944
rect 176 871 222 910
rect 176 837 182 871
rect 216 837 222 871
rect 176 798 222 837
rect 176 764 182 798
rect 216 764 222 798
rect 176 725 222 764
rect 176 691 182 725
rect 216 691 222 725
rect 176 652 222 691
rect 176 618 182 652
rect 216 618 222 652
rect 176 579 222 618
rect 176 545 182 579
rect 216 545 222 579
rect 332 2185 690 2197
rect 332 2151 338 2185
rect 372 2151 650 2185
rect 684 2151 690 2185
rect 332 2110 690 2151
rect 332 2076 338 2110
rect 372 2076 650 2110
rect 684 2076 690 2110
rect 332 2035 690 2076
rect 332 2001 338 2035
rect 372 2001 650 2035
rect 684 2001 690 2035
rect 332 1961 690 2001
rect 332 1960 418 1961
tri 418 1960 419 1961 nw
tri 602 1960 603 1961 ne
rect 603 1960 690 1961
rect 332 1926 338 1960
rect 372 1926 384 1960
tri 384 1926 418 1960 nw
tri 603 1926 637 1960 ne
rect 637 1926 650 1960
rect 684 1926 690 1960
rect 332 1885 378 1926
tri 378 1920 384 1926 nw
tri 637 1920 643 1926 ne
rect 643 1920 690 1926
tri 643 1919 644 1920 ne
rect 332 1851 338 1885
rect 372 1851 378 1885
rect 332 1810 378 1851
rect 644 1885 690 1920
rect 644 1851 650 1885
rect 684 1851 690 1885
rect 332 1776 338 1810
rect 372 1776 378 1810
rect 332 1735 378 1776
rect 332 1701 338 1735
rect 372 1701 378 1735
rect 332 1660 378 1701
rect 332 1626 338 1660
rect 372 1626 378 1660
rect 332 1585 378 1626
rect 332 1551 338 1585
rect 372 1551 378 1585
rect 332 1510 378 1551
rect 332 1476 338 1510
rect 372 1476 378 1510
rect 332 1435 378 1476
rect 332 1401 338 1435
rect 372 1401 378 1435
rect 332 1360 378 1401
rect 332 1326 338 1360
rect 372 1326 378 1360
rect 332 1285 378 1326
rect 332 1251 338 1285
rect 372 1251 378 1285
rect 332 1210 378 1251
rect 332 1176 338 1210
rect 372 1176 378 1210
rect 332 1135 378 1176
rect 332 1101 338 1135
rect 372 1101 378 1135
rect 332 1060 378 1101
rect 332 1026 338 1060
rect 372 1026 378 1060
rect 332 986 378 1026
rect 332 952 338 986
rect 372 952 378 986
rect 332 912 378 952
rect 332 878 338 912
rect 372 878 378 912
rect 332 838 378 878
rect 332 804 338 838
rect 372 804 378 838
rect 332 764 378 804
rect 332 730 338 764
rect 372 730 378 764
rect 332 690 378 730
rect 332 656 338 690
rect 372 656 378 690
rect 332 616 378 656
rect 332 582 338 616
rect 372 582 378 616
rect 332 570 378 582
rect 488 1836 534 1848
rect 488 1802 494 1836
rect 528 1802 534 1836
rect 488 1762 534 1802
rect 488 1728 494 1762
rect 528 1728 534 1762
rect 488 1688 534 1728
rect 488 1654 494 1688
rect 528 1654 534 1688
rect 488 1614 534 1654
rect 488 1580 494 1614
rect 528 1580 534 1614
rect 488 1540 534 1580
rect 488 1506 494 1540
rect 528 1506 534 1540
rect 488 1466 534 1506
rect 488 1432 494 1466
rect 528 1432 534 1466
rect 488 1392 534 1432
rect 488 1358 494 1392
rect 528 1358 534 1392
rect 488 1318 534 1358
rect 488 1284 494 1318
rect 528 1284 534 1318
rect 488 1244 534 1284
rect 488 1210 494 1244
rect 528 1210 534 1244
rect 488 1170 534 1210
rect 488 1136 494 1170
rect 528 1136 534 1170
rect 488 1096 534 1136
rect 488 1062 494 1096
rect 528 1062 534 1096
rect 488 1022 534 1062
rect 488 988 494 1022
rect 528 988 534 1022
rect 488 948 534 988
rect 488 914 494 948
rect 528 914 534 948
rect 488 874 534 914
rect 488 840 494 874
rect 528 840 534 874
rect 488 800 534 840
rect 488 766 494 800
rect 528 766 534 800
rect 488 727 534 766
rect 488 693 494 727
rect 528 693 534 727
rect 488 654 534 693
rect 488 620 494 654
rect 528 620 534 654
rect 488 581 534 620
rect 176 513 222 545
rect 488 547 494 581
rect 528 547 534 581
rect 644 1810 690 1851
rect 644 1776 650 1810
rect 684 1776 690 1810
rect 644 1735 690 1776
rect 644 1701 650 1735
rect 684 1701 690 1735
rect 644 1660 690 1701
rect 644 1626 650 1660
rect 684 1626 690 1660
rect 644 1585 690 1626
rect 644 1551 650 1585
rect 684 1551 690 1585
rect 644 1510 690 1551
rect 644 1476 650 1510
rect 684 1476 690 1510
rect 644 1435 690 1476
rect 644 1401 650 1435
rect 684 1401 690 1435
rect 644 1360 690 1401
rect 644 1326 650 1360
rect 684 1326 690 1360
rect 644 1285 690 1326
rect 644 1251 650 1285
rect 684 1251 690 1285
rect 644 1210 690 1251
rect 644 1176 650 1210
rect 684 1176 690 1210
rect 644 1135 690 1176
rect 644 1101 650 1135
rect 684 1101 690 1135
rect 644 1060 690 1101
rect 644 1026 650 1060
rect 684 1026 690 1060
rect 644 986 690 1026
rect 644 952 650 986
rect 684 952 690 986
rect 644 912 690 952
rect 644 878 650 912
rect 684 878 690 912
rect 644 838 690 878
rect 644 804 650 838
rect 684 804 690 838
rect 644 764 690 804
rect 644 730 650 764
rect 684 730 690 764
rect 644 690 690 730
rect 644 656 650 690
rect 684 656 690 690
rect 644 616 690 656
rect 644 582 650 616
rect 684 582 690 616
rect 644 570 690 582
rect 800 2185 846 2197
rect 800 2151 806 2185
rect 840 2151 846 2185
rect 800 2112 846 2151
rect 800 2078 806 2112
rect 840 2078 846 2112
rect 800 2039 846 2078
rect 800 2005 806 2039
rect 840 2005 846 2039
rect 800 1966 846 2005
rect 800 1932 806 1966
rect 840 1932 846 1966
rect 800 1893 846 1932
rect 800 1859 806 1893
rect 840 1859 846 1893
rect 800 1820 846 1859
rect 800 1786 806 1820
rect 840 1786 846 1820
rect 800 1747 846 1786
rect 800 1713 806 1747
rect 840 1713 846 1747
rect 800 1674 846 1713
rect 800 1640 806 1674
rect 840 1640 846 1674
rect 800 1601 846 1640
rect 800 1567 806 1601
rect 840 1567 846 1601
rect 800 1528 846 1567
rect 800 1494 806 1528
rect 840 1494 846 1528
rect 800 1455 846 1494
rect 800 1421 806 1455
rect 840 1421 846 1455
rect 800 1382 846 1421
rect 800 1348 806 1382
rect 840 1348 846 1382
rect 800 1309 846 1348
rect 800 1275 806 1309
rect 840 1275 846 1309
rect 800 1236 846 1275
rect 800 1202 806 1236
rect 840 1202 846 1236
rect 800 1163 846 1202
rect 800 1129 806 1163
rect 840 1129 846 1163
rect 800 1090 846 1129
rect 800 1056 806 1090
rect 840 1056 846 1090
rect 800 1017 846 1056
rect 800 983 806 1017
rect 840 983 846 1017
rect 800 944 846 983
rect 800 910 806 944
rect 840 910 846 944
rect 800 871 846 910
rect 800 837 806 871
rect 840 837 846 871
rect 800 798 846 837
rect 800 764 806 798
rect 840 764 846 798
rect 800 725 846 764
rect 800 691 806 725
rect 840 691 846 725
rect 800 652 846 691
rect 800 618 806 652
rect 840 618 846 652
rect 800 579 846 618
rect 488 534 534 547
rect 800 545 806 579
rect 840 545 846 579
rect 488 533 536 534
tri 536 533 537 534 sw
tri 222 513 237 528 sw
rect 176 508 237 513
tri 237 508 242 513 sw
tri 483 508 488 513 se
rect 488 508 537 533
rect 176 506 242 508
rect 176 472 182 506
rect 216 479 242 506
tri 242 479 271 508 sw
tri 454 479 483 508 se
rect 483 479 494 508
rect 216 474 494 479
rect 528 506 537 508
tri 537 506 564 533 sw
rect 800 506 846 545
rect 528 479 564 506
tri 564 479 591 506 sw
tri 774 479 800 505 se
rect 800 479 806 506
rect 528 474 806 479
rect 216 472 806 474
rect 840 472 846 506
rect 176 435 846 472
rect 176 433 494 435
rect 176 399 182 433
rect 216 401 494 433
rect 528 433 846 435
rect 528 401 806 433
rect 216 399 806 401
rect 840 399 846 433
rect 176 362 846 399
rect 176 361 494 362
rect 176 327 182 361
rect 216 328 494 361
rect 528 361 846 362
rect 528 328 806 361
rect 216 327 806 328
rect 840 327 846 361
rect 176 289 846 327
rect 176 255 182 289
rect 216 255 494 289
rect 528 255 806 289
rect 840 255 846 289
rect 176 243 846 255
rect 228 174 794 186
rect 228 140 240 174
rect 274 140 312 174
rect 346 140 384 174
rect 418 140 456 174
rect 490 140 529 174
rect 563 140 602 174
rect 636 140 675 174
rect 709 140 748 174
rect 782 140 794 174
rect 228 134 794 140
use pfet_CDNS_524688791851505  pfet_CDNS_524688791851505_0
timestamp 1707688321
transform 1 0 227 0 1 220
box -119 -66 687 2066
use PYL1_CDNS_524688791851504  PYL1_CDNS_524688791851504_0
timestamp 1707688321
transform 1 0 240 0 1 122
box 0 0 542 66
use PYL1_CDNS_524688791851504  PYL1_CDNS_524688791851504_1
timestamp 1707688321
transform 1 0 240 0 1 2252
box 0 0 542 66
<< labels >>
flabel comment s 498 1217 498 1217 0 FreeSans 4000 90 0 0 vpb_drvr
flabel metal1 s 423 2019 599 2154 0 FreeSans 200 0 0 0 pad
port 1 nsew
<< properties >>
string GDS_END 90881206
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 90863932
string path 2.075 60.000 2.075 17.800 
<< end >>
