magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -76 -26 10322 1026
<< nmos >>
rect 0 0 36 1000
rect 238 0 274 1000
rect 554 0 590 1000
rect 792 0 828 1000
rect 1108 0 1144 1000
rect 1346 0 1382 1000
rect 1662 0 1698 1000
rect 1900 0 1936 1000
rect 2216 0 2252 1000
rect 2454 0 2490 1000
rect 2770 0 2806 1000
rect 3008 0 3044 1000
rect 3324 0 3360 1000
rect 3562 0 3598 1000
rect 3878 0 3914 1000
rect 4116 0 4152 1000
rect 4432 0 4468 1000
rect 4670 0 4706 1000
rect 4986 0 5022 1000
rect 5224 0 5260 1000
rect 5540 0 5576 1000
rect 5778 0 5814 1000
rect 6094 0 6130 1000
rect 6332 0 6368 1000
rect 6648 0 6684 1000
rect 6886 0 6922 1000
rect 7202 0 7238 1000
rect 7440 0 7476 1000
rect 7756 0 7792 1000
rect 7994 0 8030 1000
rect 8310 0 8346 1000
rect 8548 0 8584 1000
rect 8864 0 8900 1000
rect 9102 0 9138 1000
rect 9418 0 9454 1000
rect 9656 0 9692 1000
rect 9972 0 10008 1000
rect 10210 0 10246 1000
<< ndiff >>
rect -50 0 0 1000
rect 36 0 238 1000
rect 274 0 314 1000
rect 514 0 554 1000
rect 590 0 792 1000
rect 828 0 868 1000
rect 1068 0 1108 1000
rect 1144 0 1346 1000
rect 1382 0 1422 1000
rect 1622 0 1662 1000
rect 1698 0 1900 1000
rect 1936 0 1976 1000
rect 2176 0 2216 1000
rect 2252 0 2454 1000
rect 2490 0 2530 1000
rect 2730 0 2770 1000
rect 2806 0 3008 1000
rect 3044 0 3084 1000
rect 3284 0 3324 1000
rect 3360 0 3562 1000
rect 3598 0 3638 1000
rect 3838 0 3878 1000
rect 3914 0 4116 1000
rect 4152 0 4192 1000
rect 4392 0 4432 1000
rect 4468 0 4670 1000
rect 4706 0 4746 1000
rect 4946 0 4986 1000
rect 5022 0 5224 1000
rect 5260 0 5300 1000
rect 5500 0 5540 1000
rect 5576 0 5778 1000
rect 5814 0 5854 1000
rect 6054 0 6094 1000
rect 6130 0 6332 1000
rect 6368 0 6408 1000
rect 6608 0 6648 1000
rect 6684 0 6886 1000
rect 6922 0 6962 1000
rect 7162 0 7202 1000
rect 7238 0 7440 1000
rect 7476 0 7516 1000
rect 7716 0 7756 1000
rect 7792 0 7994 1000
rect 8030 0 8070 1000
rect 8270 0 8310 1000
rect 8346 0 8548 1000
rect 8584 0 8624 1000
rect 8824 0 8864 1000
rect 8900 0 9102 1000
rect 9138 0 9178 1000
rect 9378 0 9418 1000
rect 9454 0 9656 1000
rect 9692 0 9732 1000
rect 9932 0 9972 1000
rect 10008 0 10210 1000
rect 10246 0 10296 1000
<< poly >>
rect 0 1000 36 1032
rect 238 1000 274 1032
rect 554 1000 590 1032
rect 792 1000 828 1032
rect 1108 1000 1144 1032
rect 1346 1000 1382 1032
rect 1662 1000 1698 1032
rect 1900 1000 1936 1032
rect 2216 1000 2252 1032
rect 2454 1000 2490 1032
rect 2770 1000 2806 1032
rect 3008 1000 3044 1032
rect 3324 1000 3360 1032
rect 3562 1000 3598 1032
rect 3878 1000 3914 1032
rect 4116 1000 4152 1032
rect 4432 1000 4468 1032
rect 4670 1000 4706 1032
rect 4986 1000 5022 1032
rect 5224 1000 5260 1032
rect 5540 1000 5576 1032
rect 5778 1000 5814 1032
rect 6094 1000 6130 1032
rect 6332 1000 6368 1032
rect 6648 1000 6684 1032
rect 6886 1000 6922 1032
rect 7202 1000 7238 1032
rect 7440 1000 7476 1032
rect 7756 1000 7792 1032
rect 7994 1000 8030 1032
rect 8310 1000 8346 1032
rect 8548 1000 8584 1032
rect 8864 1000 8900 1032
rect 9102 1000 9138 1032
rect 9418 1000 9454 1032
rect 9656 1000 9692 1032
rect 9972 1000 10008 1032
rect 10210 1000 10246 1032
rect 0 -32 36 0
rect 238 -32 274 0
rect 554 -32 590 0
rect 792 -32 828 0
rect 1108 -32 1144 0
rect 1346 -32 1382 0
rect 1662 -32 1698 0
rect 1900 -32 1936 0
rect 2216 -32 2252 0
rect 2454 -32 2490 0
rect 2770 -32 2806 0
rect 3008 -32 3044 0
rect 3324 -32 3360 0
rect 3562 -32 3598 0
rect 3878 -32 3914 0
rect 4116 -32 4152 0
rect 4432 -32 4468 0
rect 4670 -32 4706 0
rect 4986 -32 5022 0
rect 5224 -32 5260 0
rect 5540 -32 5576 0
rect 5778 -32 5814 0
rect 6094 -32 6130 0
rect 6332 -32 6368 0
rect 6648 -32 6684 0
rect 6886 -32 6922 0
rect 7202 -32 7238 0
rect 7440 -32 7476 0
rect 7756 -32 7792 0
rect 7994 -32 8030 0
rect 8310 -32 8346 0
rect 8548 -32 8584 0
rect 8864 -32 8900 0
rect 9102 -32 9138 0
rect 9418 -32 9454 0
rect 9656 -32 9692 0
rect 9972 -32 10008 0
rect 10210 -32 10246 0
<< locali >>
rect -229 -4 -51 946
rect 325 -4 503 946
rect 879 -4 1057 946
rect 1433 -4 1611 946
rect 1987 -4 2165 946
rect 2541 -4 2719 946
rect 3095 -4 3273 946
rect 3649 -4 3827 946
rect 4203 -4 4381 946
rect 4757 -4 4935 946
rect 5311 -4 5489 946
rect 5865 -4 6043 946
rect 6419 -4 6597 946
rect 6973 -4 7151 946
rect 7527 -4 7705 946
rect 8081 -4 8259 946
rect 8635 -4 8813 946
rect 9189 -4 9367 946
rect 9743 -4 9921 946
rect 10297 -4 10475 946
use DFTPL1s2_CDNS_55959141808694  DFTPL1s2_CDNS_55959141808694_0
timestamp 1707688321
transform -1 0 -40 0 1 0
box -26 -26 226 1026
use DFTPL1s2_CDNS_55959141808694  DFTPL1s2_CDNS_55959141808694_1
timestamp 1707688321
transform 1 0 314 0 1 0
box -26 -26 226 1026
use DFTPL1s2_CDNS_55959141808694  DFTPL1s2_CDNS_55959141808694_2
timestamp 1707688321
transform 1 0 868 0 1 0
box -26 -26 226 1026
use DFTPL1s2_CDNS_55959141808694  DFTPL1s2_CDNS_55959141808694_3
timestamp 1707688321
transform 1 0 1422 0 1 0
box -26 -26 226 1026
use DFTPL1s2_CDNS_55959141808694  DFTPL1s2_CDNS_55959141808694_4
timestamp 1707688321
transform 1 0 1976 0 1 0
box -26 -26 226 1026
use DFTPL1s2_CDNS_55959141808694  DFTPL1s2_CDNS_55959141808694_5
timestamp 1707688321
transform 1 0 2530 0 1 0
box -26 -26 226 1026
use DFTPL1s2_CDNS_55959141808694  DFTPL1s2_CDNS_55959141808694_6
timestamp 1707688321
transform 1 0 3084 0 1 0
box -26 -26 226 1026
use DFTPL1s2_CDNS_55959141808694  DFTPL1s2_CDNS_55959141808694_7
timestamp 1707688321
transform 1 0 3638 0 1 0
box -26 -26 226 1026
use DFTPL1s2_CDNS_55959141808694  DFTPL1s2_CDNS_55959141808694_8
timestamp 1707688321
transform 1 0 4192 0 1 0
box -26 -26 226 1026
use DFTPL1s2_CDNS_55959141808694  DFTPL1s2_CDNS_55959141808694_9
timestamp 1707688321
transform 1 0 4746 0 1 0
box -26 -26 226 1026
use DFTPL1s2_CDNS_55959141808694  DFTPL1s2_CDNS_55959141808694_10
timestamp 1707688321
transform 1 0 5300 0 1 0
box -26 -26 226 1026
use DFTPL1s2_CDNS_55959141808694  DFTPL1s2_CDNS_55959141808694_11
timestamp 1707688321
transform 1 0 5854 0 1 0
box -26 -26 226 1026
use DFTPL1s2_CDNS_55959141808694  DFTPL1s2_CDNS_55959141808694_12
timestamp 1707688321
transform 1 0 6408 0 1 0
box -26 -26 226 1026
use DFTPL1s2_CDNS_55959141808694  DFTPL1s2_CDNS_55959141808694_13
timestamp 1707688321
transform 1 0 6962 0 1 0
box -26 -26 226 1026
use DFTPL1s2_CDNS_55959141808694  DFTPL1s2_CDNS_55959141808694_14
timestamp 1707688321
transform 1 0 7516 0 1 0
box -26 -26 226 1026
use DFTPL1s2_CDNS_55959141808694  DFTPL1s2_CDNS_55959141808694_15
timestamp 1707688321
transform 1 0 8070 0 1 0
box -26 -26 226 1026
use DFTPL1s2_CDNS_55959141808694  DFTPL1s2_CDNS_55959141808694_16
timestamp 1707688321
transform 1 0 8624 0 1 0
box -26 -26 226 1026
use DFTPL1s2_CDNS_55959141808694  DFTPL1s2_CDNS_55959141808694_17
timestamp 1707688321
transform 1 0 9178 0 1 0
box -26 -26 226 1026
use DFTPL1s2_CDNS_55959141808694  DFTPL1s2_CDNS_55959141808694_18
timestamp 1707688321
transform 1 0 9732 0 1 0
box -26 -26 226 1026
use DFTPL1s2_CDNS_55959141808694  DFTPL1s2_CDNS_55959141808694_19
timestamp 1707688321
transform 1 0 10286 0 1 0
box -26 -26 226 1026
<< labels >>
flabel comment s 10386 471 10386 471 0 FreeSans 300 0 0 0 S
flabel comment s 10109 500 10109 500 0 FreeSans 300 0 0 0 D
flabel comment s 9832 471 9832 471 0 FreeSans 300 0 0 0 S
flabel comment s 9555 500 9555 500 0 FreeSans 300 0 0 0 D
flabel comment s 9278 471 9278 471 0 FreeSans 300 0 0 0 S
flabel comment s 9001 500 9001 500 0 FreeSans 300 0 0 0 D
flabel comment s 8724 471 8724 471 0 FreeSans 300 0 0 0 S
flabel comment s 8447 500 8447 500 0 FreeSans 300 0 0 0 D
flabel comment s 8170 471 8170 471 0 FreeSans 300 0 0 0 S
flabel comment s 7893 500 7893 500 0 FreeSans 300 0 0 0 D
flabel comment s 7616 471 7616 471 0 FreeSans 300 0 0 0 S
flabel comment s 7339 500 7339 500 0 FreeSans 300 0 0 0 D
flabel comment s 7062 471 7062 471 0 FreeSans 300 0 0 0 S
flabel comment s 6785 500 6785 500 0 FreeSans 300 0 0 0 D
flabel comment s 6508 471 6508 471 0 FreeSans 300 0 0 0 S
flabel comment s 6231 500 6231 500 0 FreeSans 300 0 0 0 D
flabel comment s 5954 471 5954 471 0 FreeSans 300 0 0 0 S
flabel comment s 5677 500 5677 500 0 FreeSans 300 0 0 0 D
flabel comment s 5400 471 5400 471 0 FreeSans 300 0 0 0 S
flabel comment s 5123 500 5123 500 0 FreeSans 300 0 0 0 D
flabel comment s 4846 471 4846 471 0 FreeSans 300 0 0 0 S
flabel comment s 4569 500 4569 500 0 FreeSans 300 0 0 0 D
flabel comment s 4292 471 4292 471 0 FreeSans 300 0 0 0 S
flabel comment s 4015 500 4015 500 0 FreeSans 300 0 0 0 D
flabel comment s 3738 471 3738 471 0 FreeSans 300 0 0 0 S
flabel comment s 3461 500 3461 500 0 FreeSans 300 0 0 0 D
flabel comment s 3184 471 3184 471 0 FreeSans 300 0 0 0 S
flabel comment s 2907 500 2907 500 0 FreeSans 300 0 0 0 D
flabel comment s 2630 471 2630 471 0 FreeSans 300 0 0 0 S
flabel comment s 2353 500 2353 500 0 FreeSans 300 0 0 0 D
flabel comment s 2076 471 2076 471 0 FreeSans 300 0 0 0 S
flabel comment s 1799 500 1799 500 0 FreeSans 300 0 0 0 D
flabel comment s 1522 471 1522 471 0 FreeSans 300 0 0 0 S
flabel comment s 1245 500 1245 500 0 FreeSans 300 0 0 0 D
flabel comment s 968 471 968 471 0 FreeSans 300 0 0 0 S
flabel comment s 691 500 691 500 0 FreeSans 300 0 0 0 D
flabel comment s 414 471 414 471 0 FreeSans 300 0 0 0 S
flabel comment s 137 500 137 500 0 FreeSans 300 0 0 0 D
flabel comment s -140 471 -140 471 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 42998392
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 42978912
<< end >>
