magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -76 -26 1676 226
<< mvnmos >>
rect 0 0 1600 200
<< mvndiff >>
rect -50 0 0 200
rect 1600 0 1650 200
<< poly >>
rect 0 200 1600 232
rect 0 -32 1600 0
<< metal1 >>
rect -51 -16 -5 186
rect 1605 -16 1651 186
use hvDFM1sd2_CDNS_52468879185104  hvDFM1sd2_CDNS_52468879185104_0
timestamp 1707688321
transform -1 0 0 0 1 0
box -26 -26 82 226
use hvDFM1sd2_CDNS_52468879185104  hvDFM1sd2_CDNS_52468879185104_1
timestamp 1707688321
transform 1 0 1600 0 1 0
box -26 -26 82 226
<< labels >>
flabel comment s -28 85 -28 85 0 FreeSans 300 0 0 0 S
flabel comment s 1628 85 1628 85 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 6110274
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 6109380
<< end >>
