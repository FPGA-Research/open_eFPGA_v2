magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< metal3 >>
rect 7582 7551 9707 7592
rect 7582 7007 7612 7551
rect 9676 7007 9707 7551
rect 7582 6966 9707 7007
rect 5196 3198 7321 3242
rect 5196 2654 5226 3198
rect 7290 2654 7321 3198
rect 5196 2610 7321 2654
<< via3 >>
rect 7612 7007 9676 7551
rect 5226 2654 7290 3198
<< metal4 >>
rect 7582 7551 9707 7592
rect 7582 7007 7612 7551
rect 9676 7007 9707 7551
rect 7582 6966 9707 7007
rect 5196 3198 7321 3242
rect 5196 2654 5226 3198
rect 7290 2654 7321 3198
rect 5196 2610 7321 2654
<< properties >>
string FIXED_BBOX 0 -406 15000 39593
string GDS_END 3034516
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io.gds
string GDS_START 3010896
<< end >>
