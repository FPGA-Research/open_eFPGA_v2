magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 821 157 1195 203
rect 1 21 1195 157
rect 29 -17 63 21
<< locali >>
rect 17 197 65 325
rect 287 191 353 265
rect 1127 334 1179 491
rect 949 199 1015 265
rect 949 69 995 199
rect 1145 149 1179 334
rect 1122 69 1179 149
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 17 393 69 493
rect 103 427 169 527
rect 17 359 155 393
rect 121 280 155 359
rect 203 337 247 493
rect 121 214 167 280
rect 121 161 155 214
rect 34 127 155 161
rect 34 69 69 127
rect 103 17 169 93
rect 203 69 237 337
rect 286 333 357 483
rect 391 367 449 527
rect 562 451 725 485
rect 580 357 653 399
rect 286 299 423 333
rect 389 219 423 299
rect 489 325 552 337
rect 601 327 653 357
rect 489 271 567 325
rect 601 219 649 327
rect 691 265 725 451
rect 786 427 889 527
rect 925 373 993 487
rect 1027 383 1093 527
rect 763 347 993 373
rect 763 307 1093 347
rect 869 301 1093 307
rect 691 233 835 265
rect 389 157 467 219
rect 302 153 467 157
rect 538 153 649 219
rect 683 199 835 233
rect 302 123 423 153
rect 302 69 341 123
rect 683 107 717 199
rect 869 161 915 301
rect 1049 265 1093 301
rect 375 17 441 89
rect 563 73 717 107
rect 751 17 805 122
rect 839 59 915 161
rect 1049 199 1111 265
rect 1031 17 1088 143
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< obsm1 >>
rect 201 388 259 397
rect 573 388 631 397
rect 201 360 631 388
rect 201 351 259 360
rect 573 351 631 360
rect 109 320 167 329
rect 477 320 535 329
rect 109 292 535 320
rect 109 283 167 292
rect 477 283 535 292
<< labels >>
rlabel locali s 287 191 353 265 6 D
port 1 nsew signal input
rlabel locali s 17 197 65 325 6 GATE
port 2 nsew clock input
rlabel locali s 949 69 995 199 6 RESET_B
port 3 nsew signal input
rlabel locali s 949 199 1015 265 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 0 -48 1196 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 1195 157 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 821 157 1195 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 1234 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 1196 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1122 69 1179 149 6 Q
port 8 nsew signal output
rlabel locali s 1145 149 1179 334 6 Q
port 8 nsew signal output
rlabel locali s 1127 334 1179 491 6 Q
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1196 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2771482
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2760744
<< end >>
