magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -210 30 2206 2082
<< mvnnmos >>
tri 578 2036 598 2056 ne
tri 578 56 598 76 se
rect 598 56 1398 2056
tri 1398 2036 1418 2056 nw
tri 1398 56 1418 76 sw
<< ndiff >>
rect -184 1957 -20 2056
rect -184 1923 -44 1957
rect -184 1889 -20 1923
rect -184 1855 -44 1889
rect -184 1821 -20 1855
rect -184 1787 -44 1821
rect -184 1753 -20 1787
rect -184 1719 -44 1753
rect -184 1685 -20 1719
rect -184 1651 -44 1685
rect -184 1617 -20 1651
rect -184 1583 -44 1617
rect -184 1549 -20 1583
rect -184 1515 -44 1549
rect -184 1481 -20 1515
rect -184 1447 -44 1481
rect -184 1413 -20 1447
rect -184 1379 -44 1413
rect -184 1345 -20 1379
rect -184 1311 -44 1345
rect -184 1277 -20 1311
rect -184 1243 -44 1277
rect -184 1209 -20 1243
rect -184 1175 -44 1209
rect -184 1141 -20 1175
rect -184 1107 -44 1141
rect -184 1073 -20 1107
rect -184 1039 -44 1073
rect -184 1005 -20 1039
rect -184 971 -44 1005
rect -184 937 -20 971
rect -184 903 -44 937
rect -184 869 -20 903
rect -184 835 -44 869
rect -184 801 -20 835
rect -184 767 -44 801
rect -184 733 -20 767
rect -184 699 -44 733
rect -184 665 -20 699
rect -184 631 -44 665
rect -184 597 -20 631
rect -184 563 -44 597
rect -184 529 -20 563
rect -184 495 -44 529
rect -184 461 -20 495
rect -184 427 -44 461
rect -184 393 -20 427
rect -184 359 -44 393
rect -184 325 -20 359
rect -184 291 -44 325
rect -184 257 -20 291
rect -184 223 -44 257
rect -184 189 -20 223
rect -184 155 -44 189
rect -184 56 -20 155
rect 1736 1957 2180 2056
rect 1736 155 1938 1957
rect 2040 155 2180 1957
rect 1736 56 2180 155
<< mvndiff >>
rect -20 2036 578 2056
tri 578 2036 598 2056 sw
rect -20 1957 598 2036
rect 58 155 598 1957
rect -20 76 598 155
rect -20 56 578 76
tri 578 56 598 76 nw
tri 1398 2036 1418 2056 se
rect 1418 2036 1736 2056
rect 1398 76 1736 2036
tri 1398 56 1418 76 ne
rect 1418 56 1736 76
<< ndiffc >>
rect -44 1923 -20 1957
rect -44 1855 -20 1889
rect -44 1787 -20 1821
rect -44 1719 -20 1753
rect -44 1651 -20 1685
rect -44 1583 -20 1617
rect -44 1515 -20 1549
rect -44 1447 -20 1481
rect -44 1379 -20 1413
rect -44 1311 -20 1345
rect -44 1243 -20 1277
rect -44 1175 -20 1209
rect -44 1107 -20 1141
rect -44 1039 -20 1073
rect -44 971 -20 1005
rect -44 903 -20 937
rect -44 835 -20 869
rect -44 767 -20 801
rect -44 699 -20 733
rect -44 631 -20 665
rect -44 563 -20 597
rect -44 495 -20 529
rect -44 427 -20 461
rect -44 359 -20 393
rect -44 291 -20 325
rect -44 223 -20 257
rect -44 155 -20 189
rect 1938 155 2040 1957
<< mvndiffc >>
rect -20 155 58 1957
<< poly >>
rect 558 2183 1438 2199
rect 558 2149 574 2183
rect 608 2149 648 2183
rect 682 2149 722 2183
rect 756 2149 796 2183
rect 830 2149 870 2183
rect 904 2149 944 2183
rect 978 2149 1018 2183
rect 1052 2149 1092 2183
rect 1126 2149 1166 2183
rect 1200 2149 1240 2183
rect 1274 2149 1314 2183
rect 1348 2149 1388 2183
rect 1422 2149 1438 2183
rect 558 2076 1438 2149
tri 558 2056 578 2076 ne
rect 578 2056 1418 2076
tri 1418 2056 1438 2076 nw
tri 558 36 578 56 se
rect 578 36 1418 56
tri 1418 36 1438 56 sw
rect 558 -87 1438 36
<< polycont >>
rect 574 2149 608 2183
rect 648 2149 682 2183
rect 722 2149 756 2183
rect 796 2149 830 2183
rect 870 2149 904 2183
rect 944 2149 978 2183
rect 1018 2149 1052 2183
rect 1092 2149 1126 2183
rect 1166 2149 1200 2183
rect 1240 2149 1274 2183
rect 1314 2149 1348 2183
rect 1388 2149 1422 2183
<< locali >>
rect 558 2149 574 2183
rect 608 2149 648 2183
rect 682 2149 722 2183
rect 756 2149 796 2183
rect 830 2149 870 2183
rect 904 2149 944 2183
rect 978 2149 1018 2183
rect 1052 2149 1092 2183
rect 1126 2149 1166 2183
rect 1200 2149 1240 2183
rect 1274 2149 1314 2183
rect 1348 2149 1388 2183
rect 1422 2149 1438 2183
rect -236 1957 307 2056
rect -236 1923 -46 1957
rect 60 1923 307 1957
rect -236 1889 -20 1923
rect -236 1884 -44 1889
rect 58 1884 307 1923
rect -236 1850 -46 1884
rect 60 1850 307 1884
rect -236 1821 -20 1850
rect -236 1811 -44 1821
rect 58 1811 307 1850
rect -236 1777 -46 1811
rect 60 1777 307 1811
rect -236 1753 -20 1777
rect -236 1738 -44 1753
rect 58 1738 307 1777
rect -236 1704 -46 1738
rect 60 1704 307 1738
rect -236 1685 -20 1704
rect -236 1665 -44 1685
rect 58 1665 307 1704
rect -236 1631 -46 1665
rect 60 1631 307 1665
rect -236 1617 -20 1631
rect -236 1592 -44 1617
rect 58 1592 307 1631
rect -236 1558 -46 1592
rect 60 1558 307 1592
rect -236 1549 -20 1558
rect -236 1519 -44 1549
rect 58 1519 307 1558
rect -236 1485 -46 1519
rect 60 1485 307 1519
rect -236 1481 -20 1485
rect -236 1447 -44 1481
rect -236 1446 -20 1447
rect 58 1446 307 1485
rect -236 1412 -46 1446
rect 60 1412 307 1446
rect -236 1379 -44 1412
rect -236 1373 -20 1379
rect 58 1373 307 1412
rect -236 1339 -46 1373
rect 60 1339 307 1373
rect -236 1311 -44 1339
rect -236 1299 -20 1311
rect 58 1299 307 1339
rect -236 1265 -46 1299
rect 60 1265 307 1299
rect -236 1243 -44 1265
rect -236 1225 -20 1243
rect 58 1225 307 1265
rect -236 1191 -46 1225
rect 60 1191 307 1225
rect -236 1175 -44 1191
rect -236 1151 -20 1175
rect 58 1151 307 1191
rect -236 1117 -46 1151
rect 60 1117 307 1151
rect -236 1107 -44 1117
rect -236 1077 -20 1107
rect 58 1077 307 1117
rect -236 1043 -46 1077
rect 60 1043 307 1077
rect -236 1039 -44 1043
rect -236 1005 -20 1039
rect -236 1003 -44 1005
rect 58 1003 307 1043
rect -236 969 -46 1003
rect 60 969 307 1003
rect -236 937 -20 969
rect -236 929 -44 937
rect 58 929 307 969
rect -236 895 -46 929
rect 60 895 307 929
rect -236 869 -20 895
rect -236 855 -44 869
rect 58 855 307 895
rect -236 821 -46 855
rect 60 821 307 855
rect -236 801 -20 821
rect -236 781 -44 801
rect 58 781 307 821
rect -236 747 -46 781
rect 60 747 307 781
rect -236 733 -20 747
rect -236 707 -44 733
rect 58 707 307 747
rect -236 673 -46 707
rect 60 673 307 707
rect -236 665 -20 673
rect -236 633 -44 665
rect 58 633 307 673
rect -236 599 -46 633
rect 60 599 307 633
rect -236 597 -20 599
rect -236 563 -44 597
rect -236 559 -20 563
rect 58 559 307 599
rect -236 525 -46 559
rect 60 525 307 559
rect -236 495 -44 525
rect -236 485 -20 495
rect 58 485 307 525
rect -236 451 -46 485
rect 60 451 307 485
rect -236 427 -44 451
rect -236 411 -20 427
rect 58 411 307 451
rect -236 377 -46 411
rect 60 377 307 411
rect -236 359 -44 377
rect -236 337 -20 359
rect 58 337 307 377
rect -236 303 -46 337
rect 60 303 307 337
rect -236 291 -44 303
rect -236 263 -20 291
rect 58 263 307 303
rect -236 229 -46 263
rect 60 229 307 263
rect -236 223 -44 229
rect -236 189 -20 223
rect 58 189 307 229
rect -236 155 -46 189
rect 60 155 307 189
rect -236 56 307 155
rect 1689 1957 2232 2056
rect 1689 1923 1936 1957
rect 2042 1923 2232 1957
rect 1689 1884 1938 1923
rect 2040 1884 2232 1923
rect 1689 1850 1936 1884
rect 2042 1850 2232 1884
rect 1689 1811 1938 1850
rect 2040 1811 2232 1850
rect 1689 1777 1936 1811
rect 2042 1777 2232 1811
rect 1689 1738 1938 1777
rect 2040 1738 2232 1777
rect 1689 1704 1936 1738
rect 2042 1704 2232 1738
rect 1689 1665 1938 1704
rect 2040 1665 2232 1704
rect 1689 1631 1936 1665
rect 2042 1631 2232 1665
rect 1689 1592 1938 1631
rect 2040 1592 2232 1631
rect 1689 1558 1936 1592
rect 2042 1558 2232 1592
rect 1689 1519 1938 1558
rect 2040 1519 2232 1558
rect 1689 1485 1936 1519
rect 2042 1485 2232 1519
rect 1689 1446 1938 1485
rect 2040 1446 2232 1485
rect 1689 1412 1936 1446
rect 2042 1412 2232 1446
rect 1689 1373 1938 1412
rect 2040 1373 2232 1412
rect 1689 1339 1936 1373
rect 2042 1339 2232 1373
rect 1689 1299 1938 1339
rect 2040 1299 2232 1339
rect 1689 1265 1936 1299
rect 2042 1265 2232 1299
rect 1689 1225 1938 1265
rect 2040 1225 2232 1265
rect 1689 1191 1936 1225
rect 2042 1191 2232 1225
rect 1689 1151 1938 1191
rect 2040 1151 2232 1191
rect 1689 1117 1936 1151
rect 2042 1117 2232 1151
rect 1689 1077 1938 1117
rect 2040 1077 2232 1117
rect 1689 1043 1936 1077
rect 2042 1043 2232 1077
rect 1689 1003 1938 1043
rect 2040 1003 2232 1043
rect 1689 969 1936 1003
rect 2042 969 2232 1003
rect 1689 929 1938 969
rect 2040 929 2232 969
rect 1689 895 1936 929
rect 2042 895 2232 929
rect 1689 855 1938 895
rect 2040 855 2232 895
rect 1689 821 1936 855
rect 2042 821 2232 855
rect 1689 781 1938 821
rect 2040 781 2232 821
rect 1689 747 1936 781
rect 2042 747 2232 781
rect 1689 707 1938 747
rect 2040 707 2232 747
rect 1689 673 1936 707
rect 2042 673 2232 707
rect 1689 633 1938 673
rect 2040 633 2232 673
rect 1689 599 1936 633
rect 2042 599 2232 633
rect 1689 559 1938 599
rect 2040 559 2232 599
rect 1689 525 1936 559
rect 2042 525 2232 559
rect 1689 485 1938 525
rect 2040 485 2232 525
rect 1689 451 1936 485
rect 2042 451 2232 485
rect 1689 411 1938 451
rect 2040 411 2232 451
rect 1689 377 1936 411
rect 2042 377 2232 411
rect 1689 337 1938 377
rect 2040 337 2232 377
rect 1689 303 1936 337
rect 2042 303 2232 337
rect 1689 263 1938 303
rect 2040 263 2232 303
rect 1689 229 1936 263
rect 2042 229 2232 263
rect 1689 189 1938 229
rect 2040 189 2232 229
rect 1689 155 1936 189
rect 2042 155 2232 189
rect 1689 56 2232 155
<< viali >>
rect -46 1923 -44 1957
rect -44 1923 -20 1957
rect -20 1923 -12 1957
rect 26 1923 58 1957
rect 58 1923 60 1957
rect -46 1855 -44 1884
rect -44 1855 -20 1884
rect -46 1850 -20 1855
rect -20 1850 -12 1884
rect 26 1850 58 1884
rect 58 1850 60 1884
rect -46 1787 -44 1811
rect -44 1787 -20 1811
rect -46 1777 -20 1787
rect -20 1777 -12 1811
rect 26 1777 58 1811
rect 58 1777 60 1811
rect -46 1719 -44 1738
rect -44 1719 -20 1738
rect -46 1704 -20 1719
rect -20 1704 -12 1738
rect 26 1704 58 1738
rect 58 1704 60 1738
rect -46 1651 -44 1665
rect -44 1651 -20 1665
rect -46 1631 -20 1651
rect -20 1631 -12 1665
rect 26 1631 58 1665
rect 58 1631 60 1665
rect -46 1583 -44 1592
rect -44 1583 -20 1592
rect -46 1558 -20 1583
rect -20 1558 -12 1592
rect 26 1558 58 1592
rect 58 1558 60 1592
rect -46 1515 -44 1519
rect -44 1515 -20 1519
rect -46 1485 -20 1515
rect -20 1485 -12 1519
rect 26 1485 58 1519
rect 58 1485 60 1519
rect -46 1413 -20 1446
rect -46 1412 -44 1413
rect -44 1412 -20 1413
rect -20 1412 -12 1446
rect 26 1412 58 1446
rect 58 1412 60 1446
rect -46 1345 -20 1373
rect -46 1339 -44 1345
rect -44 1339 -20 1345
rect -20 1339 -12 1373
rect 26 1339 58 1373
rect 58 1339 60 1373
rect -46 1277 -20 1299
rect -46 1265 -44 1277
rect -44 1265 -20 1277
rect -20 1265 -12 1299
rect 26 1265 58 1299
rect 58 1265 60 1299
rect -46 1209 -20 1225
rect -46 1191 -44 1209
rect -44 1191 -20 1209
rect -20 1191 -12 1225
rect 26 1191 58 1225
rect 58 1191 60 1225
rect -46 1141 -20 1151
rect -46 1117 -44 1141
rect -44 1117 -20 1141
rect -20 1117 -12 1151
rect 26 1117 58 1151
rect 58 1117 60 1151
rect -46 1073 -20 1077
rect -46 1043 -44 1073
rect -44 1043 -20 1073
rect -20 1043 -12 1077
rect 26 1043 58 1077
rect 58 1043 60 1077
rect -46 971 -44 1003
rect -44 971 -20 1003
rect -46 969 -20 971
rect -20 969 -12 1003
rect 26 969 58 1003
rect 58 969 60 1003
rect -46 903 -44 929
rect -44 903 -20 929
rect -46 895 -20 903
rect -20 895 -12 929
rect 26 895 58 929
rect 58 895 60 929
rect -46 835 -44 855
rect -44 835 -20 855
rect -46 821 -20 835
rect -20 821 -12 855
rect 26 821 58 855
rect 58 821 60 855
rect -46 767 -44 781
rect -44 767 -20 781
rect -46 747 -20 767
rect -20 747 -12 781
rect 26 747 58 781
rect 58 747 60 781
rect -46 699 -44 707
rect -44 699 -20 707
rect -46 673 -20 699
rect -20 673 -12 707
rect 26 673 58 707
rect 58 673 60 707
rect -46 631 -44 633
rect -44 631 -20 633
rect -46 599 -20 631
rect -20 599 -12 633
rect 26 599 58 633
rect 58 599 60 633
rect -46 529 -20 559
rect -46 525 -44 529
rect -44 525 -20 529
rect -20 525 -12 559
rect 26 525 58 559
rect 58 525 60 559
rect -46 461 -20 485
rect -46 451 -44 461
rect -44 451 -20 461
rect -20 451 -12 485
rect 26 451 58 485
rect 58 451 60 485
rect -46 393 -20 411
rect -46 377 -44 393
rect -44 377 -20 393
rect -20 377 -12 411
rect 26 377 58 411
rect 58 377 60 411
rect -46 325 -20 337
rect -46 303 -44 325
rect -44 303 -20 325
rect -20 303 -12 337
rect 26 303 58 337
rect 58 303 60 337
rect -46 257 -20 263
rect -46 229 -44 257
rect -44 229 -20 257
rect -20 229 -12 263
rect 26 229 58 263
rect 58 229 60 263
rect -46 155 -44 189
rect -44 155 -20 189
rect -20 155 -12 189
rect 26 155 58 189
rect 58 155 60 189
rect 1936 1923 1938 1957
rect 1938 1923 1970 1957
rect 2008 1923 2040 1957
rect 2040 1923 2042 1957
rect 1936 1850 1938 1884
rect 1938 1850 1970 1884
rect 2008 1850 2040 1884
rect 2040 1850 2042 1884
rect 1936 1777 1938 1811
rect 1938 1777 1970 1811
rect 2008 1777 2040 1811
rect 2040 1777 2042 1811
rect 1936 1704 1938 1738
rect 1938 1704 1970 1738
rect 2008 1704 2040 1738
rect 2040 1704 2042 1738
rect 1936 1631 1938 1665
rect 1938 1631 1970 1665
rect 2008 1631 2040 1665
rect 2040 1631 2042 1665
rect 1936 1558 1938 1592
rect 1938 1558 1970 1592
rect 2008 1558 2040 1592
rect 2040 1558 2042 1592
rect 1936 1485 1938 1519
rect 1938 1485 1970 1519
rect 2008 1485 2040 1519
rect 2040 1485 2042 1519
rect 1936 1412 1938 1446
rect 1938 1412 1970 1446
rect 2008 1412 2040 1446
rect 2040 1412 2042 1446
rect 1936 1339 1938 1373
rect 1938 1339 1970 1373
rect 2008 1339 2040 1373
rect 2040 1339 2042 1373
rect 1936 1265 1938 1299
rect 1938 1265 1970 1299
rect 2008 1265 2040 1299
rect 2040 1265 2042 1299
rect 1936 1191 1938 1225
rect 1938 1191 1970 1225
rect 2008 1191 2040 1225
rect 2040 1191 2042 1225
rect 1936 1117 1938 1151
rect 1938 1117 1970 1151
rect 2008 1117 2040 1151
rect 2040 1117 2042 1151
rect 1936 1043 1938 1077
rect 1938 1043 1970 1077
rect 2008 1043 2040 1077
rect 2040 1043 2042 1077
rect 1936 969 1938 1003
rect 1938 969 1970 1003
rect 2008 969 2040 1003
rect 2040 969 2042 1003
rect 1936 895 1938 929
rect 1938 895 1970 929
rect 2008 895 2040 929
rect 2040 895 2042 929
rect 1936 821 1938 855
rect 1938 821 1970 855
rect 2008 821 2040 855
rect 2040 821 2042 855
rect 1936 747 1938 781
rect 1938 747 1970 781
rect 2008 747 2040 781
rect 2040 747 2042 781
rect 1936 673 1938 707
rect 1938 673 1970 707
rect 2008 673 2040 707
rect 2040 673 2042 707
rect 1936 599 1938 633
rect 1938 599 1970 633
rect 2008 599 2040 633
rect 2040 599 2042 633
rect 1936 525 1938 559
rect 1938 525 1970 559
rect 2008 525 2040 559
rect 2040 525 2042 559
rect 1936 451 1938 485
rect 1938 451 1970 485
rect 2008 451 2040 485
rect 2040 451 2042 485
rect 1936 377 1938 411
rect 1938 377 1970 411
rect 2008 377 2040 411
rect 2040 377 2042 411
rect 1936 303 1938 337
rect 1938 303 1970 337
rect 2008 303 2040 337
rect 2040 303 2042 337
rect 1936 229 1938 263
rect 1938 229 1970 263
rect 2008 229 2040 263
rect 2040 229 2042 263
rect 1936 155 1938 189
rect 1938 155 1970 189
rect 2008 155 2040 189
rect 2040 155 2042 189
<< metal1 >>
tri -269 2056 -222 2103 se
rect -222 2056 236 2103
tri 236 2056 283 2103 sw
rect -269 1957 283 2056
rect -269 1923 -46 1957
rect -12 1923 26 1957
rect 60 1923 283 1957
rect -269 1884 283 1923
rect -269 1850 -46 1884
rect -12 1850 26 1884
rect 60 1850 283 1884
rect -269 1811 283 1850
rect -269 1777 -46 1811
rect -12 1777 26 1811
rect 60 1777 283 1811
rect -269 1738 283 1777
rect -269 1704 -46 1738
rect -12 1704 26 1738
rect 60 1704 283 1738
rect -269 1665 283 1704
rect -269 1631 -46 1665
rect -12 1631 26 1665
rect 60 1631 283 1665
rect -269 1592 283 1631
rect -269 1558 -46 1592
rect -12 1558 26 1592
rect 60 1558 283 1592
rect -269 1519 283 1558
rect -269 1485 -46 1519
rect -12 1485 26 1519
rect 60 1485 283 1519
rect -269 1446 283 1485
rect -269 1412 -46 1446
rect -12 1412 26 1446
rect 60 1412 283 1446
rect -269 1373 283 1412
rect -269 1339 -46 1373
rect -12 1339 26 1373
rect 60 1339 283 1373
rect -269 1299 283 1339
rect -269 1265 -46 1299
rect -12 1265 26 1299
rect 60 1265 283 1299
rect -269 1225 283 1265
rect -269 1191 -46 1225
rect -12 1191 26 1225
rect 60 1191 283 1225
rect -269 1151 283 1191
rect -269 1117 -46 1151
rect -12 1117 26 1151
rect 60 1117 283 1151
rect -269 1077 283 1117
rect -269 1043 -46 1077
rect -12 1043 26 1077
rect 60 1043 283 1077
rect -269 1003 283 1043
rect -269 969 -46 1003
rect -12 969 26 1003
rect 60 969 283 1003
rect -269 929 283 969
rect -269 895 -46 929
rect -12 895 26 929
rect 60 895 283 929
rect -269 855 283 895
rect -269 821 -46 855
rect -12 821 26 855
rect 60 821 283 855
rect -269 781 283 821
rect -269 747 -46 781
rect -12 747 26 781
rect 60 747 283 781
rect -269 707 283 747
rect -269 673 -46 707
rect -12 673 26 707
rect 60 673 283 707
rect -269 633 283 673
rect -269 599 -46 633
rect -12 599 26 633
rect 60 599 283 633
rect -269 559 283 599
rect -269 525 -46 559
rect -12 525 26 559
rect 60 525 283 559
rect -269 485 283 525
rect -269 451 -46 485
rect -12 451 26 485
rect 60 451 283 485
rect -269 411 283 451
rect -269 377 -46 411
rect -12 377 26 411
rect 60 377 283 411
rect -269 337 283 377
rect -269 303 -46 337
rect -12 303 26 337
rect 60 303 283 337
rect -269 263 283 303
rect -269 229 -46 263
rect -12 229 26 263
rect 60 229 283 263
rect -269 189 283 229
rect -269 155 -46 189
rect -12 155 26 189
rect 60 155 283 189
rect -269 56 283 155
tri -269 9 -222 56 ne
rect -222 9 236 56
tri 236 9 283 56 nw
tri 1713 2056 1760 2103 se
rect 1760 2056 2218 2103
tri 2218 2056 2265 2103 sw
rect 1713 1957 2265 2056
rect 1713 1923 1936 1957
rect 1970 1923 2008 1957
rect 2042 1923 2265 1957
rect 1713 1884 2265 1923
rect 1713 1850 1936 1884
rect 1970 1850 2008 1884
rect 2042 1850 2265 1884
rect 1713 1811 2265 1850
rect 1713 1777 1936 1811
rect 1970 1777 2008 1811
rect 2042 1777 2265 1811
rect 1713 1738 2265 1777
rect 1713 1704 1936 1738
rect 1970 1704 2008 1738
rect 2042 1704 2265 1738
rect 1713 1665 2265 1704
rect 1713 1631 1936 1665
rect 1970 1631 2008 1665
rect 2042 1631 2265 1665
rect 1713 1592 2265 1631
rect 1713 1558 1936 1592
rect 1970 1558 2008 1592
rect 2042 1558 2265 1592
rect 1713 1519 2265 1558
rect 1713 1485 1936 1519
rect 1970 1485 2008 1519
rect 2042 1485 2265 1519
rect 1713 1446 2265 1485
rect 1713 1412 1936 1446
rect 1970 1412 2008 1446
rect 2042 1412 2265 1446
rect 1713 1373 2265 1412
rect 1713 1339 1936 1373
rect 1970 1339 2008 1373
rect 2042 1339 2265 1373
rect 1713 1299 2265 1339
rect 1713 1265 1936 1299
rect 1970 1265 2008 1299
rect 2042 1265 2265 1299
rect 1713 1225 2265 1265
rect 1713 1191 1936 1225
rect 1970 1191 2008 1225
rect 2042 1191 2265 1225
rect 1713 1151 2265 1191
rect 1713 1117 1936 1151
rect 1970 1117 2008 1151
rect 2042 1117 2265 1151
rect 1713 1077 2265 1117
rect 1713 1043 1936 1077
rect 1970 1043 2008 1077
rect 2042 1043 2265 1077
rect 1713 1003 2265 1043
rect 1713 969 1936 1003
rect 1970 969 2008 1003
rect 2042 969 2265 1003
rect 1713 929 2265 969
rect 1713 895 1936 929
rect 1970 895 2008 929
rect 2042 895 2265 929
rect 1713 855 2265 895
rect 1713 821 1936 855
rect 1970 821 2008 855
rect 2042 821 2265 855
rect 1713 781 2265 821
rect 1713 747 1936 781
rect 1970 747 2008 781
rect 2042 747 2265 781
rect 1713 707 2265 747
rect 1713 673 1936 707
rect 1970 673 2008 707
rect 2042 673 2265 707
rect 1713 633 2265 673
rect 1713 599 1936 633
rect 1970 599 2008 633
rect 2042 599 2265 633
rect 1713 559 2265 599
rect 1713 525 1936 559
rect 1970 525 2008 559
rect 2042 525 2265 559
rect 1713 485 2265 525
rect 1713 451 1936 485
rect 1970 451 2008 485
rect 2042 451 2265 485
rect 1713 411 2265 451
rect 1713 377 1936 411
rect 1970 377 2008 411
rect 2042 377 2265 411
rect 1713 337 2265 377
rect 1713 303 1936 337
rect 1970 303 2008 337
rect 2042 303 2265 337
rect 1713 263 2265 303
rect 1713 229 1936 263
rect 1970 229 2008 263
rect 2042 229 2265 263
rect 1713 189 2265 229
rect 1713 155 1936 189
rect 1970 155 2008 189
rect 2042 155 2265 189
rect 1713 56 2265 155
tri 1713 9 1760 56 ne
rect 1760 9 2218 56
tri 2218 9 2265 56 nw
<< labels >>
flabel comment s 1955 1037 1955 1037 0 FreeSans 300 180 0 0 S
flabel comment s 41 1037 41 1037 0 FreeSans 300 180 0 0 D
<< properties >>
string GDS_END 94762914
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 94747472
string path 0.175 3.575 0.175 49.225 
<< end >>
