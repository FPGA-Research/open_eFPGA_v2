magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -76 -26 2360 1426
<< mvnmos >>
rect 0 0 100 1400
rect 156 0 256 1400
rect 312 0 412 1400
rect 468 0 568 1400
rect 624 0 724 1400
rect 780 0 880 1400
rect 936 0 1036 1400
rect 1092 0 1192 1400
rect 1248 0 1348 1400
rect 1404 0 1504 1400
rect 1560 0 1660 1400
rect 1716 0 1816 1400
rect 1872 0 1972 1400
rect 2028 0 2128 1400
rect 2184 0 2284 1400
<< mvndiff >>
rect -50 0 0 1400
rect 2284 0 2334 1400
<< poly >>
rect 0 1400 100 1426
rect 0 -26 100 0
rect 156 1400 256 1426
rect 156 -26 256 0
rect 312 1400 412 1426
rect 312 -26 412 0
rect 468 1400 568 1426
rect 468 -26 568 0
rect 624 1400 724 1426
rect 624 -26 724 0
rect 780 1400 880 1426
rect 780 -26 880 0
rect 936 1400 1036 1426
rect 936 -26 1036 0
rect 1092 1400 1192 1426
rect 1092 -26 1192 0
rect 1248 1400 1348 1426
rect 1248 -26 1348 0
rect 1404 1400 1504 1426
rect 1404 -26 1504 0
rect 1560 1400 1660 1426
rect 1560 -26 1660 0
rect 1716 1400 1816 1426
rect 1716 -26 1816 0
rect 1872 1400 1972 1426
rect 1872 -26 1972 0
rect 2028 1400 2128 1426
rect 2028 -26 2128 0
rect 2184 1400 2284 1426
rect 2184 -26 2284 0
<< locali >>
rect -45 -4 -11 1354
rect 111 -4 145 1354
rect 267 -4 301 1354
rect 423 -4 457 1354
rect 579 -4 613 1354
rect 735 -4 769 1354
rect 891 -4 925 1354
rect 1047 -4 1081 1354
rect 1203 -4 1237 1354
rect 1359 -4 1393 1354
rect 1515 -4 1549 1354
rect 1671 -4 1705 1354
rect 1827 -4 1861 1354
rect 1983 -4 2017 1354
rect 2139 -4 2173 1354
rect 2295 -4 2329 1354
use DFL1sd2_CDNS_52468879185839  DFL1sd2_CDNS_52468879185839_0
timestamp 1707688321
transform 1 0 2128 0 1 0
box -26 -26 82 1426
use DFL1sd2_CDNS_52468879185839  DFL1sd2_CDNS_52468879185839_1
timestamp 1707688321
transform 1 0 1972 0 1 0
box -26 -26 82 1426
use DFL1sd2_CDNS_52468879185839  DFL1sd2_CDNS_52468879185839_2
timestamp 1707688321
transform 1 0 1816 0 1 0
box -26 -26 82 1426
use DFL1sd2_CDNS_52468879185839  DFL1sd2_CDNS_52468879185839_3
timestamp 1707688321
transform 1 0 1660 0 1 0
box -26 -26 82 1426
use DFL1sd2_CDNS_52468879185839  DFL1sd2_CDNS_52468879185839_4
timestamp 1707688321
transform 1 0 1504 0 1 0
box -26 -26 82 1426
use DFL1sd2_CDNS_52468879185839  DFL1sd2_CDNS_52468879185839_5
timestamp 1707688321
transform 1 0 1348 0 1 0
box -26 -26 82 1426
use DFL1sd2_CDNS_52468879185839  DFL1sd2_CDNS_52468879185839_6
timestamp 1707688321
transform 1 0 1192 0 1 0
box -26 -26 82 1426
use DFL1sd2_CDNS_52468879185839  DFL1sd2_CDNS_52468879185839_7
timestamp 1707688321
transform 1 0 1036 0 1 0
box -26 -26 82 1426
use DFL1sd2_CDNS_52468879185839  DFL1sd2_CDNS_52468879185839_8
timestamp 1707688321
transform 1 0 880 0 1 0
box -26 -26 82 1426
use DFL1sd2_CDNS_52468879185839  DFL1sd2_CDNS_52468879185839_9
timestamp 1707688321
transform 1 0 724 0 1 0
box -26 -26 82 1426
use DFL1sd2_CDNS_52468879185839  DFL1sd2_CDNS_52468879185839_10
timestamp 1707688321
transform 1 0 568 0 1 0
box -26 -26 82 1426
use DFL1sd2_CDNS_52468879185839  DFL1sd2_CDNS_52468879185839_11
timestamp 1707688321
transform 1 0 412 0 1 0
box -26 -26 82 1426
use DFL1sd2_CDNS_52468879185839  DFL1sd2_CDNS_52468879185839_12
timestamp 1707688321
transform 1 0 256 0 1 0
box -26 -26 82 1426
use DFL1sd2_CDNS_52468879185839  DFL1sd2_CDNS_52468879185839_13
timestamp 1707688321
transform 1 0 100 0 1 0
box -26 -26 82 1426
use DFL1sd_CDNS_52468879185838  DFL1sd_CDNS_52468879185838_0
timestamp 1707688321
transform -1 0 0 0 1 0
box -26 -26 79 1426
use DFL1sd_CDNS_52468879185838  DFL1sd_CDNS_52468879185838_1
timestamp 1707688321
transform 1 0 2284 0 1 0
box -26 -26 79 1426
<< labels >>
flabel comment s -28 675 -28 675 0 FreeSans 300 0 0 0 S
flabel comment s 128 675 128 675 0 FreeSans 300 0 0 0 D
flabel comment s 284 675 284 675 0 FreeSans 300 0 0 0 S
flabel comment s 440 675 440 675 0 FreeSans 300 0 0 0 D
flabel comment s 596 675 596 675 0 FreeSans 300 0 0 0 S
flabel comment s 752 675 752 675 0 FreeSans 300 0 0 0 D
flabel comment s 908 675 908 675 0 FreeSans 300 0 0 0 S
flabel comment s 1064 675 1064 675 0 FreeSans 300 0 0 0 D
flabel comment s 1220 675 1220 675 0 FreeSans 300 0 0 0 S
flabel comment s 1376 675 1376 675 0 FreeSans 300 0 0 0 D
flabel comment s 1532 675 1532 675 0 FreeSans 300 0 0 0 S
flabel comment s 1688 675 1688 675 0 FreeSans 300 0 0 0 D
flabel comment s 1844 675 1844 675 0 FreeSans 300 0 0 0 S
flabel comment s 2000 675 2000 675 0 FreeSans 300 0 0 0 D
flabel comment s 2156 675 2156 675 0 FreeSans 300 0 0 0 S
flabel comment s 2312 675 2312 675 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 34386552
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 34378694
<< end >>
