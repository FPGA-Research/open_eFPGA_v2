magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 1 21 585 203
rect 30 -17 64 21
<< locali >>
rect 19 315 85 485
rect 19 162 57 315
rect 205 265 248 331
rect 187 199 248 265
rect 283 199 340 331
rect 379 199 432 331
rect 475 199 524 331
rect 19 60 85 162
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 119 299 169 527
rect 207 399 257 483
rect 303 433 369 527
rect 415 399 465 483
rect 207 365 465 399
rect 501 399 567 485
rect 501 365 592 399
rect 91 199 153 265
rect 119 165 153 199
rect 558 165 592 365
rect 119 131 592 165
rect 119 17 185 97
rect 395 63 461 131
rect 495 17 561 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 379 199 432 331 6 A1
port 1 nsew signal input
rlabel locali s 283 199 340 331 6 A2
port 2 nsew signal input
rlabel locali s 187 199 248 265 6 A3
port 3 nsew signal input
rlabel locali s 205 265 248 331 6 A3
port 3 nsew signal input
rlabel locali s 475 199 524 331 6 B1
port 4 nsew signal input
rlabel metal1 s 0 -48 644 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 585 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 682 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 19 60 85 162 6 X
port 9 nsew signal output
rlabel locali s 19 162 57 315 6 X
port 9 nsew signal output
rlabel locali s 19 315 85 485 6 X
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 644 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 4105602
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 4099116
<< end >>
