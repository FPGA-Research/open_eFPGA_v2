magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -89 -36 189 236
<< pmos >>
rect 0 0 100 200
<< pdiff >>
rect -53 182 0 200
rect -53 148 -45 182
rect -11 148 0 182
rect -53 114 0 148
rect -53 80 -45 114
rect -11 80 0 114
rect -53 46 0 80
rect -53 12 -45 46
rect -11 12 0 46
rect -53 0 0 12
rect 100 0 150 200
<< pdiffc >>
rect -45 148 -11 182
rect -45 80 -11 114
rect -45 12 -11 46
<< poly >>
rect 0 200 100 226
rect 0 -26 100 0
<< locali >>
rect -45 182 -11 198
rect -45 114 -11 148
rect -45 46 -11 80
rect -45 -4 -11 12
<< metal1 >>
rect 105 -16 151 186
use hvDFL1sd_CDNS_5246887918589  hvDFL1sd_CDNS_5246887918589_0
timestamp 1707688321
transform -1 0 0 0 1 0
box 0 0 1 1
use hvDFM1sd_CDNS_52468879185130  hvDFM1sd_CDNS_52468879185130_0
timestamp 1707688321
transform 1 0 100 0 1 0
box -36 -36 89 236
<< labels >>
flabel comment s -28 97 -28 97 0 FreeSans 300 0 0 0 S
flabel comment s 128 85 128 85 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 86826700
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86825810
<< end >>
