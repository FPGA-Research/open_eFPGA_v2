magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< dnwell >>
rect 2776 28094 7826 39920
rect 2776 14263 6830 18335
<< nwell >>
rect 2696 39714 7906 40000
rect 2696 28300 2982 39714
rect 7620 28300 7906 39714
rect 2696 28014 7906 28300
rect 3941 24651 6047 26183
rect 4393 18415 5959 24251
rect 7259 21418 7759 21586
rect 2696 18129 6910 18415
rect 2696 14469 2982 18129
rect 6624 14469 6910 18129
rect 2696 14183 6910 14469
<< pwell >>
rect 3056 39554 5390 39640
rect 3056 30067 3142 39554
rect 5304 30302 5390 39554
rect 5614 30137 7508 30223
rect 5614 30067 5700 30137
rect 3056 29291 3574 30067
rect 5287 29291 5700 30067
rect 3056 29083 3142 29291
rect 5614 29083 5700 29291
rect 3056 28731 3574 29083
rect 5287 28731 5700 29083
rect 3056 28460 3142 28731
rect 5614 28460 5700 28731
rect 3056 28374 5700 28460
rect 2564 25625 3758 25711
rect 3672 18511 3758 25625
rect 3056 17969 6536 18055
rect 3056 17642 3422 17969
rect 3056 15988 3142 17642
rect 3839 16889 4242 17969
rect 5488 16889 5787 17969
rect 6450 17022 6536 17969
rect 3839 16769 4208 16889
rect 6185 16769 6536 17022
rect 3056 15689 3422 15988
rect 3056 14629 3142 15689
rect 3669 14629 4208 16769
rect 5862 14629 6536 16769
rect 3056 14543 6536 14629
<< mvndiff >>
rect 3304 29741 3548 30041
rect 5313 29741 5560 30041
rect 3304 29317 3548 29617
rect 5313 29317 5560 29617
rect 3304 28757 3548 29057
rect 5313 28757 5560 29057
rect 3196 17694 3396 17915
rect 3865 16915 4190 17915
rect 5540 16915 5761 17915
rect 3935 16143 4156 16743
rect 5914 16143 6135 16743
rect 3196 15715 3396 15936
rect 3935 15413 4156 16013
rect 5914 15413 6135 16013
rect 3935 14683 4156 15283
rect 5914 14683 6135 15283
<< mvpdiff >>
rect 4098 24717 4316 26117
rect 5672 24717 5890 26117
rect 4640 23796 4840 24017
rect 5064 23830 5148 24017
rect 5064 23796 5102 23830
rect 5136 23796 5148 23830
rect 5320 23830 5404 24017
rect 5320 23796 5358 23830
rect 5392 23796 5404 23830
rect 4640 20161 4840 20382
rect 5064 19604 5102 19638
rect 5136 19604 5148 19638
rect 5064 19417 5148 19604
rect 5320 19604 5358 19638
rect 5392 19604 5404 19638
rect 5320 19417 5404 19604
rect 4742 18786 4963 18986
rect 5321 18786 5542 18986
<< mvpdiffc >>
rect 5102 23796 5136 23830
rect 5358 23796 5392 23830
rect 5102 19604 5136 19638
rect 5358 19604 5392 19638
<< mvpsubdiff >>
rect 3082 39580 3154 39614
rect 3188 39580 3222 39614
rect 3256 39580 3290 39614
rect 3324 39580 3358 39614
rect 3392 39580 3426 39614
rect 3460 39580 3494 39614
rect 3528 39580 3562 39614
rect 3596 39580 3630 39614
rect 3664 39580 3698 39614
rect 3732 39580 3766 39614
rect 3800 39580 3834 39614
rect 3868 39580 3902 39614
rect 3936 39580 3970 39614
rect 4004 39580 4038 39614
rect 4072 39580 4106 39614
rect 4140 39580 4174 39614
rect 4208 39580 4242 39614
rect 4276 39580 4310 39614
rect 4344 39580 4378 39614
rect 4412 39580 4446 39614
rect 4480 39580 4514 39614
rect 4548 39580 4582 39614
rect 4616 39580 4650 39614
rect 4684 39580 4718 39614
rect 4752 39580 4786 39614
rect 4820 39580 4854 39614
rect 4888 39580 4922 39614
rect 4956 39580 4990 39614
rect 5024 39580 5058 39614
rect 5092 39580 5126 39614
rect 5160 39580 5194 39614
rect 5228 39580 5262 39614
rect 5296 39580 5364 39614
rect 3082 39546 3116 39580
rect 3082 39478 3116 39512
rect 5330 39508 5364 39580
rect 3082 39410 3116 39444
rect 3082 39342 3116 39376
rect 3082 39274 3116 39308
rect 3082 39206 3116 39240
rect 3082 39138 3116 39172
rect 3082 39070 3116 39104
rect 3082 39002 3116 39036
rect 3082 38934 3116 38968
rect 3082 38866 3116 38900
rect 3082 38798 3116 38832
rect 3082 38730 3116 38764
rect 3082 38662 3116 38696
rect 3082 38594 3116 38628
rect 3082 38526 3116 38560
rect 3082 38458 3116 38492
rect 3082 38390 3116 38424
rect 3082 38322 3116 38356
rect 3082 38254 3116 38288
rect 3082 38186 3116 38220
rect 3082 38118 3116 38152
rect 3082 38050 3116 38084
rect 3082 37982 3116 38016
rect 3082 37914 3116 37948
rect 3082 37846 3116 37880
rect 3082 37778 3116 37812
rect 3082 37710 3116 37744
rect 3082 37642 3116 37676
rect 3082 37574 3116 37608
rect 3082 37506 3116 37540
rect 3082 37438 3116 37472
rect 3082 37370 3116 37404
rect 3082 37302 3116 37336
rect 3082 37234 3116 37268
rect 3082 37166 3116 37200
rect 3082 37098 3116 37132
rect 3082 37030 3116 37064
rect 3082 36962 3116 36996
rect 3082 36894 3116 36928
rect 3082 36826 3116 36860
rect 3082 36758 3116 36792
rect 3082 36690 3116 36724
rect 3082 36622 3116 36656
rect 3082 36554 3116 36588
rect 3082 36486 3116 36520
rect 3082 36418 3116 36452
rect 3082 36350 3116 36384
rect 3082 36282 3116 36316
rect 3082 36214 3116 36248
rect 3082 36146 3116 36180
rect 3082 36078 3116 36112
rect 3082 36010 3116 36044
rect 3082 35942 3116 35976
rect 3082 35874 3116 35908
rect 3082 35806 3116 35840
rect 3082 35738 3116 35772
rect 3082 35670 3116 35704
rect 3082 35602 3116 35636
rect 3082 35534 3116 35568
rect 3082 35466 3116 35500
rect 3082 35398 3116 35432
rect 3082 35330 3116 35364
rect 3082 35262 3116 35296
rect 3082 35194 3116 35228
rect 3082 35126 3116 35160
rect 3082 35058 3116 35092
rect 3082 34990 3116 35024
rect 3082 34922 3116 34956
rect 3082 34854 3116 34888
rect 3082 34786 3116 34820
rect 3082 34718 3116 34752
rect 3082 34650 3116 34684
rect 3082 34582 3116 34616
rect 3082 34514 3116 34548
rect 3082 34446 3116 34480
rect 3082 34378 3116 34412
rect 3082 34310 3116 34344
rect 3082 34242 3116 34276
rect 3082 34174 3116 34208
rect 3082 34106 3116 34140
rect 3082 34038 3116 34072
rect 3082 33970 3116 34004
rect 3082 33902 3116 33936
rect 3082 33834 3116 33868
rect 3082 33766 3116 33800
rect 3082 33698 3116 33732
rect 3082 33630 3116 33664
rect 3082 33562 3116 33596
rect 3082 33494 3116 33528
rect 3082 33426 3116 33460
rect 3082 33358 3116 33392
rect 3082 33290 3116 33324
rect 3082 33222 3116 33256
rect 3082 33154 3116 33188
rect 3082 33086 3116 33120
rect 3082 33018 3116 33052
rect 3082 32950 3116 32984
rect 3082 32882 3116 32916
rect 3082 32814 3116 32848
rect 3082 32746 3116 32780
rect 3082 32678 3116 32712
rect 3082 32610 3116 32644
rect 3082 32542 3116 32576
rect 3082 32474 3116 32508
rect 3082 32406 3116 32440
rect 3082 32338 3116 32372
rect 3082 32270 3116 32304
rect 3082 32202 3116 32236
rect 3082 32134 3116 32168
rect 3082 32066 3116 32100
rect 3082 31998 3116 32032
rect 3082 31930 3116 31964
rect 3082 31862 3116 31896
rect 3082 31794 3116 31828
rect 3082 31726 3116 31760
rect 3082 31658 3116 31692
rect 3082 31590 3116 31624
rect 3082 31522 3116 31556
rect 3082 31454 3116 31488
rect 3082 31386 3116 31420
rect 3082 31318 3116 31352
rect 3082 31250 3116 31284
rect 3082 31182 3116 31216
rect 3082 31114 3116 31148
rect 3082 31046 3116 31080
rect 3082 30978 3116 31012
rect 3082 30910 3116 30944
rect 3082 30842 3116 30876
rect 3082 30774 3116 30808
rect 3082 30706 3116 30740
rect 3082 30638 3116 30672
rect 3082 30570 3116 30604
rect 3082 30502 3116 30536
rect 3082 30434 3116 30468
rect 3082 30366 3116 30400
rect 5330 39440 5364 39474
rect 5330 39372 5364 39406
rect 5330 39304 5364 39338
rect 5330 39236 5364 39270
rect 5330 39168 5364 39202
rect 5330 39100 5364 39134
rect 5330 39032 5364 39066
rect 5330 38964 5364 38998
rect 5330 38896 5364 38930
rect 5330 38828 5364 38862
rect 5330 38760 5364 38794
rect 5330 38692 5364 38726
rect 5330 38624 5364 38658
rect 5330 38556 5364 38590
rect 5330 38488 5364 38522
rect 5330 38420 5364 38454
rect 5330 38352 5364 38386
rect 5330 38284 5364 38318
rect 5330 38216 5364 38250
rect 5330 38148 5364 38182
rect 5330 38080 5364 38114
rect 5330 38012 5364 38046
rect 5330 37944 5364 37978
rect 5330 37876 5364 37910
rect 5330 37808 5364 37842
rect 5330 37740 5364 37774
rect 5330 37672 5364 37706
rect 5330 37604 5364 37638
rect 5330 37536 5364 37570
rect 5330 37468 5364 37502
rect 5330 37400 5364 37434
rect 5330 37332 5364 37366
rect 5330 37264 5364 37298
rect 5330 37196 5364 37230
rect 5330 37128 5364 37162
rect 5330 37060 5364 37094
rect 5330 36992 5364 37026
rect 5330 36924 5364 36958
rect 5330 36856 5364 36890
rect 5330 36788 5364 36822
rect 5330 36720 5364 36754
rect 5330 36652 5364 36686
rect 5330 36584 5364 36618
rect 5330 36516 5364 36550
rect 5330 36448 5364 36482
rect 5330 36380 5364 36414
rect 5330 36312 5364 36346
rect 5330 36244 5364 36278
rect 5330 36176 5364 36210
rect 5330 36108 5364 36142
rect 5330 36040 5364 36074
rect 5330 35972 5364 36006
rect 5330 35904 5364 35938
rect 5330 35836 5364 35870
rect 5330 35768 5364 35802
rect 5330 35700 5364 35734
rect 5330 35632 5364 35666
rect 5330 35564 5364 35598
rect 5330 35496 5364 35530
rect 5330 35428 5364 35462
rect 5330 35360 5364 35394
rect 5330 35292 5364 35326
rect 5330 35224 5364 35258
rect 5330 35156 5364 35190
rect 5330 35088 5364 35122
rect 5330 35020 5364 35054
rect 5330 34952 5364 34986
rect 5330 34884 5364 34918
rect 5330 34816 5364 34850
rect 5330 34748 5364 34782
rect 5330 34680 5364 34714
rect 5330 34612 5364 34646
rect 5330 34544 5364 34578
rect 5330 34476 5364 34510
rect 5330 34408 5364 34442
rect 5330 34340 5364 34374
rect 5330 34272 5364 34306
rect 5330 34204 5364 34238
rect 5330 34136 5364 34170
rect 5330 34068 5364 34102
rect 5330 34000 5364 34034
rect 5330 33932 5364 33966
rect 5330 33864 5364 33898
rect 5330 33796 5364 33830
rect 5330 33728 5364 33762
rect 5330 33660 5364 33694
rect 5330 33592 5364 33626
rect 5330 33524 5364 33558
rect 5330 33456 5364 33490
rect 5330 33388 5364 33422
rect 5330 33320 5364 33354
rect 5330 33252 5364 33286
rect 5330 33184 5364 33218
rect 5330 33116 5364 33150
rect 5330 33048 5364 33082
rect 5330 32980 5364 33014
rect 5330 32912 5364 32946
rect 5330 32844 5364 32878
rect 5330 32776 5364 32810
rect 5330 32708 5364 32742
rect 5330 32640 5364 32674
rect 5330 32572 5364 32606
rect 5330 32504 5364 32538
rect 5330 32436 5364 32470
rect 5330 32368 5364 32402
rect 5330 32300 5364 32334
rect 5330 32232 5364 32266
rect 5330 32164 5364 32198
rect 5330 32096 5364 32130
rect 5330 32028 5364 32062
rect 5330 31960 5364 31994
rect 5330 31892 5364 31926
rect 5330 31824 5364 31858
rect 5330 31756 5364 31790
rect 5330 31688 5364 31722
rect 5330 31620 5364 31654
rect 5330 31552 5364 31586
rect 5330 31484 5364 31518
rect 5330 31416 5364 31450
rect 5330 31348 5364 31382
rect 5330 31280 5364 31314
rect 5330 31212 5364 31246
rect 5330 31144 5364 31178
rect 5330 31076 5364 31110
rect 5330 31008 5364 31042
rect 5330 30940 5364 30974
rect 5330 30872 5364 30906
rect 5330 30804 5364 30838
rect 5330 30736 5364 30770
rect 5330 30668 5364 30702
rect 5330 30600 5364 30634
rect 5330 30532 5364 30566
rect 5330 30464 5364 30498
rect 5330 30396 5364 30430
rect 3082 30298 3116 30332
rect 5330 30328 5364 30362
rect 3082 30230 3116 30264
rect 3082 30162 3116 30196
rect 5640 30163 5664 30197
rect 5698 30163 5735 30197
rect 5769 30163 5806 30197
rect 5840 30163 5877 30197
rect 5911 30163 5948 30197
rect 5982 30163 6019 30197
rect 6053 30163 6090 30197
rect 6124 30163 6161 30197
rect 6195 30163 6232 30197
rect 6266 30163 6303 30197
rect 6337 30163 6374 30197
rect 6408 30163 6444 30197
rect 6478 30163 6514 30197
rect 6548 30163 6584 30197
rect 6618 30163 6654 30197
rect 6688 30163 6724 30197
rect 6758 30163 6794 30197
rect 6828 30163 6864 30197
rect 6898 30163 6934 30197
rect 6968 30163 7004 30197
rect 7038 30163 7074 30197
rect 7108 30163 7144 30197
rect 7178 30163 7214 30197
rect 7248 30163 7284 30197
rect 7318 30163 7354 30197
rect 7388 30163 7424 30197
rect 7458 30163 7482 30197
rect 3082 30094 3116 30128
rect 3082 30026 3116 30060
rect 3082 29958 3116 29992
rect 3082 29890 3116 29924
rect 3082 29822 3116 29856
rect 3082 29754 3116 29788
rect 5640 29998 5674 30068
rect 5640 29930 5674 29964
rect 5640 29862 5674 29896
rect 5640 29794 5674 29828
rect 3082 29686 3116 29720
rect 3082 29618 3116 29652
rect 5640 29726 5674 29760
rect 5640 29658 5674 29692
rect 3082 29550 3116 29584
rect 3082 29482 3116 29516
rect 3082 29414 3116 29448
rect 3082 29346 3116 29380
rect 5640 29590 5674 29624
rect 5640 29522 5674 29556
rect 5640 29454 5674 29488
rect 5640 29386 5674 29420
rect 5640 29318 5674 29352
rect 3082 29278 3116 29312
rect 3082 29210 3116 29244
rect 5640 29250 5674 29284
rect 3082 29142 3116 29176
rect 5640 29182 5674 29216
rect 3082 29074 3116 29108
rect 5640 29114 5674 29148
rect 3082 29006 3116 29040
rect 3082 28938 3116 28972
rect 3082 28870 3116 28904
rect 3082 28802 3116 28836
rect 3082 28734 3116 28768
rect 5640 29046 5674 29080
rect 5640 28978 5674 29012
rect 5640 28910 5674 28944
rect 5640 28842 5674 28876
rect 5640 28774 5674 28808
rect 3082 28666 3116 28700
rect 3082 28598 3116 28632
rect 3082 28530 3116 28564
rect 3082 28434 3116 28496
rect 5640 28706 5674 28740
rect 5640 28638 5674 28672
rect 5640 28570 5674 28604
rect 5640 28502 5674 28536
rect 5640 28434 5674 28468
rect 3082 28400 3150 28434
rect 3184 28400 3218 28434
rect 3252 28400 3286 28434
rect 3320 28400 3354 28434
rect 3388 28400 3422 28434
rect 3456 28400 3490 28434
rect 3524 28400 3558 28434
rect 3592 28400 3626 28434
rect 3660 28400 3694 28434
rect 3728 28400 3762 28434
rect 3796 28400 3830 28434
rect 3864 28400 3898 28434
rect 3932 28400 3966 28434
rect 4000 28400 4034 28434
rect 4068 28400 4102 28434
rect 4136 28400 4170 28434
rect 4204 28400 4238 28434
rect 4272 28400 4306 28434
rect 4340 28400 4374 28434
rect 4408 28400 4442 28434
rect 4476 28400 4510 28434
rect 4544 28400 4578 28434
rect 4612 28400 4646 28434
rect 4680 28400 4714 28434
rect 4748 28400 4782 28434
rect 4816 28400 4850 28434
rect 4884 28400 4918 28434
rect 4952 28400 4986 28434
rect 5020 28400 5054 28434
rect 5088 28400 5122 28434
rect 5156 28400 5190 28434
rect 5224 28400 5258 28434
rect 5292 28400 5326 28434
rect 5360 28400 5394 28434
rect 5428 28400 5462 28434
rect 5496 28400 5530 28434
rect 5564 28400 5674 28434
rect 2590 25651 2678 25685
rect 2712 25651 2746 25685
rect 2780 25651 2814 25685
rect 2848 25651 2882 25685
rect 2916 25651 2950 25685
rect 2984 25651 3018 25685
rect 3052 25651 3086 25685
rect 3120 25651 3154 25685
rect 3188 25651 3222 25685
rect 3256 25651 3290 25685
rect 3324 25651 3358 25685
rect 3392 25651 3426 25685
rect 3460 25651 3494 25685
rect 3528 25651 3562 25685
rect 3596 25651 3630 25685
rect 3664 25651 3732 25685
rect 3698 25609 3732 25651
rect 3698 25541 3732 25575
rect 3698 25473 3732 25507
rect 3698 25405 3732 25439
rect 3698 25337 3732 25371
rect 3698 25269 3732 25303
rect 3698 25201 3732 25235
rect 3698 25133 3732 25167
rect 3698 25065 3732 25099
rect 3698 24997 3732 25031
rect 3698 24929 3732 24963
rect 3698 24861 3732 24895
rect 3698 24793 3732 24827
rect 3698 24725 3732 24759
rect 3698 24657 3732 24691
rect 3698 24589 3732 24623
rect 3698 24521 3732 24555
rect 3698 24453 3732 24487
rect 3698 24385 3732 24419
rect 3698 24317 3732 24351
rect 3698 24249 3732 24283
rect 3698 24181 3732 24215
rect 3698 24113 3732 24147
rect 3698 24045 3732 24079
rect 3698 23977 3732 24011
rect 3698 23909 3732 23943
rect 3698 23841 3732 23875
rect 3698 23773 3732 23807
rect 3698 23705 3732 23739
rect 3698 23637 3732 23671
rect 3698 23569 3732 23603
rect 3698 23501 3732 23535
rect 3698 23433 3732 23467
rect 3698 23365 3732 23399
rect 3698 23297 3732 23331
rect 3698 23229 3732 23263
rect 3698 23161 3732 23195
rect 3698 23093 3732 23127
rect 3698 23025 3732 23059
rect 3698 22957 3732 22991
rect 3698 22889 3732 22923
rect 3698 22821 3732 22855
rect 3698 22753 3732 22787
rect 3698 22685 3732 22719
rect 3698 22617 3732 22651
rect 3698 22549 3732 22583
rect 3698 22481 3732 22515
rect 3698 22413 3732 22447
rect 3698 22345 3732 22379
rect 3698 22277 3732 22311
rect 3698 22209 3732 22243
rect 3698 22141 3732 22175
rect 3698 22073 3732 22107
rect 3698 22005 3732 22039
rect 3698 21937 3732 21971
rect 3698 21869 3732 21903
rect 3698 21801 3732 21835
rect 3698 21733 3732 21767
rect 3698 21665 3732 21699
rect 3698 21597 3732 21631
rect 3698 21529 3732 21563
rect 3698 21461 3732 21495
rect 3698 21393 3732 21427
rect 3698 21325 3732 21359
rect 3698 21257 3732 21291
rect 3698 21189 3732 21223
rect 3698 21121 3732 21155
rect 3698 21053 3732 21087
rect 3698 20985 3732 21019
rect 3698 20917 3732 20951
rect 3698 20849 3732 20883
rect 3698 20781 3732 20815
rect 3698 20713 3732 20747
rect 3698 20645 3732 20679
rect 3698 20577 3732 20611
rect 3698 20509 3732 20543
rect 3698 20441 3732 20475
rect 3698 20373 3732 20407
rect 3698 20305 3732 20339
rect 3698 20237 3732 20271
rect 3698 20169 3732 20203
rect 3698 20101 3732 20135
rect 3698 20033 3732 20067
rect 3698 19965 3732 19999
rect 3698 19897 3732 19931
rect 3698 19829 3732 19863
rect 3698 19761 3732 19795
rect 3698 19693 3732 19727
rect 3698 19625 3732 19659
rect 3698 19557 3732 19591
rect 3698 19489 3732 19523
rect 3698 19421 3732 19455
rect 3698 19353 3732 19387
rect 3698 19285 3732 19319
rect 3698 19217 3732 19251
rect 3698 19149 3732 19183
rect 3698 19081 3732 19115
rect 3698 19013 3732 19047
rect 3698 18945 3732 18979
rect 3698 18877 3732 18911
rect 3698 18809 3732 18843
rect 3698 18741 3732 18775
rect 3698 18673 3732 18707
rect 3698 18605 3732 18639
rect 3698 18537 3732 18571
rect 3082 17995 3150 18029
rect 3184 17995 3218 18029
rect 3252 17995 3286 18029
rect 3320 17995 3354 18029
rect 3388 17995 3422 18029
rect 3456 17995 3490 18029
rect 3524 17995 3558 18029
rect 3592 17995 3626 18029
rect 3660 17995 3694 18029
rect 3728 17995 3762 18029
rect 3796 17995 3830 18029
rect 3864 17995 3898 18029
rect 3932 17995 3966 18029
rect 4000 17995 4034 18029
rect 4068 17995 4102 18029
rect 4136 17995 4170 18029
rect 4204 17995 4238 18029
rect 4272 17995 4306 18029
rect 4340 17995 4374 18029
rect 4408 17995 4442 18029
rect 4476 17995 4510 18029
rect 4544 17995 4578 18029
rect 4612 17995 4646 18029
rect 4680 17995 4714 18029
rect 4748 17995 4782 18029
rect 4816 17995 4850 18029
rect 4884 17995 4918 18029
rect 4952 17995 4986 18029
rect 5020 17995 5054 18029
rect 5088 17995 5122 18029
rect 5156 17995 5190 18029
rect 5224 17995 5258 18029
rect 5292 17995 5326 18029
rect 5360 17995 5394 18029
rect 5428 17995 5462 18029
rect 5496 17995 5530 18029
rect 5564 17995 5598 18029
rect 5632 17995 5666 18029
rect 5700 17995 5734 18029
rect 5768 17995 5802 18029
rect 5836 17995 5870 18029
rect 5904 17995 5938 18029
rect 5972 17995 6006 18029
rect 6040 17995 6074 18029
rect 6108 17995 6142 18029
rect 6176 17995 6210 18029
rect 6244 17995 6278 18029
rect 6312 17995 6346 18029
rect 6380 17995 6510 18029
rect 3082 17935 3116 17995
rect 6476 17961 6510 17995
rect 3082 17867 3116 17901
rect 3082 17799 3116 17833
rect 3082 17731 3116 17765
rect 3082 17663 3116 17697
rect 3082 17595 3116 17629
rect 3082 17527 3116 17561
rect 3082 17459 3116 17493
rect 3082 17391 3116 17425
rect 3082 17323 3116 17357
rect 3082 17255 3116 17289
rect 3082 17187 3116 17221
rect 3082 17119 3116 17153
rect 3082 17051 3116 17085
rect 3082 16983 3116 17017
rect 3082 16915 3116 16949
rect 3082 16847 3116 16881
rect 3082 16779 3116 16813
rect 3082 16711 3116 16745
rect 3082 16643 3116 16677
rect 3082 16575 3116 16609
rect 3082 16507 3116 16541
rect 3082 16439 3116 16473
rect 3082 16371 3116 16405
rect 3082 16303 3116 16337
rect 3082 16235 3116 16269
rect 3082 16167 3116 16201
rect 3082 16099 3116 16133
rect 3082 16031 3116 16065
rect 6476 17893 6510 17927
rect 6476 17825 6510 17859
rect 6476 17757 6510 17791
rect 6476 17689 6510 17723
rect 6476 17621 6510 17655
rect 6476 17553 6510 17587
rect 6476 17485 6510 17519
rect 6476 17417 6510 17451
rect 6476 17349 6510 17383
rect 6476 17281 6510 17315
rect 6476 17213 6510 17247
rect 6476 17145 6510 17179
rect 6476 17077 6510 17111
rect 6476 17009 6510 17043
rect 6211 16962 6371 16996
rect 6245 16928 6337 16962
rect 6211 16819 6371 16928
rect 6245 16785 6337 16819
rect 3695 16709 3855 16743
rect 3729 16675 3821 16709
rect 3695 16564 3855 16675
rect 3729 16530 3821 16564
rect 3695 16419 3855 16530
rect 3729 16385 3821 16419
rect 3695 16274 3855 16385
rect 3729 16240 3821 16274
rect 3695 16129 3855 16240
rect 6211 16676 6371 16785
rect 6245 16642 6337 16676
rect 6211 16533 6371 16642
rect 6245 16499 6337 16533
rect 6211 16390 6371 16499
rect 6245 16356 6337 16390
rect 6211 16247 6371 16356
rect 6245 16213 6337 16247
rect 3729 16095 3821 16129
rect 3082 15963 3116 15997
rect 3695 15984 3855 16095
rect 6211 16104 6371 16213
rect 6245 16070 6337 16104
rect 3729 15950 3821 15984
rect 3082 15895 3116 15929
rect 3082 15827 3116 15861
rect 3082 15759 3116 15793
rect 3082 15691 3116 15725
rect 3695 15839 3855 15950
rect 3729 15805 3821 15839
rect 3082 15623 3116 15657
rect 3082 15555 3116 15589
rect 3082 15487 3116 15521
rect 3082 15419 3116 15453
rect 3082 15351 3116 15385
rect 3082 15283 3116 15317
rect 3082 15215 3116 15249
rect 3082 15147 3116 15181
rect 3082 15079 3116 15113
rect 3082 15011 3116 15045
rect 3082 14943 3116 14977
rect 3082 14875 3116 14909
rect 3082 14807 3116 14841
rect 3082 14739 3116 14773
rect 3082 14671 3116 14705
rect 3082 14603 3116 14637
rect 3695 15693 3855 15805
rect 3729 15659 3821 15693
rect 3695 15547 3855 15659
rect 3729 15513 3821 15547
rect 3695 15401 3855 15513
rect 6211 15961 6371 16070
rect 6245 15927 6337 15961
rect 6211 15818 6371 15927
rect 6245 15784 6337 15818
rect 6211 15675 6371 15784
rect 6245 15641 6337 15675
rect 6211 15532 6371 15641
rect 6245 15498 6337 15532
rect 3729 15367 3821 15401
rect 6211 15389 6371 15498
rect 3695 15255 3855 15367
rect 6245 15355 6337 15389
rect 3729 15221 3821 15255
rect 3695 15109 3855 15221
rect 3729 15075 3821 15109
rect 3695 14963 3855 15075
rect 3729 14929 3821 14963
rect 3695 14817 3855 14929
rect 3729 14783 3821 14817
rect 3695 14671 3855 14783
rect 6211 15246 6371 15355
rect 6245 15212 6337 15246
rect 6211 15103 6371 15212
rect 6245 15069 6337 15103
rect 6211 14959 6371 15069
rect 6245 14925 6337 14959
rect 6211 14815 6371 14925
rect 6245 14781 6337 14815
rect 3729 14637 3821 14671
rect 3695 14603 3855 14637
rect 6211 14671 6371 14781
rect 6245 14637 6337 14671
rect 6211 14603 6371 14637
rect 6476 16941 6510 16975
rect 6476 16873 6510 16907
rect 6476 16805 6510 16839
rect 6476 16737 6510 16771
rect 6476 16669 6510 16703
rect 6476 16601 6510 16635
rect 6476 16533 6510 16567
rect 6476 16465 6510 16499
rect 6476 16397 6510 16431
rect 6476 16329 6510 16363
rect 6476 16261 6510 16295
rect 6476 16193 6510 16227
rect 6476 16125 6510 16159
rect 6476 16057 6510 16091
rect 6476 15989 6510 16023
rect 6476 15921 6510 15955
rect 6476 15853 6510 15887
rect 6476 15785 6510 15819
rect 6476 15717 6510 15751
rect 6476 15649 6510 15683
rect 6476 15581 6510 15615
rect 6476 15513 6510 15547
rect 6476 15445 6510 15479
rect 6476 15377 6510 15411
rect 6476 15309 6510 15343
rect 6476 15241 6510 15275
rect 6476 15173 6510 15207
rect 6476 15105 6510 15139
rect 6476 15037 6510 15071
rect 6476 14969 6510 15003
rect 6476 14901 6510 14935
rect 6476 14833 6510 14867
rect 6476 14765 6510 14799
rect 6476 14697 6510 14731
rect 6476 14603 6510 14663
rect 3082 14569 3212 14603
rect 3246 14569 3280 14603
rect 3314 14569 3348 14603
rect 3382 14569 3416 14603
rect 3450 14569 3484 14603
rect 3518 14569 3552 14603
rect 3586 14569 3620 14603
rect 3654 14569 3688 14603
rect 3722 14569 3756 14603
rect 3790 14569 3824 14603
rect 3858 14569 3892 14603
rect 3926 14569 3960 14603
rect 3994 14569 4028 14603
rect 4062 14569 4096 14603
rect 4130 14569 4164 14603
rect 4198 14569 4232 14603
rect 4266 14569 4300 14603
rect 4334 14569 4368 14603
rect 4402 14569 4436 14603
rect 4470 14569 4504 14603
rect 4538 14569 4572 14603
rect 4606 14569 4640 14603
rect 4674 14569 4708 14603
rect 4742 14569 4776 14603
rect 4810 14569 4844 14603
rect 4878 14569 4912 14603
rect 4946 14569 4980 14603
rect 5014 14569 5048 14603
rect 5082 14569 5116 14603
rect 5150 14569 5184 14603
rect 5218 14569 5252 14603
rect 5286 14569 5320 14603
rect 5354 14569 5388 14603
rect 5422 14569 5456 14603
rect 5490 14569 5524 14603
rect 5558 14569 5592 14603
rect 5626 14569 5660 14603
rect 5694 14569 5728 14603
rect 5762 14569 5796 14603
rect 5830 14569 5864 14603
rect 5898 14569 5932 14603
rect 5966 14569 6000 14603
rect 6034 14569 6068 14603
rect 6102 14569 6136 14603
rect 6170 14569 6204 14603
rect 6238 14569 6272 14603
rect 6306 14569 6340 14603
rect 6374 14569 6408 14603
rect 6442 14569 6510 14603
<< mvnsubdiff >>
rect 2822 39840 2918 39874
rect 2952 39840 2986 39874
rect 3020 39840 3054 39874
rect 3088 39840 3122 39874
rect 3156 39840 3190 39874
rect 3224 39840 3258 39874
rect 3292 39840 3326 39874
rect 3360 39840 3394 39874
rect 3428 39840 3462 39874
rect 3496 39840 3530 39874
rect 3564 39840 3598 39874
rect 3632 39840 3666 39874
rect 3700 39840 3734 39874
rect 3768 39840 3802 39874
rect 3836 39840 3870 39874
rect 3904 39840 3938 39874
rect 3972 39840 4006 39874
rect 4040 39840 4074 39874
rect 4108 39840 4142 39874
rect 4176 39840 4210 39874
rect 4244 39840 4278 39874
rect 4312 39840 4346 39874
rect 4380 39840 4414 39874
rect 4448 39840 4482 39874
rect 4516 39840 4550 39874
rect 4584 39840 4618 39874
rect 4652 39840 4686 39874
rect 4720 39840 4754 39874
rect 4788 39840 4822 39874
rect 4856 39840 4890 39874
rect 4924 39840 4958 39874
rect 4992 39840 5026 39874
rect 5060 39840 5094 39874
rect 5128 39840 5162 39874
rect 5196 39840 5230 39874
rect 5264 39840 5298 39874
rect 5332 39840 5366 39874
rect 5400 39840 5434 39874
rect 5468 39840 5502 39874
rect 5536 39840 5570 39874
rect 5604 39840 5638 39874
rect 5672 39840 5706 39874
rect 5740 39840 5774 39874
rect 5808 39840 5842 39874
rect 5876 39840 5910 39874
rect 5944 39840 5978 39874
rect 6012 39840 6046 39874
rect 6080 39840 6114 39874
rect 6148 39840 6182 39874
rect 6216 39840 6250 39874
rect 6284 39840 6318 39874
rect 6352 39840 6386 39874
rect 6420 39840 6454 39874
rect 6488 39840 6522 39874
rect 6556 39840 6590 39874
rect 6624 39840 6658 39874
rect 6692 39840 6726 39874
rect 6760 39840 6794 39874
rect 6828 39840 6862 39874
rect 6896 39840 6930 39874
rect 6964 39840 6998 39874
rect 7032 39840 7066 39874
rect 7100 39840 7134 39874
rect 7168 39840 7202 39874
rect 7236 39840 7270 39874
rect 7304 39840 7338 39874
rect 7372 39840 7406 39874
rect 7440 39840 7474 39874
rect 7508 39840 7542 39874
rect 7576 39840 7610 39874
rect 7644 39840 7678 39874
rect 7712 39840 7780 39874
rect 2822 39806 2856 39840
rect 2822 39738 2856 39772
rect 2822 39670 2856 39704
rect 2822 39602 2856 39636
rect 7746 39802 7780 39840
rect 7746 39734 7780 39768
rect 7746 39666 7780 39700
rect 2822 39534 2856 39568
rect 2822 39466 2856 39500
rect 2822 39398 2856 39432
rect 2822 39330 2856 39364
rect 2822 39262 2856 39296
rect 2822 39194 2856 39228
rect 2822 39126 2856 39160
rect 2822 39058 2856 39092
rect 2822 38990 2856 39024
rect 2822 38922 2856 38956
rect 2822 38854 2856 38888
rect 2822 38786 2856 38820
rect 2822 38718 2856 38752
rect 2822 38650 2856 38684
rect 2822 38582 2856 38616
rect 2822 38514 2856 38548
rect 2822 38446 2856 38480
rect 2822 38378 2856 38412
rect 2822 38310 2856 38344
rect 2822 38242 2856 38276
rect 2822 38174 2856 38208
rect 2822 38106 2856 38140
rect 2822 38038 2856 38072
rect 2822 37970 2856 38004
rect 2822 37902 2856 37936
rect 2822 37834 2856 37868
rect 2822 37766 2856 37800
rect 2822 37698 2856 37732
rect 2822 37630 2856 37664
rect 2822 37562 2856 37596
rect 2822 37494 2856 37528
rect 2822 37426 2856 37460
rect 2822 37358 2856 37392
rect 2822 37290 2856 37324
rect 2822 37222 2856 37256
rect 2822 37154 2856 37188
rect 2822 37086 2856 37120
rect 2822 37018 2856 37052
rect 2822 36950 2856 36984
rect 2822 36882 2856 36916
rect 2822 36814 2856 36848
rect 2822 36746 2856 36780
rect 2822 36678 2856 36712
rect 2822 36610 2856 36644
rect 2822 36542 2856 36576
rect 2822 36474 2856 36508
rect 2822 36406 2856 36440
rect 2822 36338 2856 36372
rect 2822 36270 2856 36304
rect 2822 36202 2856 36236
rect 2822 36134 2856 36168
rect 2822 36066 2856 36100
rect 2822 35998 2856 36032
rect 2822 35930 2856 35964
rect 2822 35862 2856 35896
rect 2822 35794 2856 35828
rect 2822 35726 2856 35760
rect 2822 35658 2856 35692
rect 2822 35590 2856 35624
rect 2822 35522 2856 35556
rect 2822 35454 2856 35488
rect 2822 35386 2856 35420
rect 2822 35318 2856 35352
rect 2822 35250 2856 35284
rect 2822 35182 2856 35216
rect 2822 35114 2856 35148
rect 2822 35046 2856 35080
rect 2822 34978 2856 35012
rect 2822 34910 2856 34944
rect 2822 34842 2856 34876
rect 2822 34774 2856 34808
rect 2822 34706 2856 34740
rect 2822 34638 2856 34672
rect 2822 34570 2856 34604
rect 2822 34502 2856 34536
rect 2822 34434 2856 34468
rect 2822 34366 2856 34400
rect 2822 34298 2856 34332
rect 2822 34230 2856 34264
rect 2822 34162 2856 34196
rect 2822 34094 2856 34128
rect 2822 34026 2856 34060
rect 2822 33958 2856 33992
rect 2822 33890 2856 33924
rect 2822 33822 2856 33856
rect 2822 33754 2856 33788
rect 2822 33686 2856 33720
rect 2822 33618 2856 33652
rect 2822 33550 2856 33584
rect 2822 33482 2856 33516
rect 2822 33414 2856 33448
rect 2822 33346 2856 33380
rect 2822 33278 2856 33312
rect 2822 33210 2856 33244
rect 2822 33142 2856 33176
rect 2822 33074 2856 33108
rect 2822 33006 2856 33040
rect 2822 32938 2856 32972
rect 2822 32870 2856 32904
rect 2822 32802 2856 32836
rect 2822 32734 2856 32768
rect 2822 32666 2856 32700
rect 2822 32598 2856 32632
rect 2822 32530 2856 32564
rect 2822 32462 2856 32496
rect 2822 32394 2856 32428
rect 2822 32326 2856 32360
rect 2822 32258 2856 32292
rect 2822 32190 2856 32224
rect 2822 32122 2856 32156
rect 2822 32054 2856 32088
rect 2822 31986 2856 32020
rect 2822 31918 2856 31952
rect 2822 31850 2856 31884
rect 2822 31782 2856 31816
rect 2822 31714 2856 31748
rect 2822 31646 2856 31680
rect 2822 31578 2856 31612
rect 2822 31510 2856 31544
rect 2822 31442 2856 31476
rect 2822 31374 2856 31408
rect 2822 31306 2856 31340
rect 2822 31238 2856 31272
rect 2822 31170 2856 31204
rect 2822 31102 2856 31136
rect 2822 31034 2856 31068
rect 2822 30966 2856 31000
rect 2822 30898 2856 30932
rect 2822 30830 2856 30864
rect 2822 30762 2856 30796
rect 2822 30694 2856 30728
rect 2822 30626 2856 30660
rect 2822 30558 2856 30592
rect 2822 30490 2856 30524
rect 2822 30422 2856 30456
rect 2822 30354 2856 30388
rect 2822 30286 2856 30320
rect 2822 30218 2856 30252
rect 2822 30150 2856 30184
rect 2822 30082 2856 30116
rect 2822 30014 2856 30048
rect 2822 29946 2856 29980
rect 2822 29878 2856 29912
rect 2822 29810 2856 29844
rect 2822 29742 2856 29776
rect 2822 29674 2856 29708
rect 2822 29606 2856 29640
rect 2822 29538 2856 29572
rect 2822 29470 2856 29504
rect 2822 29402 2856 29436
rect 2822 29334 2856 29368
rect 2822 29266 2856 29300
rect 2822 29198 2856 29232
rect 2822 29130 2856 29164
rect 2822 29062 2856 29096
rect 2822 28994 2856 29028
rect 2822 28926 2856 28960
rect 2822 28858 2856 28892
rect 2822 28790 2856 28824
rect 2822 28722 2856 28756
rect 2822 28654 2856 28688
rect 2822 28586 2856 28620
rect 2822 28518 2856 28552
rect 2822 28450 2856 28484
rect 2822 28382 2856 28416
rect 7746 39598 7780 39632
rect 7746 39530 7780 39564
rect 7746 39462 7780 39496
rect 7746 39394 7780 39428
rect 7746 39326 7780 39360
rect 7746 39258 7780 39292
rect 7746 39190 7780 39224
rect 7746 39122 7780 39156
rect 7746 39054 7780 39088
rect 7746 38986 7780 39020
rect 7746 38918 7780 38952
rect 7746 38850 7780 38884
rect 7746 38782 7780 38816
rect 7746 38714 7780 38748
rect 7746 38646 7780 38680
rect 7746 38578 7780 38612
rect 7746 38510 7780 38544
rect 7746 38442 7780 38476
rect 7746 38374 7780 38408
rect 7746 38306 7780 38340
rect 7746 38238 7780 38272
rect 7746 38170 7780 38204
rect 7746 38102 7780 38136
rect 7746 38034 7780 38068
rect 7746 37966 7780 38000
rect 7746 37898 7780 37932
rect 7746 37830 7780 37864
rect 7746 37762 7780 37796
rect 7746 37694 7780 37728
rect 7746 37626 7780 37660
rect 7746 37558 7780 37592
rect 7746 37490 7780 37524
rect 7746 37422 7780 37456
rect 7746 37354 7780 37388
rect 7746 37286 7780 37320
rect 7746 37218 7780 37252
rect 7746 37150 7780 37184
rect 7746 37082 7780 37116
rect 7746 37014 7780 37048
rect 7746 36946 7780 36980
rect 7746 36878 7780 36912
rect 7746 36810 7780 36844
rect 7746 36742 7780 36776
rect 7746 36674 7780 36708
rect 7746 36606 7780 36640
rect 7746 36538 7780 36572
rect 7746 36470 7780 36504
rect 7746 36402 7780 36436
rect 7746 36334 7780 36368
rect 7746 36266 7780 36300
rect 7746 36198 7780 36232
rect 7746 36130 7780 36164
rect 7746 36062 7780 36096
rect 7746 35994 7780 36028
rect 7746 35926 7780 35960
rect 7746 35858 7780 35892
rect 7746 35790 7780 35824
rect 7746 35722 7780 35756
rect 7746 35654 7780 35688
rect 7746 35586 7780 35620
rect 7746 35518 7780 35552
rect 7746 35450 7780 35484
rect 7746 35382 7780 35416
rect 7746 35314 7780 35348
rect 7746 35246 7780 35280
rect 7746 35178 7780 35212
rect 7746 35110 7780 35144
rect 7746 35042 7780 35076
rect 7746 34974 7780 35008
rect 7746 34906 7780 34940
rect 7746 34838 7780 34872
rect 7746 34770 7780 34804
rect 7746 34702 7780 34736
rect 7746 34634 7780 34668
rect 7746 34566 7780 34600
rect 7746 34498 7780 34532
rect 7746 34430 7780 34464
rect 7746 34362 7780 34396
rect 7746 34294 7780 34328
rect 7746 34226 7780 34260
rect 7746 34158 7780 34192
rect 7746 34090 7780 34124
rect 7746 34022 7780 34056
rect 7746 33954 7780 33988
rect 7746 33886 7780 33920
rect 7746 33818 7780 33852
rect 7746 33750 7780 33784
rect 7746 33682 7780 33716
rect 7746 33614 7780 33648
rect 7746 33546 7780 33580
rect 7746 33478 7780 33512
rect 7746 33410 7780 33444
rect 7746 33342 7780 33376
rect 7746 33274 7780 33308
rect 7746 33206 7780 33240
rect 7746 33138 7780 33172
rect 7746 33070 7780 33104
rect 7746 33002 7780 33036
rect 7746 32934 7780 32968
rect 7746 32866 7780 32900
rect 7746 32798 7780 32832
rect 7746 32730 7780 32764
rect 7746 32662 7780 32696
rect 7746 32594 7780 32628
rect 7746 32526 7780 32560
rect 7746 32458 7780 32492
rect 7746 32390 7780 32424
rect 7746 32322 7780 32356
rect 7746 32254 7780 32288
rect 7746 32186 7780 32220
rect 7746 32118 7780 32152
rect 7746 32050 7780 32084
rect 7746 31982 7780 32016
rect 7746 31914 7780 31948
rect 7746 31846 7780 31880
rect 7746 31778 7780 31812
rect 7746 31710 7780 31744
rect 7746 31642 7780 31676
rect 7746 31574 7780 31608
rect 7746 31506 7780 31540
rect 7746 31438 7780 31472
rect 7746 31370 7780 31404
rect 7746 31302 7780 31336
rect 7746 31234 7780 31268
rect 7746 31166 7780 31200
rect 7746 31098 7780 31132
rect 7746 31030 7780 31064
rect 7746 30962 7780 30996
rect 7746 30894 7780 30928
rect 7746 30826 7780 30860
rect 7746 30758 7780 30792
rect 7746 30690 7780 30724
rect 7746 30622 7780 30656
rect 7746 30554 7780 30588
rect 7746 30486 7780 30520
rect 7746 30418 7780 30452
rect 7746 30350 7780 30384
rect 7746 30282 7780 30316
rect 7746 30214 7780 30248
rect 7746 30146 7780 30180
rect 7746 30078 7780 30112
rect 7746 30010 7780 30044
rect 7746 29942 7780 29976
rect 7746 29874 7780 29908
rect 7746 29806 7780 29840
rect 7746 29738 7780 29772
rect 7746 29670 7780 29704
rect 7746 29602 7780 29636
rect 7746 29534 7780 29568
rect 7746 29466 7780 29500
rect 7746 29398 7780 29432
rect 7746 29330 7780 29364
rect 7746 29262 7780 29296
rect 7746 29194 7780 29228
rect 7746 29126 7780 29160
rect 7746 29058 7780 29092
rect 7746 28990 7780 29024
rect 7746 28922 7780 28956
rect 7746 28854 7780 28888
rect 7746 28786 7780 28820
rect 7746 28718 7780 28752
rect 7746 28650 7780 28684
rect 7746 28582 7780 28616
rect 7746 28514 7780 28548
rect 7746 28446 7780 28480
rect 2822 28266 2856 28348
rect 2822 28174 2856 28232
rect 7746 28378 7780 28412
rect 7746 28310 7780 28344
rect 7746 28242 7780 28276
rect 7746 28174 7780 28208
rect 2822 28140 2890 28174
rect 2924 28140 2958 28174
rect 2992 28140 3026 28174
rect 3060 28140 3094 28174
rect 3128 28140 3162 28174
rect 3196 28140 3230 28174
rect 3264 28140 3298 28174
rect 3332 28140 3366 28174
rect 3400 28140 3434 28174
rect 3468 28140 3502 28174
rect 3536 28140 3570 28174
rect 3604 28140 3638 28174
rect 3672 28140 3706 28174
rect 3740 28140 3774 28174
rect 3808 28140 3842 28174
rect 3876 28140 3910 28174
rect 3944 28140 3978 28174
rect 4012 28140 4046 28174
rect 4080 28140 4114 28174
rect 4148 28140 4182 28174
rect 4216 28140 4250 28174
rect 4284 28140 4318 28174
rect 4352 28140 4386 28174
rect 4420 28140 4454 28174
rect 4488 28140 4522 28174
rect 4556 28140 4590 28174
rect 4624 28140 4658 28174
rect 4692 28140 4726 28174
rect 4760 28140 4794 28174
rect 4828 28140 4862 28174
rect 4896 28140 4930 28174
rect 4964 28140 4998 28174
rect 5032 28140 5066 28174
rect 5100 28140 5134 28174
rect 5168 28140 5202 28174
rect 5236 28140 5270 28174
rect 5304 28140 5338 28174
rect 5372 28140 5406 28174
rect 5440 28140 5474 28174
rect 5508 28140 5542 28174
rect 5576 28140 5610 28174
rect 5644 28140 5678 28174
rect 5712 28140 5746 28174
rect 5780 28140 5814 28174
rect 5848 28140 5882 28174
rect 5916 28140 5950 28174
rect 5984 28140 6018 28174
rect 6052 28140 6086 28174
rect 6120 28140 6154 28174
rect 6188 28140 6222 28174
rect 6256 28140 6290 28174
rect 6324 28140 6358 28174
rect 6392 28140 6426 28174
rect 6460 28140 6494 28174
rect 6528 28140 6562 28174
rect 6596 28140 6630 28174
rect 6664 28140 6698 28174
rect 6732 28140 6766 28174
rect 6800 28140 6834 28174
rect 6868 28140 6902 28174
rect 6936 28140 6970 28174
rect 7004 28140 7038 28174
rect 7072 28140 7106 28174
rect 7140 28140 7174 28174
rect 7208 28140 7242 28174
rect 7276 28140 7310 28174
rect 7344 28140 7378 28174
rect 7412 28140 7446 28174
rect 7480 28140 7514 28174
rect 7548 28140 7582 28174
rect 7616 28140 7650 28174
rect 7684 28140 7780 28174
rect 4008 26082 4042 26116
rect 4008 26014 4042 26048
rect 4008 25946 4042 25980
rect 4008 25878 4042 25912
rect 4008 25810 4042 25844
rect 4008 25742 4042 25776
rect 4008 25674 4042 25708
rect 4008 25606 4042 25640
rect 4008 25538 4042 25572
rect 4008 25470 4042 25504
rect 4008 25402 4042 25436
rect 4008 25334 4042 25368
rect 4008 25266 4042 25300
rect 4008 25198 4042 25232
rect 4008 25130 4042 25164
rect 4008 25062 4042 25096
rect 4008 24994 4042 25028
rect 4008 24926 4042 24960
rect 4008 24858 4042 24892
rect 4008 24790 4042 24824
rect 4008 24718 4042 24756
rect 5946 26082 5980 26116
rect 5946 26014 5980 26048
rect 5946 25946 5980 25980
rect 5946 25878 5980 25912
rect 5946 25810 5980 25844
rect 5946 25742 5980 25776
rect 5946 25674 5980 25708
rect 5946 25606 5980 25640
rect 5946 25538 5980 25572
rect 5946 25470 5980 25504
rect 5946 25402 5980 25436
rect 5946 25334 5980 25368
rect 5946 25266 5980 25300
rect 5946 25198 5980 25232
rect 5946 25130 5980 25164
rect 5946 25062 5980 25096
rect 5946 24994 5980 25028
rect 5946 24926 5980 24960
rect 5946 24858 5980 24892
rect 5946 24790 5980 24824
rect 5946 24718 5980 24756
rect 4460 24150 4528 24184
rect 4562 24150 4596 24184
rect 4630 24150 4664 24184
rect 4698 24150 4732 24184
rect 4766 24150 4800 24184
rect 4834 24150 4868 24184
rect 4902 24150 4936 24184
rect 4970 24150 5004 24184
rect 5038 24150 5072 24184
rect 5106 24150 5140 24184
rect 5174 24150 5208 24184
rect 5242 24150 5276 24184
rect 5310 24150 5344 24184
rect 5378 24150 5412 24184
rect 5446 24150 5480 24184
rect 5514 24150 5548 24184
rect 5582 24150 5616 24184
rect 5650 24150 5684 24184
rect 5718 24150 5752 24184
rect 5786 24150 5892 24184
rect 4460 24110 4494 24150
rect 4460 23956 4494 24076
rect 5858 24116 5892 24150
rect 5858 24048 5892 24082
rect 4460 23888 4494 23922
rect 4460 23820 4494 23854
rect 5858 23980 5892 24014
rect 5858 23912 5892 23946
rect 5858 23844 5892 23878
rect 4460 23752 4494 23786
rect 4460 23684 4494 23718
rect 5858 23776 5892 23810
rect 4460 23616 4494 23650
rect 4460 23548 4494 23582
rect 4460 23480 4494 23514
rect 4460 23412 4494 23446
rect 4460 23344 4494 23378
rect 4460 23276 4494 23310
rect 4460 23208 4494 23242
rect 4460 23140 4494 23174
rect 4460 23072 4494 23106
rect 4460 23004 4494 23038
rect 4460 22936 4494 22970
rect 4460 22868 4494 22902
rect 4460 22800 4494 22834
rect 4460 22732 4494 22766
rect 4460 22664 4494 22698
rect 4460 22596 4494 22630
rect 4460 22528 4494 22562
rect 4460 22460 4494 22494
rect 4460 22392 4494 22426
rect 4460 22324 4494 22358
rect 4460 22256 4494 22290
rect 4460 22188 4494 22222
rect 4460 22120 4494 22154
rect 4460 22052 4494 22086
rect 4460 21984 4494 22018
rect 4460 21916 4494 21950
rect 4460 21848 4494 21882
rect 4460 21780 4494 21814
rect 4460 21712 4494 21746
rect 4460 21644 4494 21678
rect 4460 21576 4494 21610
rect 4460 21508 4494 21542
rect 4460 21440 4494 21474
rect 4460 21372 4494 21406
rect 4460 21304 4494 21338
rect 4460 21236 4494 21270
rect 4460 21168 4494 21202
rect 4460 21100 4494 21134
rect 4460 21032 4494 21066
rect 4460 20964 4494 20998
rect 4460 20896 4494 20930
rect 4460 20828 4494 20862
rect 4460 20760 4494 20794
rect 4460 20692 4494 20726
rect 4460 20624 4494 20658
rect 4460 20556 4494 20590
rect 4460 20488 4494 20522
rect 4460 20420 4494 20454
rect 4460 20352 4494 20386
rect 4460 20284 4494 20318
rect 4460 20216 4494 20250
rect 4460 20148 4494 20182
rect 4460 20080 4494 20114
rect 4460 20012 4494 20046
rect 4460 19944 4494 19978
rect 4460 19876 4494 19910
rect 4460 19808 4494 19842
rect 4460 19740 4494 19774
rect 4460 19672 4494 19706
rect 4460 19604 4494 19638
rect 4460 19536 4494 19570
rect 4460 19468 4494 19502
rect 5858 23708 5892 23742
rect 5858 23640 5892 23674
rect 5858 23572 5892 23606
rect 5858 23504 5892 23538
rect 5858 23436 5892 23470
rect 5858 23368 5892 23402
rect 5858 23300 5892 23334
rect 5858 23232 5892 23266
rect 5858 23164 5892 23198
rect 5858 23096 5892 23130
rect 5858 23028 5892 23062
rect 5858 22960 5892 22994
rect 5858 22892 5892 22926
rect 5858 22824 5892 22858
rect 5858 22756 5892 22790
rect 5858 22688 5892 22722
rect 5858 22620 5892 22654
rect 5858 22552 5892 22586
rect 5858 22484 5892 22518
rect 5858 22416 5892 22450
rect 5858 22348 5892 22382
rect 5858 22280 5892 22314
rect 5858 22212 5892 22246
rect 5858 22144 5892 22178
rect 5858 22076 5892 22110
rect 5858 22008 5892 22042
rect 5858 21940 5892 21974
rect 5858 21872 5892 21906
rect 5858 21804 5892 21838
rect 5858 21736 5892 21770
rect 5858 21668 5892 21702
rect 5858 21600 5892 21634
rect 5858 21532 5892 21566
rect 5858 21464 5892 21498
rect 7326 21485 7420 21519
rect 7454 21485 7488 21519
rect 7522 21485 7556 21519
rect 7590 21485 7624 21519
rect 7658 21485 7692 21519
rect 5858 21396 5892 21430
rect 5858 21328 5892 21362
rect 5858 21260 5892 21294
rect 5858 21192 5892 21226
rect 5858 21124 5892 21158
rect 5858 21056 5892 21090
rect 5858 20988 5892 21022
rect 5858 20920 5892 20954
rect 5858 20852 5892 20886
rect 5858 20784 5892 20818
rect 5858 20716 5892 20750
rect 5858 20648 5892 20682
rect 5858 20580 5892 20614
rect 5858 20512 5892 20546
rect 5858 20444 5892 20478
rect 5858 20376 5892 20410
rect 5858 20308 5892 20342
rect 5858 20240 5892 20274
rect 5858 20172 5892 20206
rect 5858 20104 5892 20138
rect 5858 20036 5892 20070
rect 5858 19968 5892 20002
rect 5858 19900 5892 19934
rect 5858 19832 5892 19866
rect 5858 19764 5892 19798
rect 5858 19696 5892 19730
rect 4460 19400 4494 19434
rect 5858 19628 5892 19662
rect 5858 19560 5892 19594
rect 5858 19492 5892 19526
rect 5858 19424 5892 19458
rect 4460 19332 4494 19366
rect 4460 19264 4494 19298
rect 4460 19196 4494 19230
rect 4460 19128 4494 19162
rect 4460 19060 4494 19094
rect 5858 19356 5892 19390
rect 5858 19288 5892 19322
rect 5858 19220 5892 19254
rect 5858 19152 5892 19186
rect 5858 19084 5892 19118
rect 4460 18992 4494 19026
rect 5858 19016 5892 19050
rect 4460 18924 4494 18958
rect 4460 18856 4494 18890
rect 4460 18788 4494 18822
rect 5858 18948 5892 18982
rect 5858 18880 5892 18914
rect 5858 18812 5892 18846
rect 4460 18720 4494 18754
rect 4460 18652 4494 18686
rect 4460 18584 4494 18618
rect 4460 18516 4494 18550
rect 5858 18744 5892 18778
rect 5858 18676 5892 18710
rect 5858 18608 5892 18642
rect 5858 18516 5892 18574
rect 4460 18482 4566 18516
rect 4600 18482 4634 18516
rect 4668 18482 4702 18516
rect 4736 18482 4770 18516
rect 4804 18482 4838 18516
rect 4872 18482 4906 18516
rect 4940 18482 4974 18516
rect 5008 18482 5042 18516
rect 5076 18482 5110 18516
rect 5144 18482 5178 18516
rect 5212 18482 5246 18516
rect 5280 18482 5314 18516
rect 5348 18482 5382 18516
rect 5416 18482 5450 18516
rect 5484 18482 5518 18516
rect 5552 18482 5586 18516
rect 5620 18482 5654 18516
rect 5688 18482 5722 18516
rect 5756 18482 5790 18516
rect 5824 18482 5892 18516
rect 2822 18255 2890 18289
rect 2924 18255 2958 18289
rect 2992 18255 3026 18289
rect 3060 18255 3094 18289
rect 3128 18255 3162 18289
rect 3196 18255 3230 18289
rect 3264 18255 3298 18289
rect 3332 18255 3366 18289
rect 3400 18255 3434 18289
rect 3468 18255 3502 18289
rect 3536 18255 3570 18289
rect 3604 18255 3638 18289
rect 3672 18255 3706 18289
rect 3740 18255 3774 18289
rect 3808 18255 3842 18289
rect 3876 18255 3910 18289
rect 3944 18255 3978 18289
rect 4012 18255 4046 18289
rect 4080 18255 4114 18289
rect 4148 18255 4182 18289
rect 4216 18255 4250 18289
rect 4284 18255 4318 18289
rect 4352 18255 4386 18289
rect 4420 18255 4454 18289
rect 4488 18255 4522 18289
rect 4556 18255 4590 18289
rect 4624 18255 4658 18289
rect 4692 18255 4726 18289
rect 4760 18255 4794 18289
rect 4828 18255 4862 18289
rect 4896 18255 4930 18289
rect 4964 18255 4998 18289
rect 5032 18255 5066 18289
rect 5100 18255 5134 18289
rect 5168 18255 5202 18289
rect 5236 18255 5270 18289
rect 5304 18255 5338 18289
rect 5372 18255 5406 18289
rect 5440 18255 5474 18289
rect 5508 18255 5542 18289
rect 5576 18255 5610 18289
rect 5644 18255 5678 18289
rect 5712 18255 5746 18289
rect 5780 18255 5814 18289
rect 5848 18255 5882 18289
rect 5916 18255 5950 18289
rect 5984 18255 6018 18289
rect 6052 18255 6086 18289
rect 6120 18255 6154 18289
rect 6188 18255 6222 18289
rect 6256 18255 6290 18289
rect 6324 18255 6358 18289
rect 6392 18255 6426 18289
rect 6460 18255 6494 18289
rect 6528 18255 6562 18289
rect 6596 18255 6630 18289
rect 6664 18255 6784 18289
rect 2822 18197 2856 18255
rect 2822 18083 2856 18163
rect 2822 18015 2856 18049
rect 6750 18221 6784 18255
rect 6750 18153 6784 18187
rect 6750 18085 6784 18119
rect 2822 17947 2856 17981
rect 2822 17879 2856 17913
rect 2822 17811 2856 17845
rect 2822 17743 2856 17777
rect 2822 17675 2856 17709
rect 2822 17607 2856 17641
rect 2822 17539 2856 17573
rect 2822 17471 2856 17505
rect 2822 17403 2856 17437
rect 2822 17335 2856 17369
rect 2822 17267 2856 17301
rect 2822 17199 2856 17233
rect 2822 17131 2856 17165
rect 2822 17063 2856 17097
rect 2822 16995 2856 17029
rect 2822 16927 2856 16961
rect 2822 16859 2856 16893
rect 2822 16791 2856 16825
rect 2822 16723 2856 16757
rect 2822 16655 2856 16689
rect 2822 16587 2856 16621
rect 2822 16519 2856 16553
rect 2822 16451 2856 16485
rect 2822 16383 2856 16417
rect 2822 16315 2856 16349
rect 2822 16247 2856 16281
rect 2822 16179 2856 16213
rect 2822 16111 2856 16145
rect 2822 16043 2856 16077
rect 2822 15975 2856 16009
rect 2822 15907 2856 15941
rect 2822 15839 2856 15873
rect 2822 15771 2856 15805
rect 2822 15703 2856 15737
rect 2822 15635 2856 15669
rect 2822 15567 2856 15601
rect 2822 15499 2856 15533
rect 2822 15431 2856 15465
rect 2822 15363 2856 15397
rect 2822 15295 2856 15329
rect 2822 15227 2856 15261
rect 2822 15159 2856 15193
rect 2822 15091 2856 15125
rect 2822 15023 2856 15057
rect 2822 14955 2856 14989
rect 2822 14887 2856 14921
rect 2822 14819 2856 14853
rect 2822 14751 2856 14785
rect 2822 14683 2856 14717
rect 2822 14615 2856 14649
rect 2822 14547 2856 14581
rect 6750 18017 6784 18051
rect 6750 17949 6784 17983
rect 6750 17881 6784 17915
rect 6750 17813 6784 17847
rect 6750 17745 6784 17779
rect 6750 17677 6784 17711
rect 6750 17609 6784 17643
rect 6750 17541 6784 17575
rect 6750 17473 6784 17507
rect 6750 17405 6784 17439
rect 6750 17337 6784 17371
rect 6750 17269 6784 17303
rect 6750 17201 6784 17235
rect 6750 17133 6784 17167
rect 6750 17065 6784 17099
rect 6750 16997 6784 17031
rect 6750 16929 6784 16963
rect 6750 16861 6784 16895
rect 6750 16793 6784 16827
rect 6750 16725 6784 16759
rect 6750 16657 6784 16691
rect 6750 16589 6784 16623
rect 6750 16521 6784 16555
rect 6750 16453 6784 16487
rect 6750 16385 6784 16419
rect 6750 16317 6784 16351
rect 6750 16249 6784 16283
rect 6750 16181 6784 16215
rect 6750 16113 6784 16147
rect 6750 16045 6784 16079
rect 6750 15977 6784 16011
rect 6750 15909 6784 15943
rect 6750 15841 6784 15875
rect 6750 15773 6784 15807
rect 6750 15705 6784 15739
rect 6750 15637 6784 15671
rect 6750 15569 6784 15603
rect 6750 15501 6784 15535
rect 6750 15433 6784 15467
rect 6750 15365 6784 15399
rect 6750 15297 6784 15331
rect 6750 15229 6784 15263
rect 6750 15161 6784 15195
rect 6750 15093 6784 15127
rect 6750 15025 6784 15059
rect 6750 14957 6784 14991
rect 6750 14889 6784 14923
rect 6750 14821 6784 14855
rect 6750 14753 6784 14787
rect 6750 14685 6784 14719
rect 6750 14617 6784 14651
rect 2822 14479 2856 14513
rect 2822 14411 2856 14445
rect 2822 14343 2856 14377
rect 6750 14549 6784 14583
rect 6750 14481 6784 14515
rect 6750 14413 6784 14447
rect 6750 14343 6784 14379
rect 2822 14309 2942 14343
rect 2976 14309 3010 14343
rect 3044 14309 3078 14343
rect 3112 14309 3146 14343
rect 3180 14309 3214 14343
rect 3248 14309 3282 14343
rect 3316 14309 3350 14343
rect 3384 14309 3418 14343
rect 3452 14309 3486 14343
rect 3520 14309 3554 14343
rect 3588 14309 3622 14343
rect 3656 14309 3690 14343
rect 3724 14309 3758 14343
rect 3792 14309 3826 14343
rect 3860 14309 3894 14343
rect 3928 14309 3962 14343
rect 3996 14309 4030 14343
rect 4064 14309 4098 14343
rect 4132 14309 4166 14343
rect 4200 14309 4234 14343
rect 4268 14309 4302 14343
rect 4336 14309 4370 14343
rect 4404 14309 4438 14343
rect 4472 14309 4506 14343
rect 4540 14309 4574 14343
rect 4608 14309 4642 14343
rect 4676 14309 4710 14343
rect 4744 14309 4778 14343
rect 4812 14309 4846 14343
rect 4880 14309 4914 14343
rect 4948 14309 4982 14343
rect 5016 14309 5050 14343
rect 5084 14309 5118 14343
rect 5152 14309 5186 14343
rect 5220 14309 5254 14343
rect 5288 14309 5322 14343
rect 5356 14309 5390 14343
rect 5424 14309 5458 14343
rect 5492 14309 5526 14343
rect 5560 14309 5594 14343
rect 5628 14309 5662 14343
rect 5696 14309 5730 14343
rect 5764 14309 5798 14343
rect 5832 14309 5866 14343
rect 5900 14309 5934 14343
rect 5968 14309 6002 14343
rect 6036 14309 6070 14343
rect 6104 14309 6138 14343
rect 6172 14309 6206 14343
rect 6240 14309 6274 14343
rect 6308 14309 6342 14343
rect 6376 14309 6410 14343
rect 6444 14309 6478 14343
rect 6512 14309 6546 14343
rect 6580 14309 6614 14343
rect 6648 14309 6682 14343
rect 6716 14309 6784 14343
<< mvpsubdiffcont >>
rect 3154 39580 3188 39614
rect 3222 39580 3256 39614
rect 3290 39580 3324 39614
rect 3358 39580 3392 39614
rect 3426 39580 3460 39614
rect 3494 39580 3528 39614
rect 3562 39580 3596 39614
rect 3630 39580 3664 39614
rect 3698 39580 3732 39614
rect 3766 39580 3800 39614
rect 3834 39580 3868 39614
rect 3902 39580 3936 39614
rect 3970 39580 4004 39614
rect 4038 39580 4072 39614
rect 4106 39580 4140 39614
rect 4174 39580 4208 39614
rect 4242 39580 4276 39614
rect 4310 39580 4344 39614
rect 4378 39580 4412 39614
rect 4446 39580 4480 39614
rect 4514 39580 4548 39614
rect 4582 39580 4616 39614
rect 4650 39580 4684 39614
rect 4718 39580 4752 39614
rect 4786 39580 4820 39614
rect 4854 39580 4888 39614
rect 4922 39580 4956 39614
rect 4990 39580 5024 39614
rect 5058 39580 5092 39614
rect 5126 39580 5160 39614
rect 5194 39580 5228 39614
rect 5262 39580 5296 39614
rect 3082 39512 3116 39546
rect 3082 39444 3116 39478
rect 5330 39474 5364 39508
rect 3082 39376 3116 39410
rect 3082 39308 3116 39342
rect 3082 39240 3116 39274
rect 3082 39172 3116 39206
rect 3082 39104 3116 39138
rect 3082 39036 3116 39070
rect 3082 38968 3116 39002
rect 3082 38900 3116 38934
rect 3082 38832 3116 38866
rect 3082 38764 3116 38798
rect 3082 38696 3116 38730
rect 3082 38628 3116 38662
rect 3082 38560 3116 38594
rect 3082 38492 3116 38526
rect 3082 38424 3116 38458
rect 3082 38356 3116 38390
rect 3082 38288 3116 38322
rect 3082 38220 3116 38254
rect 3082 38152 3116 38186
rect 3082 38084 3116 38118
rect 3082 38016 3116 38050
rect 3082 37948 3116 37982
rect 3082 37880 3116 37914
rect 3082 37812 3116 37846
rect 3082 37744 3116 37778
rect 3082 37676 3116 37710
rect 3082 37608 3116 37642
rect 3082 37540 3116 37574
rect 3082 37472 3116 37506
rect 3082 37404 3116 37438
rect 3082 37336 3116 37370
rect 3082 37268 3116 37302
rect 3082 37200 3116 37234
rect 3082 37132 3116 37166
rect 3082 37064 3116 37098
rect 3082 36996 3116 37030
rect 3082 36928 3116 36962
rect 3082 36860 3116 36894
rect 3082 36792 3116 36826
rect 3082 36724 3116 36758
rect 3082 36656 3116 36690
rect 3082 36588 3116 36622
rect 3082 36520 3116 36554
rect 3082 36452 3116 36486
rect 3082 36384 3116 36418
rect 3082 36316 3116 36350
rect 3082 36248 3116 36282
rect 3082 36180 3116 36214
rect 3082 36112 3116 36146
rect 3082 36044 3116 36078
rect 3082 35976 3116 36010
rect 3082 35908 3116 35942
rect 3082 35840 3116 35874
rect 3082 35772 3116 35806
rect 3082 35704 3116 35738
rect 3082 35636 3116 35670
rect 3082 35568 3116 35602
rect 3082 35500 3116 35534
rect 3082 35432 3116 35466
rect 3082 35364 3116 35398
rect 3082 35296 3116 35330
rect 3082 35228 3116 35262
rect 3082 35160 3116 35194
rect 3082 35092 3116 35126
rect 3082 35024 3116 35058
rect 3082 34956 3116 34990
rect 3082 34888 3116 34922
rect 3082 34820 3116 34854
rect 3082 34752 3116 34786
rect 3082 34684 3116 34718
rect 3082 34616 3116 34650
rect 3082 34548 3116 34582
rect 3082 34480 3116 34514
rect 3082 34412 3116 34446
rect 3082 34344 3116 34378
rect 3082 34276 3116 34310
rect 3082 34208 3116 34242
rect 3082 34140 3116 34174
rect 3082 34072 3116 34106
rect 3082 34004 3116 34038
rect 3082 33936 3116 33970
rect 3082 33868 3116 33902
rect 3082 33800 3116 33834
rect 3082 33732 3116 33766
rect 3082 33664 3116 33698
rect 3082 33596 3116 33630
rect 3082 33528 3116 33562
rect 3082 33460 3116 33494
rect 3082 33392 3116 33426
rect 3082 33324 3116 33358
rect 3082 33256 3116 33290
rect 3082 33188 3116 33222
rect 3082 33120 3116 33154
rect 3082 33052 3116 33086
rect 3082 32984 3116 33018
rect 3082 32916 3116 32950
rect 3082 32848 3116 32882
rect 3082 32780 3116 32814
rect 3082 32712 3116 32746
rect 3082 32644 3116 32678
rect 3082 32576 3116 32610
rect 3082 32508 3116 32542
rect 3082 32440 3116 32474
rect 3082 32372 3116 32406
rect 3082 32304 3116 32338
rect 3082 32236 3116 32270
rect 3082 32168 3116 32202
rect 3082 32100 3116 32134
rect 3082 32032 3116 32066
rect 3082 31964 3116 31998
rect 3082 31896 3116 31930
rect 3082 31828 3116 31862
rect 3082 31760 3116 31794
rect 3082 31692 3116 31726
rect 3082 31624 3116 31658
rect 3082 31556 3116 31590
rect 3082 31488 3116 31522
rect 3082 31420 3116 31454
rect 3082 31352 3116 31386
rect 3082 31284 3116 31318
rect 3082 31216 3116 31250
rect 3082 31148 3116 31182
rect 3082 31080 3116 31114
rect 3082 31012 3116 31046
rect 3082 30944 3116 30978
rect 3082 30876 3116 30910
rect 3082 30808 3116 30842
rect 3082 30740 3116 30774
rect 3082 30672 3116 30706
rect 3082 30604 3116 30638
rect 3082 30536 3116 30570
rect 3082 30468 3116 30502
rect 3082 30400 3116 30434
rect 5330 39406 5364 39440
rect 5330 39338 5364 39372
rect 5330 39270 5364 39304
rect 5330 39202 5364 39236
rect 5330 39134 5364 39168
rect 5330 39066 5364 39100
rect 5330 38998 5364 39032
rect 5330 38930 5364 38964
rect 5330 38862 5364 38896
rect 5330 38794 5364 38828
rect 5330 38726 5364 38760
rect 5330 38658 5364 38692
rect 5330 38590 5364 38624
rect 5330 38522 5364 38556
rect 5330 38454 5364 38488
rect 5330 38386 5364 38420
rect 5330 38318 5364 38352
rect 5330 38250 5364 38284
rect 5330 38182 5364 38216
rect 5330 38114 5364 38148
rect 5330 38046 5364 38080
rect 5330 37978 5364 38012
rect 5330 37910 5364 37944
rect 5330 37842 5364 37876
rect 5330 37774 5364 37808
rect 5330 37706 5364 37740
rect 5330 37638 5364 37672
rect 5330 37570 5364 37604
rect 5330 37502 5364 37536
rect 5330 37434 5364 37468
rect 5330 37366 5364 37400
rect 5330 37298 5364 37332
rect 5330 37230 5364 37264
rect 5330 37162 5364 37196
rect 5330 37094 5364 37128
rect 5330 37026 5364 37060
rect 5330 36958 5364 36992
rect 5330 36890 5364 36924
rect 5330 36822 5364 36856
rect 5330 36754 5364 36788
rect 5330 36686 5364 36720
rect 5330 36618 5364 36652
rect 5330 36550 5364 36584
rect 5330 36482 5364 36516
rect 5330 36414 5364 36448
rect 5330 36346 5364 36380
rect 5330 36278 5364 36312
rect 5330 36210 5364 36244
rect 5330 36142 5364 36176
rect 5330 36074 5364 36108
rect 5330 36006 5364 36040
rect 5330 35938 5364 35972
rect 5330 35870 5364 35904
rect 5330 35802 5364 35836
rect 5330 35734 5364 35768
rect 5330 35666 5364 35700
rect 5330 35598 5364 35632
rect 5330 35530 5364 35564
rect 5330 35462 5364 35496
rect 5330 35394 5364 35428
rect 5330 35326 5364 35360
rect 5330 35258 5364 35292
rect 5330 35190 5364 35224
rect 5330 35122 5364 35156
rect 5330 35054 5364 35088
rect 5330 34986 5364 35020
rect 5330 34918 5364 34952
rect 5330 34850 5364 34884
rect 5330 34782 5364 34816
rect 5330 34714 5364 34748
rect 5330 34646 5364 34680
rect 5330 34578 5364 34612
rect 5330 34510 5364 34544
rect 5330 34442 5364 34476
rect 5330 34374 5364 34408
rect 5330 34306 5364 34340
rect 5330 34238 5364 34272
rect 5330 34170 5364 34204
rect 5330 34102 5364 34136
rect 5330 34034 5364 34068
rect 5330 33966 5364 34000
rect 5330 33898 5364 33932
rect 5330 33830 5364 33864
rect 5330 33762 5364 33796
rect 5330 33694 5364 33728
rect 5330 33626 5364 33660
rect 5330 33558 5364 33592
rect 5330 33490 5364 33524
rect 5330 33422 5364 33456
rect 5330 33354 5364 33388
rect 5330 33286 5364 33320
rect 5330 33218 5364 33252
rect 5330 33150 5364 33184
rect 5330 33082 5364 33116
rect 5330 33014 5364 33048
rect 5330 32946 5364 32980
rect 5330 32878 5364 32912
rect 5330 32810 5364 32844
rect 5330 32742 5364 32776
rect 5330 32674 5364 32708
rect 5330 32606 5364 32640
rect 5330 32538 5364 32572
rect 5330 32470 5364 32504
rect 5330 32402 5364 32436
rect 5330 32334 5364 32368
rect 5330 32266 5364 32300
rect 5330 32198 5364 32232
rect 5330 32130 5364 32164
rect 5330 32062 5364 32096
rect 5330 31994 5364 32028
rect 5330 31926 5364 31960
rect 5330 31858 5364 31892
rect 5330 31790 5364 31824
rect 5330 31722 5364 31756
rect 5330 31654 5364 31688
rect 5330 31586 5364 31620
rect 5330 31518 5364 31552
rect 5330 31450 5364 31484
rect 5330 31382 5364 31416
rect 5330 31314 5364 31348
rect 5330 31246 5364 31280
rect 5330 31178 5364 31212
rect 5330 31110 5364 31144
rect 5330 31042 5364 31076
rect 5330 30974 5364 31008
rect 5330 30906 5364 30940
rect 5330 30838 5364 30872
rect 5330 30770 5364 30804
rect 5330 30702 5364 30736
rect 5330 30634 5364 30668
rect 5330 30566 5364 30600
rect 5330 30498 5364 30532
rect 5330 30430 5364 30464
rect 3082 30332 3116 30366
rect 5330 30362 5364 30396
rect 3082 30264 3116 30298
rect 3082 30196 3116 30230
rect 5664 30163 5698 30197
rect 5735 30163 5769 30197
rect 5806 30163 5840 30197
rect 5877 30163 5911 30197
rect 5948 30163 5982 30197
rect 6019 30163 6053 30197
rect 6090 30163 6124 30197
rect 6161 30163 6195 30197
rect 6232 30163 6266 30197
rect 6303 30163 6337 30197
rect 6374 30163 6408 30197
rect 6444 30163 6478 30197
rect 6514 30163 6548 30197
rect 6584 30163 6618 30197
rect 6654 30163 6688 30197
rect 6724 30163 6758 30197
rect 6794 30163 6828 30197
rect 6864 30163 6898 30197
rect 6934 30163 6968 30197
rect 7004 30163 7038 30197
rect 7074 30163 7108 30197
rect 7144 30163 7178 30197
rect 7214 30163 7248 30197
rect 7284 30163 7318 30197
rect 7354 30163 7388 30197
rect 7424 30163 7458 30197
rect 3082 30128 3116 30162
rect 3082 30060 3116 30094
rect 3082 29992 3116 30026
rect 3082 29924 3116 29958
rect 3082 29856 3116 29890
rect 3082 29788 3116 29822
rect 3082 29720 3116 29754
rect 5640 29964 5674 29998
rect 5640 29896 5674 29930
rect 5640 29828 5674 29862
rect 5640 29760 5674 29794
rect 3082 29652 3116 29686
rect 3082 29584 3116 29618
rect 5640 29692 5674 29726
rect 5640 29624 5674 29658
rect 3082 29516 3116 29550
rect 3082 29448 3116 29482
rect 3082 29380 3116 29414
rect 3082 29312 3116 29346
rect 5640 29556 5674 29590
rect 5640 29488 5674 29522
rect 5640 29420 5674 29454
rect 5640 29352 5674 29386
rect 3082 29244 3116 29278
rect 5640 29284 5674 29318
rect 3082 29176 3116 29210
rect 5640 29216 5674 29250
rect 3082 29108 3116 29142
rect 5640 29148 5674 29182
rect 3082 29040 3116 29074
rect 5640 29080 5674 29114
rect 3082 28972 3116 29006
rect 3082 28904 3116 28938
rect 3082 28836 3116 28870
rect 3082 28768 3116 28802
rect 5640 29012 5674 29046
rect 5640 28944 5674 28978
rect 5640 28876 5674 28910
rect 5640 28808 5674 28842
rect 3082 28700 3116 28734
rect 3082 28632 3116 28666
rect 3082 28564 3116 28598
rect 3082 28496 3116 28530
rect 5640 28740 5674 28774
rect 5640 28672 5674 28706
rect 5640 28604 5674 28638
rect 5640 28536 5674 28570
rect 5640 28468 5674 28502
rect 3150 28400 3184 28434
rect 3218 28400 3252 28434
rect 3286 28400 3320 28434
rect 3354 28400 3388 28434
rect 3422 28400 3456 28434
rect 3490 28400 3524 28434
rect 3558 28400 3592 28434
rect 3626 28400 3660 28434
rect 3694 28400 3728 28434
rect 3762 28400 3796 28434
rect 3830 28400 3864 28434
rect 3898 28400 3932 28434
rect 3966 28400 4000 28434
rect 4034 28400 4068 28434
rect 4102 28400 4136 28434
rect 4170 28400 4204 28434
rect 4238 28400 4272 28434
rect 4306 28400 4340 28434
rect 4374 28400 4408 28434
rect 4442 28400 4476 28434
rect 4510 28400 4544 28434
rect 4578 28400 4612 28434
rect 4646 28400 4680 28434
rect 4714 28400 4748 28434
rect 4782 28400 4816 28434
rect 4850 28400 4884 28434
rect 4918 28400 4952 28434
rect 4986 28400 5020 28434
rect 5054 28400 5088 28434
rect 5122 28400 5156 28434
rect 5190 28400 5224 28434
rect 5258 28400 5292 28434
rect 5326 28400 5360 28434
rect 5394 28400 5428 28434
rect 5462 28400 5496 28434
rect 5530 28400 5564 28434
rect 2678 25651 2712 25685
rect 2746 25651 2780 25685
rect 2814 25651 2848 25685
rect 2882 25651 2916 25685
rect 2950 25651 2984 25685
rect 3018 25651 3052 25685
rect 3086 25651 3120 25685
rect 3154 25651 3188 25685
rect 3222 25651 3256 25685
rect 3290 25651 3324 25685
rect 3358 25651 3392 25685
rect 3426 25651 3460 25685
rect 3494 25651 3528 25685
rect 3562 25651 3596 25685
rect 3630 25651 3664 25685
rect 3698 25575 3732 25609
rect 3698 25507 3732 25541
rect 3698 25439 3732 25473
rect 3698 25371 3732 25405
rect 3698 25303 3732 25337
rect 3698 25235 3732 25269
rect 3698 25167 3732 25201
rect 3698 25099 3732 25133
rect 3698 25031 3732 25065
rect 3698 24963 3732 24997
rect 3698 24895 3732 24929
rect 3698 24827 3732 24861
rect 3698 24759 3732 24793
rect 3698 24691 3732 24725
rect 3698 24623 3732 24657
rect 3698 24555 3732 24589
rect 3698 24487 3732 24521
rect 3698 24419 3732 24453
rect 3698 24351 3732 24385
rect 3698 24283 3732 24317
rect 3698 24215 3732 24249
rect 3698 24147 3732 24181
rect 3698 24079 3732 24113
rect 3698 24011 3732 24045
rect 3698 23943 3732 23977
rect 3698 23875 3732 23909
rect 3698 23807 3732 23841
rect 3698 23739 3732 23773
rect 3698 23671 3732 23705
rect 3698 23603 3732 23637
rect 3698 23535 3732 23569
rect 3698 23467 3732 23501
rect 3698 23399 3732 23433
rect 3698 23331 3732 23365
rect 3698 23263 3732 23297
rect 3698 23195 3732 23229
rect 3698 23127 3732 23161
rect 3698 23059 3732 23093
rect 3698 22991 3732 23025
rect 3698 22923 3732 22957
rect 3698 22855 3732 22889
rect 3698 22787 3732 22821
rect 3698 22719 3732 22753
rect 3698 22651 3732 22685
rect 3698 22583 3732 22617
rect 3698 22515 3732 22549
rect 3698 22447 3732 22481
rect 3698 22379 3732 22413
rect 3698 22311 3732 22345
rect 3698 22243 3732 22277
rect 3698 22175 3732 22209
rect 3698 22107 3732 22141
rect 3698 22039 3732 22073
rect 3698 21971 3732 22005
rect 3698 21903 3732 21937
rect 3698 21835 3732 21869
rect 3698 21767 3732 21801
rect 3698 21699 3732 21733
rect 3698 21631 3732 21665
rect 3698 21563 3732 21597
rect 3698 21495 3732 21529
rect 3698 21427 3732 21461
rect 3698 21359 3732 21393
rect 3698 21291 3732 21325
rect 3698 21223 3732 21257
rect 3698 21155 3732 21189
rect 3698 21087 3732 21121
rect 3698 21019 3732 21053
rect 3698 20951 3732 20985
rect 3698 20883 3732 20917
rect 3698 20815 3732 20849
rect 3698 20747 3732 20781
rect 3698 20679 3732 20713
rect 3698 20611 3732 20645
rect 3698 20543 3732 20577
rect 3698 20475 3732 20509
rect 3698 20407 3732 20441
rect 3698 20339 3732 20373
rect 3698 20271 3732 20305
rect 3698 20203 3732 20237
rect 3698 20135 3732 20169
rect 3698 20067 3732 20101
rect 3698 19999 3732 20033
rect 3698 19931 3732 19965
rect 3698 19863 3732 19897
rect 3698 19795 3732 19829
rect 3698 19727 3732 19761
rect 3698 19659 3732 19693
rect 3698 19591 3732 19625
rect 3698 19523 3732 19557
rect 3698 19455 3732 19489
rect 3698 19387 3732 19421
rect 3698 19319 3732 19353
rect 3698 19251 3732 19285
rect 3698 19183 3732 19217
rect 3698 19115 3732 19149
rect 3698 19047 3732 19081
rect 3698 18979 3732 19013
rect 3698 18911 3732 18945
rect 3698 18843 3732 18877
rect 3698 18775 3732 18809
rect 3698 18707 3732 18741
rect 3698 18639 3732 18673
rect 3698 18571 3732 18605
rect 3150 17995 3184 18029
rect 3218 17995 3252 18029
rect 3286 17995 3320 18029
rect 3354 17995 3388 18029
rect 3422 17995 3456 18029
rect 3490 17995 3524 18029
rect 3558 17995 3592 18029
rect 3626 17995 3660 18029
rect 3694 17995 3728 18029
rect 3762 17995 3796 18029
rect 3830 17995 3864 18029
rect 3898 17995 3932 18029
rect 3966 17995 4000 18029
rect 4034 17995 4068 18029
rect 4102 17995 4136 18029
rect 4170 17995 4204 18029
rect 4238 17995 4272 18029
rect 4306 17995 4340 18029
rect 4374 17995 4408 18029
rect 4442 17995 4476 18029
rect 4510 17995 4544 18029
rect 4578 17995 4612 18029
rect 4646 17995 4680 18029
rect 4714 17995 4748 18029
rect 4782 17995 4816 18029
rect 4850 17995 4884 18029
rect 4918 17995 4952 18029
rect 4986 17995 5020 18029
rect 5054 17995 5088 18029
rect 5122 17995 5156 18029
rect 5190 17995 5224 18029
rect 5258 17995 5292 18029
rect 5326 17995 5360 18029
rect 5394 17995 5428 18029
rect 5462 17995 5496 18029
rect 5530 17995 5564 18029
rect 5598 17995 5632 18029
rect 5666 17995 5700 18029
rect 5734 17995 5768 18029
rect 5802 17995 5836 18029
rect 5870 17995 5904 18029
rect 5938 17995 5972 18029
rect 6006 17995 6040 18029
rect 6074 17995 6108 18029
rect 6142 17995 6176 18029
rect 6210 17995 6244 18029
rect 6278 17995 6312 18029
rect 6346 17995 6380 18029
rect 3082 17901 3116 17935
rect 6476 17927 6510 17961
rect 3082 17833 3116 17867
rect 3082 17765 3116 17799
rect 3082 17697 3116 17731
rect 3082 17629 3116 17663
rect 3082 17561 3116 17595
rect 3082 17493 3116 17527
rect 3082 17425 3116 17459
rect 3082 17357 3116 17391
rect 3082 17289 3116 17323
rect 3082 17221 3116 17255
rect 3082 17153 3116 17187
rect 3082 17085 3116 17119
rect 3082 17017 3116 17051
rect 3082 16949 3116 16983
rect 3082 16881 3116 16915
rect 3082 16813 3116 16847
rect 3082 16745 3116 16779
rect 3082 16677 3116 16711
rect 3082 16609 3116 16643
rect 3082 16541 3116 16575
rect 3082 16473 3116 16507
rect 3082 16405 3116 16439
rect 3082 16337 3116 16371
rect 3082 16269 3116 16303
rect 3082 16201 3116 16235
rect 3082 16133 3116 16167
rect 3082 16065 3116 16099
rect 3082 15997 3116 16031
rect 6476 17859 6510 17893
rect 6476 17791 6510 17825
rect 6476 17723 6510 17757
rect 6476 17655 6510 17689
rect 6476 17587 6510 17621
rect 6476 17519 6510 17553
rect 6476 17451 6510 17485
rect 6476 17383 6510 17417
rect 6476 17315 6510 17349
rect 6476 17247 6510 17281
rect 6476 17179 6510 17213
rect 6476 17111 6510 17145
rect 6476 17043 6510 17077
rect 6211 16928 6245 16962
rect 6337 16928 6371 16962
rect 6211 16785 6245 16819
rect 6337 16785 6371 16819
rect 3695 16675 3729 16709
rect 3821 16675 3855 16709
rect 3695 16530 3729 16564
rect 3821 16530 3855 16564
rect 3695 16385 3729 16419
rect 3821 16385 3855 16419
rect 3695 16240 3729 16274
rect 3821 16240 3855 16274
rect 6211 16642 6245 16676
rect 6337 16642 6371 16676
rect 6211 16499 6245 16533
rect 6337 16499 6371 16533
rect 6211 16356 6245 16390
rect 6337 16356 6371 16390
rect 6211 16213 6245 16247
rect 6337 16213 6371 16247
rect 3695 16095 3729 16129
rect 3821 16095 3855 16129
rect 3082 15929 3116 15963
rect 6211 16070 6245 16104
rect 6337 16070 6371 16104
rect 3695 15950 3729 15984
rect 3821 15950 3855 15984
rect 3082 15861 3116 15895
rect 3082 15793 3116 15827
rect 3082 15725 3116 15759
rect 3695 15805 3729 15839
rect 3821 15805 3855 15839
rect 3082 15657 3116 15691
rect 3082 15589 3116 15623
rect 3082 15521 3116 15555
rect 3082 15453 3116 15487
rect 3082 15385 3116 15419
rect 3082 15317 3116 15351
rect 3082 15249 3116 15283
rect 3082 15181 3116 15215
rect 3082 15113 3116 15147
rect 3082 15045 3116 15079
rect 3082 14977 3116 15011
rect 3082 14909 3116 14943
rect 3082 14841 3116 14875
rect 3082 14773 3116 14807
rect 3082 14705 3116 14739
rect 3082 14637 3116 14671
rect 3695 15659 3729 15693
rect 3821 15659 3855 15693
rect 3695 15513 3729 15547
rect 3821 15513 3855 15547
rect 6211 15927 6245 15961
rect 6337 15927 6371 15961
rect 6211 15784 6245 15818
rect 6337 15784 6371 15818
rect 6211 15641 6245 15675
rect 6337 15641 6371 15675
rect 6211 15498 6245 15532
rect 6337 15498 6371 15532
rect 3695 15367 3729 15401
rect 3821 15367 3855 15401
rect 6211 15355 6245 15389
rect 6337 15355 6371 15389
rect 3695 15221 3729 15255
rect 3821 15221 3855 15255
rect 3695 15075 3729 15109
rect 3821 15075 3855 15109
rect 3695 14929 3729 14963
rect 3821 14929 3855 14963
rect 3695 14783 3729 14817
rect 3821 14783 3855 14817
rect 6211 15212 6245 15246
rect 6337 15212 6371 15246
rect 6211 15069 6245 15103
rect 6337 15069 6371 15103
rect 6211 14925 6245 14959
rect 6337 14925 6371 14959
rect 6211 14781 6245 14815
rect 6337 14781 6371 14815
rect 3695 14637 3729 14671
rect 3821 14637 3855 14671
rect 6211 14637 6245 14671
rect 6337 14637 6371 14671
rect 6476 16975 6510 17009
rect 6476 16907 6510 16941
rect 6476 16839 6510 16873
rect 6476 16771 6510 16805
rect 6476 16703 6510 16737
rect 6476 16635 6510 16669
rect 6476 16567 6510 16601
rect 6476 16499 6510 16533
rect 6476 16431 6510 16465
rect 6476 16363 6510 16397
rect 6476 16295 6510 16329
rect 6476 16227 6510 16261
rect 6476 16159 6510 16193
rect 6476 16091 6510 16125
rect 6476 16023 6510 16057
rect 6476 15955 6510 15989
rect 6476 15887 6510 15921
rect 6476 15819 6510 15853
rect 6476 15751 6510 15785
rect 6476 15683 6510 15717
rect 6476 15615 6510 15649
rect 6476 15547 6510 15581
rect 6476 15479 6510 15513
rect 6476 15411 6510 15445
rect 6476 15343 6510 15377
rect 6476 15275 6510 15309
rect 6476 15207 6510 15241
rect 6476 15139 6510 15173
rect 6476 15071 6510 15105
rect 6476 15003 6510 15037
rect 6476 14935 6510 14969
rect 6476 14867 6510 14901
rect 6476 14799 6510 14833
rect 6476 14731 6510 14765
rect 6476 14663 6510 14697
rect 3212 14569 3246 14603
rect 3280 14569 3314 14603
rect 3348 14569 3382 14603
rect 3416 14569 3450 14603
rect 3484 14569 3518 14603
rect 3552 14569 3586 14603
rect 3620 14569 3654 14603
rect 3688 14569 3722 14603
rect 3756 14569 3790 14603
rect 3824 14569 3858 14603
rect 3892 14569 3926 14603
rect 3960 14569 3994 14603
rect 4028 14569 4062 14603
rect 4096 14569 4130 14603
rect 4164 14569 4198 14603
rect 4232 14569 4266 14603
rect 4300 14569 4334 14603
rect 4368 14569 4402 14603
rect 4436 14569 4470 14603
rect 4504 14569 4538 14603
rect 4572 14569 4606 14603
rect 4640 14569 4674 14603
rect 4708 14569 4742 14603
rect 4776 14569 4810 14603
rect 4844 14569 4878 14603
rect 4912 14569 4946 14603
rect 4980 14569 5014 14603
rect 5048 14569 5082 14603
rect 5116 14569 5150 14603
rect 5184 14569 5218 14603
rect 5252 14569 5286 14603
rect 5320 14569 5354 14603
rect 5388 14569 5422 14603
rect 5456 14569 5490 14603
rect 5524 14569 5558 14603
rect 5592 14569 5626 14603
rect 5660 14569 5694 14603
rect 5728 14569 5762 14603
rect 5796 14569 5830 14603
rect 5864 14569 5898 14603
rect 5932 14569 5966 14603
rect 6000 14569 6034 14603
rect 6068 14569 6102 14603
rect 6136 14569 6170 14603
rect 6204 14569 6238 14603
rect 6272 14569 6306 14603
rect 6340 14569 6374 14603
rect 6408 14569 6442 14603
<< mvnsubdiffcont >>
rect 2918 39840 2952 39874
rect 2986 39840 3020 39874
rect 3054 39840 3088 39874
rect 3122 39840 3156 39874
rect 3190 39840 3224 39874
rect 3258 39840 3292 39874
rect 3326 39840 3360 39874
rect 3394 39840 3428 39874
rect 3462 39840 3496 39874
rect 3530 39840 3564 39874
rect 3598 39840 3632 39874
rect 3666 39840 3700 39874
rect 3734 39840 3768 39874
rect 3802 39840 3836 39874
rect 3870 39840 3904 39874
rect 3938 39840 3972 39874
rect 4006 39840 4040 39874
rect 4074 39840 4108 39874
rect 4142 39840 4176 39874
rect 4210 39840 4244 39874
rect 4278 39840 4312 39874
rect 4346 39840 4380 39874
rect 4414 39840 4448 39874
rect 4482 39840 4516 39874
rect 4550 39840 4584 39874
rect 4618 39840 4652 39874
rect 4686 39840 4720 39874
rect 4754 39840 4788 39874
rect 4822 39840 4856 39874
rect 4890 39840 4924 39874
rect 4958 39840 4992 39874
rect 5026 39840 5060 39874
rect 5094 39840 5128 39874
rect 5162 39840 5196 39874
rect 5230 39840 5264 39874
rect 5298 39840 5332 39874
rect 5366 39840 5400 39874
rect 5434 39840 5468 39874
rect 5502 39840 5536 39874
rect 5570 39840 5604 39874
rect 5638 39840 5672 39874
rect 5706 39840 5740 39874
rect 5774 39840 5808 39874
rect 5842 39840 5876 39874
rect 5910 39840 5944 39874
rect 5978 39840 6012 39874
rect 6046 39840 6080 39874
rect 6114 39840 6148 39874
rect 6182 39840 6216 39874
rect 6250 39840 6284 39874
rect 6318 39840 6352 39874
rect 6386 39840 6420 39874
rect 6454 39840 6488 39874
rect 6522 39840 6556 39874
rect 6590 39840 6624 39874
rect 6658 39840 6692 39874
rect 6726 39840 6760 39874
rect 6794 39840 6828 39874
rect 6862 39840 6896 39874
rect 6930 39840 6964 39874
rect 6998 39840 7032 39874
rect 7066 39840 7100 39874
rect 7134 39840 7168 39874
rect 7202 39840 7236 39874
rect 7270 39840 7304 39874
rect 7338 39840 7372 39874
rect 7406 39840 7440 39874
rect 7474 39840 7508 39874
rect 7542 39840 7576 39874
rect 7610 39840 7644 39874
rect 7678 39840 7712 39874
rect 2822 39772 2856 39806
rect 2822 39704 2856 39738
rect 2822 39636 2856 39670
rect 7746 39768 7780 39802
rect 7746 39700 7780 39734
rect 7746 39632 7780 39666
rect 2822 39568 2856 39602
rect 2822 39500 2856 39534
rect 2822 39432 2856 39466
rect 2822 39364 2856 39398
rect 2822 39296 2856 39330
rect 2822 39228 2856 39262
rect 2822 39160 2856 39194
rect 2822 39092 2856 39126
rect 2822 39024 2856 39058
rect 2822 38956 2856 38990
rect 2822 38888 2856 38922
rect 2822 38820 2856 38854
rect 2822 38752 2856 38786
rect 2822 38684 2856 38718
rect 2822 38616 2856 38650
rect 2822 38548 2856 38582
rect 2822 38480 2856 38514
rect 2822 38412 2856 38446
rect 2822 38344 2856 38378
rect 2822 38276 2856 38310
rect 2822 38208 2856 38242
rect 2822 38140 2856 38174
rect 2822 38072 2856 38106
rect 2822 38004 2856 38038
rect 2822 37936 2856 37970
rect 2822 37868 2856 37902
rect 2822 37800 2856 37834
rect 2822 37732 2856 37766
rect 2822 37664 2856 37698
rect 2822 37596 2856 37630
rect 2822 37528 2856 37562
rect 2822 37460 2856 37494
rect 2822 37392 2856 37426
rect 2822 37324 2856 37358
rect 2822 37256 2856 37290
rect 2822 37188 2856 37222
rect 2822 37120 2856 37154
rect 2822 37052 2856 37086
rect 2822 36984 2856 37018
rect 2822 36916 2856 36950
rect 2822 36848 2856 36882
rect 2822 36780 2856 36814
rect 2822 36712 2856 36746
rect 2822 36644 2856 36678
rect 2822 36576 2856 36610
rect 2822 36508 2856 36542
rect 2822 36440 2856 36474
rect 2822 36372 2856 36406
rect 2822 36304 2856 36338
rect 2822 36236 2856 36270
rect 2822 36168 2856 36202
rect 2822 36100 2856 36134
rect 2822 36032 2856 36066
rect 2822 35964 2856 35998
rect 2822 35896 2856 35930
rect 2822 35828 2856 35862
rect 2822 35760 2856 35794
rect 2822 35692 2856 35726
rect 2822 35624 2856 35658
rect 2822 35556 2856 35590
rect 2822 35488 2856 35522
rect 2822 35420 2856 35454
rect 2822 35352 2856 35386
rect 2822 35284 2856 35318
rect 2822 35216 2856 35250
rect 2822 35148 2856 35182
rect 2822 35080 2856 35114
rect 2822 35012 2856 35046
rect 2822 34944 2856 34978
rect 2822 34876 2856 34910
rect 2822 34808 2856 34842
rect 2822 34740 2856 34774
rect 2822 34672 2856 34706
rect 2822 34604 2856 34638
rect 2822 34536 2856 34570
rect 2822 34468 2856 34502
rect 2822 34400 2856 34434
rect 2822 34332 2856 34366
rect 2822 34264 2856 34298
rect 2822 34196 2856 34230
rect 2822 34128 2856 34162
rect 2822 34060 2856 34094
rect 2822 33992 2856 34026
rect 2822 33924 2856 33958
rect 2822 33856 2856 33890
rect 2822 33788 2856 33822
rect 2822 33720 2856 33754
rect 2822 33652 2856 33686
rect 2822 33584 2856 33618
rect 2822 33516 2856 33550
rect 2822 33448 2856 33482
rect 2822 33380 2856 33414
rect 2822 33312 2856 33346
rect 2822 33244 2856 33278
rect 2822 33176 2856 33210
rect 2822 33108 2856 33142
rect 2822 33040 2856 33074
rect 2822 32972 2856 33006
rect 2822 32904 2856 32938
rect 2822 32836 2856 32870
rect 2822 32768 2856 32802
rect 2822 32700 2856 32734
rect 2822 32632 2856 32666
rect 2822 32564 2856 32598
rect 2822 32496 2856 32530
rect 2822 32428 2856 32462
rect 2822 32360 2856 32394
rect 2822 32292 2856 32326
rect 2822 32224 2856 32258
rect 2822 32156 2856 32190
rect 2822 32088 2856 32122
rect 2822 32020 2856 32054
rect 2822 31952 2856 31986
rect 2822 31884 2856 31918
rect 2822 31816 2856 31850
rect 2822 31748 2856 31782
rect 2822 31680 2856 31714
rect 2822 31612 2856 31646
rect 2822 31544 2856 31578
rect 2822 31476 2856 31510
rect 2822 31408 2856 31442
rect 2822 31340 2856 31374
rect 2822 31272 2856 31306
rect 2822 31204 2856 31238
rect 2822 31136 2856 31170
rect 2822 31068 2856 31102
rect 2822 31000 2856 31034
rect 2822 30932 2856 30966
rect 2822 30864 2856 30898
rect 2822 30796 2856 30830
rect 2822 30728 2856 30762
rect 2822 30660 2856 30694
rect 2822 30592 2856 30626
rect 2822 30524 2856 30558
rect 2822 30456 2856 30490
rect 2822 30388 2856 30422
rect 2822 30320 2856 30354
rect 2822 30252 2856 30286
rect 2822 30184 2856 30218
rect 2822 30116 2856 30150
rect 2822 30048 2856 30082
rect 2822 29980 2856 30014
rect 2822 29912 2856 29946
rect 2822 29844 2856 29878
rect 2822 29776 2856 29810
rect 2822 29708 2856 29742
rect 2822 29640 2856 29674
rect 2822 29572 2856 29606
rect 2822 29504 2856 29538
rect 2822 29436 2856 29470
rect 2822 29368 2856 29402
rect 2822 29300 2856 29334
rect 2822 29232 2856 29266
rect 2822 29164 2856 29198
rect 2822 29096 2856 29130
rect 2822 29028 2856 29062
rect 2822 28960 2856 28994
rect 2822 28892 2856 28926
rect 2822 28824 2856 28858
rect 2822 28756 2856 28790
rect 2822 28688 2856 28722
rect 2822 28620 2856 28654
rect 2822 28552 2856 28586
rect 2822 28484 2856 28518
rect 2822 28416 2856 28450
rect 7746 39564 7780 39598
rect 7746 39496 7780 39530
rect 7746 39428 7780 39462
rect 7746 39360 7780 39394
rect 7746 39292 7780 39326
rect 7746 39224 7780 39258
rect 7746 39156 7780 39190
rect 7746 39088 7780 39122
rect 7746 39020 7780 39054
rect 7746 38952 7780 38986
rect 7746 38884 7780 38918
rect 7746 38816 7780 38850
rect 7746 38748 7780 38782
rect 7746 38680 7780 38714
rect 7746 38612 7780 38646
rect 7746 38544 7780 38578
rect 7746 38476 7780 38510
rect 7746 38408 7780 38442
rect 7746 38340 7780 38374
rect 7746 38272 7780 38306
rect 7746 38204 7780 38238
rect 7746 38136 7780 38170
rect 7746 38068 7780 38102
rect 7746 38000 7780 38034
rect 7746 37932 7780 37966
rect 7746 37864 7780 37898
rect 7746 37796 7780 37830
rect 7746 37728 7780 37762
rect 7746 37660 7780 37694
rect 7746 37592 7780 37626
rect 7746 37524 7780 37558
rect 7746 37456 7780 37490
rect 7746 37388 7780 37422
rect 7746 37320 7780 37354
rect 7746 37252 7780 37286
rect 7746 37184 7780 37218
rect 7746 37116 7780 37150
rect 7746 37048 7780 37082
rect 7746 36980 7780 37014
rect 7746 36912 7780 36946
rect 7746 36844 7780 36878
rect 7746 36776 7780 36810
rect 7746 36708 7780 36742
rect 7746 36640 7780 36674
rect 7746 36572 7780 36606
rect 7746 36504 7780 36538
rect 7746 36436 7780 36470
rect 7746 36368 7780 36402
rect 7746 36300 7780 36334
rect 7746 36232 7780 36266
rect 7746 36164 7780 36198
rect 7746 36096 7780 36130
rect 7746 36028 7780 36062
rect 7746 35960 7780 35994
rect 7746 35892 7780 35926
rect 7746 35824 7780 35858
rect 7746 35756 7780 35790
rect 7746 35688 7780 35722
rect 7746 35620 7780 35654
rect 7746 35552 7780 35586
rect 7746 35484 7780 35518
rect 7746 35416 7780 35450
rect 7746 35348 7780 35382
rect 7746 35280 7780 35314
rect 7746 35212 7780 35246
rect 7746 35144 7780 35178
rect 7746 35076 7780 35110
rect 7746 35008 7780 35042
rect 7746 34940 7780 34974
rect 7746 34872 7780 34906
rect 7746 34804 7780 34838
rect 7746 34736 7780 34770
rect 7746 34668 7780 34702
rect 7746 34600 7780 34634
rect 7746 34532 7780 34566
rect 7746 34464 7780 34498
rect 7746 34396 7780 34430
rect 7746 34328 7780 34362
rect 7746 34260 7780 34294
rect 7746 34192 7780 34226
rect 7746 34124 7780 34158
rect 7746 34056 7780 34090
rect 7746 33988 7780 34022
rect 7746 33920 7780 33954
rect 7746 33852 7780 33886
rect 7746 33784 7780 33818
rect 7746 33716 7780 33750
rect 7746 33648 7780 33682
rect 7746 33580 7780 33614
rect 7746 33512 7780 33546
rect 7746 33444 7780 33478
rect 7746 33376 7780 33410
rect 7746 33308 7780 33342
rect 7746 33240 7780 33274
rect 7746 33172 7780 33206
rect 7746 33104 7780 33138
rect 7746 33036 7780 33070
rect 7746 32968 7780 33002
rect 7746 32900 7780 32934
rect 7746 32832 7780 32866
rect 7746 32764 7780 32798
rect 7746 32696 7780 32730
rect 7746 32628 7780 32662
rect 7746 32560 7780 32594
rect 7746 32492 7780 32526
rect 7746 32424 7780 32458
rect 7746 32356 7780 32390
rect 7746 32288 7780 32322
rect 7746 32220 7780 32254
rect 7746 32152 7780 32186
rect 7746 32084 7780 32118
rect 7746 32016 7780 32050
rect 7746 31948 7780 31982
rect 7746 31880 7780 31914
rect 7746 31812 7780 31846
rect 7746 31744 7780 31778
rect 7746 31676 7780 31710
rect 7746 31608 7780 31642
rect 7746 31540 7780 31574
rect 7746 31472 7780 31506
rect 7746 31404 7780 31438
rect 7746 31336 7780 31370
rect 7746 31268 7780 31302
rect 7746 31200 7780 31234
rect 7746 31132 7780 31166
rect 7746 31064 7780 31098
rect 7746 30996 7780 31030
rect 7746 30928 7780 30962
rect 7746 30860 7780 30894
rect 7746 30792 7780 30826
rect 7746 30724 7780 30758
rect 7746 30656 7780 30690
rect 7746 30588 7780 30622
rect 7746 30520 7780 30554
rect 7746 30452 7780 30486
rect 7746 30384 7780 30418
rect 7746 30316 7780 30350
rect 7746 30248 7780 30282
rect 7746 30180 7780 30214
rect 7746 30112 7780 30146
rect 7746 30044 7780 30078
rect 7746 29976 7780 30010
rect 7746 29908 7780 29942
rect 7746 29840 7780 29874
rect 7746 29772 7780 29806
rect 7746 29704 7780 29738
rect 7746 29636 7780 29670
rect 7746 29568 7780 29602
rect 7746 29500 7780 29534
rect 7746 29432 7780 29466
rect 7746 29364 7780 29398
rect 7746 29296 7780 29330
rect 7746 29228 7780 29262
rect 7746 29160 7780 29194
rect 7746 29092 7780 29126
rect 7746 29024 7780 29058
rect 7746 28956 7780 28990
rect 7746 28888 7780 28922
rect 7746 28820 7780 28854
rect 7746 28752 7780 28786
rect 7746 28684 7780 28718
rect 7746 28616 7780 28650
rect 7746 28548 7780 28582
rect 7746 28480 7780 28514
rect 7746 28412 7780 28446
rect 2822 28348 2856 28382
rect 2822 28232 2856 28266
rect 7746 28344 7780 28378
rect 7746 28276 7780 28310
rect 7746 28208 7780 28242
rect 2890 28140 2924 28174
rect 2958 28140 2992 28174
rect 3026 28140 3060 28174
rect 3094 28140 3128 28174
rect 3162 28140 3196 28174
rect 3230 28140 3264 28174
rect 3298 28140 3332 28174
rect 3366 28140 3400 28174
rect 3434 28140 3468 28174
rect 3502 28140 3536 28174
rect 3570 28140 3604 28174
rect 3638 28140 3672 28174
rect 3706 28140 3740 28174
rect 3774 28140 3808 28174
rect 3842 28140 3876 28174
rect 3910 28140 3944 28174
rect 3978 28140 4012 28174
rect 4046 28140 4080 28174
rect 4114 28140 4148 28174
rect 4182 28140 4216 28174
rect 4250 28140 4284 28174
rect 4318 28140 4352 28174
rect 4386 28140 4420 28174
rect 4454 28140 4488 28174
rect 4522 28140 4556 28174
rect 4590 28140 4624 28174
rect 4658 28140 4692 28174
rect 4726 28140 4760 28174
rect 4794 28140 4828 28174
rect 4862 28140 4896 28174
rect 4930 28140 4964 28174
rect 4998 28140 5032 28174
rect 5066 28140 5100 28174
rect 5134 28140 5168 28174
rect 5202 28140 5236 28174
rect 5270 28140 5304 28174
rect 5338 28140 5372 28174
rect 5406 28140 5440 28174
rect 5474 28140 5508 28174
rect 5542 28140 5576 28174
rect 5610 28140 5644 28174
rect 5678 28140 5712 28174
rect 5746 28140 5780 28174
rect 5814 28140 5848 28174
rect 5882 28140 5916 28174
rect 5950 28140 5984 28174
rect 6018 28140 6052 28174
rect 6086 28140 6120 28174
rect 6154 28140 6188 28174
rect 6222 28140 6256 28174
rect 6290 28140 6324 28174
rect 6358 28140 6392 28174
rect 6426 28140 6460 28174
rect 6494 28140 6528 28174
rect 6562 28140 6596 28174
rect 6630 28140 6664 28174
rect 6698 28140 6732 28174
rect 6766 28140 6800 28174
rect 6834 28140 6868 28174
rect 6902 28140 6936 28174
rect 6970 28140 7004 28174
rect 7038 28140 7072 28174
rect 7106 28140 7140 28174
rect 7174 28140 7208 28174
rect 7242 28140 7276 28174
rect 7310 28140 7344 28174
rect 7378 28140 7412 28174
rect 7446 28140 7480 28174
rect 7514 28140 7548 28174
rect 7582 28140 7616 28174
rect 7650 28140 7684 28174
rect 4008 26048 4042 26082
rect 4008 25980 4042 26014
rect 4008 25912 4042 25946
rect 4008 25844 4042 25878
rect 4008 25776 4042 25810
rect 4008 25708 4042 25742
rect 4008 25640 4042 25674
rect 4008 25572 4042 25606
rect 4008 25504 4042 25538
rect 4008 25436 4042 25470
rect 4008 25368 4042 25402
rect 4008 25300 4042 25334
rect 4008 25232 4042 25266
rect 4008 25164 4042 25198
rect 4008 25096 4042 25130
rect 4008 25028 4042 25062
rect 4008 24960 4042 24994
rect 4008 24892 4042 24926
rect 4008 24824 4042 24858
rect 4008 24756 4042 24790
rect 5946 26048 5980 26082
rect 5946 25980 5980 26014
rect 5946 25912 5980 25946
rect 5946 25844 5980 25878
rect 5946 25776 5980 25810
rect 5946 25708 5980 25742
rect 5946 25640 5980 25674
rect 5946 25572 5980 25606
rect 5946 25504 5980 25538
rect 5946 25436 5980 25470
rect 5946 25368 5980 25402
rect 5946 25300 5980 25334
rect 5946 25232 5980 25266
rect 5946 25164 5980 25198
rect 5946 25096 5980 25130
rect 5946 25028 5980 25062
rect 5946 24960 5980 24994
rect 5946 24892 5980 24926
rect 5946 24824 5980 24858
rect 5946 24756 5980 24790
rect 4528 24150 4562 24184
rect 4596 24150 4630 24184
rect 4664 24150 4698 24184
rect 4732 24150 4766 24184
rect 4800 24150 4834 24184
rect 4868 24150 4902 24184
rect 4936 24150 4970 24184
rect 5004 24150 5038 24184
rect 5072 24150 5106 24184
rect 5140 24150 5174 24184
rect 5208 24150 5242 24184
rect 5276 24150 5310 24184
rect 5344 24150 5378 24184
rect 5412 24150 5446 24184
rect 5480 24150 5514 24184
rect 5548 24150 5582 24184
rect 5616 24150 5650 24184
rect 5684 24150 5718 24184
rect 5752 24150 5786 24184
rect 4460 24076 4494 24110
rect 5858 24082 5892 24116
rect 4460 23922 4494 23956
rect 4460 23854 4494 23888
rect 4460 23786 4494 23820
rect 5858 24014 5892 24048
rect 5858 23946 5892 23980
rect 5858 23878 5892 23912
rect 5858 23810 5892 23844
rect 4460 23718 4494 23752
rect 5858 23742 5892 23776
rect 4460 23650 4494 23684
rect 4460 23582 4494 23616
rect 4460 23514 4494 23548
rect 4460 23446 4494 23480
rect 4460 23378 4494 23412
rect 4460 23310 4494 23344
rect 4460 23242 4494 23276
rect 4460 23174 4494 23208
rect 4460 23106 4494 23140
rect 4460 23038 4494 23072
rect 4460 22970 4494 23004
rect 4460 22902 4494 22936
rect 4460 22834 4494 22868
rect 4460 22766 4494 22800
rect 4460 22698 4494 22732
rect 4460 22630 4494 22664
rect 4460 22562 4494 22596
rect 4460 22494 4494 22528
rect 4460 22426 4494 22460
rect 4460 22358 4494 22392
rect 4460 22290 4494 22324
rect 4460 22222 4494 22256
rect 4460 22154 4494 22188
rect 4460 22086 4494 22120
rect 4460 22018 4494 22052
rect 4460 21950 4494 21984
rect 4460 21882 4494 21916
rect 4460 21814 4494 21848
rect 4460 21746 4494 21780
rect 4460 21678 4494 21712
rect 4460 21610 4494 21644
rect 4460 21542 4494 21576
rect 4460 21474 4494 21508
rect 4460 21406 4494 21440
rect 4460 21338 4494 21372
rect 4460 21270 4494 21304
rect 4460 21202 4494 21236
rect 4460 21134 4494 21168
rect 4460 21066 4494 21100
rect 4460 20998 4494 21032
rect 4460 20930 4494 20964
rect 4460 20862 4494 20896
rect 4460 20794 4494 20828
rect 4460 20726 4494 20760
rect 4460 20658 4494 20692
rect 4460 20590 4494 20624
rect 4460 20522 4494 20556
rect 4460 20454 4494 20488
rect 4460 20386 4494 20420
rect 4460 20318 4494 20352
rect 4460 20250 4494 20284
rect 4460 20182 4494 20216
rect 4460 20114 4494 20148
rect 4460 20046 4494 20080
rect 4460 19978 4494 20012
rect 4460 19910 4494 19944
rect 4460 19842 4494 19876
rect 4460 19774 4494 19808
rect 4460 19706 4494 19740
rect 4460 19638 4494 19672
rect 4460 19570 4494 19604
rect 4460 19502 4494 19536
rect 5858 23674 5892 23708
rect 5858 23606 5892 23640
rect 5858 23538 5892 23572
rect 5858 23470 5892 23504
rect 5858 23402 5892 23436
rect 5858 23334 5892 23368
rect 5858 23266 5892 23300
rect 5858 23198 5892 23232
rect 5858 23130 5892 23164
rect 5858 23062 5892 23096
rect 5858 22994 5892 23028
rect 5858 22926 5892 22960
rect 5858 22858 5892 22892
rect 5858 22790 5892 22824
rect 5858 22722 5892 22756
rect 5858 22654 5892 22688
rect 5858 22586 5892 22620
rect 5858 22518 5892 22552
rect 5858 22450 5892 22484
rect 5858 22382 5892 22416
rect 5858 22314 5892 22348
rect 5858 22246 5892 22280
rect 5858 22178 5892 22212
rect 5858 22110 5892 22144
rect 5858 22042 5892 22076
rect 5858 21974 5892 22008
rect 5858 21906 5892 21940
rect 5858 21838 5892 21872
rect 5858 21770 5892 21804
rect 5858 21702 5892 21736
rect 5858 21634 5892 21668
rect 5858 21566 5892 21600
rect 5858 21498 5892 21532
rect 7420 21485 7454 21519
rect 7488 21485 7522 21519
rect 7556 21485 7590 21519
rect 7624 21485 7658 21519
rect 5858 21430 5892 21464
rect 5858 21362 5892 21396
rect 5858 21294 5892 21328
rect 5858 21226 5892 21260
rect 5858 21158 5892 21192
rect 5858 21090 5892 21124
rect 5858 21022 5892 21056
rect 5858 20954 5892 20988
rect 5858 20886 5892 20920
rect 5858 20818 5892 20852
rect 5858 20750 5892 20784
rect 5858 20682 5892 20716
rect 5858 20614 5892 20648
rect 5858 20546 5892 20580
rect 5858 20478 5892 20512
rect 5858 20410 5892 20444
rect 5858 20342 5892 20376
rect 5858 20274 5892 20308
rect 5858 20206 5892 20240
rect 5858 20138 5892 20172
rect 5858 20070 5892 20104
rect 5858 20002 5892 20036
rect 5858 19934 5892 19968
rect 5858 19866 5892 19900
rect 5858 19798 5892 19832
rect 5858 19730 5892 19764
rect 5858 19662 5892 19696
rect 4460 19434 4494 19468
rect 5858 19594 5892 19628
rect 5858 19526 5892 19560
rect 5858 19458 5892 19492
rect 4460 19366 4494 19400
rect 4460 19298 4494 19332
rect 4460 19230 4494 19264
rect 4460 19162 4494 19196
rect 4460 19094 4494 19128
rect 5858 19390 5892 19424
rect 5858 19322 5892 19356
rect 5858 19254 5892 19288
rect 5858 19186 5892 19220
rect 5858 19118 5892 19152
rect 4460 19026 4494 19060
rect 5858 19050 5892 19084
rect 4460 18958 4494 18992
rect 4460 18890 4494 18924
rect 4460 18822 4494 18856
rect 4460 18754 4494 18788
rect 5858 18982 5892 19016
rect 5858 18914 5892 18948
rect 5858 18846 5892 18880
rect 4460 18686 4494 18720
rect 4460 18618 4494 18652
rect 4460 18550 4494 18584
rect 5858 18778 5892 18812
rect 5858 18710 5892 18744
rect 5858 18642 5892 18676
rect 5858 18574 5892 18608
rect 4566 18482 4600 18516
rect 4634 18482 4668 18516
rect 4702 18482 4736 18516
rect 4770 18482 4804 18516
rect 4838 18482 4872 18516
rect 4906 18482 4940 18516
rect 4974 18482 5008 18516
rect 5042 18482 5076 18516
rect 5110 18482 5144 18516
rect 5178 18482 5212 18516
rect 5246 18482 5280 18516
rect 5314 18482 5348 18516
rect 5382 18482 5416 18516
rect 5450 18482 5484 18516
rect 5518 18482 5552 18516
rect 5586 18482 5620 18516
rect 5654 18482 5688 18516
rect 5722 18482 5756 18516
rect 5790 18482 5824 18516
rect 2890 18255 2924 18289
rect 2958 18255 2992 18289
rect 3026 18255 3060 18289
rect 3094 18255 3128 18289
rect 3162 18255 3196 18289
rect 3230 18255 3264 18289
rect 3298 18255 3332 18289
rect 3366 18255 3400 18289
rect 3434 18255 3468 18289
rect 3502 18255 3536 18289
rect 3570 18255 3604 18289
rect 3638 18255 3672 18289
rect 3706 18255 3740 18289
rect 3774 18255 3808 18289
rect 3842 18255 3876 18289
rect 3910 18255 3944 18289
rect 3978 18255 4012 18289
rect 4046 18255 4080 18289
rect 4114 18255 4148 18289
rect 4182 18255 4216 18289
rect 4250 18255 4284 18289
rect 4318 18255 4352 18289
rect 4386 18255 4420 18289
rect 4454 18255 4488 18289
rect 4522 18255 4556 18289
rect 4590 18255 4624 18289
rect 4658 18255 4692 18289
rect 4726 18255 4760 18289
rect 4794 18255 4828 18289
rect 4862 18255 4896 18289
rect 4930 18255 4964 18289
rect 4998 18255 5032 18289
rect 5066 18255 5100 18289
rect 5134 18255 5168 18289
rect 5202 18255 5236 18289
rect 5270 18255 5304 18289
rect 5338 18255 5372 18289
rect 5406 18255 5440 18289
rect 5474 18255 5508 18289
rect 5542 18255 5576 18289
rect 5610 18255 5644 18289
rect 5678 18255 5712 18289
rect 5746 18255 5780 18289
rect 5814 18255 5848 18289
rect 5882 18255 5916 18289
rect 5950 18255 5984 18289
rect 6018 18255 6052 18289
rect 6086 18255 6120 18289
rect 6154 18255 6188 18289
rect 6222 18255 6256 18289
rect 6290 18255 6324 18289
rect 6358 18255 6392 18289
rect 6426 18255 6460 18289
rect 6494 18255 6528 18289
rect 6562 18255 6596 18289
rect 6630 18255 6664 18289
rect 2822 18163 2856 18197
rect 2822 18049 2856 18083
rect 6750 18187 6784 18221
rect 6750 18119 6784 18153
rect 6750 18051 6784 18085
rect 2822 17981 2856 18015
rect 2822 17913 2856 17947
rect 2822 17845 2856 17879
rect 2822 17777 2856 17811
rect 2822 17709 2856 17743
rect 2822 17641 2856 17675
rect 2822 17573 2856 17607
rect 2822 17505 2856 17539
rect 2822 17437 2856 17471
rect 2822 17369 2856 17403
rect 2822 17301 2856 17335
rect 2822 17233 2856 17267
rect 2822 17165 2856 17199
rect 2822 17097 2856 17131
rect 2822 17029 2856 17063
rect 2822 16961 2856 16995
rect 2822 16893 2856 16927
rect 2822 16825 2856 16859
rect 2822 16757 2856 16791
rect 2822 16689 2856 16723
rect 2822 16621 2856 16655
rect 2822 16553 2856 16587
rect 2822 16485 2856 16519
rect 2822 16417 2856 16451
rect 2822 16349 2856 16383
rect 2822 16281 2856 16315
rect 2822 16213 2856 16247
rect 2822 16145 2856 16179
rect 2822 16077 2856 16111
rect 2822 16009 2856 16043
rect 2822 15941 2856 15975
rect 2822 15873 2856 15907
rect 2822 15805 2856 15839
rect 2822 15737 2856 15771
rect 2822 15669 2856 15703
rect 2822 15601 2856 15635
rect 2822 15533 2856 15567
rect 2822 15465 2856 15499
rect 2822 15397 2856 15431
rect 2822 15329 2856 15363
rect 2822 15261 2856 15295
rect 2822 15193 2856 15227
rect 2822 15125 2856 15159
rect 2822 15057 2856 15091
rect 2822 14989 2856 15023
rect 2822 14921 2856 14955
rect 2822 14853 2856 14887
rect 2822 14785 2856 14819
rect 2822 14717 2856 14751
rect 2822 14649 2856 14683
rect 2822 14581 2856 14615
rect 6750 17983 6784 18017
rect 6750 17915 6784 17949
rect 6750 17847 6784 17881
rect 6750 17779 6784 17813
rect 6750 17711 6784 17745
rect 6750 17643 6784 17677
rect 6750 17575 6784 17609
rect 6750 17507 6784 17541
rect 6750 17439 6784 17473
rect 6750 17371 6784 17405
rect 6750 17303 6784 17337
rect 6750 17235 6784 17269
rect 6750 17167 6784 17201
rect 6750 17099 6784 17133
rect 6750 17031 6784 17065
rect 6750 16963 6784 16997
rect 6750 16895 6784 16929
rect 6750 16827 6784 16861
rect 6750 16759 6784 16793
rect 6750 16691 6784 16725
rect 6750 16623 6784 16657
rect 6750 16555 6784 16589
rect 6750 16487 6784 16521
rect 6750 16419 6784 16453
rect 6750 16351 6784 16385
rect 6750 16283 6784 16317
rect 6750 16215 6784 16249
rect 6750 16147 6784 16181
rect 6750 16079 6784 16113
rect 6750 16011 6784 16045
rect 6750 15943 6784 15977
rect 6750 15875 6784 15909
rect 6750 15807 6784 15841
rect 6750 15739 6784 15773
rect 6750 15671 6784 15705
rect 6750 15603 6784 15637
rect 6750 15535 6784 15569
rect 6750 15467 6784 15501
rect 6750 15399 6784 15433
rect 6750 15331 6784 15365
rect 6750 15263 6784 15297
rect 6750 15195 6784 15229
rect 6750 15127 6784 15161
rect 6750 15059 6784 15093
rect 6750 14991 6784 15025
rect 6750 14923 6784 14957
rect 6750 14855 6784 14889
rect 6750 14787 6784 14821
rect 6750 14719 6784 14753
rect 6750 14651 6784 14685
rect 6750 14583 6784 14617
rect 2822 14513 2856 14547
rect 2822 14445 2856 14479
rect 2822 14377 2856 14411
rect 6750 14515 6784 14549
rect 6750 14447 6784 14481
rect 6750 14379 6784 14413
rect 2942 14309 2976 14343
rect 3010 14309 3044 14343
rect 3078 14309 3112 14343
rect 3146 14309 3180 14343
rect 3214 14309 3248 14343
rect 3282 14309 3316 14343
rect 3350 14309 3384 14343
rect 3418 14309 3452 14343
rect 3486 14309 3520 14343
rect 3554 14309 3588 14343
rect 3622 14309 3656 14343
rect 3690 14309 3724 14343
rect 3758 14309 3792 14343
rect 3826 14309 3860 14343
rect 3894 14309 3928 14343
rect 3962 14309 3996 14343
rect 4030 14309 4064 14343
rect 4098 14309 4132 14343
rect 4166 14309 4200 14343
rect 4234 14309 4268 14343
rect 4302 14309 4336 14343
rect 4370 14309 4404 14343
rect 4438 14309 4472 14343
rect 4506 14309 4540 14343
rect 4574 14309 4608 14343
rect 4642 14309 4676 14343
rect 4710 14309 4744 14343
rect 4778 14309 4812 14343
rect 4846 14309 4880 14343
rect 4914 14309 4948 14343
rect 4982 14309 5016 14343
rect 5050 14309 5084 14343
rect 5118 14309 5152 14343
rect 5186 14309 5220 14343
rect 5254 14309 5288 14343
rect 5322 14309 5356 14343
rect 5390 14309 5424 14343
rect 5458 14309 5492 14343
rect 5526 14309 5560 14343
rect 5594 14309 5628 14343
rect 5662 14309 5696 14343
rect 5730 14309 5764 14343
rect 5798 14309 5832 14343
rect 5866 14309 5900 14343
rect 5934 14309 5968 14343
rect 6002 14309 6036 14343
rect 6070 14309 6104 14343
rect 6138 14309 6172 14343
rect 6206 14309 6240 14343
rect 6274 14309 6308 14343
rect 6342 14309 6376 14343
rect 6410 14309 6444 14343
rect 6478 14309 6512 14343
rect 6546 14309 6580 14343
rect 6614 14309 6648 14343
rect 6682 14309 6716 14343
<< poly >>
rect 3158 39431 3224 39447
rect 3158 39397 3174 39431
rect 3208 39397 3224 39431
rect 3158 39363 3224 39397
rect 3158 39329 3174 39363
rect 3208 39329 3224 39363
rect 3158 39295 3224 39329
rect 3158 39261 3174 39295
rect 3208 39261 3224 39295
rect 3158 39227 3224 39261
rect 3158 39193 3174 39227
rect 3208 39193 3224 39227
rect 3158 39159 3224 39193
rect 3158 39125 3174 39159
rect 3208 39125 3224 39159
rect 3158 39091 3224 39125
rect 3158 39057 3174 39091
rect 3208 39057 3224 39091
rect 3158 39023 3224 39057
rect 3158 38989 3174 39023
rect 3208 38989 3224 39023
rect 3158 38955 3224 38989
rect 3158 38921 3174 38955
rect 3208 38921 3224 38955
rect 3158 38887 3224 38921
rect 3158 38853 3174 38887
rect 3208 38853 3224 38887
rect 3158 38819 3224 38853
rect 3158 38785 3174 38819
rect 3208 38785 3224 38819
rect 3158 38751 3224 38785
rect 3158 38717 3174 38751
rect 3208 38717 3224 38751
rect 3158 38683 3224 38717
rect 3158 38649 3174 38683
rect 3208 38649 3224 38683
rect 3158 38615 3224 38649
rect 3158 38581 3174 38615
rect 3208 38581 3224 38615
rect 3158 38547 3224 38581
rect 3158 38513 3174 38547
rect 3208 38513 3224 38547
rect 3158 38479 3224 38513
rect 3158 38445 3174 38479
rect 3208 38445 3224 38479
rect 3158 38411 3224 38445
rect 3158 38377 3174 38411
rect 3208 38377 3224 38411
rect 3158 38343 3224 38377
rect 3158 38309 3174 38343
rect 3208 38309 3224 38343
rect 3158 38275 3224 38309
rect 3158 38241 3174 38275
rect 3208 38241 3224 38275
rect 3158 38207 3224 38241
rect 3158 38173 3174 38207
rect 3208 38173 3224 38207
rect 3158 38139 3224 38173
rect 3158 38105 3174 38139
rect 3208 38105 3224 38139
rect 3158 38071 3224 38105
rect 3158 38037 3174 38071
rect 3208 38037 3224 38071
rect 3158 38003 3224 38037
rect 3158 37969 3174 38003
rect 3208 37969 3224 38003
rect 3158 37935 3224 37969
rect 3158 37901 3174 37935
rect 3208 37901 3224 37935
rect 3158 37867 3224 37901
rect 3158 37833 3174 37867
rect 3208 37833 3224 37867
rect 3158 37799 3224 37833
rect 3158 37765 3174 37799
rect 3208 37765 3224 37799
rect 3158 37731 3224 37765
rect 3158 37697 3174 37731
rect 3208 37697 3224 37731
rect 3158 37663 3224 37697
rect 3158 37629 3174 37663
rect 3208 37629 3224 37663
rect 3158 37595 3224 37629
rect 3158 37561 3174 37595
rect 3208 37561 3224 37595
rect 3158 37527 3224 37561
rect 3158 37493 3174 37527
rect 3208 37493 3224 37527
rect 3158 37459 3224 37493
rect 3158 37425 3174 37459
rect 3208 37425 3224 37459
rect 3158 37391 3224 37425
rect 3158 37357 3174 37391
rect 3208 37357 3224 37391
rect 3158 37323 3224 37357
rect 3158 37289 3174 37323
rect 3208 37289 3224 37323
rect 3158 37255 3224 37289
rect 3158 37221 3174 37255
rect 3208 37221 3224 37255
rect 3158 37187 3224 37221
rect 3158 37153 3174 37187
rect 3208 37153 3224 37187
rect 3158 37119 3224 37153
rect 3158 37085 3174 37119
rect 3208 37085 3224 37119
rect 3158 37051 3224 37085
rect 3158 37017 3174 37051
rect 3208 37017 3224 37051
rect 3158 36983 3224 37017
rect 3158 36949 3174 36983
rect 3208 36949 3224 36983
rect 3158 36915 3224 36949
rect 3158 36881 3174 36915
rect 3208 36881 3224 36915
rect 3158 36847 3224 36881
rect 3158 36813 3174 36847
rect 3208 36813 3224 36847
rect 3158 36779 3224 36813
rect 3158 36745 3174 36779
rect 3208 36745 3224 36779
rect 3158 36711 3224 36745
rect 3158 36677 3174 36711
rect 3208 36677 3224 36711
rect 3158 36643 3224 36677
rect 3158 36609 3174 36643
rect 3208 36609 3224 36643
rect 3158 36575 3224 36609
rect 3158 36541 3174 36575
rect 3208 36541 3224 36575
rect 3158 36507 3224 36541
rect 3158 36473 3174 36507
rect 3208 36473 3224 36507
rect 3158 36439 3224 36473
rect 3158 36405 3174 36439
rect 3208 36405 3224 36439
rect 3158 36371 3224 36405
rect 3158 36337 3174 36371
rect 3208 36337 3224 36371
rect 3158 36303 3224 36337
rect 3158 36269 3174 36303
rect 3208 36269 3224 36303
rect 3158 36235 3224 36269
rect 3158 36201 3174 36235
rect 3208 36201 3224 36235
rect 3158 36167 3224 36201
rect 3158 36133 3174 36167
rect 3208 36133 3224 36167
rect 3158 36099 3224 36133
rect 3158 36065 3174 36099
rect 3208 36065 3224 36099
rect 3158 36031 3224 36065
rect 3158 35997 3174 36031
rect 3208 35997 3224 36031
rect 3158 35963 3224 35997
rect 3158 35929 3174 35963
rect 3208 35929 3224 35963
rect 3158 35895 3224 35929
rect 3158 35861 3174 35895
rect 3208 35861 3224 35895
rect 3158 35827 3224 35861
rect 3158 35793 3174 35827
rect 3208 35793 3224 35827
rect 3158 35759 3224 35793
rect 3158 35725 3174 35759
rect 3208 35725 3224 35759
rect 3158 35691 3224 35725
rect 3158 35657 3174 35691
rect 3208 35657 3224 35691
rect 3158 35623 3224 35657
rect 3158 35589 3174 35623
rect 3208 35589 3224 35623
rect 3158 35555 3224 35589
rect 3158 35521 3174 35555
rect 3208 35521 3224 35555
rect 3158 35487 3224 35521
rect 3158 35453 3174 35487
rect 3208 35453 3224 35487
rect 3158 35419 3224 35453
rect 3158 35385 3174 35419
rect 3208 35385 3224 35419
rect 3158 35351 3224 35385
rect 3158 35317 3174 35351
rect 3208 35317 3224 35351
rect 3158 35283 3224 35317
rect 3158 35249 3174 35283
rect 3208 35249 3224 35283
rect 3158 35215 3224 35249
rect 3158 35181 3174 35215
rect 3208 35181 3224 35215
rect 3158 35147 3224 35181
rect 3158 35113 3174 35147
rect 3208 35113 3224 35147
rect 3158 35079 3224 35113
rect 3158 35045 3174 35079
rect 3208 35045 3224 35079
rect 3158 35011 3224 35045
rect 3158 34977 3174 35011
rect 3208 34977 3224 35011
rect 3158 34943 3224 34977
rect 3158 34909 3174 34943
rect 3208 34909 3224 34943
rect 3158 34875 3224 34909
rect 3158 34841 3174 34875
rect 3208 34841 3224 34875
rect 3158 34807 3224 34841
rect 3158 34773 3174 34807
rect 3208 34773 3224 34807
rect 3158 34739 3224 34773
rect 3158 34705 3174 34739
rect 3208 34705 3224 34739
rect 3158 34671 3224 34705
rect 3158 34637 3174 34671
rect 3208 34637 3224 34671
rect 3158 34603 3224 34637
rect 3158 34569 3174 34603
rect 3208 34569 3224 34603
rect 3158 34535 3224 34569
rect 3158 34501 3174 34535
rect 3208 34501 3224 34535
rect 3158 34467 3224 34501
rect 3158 34433 3174 34467
rect 3208 34433 3224 34467
rect 3158 34399 3224 34433
rect 3158 34365 3174 34399
rect 3208 34365 3224 34399
rect 3158 34331 3224 34365
rect 3158 34297 3174 34331
rect 3208 34297 3224 34331
rect 3158 34263 3224 34297
rect 3158 34229 3174 34263
rect 3208 34229 3224 34263
rect 3158 34195 3224 34229
rect 3158 34161 3174 34195
rect 3208 34161 3224 34195
rect 3158 34127 3224 34161
rect 3158 34093 3174 34127
rect 3208 34093 3224 34127
rect 3158 34059 3224 34093
rect 3158 34025 3174 34059
rect 3208 34025 3224 34059
rect 3158 33991 3224 34025
rect 3158 33957 3174 33991
rect 3208 33957 3224 33991
rect 3158 33923 3224 33957
rect 3158 33889 3174 33923
rect 3208 33889 3224 33923
rect 3158 33855 3224 33889
rect 3158 33821 3174 33855
rect 3208 33821 3224 33855
rect 3158 33787 3224 33821
rect 3158 33753 3174 33787
rect 3208 33753 3224 33787
rect 3158 33719 3224 33753
rect 3158 33685 3174 33719
rect 3208 33685 3224 33719
rect 3158 33651 3224 33685
rect 3158 33617 3174 33651
rect 3208 33617 3224 33651
rect 3158 33583 3224 33617
rect 3158 33549 3174 33583
rect 3208 33549 3224 33583
rect 3158 33515 3224 33549
rect 3158 33481 3174 33515
rect 3208 33481 3224 33515
rect 3158 33447 3224 33481
rect 3158 33413 3174 33447
rect 3208 33413 3224 33447
rect 3158 33379 3224 33413
rect 3158 33345 3174 33379
rect 3208 33345 3224 33379
rect 3158 33311 3224 33345
rect 3158 33277 3174 33311
rect 3208 33277 3224 33311
rect 3158 33243 3224 33277
rect 3158 33209 3174 33243
rect 3208 33209 3224 33243
rect 3158 33175 3224 33209
rect 3158 33141 3174 33175
rect 3208 33141 3224 33175
rect 3158 33107 3224 33141
rect 3158 33073 3174 33107
rect 3208 33073 3224 33107
rect 3158 33039 3224 33073
rect 3158 33005 3174 33039
rect 3208 33005 3224 33039
rect 3158 32971 3224 33005
rect 3158 32937 3174 32971
rect 3208 32937 3224 32971
rect 3158 32903 3224 32937
rect 3158 32869 3174 32903
rect 3208 32869 3224 32903
rect 3158 32835 3224 32869
rect 3158 32801 3174 32835
rect 3208 32801 3224 32835
rect 3158 32767 3224 32801
rect 3158 32733 3174 32767
rect 3208 32733 3224 32767
rect 3158 32699 3224 32733
rect 3158 32665 3174 32699
rect 3208 32665 3224 32699
rect 3158 32631 3224 32665
rect 3158 32597 3174 32631
rect 3208 32597 3224 32631
rect 3158 32563 3224 32597
rect 3158 32529 3174 32563
rect 3208 32529 3224 32563
rect 3158 32495 3224 32529
rect 3158 32461 3174 32495
rect 3208 32461 3224 32495
rect 3158 32427 3224 32461
rect 3158 32393 3174 32427
rect 3208 32393 3224 32427
rect 3158 32359 3224 32393
rect 3158 32325 3174 32359
rect 3208 32325 3224 32359
rect 3158 32291 3224 32325
rect 3158 32257 3174 32291
rect 3208 32257 3224 32291
rect 3158 32223 3224 32257
rect 3158 32189 3174 32223
rect 3208 32189 3224 32223
rect 3158 32155 3224 32189
rect 3158 32121 3174 32155
rect 3208 32121 3224 32155
rect 3158 32087 3224 32121
rect 3158 32053 3174 32087
rect 3208 32053 3224 32087
rect 3158 32019 3224 32053
rect 3158 31985 3174 32019
rect 3208 31985 3224 32019
rect 3158 31951 3224 31985
rect 3158 31917 3174 31951
rect 3208 31917 3224 31951
rect 3158 31882 3224 31917
rect 3158 31848 3174 31882
rect 3208 31848 3224 31882
rect 3158 31813 3224 31848
rect 3158 31779 3174 31813
rect 3208 31779 3224 31813
rect 3158 31744 3224 31779
rect 3158 31710 3174 31744
rect 3208 31710 3224 31744
rect 3158 31675 3224 31710
rect 3158 31641 3174 31675
rect 3208 31641 3224 31675
rect 3158 31606 3224 31641
rect 3158 31572 3174 31606
rect 3208 31572 3224 31606
rect 3158 31537 3224 31572
rect 3158 31503 3174 31537
rect 3208 31503 3224 31537
rect 3158 31468 3224 31503
rect 3158 31434 3174 31468
rect 3208 31434 3224 31468
rect 3158 31399 3224 31434
rect 3158 31365 3174 31399
rect 3208 31365 3224 31399
rect 3158 31330 3224 31365
rect 3158 31296 3174 31330
rect 3208 31296 3224 31330
rect 3158 31261 3224 31296
rect 3158 31227 3174 31261
rect 3208 31227 3224 31261
rect 3158 31192 3224 31227
rect 3158 31158 3174 31192
rect 3208 31158 3224 31192
rect 3158 31123 3224 31158
rect 3158 31089 3174 31123
rect 3208 31089 3224 31123
rect 3158 31054 3224 31089
rect 3158 31020 3174 31054
rect 3208 31020 3224 31054
rect 3158 30985 3224 31020
rect 3158 30951 3174 30985
rect 3208 30951 3224 30985
rect 3158 30916 3224 30951
rect 3158 30882 3174 30916
rect 3208 30882 3224 30916
rect 3158 30847 3224 30882
rect 3158 30813 3174 30847
rect 3208 30813 3224 30847
rect 3158 30778 3224 30813
rect 3158 30744 3174 30778
rect 3208 30744 3224 30778
rect 3158 30709 3224 30744
rect 3158 30675 3174 30709
rect 3208 30675 3224 30709
rect 3158 30640 3224 30675
rect 3158 30606 3174 30640
rect 3208 30606 3224 30640
rect 3158 30571 3224 30606
rect 3158 30537 3174 30571
rect 3208 30537 3224 30571
rect 3158 30502 3224 30537
rect 3158 30468 3174 30502
rect 3208 30468 3224 30502
rect 3158 30433 3224 30468
rect 3158 30399 3174 30433
rect 3208 30399 3224 30433
rect 3158 30383 3224 30399
rect 3604 30123 5260 30139
rect 3604 30089 3620 30123
rect 3654 30089 3690 30123
rect 3724 30089 3760 30123
rect 3794 30089 3830 30123
rect 3864 30089 3899 30123
rect 3933 30089 3968 30123
rect 4002 30089 4037 30123
rect 4071 30089 4106 30123
rect 4140 30089 4175 30123
rect 4209 30089 4244 30123
rect 4278 30089 4313 30123
rect 4347 30089 4382 30123
rect 4416 30089 4451 30123
rect 4485 30089 4520 30123
rect 4554 30089 4589 30123
rect 4623 30089 4658 30123
rect 4692 30089 4727 30123
rect 4761 30089 4796 30123
rect 4830 30089 4865 30123
rect 4899 30089 4934 30123
rect 4968 30089 5003 30123
rect 5037 30089 5072 30123
rect 5106 30089 5141 30123
rect 5175 30089 5210 30123
rect 5244 30089 5260 30123
rect 3604 30073 5260 30089
rect 6221 29888 6355 29904
rect 6221 29854 6237 29888
rect 6271 29854 6305 29888
rect 6339 29854 6355 29888
rect 6221 29838 6355 29854
rect 6411 29888 6545 29904
rect 6411 29854 6427 29888
rect 6461 29854 6495 29888
rect 6529 29854 6545 29888
rect 6411 29838 6545 29854
rect 3604 29269 5260 29285
rect 3604 29235 3620 29269
rect 3654 29235 3690 29269
rect 3724 29235 3760 29269
rect 3794 29235 3830 29269
rect 3864 29235 3899 29269
rect 3933 29235 3968 29269
rect 4002 29235 4037 29269
rect 4071 29235 4106 29269
rect 4140 29235 4175 29269
rect 4209 29235 4244 29269
rect 4278 29235 4313 29269
rect 4347 29235 4382 29269
rect 4416 29235 4451 29269
rect 4485 29235 4520 29269
rect 4554 29235 4589 29269
rect 4623 29235 4658 29269
rect 4692 29235 4727 29269
rect 4761 29235 4796 29269
rect 4830 29235 4865 29269
rect 4899 29235 4934 29269
rect 4968 29235 5003 29269
rect 5037 29235 5072 29269
rect 5106 29235 5141 29269
rect 5175 29235 5210 29269
rect 5244 29235 5260 29269
rect 3604 29219 5260 29235
rect 3604 29139 5260 29155
rect 3604 29105 3620 29139
rect 3654 29105 3690 29139
rect 3724 29105 3760 29139
rect 3794 29105 3830 29139
rect 3864 29105 3899 29139
rect 3933 29105 3968 29139
rect 4002 29105 4037 29139
rect 4071 29105 4106 29139
rect 4140 29105 4175 29139
rect 4209 29105 4244 29139
rect 4278 29105 4313 29139
rect 4347 29105 4382 29139
rect 4416 29105 4451 29139
rect 4485 29105 4520 29139
rect 4554 29105 4589 29139
rect 4623 29105 4658 29139
rect 4692 29105 4727 29139
rect 4761 29105 4796 29139
rect 4830 29105 4865 29139
rect 4899 29105 4934 29139
rect 4968 29105 5003 29139
rect 5037 29105 5072 29139
rect 5106 29105 5141 29139
rect 5175 29105 5210 29139
rect 5244 29105 5260 29139
rect 3604 29089 5260 29105
rect 4398 26199 5590 26215
rect 4398 26165 4414 26199
rect 4448 26165 4485 26199
rect 4519 26165 4556 26199
rect 4590 26165 4627 26199
rect 4661 26165 4698 26199
rect 4732 26165 4769 26199
rect 4803 26165 4840 26199
rect 4874 26165 4910 26199
rect 4944 26165 4980 26199
rect 5014 26165 5050 26199
rect 5084 26165 5120 26199
rect 5154 26165 5190 26199
rect 5224 26165 5260 26199
rect 5294 26165 5330 26199
rect 5364 26165 5400 26199
rect 5434 26165 5470 26199
rect 5504 26165 5540 26199
rect 5574 26165 5590 26199
rect 4398 26149 5590 26165
rect 4872 23701 4938 23717
rect 4872 23667 4888 23701
rect 4922 23667 4938 23701
rect 4872 23631 4938 23667
rect 4872 23597 4888 23631
rect 4922 23597 4938 23631
rect 4872 23561 4938 23597
rect 4872 23527 4888 23561
rect 4922 23527 4938 23561
rect 4872 23491 4938 23527
rect 4872 23457 4888 23491
rect 4922 23457 4938 23491
rect 4872 23421 4938 23457
rect 4872 23387 4888 23421
rect 4922 23387 4938 23421
rect 4872 23351 4938 23387
rect 4872 23317 4888 23351
rect 4922 23317 4938 23351
rect 4872 23281 4938 23317
rect 4872 23247 4888 23281
rect 4922 23247 4938 23281
rect 4872 23211 4938 23247
rect 4872 23177 4888 23211
rect 4922 23177 4938 23211
rect 4872 23141 4938 23177
rect 4872 23107 4888 23141
rect 4922 23107 4938 23141
rect 4872 23071 4938 23107
rect 4872 23037 4888 23071
rect 4922 23037 4938 23071
rect 4872 23001 4938 23037
rect 4872 22967 4888 23001
rect 4922 22967 4938 23001
rect 4872 22931 4938 22967
rect 4872 22897 4888 22931
rect 4922 22897 4938 22931
rect 4872 22861 4938 22897
rect 4872 22827 4888 22861
rect 4922 22827 4938 22861
rect 4872 22791 4938 22827
rect 4872 22757 4888 22791
rect 4922 22757 4938 22791
rect 4872 22721 4938 22757
rect 4872 22687 4888 22721
rect 4922 22687 4938 22721
rect 4872 22651 4938 22687
rect 4872 22617 4888 22651
rect 4922 22617 4938 22651
rect 4872 22581 4938 22617
rect 4872 22547 4888 22581
rect 4922 22547 4938 22581
rect 4872 22512 4938 22547
rect 4872 22478 4888 22512
rect 4922 22478 4938 22512
rect 4872 22443 4938 22478
rect 4872 22409 4888 22443
rect 4922 22409 4938 22443
rect 4872 22374 4938 22409
rect 4872 22340 4888 22374
rect 4922 22340 4938 22374
rect 4872 22305 4938 22340
rect 4872 22271 4888 22305
rect 4922 22271 4938 22305
rect 4872 22236 4938 22271
rect 4872 22202 4888 22236
rect 4922 22202 4938 22236
rect 4872 22167 4938 22202
rect 4872 22133 4888 22167
rect 4922 22133 4938 22167
rect 4872 22098 4938 22133
rect 4872 22064 4888 22098
rect 4922 22064 4938 22098
rect 4872 22029 4938 22064
rect 4872 21995 4888 22029
rect 4922 21995 4938 22029
rect 4872 21960 4938 21995
rect 4872 21926 4888 21960
rect 4922 21926 4938 21960
rect 4872 21891 4938 21926
rect 4872 21857 4888 21891
rect 4922 21857 4938 21891
rect 4872 21822 4938 21857
rect 4872 21788 4888 21822
rect 4922 21788 4938 21822
rect 4872 21753 4938 21788
rect 4872 21719 4888 21753
rect 4922 21719 4938 21753
rect 4872 21684 4938 21719
rect 4872 21650 4888 21684
rect 4922 21650 4938 21684
rect 4872 21615 4938 21650
rect 4872 21581 4888 21615
rect 4922 21581 4938 21615
rect 4872 21546 4938 21581
rect 4872 21512 4888 21546
rect 4922 21512 4938 21546
rect 4872 21477 4938 21512
rect 4872 21443 4888 21477
rect 4922 21443 4938 21477
rect 4872 21408 4938 21443
rect 4872 21374 4888 21408
rect 4922 21374 4938 21408
rect 4872 21339 4938 21374
rect 4872 21305 4888 21339
rect 4922 21305 4938 21339
rect 4872 21270 4938 21305
rect 4872 21236 4888 21270
rect 4922 21236 4938 21270
rect 4872 21201 4938 21236
rect 4872 21167 4888 21201
rect 4922 21167 4938 21201
rect 4872 21132 4938 21167
rect 4872 21098 4888 21132
rect 4922 21098 4938 21132
rect 4872 21063 4938 21098
rect 4872 21029 4888 21063
rect 4922 21029 4938 21063
rect 4872 20994 4938 21029
rect 4872 20960 4888 20994
rect 4922 20960 4938 20994
rect 4872 20925 4938 20960
rect 4872 20891 4888 20925
rect 4922 20891 4938 20925
rect 4872 20856 4938 20891
rect 4872 20822 4888 20856
rect 4922 20822 4938 20856
rect 4872 20787 4938 20822
rect 4872 20753 4888 20787
rect 4922 20753 4938 20787
rect 4872 20718 4938 20753
rect 4872 20684 4888 20718
rect 4922 20684 4938 20718
rect 4872 20649 4938 20684
rect 4872 20615 4888 20649
rect 4922 20615 4938 20649
rect 4872 20580 4938 20615
rect 4872 20546 4888 20580
rect 4922 20546 4938 20580
rect 4872 20511 4938 20546
rect 4872 20477 4888 20511
rect 4922 20477 4938 20511
rect 4872 20461 4938 20477
rect 5180 23701 5246 23717
rect 5180 23667 5196 23701
rect 5230 23667 5246 23701
rect 5180 23631 5246 23667
rect 5180 23597 5196 23631
rect 5230 23597 5246 23631
rect 5180 23562 5246 23597
rect 5180 23528 5196 23562
rect 5230 23528 5246 23562
rect 5180 23493 5246 23528
rect 5180 23459 5196 23493
rect 5230 23459 5246 23493
rect 5180 23424 5246 23459
rect 5180 23390 5196 23424
rect 5230 23390 5246 23424
rect 5180 23355 5246 23390
rect 5180 23321 5196 23355
rect 5230 23321 5246 23355
rect 5180 23286 5246 23321
rect 5180 23252 5196 23286
rect 5230 23252 5246 23286
rect 5180 23217 5246 23252
rect 5180 23183 5196 23217
rect 5230 23183 5246 23217
rect 5180 23148 5246 23183
rect 5180 23114 5196 23148
rect 5230 23114 5246 23148
rect 5180 23079 5246 23114
rect 5180 23045 5196 23079
rect 5230 23045 5246 23079
rect 5180 23010 5246 23045
rect 5180 22976 5196 23010
rect 5230 22976 5246 23010
rect 5180 22941 5246 22976
rect 5180 22907 5196 22941
rect 5230 22907 5246 22941
rect 5180 22872 5246 22907
rect 5180 22838 5196 22872
rect 5230 22838 5246 22872
rect 5180 22803 5246 22838
rect 5180 22769 5196 22803
rect 5230 22769 5246 22803
rect 5180 22734 5246 22769
rect 5180 22700 5196 22734
rect 5230 22700 5246 22734
rect 5180 22665 5246 22700
rect 5180 22631 5196 22665
rect 5230 22631 5246 22665
rect 5180 22596 5246 22631
rect 5180 22562 5196 22596
rect 5230 22562 5246 22596
rect 5180 22527 5246 22562
rect 5180 22493 5196 22527
rect 5230 22493 5246 22527
rect 5180 22458 5246 22493
rect 5180 22424 5196 22458
rect 5230 22424 5246 22458
rect 5180 22389 5246 22424
rect 5180 22355 5196 22389
rect 5230 22355 5246 22389
rect 5180 22320 5246 22355
rect 5180 22286 5196 22320
rect 5230 22286 5246 22320
rect 5180 22251 5246 22286
rect 5180 22217 5196 22251
rect 5230 22217 5246 22251
rect 5180 22182 5246 22217
rect 5180 22148 5196 22182
rect 5230 22148 5246 22182
rect 5180 22113 5246 22148
rect 5180 22079 5196 22113
rect 5230 22079 5246 22113
rect 5180 22044 5246 22079
rect 5180 22010 5196 22044
rect 5230 22010 5246 22044
rect 5180 21975 5246 22010
rect 5180 21941 5196 21975
rect 5230 21941 5246 21975
rect 5180 21906 5246 21941
rect 5180 21872 5196 21906
rect 5230 21872 5246 21906
rect 5180 21837 5246 21872
rect 5180 21803 5196 21837
rect 5230 21803 5246 21837
rect 5180 21768 5246 21803
rect 5180 21734 5196 21768
rect 5230 21734 5246 21768
rect 5180 21699 5246 21734
rect 5180 21665 5196 21699
rect 5230 21665 5246 21699
rect 5180 21630 5246 21665
rect 5180 21596 5196 21630
rect 5230 21596 5246 21630
rect 5180 21561 5246 21596
rect 5180 21527 5196 21561
rect 5230 21527 5246 21561
rect 5180 21492 5246 21527
rect 5180 21458 5196 21492
rect 5230 21458 5246 21492
rect 5180 21423 5246 21458
rect 5180 21389 5196 21423
rect 5230 21389 5246 21423
rect 5180 21354 5246 21389
rect 5180 21320 5196 21354
rect 5230 21320 5246 21354
rect 5180 21285 5246 21320
rect 5180 21251 5196 21285
rect 5230 21251 5246 21285
rect 5180 21216 5246 21251
rect 5180 21182 5196 21216
rect 5230 21182 5246 21216
rect 5180 21147 5246 21182
rect 5180 21113 5196 21147
rect 5230 21113 5246 21147
rect 5180 21078 5246 21113
rect 5180 21044 5196 21078
rect 5230 21044 5246 21078
rect 5180 21009 5246 21044
rect 5180 20975 5196 21009
rect 5230 20975 5246 21009
rect 5180 20940 5246 20975
rect 5180 20906 5196 20940
rect 5230 20906 5246 20940
rect 5180 20871 5246 20906
rect 5180 20837 5196 20871
rect 5230 20837 5246 20871
rect 5180 20802 5246 20837
rect 5180 20768 5196 20802
rect 5230 20768 5246 20802
rect 5180 20733 5246 20768
rect 5180 20699 5196 20733
rect 5230 20699 5246 20733
rect 5180 20664 5246 20699
rect 5180 20630 5196 20664
rect 5230 20630 5246 20664
rect 5180 20595 5246 20630
rect 5180 20561 5196 20595
rect 5230 20561 5246 20595
rect 5180 20526 5246 20561
rect 5180 20492 5196 20526
rect 5230 20492 5246 20526
rect 5180 20457 5246 20492
rect 5180 20423 5196 20457
rect 5230 20423 5246 20457
rect 5180 20388 5246 20423
rect 5180 20354 5196 20388
rect 5230 20354 5246 20388
rect 5180 20319 5246 20354
rect 5180 20285 5196 20319
rect 5230 20285 5246 20319
rect 5180 20250 5246 20285
rect 5180 20216 5196 20250
rect 5230 20216 5246 20250
rect 5180 20181 5246 20216
rect 5180 20147 5196 20181
rect 5230 20147 5246 20181
rect 5180 20112 5246 20147
rect 5180 20078 5196 20112
rect 5230 20078 5246 20112
rect 4883 20032 4949 20048
rect 4883 19998 4899 20032
rect 4933 19998 4949 20032
rect 4883 19961 4949 19998
rect 4883 19927 4899 19961
rect 4933 19927 4949 19961
rect 4883 19890 4949 19927
rect 4883 19856 4899 19890
rect 4933 19856 4949 19890
rect 4883 19818 4949 19856
rect 4883 19784 4899 19818
rect 4933 19784 4949 19818
rect 4883 19746 4949 19784
rect 4883 19712 4899 19746
rect 4933 19712 4949 19746
rect 5180 20043 5246 20078
rect 5180 20009 5196 20043
rect 5230 20009 5246 20043
rect 5180 19974 5246 20009
rect 5180 19940 5196 19974
rect 5230 19940 5246 19974
rect 5180 19905 5246 19940
rect 5180 19871 5196 19905
rect 5230 19871 5246 19905
rect 5180 19836 5246 19871
rect 5180 19802 5196 19836
rect 5230 19802 5246 19836
rect 5180 19767 5246 19802
rect 5180 19733 5196 19767
rect 5230 19733 5246 19767
rect 5180 19717 5246 19733
rect 5436 23701 5502 23717
rect 5436 23667 5452 23701
rect 5486 23667 5502 23701
rect 5436 23631 5502 23667
rect 5436 23597 5452 23631
rect 5486 23597 5502 23631
rect 5436 23562 5502 23597
rect 5436 23528 5452 23562
rect 5486 23528 5502 23562
rect 5436 23493 5502 23528
rect 5436 23459 5452 23493
rect 5486 23459 5502 23493
rect 5436 23424 5502 23459
rect 5436 23390 5452 23424
rect 5486 23390 5502 23424
rect 5436 23355 5502 23390
rect 5436 23321 5452 23355
rect 5486 23321 5502 23355
rect 5436 23286 5502 23321
rect 5436 23252 5452 23286
rect 5486 23252 5502 23286
rect 5436 23217 5502 23252
rect 5436 23183 5452 23217
rect 5486 23183 5502 23217
rect 5436 23148 5502 23183
rect 5436 23114 5452 23148
rect 5486 23114 5502 23148
rect 5436 23079 5502 23114
rect 5436 23045 5452 23079
rect 5486 23045 5502 23079
rect 5436 23010 5502 23045
rect 5436 22976 5452 23010
rect 5486 22976 5502 23010
rect 5436 22941 5502 22976
rect 5436 22907 5452 22941
rect 5486 22907 5502 22941
rect 5436 22872 5502 22907
rect 5436 22838 5452 22872
rect 5486 22838 5502 22872
rect 5436 22803 5502 22838
rect 5436 22769 5452 22803
rect 5486 22769 5502 22803
rect 5436 22734 5502 22769
rect 5436 22700 5452 22734
rect 5486 22700 5502 22734
rect 5436 22665 5502 22700
rect 5436 22631 5452 22665
rect 5486 22631 5502 22665
rect 5436 22596 5502 22631
rect 5436 22562 5452 22596
rect 5486 22562 5502 22596
rect 5436 22527 5502 22562
rect 5436 22493 5452 22527
rect 5486 22493 5502 22527
rect 5436 22458 5502 22493
rect 5436 22424 5452 22458
rect 5486 22424 5502 22458
rect 5436 22389 5502 22424
rect 5436 22355 5452 22389
rect 5486 22355 5502 22389
rect 5436 22320 5502 22355
rect 5436 22286 5452 22320
rect 5486 22286 5502 22320
rect 5436 22251 5502 22286
rect 5436 22217 5452 22251
rect 5486 22217 5502 22251
rect 5436 22182 5502 22217
rect 5436 22148 5452 22182
rect 5486 22148 5502 22182
rect 5436 22113 5502 22148
rect 5436 22079 5452 22113
rect 5486 22079 5502 22113
rect 5436 22044 5502 22079
rect 5436 22010 5452 22044
rect 5486 22010 5502 22044
rect 5436 21975 5502 22010
rect 5436 21941 5452 21975
rect 5486 21941 5502 21975
rect 5436 21906 5502 21941
rect 5436 21872 5452 21906
rect 5486 21872 5502 21906
rect 5436 21837 5502 21872
rect 5436 21803 5452 21837
rect 5486 21803 5502 21837
rect 5436 21768 5502 21803
rect 5436 21734 5452 21768
rect 5486 21734 5502 21768
rect 5436 21699 5502 21734
rect 5436 21665 5452 21699
rect 5486 21665 5502 21699
rect 5436 21630 5502 21665
rect 5436 21596 5452 21630
rect 5486 21596 5502 21630
rect 5436 21561 5502 21596
rect 5436 21527 5452 21561
rect 5486 21527 5502 21561
rect 5436 21492 5502 21527
rect 5436 21458 5452 21492
rect 5486 21458 5502 21492
rect 5436 21423 5502 21458
rect 5436 21389 5452 21423
rect 5486 21389 5502 21423
rect 5436 21354 5502 21389
rect 5436 21320 5452 21354
rect 5486 21320 5502 21354
rect 5436 21285 5502 21320
rect 5436 21251 5452 21285
rect 5486 21251 5502 21285
rect 5436 21216 5502 21251
rect 5436 21182 5452 21216
rect 5486 21182 5502 21216
rect 5436 21147 5502 21182
rect 5436 21113 5452 21147
rect 5486 21113 5502 21147
rect 5436 21078 5502 21113
rect 5436 21044 5452 21078
rect 5486 21044 5502 21078
rect 5436 21009 5502 21044
rect 5436 20975 5452 21009
rect 5486 20975 5502 21009
rect 5436 20940 5502 20975
rect 5436 20906 5452 20940
rect 5486 20906 5502 20940
rect 5436 20871 5502 20906
rect 5436 20837 5452 20871
rect 5486 20837 5502 20871
rect 5436 20802 5502 20837
rect 5436 20768 5452 20802
rect 5486 20768 5502 20802
rect 5436 20733 5502 20768
rect 5436 20699 5452 20733
rect 5486 20699 5502 20733
rect 5436 20664 5502 20699
rect 5436 20630 5452 20664
rect 5486 20630 5502 20664
rect 5436 20595 5502 20630
rect 5436 20561 5452 20595
rect 5486 20561 5502 20595
rect 5436 20526 5502 20561
rect 5436 20492 5452 20526
rect 5486 20492 5502 20526
rect 5436 20457 5502 20492
rect 5436 20423 5452 20457
rect 5486 20423 5502 20457
rect 5436 20388 5502 20423
rect 5436 20354 5452 20388
rect 5486 20354 5502 20388
rect 5436 20319 5502 20354
rect 5436 20285 5452 20319
rect 5486 20285 5502 20319
rect 5436 20250 5502 20285
rect 5436 20216 5452 20250
rect 5486 20216 5502 20250
rect 5436 20181 5502 20216
rect 5436 20147 5452 20181
rect 5486 20147 5502 20181
rect 5436 20112 5502 20147
rect 5436 20078 5452 20112
rect 5486 20078 5502 20112
rect 5436 20043 5502 20078
rect 5436 20009 5452 20043
rect 5486 20009 5502 20043
rect 5436 19974 5502 20009
rect 5436 19940 5452 19974
rect 5486 19940 5502 19974
rect 5436 19905 5502 19940
rect 5436 19871 5452 19905
rect 5486 19871 5502 19905
rect 5436 19836 5502 19871
rect 5436 19802 5452 19836
rect 5486 19802 5502 19836
rect 5436 19767 5502 19802
rect 5436 19733 5452 19767
rect 5486 19733 5502 19767
rect 5436 19717 5502 19733
rect 7347 22034 7481 22050
rect 7347 22000 7363 22034
rect 7397 22000 7431 22034
rect 7465 22000 7481 22034
rect 7347 21984 7481 22000
rect 7537 22034 7671 22050
rect 7537 22000 7553 22034
rect 7587 22000 7621 22034
rect 7655 22000 7671 22034
rect 7537 21984 7671 22000
rect 4883 19674 4949 19712
rect 4883 19640 4899 19674
rect 4933 19640 4949 19674
rect 4883 19602 4949 19640
rect 4883 19568 4899 19602
rect 4933 19568 4949 19602
rect 4883 19530 4949 19568
rect 4883 19496 4899 19530
rect 4933 19496 4949 19530
rect 4883 19480 4949 19496
rect 5042 19068 5242 19084
rect 5042 19034 5058 19068
rect 5092 19034 5192 19068
rect 5226 19034 5242 19068
rect 5042 19018 5242 19034
rect 3536 17684 3602 17700
rect 3536 17650 3552 17684
rect 3586 17650 3602 17684
rect 3428 17599 3494 17615
rect 3428 17565 3444 17599
rect 3478 17565 3494 17599
rect 3428 17530 3494 17565
rect 3428 17496 3444 17530
rect 3478 17496 3494 17530
rect 3428 17461 3494 17496
rect 3428 17427 3444 17461
rect 3478 17427 3494 17461
rect 3428 17392 3494 17427
rect 3428 17358 3444 17392
rect 3478 17358 3494 17392
rect 3428 17323 3494 17358
rect 3428 17289 3444 17323
rect 3478 17289 3494 17323
rect 3428 17254 3494 17289
rect 3428 17220 3444 17254
rect 3478 17220 3494 17254
rect 3428 17185 3494 17220
rect 3428 17151 3444 17185
rect 3478 17151 3494 17185
rect 3428 17115 3494 17151
rect 3536 17613 3602 17650
rect 3536 17579 3552 17613
rect 3586 17579 3602 17613
rect 3536 17542 3602 17579
rect 3536 17508 3552 17542
rect 3586 17508 3602 17542
rect 3536 17470 3602 17508
rect 3536 17436 3552 17470
rect 3586 17436 3602 17470
rect 3536 17398 3602 17436
rect 3536 17364 3552 17398
rect 3586 17364 3602 17398
rect 3536 17326 3602 17364
rect 3536 17292 3552 17326
rect 3586 17292 3602 17326
rect 3536 17254 3602 17292
rect 3536 17220 3552 17254
rect 3586 17220 3602 17254
rect 3536 17182 3602 17220
rect 3536 17148 3552 17182
rect 3586 17148 3602 17182
rect 3536 17132 3602 17148
rect 3428 17081 3444 17115
rect 3478 17081 3494 17115
rect 3428 17045 3494 17081
rect 3428 17011 3444 17045
rect 3478 17011 3494 17045
rect 3428 16975 3494 17011
rect 3428 16941 3444 16975
rect 3478 16941 3494 16975
rect 3428 16905 3494 16941
rect 3428 16871 3444 16905
rect 3478 16871 3494 16905
rect 3428 16835 3494 16871
rect 3428 16801 3444 16835
rect 3478 16801 3494 16835
rect 4269 16867 4837 16883
rect 4269 16833 4285 16867
rect 4319 16833 4357 16867
rect 4391 16833 4429 16867
rect 4463 16833 4501 16867
rect 4535 16833 4573 16867
rect 4607 16833 4645 16867
rect 4679 16833 4716 16867
rect 4750 16833 4787 16867
rect 4821 16833 4837 16867
rect 4269 16817 4837 16833
rect 4893 16867 5461 16883
rect 4893 16833 4909 16867
rect 4943 16833 4981 16867
rect 5015 16833 5053 16867
rect 5087 16833 5125 16867
rect 5159 16833 5197 16867
rect 5231 16833 5269 16867
rect 5303 16833 5340 16867
rect 5374 16833 5411 16867
rect 5445 16833 5461 16867
rect 4893 16817 5461 16833
rect 3428 16765 3494 16801
rect 3428 16731 3444 16765
rect 3478 16731 3494 16765
rect 3428 16695 3494 16731
rect 3428 16661 3444 16695
rect 3478 16661 3494 16695
rect 3428 16625 3494 16661
rect 3428 16591 3444 16625
rect 3478 16591 3494 16625
rect 3428 16555 3494 16591
rect 3428 16521 3444 16555
rect 3478 16521 3494 16555
rect 3428 16485 3494 16521
rect 3428 16451 3444 16485
rect 3478 16451 3494 16485
rect 3428 16415 3494 16451
rect 3428 16381 3444 16415
rect 3478 16381 3494 16415
rect 3428 16345 3494 16381
rect 3428 16311 3444 16345
rect 3478 16311 3494 16345
rect 3428 16275 3494 16311
rect 3428 16241 3444 16275
rect 3478 16241 3494 16275
rect 3428 16205 3494 16241
rect 3428 16171 3444 16205
rect 3478 16171 3494 16205
rect 3428 16135 3494 16171
rect 3428 16101 3444 16135
rect 3478 16101 3494 16135
rect 3428 16065 3494 16101
rect 3428 16031 3444 16065
rect 3478 16031 3494 16065
rect 3428 16015 3494 16031
rect 4235 16095 5835 16111
rect 4235 16061 4251 16095
rect 4285 16061 4320 16095
rect 4354 16061 4389 16095
rect 4423 16061 4458 16095
rect 4492 16061 4527 16095
rect 4561 16061 4596 16095
rect 4630 16061 4665 16095
rect 4699 16061 4735 16095
rect 4769 16061 4805 16095
rect 4839 16061 4875 16095
rect 4909 16061 4945 16095
rect 4979 16061 5015 16095
rect 5049 16061 5085 16095
rect 5119 16061 5155 16095
rect 5189 16061 5225 16095
rect 5259 16061 5295 16095
rect 5329 16061 5365 16095
rect 5399 16061 5435 16095
rect 5469 16061 5505 16095
rect 5539 16061 5575 16095
rect 5609 16061 5645 16095
rect 5679 16061 5715 16095
rect 5749 16061 5785 16095
rect 5819 16061 5835 16095
rect 4235 16045 5835 16061
rect 4235 15365 5835 15381
rect 4235 15331 4251 15365
rect 4285 15331 4320 15365
rect 4354 15331 4389 15365
rect 4423 15331 4458 15365
rect 4492 15331 4527 15365
rect 4561 15331 4596 15365
rect 4630 15331 4665 15365
rect 4699 15331 4735 15365
rect 4769 15331 4805 15365
rect 4839 15331 4875 15365
rect 4909 15331 4945 15365
rect 4979 15331 5015 15365
rect 5049 15331 5085 15365
rect 5119 15331 5155 15365
rect 5189 15331 5225 15365
rect 5259 15331 5295 15365
rect 5329 15331 5365 15365
rect 5399 15331 5435 15365
rect 5469 15331 5505 15365
rect 5539 15331 5575 15365
rect 5609 15331 5645 15365
rect 5679 15331 5715 15365
rect 5749 15331 5785 15365
rect 5819 15331 5835 15365
rect 4235 15315 5835 15331
<< polycont >>
rect 3174 39397 3208 39431
rect 3174 39329 3208 39363
rect 3174 39261 3208 39295
rect 3174 39193 3208 39227
rect 3174 39125 3208 39159
rect 3174 39057 3208 39091
rect 3174 38989 3208 39023
rect 3174 38921 3208 38955
rect 3174 38853 3208 38887
rect 3174 38785 3208 38819
rect 3174 38717 3208 38751
rect 3174 38649 3208 38683
rect 3174 38581 3208 38615
rect 3174 38513 3208 38547
rect 3174 38445 3208 38479
rect 3174 38377 3208 38411
rect 3174 38309 3208 38343
rect 3174 38241 3208 38275
rect 3174 38173 3208 38207
rect 3174 38105 3208 38139
rect 3174 38037 3208 38071
rect 3174 37969 3208 38003
rect 3174 37901 3208 37935
rect 3174 37833 3208 37867
rect 3174 37765 3208 37799
rect 3174 37697 3208 37731
rect 3174 37629 3208 37663
rect 3174 37561 3208 37595
rect 3174 37493 3208 37527
rect 3174 37425 3208 37459
rect 3174 37357 3208 37391
rect 3174 37289 3208 37323
rect 3174 37221 3208 37255
rect 3174 37153 3208 37187
rect 3174 37085 3208 37119
rect 3174 37017 3208 37051
rect 3174 36949 3208 36983
rect 3174 36881 3208 36915
rect 3174 36813 3208 36847
rect 3174 36745 3208 36779
rect 3174 36677 3208 36711
rect 3174 36609 3208 36643
rect 3174 36541 3208 36575
rect 3174 36473 3208 36507
rect 3174 36405 3208 36439
rect 3174 36337 3208 36371
rect 3174 36269 3208 36303
rect 3174 36201 3208 36235
rect 3174 36133 3208 36167
rect 3174 36065 3208 36099
rect 3174 35997 3208 36031
rect 3174 35929 3208 35963
rect 3174 35861 3208 35895
rect 3174 35793 3208 35827
rect 3174 35725 3208 35759
rect 3174 35657 3208 35691
rect 3174 35589 3208 35623
rect 3174 35521 3208 35555
rect 3174 35453 3208 35487
rect 3174 35385 3208 35419
rect 3174 35317 3208 35351
rect 3174 35249 3208 35283
rect 3174 35181 3208 35215
rect 3174 35113 3208 35147
rect 3174 35045 3208 35079
rect 3174 34977 3208 35011
rect 3174 34909 3208 34943
rect 3174 34841 3208 34875
rect 3174 34773 3208 34807
rect 3174 34705 3208 34739
rect 3174 34637 3208 34671
rect 3174 34569 3208 34603
rect 3174 34501 3208 34535
rect 3174 34433 3208 34467
rect 3174 34365 3208 34399
rect 3174 34297 3208 34331
rect 3174 34229 3208 34263
rect 3174 34161 3208 34195
rect 3174 34093 3208 34127
rect 3174 34025 3208 34059
rect 3174 33957 3208 33991
rect 3174 33889 3208 33923
rect 3174 33821 3208 33855
rect 3174 33753 3208 33787
rect 3174 33685 3208 33719
rect 3174 33617 3208 33651
rect 3174 33549 3208 33583
rect 3174 33481 3208 33515
rect 3174 33413 3208 33447
rect 3174 33345 3208 33379
rect 3174 33277 3208 33311
rect 3174 33209 3208 33243
rect 3174 33141 3208 33175
rect 3174 33073 3208 33107
rect 3174 33005 3208 33039
rect 3174 32937 3208 32971
rect 3174 32869 3208 32903
rect 3174 32801 3208 32835
rect 3174 32733 3208 32767
rect 3174 32665 3208 32699
rect 3174 32597 3208 32631
rect 3174 32529 3208 32563
rect 3174 32461 3208 32495
rect 3174 32393 3208 32427
rect 3174 32325 3208 32359
rect 3174 32257 3208 32291
rect 3174 32189 3208 32223
rect 3174 32121 3208 32155
rect 3174 32053 3208 32087
rect 3174 31985 3208 32019
rect 3174 31917 3208 31951
rect 3174 31848 3208 31882
rect 3174 31779 3208 31813
rect 3174 31710 3208 31744
rect 3174 31641 3208 31675
rect 3174 31572 3208 31606
rect 3174 31503 3208 31537
rect 3174 31434 3208 31468
rect 3174 31365 3208 31399
rect 3174 31296 3208 31330
rect 3174 31227 3208 31261
rect 3174 31158 3208 31192
rect 3174 31089 3208 31123
rect 3174 31020 3208 31054
rect 3174 30951 3208 30985
rect 3174 30882 3208 30916
rect 3174 30813 3208 30847
rect 3174 30744 3208 30778
rect 3174 30675 3208 30709
rect 3174 30606 3208 30640
rect 3174 30537 3208 30571
rect 3174 30468 3208 30502
rect 3174 30399 3208 30433
rect 3620 30089 3654 30123
rect 3690 30089 3724 30123
rect 3760 30089 3794 30123
rect 3830 30089 3864 30123
rect 3899 30089 3933 30123
rect 3968 30089 4002 30123
rect 4037 30089 4071 30123
rect 4106 30089 4140 30123
rect 4175 30089 4209 30123
rect 4244 30089 4278 30123
rect 4313 30089 4347 30123
rect 4382 30089 4416 30123
rect 4451 30089 4485 30123
rect 4520 30089 4554 30123
rect 4589 30089 4623 30123
rect 4658 30089 4692 30123
rect 4727 30089 4761 30123
rect 4796 30089 4830 30123
rect 4865 30089 4899 30123
rect 4934 30089 4968 30123
rect 5003 30089 5037 30123
rect 5072 30089 5106 30123
rect 5141 30089 5175 30123
rect 5210 30089 5244 30123
rect 6237 29854 6271 29888
rect 6305 29854 6339 29888
rect 6427 29854 6461 29888
rect 6495 29854 6529 29888
rect 3620 29235 3654 29269
rect 3690 29235 3724 29269
rect 3760 29235 3794 29269
rect 3830 29235 3864 29269
rect 3899 29235 3933 29269
rect 3968 29235 4002 29269
rect 4037 29235 4071 29269
rect 4106 29235 4140 29269
rect 4175 29235 4209 29269
rect 4244 29235 4278 29269
rect 4313 29235 4347 29269
rect 4382 29235 4416 29269
rect 4451 29235 4485 29269
rect 4520 29235 4554 29269
rect 4589 29235 4623 29269
rect 4658 29235 4692 29269
rect 4727 29235 4761 29269
rect 4796 29235 4830 29269
rect 4865 29235 4899 29269
rect 4934 29235 4968 29269
rect 5003 29235 5037 29269
rect 5072 29235 5106 29269
rect 5141 29235 5175 29269
rect 5210 29235 5244 29269
rect 3620 29105 3654 29139
rect 3690 29105 3724 29139
rect 3760 29105 3794 29139
rect 3830 29105 3864 29139
rect 3899 29105 3933 29139
rect 3968 29105 4002 29139
rect 4037 29105 4071 29139
rect 4106 29105 4140 29139
rect 4175 29105 4209 29139
rect 4244 29105 4278 29139
rect 4313 29105 4347 29139
rect 4382 29105 4416 29139
rect 4451 29105 4485 29139
rect 4520 29105 4554 29139
rect 4589 29105 4623 29139
rect 4658 29105 4692 29139
rect 4727 29105 4761 29139
rect 4796 29105 4830 29139
rect 4865 29105 4899 29139
rect 4934 29105 4968 29139
rect 5003 29105 5037 29139
rect 5072 29105 5106 29139
rect 5141 29105 5175 29139
rect 5210 29105 5244 29139
rect 4414 26165 4448 26199
rect 4485 26165 4519 26199
rect 4556 26165 4590 26199
rect 4627 26165 4661 26199
rect 4698 26165 4732 26199
rect 4769 26165 4803 26199
rect 4840 26165 4874 26199
rect 4910 26165 4944 26199
rect 4980 26165 5014 26199
rect 5050 26165 5084 26199
rect 5120 26165 5154 26199
rect 5190 26165 5224 26199
rect 5260 26165 5294 26199
rect 5330 26165 5364 26199
rect 5400 26165 5434 26199
rect 5470 26165 5504 26199
rect 5540 26165 5574 26199
rect 4888 23667 4922 23701
rect 4888 23597 4922 23631
rect 4888 23527 4922 23561
rect 4888 23457 4922 23491
rect 4888 23387 4922 23421
rect 4888 23317 4922 23351
rect 4888 23247 4922 23281
rect 4888 23177 4922 23211
rect 4888 23107 4922 23141
rect 4888 23037 4922 23071
rect 4888 22967 4922 23001
rect 4888 22897 4922 22931
rect 4888 22827 4922 22861
rect 4888 22757 4922 22791
rect 4888 22687 4922 22721
rect 4888 22617 4922 22651
rect 4888 22547 4922 22581
rect 4888 22478 4922 22512
rect 4888 22409 4922 22443
rect 4888 22340 4922 22374
rect 4888 22271 4922 22305
rect 4888 22202 4922 22236
rect 4888 22133 4922 22167
rect 4888 22064 4922 22098
rect 4888 21995 4922 22029
rect 4888 21926 4922 21960
rect 4888 21857 4922 21891
rect 4888 21788 4922 21822
rect 4888 21719 4922 21753
rect 4888 21650 4922 21684
rect 4888 21581 4922 21615
rect 4888 21512 4922 21546
rect 4888 21443 4922 21477
rect 4888 21374 4922 21408
rect 4888 21305 4922 21339
rect 4888 21236 4922 21270
rect 4888 21167 4922 21201
rect 4888 21098 4922 21132
rect 4888 21029 4922 21063
rect 4888 20960 4922 20994
rect 4888 20891 4922 20925
rect 4888 20822 4922 20856
rect 4888 20753 4922 20787
rect 4888 20684 4922 20718
rect 4888 20615 4922 20649
rect 4888 20546 4922 20580
rect 4888 20477 4922 20511
rect 5196 23667 5230 23701
rect 5196 23597 5230 23631
rect 5196 23528 5230 23562
rect 5196 23459 5230 23493
rect 5196 23390 5230 23424
rect 5196 23321 5230 23355
rect 5196 23252 5230 23286
rect 5196 23183 5230 23217
rect 5196 23114 5230 23148
rect 5196 23045 5230 23079
rect 5196 22976 5230 23010
rect 5196 22907 5230 22941
rect 5196 22838 5230 22872
rect 5196 22769 5230 22803
rect 5196 22700 5230 22734
rect 5196 22631 5230 22665
rect 5196 22562 5230 22596
rect 5196 22493 5230 22527
rect 5196 22424 5230 22458
rect 5196 22355 5230 22389
rect 5196 22286 5230 22320
rect 5196 22217 5230 22251
rect 5196 22148 5230 22182
rect 5196 22079 5230 22113
rect 5196 22010 5230 22044
rect 5196 21941 5230 21975
rect 5196 21872 5230 21906
rect 5196 21803 5230 21837
rect 5196 21734 5230 21768
rect 5196 21665 5230 21699
rect 5196 21596 5230 21630
rect 5196 21527 5230 21561
rect 5196 21458 5230 21492
rect 5196 21389 5230 21423
rect 5196 21320 5230 21354
rect 5196 21251 5230 21285
rect 5196 21182 5230 21216
rect 5196 21113 5230 21147
rect 5196 21044 5230 21078
rect 5196 20975 5230 21009
rect 5196 20906 5230 20940
rect 5196 20837 5230 20871
rect 5196 20768 5230 20802
rect 5196 20699 5230 20733
rect 5196 20630 5230 20664
rect 5196 20561 5230 20595
rect 5196 20492 5230 20526
rect 5196 20423 5230 20457
rect 5196 20354 5230 20388
rect 5196 20285 5230 20319
rect 5196 20216 5230 20250
rect 5196 20147 5230 20181
rect 5196 20078 5230 20112
rect 4899 19998 4933 20032
rect 4899 19927 4933 19961
rect 4899 19856 4933 19890
rect 4899 19784 4933 19818
rect 4899 19712 4933 19746
rect 5196 20009 5230 20043
rect 5196 19940 5230 19974
rect 5196 19871 5230 19905
rect 5196 19802 5230 19836
rect 5196 19733 5230 19767
rect 5452 23667 5486 23701
rect 5452 23597 5486 23631
rect 5452 23528 5486 23562
rect 5452 23459 5486 23493
rect 5452 23390 5486 23424
rect 5452 23321 5486 23355
rect 5452 23252 5486 23286
rect 5452 23183 5486 23217
rect 5452 23114 5486 23148
rect 5452 23045 5486 23079
rect 5452 22976 5486 23010
rect 5452 22907 5486 22941
rect 5452 22838 5486 22872
rect 5452 22769 5486 22803
rect 5452 22700 5486 22734
rect 5452 22631 5486 22665
rect 5452 22562 5486 22596
rect 5452 22493 5486 22527
rect 5452 22424 5486 22458
rect 5452 22355 5486 22389
rect 5452 22286 5486 22320
rect 5452 22217 5486 22251
rect 5452 22148 5486 22182
rect 5452 22079 5486 22113
rect 5452 22010 5486 22044
rect 5452 21941 5486 21975
rect 5452 21872 5486 21906
rect 5452 21803 5486 21837
rect 5452 21734 5486 21768
rect 5452 21665 5486 21699
rect 5452 21596 5486 21630
rect 5452 21527 5486 21561
rect 5452 21458 5486 21492
rect 5452 21389 5486 21423
rect 5452 21320 5486 21354
rect 5452 21251 5486 21285
rect 5452 21182 5486 21216
rect 5452 21113 5486 21147
rect 5452 21044 5486 21078
rect 5452 20975 5486 21009
rect 5452 20906 5486 20940
rect 5452 20837 5486 20871
rect 5452 20768 5486 20802
rect 5452 20699 5486 20733
rect 5452 20630 5486 20664
rect 5452 20561 5486 20595
rect 5452 20492 5486 20526
rect 5452 20423 5486 20457
rect 5452 20354 5486 20388
rect 5452 20285 5486 20319
rect 5452 20216 5486 20250
rect 5452 20147 5486 20181
rect 5452 20078 5486 20112
rect 5452 20009 5486 20043
rect 5452 19940 5486 19974
rect 5452 19871 5486 19905
rect 5452 19802 5486 19836
rect 5452 19733 5486 19767
rect 7363 22000 7397 22034
rect 7431 22000 7465 22034
rect 7553 22000 7587 22034
rect 7621 22000 7655 22034
rect 4899 19640 4933 19674
rect 4899 19568 4933 19602
rect 4899 19496 4933 19530
rect 5058 19034 5092 19068
rect 5192 19034 5226 19068
rect 3552 17650 3586 17684
rect 3444 17565 3478 17599
rect 3444 17496 3478 17530
rect 3444 17427 3478 17461
rect 3444 17358 3478 17392
rect 3444 17289 3478 17323
rect 3444 17220 3478 17254
rect 3444 17151 3478 17185
rect 3552 17579 3586 17613
rect 3552 17508 3586 17542
rect 3552 17436 3586 17470
rect 3552 17364 3586 17398
rect 3552 17292 3586 17326
rect 3552 17220 3586 17254
rect 3552 17148 3586 17182
rect 3444 17081 3478 17115
rect 3444 17011 3478 17045
rect 3444 16941 3478 16975
rect 3444 16871 3478 16905
rect 3444 16801 3478 16835
rect 4285 16833 4319 16867
rect 4357 16833 4391 16867
rect 4429 16833 4463 16867
rect 4501 16833 4535 16867
rect 4573 16833 4607 16867
rect 4645 16833 4679 16867
rect 4716 16833 4750 16867
rect 4787 16833 4821 16867
rect 4909 16833 4943 16867
rect 4981 16833 5015 16867
rect 5053 16833 5087 16867
rect 5125 16833 5159 16867
rect 5197 16833 5231 16867
rect 5269 16833 5303 16867
rect 5340 16833 5374 16867
rect 5411 16833 5445 16867
rect 3444 16731 3478 16765
rect 3444 16661 3478 16695
rect 3444 16591 3478 16625
rect 3444 16521 3478 16555
rect 3444 16451 3478 16485
rect 3444 16381 3478 16415
rect 3444 16311 3478 16345
rect 3444 16241 3478 16275
rect 3444 16171 3478 16205
rect 3444 16101 3478 16135
rect 3444 16031 3478 16065
rect 4251 16061 4285 16095
rect 4320 16061 4354 16095
rect 4389 16061 4423 16095
rect 4458 16061 4492 16095
rect 4527 16061 4561 16095
rect 4596 16061 4630 16095
rect 4665 16061 4699 16095
rect 4735 16061 4769 16095
rect 4805 16061 4839 16095
rect 4875 16061 4909 16095
rect 4945 16061 4979 16095
rect 5015 16061 5049 16095
rect 5085 16061 5119 16095
rect 5155 16061 5189 16095
rect 5225 16061 5259 16095
rect 5295 16061 5329 16095
rect 5365 16061 5399 16095
rect 5435 16061 5469 16095
rect 5505 16061 5539 16095
rect 5575 16061 5609 16095
rect 5645 16061 5679 16095
rect 5715 16061 5749 16095
rect 5785 16061 5819 16095
rect 4251 15331 4285 15365
rect 4320 15331 4354 15365
rect 4389 15331 4423 15365
rect 4458 15331 4492 15365
rect 4527 15331 4561 15365
rect 4596 15331 4630 15365
rect 4665 15331 4699 15365
rect 4735 15331 4769 15365
rect 4805 15331 4839 15365
rect 4875 15331 4909 15365
rect 4945 15331 4979 15365
rect 5015 15331 5049 15365
rect 5085 15331 5119 15365
rect 5155 15331 5189 15365
rect 5225 15331 5259 15365
rect 5295 15331 5329 15365
rect 5365 15331 5399 15365
rect 5435 15331 5469 15365
rect 5505 15331 5539 15365
rect 5575 15331 5609 15365
rect 5645 15331 5679 15365
rect 5715 15331 5749 15365
rect 5785 15331 5819 15365
<< locali >>
rect 2816 39874 7786 39880
rect 2816 39840 2897 39874
rect 2952 39840 2972 39874
rect 3020 39840 3047 39874
rect 3088 39840 3122 39874
rect 3157 39840 3190 39874
rect 3233 39840 3258 39874
rect 3309 39840 3326 39874
rect 3385 39840 3394 39874
rect 3461 39840 3462 39874
rect 3496 39840 3503 39874
rect 3564 39840 3579 39874
rect 3632 39840 3655 39874
rect 3700 39840 3731 39874
rect 3768 39840 3802 39874
rect 3841 39840 3870 39874
rect 3917 39840 3938 39874
rect 3993 39840 4006 39874
rect 4069 39840 4074 39874
rect 4108 39840 4111 39874
rect 4176 39840 4210 39874
rect 4255 39840 4278 39874
rect 4328 39840 4346 39874
rect 4401 39840 4414 39874
rect 4474 39840 4482 39874
rect 4547 39840 4550 39874
rect 4584 39840 4586 39874
rect 4652 39840 4659 39874
rect 4720 39840 4732 39874
rect 4788 39840 4805 39874
rect 4856 39840 4878 39874
rect 4924 39840 4951 39874
rect 4992 39840 5024 39874
rect 5060 39840 5094 39874
rect 5131 39840 5162 39874
rect 5204 39840 5230 39874
rect 5277 39840 5298 39874
rect 5350 39840 5366 39874
rect 5423 39840 5434 39874
rect 5496 39840 5502 39874
rect 5569 39840 5570 39874
rect 5604 39840 5608 39874
rect 5672 39840 5681 39874
rect 5740 39840 5754 39874
rect 5808 39840 5827 39874
rect 5876 39840 5900 39874
rect 5944 39840 5973 39874
rect 6012 39840 6046 39874
rect 6080 39840 6114 39874
rect 6154 39840 6182 39874
rect 6228 39840 6250 39874
rect 6302 39840 6318 39874
rect 6376 39840 6386 39874
rect 6450 39840 6454 39874
rect 6488 39840 6490 39874
rect 6556 39840 6564 39874
rect 6624 39840 6638 39874
rect 6692 39840 6712 39874
rect 6760 39840 6786 39874
rect 6828 39840 6860 39874
rect 6896 39840 6930 39874
rect 6968 39840 6998 39874
rect 7042 39840 7066 39874
rect 7116 39840 7134 39874
rect 7190 39840 7202 39874
rect 7264 39840 7270 39874
rect 7372 39840 7378 39874
rect 7440 39840 7452 39874
rect 7508 39840 7526 39874
rect 7576 39840 7600 39874
rect 7644 39840 7674 39874
rect 7712 39840 7786 39874
rect 2816 39834 7786 39840
rect 2816 39806 2862 39834
rect 2816 39768 2822 39806
rect 2856 39768 2862 39806
rect 2816 39738 2862 39768
rect 2816 39695 2822 39738
rect 2856 39695 2862 39738
rect 2816 39670 2862 39695
rect 2816 39622 2822 39670
rect 2856 39622 2862 39670
rect 2816 39602 2862 39622
rect 7740 39802 7786 39834
rect 7740 39768 7746 39802
rect 7780 39768 7786 39802
rect 7740 39734 7786 39768
rect 7740 39696 7746 39734
rect 7780 39696 7786 39734
rect 7740 39666 7786 39696
rect 7740 39624 7746 39666
rect 7780 39624 7786 39666
rect 2816 39549 2822 39602
rect 2856 39549 2862 39602
rect 2816 39534 2862 39549
rect 2816 39476 2822 39534
rect 2856 39476 2862 39534
rect 2816 39466 2862 39476
rect 2816 39403 2822 39466
rect 2856 39403 2862 39466
rect 2816 39398 2862 39403
rect 2816 39296 2822 39398
rect 2856 39296 2862 39398
rect 2816 39291 2862 39296
rect 2816 39228 2822 39291
rect 2856 39228 2862 39291
rect 2816 39218 2862 39228
rect 2816 39160 2822 39218
rect 2856 39160 2862 39218
rect 2816 39145 2862 39160
rect 2816 39092 2822 39145
rect 2856 39092 2862 39145
rect 2816 39072 2862 39092
rect 2816 39024 2822 39072
rect 2856 39024 2862 39072
rect 2816 38999 2862 39024
rect 2816 38956 2822 38999
rect 2856 38956 2862 38999
rect 2816 38926 2862 38956
rect 2816 38888 2822 38926
rect 2856 38888 2862 38926
rect 2816 38854 2862 38888
rect 2816 38819 2822 38854
rect 2856 38819 2862 38854
rect 2816 38786 2862 38819
rect 2816 38746 2822 38786
rect 2856 38746 2862 38786
rect 2816 38718 2862 38746
rect 2816 38673 2822 38718
rect 2856 38673 2862 38718
rect 2816 38650 2862 38673
rect 2816 38600 2822 38650
rect 2856 38600 2862 38650
rect 2816 38582 2862 38600
rect 2816 38527 2822 38582
rect 2856 38527 2862 38582
rect 2816 38514 2862 38527
rect 2816 38454 2822 38514
rect 2856 38454 2862 38514
rect 2816 38446 2862 38454
rect 2816 38381 2822 38446
rect 2856 38381 2862 38446
rect 2816 38378 2862 38381
rect 2816 38344 2822 38378
rect 2856 38344 2862 38378
rect 2816 38342 2862 38344
rect 2816 38276 2822 38342
rect 2856 38276 2862 38342
rect 2816 38269 2862 38276
rect 2816 38208 2822 38269
rect 2856 38208 2862 38269
rect 2816 38196 2862 38208
rect 2816 38140 2822 38196
rect 2856 38140 2862 38196
rect 2816 38123 2862 38140
rect 2816 38072 2822 38123
rect 2856 38072 2862 38123
rect 2816 38050 2862 38072
rect 2816 38004 2822 38050
rect 2856 38004 2862 38050
rect 2816 37977 2862 38004
rect 2816 37936 2822 37977
rect 2856 37936 2862 37977
rect 2816 37904 2862 37936
rect 2816 37868 2822 37904
rect 2856 37868 2862 37904
rect 2816 37834 2862 37868
rect 2816 37797 2822 37834
rect 2856 37797 2862 37834
rect 2816 37766 2862 37797
rect 2816 37724 2822 37766
rect 2856 37724 2862 37766
rect 2816 37698 2862 37724
rect 2816 37651 2822 37698
rect 2856 37651 2862 37698
rect 2816 37630 2862 37651
rect 2816 37578 2822 37630
rect 2856 37578 2862 37630
rect 2816 37562 2862 37578
rect 2816 37505 2822 37562
rect 2856 37505 2862 37562
rect 2816 37494 2862 37505
rect 2816 37432 2822 37494
rect 2856 37432 2862 37494
rect 2816 37426 2862 37432
rect 2816 37359 2822 37426
rect 2856 37359 2862 37426
rect 2816 37358 2862 37359
rect 2816 37324 2822 37358
rect 2856 37324 2862 37358
rect 2816 37320 2862 37324
rect 2816 37256 2822 37320
rect 2856 37256 2862 37320
rect 2816 37247 2862 37256
rect 2816 37188 2822 37247
rect 2856 37188 2862 37247
rect 2816 37174 2862 37188
rect 2816 37120 2822 37174
rect 2856 37120 2862 37174
rect 2816 37102 2862 37120
rect 2816 37052 2822 37102
rect 2856 37052 2862 37102
rect 2816 37030 2862 37052
rect 2816 36984 2822 37030
rect 2856 36984 2862 37030
rect 2816 36958 2862 36984
rect 2816 36916 2822 36958
rect 2856 36916 2862 36958
rect 2816 36886 2862 36916
rect 2816 36848 2822 36886
rect 2856 36848 2862 36886
rect 2816 36814 2862 36848
rect 2816 36780 2822 36814
rect 2856 36780 2862 36814
rect 2816 36746 2862 36780
rect 2816 36708 2822 36746
rect 2856 36708 2862 36746
rect 2816 36678 2862 36708
rect 2816 36636 2822 36678
rect 2856 36636 2862 36678
rect 2816 36610 2862 36636
rect 2816 36564 2822 36610
rect 2856 36564 2862 36610
rect 2816 36542 2862 36564
rect 2816 36492 2822 36542
rect 2856 36492 2862 36542
rect 2816 36474 2862 36492
rect 2816 36420 2822 36474
rect 2856 36420 2862 36474
rect 2816 36406 2862 36420
rect 2816 36348 2822 36406
rect 2856 36348 2862 36406
rect 2816 36338 2862 36348
rect 2816 36276 2822 36338
rect 2856 36276 2862 36338
rect 2816 36270 2862 36276
rect 2816 36204 2822 36270
rect 2856 36204 2862 36270
rect 2816 36202 2862 36204
rect 2816 36168 2822 36202
rect 2856 36168 2862 36202
rect 2816 36166 2862 36168
rect 2816 36100 2822 36166
rect 2856 36100 2862 36166
rect 2816 36094 2862 36100
rect 2816 36032 2822 36094
rect 2856 36032 2862 36094
rect 2816 36022 2862 36032
rect 2816 35964 2822 36022
rect 2856 35964 2862 36022
rect 2816 35950 2862 35964
rect 2816 35896 2822 35950
rect 2856 35896 2862 35950
rect 2816 35878 2862 35896
rect 2816 35828 2822 35878
rect 2856 35828 2862 35878
rect 2816 35806 2862 35828
rect 2816 35760 2822 35806
rect 2856 35760 2862 35806
rect 2816 35734 2862 35760
rect 2816 35692 2822 35734
rect 2856 35692 2862 35734
rect 2816 35662 2862 35692
rect 2816 35624 2822 35662
rect 2856 35624 2862 35662
rect 2816 35590 2862 35624
rect 2816 35556 2822 35590
rect 2856 35556 2862 35590
rect 2816 35522 2862 35556
rect 2816 35484 2822 35522
rect 2856 35484 2862 35522
rect 2816 35454 2862 35484
rect 2816 35412 2822 35454
rect 2856 35412 2862 35454
rect 2816 35386 2862 35412
rect 2816 35340 2822 35386
rect 2856 35340 2862 35386
rect 2816 35318 2862 35340
rect 2816 35268 2822 35318
rect 2856 35268 2862 35318
rect 2816 35250 2862 35268
rect 2816 35196 2822 35250
rect 2856 35196 2862 35250
rect 2816 35182 2862 35196
rect 2816 35124 2822 35182
rect 2856 35124 2862 35182
rect 2816 35114 2862 35124
rect 2816 35052 2822 35114
rect 2856 35052 2862 35114
rect 2816 35046 2862 35052
rect 2816 34980 2822 35046
rect 2856 34980 2862 35046
rect 2816 34978 2862 34980
rect 2816 34944 2822 34978
rect 2856 34944 2862 34978
rect 2816 34942 2862 34944
rect 2816 34876 2822 34942
rect 2856 34876 2862 34942
rect 2816 34870 2862 34876
rect 2816 34808 2822 34870
rect 2856 34808 2862 34870
rect 2816 34798 2862 34808
rect 2816 34740 2822 34798
rect 2856 34740 2862 34798
rect 2816 34726 2862 34740
rect 2816 34672 2822 34726
rect 2856 34672 2862 34726
rect 2816 34654 2862 34672
rect 2816 34604 2822 34654
rect 2856 34604 2862 34654
rect 2816 34582 2862 34604
rect 2816 34536 2822 34582
rect 2856 34536 2862 34582
rect 2816 34510 2862 34536
rect 2816 34468 2822 34510
rect 2856 34468 2862 34510
rect 2816 34438 2862 34468
rect 2816 34400 2822 34438
rect 2856 34400 2862 34438
rect 2816 34366 2862 34400
rect 2816 34332 2822 34366
rect 2856 34332 2862 34366
rect 2816 34298 2862 34332
rect 2816 34260 2822 34298
rect 2856 34260 2862 34298
rect 2816 34230 2862 34260
rect 2816 34188 2822 34230
rect 2856 34188 2862 34230
rect 2816 34162 2862 34188
rect 2816 34116 2822 34162
rect 2856 34116 2862 34162
rect 2816 34094 2862 34116
rect 2816 34044 2822 34094
rect 2856 34044 2862 34094
rect 2816 34026 2862 34044
rect 2816 33972 2822 34026
rect 2856 33972 2862 34026
rect 2816 33958 2862 33972
rect 2816 33900 2822 33958
rect 2856 33900 2862 33958
rect 2816 33890 2862 33900
rect 2816 33828 2822 33890
rect 2856 33828 2862 33890
rect 2816 33822 2862 33828
rect 2816 33756 2822 33822
rect 2856 33756 2862 33822
rect 2816 33754 2862 33756
rect 2816 33720 2822 33754
rect 2856 33720 2862 33754
rect 2816 33718 2862 33720
rect 2816 33652 2822 33718
rect 2856 33652 2862 33718
rect 2816 33646 2862 33652
rect 2816 33584 2822 33646
rect 2856 33584 2862 33646
rect 2816 33574 2862 33584
rect 2816 33516 2822 33574
rect 2856 33516 2862 33574
rect 2816 33502 2862 33516
rect 2816 33448 2822 33502
rect 2856 33448 2862 33502
rect 2816 33430 2862 33448
rect 2816 33380 2822 33430
rect 2856 33380 2862 33430
rect 2816 33358 2862 33380
rect 2816 33312 2822 33358
rect 2856 33312 2862 33358
rect 2816 33286 2862 33312
rect 2816 33244 2822 33286
rect 2856 33244 2862 33286
rect 2816 33214 2862 33244
rect 2816 33176 2822 33214
rect 2856 33176 2862 33214
rect 2816 33142 2862 33176
rect 2816 33108 2822 33142
rect 2856 33108 2862 33142
rect 2816 33074 2862 33108
rect 2816 33036 2822 33074
rect 2856 33036 2862 33074
rect 2816 33006 2862 33036
rect 2816 32964 2822 33006
rect 2856 32964 2862 33006
rect 2816 32938 2862 32964
rect 2816 32892 2822 32938
rect 2856 32892 2862 32938
rect 2816 32870 2862 32892
rect 2816 32820 2822 32870
rect 2856 32820 2862 32870
rect 2816 32802 2862 32820
rect 2816 32748 2822 32802
rect 2856 32748 2862 32802
rect 2816 32734 2862 32748
rect 2816 32676 2822 32734
rect 2856 32676 2862 32734
rect 2816 32666 2862 32676
rect 2816 32604 2822 32666
rect 2856 32604 2862 32666
rect 2816 32598 2862 32604
rect 2816 32532 2822 32598
rect 2856 32532 2862 32598
rect 2816 32530 2862 32532
rect 2816 32496 2822 32530
rect 2856 32496 2862 32530
rect 2816 32494 2862 32496
rect 2816 32428 2822 32494
rect 2856 32428 2862 32494
rect 2816 32422 2862 32428
rect 2816 32360 2822 32422
rect 2856 32360 2862 32422
rect 2816 32350 2862 32360
rect 2816 32292 2822 32350
rect 2856 32292 2862 32350
rect 2816 32278 2862 32292
rect 2816 32224 2822 32278
rect 2856 32224 2862 32278
rect 2816 32206 2862 32224
rect 2816 32156 2822 32206
rect 2856 32156 2862 32206
rect 2816 32134 2862 32156
rect 2816 32088 2822 32134
rect 2856 32088 2862 32134
rect 2816 32062 2862 32088
rect 2816 32020 2822 32062
rect 2856 32020 2862 32062
rect 2816 31990 2862 32020
rect 2816 31952 2822 31990
rect 2856 31952 2862 31990
rect 2816 31918 2862 31952
rect 2816 31884 2822 31918
rect 2856 31884 2862 31918
rect 2816 31850 2862 31884
rect 2816 31812 2822 31850
rect 2856 31812 2862 31850
rect 2816 31782 2862 31812
rect 2816 31740 2822 31782
rect 2856 31740 2862 31782
rect 2816 31714 2862 31740
rect 2816 31668 2822 31714
rect 2856 31668 2862 31714
rect 2816 31646 2862 31668
rect 2816 31596 2822 31646
rect 2856 31596 2862 31646
rect 2816 31578 2862 31596
rect 2816 31524 2822 31578
rect 2856 31524 2862 31578
rect 2816 31510 2862 31524
rect 2816 31452 2822 31510
rect 2856 31452 2862 31510
rect 2816 31442 2862 31452
rect 2816 31380 2822 31442
rect 2856 31380 2862 31442
rect 2816 31374 2862 31380
rect 2816 31308 2822 31374
rect 2856 31308 2862 31374
rect 2816 31306 2862 31308
rect 2816 31272 2822 31306
rect 2856 31272 2862 31306
rect 2816 31270 2862 31272
rect 2816 31204 2822 31270
rect 2856 31204 2862 31270
rect 2816 31198 2862 31204
rect 2816 31136 2822 31198
rect 2856 31136 2862 31198
rect 2816 31126 2862 31136
rect 2816 31068 2822 31126
rect 2856 31068 2862 31126
rect 2816 31054 2862 31068
rect 2816 31000 2822 31054
rect 2856 31000 2862 31054
rect 2816 30982 2862 31000
rect 2816 30932 2822 30982
rect 2856 30932 2862 30982
rect 2816 30910 2862 30932
rect 2816 30864 2822 30910
rect 2856 30864 2862 30910
rect 2816 30838 2862 30864
rect 2816 30796 2822 30838
rect 2856 30796 2862 30838
rect 2816 30766 2862 30796
rect 2816 30728 2822 30766
rect 2856 30728 2862 30766
rect 2816 30694 2862 30728
rect 2816 30660 2822 30694
rect 2856 30660 2862 30694
rect 2816 30626 2862 30660
rect 2816 30588 2822 30626
rect 2856 30588 2862 30626
rect 2816 30558 2862 30588
rect 2816 30516 2822 30558
rect 2856 30516 2862 30558
rect 2816 30490 2862 30516
rect 2816 30444 2822 30490
rect 2856 30444 2862 30490
rect 2816 30422 2862 30444
rect 2816 30372 2822 30422
rect 2856 30372 2862 30422
rect 2816 30354 2862 30372
rect 2816 30300 2822 30354
rect 2856 30300 2862 30354
rect 2816 30286 2862 30300
rect 2816 30228 2822 30286
rect 2856 30228 2862 30286
rect 2816 30218 2862 30228
rect 2816 30156 2822 30218
rect 2856 30156 2862 30218
rect 2816 30150 2862 30156
rect 2816 30084 2822 30150
rect 2856 30084 2862 30150
rect 2816 30082 2862 30084
rect 2816 30048 2822 30082
rect 2856 30048 2862 30082
rect 2816 30046 2862 30048
rect 2816 29980 2822 30046
rect 2856 29980 2862 30046
rect 2816 29974 2862 29980
rect 2816 29912 2822 29974
rect 2856 29912 2862 29974
rect 2816 29902 2862 29912
rect 2816 29844 2822 29902
rect 2856 29844 2862 29902
rect 2816 29830 2862 29844
rect 2816 29776 2822 29830
rect 2856 29776 2862 29830
rect 2816 29758 2862 29776
rect 2816 29708 2822 29758
rect 2856 29708 2862 29758
rect 2816 29686 2862 29708
rect 2816 29640 2822 29686
rect 2856 29640 2862 29686
rect 2816 29614 2862 29640
rect 2816 29572 2822 29614
rect 2856 29572 2862 29614
rect 2816 29542 2862 29572
rect 2816 29504 2822 29542
rect 2856 29504 2862 29542
rect 2816 29470 2862 29504
rect 2816 29436 2822 29470
rect 2856 29436 2862 29470
rect 2816 29402 2862 29436
rect 2816 29364 2822 29402
rect 2856 29364 2862 29402
rect 2816 29334 2862 29364
rect 2816 29292 2822 29334
rect 2856 29292 2862 29334
rect 2816 29266 2862 29292
rect 2816 29220 2822 29266
rect 2856 29220 2862 29266
rect 2816 29198 2862 29220
rect 2816 29148 2822 29198
rect 2856 29148 2862 29198
rect 2816 29130 2862 29148
rect 2816 29076 2822 29130
rect 2856 29076 2862 29130
rect 2816 29062 2862 29076
rect 2816 29004 2822 29062
rect 2856 29004 2862 29062
rect 2816 28994 2862 29004
rect 2816 28932 2822 28994
rect 2856 28932 2862 28994
rect 2816 28926 2862 28932
rect 2816 28860 2822 28926
rect 2856 28860 2862 28926
rect 2816 28858 2862 28860
rect 2816 28824 2822 28858
rect 2856 28824 2862 28858
rect 2816 28822 2862 28824
rect 2816 28756 2822 28822
rect 2856 28756 2862 28822
rect 2816 28750 2862 28756
rect 2816 28688 2822 28750
rect 2856 28688 2862 28750
rect 2816 28678 2862 28688
rect 2816 28620 2822 28678
rect 2856 28620 2862 28678
rect 2816 28606 2862 28620
rect 2816 28552 2822 28606
rect 2856 28552 2862 28606
rect 2816 28534 2862 28552
rect 2816 28484 2822 28534
rect 2856 28484 2862 28534
rect 2816 28462 2862 28484
rect 2816 28416 2822 28462
rect 2856 28416 2862 28462
rect 2816 28390 2862 28416
rect 3076 39614 5370 39620
rect 3076 39580 3154 39614
rect 3191 39580 3222 39614
rect 3266 39580 3290 39614
rect 3341 39580 3358 39614
rect 3416 39580 3426 39614
rect 3491 39580 3494 39614
rect 3528 39580 3532 39614
rect 3596 39580 3607 39614
rect 3664 39580 3682 39614
rect 3732 39580 3757 39614
rect 3800 39580 3832 39614
rect 3868 39580 3902 39614
rect 3941 39580 3970 39614
rect 4016 39580 4038 39614
rect 4091 39580 4106 39614
rect 4166 39580 4174 39614
rect 4241 39580 4242 39614
rect 4276 39580 4282 39614
rect 4344 39580 4357 39614
rect 4412 39580 4433 39614
rect 4480 39580 4509 39614
rect 4548 39580 4582 39614
rect 4616 39580 4619 39614
rect 4684 39580 4698 39614
rect 4752 39580 4778 39614
rect 4820 39580 4854 39614
rect 4892 39580 4922 39614
rect 4972 39580 4990 39614
rect 5052 39580 5058 39614
rect 5092 39580 5098 39614
rect 5160 39580 5178 39614
rect 5228 39580 5258 39614
rect 5296 39580 5370 39614
rect 3076 39574 5370 39580
rect 3076 39546 3122 39574
rect 3076 39508 3082 39546
rect 3116 39508 3122 39546
rect 3076 39478 3122 39508
rect 3076 39435 3082 39478
rect 3116 39435 3122 39478
rect 5324 39542 5370 39574
rect 5324 39474 5330 39542
rect 5364 39474 5370 39542
rect 5324 39470 5370 39474
rect 3076 39410 3122 39435
rect 3076 39362 3082 39410
rect 3116 39362 3122 39410
rect 3076 39342 3122 39362
rect 3076 39289 3082 39342
rect 3116 39289 3122 39342
rect 3076 39274 3122 39289
rect 3076 39216 3082 39274
rect 3116 39216 3122 39274
rect 3076 39206 3122 39216
rect 3076 39143 3082 39206
rect 3116 39143 3122 39206
rect 3076 39138 3122 39143
rect 3076 39036 3082 39138
rect 3116 39036 3122 39138
rect 3076 39031 3122 39036
rect 3076 38968 3082 39031
rect 3116 38968 3122 39031
rect 3076 38958 3122 38968
rect 3076 38900 3082 38958
rect 3116 38900 3122 38958
rect 3076 38885 3122 38900
rect 3076 38832 3082 38885
rect 3116 38832 3122 38885
rect 3076 38812 3122 38832
rect 3076 38764 3082 38812
rect 3116 38764 3122 38812
rect 3076 38739 3122 38764
rect 3076 38696 3082 38739
rect 3116 38696 3122 38739
rect 3076 38666 3122 38696
rect 3076 38628 3082 38666
rect 3116 38628 3122 38666
rect 3076 38594 3122 38628
rect 3076 38559 3082 38594
rect 3116 38559 3122 38594
rect 3076 38526 3122 38559
rect 3076 38486 3082 38526
rect 3116 38486 3122 38526
rect 3076 38458 3122 38486
rect 3076 38413 3082 38458
rect 3116 38413 3122 38458
rect 3076 38390 3122 38413
rect 3076 38340 3082 38390
rect 3116 38340 3122 38390
rect 3076 38322 3122 38340
rect 3076 38267 3082 38322
rect 3116 38267 3122 38322
rect 3076 38254 3122 38267
rect 3076 38194 3082 38254
rect 3116 38194 3122 38254
rect 3076 38186 3122 38194
rect 3076 38121 3082 38186
rect 3116 38121 3122 38186
rect 3076 38118 3122 38121
rect 3076 38084 3082 38118
rect 3116 38084 3122 38118
rect 3076 38082 3122 38084
rect 3076 38016 3082 38082
rect 3116 38016 3122 38082
rect 3076 38010 3122 38016
rect 3076 37948 3082 38010
rect 3116 37948 3122 38010
rect 3076 37938 3122 37948
rect 3076 37880 3082 37938
rect 3116 37880 3122 37938
rect 3076 37866 3122 37880
rect 3076 37812 3082 37866
rect 3116 37812 3122 37866
rect 3076 37794 3122 37812
rect 3076 37744 3082 37794
rect 3116 37744 3122 37794
rect 3076 37722 3122 37744
rect 3076 37676 3082 37722
rect 3116 37676 3122 37722
rect 3076 37650 3122 37676
rect 3076 37608 3082 37650
rect 3116 37608 3122 37650
rect 3076 37578 3122 37608
rect 3076 37540 3082 37578
rect 3116 37540 3122 37578
rect 3076 37506 3122 37540
rect 3076 37472 3082 37506
rect 3116 37472 3122 37506
rect 3076 37438 3122 37472
rect 3076 37400 3082 37438
rect 3116 37400 3122 37438
rect 3076 37370 3122 37400
rect 3076 37328 3082 37370
rect 3116 37328 3122 37370
rect 3076 37302 3122 37328
rect 3076 37256 3082 37302
rect 3116 37256 3122 37302
rect 3076 37234 3122 37256
rect 3076 37184 3082 37234
rect 3116 37184 3122 37234
rect 3076 37166 3122 37184
rect 3076 37112 3082 37166
rect 3116 37112 3122 37166
rect 3076 37098 3122 37112
rect 3076 37040 3082 37098
rect 3116 37040 3122 37098
rect 3076 37030 3122 37040
rect 3076 36968 3082 37030
rect 3116 36968 3122 37030
rect 3076 36962 3122 36968
rect 3076 36896 3082 36962
rect 3116 36896 3122 36962
rect 3076 36894 3122 36896
rect 3076 36860 3082 36894
rect 3116 36860 3122 36894
rect 3076 36858 3122 36860
rect 3076 36792 3082 36858
rect 3116 36792 3122 36858
rect 3076 36786 3122 36792
rect 3076 36724 3082 36786
rect 3116 36724 3122 36786
rect 3076 36714 3122 36724
rect 3076 36656 3082 36714
rect 3116 36656 3122 36714
rect 3076 36642 3122 36656
rect 3076 36588 3082 36642
rect 3116 36588 3122 36642
rect 3076 36570 3122 36588
rect 3076 36520 3082 36570
rect 3116 36520 3122 36570
rect 3076 36498 3122 36520
rect 3076 36452 3082 36498
rect 3116 36452 3122 36498
rect 3076 36426 3122 36452
rect 3076 36384 3082 36426
rect 3116 36384 3122 36426
rect 3076 36354 3122 36384
rect 3076 36316 3082 36354
rect 3116 36316 3122 36354
rect 3076 36282 3122 36316
rect 3076 36248 3082 36282
rect 3116 36248 3122 36282
rect 3076 36214 3122 36248
rect 3076 36176 3082 36214
rect 3116 36176 3122 36214
rect 3076 36146 3122 36176
rect 3076 36104 3082 36146
rect 3116 36104 3122 36146
rect 3076 36078 3122 36104
rect 3076 36032 3082 36078
rect 3116 36032 3122 36078
rect 3076 36010 3122 36032
rect 3076 35960 3082 36010
rect 3116 35960 3122 36010
rect 3076 35942 3122 35960
rect 3076 35888 3082 35942
rect 3116 35888 3122 35942
rect 3076 35874 3122 35888
rect 3076 35816 3082 35874
rect 3116 35816 3122 35874
rect 3076 35806 3122 35816
rect 3076 35744 3082 35806
rect 3116 35744 3122 35806
rect 3076 35738 3122 35744
rect 3076 35672 3082 35738
rect 3116 35672 3122 35738
rect 3076 35670 3122 35672
rect 3076 35636 3082 35670
rect 3116 35636 3122 35670
rect 3076 35634 3122 35636
rect 3076 35568 3082 35634
rect 3116 35568 3122 35634
rect 3076 35562 3122 35568
rect 3076 35500 3082 35562
rect 3116 35500 3122 35562
rect 3076 35490 3122 35500
rect 3076 35432 3082 35490
rect 3116 35432 3122 35490
rect 3076 35418 3122 35432
rect 3076 35364 3082 35418
rect 3116 35364 3122 35418
rect 3076 35346 3122 35364
rect 3076 35296 3082 35346
rect 3116 35296 3122 35346
rect 3076 35274 3122 35296
rect 3076 35228 3082 35274
rect 3116 35228 3122 35274
rect 3076 35202 3122 35228
rect 3076 35160 3082 35202
rect 3116 35160 3122 35202
rect 3076 35130 3122 35160
rect 3076 35092 3082 35130
rect 3116 35092 3122 35130
rect 3076 35058 3122 35092
rect 3076 35024 3082 35058
rect 3116 35024 3122 35058
rect 3076 34990 3122 35024
rect 3076 34952 3082 34990
rect 3116 34952 3122 34990
rect 3076 34922 3122 34952
rect 3076 34880 3082 34922
rect 3116 34880 3122 34922
rect 3076 34854 3122 34880
rect 3076 34808 3082 34854
rect 3116 34808 3122 34854
rect 3076 34786 3122 34808
rect 3076 34736 3082 34786
rect 3116 34736 3122 34786
rect 3076 34718 3122 34736
rect 3076 34664 3082 34718
rect 3116 34664 3122 34718
rect 3076 34650 3122 34664
rect 3076 34592 3082 34650
rect 3116 34592 3122 34650
rect 3076 34582 3122 34592
rect 3076 34520 3082 34582
rect 3116 34520 3122 34582
rect 3076 34514 3122 34520
rect 3076 34448 3082 34514
rect 3116 34448 3122 34514
rect 3076 34446 3122 34448
rect 3076 34412 3082 34446
rect 3116 34412 3122 34446
rect 3076 34410 3122 34412
rect 3076 34344 3082 34410
rect 3116 34344 3122 34410
rect 3076 34338 3122 34344
rect 3076 34276 3082 34338
rect 3116 34276 3122 34338
rect 3076 34266 3122 34276
rect 3076 34208 3082 34266
rect 3116 34208 3122 34266
rect 3076 34194 3122 34208
rect 3076 34140 3082 34194
rect 3116 34140 3122 34194
rect 3076 34122 3122 34140
rect 3076 34072 3082 34122
rect 3116 34072 3122 34122
rect 3076 34050 3122 34072
rect 3076 34004 3082 34050
rect 3116 34004 3122 34050
rect 3076 33978 3122 34004
rect 3076 33936 3082 33978
rect 3116 33936 3122 33978
rect 3076 33906 3122 33936
rect 3076 33868 3082 33906
rect 3116 33868 3122 33906
rect 3076 33834 3122 33868
rect 3076 33800 3082 33834
rect 3116 33800 3122 33834
rect 3076 33766 3122 33800
rect 3076 33728 3082 33766
rect 3116 33728 3122 33766
rect 3076 33698 3122 33728
rect 3076 33656 3082 33698
rect 3116 33656 3122 33698
rect 3076 33630 3122 33656
rect 3076 33584 3082 33630
rect 3116 33584 3122 33630
rect 3076 33562 3122 33584
rect 3076 33512 3082 33562
rect 3116 33512 3122 33562
rect 3076 33494 3122 33512
rect 3076 33440 3082 33494
rect 3116 33440 3122 33494
rect 3076 33426 3122 33440
rect 3076 33368 3082 33426
rect 3116 33368 3122 33426
rect 3076 33358 3122 33368
rect 3076 33296 3082 33358
rect 3116 33296 3122 33358
rect 3076 33290 3122 33296
rect 3076 33224 3082 33290
rect 3116 33224 3122 33290
rect 3076 33222 3122 33224
rect 3076 33188 3082 33222
rect 3116 33188 3122 33222
rect 3076 33186 3122 33188
rect 3076 33120 3082 33186
rect 3116 33120 3122 33186
rect 3076 33114 3122 33120
rect 3076 33052 3082 33114
rect 3116 33052 3122 33114
rect 3076 33042 3122 33052
rect 3076 32984 3082 33042
rect 3116 32984 3122 33042
rect 3076 32970 3122 32984
rect 3076 32916 3082 32970
rect 3116 32916 3122 32970
rect 3076 32898 3122 32916
rect 3076 32848 3082 32898
rect 3116 32848 3122 32898
rect 3076 32826 3122 32848
rect 3076 32780 3082 32826
rect 3116 32780 3122 32826
rect 3076 32754 3122 32780
rect 3076 32712 3082 32754
rect 3116 32712 3122 32754
rect 3076 32682 3122 32712
rect 3076 32644 3082 32682
rect 3116 32644 3122 32682
rect 3076 32610 3122 32644
rect 3076 32576 3082 32610
rect 3116 32576 3122 32610
rect 3076 32542 3122 32576
rect 3076 32504 3082 32542
rect 3116 32504 3122 32542
rect 3076 32474 3122 32504
rect 3076 32432 3082 32474
rect 3116 32432 3122 32474
rect 3076 32406 3122 32432
rect 3076 32360 3082 32406
rect 3116 32360 3122 32406
rect 3076 32338 3122 32360
rect 3076 32288 3082 32338
rect 3116 32288 3122 32338
rect 3076 32270 3122 32288
rect 3076 32216 3082 32270
rect 3116 32216 3122 32270
rect 3076 32202 3122 32216
rect 3076 32144 3082 32202
rect 3116 32144 3122 32202
rect 3076 32134 3122 32144
rect 3076 32072 3082 32134
rect 3116 32072 3122 32134
rect 3076 32066 3122 32072
rect 3076 32000 3082 32066
rect 3116 32000 3122 32066
rect 3076 31998 3122 32000
rect 3076 31964 3082 31998
rect 3116 31964 3122 31998
rect 3076 31962 3122 31964
rect 3076 31896 3082 31962
rect 3116 31896 3122 31962
rect 3076 31890 3122 31896
rect 3076 31828 3082 31890
rect 3116 31828 3122 31890
rect 3076 31818 3122 31828
rect 3076 31760 3082 31818
rect 3116 31760 3122 31818
rect 3076 31746 3122 31760
rect 3076 31692 3082 31746
rect 3116 31692 3122 31746
rect 3076 31674 3122 31692
rect 3076 31624 3082 31674
rect 3116 31624 3122 31674
rect 3076 31602 3122 31624
rect 3076 31556 3082 31602
rect 3116 31556 3122 31602
rect 3076 31530 3122 31556
rect 3076 31488 3082 31530
rect 3116 31488 3122 31530
rect 3076 31458 3122 31488
rect 3076 31420 3082 31458
rect 3116 31420 3122 31458
rect 3076 31386 3122 31420
rect 3076 31352 3082 31386
rect 3116 31352 3122 31386
rect 3076 31318 3122 31352
rect 3076 31280 3082 31318
rect 3116 31280 3122 31318
rect 3076 31250 3122 31280
rect 3076 31208 3082 31250
rect 3116 31208 3122 31250
rect 3076 31182 3122 31208
rect 3076 31136 3082 31182
rect 3116 31136 3122 31182
rect 3076 31114 3122 31136
rect 3076 31064 3082 31114
rect 3116 31064 3122 31114
rect 3076 31046 3122 31064
rect 3076 30992 3082 31046
rect 3116 30992 3122 31046
rect 3076 30978 3122 30992
rect 3076 30920 3082 30978
rect 3116 30920 3122 30978
rect 3076 30910 3122 30920
rect 3076 30848 3082 30910
rect 3116 30848 3122 30910
rect 3076 30842 3122 30848
rect 3076 30776 3082 30842
rect 3116 30776 3122 30842
rect 3076 30774 3122 30776
rect 3076 30740 3082 30774
rect 3116 30740 3122 30774
rect 3076 30738 3122 30740
rect 3076 30672 3082 30738
rect 3116 30672 3122 30738
rect 3076 30666 3122 30672
rect 3076 30604 3082 30666
rect 3116 30604 3122 30666
rect 3076 30594 3122 30604
rect 3076 30536 3082 30594
rect 3116 30536 3122 30594
rect 3076 30522 3122 30536
rect 3076 30468 3082 30522
rect 3116 30468 3122 30522
rect 3076 30450 3122 30468
rect 3076 30400 3082 30450
rect 3116 30400 3122 30450
rect 3076 30378 3122 30400
rect 3174 39431 3208 39447
rect 3174 39363 3208 39397
rect 3174 39295 3208 39319
rect 3174 39227 3208 39247
rect 3174 39159 3208 39175
rect 3174 39091 3208 39103
rect 3174 39023 3208 39031
rect 3174 38955 3208 38959
rect 3174 38849 3208 38853
rect 3174 38777 3208 38785
rect 3174 38705 3208 38717
rect 3174 38633 3208 38649
rect 3174 38561 3208 38581
rect 3174 38489 3208 38513
rect 3174 38417 3208 38445
rect 3174 38345 3208 38377
rect 3174 38275 3208 38309
rect 3174 38207 3208 38239
rect 3174 38139 3208 38167
rect 3174 38071 3208 38095
rect 3174 38003 3208 38023
rect 3174 37935 3208 37951
rect 3174 37867 3208 37879
rect 3174 37799 3208 37807
rect 3174 37731 3208 37735
rect 3174 37625 3208 37629
rect 3174 37553 3208 37561
rect 3174 37481 3208 37493
rect 3174 37409 3208 37425
rect 3174 37337 3208 37357
rect 3174 37265 3208 37289
rect 3174 37193 3208 37221
rect 3174 37121 3208 37153
rect 3174 37051 3208 37085
rect 3174 36983 3208 37015
rect 3174 36915 3208 36943
rect 3174 36847 3208 36871
rect 3174 36779 3208 36799
rect 3174 36711 3208 36727
rect 3174 36643 3208 36655
rect 3174 36575 3208 36583
rect 3174 36507 3208 36511
rect 3174 36401 3208 36405
rect 3174 36329 3208 36337
rect 3174 36257 3208 36269
rect 3174 36185 3208 36201
rect 3174 36113 3208 36133
rect 3174 36041 3208 36065
rect 3174 35969 3208 35997
rect 3174 35897 3208 35929
rect 3174 35827 3208 35861
rect 3174 35759 3208 35791
rect 3174 35691 3208 35719
rect 3174 35623 3208 35647
rect 3174 35555 3208 35575
rect 3174 35487 3208 35503
rect 3174 35419 3208 35431
rect 3174 35351 3208 35359
rect 3174 35283 3208 35287
rect 3174 35177 3208 35181
rect 3174 35105 3208 35113
rect 3174 35033 3208 35045
rect 3174 34961 3208 34977
rect 3174 34889 3208 34909
rect 3174 34817 3208 34841
rect 3174 34745 3208 34773
rect 3174 34673 3208 34705
rect 3174 34603 3208 34637
rect 3174 34535 3208 34567
rect 3174 34467 3208 34495
rect 3174 34399 3208 34423
rect 3174 34331 3208 34351
rect 3174 34263 3208 34279
rect 3174 34195 3208 34207
rect 3174 34127 3208 34135
rect 3174 34059 3208 34063
rect 3174 33953 3208 33957
rect 3174 33881 3208 33889
rect 3174 33809 3208 33821
rect 3174 33737 3208 33753
rect 3174 33665 3208 33685
rect 3174 33593 3208 33617
rect 3174 33521 3208 33549
rect 3174 33449 3208 33481
rect 3174 33379 3208 33413
rect 3174 33311 3208 33343
rect 3174 33243 3208 33271
rect 3174 33175 3208 33199
rect 3174 33107 3208 33127
rect 3174 33039 3208 33055
rect 3174 32971 3208 32983
rect 3174 32903 3208 32911
rect 3174 32835 3208 32839
rect 3174 32729 3208 32733
rect 3174 32657 3208 32665
rect 3174 32585 3208 32597
rect 3174 32513 3208 32529
rect 3174 32441 3208 32461
rect 3174 32369 3208 32393
rect 3174 32296 3208 32325
rect 3174 32223 3208 32257
rect 3174 32155 3208 32189
rect 3174 32087 3208 32116
rect 3174 32019 3208 32043
rect 3174 31951 3208 31970
rect 3174 31882 3208 31897
rect 3174 31813 3208 31824
rect 3174 31744 3208 31751
rect 3174 31675 3208 31678
rect 3174 31639 3208 31641
rect 3174 31566 3208 31572
rect 3174 31493 3208 31503
rect 3174 31420 3208 31434
rect 3174 31347 3208 31365
rect 3174 31274 3208 31296
rect 3174 31201 3208 31227
rect 3174 31128 3208 31158
rect 3174 31055 3208 31089
rect 3174 30985 3208 31020
rect 3174 30916 3208 30948
rect 3174 30847 3208 30875
rect 3174 30778 3208 30802
rect 3174 30709 3208 30729
rect 3174 30640 3208 30656
rect 3174 30571 3208 30583
rect 3174 30502 3208 30510
rect 3174 30433 3208 30437
rect 3174 30383 3208 30399
rect 5324 39406 5330 39470
rect 5364 39406 5370 39470
rect 5324 39398 5370 39406
rect 5324 39338 5330 39398
rect 5364 39338 5370 39398
rect 5324 39326 5370 39338
rect 5324 39270 5330 39326
rect 5364 39270 5370 39326
rect 5324 39254 5370 39270
rect 5324 39202 5330 39254
rect 5364 39202 5370 39254
rect 5324 39182 5370 39202
rect 5324 39134 5330 39182
rect 5364 39134 5370 39182
rect 5324 39110 5370 39134
rect 5324 39066 5330 39110
rect 5364 39066 5370 39110
rect 5324 39038 5370 39066
rect 5324 38998 5330 39038
rect 5364 38998 5370 39038
rect 5324 38966 5370 38998
rect 5324 38930 5330 38966
rect 5364 38930 5370 38966
rect 5324 38896 5370 38930
rect 5324 38860 5330 38896
rect 5364 38860 5370 38896
rect 5324 38828 5370 38860
rect 5324 38788 5330 38828
rect 5364 38788 5370 38828
rect 5324 38760 5370 38788
rect 5324 38716 5330 38760
rect 5364 38716 5370 38760
rect 5324 38692 5370 38716
rect 5324 38644 5330 38692
rect 5364 38644 5370 38692
rect 5324 38624 5370 38644
rect 5324 38572 5330 38624
rect 5364 38572 5370 38624
rect 5324 38556 5370 38572
rect 5324 38500 5330 38556
rect 5364 38500 5370 38556
rect 5324 38488 5370 38500
rect 5324 38428 5330 38488
rect 5364 38428 5370 38488
rect 5324 38420 5370 38428
rect 5324 38356 5330 38420
rect 5364 38356 5370 38420
rect 5324 38352 5370 38356
rect 5324 38250 5330 38352
rect 5364 38250 5370 38352
rect 5324 38246 5370 38250
rect 5324 38182 5330 38246
rect 5364 38182 5370 38246
rect 5324 38174 5370 38182
rect 5324 38114 5330 38174
rect 5364 38114 5370 38174
rect 5324 38102 5370 38114
rect 5324 38046 5330 38102
rect 5364 38046 5370 38102
rect 5324 38030 5370 38046
rect 5324 37978 5330 38030
rect 5364 37978 5370 38030
rect 5324 37958 5370 37978
rect 5324 37910 5330 37958
rect 5364 37910 5370 37958
rect 5324 37886 5370 37910
rect 5324 37842 5330 37886
rect 5364 37842 5370 37886
rect 5324 37814 5370 37842
rect 5324 37774 5330 37814
rect 5364 37774 5370 37814
rect 5324 37742 5370 37774
rect 5324 37706 5330 37742
rect 5364 37706 5370 37742
rect 5324 37672 5370 37706
rect 5324 37636 5330 37672
rect 5364 37636 5370 37672
rect 5324 37604 5370 37636
rect 5324 37564 5330 37604
rect 5364 37564 5370 37604
rect 5324 37536 5370 37564
rect 5324 37492 5330 37536
rect 5364 37492 5370 37536
rect 5324 37468 5370 37492
rect 5324 37420 5330 37468
rect 5364 37420 5370 37468
rect 5324 37400 5370 37420
rect 5324 37348 5330 37400
rect 5364 37348 5370 37400
rect 5324 37332 5370 37348
rect 5324 37276 5330 37332
rect 5364 37276 5370 37332
rect 5324 37264 5370 37276
rect 5324 37204 5330 37264
rect 5364 37204 5370 37264
rect 5324 37196 5370 37204
rect 5324 37132 5330 37196
rect 5364 37132 5370 37196
rect 5324 37128 5370 37132
rect 5324 37026 5330 37128
rect 5364 37026 5370 37128
rect 5324 37022 5370 37026
rect 5324 36958 5330 37022
rect 5364 36958 5370 37022
rect 5324 36950 5370 36958
rect 5324 36890 5330 36950
rect 5364 36890 5370 36950
rect 5324 36878 5370 36890
rect 5324 36822 5330 36878
rect 5364 36822 5370 36878
rect 5324 36806 5370 36822
rect 5324 36754 5330 36806
rect 5364 36754 5370 36806
rect 5324 36734 5370 36754
rect 5324 36686 5330 36734
rect 5364 36686 5370 36734
rect 5324 36662 5370 36686
rect 5324 36618 5330 36662
rect 5364 36618 5370 36662
rect 5324 36590 5370 36618
rect 5324 36550 5330 36590
rect 5364 36550 5370 36590
rect 5324 36518 5370 36550
rect 5324 36482 5330 36518
rect 5364 36482 5370 36518
rect 5324 36448 5370 36482
rect 5324 36412 5330 36448
rect 5364 36412 5370 36448
rect 5324 36380 5370 36412
rect 5324 36340 5330 36380
rect 5364 36340 5370 36380
rect 5324 36312 5370 36340
rect 5324 36268 5330 36312
rect 5364 36268 5370 36312
rect 5324 36244 5370 36268
rect 5324 36196 5330 36244
rect 5364 36196 5370 36244
rect 5324 36176 5370 36196
rect 5324 36124 5330 36176
rect 5364 36124 5370 36176
rect 5324 36108 5370 36124
rect 5324 36052 5330 36108
rect 5364 36052 5370 36108
rect 5324 36040 5370 36052
rect 5324 35980 5330 36040
rect 5364 35980 5370 36040
rect 5324 35972 5370 35980
rect 5324 35908 5330 35972
rect 5364 35908 5370 35972
rect 5324 35904 5370 35908
rect 5324 35802 5330 35904
rect 5364 35802 5370 35904
rect 5324 35798 5370 35802
rect 5324 35734 5330 35798
rect 5364 35734 5370 35798
rect 5324 35726 5370 35734
rect 5324 35666 5330 35726
rect 5364 35666 5370 35726
rect 5324 35654 5370 35666
rect 5324 35598 5330 35654
rect 5364 35598 5370 35654
rect 5324 35582 5370 35598
rect 5324 35530 5330 35582
rect 5364 35530 5370 35582
rect 5324 35510 5370 35530
rect 5324 35462 5330 35510
rect 5364 35462 5370 35510
rect 5324 35438 5370 35462
rect 5324 35394 5330 35438
rect 5364 35394 5370 35438
rect 5324 35366 5370 35394
rect 5324 35326 5330 35366
rect 5364 35326 5370 35366
rect 5324 35294 5370 35326
rect 5324 35258 5330 35294
rect 5364 35258 5370 35294
rect 5324 35224 5370 35258
rect 5324 35188 5330 35224
rect 5364 35188 5370 35224
rect 5324 35156 5370 35188
rect 5324 35115 5330 35156
rect 5364 35115 5370 35156
rect 5324 35088 5370 35115
rect 5324 35042 5330 35088
rect 5364 35042 5370 35088
rect 5324 35020 5370 35042
rect 5324 34969 5330 35020
rect 5364 34969 5370 35020
rect 5324 34952 5370 34969
rect 5324 34896 5330 34952
rect 5364 34896 5370 34952
rect 5324 34884 5370 34896
rect 5324 34823 5330 34884
rect 5364 34823 5370 34884
rect 5324 34816 5370 34823
rect 5324 34750 5330 34816
rect 5364 34750 5370 34816
rect 5324 34748 5370 34750
rect 5324 34714 5330 34748
rect 5364 34714 5370 34748
rect 5324 34711 5370 34714
rect 5324 34646 5330 34711
rect 5364 34646 5370 34711
rect 5324 34638 5370 34646
rect 5324 34578 5330 34638
rect 5364 34578 5370 34638
rect 5324 34565 5370 34578
rect 5324 34510 5330 34565
rect 5364 34510 5370 34565
rect 5324 34492 5370 34510
rect 5324 34442 5330 34492
rect 5364 34442 5370 34492
rect 5324 34419 5370 34442
rect 5324 34374 5330 34419
rect 5364 34374 5370 34419
rect 5324 34346 5370 34374
rect 5324 34306 5330 34346
rect 5364 34306 5370 34346
rect 5324 34273 5370 34306
rect 5324 34238 5330 34273
rect 5364 34238 5370 34273
rect 5324 34204 5370 34238
rect 5324 34166 5330 34204
rect 5364 34166 5370 34204
rect 5324 34136 5370 34166
rect 5324 34093 5330 34136
rect 5364 34093 5370 34136
rect 5324 34068 5370 34093
rect 5324 34020 5330 34068
rect 5364 34020 5370 34068
rect 5324 34000 5370 34020
rect 5324 33947 5330 34000
rect 5364 33947 5370 34000
rect 5324 33932 5370 33947
rect 5324 33874 5330 33932
rect 5364 33874 5370 33932
rect 5324 33864 5370 33874
rect 5324 33801 5330 33864
rect 5364 33801 5370 33864
rect 5324 33796 5370 33801
rect 5324 33694 5330 33796
rect 5364 33694 5370 33796
rect 5324 33689 5370 33694
rect 5324 33626 5330 33689
rect 5364 33626 5370 33689
rect 5324 33616 5370 33626
rect 5324 33558 5330 33616
rect 5364 33558 5370 33616
rect 5324 33543 5370 33558
rect 5324 33490 5330 33543
rect 5364 33490 5370 33543
rect 5324 33470 5370 33490
rect 5324 33422 5330 33470
rect 5364 33422 5370 33470
rect 5324 33397 5370 33422
rect 5324 33354 5330 33397
rect 5364 33354 5370 33397
rect 5324 33324 5370 33354
rect 5324 33286 5330 33324
rect 5364 33286 5370 33324
rect 5324 33252 5370 33286
rect 5324 33217 5330 33252
rect 5364 33217 5370 33252
rect 5324 33184 5370 33217
rect 5324 33144 5330 33184
rect 5364 33144 5370 33184
rect 5324 33116 5370 33144
rect 5324 33071 5330 33116
rect 5364 33071 5370 33116
rect 5324 33048 5370 33071
rect 5324 32998 5330 33048
rect 5364 32998 5370 33048
rect 5324 32980 5370 32998
rect 5324 32925 5330 32980
rect 5364 32925 5370 32980
rect 5324 32912 5370 32925
rect 5324 32852 5330 32912
rect 5364 32852 5370 32912
rect 5324 32844 5370 32852
rect 5324 32779 5330 32844
rect 5364 32779 5370 32844
rect 5324 32776 5370 32779
rect 5324 32742 5330 32776
rect 5364 32742 5370 32776
rect 5324 32740 5370 32742
rect 5324 32674 5330 32740
rect 5364 32674 5370 32740
rect 5324 32667 5370 32674
rect 5324 32606 5330 32667
rect 5364 32606 5370 32667
rect 5324 32594 5370 32606
rect 5324 32538 5330 32594
rect 5364 32538 5370 32594
rect 5324 32521 5370 32538
rect 5324 32470 5330 32521
rect 5364 32470 5370 32521
rect 5324 32448 5370 32470
rect 5324 32402 5330 32448
rect 5364 32402 5370 32448
rect 5324 32375 5370 32402
rect 5324 32334 5330 32375
rect 5364 32334 5370 32375
rect 5324 32302 5370 32334
rect 5324 32266 5330 32302
rect 5364 32266 5370 32302
rect 5324 32232 5370 32266
rect 5324 32195 5330 32232
rect 5364 32195 5370 32232
rect 5324 32164 5370 32195
rect 5324 32122 5330 32164
rect 5364 32122 5370 32164
rect 5324 32096 5370 32122
rect 5324 32049 5330 32096
rect 5364 32049 5370 32096
rect 5324 32028 5370 32049
rect 5324 31976 5330 32028
rect 5364 31976 5370 32028
rect 5324 31960 5370 31976
rect 5324 31903 5330 31960
rect 5364 31903 5370 31960
rect 5324 31892 5370 31903
rect 5324 31830 5330 31892
rect 5364 31830 5370 31892
rect 5324 31824 5370 31830
rect 5324 31757 5330 31824
rect 5364 31757 5370 31824
rect 5324 31756 5370 31757
rect 5324 31722 5330 31756
rect 5364 31722 5370 31756
rect 5324 31718 5370 31722
rect 5324 31654 5330 31718
rect 5364 31654 5370 31718
rect 5324 31645 5370 31654
rect 5324 31586 5330 31645
rect 5364 31586 5370 31645
rect 5324 31572 5370 31586
rect 5324 31518 5330 31572
rect 5364 31518 5370 31572
rect 5324 31499 5370 31518
rect 5324 31450 5330 31499
rect 5364 31450 5370 31499
rect 5324 31426 5370 31450
rect 5324 31382 5330 31426
rect 5364 31382 5370 31426
rect 5324 31353 5370 31382
rect 5324 31314 5330 31353
rect 5364 31314 5370 31353
rect 5324 31280 5370 31314
rect 5324 31246 5330 31280
rect 5364 31246 5370 31280
rect 5324 31212 5370 31246
rect 5324 31173 5330 31212
rect 5364 31173 5370 31212
rect 5324 31144 5370 31173
rect 5324 31100 5330 31144
rect 5364 31100 5370 31144
rect 5324 31076 5370 31100
rect 5324 31027 5330 31076
rect 5364 31027 5370 31076
rect 5324 31008 5370 31027
rect 5324 30954 5330 31008
rect 5364 30954 5370 31008
rect 5324 30940 5370 30954
rect 5324 30881 5330 30940
rect 5364 30881 5370 30940
rect 5324 30872 5370 30881
rect 5324 30808 5330 30872
rect 5364 30808 5370 30872
rect 5324 30804 5370 30808
rect 5324 30770 5330 30804
rect 5364 30770 5370 30804
rect 5324 30769 5370 30770
rect 5324 30702 5330 30769
rect 5364 30702 5370 30769
rect 5324 30696 5370 30702
rect 5324 30634 5330 30696
rect 5364 30634 5370 30696
rect 5324 30623 5370 30634
rect 5324 30566 5330 30623
rect 5364 30566 5370 30623
rect 5324 30550 5370 30566
rect 5324 30498 5330 30550
rect 5364 30498 5370 30550
rect 5324 30477 5370 30498
rect 5324 30430 5330 30477
rect 5364 30430 5370 30477
rect 5324 30404 5370 30430
rect 3076 30332 3082 30378
rect 3116 30332 3122 30378
rect 5324 30362 5330 30404
rect 5364 30362 5370 30404
rect 5324 30332 5370 30362
rect 7740 39598 7786 39624
rect 7740 39552 7746 39598
rect 7780 39552 7786 39598
rect 7740 39530 7786 39552
rect 7740 39480 7746 39530
rect 7780 39480 7786 39530
rect 7740 39462 7786 39480
rect 7740 39408 7746 39462
rect 7780 39408 7786 39462
rect 7740 39394 7786 39408
rect 7740 39336 7746 39394
rect 7780 39336 7786 39394
rect 7740 39326 7786 39336
rect 7740 39264 7746 39326
rect 7780 39264 7786 39326
rect 7740 39258 7786 39264
rect 7740 39192 7746 39258
rect 7780 39192 7786 39258
rect 7740 39190 7786 39192
rect 7740 39156 7746 39190
rect 7780 39156 7786 39190
rect 7740 39154 7786 39156
rect 7740 39088 7746 39154
rect 7780 39088 7786 39154
rect 7740 39082 7786 39088
rect 7740 39020 7746 39082
rect 7780 39020 7786 39082
rect 7740 39010 7786 39020
rect 7740 38952 7746 39010
rect 7780 38952 7786 39010
rect 7740 38938 7786 38952
rect 7740 38884 7746 38938
rect 7780 38884 7786 38938
rect 7740 38866 7786 38884
rect 7740 38816 7746 38866
rect 7780 38816 7786 38866
rect 7740 38794 7786 38816
rect 7740 38748 7746 38794
rect 7780 38748 7786 38794
rect 7740 38722 7786 38748
rect 7740 38680 7746 38722
rect 7780 38680 7786 38722
rect 7740 38650 7786 38680
rect 7740 38612 7746 38650
rect 7780 38612 7786 38650
rect 7740 38578 7786 38612
rect 7740 38544 7746 38578
rect 7780 38544 7786 38578
rect 7740 38510 7786 38544
rect 7740 38472 7746 38510
rect 7780 38472 7786 38510
rect 7740 38442 7786 38472
rect 7740 38400 7746 38442
rect 7780 38400 7786 38442
rect 7740 38374 7786 38400
rect 7740 38328 7746 38374
rect 7780 38328 7786 38374
rect 7740 38306 7786 38328
rect 7740 38256 7746 38306
rect 7780 38256 7786 38306
rect 7740 38238 7786 38256
rect 7740 38184 7746 38238
rect 7780 38184 7786 38238
rect 7740 38170 7786 38184
rect 7740 38112 7746 38170
rect 7780 38112 7786 38170
rect 7740 38102 7786 38112
rect 7740 38040 7746 38102
rect 7780 38040 7786 38102
rect 7740 38034 7786 38040
rect 7740 37968 7746 38034
rect 7780 37968 7786 38034
rect 7740 37966 7786 37968
rect 7740 37932 7746 37966
rect 7780 37932 7786 37966
rect 7740 37930 7786 37932
rect 7740 37864 7746 37930
rect 7780 37864 7786 37930
rect 7740 37858 7786 37864
rect 7740 37796 7746 37858
rect 7780 37796 7786 37858
rect 7740 37786 7786 37796
rect 7740 37728 7746 37786
rect 7780 37728 7786 37786
rect 7740 37714 7786 37728
rect 7740 37660 7746 37714
rect 7780 37660 7786 37714
rect 7740 37642 7786 37660
rect 7740 37592 7746 37642
rect 7780 37592 7786 37642
rect 7740 37570 7786 37592
rect 7740 37524 7746 37570
rect 7780 37524 7786 37570
rect 7740 37498 7786 37524
rect 7740 37456 7746 37498
rect 7780 37456 7786 37498
rect 7740 37426 7786 37456
rect 7740 37388 7746 37426
rect 7780 37388 7786 37426
rect 7740 37354 7786 37388
rect 7740 37320 7746 37354
rect 7780 37320 7786 37354
rect 7740 37286 7786 37320
rect 7740 37248 7746 37286
rect 7780 37248 7786 37286
rect 7740 37218 7786 37248
rect 7740 37176 7746 37218
rect 7780 37176 7786 37218
rect 7740 37150 7786 37176
rect 7740 37104 7746 37150
rect 7780 37104 7786 37150
rect 7740 37082 7786 37104
rect 7740 37032 7746 37082
rect 7780 37032 7786 37082
rect 7740 37014 7786 37032
rect 7740 36960 7746 37014
rect 7780 36960 7786 37014
rect 7740 36946 7786 36960
rect 7740 36888 7746 36946
rect 7780 36888 7786 36946
rect 7740 36878 7786 36888
rect 7740 36816 7746 36878
rect 7780 36816 7786 36878
rect 7740 36810 7786 36816
rect 7740 36744 7746 36810
rect 7780 36744 7786 36810
rect 7740 36742 7786 36744
rect 7740 36708 7746 36742
rect 7780 36708 7786 36742
rect 7740 36706 7786 36708
rect 7740 36640 7746 36706
rect 7780 36640 7786 36706
rect 7740 36634 7786 36640
rect 7740 36572 7746 36634
rect 7780 36572 7786 36634
rect 7740 36562 7786 36572
rect 7740 36504 7746 36562
rect 7780 36504 7786 36562
rect 7740 36490 7786 36504
rect 7740 36436 7746 36490
rect 7780 36436 7786 36490
rect 7740 36418 7786 36436
rect 7740 36368 7746 36418
rect 7780 36368 7786 36418
rect 7740 36346 7786 36368
rect 7740 36300 7746 36346
rect 7780 36300 7786 36346
rect 7740 36274 7786 36300
rect 7740 36232 7746 36274
rect 7780 36232 7786 36274
rect 7740 36202 7786 36232
rect 7740 36164 7746 36202
rect 7780 36164 7786 36202
rect 7740 36130 7786 36164
rect 7740 36096 7746 36130
rect 7780 36096 7786 36130
rect 7740 36062 7786 36096
rect 7740 36024 7746 36062
rect 7780 36024 7786 36062
rect 7740 35994 7786 36024
rect 7740 35952 7746 35994
rect 7780 35952 7786 35994
rect 7740 35926 7786 35952
rect 7740 35880 7746 35926
rect 7780 35880 7786 35926
rect 7740 35858 7786 35880
rect 7740 35808 7746 35858
rect 7780 35808 7786 35858
rect 7740 35790 7786 35808
rect 7740 35736 7746 35790
rect 7780 35736 7786 35790
rect 7740 35722 7786 35736
rect 7740 35664 7746 35722
rect 7780 35664 7786 35722
rect 7740 35654 7786 35664
rect 7740 35592 7746 35654
rect 7780 35592 7786 35654
rect 7740 35586 7786 35592
rect 7740 35520 7746 35586
rect 7780 35520 7786 35586
rect 7740 35518 7786 35520
rect 7740 35484 7746 35518
rect 7780 35484 7786 35518
rect 7740 35482 7786 35484
rect 7740 35416 7746 35482
rect 7780 35416 7786 35482
rect 7740 35410 7786 35416
rect 7740 35348 7746 35410
rect 7780 35348 7786 35410
rect 7740 35338 7786 35348
rect 7740 35280 7746 35338
rect 7780 35280 7786 35338
rect 7740 35266 7786 35280
rect 7740 35212 7746 35266
rect 7780 35212 7786 35266
rect 7740 35194 7786 35212
rect 7740 35144 7746 35194
rect 7780 35144 7786 35194
rect 7740 35122 7786 35144
rect 7740 35076 7746 35122
rect 7780 35076 7786 35122
rect 7740 35050 7786 35076
rect 7740 35008 7746 35050
rect 7780 35008 7786 35050
rect 7740 34978 7786 35008
rect 7740 34940 7746 34978
rect 7780 34940 7786 34978
rect 7740 34906 7786 34940
rect 7740 34872 7746 34906
rect 7780 34872 7786 34906
rect 7740 34838 7786 34872
rect 7740 34800 7746 34838
rect 7780 34800 7786 34838
rect 7740 34770 7786 34800
rect 7740 34728 7746 34770
rect 7780 34728 7786 34770
rect 7740 34702 7786 34728
rect 7740 34656 7746 34702
rect 7780 34656 7786 34702
rect 7740 34634 7786 34656
rect 7740 34584 7746 34634
rect 7780 34584 7786 34634
rect 7740 34566 7786 34584
rect 7740 34512 7746 34566
rect 7780 34512 7786 34566
rect 7740 34498 7786 34512
rect 7740 34440 7746 34498
rect 7780 34440 7786 34498
rect 7740 34430 7786 34440
rect 7740 34368 7746 34430
rect 7780 34368 7786 34430
rect 7740 34362 7786 34368
rect 7740 34296 7746 34362
rect 7780 34296 7786 34362
rect 7740 34294 7786 34296
rect 7740 34260 7746 34294
rect 7780 34260 7786 34294
rect 7740 34258 7786 34260
rect 7740 34192 7746 34258
rect 7780 34192 7786 34258
rect 7740 34186 7786 34192
rect 7740 34124 7746 34186
rect 7780 34124 7786 34186
rect 7740 34114 7786 34124
rect 7740 34056 7746 34114
rect 7780 34056 7786 34114
rect 7740 34042 7786 34056
rect 7740 33988 7746 34042
rect 7780 33988 7786 34042
rect 7740 33970 7786 33988
rect 7740 33920 7746 33970
rect 7780 33920 7786 33970
rect 7740 33898 7786 33920
rect 7740 33852 7746 33898
rect 7780 33852 7786 33898
rect 7740 33826 7786 33852
rect 7740 33784 7746 33826
rect 7780 33784 7786 33826
rect 7740 33754 7786 33784
rect 7740 33716 7746 33754
rect 7780 33716 7786 33754
rect 7740 33682 7786 33716
rect 7740 33648 7746 33682
rect 7780 33648 7786 33682
rect 7740 33614 7786 33648
rect 7740 33576 7746 33614
rect 7780 33576 7786 33614
rect 7740 33546 7786 33576
rect 7740 33504 7746 33546
rect 7780 33504 7786 33546
rect 7740 33478 7786 33504
rect 7740 33432 7746 33478
rect 7780 33432 7786 33478
rect 7740 33410 7786 33432
rect 7740 33360 7746 33410
rect 7780 33360 7786 33410
rect 7740 33342 7786 33360
rect 7740 33288 7746 33342
rect 7780 33288 7786 33342
rect 7740 33274 7786 33288
rect 7740 33216 7746 33274
rect 7780 33216 7786 33274
rect 7740 33206 7786 33216
rect 7740 33144 7746 33206
rect 7780 33144 7786 33206
rect 7740 33138 7786 33144
rect 7740 33072 7746 33138
rect 7780 33072 7786 33138
rect 7740 33070 7786 33072
rect 7740 33036 7746 33070
rect 7780 33036 7786 33070
rect 7740 33034 7786 33036
rect 7740 32968 7746 33034
rect 7780 32968 7786 33034
rect 7740 32962 7786 32968
rect 7740 32900 7746 32962
rect 7780 32900 7786 32962
rect 7740 32890 7786 32900
rect 7740 32832 7746 32890
rect 7780 32832 7786 32890
rect 7740 32818 7786 32832
rect 7740 32764 7746 32818
rect 7780 32764 7786 32818
rect 7740 32746 7786 32764
rect 7740 32696 7746 32746
rect 7780 32696 7786 32746
rect 7740 32674 7786 32696
rect 7740 32628 7746 32674
rect 7780 32628 7786 32674
rect 7740 32602 7786 32628
rect 7740 32560 7746 32602
rect 7780 32560 7786 32602
rect 7740 32530 7786 32560
rect 7740 32492 7746 32530
rect 7780 32492 7786 32530
rect 7740 32458 7786 32492
rect 7740 32424 7746 32458
rect 7780 32424 7786 32458
rect 7740 32390 7786 32424
rect 7740 32352 7746 32390
rect 7780 32352 7786 32390
rect 7740 32322 7786 32352
rect 7740 32280 7746 32322
rect 7780 32280 7786 32322
rect 7740 32254 7786 32280
rect 7740 32208 7746 32254
rect 7780 32208 7786 32254
rect 7740 32186 7786 32208
rect 7740 32136 7746 32186
rect 7780 32136 7786 32186
rect 7740 32118 7786 32136
rect 7740 32064 7746 32118
rect 7780 32064 7786 32118
rect 7740 32050 7786 32064
rect 7740 31992 7746 32050
rect 7780 31992 7786 32050
rect 7740 31982 7786 31992
rect 7740 31920 7746 31982
rect 7780 31920 7786 31982
rect 7740 31914 7786 31920
rect 7740 31848 7746 31914
rect 7780 31848 7786 31914
rect 7740 31846 7786 31848
rect 7740 31812 7746 31846
rect 7780 31812 7786 31846
rect 7740 31810 7786 31812
rect 7740 31744 7746 31810
rect 7780 31744 7786 31810
rect 7740 31738 7786 31744
rect 7740 31676 7746 31738
rect 7780 31676 7786 31738
rect 7740 31666 7786 31676
rect 7740 31608 7746 31666
rect 7780 31608 7786 31666
rect 7740 31594 7786 31608
rect 7740 31540 7746 31594
rect 7780 31540 7786 31594
rect 7740 31522 7786 31540
rect 7740 31472 7746 31522
rect 7780 31472 7786 31522
rect 7740 31450 7786 31472
rect 7740 31404 7746 31450
rect 7780 31404 7786 31450
rect 7740 31378 7786 31404
rect 7740 31336 7746 31378
rect 7780 31336 7786 31378
rect 7740 31306 7786 31336
rect 7740 31268 7746 31306
rect 7780 31268 7786 31306
rect 7740 31234 7786 31268
rect 7740 31200 7746 31234
rect 7780 31200 7786 31234
rect 7740 31166 7786 31200
rect 7740 31128 7746 31166
rect 7780 31128 7786 31166
rect 7740 31098 7786 31128
rect 7740 31056 7746 31098
rect 7780 31056 7786 31098
rect 7740 31030 7786 31056
rect 7740 30984 7746 31030
rect 7780 30984 7786 31030
rect 7740 30962 7786 30984
rect 7740 30912 7746 30962
rect 7780 30912 7786 30962
rect 7740 30894 7786 30912
rect 7740 30840 7746 30894
rect 7780 30840 7786 30894
rect 7740 30826 7786 30840
rect 7740 30767 7746 30826
rect 7780 30767 7786 30826
rect 7740 30758 7786 30767
rect 7740 30694 7746 30758
rect 7780 30694 7786 30758
rect 7740 30690 7786 30694
rect 7740 30656 7746 30690
rect 7780 30656 7786 30690
rect 7740 30655 7786 30656
rect 7740 30588 7746 30655
rect 7780 30588 7786 30655
rect 7740 30582 7786 30588
rect 7740 30520 7746 30582
rect 7780 30520 7786 30582
rect 7740 30509 7786 30520
rect 7740 30452 7746 30509
rect 7780 30452 7786 30509
rect 7740 30436 7786 30452
rect 7740 30384 7746 30436
rect 7780 30384 7786 30436
rect 7740 30363 7786 30384
rect 3076 30306 3122 30332
rect 5330 30328 5364 30332
rect 3076 30264 3082 30306
rect 3116 30264 3122 30306
rect 3076 30234 3122 30264
rect 3076 30196 3082 30234
rect 3116 30196 3122 30234
rect 7740 30316 7746 30363
rect 7780 30316 7786 30363
rect 7740 30290 7786 30316
rect 7740 30248 7746 30290
rect 7780 30248 7786 30290
rect 7740 30217 7786 30248
rect 3076 30162 3122 30196
rect 5640 30163 5646 30197
rect 5698 30163 5721 30197
rect 5769 30163 5796 30197
rect 5840 30163 5871 30197
rect 5911 30163 5946 30197
rect 5982 30163 6019 30197
rect 6055 30163 6090 30197
rect 6130 30163 6161 30197
rect 6205 30163 6232 30197
rect 6280 30163 6303 30197
rect 6355 30163 6374 30197
rect 6430 30163 6444 30197
rect 6505 30163 6514 30197
rect 6580 30163 6584 30197
rect 6618 30163 6621 30197
rect 6688 30163 6696 30197
rect 6758 30163 6770 30197
rect 6828 30163 6844 30197
rect 6898 30163 6918 30197
rect 6968 30163 6992 30197
rect 7038 30163 7066 30197
rect 7108 30163 7140 30197
rect 7178 30163 7214 30197
rect 7248 30163 7284 30197
rect 7322 30163 7354 30197
rect 7396 30163 7424 30197
rect 7470 30163 7482 30197
rect 7740 30180 7746 30217
rect 7780 30180 7786 30217
rect 3076 30128 3082 30162
rect 3116 30128 3122 30162
rect 3076 30094 3122 30128
rect 7740 30146 7786 30180
rect 3723 30123 3764 30125
rect 3798 30123 3839 30125
rect 3873 30123 3914 30125
rect 3948 30123 3989 30125
rect 4023 30123 4064 30125
rect 4098 30123 4139 30125
rect 4173 30123 4214 30125
rect 4248 30123 4289 30125
rect 4323 30123 4364 30125
rect 4398 30123 4439 30125
rect 4473 30123 4514 30125
rect 4548 30123 4589 30125
rect 4623 30123 4664 30125
rect 4698 30123 4739 30125
rect 4773 30123 4814 30125
rect 4848 30123 4889 30125
rect 4923 30123 4964 30125
rect 4998 30123 5038 30125
rect 3076 30056 3082 30094
rect 3116 30056 3122 30094
rect 3604 30089 3620 30123
rect 3654 30091 3689 30123
rect 3654 30089 3690 30091
rect 3724 30089 3760 30123
rect 3798 30091 3830 30123
rect 3873 30091 3899 30123
rect 3948 30091 3968 30123
rect 4023 30091 4037 30123
rect 4098 30091 4106 30123
rect 4173 30091 4175 30123
rect 3794 30089 3830 30091
rect 3864 30089 3899 30091
rect 3933 30089 3968 30091
rect 4002 30089 4037 30091
rect 4071 30089 4106 30091
rect 4140 30089 4175 30091
rect 4209 30091 4214 30123
rect 4278 30091 4289 30123
rect 4347 30091 4364 30123
rect 4416 30091 4439 30123
rect 4485 30091 4514 30123
rect 4209 30089 4244 30091
rect 4278 30089 4313 30091
rect 4347 30089 4382 30091
rect 4416 30089 4451 30091
rect 4485 30089 4520 30091
rect 4554 30089 4589 30123
rect 4623 30089 4658 30123
rect 4698 30091 4727 30123
rect 4773 30091 4796 30123
rect 4848 30091 4865 30123
rect 4923 30091 4934 30123
rect 4998 30091 5003 30123
rect 4692 30089 4727 30091
rect 4761 30089 4796 30091
rect 4830 30089 4865 30091
rect 4899 30089 4934 30091
rect 4968 30089 5003 30091
rect 5037 30091 5038 30123
rect 5072 30123 5112 30125
rect 5146 30123 5186 30125
rect 5037 30089 5072 30091
rect 5106 30091 5112 30123
rect 5175 30091 5186 30123
rect 5106 30089 5141 30091
rect 5175 30089 5210 30091
rect 5244 30089 5260 30123
rect 7740 30110 7746 30146
rect 7780 30110 7786 30146
rect 7740 30078 7786 30110
rect 3076 30026 3122 30056
rect 5640 30040 5674 30068
rect 3076 29984 3082 30026
rect 3116 29984 3122 30026
rect 3076 29958 3122 29984
rect 3076 29912 3082 29958
rect 3116 29912 3122 29958
rect 3076 29890 3122 29912
rect 3076 29840 3082 29890
rect 3116 29840 3122 29890
rect 3076 29822 3122 29840
rect 3076 29768 3082 29822
rect 3116 29768 3122 29822
rect 3076 29754 3122 29768
rect 3076 29696 3082 29754
rect 3116 29696 3122 29754
rect 3076 29686 3122 29696
rect 3076 29624 3082 29686
rect 3116 29624 3122 29686
rect 3076 29618 3122 29624
rect 3076 29552 3082 29618
rect 3116 29552 3122 29618
rect 3076 29550 3122 29552
rect 3076 29516 3082 29550
rect 3116 29516 3122 29550
rect 3076 29514 3122 29516
rect 3076 29448 3082 29514
rect 3116 29448 3122 29514
rect 3076 29442 3122 29448
rect 3076 29380 3082 29442
rect 3116 29380 3122 29442
rect 3076 29370 3122 29380
rect 3076 29312 3082 29370
rect 3116 29312 3122 29370
rect 3076 29298 3122 29312
rect 3076 29244 3082 29298
rect 3116 29244 3122 29298
rect 5634 30002 5680 30040
rect 5634 29964 5640 30002
rect 5674 29964 5680 30002
rect 5634 29930 5680 29964
rect 5634 29894 5640 29930
rect 5674 29894 5680 29930
rect 5634 29862 5680 29894
rect 7740 30037 7746 30078
rect 7780 30037 7786 30078
rect 7740 30010 7786 30037
rect 7740 29964 7746 30010
rect 7780 29964 7786 30010
rect 7740 29942 7786 29964
rect 7740 29891 7746 29942
rect 7780 29891 7786 29942
rect 5634 29820 5640 29862
rect 5674 29820 5680 29862
rect 6271 29854 6286 29888
rect 6339 29854 6355 29888
rect 6411 29854 6427 29888
rect 6480 29854 6495 29888
rect 7740 29874 7786 29891
rect 5634 29794 5680 29820
rect 5634 29746 5640 29794
rect 5674 29746 5680 29794
rect 5634 29726 5680 29746
rect 5634 29672 5640 29726
rect 5674 29672 5680 29726
rect 5634 29658 5680 29672
rect 5634 29597 5640 29658
rect 5674 29597 5680 29658
rect 5634 29590 5680 29597
rect 5634 29488 5640 29590
rect 5674 29488 5680 29590
rect 5634 29481 5680 29488
rect 5634 29420 5640 29481
rect 5674 29420 5680 29481
rect 5634 29406 5680 29420
rect 5634 29352 5640 29406
rect 5674 29352 5680 29406
rect 5634 29331 5680 29352
rect 5634 29284 5640 29331
rect 5674 29284 5680 29331
rect 3076 29226 3122 29244
rect 3604 29235 3620 29269
rect 3654 29235 3690 29269
rect 3749 29235 3760 29269
rect 3823 29235 3830 29269
rect 3897 29235 3899 29269
rect 3933 29235 3937 29269
rect 4002 29235 4011 29269
rect 4071 29235 4085 29269
rect 4140 29235 4159 29269
rect 4209 29235 4232 29269
rect 4278 29235 4305 29269
rect 4347 29235 4378 29269
rect 4416 29235 4451 29269
rect 4485 29235 4520 29269
rect 4558 29235 4589 29269
rect 4631 29235 4658 29269
rect 4704 29235 4727 29269
rect 4777 29235 4796 29269
rect 4850 29235 4865 29269
rect 4923 29235 4934 29269
rect 4996 29235 5003 29269
rect 5069 29235 5072 29269
rect 5106 29235 5108 29269
rect 5175 29235 5181 29269
rect 5244 29235 5260 29269
rect 5634 29256 5680 29284
rect 3076 29176 3082 29226
rect 3116 29176 3122 29226
rect 3076 29154 3122 29176
rect 3076 29108 3082 29154
rect 3116 29108 3122 29154
rect 5634 29216 5640 29256
rect 5674 29216 5680 29256
rect 5634 29182 5680 29216
rect 5634 29147 5640 29182
rect 5674 29147 5680 29182
rect 3076 29082 3122 29108
rect 3604 29105 3620 29139
rect 3654 29105 3690 29139
rect 3749 29105 3760 29139
rect 3826 29105 3830 29139
rect 3864 29105 3869 29139
rect 3933 29105 3946 29139
rect 4002 29105 4023 29139
rect 4071 29105 4100 29139
rect 4140 29105 4175 29139
rect 4211 29105 4244 29139
rect 4288 29105 4313 29139
rect 4364 29105 4382 29139
rect 4416 29105 4451 29139
rect 4485 29105 4515 29139
rect 4554 29105 4589 29139
rect 4624 29105 4658 29139
rect 4699 29105 4727 29139
rect 4774 29105 4796 29139
rect 4849 29105 4865 29139
rect 4924 29105 4934 29139
rect 4999 29105 5003 29139
rect 5037 29105 5040 29139
rect 5106 29105 5115 29139
rect 5175 29105 5189 29139
rect 5244 29105 5260 29139
rect 5634 29114 5680 29147
rect 3076 29040 3082 29082
rect 3116 29040 3122 29082
rect 3076 29010 3122 29040
rect 3076 28972 3082 29010
rect 3116 28972 3122 29010
rect 3076 28938 3122 28972
rect 3076 28904 3082 28938
rect 3116 28904 3122 28938
rect 3076 28870 3122 28904
rect 3076 28832 3082 28870
rect 3116 28832 3122 28870
rect 3076 28802 3122 28832
rect 3076 28760 3082 28802
rect 3116 28760 3122 28802
rect 3076 28734 3122 28760
rect 3076 28688 3082 28734
rect 3116 28688 3122 28734
rect 3076 28666 3122 28688
rect 3076 28616 3082 28666
rect 3116 28616 3122 28666
rect 3076 28598 3122 28616
rect 3076 28544 3082 28598
rect 3116 28544 3122 28598
rect 3076 28530 3122 28544
rect 3076 28472 3082 28530
rect 3116 28472 3122 28530
rect 3076 28440 3122 28472
rect 5634 29072 5640 29114
rect 5674 29072 5680 29114
rect 5634 29046 5680 29072
rect 5634 28997 5640 29046
rect 5674 28997 5680 29046
rect 5634 28978 5680 28997
rect 5634 28922 5640 28978
rect 5674 28922 5680 28978
rect 5634 28910 5680 28922
rect 5634 28847 5640 28910
rect 5674 28847 5680 28910
rect 5634 28842 5680 28847
rect 5634 28808 5640 28842
rect 5674 28808 5680 28842
rect 5634 28806 5680 28808
rect 5634 28740 5640 28806
rect 5674 28740 5680 28806
rect 5634 28731 5680 28740
rect 5634 28672 5640 28731
rect 5674 28672 5680 28731
rect 5634 28656 5680 28672
rect 5634 28604 5640 28656
rect 5674 28604 5680 28656
rect 5634 28581 5680 28604
rect 5634 28536 5640 28581
rect 5674 28536 5680 28581
rect 5634 28506 5680 28536
rect 5634 28468 5640 28506
rect 5674 28468 5680 28506
rect 5634 28440 5680 28468
rect 3076 28434 5680 28440
rect 3076 28400 3150 28434
rect 3188 28400 3218 28434
rect 3262 28400 3286 28434
rect 3336 28400 3354 28434
rect 3410 28400 3422 28434
rect 3484 28400 3490 28434
rect 3557 28400 3558 28434
rect 3592 28400 3596 28434
rect 3660 28400 3669 28434
rect 3728 28400 3742 28434
rect 3796 28400 3815 28434
rect 3864 28400 3888 28434
rect 3932 28400 3961 28434
rect 4000 28400 4034 28434
rect 4068 28400 4102 28434
rect 4141 28400 4170 28434
rect 4214 28400 4238 28434
rect 4287 28400 4306 28434
rect 4360 28400 4374 28434
rect 4433 28400 4442 28434
rect 4506 28400 4510 28434
rect 4544 28400 4545 28434
rect 4612 28400 4618 28434
rect 4680 28400 4691 28434
rect 4748 28400 4764 28434
rect 4816 28400 4837 28434
rect 4884 28400 4910 28434
rect 4952 28400 4983 28434
rect 5020 28400 5054 28434
rect 5090 28400 5122 28434
rect 5163 28400 5190 28434
rect 5236 28400 5258 28434
rect 5309 28400 5326 28434
rect 5382 28400 5394 28434
rect 5455 28400 5462 28434
rect 5528 28400 5530 28434
rect 5564 28400 5567 28434
rect 5601 28400 5680 28434
rect 3076 28394 5680 28400
rect 7740 29818 7746 29874
rect 7780 29818 7786 29874
rect 7740 29806 7786 29818
rect 7740 29745 7746 29806
rect 7780 29745 7786 29806
rect 7740 29738 7786 29745
rect 7740 29672 7746 29738
rect 7780 29672 7786 29738
rect 7740 29670 7786 29672
rect 7740 29636 7746 29670
rect 7780 29636 7786 29670
rect 7740 29633 7786 29636
rect 7740 29568 7746 29633
rect 7780 29568 7786 29633
rect 7740 29560 7786 29568
rect 7740 29500 7746 29560
rect 7780 29500 7786 29560
rect 7740 29487 7786 29500
rect 7740 29432 7746 29487
rect 7780 29432 7786 29487
rect 7740 29414 7786 29432
rect 7740 29364 7746 29414
rect 7780 29364 7786 29414
rect 7740 29341 7786 29364
rect 7740 29296 7746 29341
rect 7780 29296 7786 29341
rect 7740 29268 7786 29296
rect 7740 29228 7746 29268
rect 7780 29228 7786 29268
rect 7740 29195 7786 29228
rect 7740 29160 7746 29195
rect 7780 29160 7786 29195
rect 7740 29126 7786 29160
rect 7740 29088 7746 29126
rect 7780 29088 7786 29126
rect 7740 29058 7786 29088
rect 7740 29015 7746 29058
rect 7780 29015 7786 29058
rect 7740 28990 7786 29015
rect 7740 28942 7746 28990
rect 7780 28942 7786 28990
rect 7740 28922 7786 28942
rect 7740 28869 7746 28922
rect 7780 28869 7786 28922
rect 7740 28854 7786 28869
rect 7740 28796 7746 28854
rect 7780 28796 7786 28854
rect 7740 28786 7786 28796
rect 7740 28723 7746 28786
rect 7780 28723 7786 28786
rect 7740 28718 7786 28723
rect 7740 28616 7746 28718
rect 7780 28616 7786 28718
rect 7740 28611 7786 28616
rect 7740 28548 7746 28611
rect 7780 28548 7786 28611
rect 7740 28538 7786 28548
rect 7740 28480 7746 28538
rect 7780 28480 7786 28538
rect 7740 28465 7786 28480
rect 7740 28412 7746 28465
rect 7780 28412 7786 28465
rect 2816 28348 2822 28390
rect 2856 28348 2862 28390
rect 2816 28318 2862 28348
rect 2816 28284 2822 28318
rect 2856 28284 2862 28318
rect 2816 28266 2862 28284
rect 2816 28212 2822 28266
rect 2856 28212 2862 28266
rect 2816 28180 2862 28212
rect 7740 28392 7786 28412
rect 7740 28344 7746 28392
rect 7780 28344 7786 28392
rect 7740 28319 7786 28344
rect 7740 28276 7746 28319
rect 7780 28276 7786 28319
rect 7740 28246 7786 28276
rect 7740 28208 7746 28246
rect 7780 28208 7786 28246
rect 7740 28180 7786 28208
rect 2816 28174 7786 28180
rect 2816 28140 2890 28174
rect 2928 28140 2958 28174
rect 3001 28140 3026 28174
rect 3074 28140 3094 28174
rect 3147 28140 3162 28174
rect 3220 28140 3230 28174
rect 3293 28140 3298 28174
rect 3400 28140 3405 28174
rect 3468 28140 3478 28174
rect 3536 28140 3551 28174
rect 3604 28140 3624 28174
rect 3672 28140 3697 28174
rect 3740 28140 3770 28174
rect 3808 28140 3842 28174
rect 3877 28140 3910 28174
rect 3950 28140 3978 28174
rect 4023 28140 4046 28174
rect 4096 28140 4114 28174
rect 4169 28140 4182 28174
rect 4242 28140 4250 28174
rect 4315 28140 4318 28174
rect 4352 28140 4354 28174
rect 4420 28140 4427 28174
rect 4488 28140 4500 28174
rect 4556 28140 4573 28174
rect 4624 28140 4646 28174
rect 4692 28140 4719 28174
rect 4760 28140 4792 28174
rect 4828 28140 4862 28174
rect 4899 28140 4930 28174
rect 4972 28140 4998 28174
rect 5044 28140 5066 28174
rect 5116 28140 5134 28174
rect 5188 28140 5202 28174
rect 5260 28140 5270 28174
rect 5332 28140 5338 28174
rect 5404 28140 5406 28174
rect 5440 28140 5442 28174
rect 5508 28140 5514 28174
rect 5576 28140 5586 28174
rect 5644 28140 5658 28174
rect 5712 28140 5730 28174
rect 5780 28140 5802 28174
rect 5848 28140 5874 28174
rect 5916 28140 5946 28174
rect 5984 28140 6018 28174
rect 6052 28140 6086 28174
rect 6124 28140 6154 28174
rect 6196 28140 6222 28174
rect 6268 28140 6290 28174
rect 6340 28140 6358 28174
rect 6412 28140 6426 28174
rect 6484 28140 6494 28174
rect 6556 28140 6562 28174
rect 6628 28140 6630 28174
rect 6664 28140 6666 28174
rect 6732 28140 6738 28174
rect 6800 28140 6810 28174
rect 6868 28140 6882 28174
rect 6936 28140 6954 28174
rect 7004 28140 7026 28174
rect 7072 28140 7098 28174
rect 7140 28140 7170 28174
rect 7208 28140 7242 28174
rect 7276 28140 7310 28174
rect 7348 28140 7378 28174
rect 7420 28140 7446 28174
rect 7492 28140 7514 28174
rect 7564 28140 7582 28174
rect 7636 28140 7650 28174
rect 7708 28140 7786 28174
rect 2816 28134 7786 28140
rect 4398 26165 4414 26199
rect 4448 26165 4485 26199
rect 4519 26165 4556 26199
rect 4590 26165 4627 26199
rect 4661 26165 4698 26199
rect 4732 26165 4769 26199
rect 4803 26165 4840 26199
rect 4874 26165 4910 26199
rect 4944 26165 4980 26199
rect 5014 26165 5050 26199
rect 5093 26165 5120 26199
rect 5172 26165 5190 26199
rect 5251 26165 5260 26199
rect 5294 26165 5295 26199
rect 5329 26165 5330 26199
rect 5364 26165 5373 26199
rect 5434 26165 5451 26199
rect 5504 26165 5529 26199
rect 5574 26165 5590 26199
rect 5946 26082 5980 26116
rect 4008 26041 4042 26048
rect 4008 25966 4042 25980
rect 4008 25891 4042 25912
rect 4008 25816 4042 25844
rect 4008 25742 4042 25776
rect 2590 25651 2678 25685
rect 2712 25651 2746 25685
rect 2780 25651 2814 25685
rect 2848 25651 2850 25685
rect 2916 25651 2928 25685
rect 2984 25651 3005 25685
rect 3052 25651 3082 25685
rect 3120 25651 3154 25685
rect 3193 25651 3222 25685
rect 3270 25651 3290 25685
rect 3347 25651 3358 25685
rect 3424 25651 3426 25685
rect 3460 25651 3467 25685
rect 3528 25651 3544 25685
rect 3596 25651 3621 25685
rect 3664 25651 3732 25685
rect 3698 25613 3732 25651
rect 3698 25541 3732 25575
rect 2745 25472 2832 25506
rect 2866 25472 2904 25506
rect 2745 25404 2938 25472
rect 3570 25472 3608 25506
rect 3536 25398 3642 25472
rect 3698 25473 3732 25506
rect 3698 25405 3732 25433
rect 3698 25337 3732 25360
rect 3698 25269 3732 25287
rect 3698 25201 3732 25214
rect 3698 25133 3732 25141
rect 3698 25065 3732 25068
rect 3698 25029 3732 25031
rect 3698 24956 3732 24963
rect 3698 24883 3732 24895
rect 3698 24810 3732 24827
rect 3698 24737 3732 24759
rect 4008 25674 4042 25706
rect 4008 25606 4042 25630
rect 4008 25538 4042 25554
rect 4008 25470 4042 25478
rect 4008 25360 4042 25368
rect 4008 25284 4042 25300
rect 4008 25208 4042 25232
rect 4008 25132 4042 25164
rect 4008 25062 4042 25096
rect 4008 24994 4042 25022
rect 4008 24926 4042 24946
rect 4008 24858 4042 24870
rect 4008 24790 4042 24794
rect 4008 24752 4042 24756
rect 4353 25998 4387 26037
rect 4353 25925 4387 25964
rect 4353 25852 4387 25891
rect 4353 25779 4387 25818
rect 4353 25706 4387 25745
rect 4353 25633 4387 25672
rect 4353 25560 4387 25599
rect 4353 25487 4387 25526
rect 4353 25413 4387 25453
rect 4353 25339 4387 25379
rect 4353 25265 4387 25305
rect 4353 25191 4387 25231
rect 4353 25117 4387 25157
rect 4353 25043 4387 25083
rect 4353 24969 4387 25009
rect 4353 24895 4387 24935
rect 4353 24821 4387 24861
rect 4353 24747 4387 24787
rect 4509 25998 4543 26037
rect 4509 25925 4543 25964
rect 4509 25852 4543 25891
rect 4509 25779 4543 25818
rect 4509 25706 4543 25745
rect 4509 25633 4543 25672
rect 4509 25560 4543 25599
rect 4509 25487 4543 25526
rect 4509 25413 4543 25453
rect 4509 25339 4543 25379
rect 4509 25265 4543 25305
rect 4509 25191 4543 25231
rect 4509 25117 4543 25157
rect 4509 25043 4543 25083
rect 4509 24969 4543 25009
rect 4509 24895 4543 24935
rect 4509 24821 4543 24861
rect 4509 24747 4543 24787
rect 4665 25998 4699 26037
rect 4665 25925 4699 25964
rect 4665 25852 4699 25891
rect 4665 25779 4699 25818
rect 4665 25706 4699 25745
rect 4665 25633 4699 25672
rect 4665 25560 4699 25599
rect 4665 25487 4699 25526
rect 4665 25413 4699 25453
rect 4665 25339 4699 25379
rect 4665 25265 4699 25305
rect 4665 25191 4699 25231
rect 4665 25117 4699 25157
rect 4665 25043 4699 25083
rect 4665 24969 4699 25009
rect 4665 24895 4699 24935
rect 4665 24821 4699 24861
rect 4665 24747 4699 24787
rect 4821 25998 4855 26037
rect 4821 25925 4855 25964
rect 4821 25852 4855 25891
rect 4821 25779 4855 25818
rect 4821 25706 4855 25745
rect 4821 25633 4855 25672
rect 4821 25560 4855 25599
rect 4821 25487 4855 25526
rect 4821 25413 4855 25453
rect 4821 25339 4855 25379
rect 4821 25265 4855 25305
rect 4821 25191 4855 25231
rect 4821 25117 4855 25157
rect 4821 25043 4855 25083
rect 4821 24969 4855 25009
rect 4821 24895 4855 24935
rect 4821 24821 4855 24861
rect 4821 24747 4855 24787
rect 4977 25998 5011 26037
rect 4977 25925 5011 25964
rect 4977 25852 5011 25891
rect 4977 25779 5011 25818
rect 4977 25706 5011 25745
rect 4977 25633 5011 25672
rect 4977 25560 5011 25599
rect 4977 25487 5011 25526
rect 4977 25413 5011 25453
rect 4977 25339 5011 25379
rect 4977 25265 5011 25305
rect 4977 25191 5011 25231
rect 4977 25117 5011 25157
rect 4977 25043 5011 25083
rect 4977 24969 5011 25009
rect 4977 24895 5011 24935
rect 4977 24821 5011 24861
rect 4977 24747 5011 24787
rect 5133 25998 5167 26037
rect 5133 25925 5167 25964
rect 5133 25852 5167 25891
rect 5133 25779 5167 25818
rect 5133 25706 5167 25745
rect 5133 25633 5167 25672
rect 5133 25560 5167 25599
rect 5133 25487 5167 25526
rect 5133 25413 5167 25453
rect 5133 25339 5167 25379
rect 5133 25265 5167 25305
rect 5133 25191 5167 25231
rect 5133 25117 5167 25157
rect 5133 25043 5167 25083
rect 5133 24969 5167 25009
rect 5133 24895 5167 24935
rect 5133 24821 5167 24861
rect 5133 24747 5167 24787
rect 5289 25998 5323 26037
rect 5289 25925 5323 25964
rect 5289 25852 5323 25891
rect 5289 25779 5323 25818
rect 5289 25706 5323 25745
rect 5289 25633 5323 25672
rect 5289 25560 5323 25599
rect 5289 25487 5323 25526
rect 5289 25413 5323 25453
rect 5289 25339 5323 25379
rect 5289 25265 5323 25305
rect 5289 25191 5323 25231
rect 5289 25117 5323 25157
rect 5289 25043 5323 25083
rect 5289 24969 5323 25009
rect 5289 24895 5323 24935
rect 5289 24821 5323 24861
rect 5289 24747 5323 24787
rect 5445 25998 5479 26037
rect 5445 25925 5479 25964
rect 5445 25852 5479 25891
rect 5445 25779 5479 25818
rect 5445 25706 5479 25745
rect 5445 25633 5479 25672
rect 5445 25560 5479 25599
rect 5445 25487 5479 25526
rect 5445 25413 5479 25453
rect 5445 25339 5479 25379
rect 5445 25265 5479 25305
rect 5445 25191 5479 25231
rect 5445 25117 5479 25157
rect 5445 25043 5479 25083
rect 5445 24969 5479 25009
rect 5445 24895 5479 24935
rect 5445 24821 5479 24861
rect 5445 24747 5479 24787
rect 5601 25998 5635 26037
rect 5601 25925 5635 25964
rect 5601 25852 5635 25891
rect 5601 25779 5635 25818
rect 5601 25706 5635 25745
rect 5601 25633 5635 25672
rect 5601 25560 5635 25599
rect 5601 25487 5635 25526
rect 5601 25413 5635 25453
rect 5601 25339 5635 25379
rect 5601 25265 5635 25305
rect 5601 25191 5635 25231
rect 5601 25117 5635 25157
rect 5601 25043 5635 25083
rect 5601 24969 5635 25009
rect 5601 24895 5635 24935
rect 5601 24821 5635 24861
rect 5601 24747 5635 24787
rect 5946 26014 5980 26037
rect 5946 25946 5980 25964
rect 5946 25878 5980 25891
rect 5946 25810 5980 25818
rect 5946 25742 5980 25745
rect 5946 25706 5980 25708
rect 5946 25633 5980 25640
rect 5946 25560 5980 25572
rect 5946 25487 5980 25504
rect 5946 25413 5980 25436
rect 5946 25339 5980 25368
rect 5946 25266 5980 25300
rect 5946 25198 5980 25231
rect 5946 25130 5980 25157
rect 5946 25062 5980 25083
rect 5946 24994 5980 25009
rect 5946 24926 5980 24935
rect 5946 24858 5980 24861
rect 5946 24821 5980 24824
rect 5946 24747 5980 24756
rect 3698 24664 3732 24691
rect 3698 24591 3732 24623
rect 3698 24521 3732 24555
rect 3698 24453 3732 24484
rect 3698 24385 3732 24411
rect 3698 24317 3732 24338
rect 3698 24249 3732 24265
rect 3698 24181 3732 24192
rect 3698 24113 3732 24119
rect 3698 24045 3732 24046
rect 3698 24007 3732 24011
rect 3698 23934 3732 23943
rect 3698 23861 3732 23875
rect 3698 23788 3732 23807
rect 3698 23715 3732 23739
rect 3698 23642 3732 23671
rect 3698 23569 3732 23603
rect 3698 23501 3732 23535
rect 3698 23433 3732 23462
rect 3698 23365 3732 23389
rect 3698 23297 3732 23316
rect 3698 23229 3732 23243
rect 3698 23161 3732 23170
rect 3698 23093 3732 23097
rect 3698 23058 3732 23059
rect 3698 22985 3732 22991
rect 3698 22912 3732 22923
rect 3698 22839 3732 22855
rect 3698 22766 3732 22787
rect 3698 22693 3732 22719
rect 3698 22621 3732 22651
rect 3698 22549 3732 22583
rect 3698 22481 3732 22515
rect 3698 22413 3732 22443
rect 3698 22345 3732 22371
rect 3698 22277 3732 22299
rect 3698 22209 3732 22227
rect 3698 22141 3732 22155
rect 3698 22073 3732 22083
rect 3698 22005 3732 22011
rect 3698 21937 3732 21939
rect 3698 21901 3732 21903
rect 3698 21829 3732 21835
rect 3698 21757 3732 21767
rect 3698 21685 3732 21699
rect 3698 21613 3732 21631
rect 3698 21541 3732 21563
rect 3698 21469 3732 21495
rect 3698 21397 3732 21427
rect 3698 21325 3732 21359
rect 3698 21257 3732 21291
rect 3698 21189 3732 21219
rect 3698 21121 3732 21147
rect 3698 21053 3732 21075
rect 3698 20985 3732 21003
rect 3698 20917 3732 20931
rect 3698 20849 3732 20859
rect 3698 20781 3732 20787
rect 3698 20713 3732 20715
rect 3698 20677 3732 20679
rect 3698 20605 3732 20611
rect 3698 20533 3732 20543
rect 3698 20461 3732 20475
rect 3698 20389 3732 20407
rect 3698 20317 3732 20339
rect 3698 20245 3732 20271
rect 3698 20173 3732 20203
rect 3698 20101 3732 20135
rect 3698 20033 3732 20067
rect 3698 19965 3732 19995
rect 3698 19897 3732 19923
rect 3698 19829 3732 19851
rect 3698 19761 3732 19779
rect 3698 19693 3732 19707
rect 3698 19625 3732 19635
rect 3698 19557 3732 19563
rect 3698 19489 3732 19491
rect 3698 19453 3732 19455
rect 3698 19381 3732 19387
rect 3698 19309 3732 19319
rect 3698 19237 3732 19251
rect 3698 19165 3732 19183
rect 3698 19093 3732 19115
rect 3698 19021 3732 19047
rect 3698 18949 3732 18979
rect 3698 18877 3732 18911
rect 3698 18809 3732 18843
rect 3698 18741 3732 18771
rect 3698 18673 3732 18699
rect 3698 18605 3732 18627
rect 3698 18537 3732 18555
rect 4454 24184 5898 24190
rect 4454 24150 4528 24184
rect 4589 24150 4596 24184
rect 4630 24150 4664 24184
rect 4721 24150 4732 24184
rect 4794 24150 4800 24184
rect 4867 24150 4868 24184
rect 4902 24150 4906 24184
rect 4970 24150 4979 24184
rect 5038 24150 5052 24184
rect 5106 24150 5125 24184
rect 5174 24150 5198 24184
rect 5242 24150 5271 24184
rect 5310 24150 5344 24184
rect 5378 24150 5412 24184
rect 5451 24150 5480 24184
rect 5524 24150 5548 24184
rect 5598 24150 5616 24184
rect 5672 24150 5684 24184
rect 5746 24150 5752 24184
rect 5820 24150 5898 24184
rect 4454 24144 5898 24150
rect 4454 24112 4500 24144
rect 4454 24076 4460 24112
rect 4494 24076 4500 24112
rect 4454 24039 4500 24076
rect 4454 24005 4460 24039
rect 4494 24005 4500 24039
rect 4454 23966 4500 24005
rect 4454 23922 4460 23966
rect 4494 23922 4500 23966
rect 4454 23893 4500 23922
rect 4454 23854 4460 23893
rect 4494 23854 4500 23893
rect 5852 24116 5898 24144
rect 5852 24078 5858 24116
rect 5892 24078 5898 24116
rect 5852 24048 5898 24078
rect 5852 24006 5858 24048
rect 5892 24006 5898 24048
rect 5852 23980 5898 24006
rect 5852 23934 5858 23980
rect 5892 23934 5898 23980
rect 5852 23912 5898 23934
rect 5852 23862 5858 23912
rect 5892 23862 5898 23912
rect 4454 23820 4500 23854
rect 4454 23786 4460 23820
rect 4494 23786 4500 23820
rect 4454 23752 4500 23786
rect 4454 23713 4460 23752
rect 4494 23713 4500 23752
rect 4685 23800 4731 23834
rect 4765 23800 4810 23834
rect 4651 23762 4844 23800
rect 4685 23728 4731 23762
rect 4765 23728 4810 23762
rect 5852 23844 5898 23862
rect 5852 23790 5858 23844
rect 5892 23790 5898 23844
rect 5852 23776 5898 23790
rect 5852 23718 5858 23776
rect 5892 23718 5898 23776
rect 4454 23684 4500 23713
rect 4454 23640 4460 23684
rect 4494 23640 4500 23684
rect 4454 23616 4500 23640
rect 4454 23567 4460 23616
rect 4494 23567 4500 23616
rect 4454 23548 4500 23567
rect 4454 23494 4460 23548
rect 4494 23494 4500 23548
rect 4454 23480 4500 23494
rect 4454 23421 4460 23480
rect 4494 23421 4500 23480
rect 4454 23412 4500 23421
rect 4454 23348 4460 23412
rect 4494 23348 4500 23412
rect 4454 23344 4500 23348
rect 4454 23310 4460 23344
rect 4494 23310 4500 23344
rect 4454 23309 4500 23310
rect 4454 23242 4460 23309
rect 4494 23242 4500 23309
rect 4454 23236 4500 23242
rect 4454 23174 4460 23236
rect 4494 23174 4500 23236
rect 4454 23163 4500 23174
rect 4454 23106 4460 23163
rect 4494 23106 4500 23163
rect 4454 23090 4500 23106
rect 4454 23038 4460 23090
rect 4494 23038 4500 23090
rect 4454 23017 4500 23038
rect 4454 22970 4460 23017
rect 4494 22970 4500 23017
rect 4454 22944 4500 22970
rect 4454 22902 4460 22944
rect 4494 22902 4500 22944
rect 4454 22871 4500 22902
rect 4454 22834 4460 22871
rect 4494 22834 4500 22871
rect 4454 22800 4500 22834
rect 4454 22764 4460 22800
rect 4494 22764 4500 22800
rect 4454 22732 4500 22764
rect 4454 22691 4460 22732
rect 4494 22691 4500 22732
rect 4454 22664 4500 22691
rect 4454 22618 4460 22664
rect 4494 22618 4500 22664
rect 4454 22596 4500 22618
rect 4454 22545 4460 22596
rect 4494 22545 4500 22596
rect 4454 22528 4500 22545
rect 4454 22472 4460 22528
rect 4494 22472 4500 22528
rect 4454 22460 4500 22472
rect 4454 22399 4460 22460
rect 4494 22399 4500 22460
rect 4454 22392 4500 22399
rect 4454 22326 4460 22392
rect 4494 22326 4500 22392
rect 4454 22324 4500 22326
rect 4454 22290 4460 22324
rect 4494 22290 4500 22324
rect 4454 22287 4500 22290
rect 4454 22222 4460 22287
rect 4494 22222 4500 22287
rect 4454 22214 4500 22222
rect 4454 22154 4460 22214
rect 4494 22154 4500 22214
rect 4454 22141 4500 22154
rect 4454 22086 4460 22141
rect 4494 22086 4500 22141
rect 4888 23701 4922 23717
rect 4888 23660 4922 23667
rect 4888 23587 4922 23597
rect 4888 23514 4922 23527
rect 4888 23441 4922 23457
rect 4888 23368 4922 23387
rect 4888 23295 4922 23317
rect 4888 23222 4922 23247
rect 4888 23149 4922 23177
rect 4888 23076 4922 23107
rect 4888 23003 4922 23037
rect 4888 22931 4922 22967
rect 4888 22861 4922 22896
rect 4888 22791 4922 22823
rect 4888 22721 4922 22750
rect 4888 22651 4922 22677
rect 4888 22581 4922 22604
rect 4888 22512 4922 22531
rect 4888 22443 4922 22458
rect 4888 22374 4922 22385
rect 4888 22305 4922 22312
rect 4888 22236 4922 22239
rect 4888 22200 4922 22202
rect 4888 22127 4922 22133
rect 4454 22068 4500 22086
rect 4676 22072 4715 22106
rect 4749 22072 4788 22106
rect 4454 22018 4460 22068
rect 4494 22018 4500 22068
rect 4454 21995 4500 22018
rect 4454 21950 4460 21995
rect 4494 21950 4500 21995
rect 4454 21922 4500 21950
rect 4454 21882 4460 21922
rect 4494 21882 4500 21922
rect 4454 21849 4500 21882
rect 4454 21814 4460 21849
rect 4494 21814 4500 21849
rect 4454 21780 4500 21814
rect 4454 21742 4460 21780
rect 4494 21742 4500 21780
rect 4454 21712 4500 21742
rect 4454 21669 4460 21712
rect 4494 21669 4500 21712
rect 4454 21644 4500 21669
rect 4454 21596 4460 21644
rect 4494 21596 4500 21644
rect 4454 21576 4500 21596
rect 4454 21523 4460 21576
rect 4494 21523 4500 21576
rect 4454 21508 4500 21523
rect 4454 21450 4460 21508
rect 4494 21450 4500 21508
rect 4454 21440 4500 21450
rect 4454 21377 4460 21440
rect 4494 21377 4500 21440
rect 4454 21372 4500 21377
rect 4454 21270 4460 21372
rect 4494 21270 4500 21372
rect 4454 21265 4500 21270
rect 4454 21202 4460 21265
rect 4494 21202 4500 21265
rect 4454 21192 4500 21202
rect 4454 21134 4460 21192
rect 4494 21134 4500 21192
rect 4454 21119 4500 21134
rect 4454 21066 4460 21119
rect 4494 21066 4500 21119
rect 4454 21046 4500 21066
rect 4454 20998 4460 21046
rect 4494 20998 4500 21046
rect 4454 20973 4500 20998
rect 4454 20930 4460 20973
rect 4494 20930 4500 20973
rect 4454 20900 4500 20930
rect 4454 20862 4460 20900
rect 4494 20862 4500 20900
rect 4454 20828 4500 20862
rect 4454 20793 4460 20828
rect 4494 20793 4500 20828
rect 4454 20760 4500 20793
rect 4454 20720 4460 20760
rect 4494 20720 4500 20760
rect 4454 20692 4500 20720
rect 4454 20647 4460 20692
rect 4494 20647 4500 20692
rect 4454 20624 4500 20647
rect 4454 20574 4460 20624
rect 4494 20574 4500 20624
rect 4454 20556 4500 20574
rect 4454 20501 4460 20556
rect 4494 20501 4500 20556
rect 4454 20488 4500 20501
rect 4454 20428 4460 20488
rect 4494 20428 4500 20488
rect 4888 22054 4922 22064
rect 4888 21981 4922 21995
rect 4888 21908 4922 21926
rect 4888 21835 4922 21857
rect 4888 21762 4922 21788
rect 4888 21689 4922 21719
rect 4888 21616 4922 21650
rect 4888 21546 4922 21581
rect 4888 21477 4922 21509
rect 4888 21408 4922 21436
rect 4888 21339 4922 21363
rect 4888 21270 4922 21290
rect 4888 21201 4922 21217
rect 4888 21132 4922 21144
rect 4888 21063 4922 21071
rect 4888 20994 4922 20998
rect 4888 20959 4922 20960
rect 4888 20886 4922 20891
rect 4888 20813 4922 20822
rect 4888 20740 4922 20753
rect 4888 20667 4922 20684
rect 4888 20594 4922 20615
rect 4888 20520 4922 20546
rect 4888 20461 4922 20477
rect 5196 23701 5230 23717
rect 5196 23637 5230 23667
rect 5196 23564 5230 23597
rect 5196 23493 5230 23528
rect 5196 23424 5230 23457
rect 5196 23355 5230 23384
rect 5196 23286 5230 23311
rect 5196 23217 5230 23238
rect 5196 23148 5230 23165
rect 5196 23079 5230 23092
rect 5196 23010 5230 23019
rect 5196 22941 5230 22946
rect 5196 22872 5230 22873
rect 5196 22834 5230 22838
rect 5196 22761 5230 22769
rect 5196 22688 5230 22700
rect 5196 22615 5230 22631
rect 5196 22542 5230 22562
rect 5196 22469 5230 22493
rect 5196 22396 5230 22424
rect 5196 22323 5230 22355
rect 5196 22251 5230 22286
rect 5196 22182 5230 22216
rect 5196 22113 5230 22143
rect 5196 22044 5230 22070
rect 5196 21975 5230 21997
rect 5196 21906 5230 21924
rect 5196 21837 5230 21851
rect 5196 21768 5230 21778
rect 5196 21699 5230 21705
rect 5196 21630 5230 21632
rect 5196 21593 5230 21596
rect 5196 21520 5230 21527
rect 5196 21447 5230 21458
rect 5196 21374 5230 21389
rect 5196 21301 5230 21320
rect 5196 21228 5230 21251
rect 5196 21155 5230 21182
rect 5196 21082 5230 21113
rect 5196 21009 5230 21044
rect 5196 20940 5230 20975
rect 5196 20871 5230 20902
rect 5196 20802 5230 20829
rect 5196 20733 5230 20756
rect 5196 20664 5230 20683
rect 5196 20595 5230 20610
rect 5196 20526 5230 20537
rect 5196 20457 5230 20464
rect 4454 20420 4500 20428
rect 4454 20355 4460 20420
rect 4494 20355 4500 20420
rect 4454 20352 4500 20355
rect 4454 20318 4460 20352
rect 4494 20318 4500 20352
rect 4676 20411 4726 20445
rect 4760 20411 4810 20445
rect 4642 20373 4844 20411
rect 4676 20339 4726 20373
rect 4760 20339 4810 20373
rect 5196 20388 5230 20391
rect 5196 20352 5230 20354
rect 4454 20316 4500 20318
rect 4454 20250 4460 20316
rect 4494 20250 4500 20316
rect 4454 20244 4500 20250
rect 4454 20182 4460 20244
rect 4494 20182 4500 20244
rect 4454 20172 4500 20182
rect 4454 20114 4460 20172
rect 4494 20114 4500 20172
rect 4454 20100 4500 20114
rect 4454 20046 4460 20100
rect 4494 20046 4500 20100
rect 5196 20278 5230 20285
rect 5196 20204 5230 20216
rect 5196 20130 5230 20147
rect 4619 20059 4660 20093
rect 4694 20059 4735 20093
rect 4769 20059 4809 20093
rect 5196 20056 5230 20078
rect 4454 20028 4500 20046
rect 4454 19978 4460 20028
rect 4494 19978 4500 20028
rect 4454 19956 4500 19978
rect 4454 19910 4460 19956
rect 4494 19910 4500 19956
rect 4899 20036 4933 20048
rect 4899 19964 4933 19998
rect 4454 19884 4500 19910
rect 4676 19903 4726 19937
rect 4760 19903 4809 19937
rect 4454 19842 4460 19884
rect 4494 19842 4500 19884
rect 4454 19812 4500 19842
rect 4454 19774 4460 19812
rect 4494 19774 4500 19812
rect 4899 19891 4933 19927
rect 4899 19818 4933 19856
rect 4454 19740 4500 19774
rect 4619 19747 4657 19781
rect 4691 19747 4729 19781
rect 4454 19706 4460 19740
rect 4494 19706 4500 19740
rect 4454 19672 4500 19706
rect 4454 19634 4460 19672
rect 4494 19634 4500 19672
rect 4454 19604 4500 19634
rect 4899 19746 4933 19784
rect 5196 19982 5230 20009
rect 5196 19908 5230 19940
rect 5196 19836 5230 19871
rect 5196 19767 5230 19800
rect 5196 19717 5230 19733
rect 5452 23701 5486 23717
rect 5452 23637 5486 23667
rect 5452 23564 5486 23597
rect 5452 23493 5486 23528
rect 5452 23424 5486 23457
rect 5452 23355 5486 23384
rect 5452 23286 5486 23311
rect 5452 23217 5486 23238
rect 5452 23148 5486 23165
rect 5452 23079 5486 23092
rect 5452 23010 5486 23019
rect 5452 22941 5486 22946
rect 5452 22872 5486 22873
rect 5452 22834 5486 22838
rect 5452 22761 5486 22769
rect 5452 22688 5486 22700
rect 5452 22615 5486 22631
rect 5452 22542 5486 22562
rect 5452 22469 5486 22493
rect 5452 22396 5486 22424
rect 5452 22323 5486 22355
rect 5452 22251 5486 22286
rect 5452 22182 5486 22216
rect 5452 22113 5486 22143
rect 5452 22044 5486 22070
rect 5452 21975 5486 21997
rect 5452 21906 5486 21924
rect 5452 21837 5486 21851
rect 5452 21768 5486 21778
rect 5452 21699 5486 21705
rect 5452 21630 5486 21632
rect 5452 21593 5486 21596
rect 5452 21520 5486 21527
rect 5452 21447 5486 21458
rect 5452 21374 5486 21389
rect 5452 21301 5486 21320
rect 5452 21228 5486 21251
rect 5452 21155 5486 21182
rect 5452 21082 5486 21113
rect 5452 21009 5486 21044
rect 5452 20940 5486 20975
rect 5452 20871 5486 20902
rect 5452 20802 5486 20829
rect 5452 20733 5486 20756
rect 5452 20664 5486 20683
rect 5452 20595 5486 20610
rect 5452 20526 5486 20537
rect 5452 20457 5486 20464
rect 5452 20388 5486 20391
rect 5452 20352 5486 20354
rect 5452 20278 5486 20285
rect 5452 20204 5486 20216
rect 5452 20130 5486 20147
rect 5452 20056 5486 20078
rect 5452 19982 5486 20009
rect 5452 19908 5486 19940
rect 5452 19836 5486 19871
rect 5452 19767 5486 19800
rect 5452 19717 5486 19733
rect 5852 23708 5898 23718
rect 5852 23646 5858 23708
rect 5892 23646 5898 23708
rect 5852 23640 5898 23646
rect 5852 23574 5858 23640
rect 5892 23574 5898 23640
rect 5852 23572 5898 23574
rect 5852 23538 5858 23572
rect 5892 23538 5898 23572
rect 5852 23536 5898 23538
rect 5852 23470 5858 23536
rect 5892 23470 5898 23536
rect 5852 23464 5898 23470
rect 5852 23402 5858 23464
rect 5892 23402 5898 23464
rect 5852 23392 5898 23402
rect 5852 23334 5858 23392
rect 5892 23334 5898 23392
rect 5852 23320 5898 23334
rect 5852 23266 5858 23320
rect 5892 23266 5898 23320
rect 5852 23248 5898 23266
rect 5852 23198 5858 23248
rect 5892 23198 5898 23248
rect 5852 23176 5898 23198
rect 5852 23130 5858 23176
rect 5892 23130 5898 23176
rect 5852 23104 5898 23130
rect 5852 23062 5858 23104
rect 5892 23062 5898 23104
rect 5852 23032 5898 23062
rect 5852 22994 5858 23032
rect 5892 22994 5898 23032
rect 5852 22960 5898 22994
rect 5852 22926 5858 22960
rect 5892 22926 5898 22960
rect 5852 22892 5898 22926
rect 5852 22854 5858 22892
rect 5892 22854 5898 22892
rect 5852 22824 5898 22854
rect 5852 22782 5858 22824
rect 5892 22782 5898 22824
rect 5852 22756 5898 22782
rect 5852 22710 5858 22756
rect 5892 22710 5898 22756
rect 5852 22688 5898 22710
rect 5852 22638 5858 22688
rect 5892 22638 5898 22688
rect 5852 22620 5898 22638
rect 5852 22566 5858 22620
rect 5892 22566 5898 22620
rect 5852 22552 5898 22566
rect 5852 22494 5858 22552
rect 5892 22494 5898 22552
rect 5852 22484 5898 22494
rect 5852 22422 5858 22484
rect 5892 22422 5898 22484
rect 5852 22416 5898 22422
rect 5852 22350 5858 22416
rect 5892 22350 5898 22416
rect 5852 22348 5898 22350
rect 5852 22314 5858 22348
rect 5892 22314 5898 22348
rect 5852 22311 5898 22314
rect 5852 22246 5858 22311
rect 5892 22246 5898 22311
rect 5852 22238 5898 22246
rect 5852 22178 5858 22238
rect 5892 22178 5898 22238
rect 5852 22165 5898 22178
rect 5852 22110 5858 22165
rect 5892 22110 5898 22165
rect 5852 22092 5898 22110
rect 5852 22042 5858 22092
rect 5892 22042 5898 22092
rect 5852 22019 5898 22042
rect 5852 21974 5858 22019
rect 5892 21974 5898 22019
rect 7397 22000 7412 22034
rect 7465 22000 7481 22034
rect 7537 22000 7553 22034
rect 7606 22000 7621 22034
rect 5852 21946 5898 21974
rect 5852 21906 5858 21946
rect 5892 21906 5898 21946
rect 5852 21873 5898 21906
rect 5852 21838 5858 21873
rect 5892 21838 5898 21873
rect 5852 21804 5898 21838
rect 5852 21766 5858 21804
rect 5892 21766 5898 21804
rect 5852 21736 5898 21766
rect 5852 21693 5858 21736
rect 5892 21693 5898 21736
rect 5852 21668 5898 21693
rect 5852 21620 5858 21668
rect 5892 21620 5898 21668
rect 5852 21600 5898 21620
rect 5852 21547 5858 21600
rect 5892 21547 5898 21600
rect 5852 21532 5898 21547
rect 5852 21474 5858 21532
rect 5892 21474 5898 21532
rect 7326 21485 7342 21519
rect 7376 21485 7417 21519
rect 7454 21485 7488 21519
rect 7526 21485 7556 21519
rect 7601 21485 7624 21519
rect 7676 21485 7692 21519
rect 5852 21464 5898 21474
rect 5852 21401 5858 21464
rect 5892 21401 5898 21464
rect 5852 21396 5898 21401
rect 5852 21294 5858 21396
rect 5892 21294 5898 21396
rect 5852 21289 5898 21294
rect 5852 21226 5858 21289
rect 5892 21226 5898 21289
rect 5852 21216 5898 21226
rect 5852 21158 5858 21216
rect 5892 21158 5898 21216
rect 5852 21143 5898 21158
rect 5852 21090 5858 21143
rect 5892 21090 5898 21143
rect 5852 21070 5898 21090
rect 5852 21022 5858 21070
rect 5892 21022 5898 21070
rect 5852 20997 5898 21022
rect 5852 20954 5858 20997
rect 5892 20954 5898 20997
rect 5852 20924 5898 20954
rect 5852 20886 5858 20924
rect 5892 20886 5898 20924
rect 5852 20852 5898 20886
rect 5852 20817 5858 20852
rect 5892 20817 5898 20852
rect 5852 20784 5898 20817
rect 5852 20744 5858 20784
rect 5892 20744 5898 20784
rect 5852 20716 5898 20744
rect 5852 20671 5858 20716
rect 5892 20671 5898 20716
rect 5852 20648 5898 20671
rect 5852 20598 5858 20648
rect 5892 20598 5898 20648
rect 5852 20580 5898 20598
rect 5852 20525 5858 20580
rect 5892 20525 5898 20580
rect 5852 20512 5898 20525
rect 5852 20452 5858 20512
rect 5892 20452 5898 20512
rect 5852 20444 5898 20452
rect 5852 20379 5858 20444
rect 5892 20379 5898 20444
rect 5852 20376 5898 20379
rect 5852 20342 5858 20376
rect 5892 20342 5898 20376
rect 5852 20340 5898 20342
rect 5852 20274 5858 20340
rect 5892 20274 5898 20340
rect 5852 20267 5898 20274
rect 5852 20206 5858 20267
rect 5892 20206 5898 20267
rect 5852 20194 5898 20206
rect 5852 20138 5858 20194
rect 5892 20138 5898 20194
rect 5852 20121 5898 20138
rect 5852 20070 5858 20121
rect 5892 20070 5898 20121
rect 5852 20048 5898 20070
rect 5852 20002 5858 20048
rect 5892 20002 5898 20048
rect 5852 19975 5898 20002
rect 5852 19934 5858 19975
rect 5892 19934 5898 19975
rect 5852 19902 5898 19934
rect 5852 19866 5858 19902
rect 5892 19866 5898 19902
rect 5852 19832 5898 19866
rect 5852 19795 5858 19832
rect 5892 19795 5898 19832
rect 5852 19764 5898 19795
rect 5852 19722 5858 19764
rect 5892 19722 5898 19764
rect 4899 19674 4933 19711
rect 4454 19562 4460 19604
rect 4494 19562 4500 19604
rect 4676 19591 4726 19625
rect 4760 19591 4809 19625
rect 4899 19602 4933 19638
rect 4454 19536 4500 19562
rect 4454 19490 4460 19536
rect 4494 19490 4500 19536
rect 4454 19468 4500 19490
rect 5120 19666 5152 19684
rect 5086 19638 5152 19666
rect 5086 19628 5102 19638
rect 5136 19604 5152 19638
rect 5342 19666 5362 19677
rect 5852 19696 5898 19722
rect 5396 19666 5408 19677
rect 5342 19638 5408 19666
rect 5342 19604 5358 19638
rect 5392 19628 5408 19638
rect 5396 19604 5408 19628
rect 5852 19649 5858 19696
rect 5892 19649 5898 19696
rect 5852 19628 5898 19649
rect 5120 19594 5152 19604
rect 4899 19530 4933 19565
rect 4899 19480 4933 19492
rect 5852 19576 5858 19628
rect 5892 19576 5898 19628
rect 5852 19560 5898 19576
rect 5852 19503 5858 19560
rect 5892 19503 5898 19560
rect 5852 19492 5898 19503
rect 4454 19418 4460 19468
rect 4494 19418 4500 19468
rect 4619 19435 4660 19469
rect 4694 19435 4735 19469
rect 4769 19435 4809 19469
rect 4454 19400 4500 19418
rect 4454 19346 4460 19400
rect 4494 19346 4500 19400
rect 4454 19332 4500 19346
rect 4454 19274 4460 19332
rect 4494 19274 4500 19332
rect 4454 19264 4500 19274
rect 4454 19202 4460 19264
rect 4494 19202 4500 19264
rect 4454 19196 4500 19202
rect 4454 19130 4460 19196
rect 4494 19130 4500 19196
rect 4454 19128 4500 19130
rect 4454 19094 4460 19128
rect 4494 19094 4500 19128
rect 4454 19092 4500 19094
rect 4454 19026 4460 19092
rect 4494 19026 4500 19092
rect 5852 19430 5858 19492
rect 5892 19430 5898 19492
rect 5852 19424 5898 19430
rect 5852 19357 5858 19424
rect 5892 19357 5898 19424
rect 5852 19356 5898 19357
rect 5852 19322 5858 19356
rect 5892 19322 5898 19356
rect 5852 19318 5898 19322
rect 5852 19254 5858 19318
rect 5892 19254 5898 19318
rect 5852 19245 5898 19254
rect 5852 19186 5858 19245
rect 5892 19186 5898 19245
rect 5852 19172 5898 19186
rect 5852 19118 5858 19172
rect 5892 19118 5898 19172
rect 5852 19099 5898 19118
rect 5042 19034 5058 19068
rect 5114 19034 5152 19068
rect 5186 19034 5192 19068
rect 5226 19034 5242 19068
rect 5852 19050 5858 19099
rect 5892 19050 5898 19099
rect 4454 19020 4500 19026
rect 4454 18958 4460 19020
rect 4494 18958 4500 19020
rect 4454 18948 4500 18958
rect 4454 18890 4460 18948
rect 4494 18890 4500 18948
rect 4454 18876 4500 18890
rect 4454 18822 4460 18876
rect 4494 18822 4500 18876
rect 4454 18804 4500 18822
rect 4454 18754 4460 18804
rect 4494 18754 4500 18804
rect 4454 18732 4500 18754
rect 4454 18686 4460 18732
rect 4494 18686 4500 18732
rect 4454 18660 4500 18686
rect 4454 18618 4460 18660
rect 4494 18618 4500 18660
rect 4454 18588 4500 18618
rect 4454 18550 4460 18588
rect 4494 18550 4500 18588
rect 4454 18522 4500 18550
rect 5852 19026 5898 19050
rect 5852 18982 5858 19026
rect 5892 18982 5898 19026
rect 5852 18953 5898 18982
rect 5852 18914 5858 18953
rect 5892 18914 5898 18953
rect 5852 18880 5898 18914
rect 5852 18846 5858 18880
rect 5892 18846 5898 18880
rect 5852 18812 5898 18846
rect 5852 18773 5858 18812
rect 5892 18773 5898 18812
rect 5852 18744 5898 18773
rect 5852 18700 5858 18744
rect 5892 18700 5898 18744
rect 5852 18676 5898 18700
rect 5852 18627 5858 18676
rect 5892 18627 5898 18676
rect 5852 18608 5898 18627
rect 5852 18554 5858 18608
rect 5892 18554 5898 18608
rect 5852 18522 5898 18554
rect 4454 18516 5898 18522
rect 4454 18482 4532 18516
rect 4600 18482 4606 18516
rect 4668 18482 4680 18516
rect 4736 18482 4754 18516
rect 4804 18482 4828 18516
rect 4872 18482 4902 18516
rect 4940 18482 4974 18516
rect 5010 18482 5042 18516
rect 5084 18482 5110 18516
rect 5158 18482 5178 18516
rect 5232 18482 5246 18516
rect 5306 18482 5314 18516
rect 5380 18482 5382 18516
rect 5416 18482 5420 18516
rect 5484 18482 5493 18516
rect 5552 18482 5566 18516
rect 5620 18482 5639 18516
rect 5688 18482 5712 18516
rect 5756 18482 5785 18516
rect 5824 18482 5898 18516
rect 4454 18476 5898 18482
rect 2816 18289 6790 18295
rect 2816 18255 2890 18289
rect 2933 18255 2958 18289
rect 3011 18255 3026 18289
rect 3089 18255 3094 18289
rect 3128 18255 3133 18289
rect 3196 18255 3211 18289
rect 3264 18255 3289 18289
rect 3332 18255 3366 18289
rect 3401 18255 3434 18289
rect 3479 18255 3502 18289
rect 3557 18255 3570 18289
rect 3635 18255 3638 18289
rect 3672 18255 3679 18289
rect 3740 18255 3774 18289
rect 3823 18255 3842 18289
rect 3895 18255 3910 18289
rect 3967 18255 3978 18289
rect 4039 18255 4046 18289
rect 4111 18255 4114 18289
rect 4148 18255 4149 18289
rect 4216 18255 4221 18289
rect 4284 18255 4293 18289
rect 4352 18255 4365 18289
rect 4420 18255 4437 18289
rect 4488 18255 4509 18289
rect 4556 18255 4581 18289
rect 4624 18255 4653 18289
rect 4692 18255 4725 18289
rect 4760 18255 4794 18289
rect 4831 18255 4862 18289
rect 4903 18255 4930 18289
rect 4975 18255 4998 18289
rect 5047 18255 5066 18289
rect 5119 18255 5134 18289
rect 5191 18255 5202 18289
rect 5263 18255 5270 18289
rect 5335 18255 5338 18289
rect 5372 18255 5373 18289
rect 5440 18255 5445 18289
rect 5508 18255 5517 18289
rect 5576 18255 5589 18289
rect 5644 18255 5661 18289
rect 5712 18255 5733 18289
rect 5780 18255 5805 18289
rect 5848 18255 5877 18289
rect 5916 18255 5949 18289
rect 5984 18255 6018 18289
rect 6055 18255 6086 18289
rect 6128 18255 6154 18289
rect 6201 18255 6222 18289
rect 6274 18255 6290 18289
rect 6347 18255 6358 18289
rect 6420 18255 6426 18289
rect 6493 18255 6494 18289
rect 6528 18255 6532 18289
rect 6596 18255 6605 18289
rect 6664 18255 6678 18289
rect 6712 18255 6790 18289
rect 2816 18249 6790 18255
rect 2816 18217 2862 18249
rect 2816 18163 2822 18217
rect 2856 18163 2862 18217
rect 2816 18143 2862 18163
rect 2816 18109 2822 18143
rect 2856 18109 2862 18143
rect 2816 18083 2862 18109
rect 2816 18035 2822 18083
rect 2856 18035 2862 18083
rect 6744 18221 6790 18249
rect 6744 18182 6750 18221
rect 6784 18182 6790 18221
rect 6744 18153 6790 18182
rect 6744 18109 6750 18153
rect 6784 18109 6790 18153
rect 6744 18085 6790 18109
rect 6744 18036 6750 18085
rect 6784 18036 6790 18085
rect 2816 18015 2862 18035
rect 2816 17961 2822 18015
rect 2856 17961 2862 18015
rect 2816 17947 2862 17961
rect 2816 17887 2822 17947
rect 2856 17887 2862 17947
rect 2816 17879 2862 17887
rect 2816 17813 2822 17879
rect 2856 17813 2862 17879
rect 2816 17811 2862 17813
rect 2816 17777 2822 17811
rect 2856 17777 2862 17811
rect 2816 17774 2862 17777
rect 2816 17709 2822 17774
rect 2856 17709 2862 17774
rect 2816 17701 2862 17709
rect 2816 17641 2822 17701
rect 2856 17641 2862 17701
rect 2816 17628 2862 17641
rect 2816 17573 2822 17628
rect 2856 17573 2862 17628
rect 2816 17555 2862 17573
rect 2816 17505 2822 17555
rect 2856 17505 2862 17555
rect 2816 17482 2862 17505
rect 2816 17437 2822 17482
rect 2856 17437 2862 17482
rect 2816 17409 2862 17437
rect 2816 17369 2822 17409
rect 2856 17369 2862 17409
rect 2816 17336 2862 17369
rect 2816 17301 2822 17336
rect 2856 17301 2862 17336
rect 2816 17267 2862 17301
rect 2816 17229 2822 17267
rect 2856 17229 2862 17267
rect 2816 17199 2862 17229
rect 2816 17156 2822 17199
rect 2856 17156 2862 17199
rect 2816 17131 2862 17156
rect 2816 17083 2822 17131
rect 2856 17083 2862 17131
rect 2816 17063 2862 17083
rect 2816 17010 2822 17063
rect 2856 17010 2862 17063
rect 2816 16995 2862 17010
rect 2816 16937 2822 16995
rect 2856 16937 2862 16995
rect 2816 16927 2862 16937
rect 2816 16864 2822 16927
rect 2856 16864 2862 16927
rect 2816 16859 2862 16864
rect 2816 16757 2822 16859
rect 2856 16757 2862 16859
rect 2816 16752 2862 16757
rect 2816 16689 2822 16752
rect 2856 16689 2862 16752
rect 2816 16679 2862 16689
rect 2816 16621 2822 16679
rect 2856 16621 2862 16679
rect 2816 16606 2862 16621
rect 2816 16553 2822 16606
rect 2856 16553 2862 16606
rect 2816 16533 2862 16553
rect 2816 16485 2822 16533
rect 2856 16485 2862 16533
rect 2816 16460 2862 16485
rect 2816 16417 2822 16460
rect 2856 16417 2862 16460
rect 2816 16387 2862 16417
rect 2816 16349 2822 16387
rect 2856 16349 2862 16387
rect 2816 16315 2862 16349
rect 2816 16280 2822 16315
rect 2856 16280 2862 16315
rect 2816 16247 2862 16280
rect 2816 16207 2822 16247
rect 2856 16207 2862 16247
rect 2816 16179 2862 16207
rect 2816 16134 2822 16179
rect 2856 16134 2862 16179
rect 2816 16111 2862 16134
rect 2816 16061 2822 16111
rect 2856 16061 2862 16111
rect 2816 16043 2862 16061
rect 2816 15988 2822 16043
rect 2856 15988 2862 16043
rect 2816 15975 2862 15988
rect 2816 15915 2822 15975
rect 2856 15915 2862 15975
rect 2816 15907 2862 15915
rect 2816 15842 2822 15907
rect 2856 15842 2862 15907
rect 2816 15839 2862 15842
rect 2816 15805 2822 15839
rect 2856 15805 2862 15839
rect 2816 15803 2862 15805
rect 2816 15737 2822 15803
rect 2856 15737 2862 15803
rect 2816 15730 2862 15737
rect 2816 15669 2822 15730
rect 2856 15669 2862 15730
rect 2816 15657 2862 15669
rect 2816 15601 2822 15657
rect 2856 15601 2862 15657
rect 2816 15584 2862 15601
rect 2816 15533 2822 15584
rect 2856 15533 2862 15584
rect 2816 15511 2862 15533
rect 2816 15465 2822 15511
rect 2856 15465 2862 15511
rect 2816 15438 2862 15465
rect 2816 15397 2822 15438
rect 2856 15397 2862 15438
rect 2816 15365 2862 15397
rect 2816 15329 2822 15365
rect 2856 15329 2862 15365
rect 2816 15295 2862 15329
rect 2816 15258 2822 15295
rect 2856 15258 2862 15295
rect 2816 15227 2862 15258
rect 2816 15185 2822 15227
rect 2856 15185 2862 15227
rect 2816 15159 2862 15185
rect 2816 15112 2822 15159
rect 2856 15112 2862 15159
rect 2816 15091 2862 15112
rect 2816 15039 2822 15091
rect 2856 15039 2862 15091
rect 2816 15023 2862 15039
rect 2816 14966 2822 15023
rect 2856 14966 2862 15023
rect 2816 14955 2862 14966
rect 2816 14893 2822 14955
rect 2856 14893 2862 14955
rect 2816 14887 2862 14893
rect 2816 14820 2822 14887
rect 2856 14820 2862 14887
rect 2816 14819 2862 14820
rect 2816 14785 2822 14819
rect 2856 14785 2862 14819
rect 2816 14781 2862 14785
rect 2816 14717 2822 14781
rect 2856 14717 2862 14781
rect 2816 14708 2862 14717
rect 2816 14649 2822 14708
rect 2856 14649 2862 14708
rect 2816 14635 2862 14649
rect 2816 14581 2822 14635
rect 2856 14581 2862 14635
rect 2816 14562 2862 14581
rect 3076 18029 6516 18035
rect 3076 17995 3150 18029
rect 3195 17995 3218 18029
rect 3274 17995 3286 18029
rect 3353 17995 3354 18029
rect 3388 17995 3398 18029
rect 3456 17995 3478 18029
rect 3524 17995 3558 18029
rect 3592 17995 3626 18029
rect 3672 17995 3694 18029
rect 3752 17995 3762 18029
rect 3796 17995 3798 18029
rect 3864 17995 3898 18029
rect 3942 17995 3966 18029
rect 4015 17995 4034 18029
rect 4088 17995 4102 18029
rect 4161 17995 4170 18029
rect 4234 17995 4238 18029
rect 4272 17995 4273 18029
rect 4340 17995 4346 18029
rect 4408 17995 4419 18029
rect 4476 17995 4492 18029
rect 4544 17995 4565 18029
rect 4612 17995 4638 18029
rect 4680 17995 4711 18029
rect 4748 17995 4782 18029
rect 4818 17995 4850 18029
rect 4891 17995 4918 18029
rect 4964 17995 4986 18029
rect 5037 17995 5054 18029
rect 5110 17995 5122 18029
rect 5183 17995 5190 18029
rect 5256 17995 5258 18029
rect 5292 17995 5295 18029
rect 5360 17995 5368 18029
rect 5428 17995 5442 18029
rect 5496 17995 5516 18029
rect 5564 17995 5590 18029
rect 5632 17995 5664 18029
rect 5700 17995 5734 18029
rect 5772 17995 5802 18029
rect 5846 17995 5870 18029
rect 5920 17995 5938 18029
rect 5994 17995 6006 18029
rect 6068 17995 6074 18029
rect 6176 17995 6182 18029
rect 6244 17995 6256 18029
rect 6312 17995 6330 18029
rect 6380 17995 6404 18029
rect 6438 17995 6516 18029
rect 3076 17989 6516 17995
rect 3076 17957 3122 17989
rect 3076 17901 3082 17957
rect 3116 17901 3122 17957
rect 3076 17884 3122 17901
rect 3076 17833 3082 17884
rect 3116 17833 3122 17884
rect 3076 17811 3122 17833
rect 3076 17765 3082 17811
rect 3116 17765 3122 17811
rect 3076 17738 3122 17765
rect 6470 17961 6516 17989
rect 6470 17923 6476 17961
rect 6510 17923 6516 17961
rect 6470 17893 6516 17923
rect 6470 17851 6476 17893
rect 6510 17851 6516 17893
rect 6470 17825 6516 17851
rect 6470 17779 6476 17825
rect 6510 17779 6516 17825
rect 6470 17757 6516 17779
rect 3076 17697 3082 17738
rect 3116 17697 3122 17738
rect 3688 17711 3745 17745
rect 3779 17711 3836 17745
rect 6470 17707 6476 17757
rect 6510 17707 6516 17757
rect 3076 17665 3122 17697
rect 3076 17629 3082 17665
rect 3116 17629 3122 17665
rect 3076 17595 3122 17629
rect 3552 17684 3586 17700
rect 3076 17558 3082 17595
rect 3116 17558 3122 17595
rect 3076 17527 3122 17558
rect 3076 17485 3082 17527
rect 3116 17485 3122 17527
rect 3076 17459 3122 17485
rect 3076 17412 3082 17459
rect 3116 17412 3122 17459
rect 3076 17391 3122 17412
rect 3076 17339 3082 17391
rect 3116 17339 3122 17391
rect 3076 17323 3122 17339
rect 3076 17266 3082 17323
rect 3116 17266 3122 17323
rect 3076 17255 3122 17266
rect 3076 17193 3082 17255
rect 3116 17193 3122 17255
rect 3076 17187 3122 17193
rect 3076 17120 3082 17187
rect 3116 17120 3122 17187
rect 3076 17119 3122 17120
rect 3076 17085 3082 17119
rect 3116 17085 3122 17119
rect 3076 17081 3122 17085
rect 3076 17017 3082 17081
rect 3116 17017 3122 17081
rect 3076 17008 3122 17017
rect 3076 16949 3082 17008
rect 3116 16949 3122 17008
rect 3076 16935 3122 16949
rect 3076 16881 3082 16935
rect 3116 16881 3122 16935
rect 3076 16862 3122 16881
rect 3076 16813 3082 16862
rect 3116 16813 3122 16862
rect 3076 16789 3122 16813
rect 3076 16745 3082 16789
rect 3116 16745 3122 16789
rect 3076 16716 3122 16745
rect 3076 16677 3082 16716
rect 3116 16677 3122 16716
rect 3076 16643 3122 16677
rect 3076 16609 3082 16643
rect 3116 16609 3122 16643
rect 3076 16575 3122 16609
rect 3076 16536 3082 16575
rect 3116 16536 3122 16575
rect 3076 16507 3122 16536
rect 3076 16463 3082 16507
rect 3116 16463 3122 16507
rect 3076 16439 3122 16463
rect 3076 16390 3082 16439
rect 3116 16390 3122 16439
rect 3076 16371 3122 16390
rect 3076 16317 3082 16371
rect 3116 16317 3122 16371
rect 3076 16303 3122 16317
rect 3076 16244 3082 16303
rect 3116 16244 3122 16303
rect 3076 16235 3122 16244
rect 3076 16171 3082 16235
rect 3116 16171 3122 16235
rect 3076 16167 3122 16171
rect 3076 16133 3082 16167
rect 3116 16133 3122 16167
rect 3076 16132 3122 16133
rect 3076 16065 3082 16132
rect 3116 16065 3122 16132
rect 3076 16059 3122 16065
rect 3076 15997 3082 16059
rect 3116 15997 3122 16059
rect 3444 17603 3478 17615
rect 3444 17530 3478 17565
rect 3444 17461 3478 17495
rect 3444 17392 3478 17421
rect 3444 17323 3478 17347
rect 3444 17254 3478 17272
rect 3444 17185 3478 17197
rect 3552 17613 3586 17636
rect 6470 17689 6516 17707
rect 6470 17634 6476 17689
rect 6510 17634 6516 17689
rect 6470 17621 6516 17634
rect 3688 17555 3728 17589
rect 6470 17561 6476 17621
rect 6510 17561 6516 17621
rect 3552 17542 3586 17555
rect 3552 17470 3586 17474
rect 3552 17427 3586 17436
rect 6470 17553 6516 17561
rect 6470 17488 6476 17553
rect 6510 17488 6516 17553
rect 6470 17485 6516 17488
rect 6470 17451 6476 17485
rect 6510 17451 6516 17485
rect 6470 17449 6516 17451
rect 3746 17399 3786 17433
rect 3552 17345 3586 17364
rect 3552 17263 3586 17292
rect 6470 17383 6476 17449
rect 6510 17383 6516 17449
rect 6470 17376 6516 17383
rect 6470 17315 6476 17376
rect 6510 17315 6516 17376
rect 6470 17303 6516 17315
rect 3688 17243 3728 17277
rect 6470 17247 6476 17303
rect 6510 17247 6516 17303
rect 3552 17182 3586 17220
rect 3552 17132 3586 17147
rect 6470 17230 6516 17247
rect 6470 17179 6476 17230
rect 6510 17179 6516 17230
rect 6470 17157 6516 17179
rect 3444 17115 3478 17122
rect 3688 17087 3745 17121
rect 3779 17087 3836 17121
rect 6470 17111 6476 17157
rect 6510 17111 6516 17157
rect 3444 17045 3478 17047
rect 3444 17006 3478 17011
rect 6470 17084 6516 17111
rect 6470 17043 6476 17084
rect 6510 17043 6516 17084
rect 6470 17011 6516 17043
rect 3444 16931 3478 16941
rect 3444 16856 3478 16871
rect 6211 16964 6371 16996
rect 6211 16962 6237 16964
rect 6271 16930 6309 16964
rect 6343 16962 6371 16964
rect 6245 16928 6337 16930
rect 6211 16891 6371 16928
rect 4269 16833 4285 16867
rect 4348 16833 4357 16867
rect 4421 16833 4429 16867
rect 4494 16833 4501 16867
rect 4567 16833 4573 16867
rect 4640 16833 4645 16867
rect 4713 16833 4716 16867
rect 4750 16833 4752 16867
rect 4786 16833 4787 16867
rect 4821 16833 4837 16867
rect 4893 16833 4909 16867
rect 4943 16833 4958 16867
rect 5015 16833 5041 16867
rect 5087 16833 5124 16867
rect 5159 16833 5197 16867
rect 5241 16833 5269 16867
rect 5323 16833 5340 16867
rect 5405 16833 5411 16867
rect 5445 16833 5461 16867
rect 6211 16857 6237 16891
rect 6271 16857 6309 16891
rect 6343 16857 6371 16891
rect 3444 16781 3478 16801
rect 6211 16819 6371 16857
rect 6245 16818 6337 16819
rect 6211 16784 6237 16785
rect 6271 16784 6309 16818
rect 6343 16784 6371 16785
rect 6211 16745 6371 16784
rect 3444 16706 3478 16731
rect 3444 16631 3478 16661
rect 3444 16556 3478 16591
rect 3444 16485 3478 16521
rect 3444 16415 3478 16447
rect 3444 16345 3478 16372
rect 3444 16275 3478 16297
rect 3444 16205 3478 16222
rect 3444 16135 3478 16147
rect 3444 16065 3478 16072
rect 3444 16015 3478 16031
rect 3695 16711 3855 16743
rect 3695 16709 3721 16711
rect 3827 16709 3855 16711
rect 3695 16564 3721 16675
rect 3827 16564 3855 16675
rect 3695 16419 3721 16530
rect 3827 16419 3855 16530
rect 3695 16274 3721 16385
rect 3827 16274 3855 16385
rect 3695 16129 3721 16240
rect 3827 16129 3855 16240
rect 3729 16095 3821 16101
rect 6211 16711 6237 16745
rect 6271 16711 6309 16745
rect 6343 16711 6371 16745
rect 6211 16676 6371 16711
rect 6245 16672 6337 16676
rect 6211 16638 6237 16642
rect 6271 16638 6309 16672
rect 6343 16638 6371 16642
rect 6211 16599 6371 16638
rect 6211 16565 6237 16599
rect 6271 16565 6309 16599
rect 6343 16565 6371 16599
rect 6211 16533 6371 16565
rect 6245 16525 6337 16533
rect 6211 16491 6237 16499
rect 6271 16491 6309 16525
rect 6343 16491 6371 16499
rect 6211 16451 6371 16491
rect 6211 16417 6237 16451
rect 6271 16417 6309 16451
rect 6343 16417 6371 16451
rect 6211 16390 6371 16417
rect 6245 16377 6337 16390
rect 6211 16343 6237 16356
rect 6271 16343 6309 16377
rect 6343 16343 6371 16356
rect 6211 16303 6371 16343
rect 6211 16269 6237 16303
rect 6271 16269 6309 16303
rect 6343 16269 6371 16303
rect 6211 16247 6371 16269
rect 6245 16229 6337 16247
rect 6211 16195 6237 16213
rect 6271 16195 6309 16229
rect 6343 16195 6371 16213
rect 6211 16155 6371 16195
rect 6211 16121 6237 16155
rect 6271 16121 6309 16155
rect 6343 16121 6371 16155
rect 6211 16104 6371 16121
rect 3695 16062 3855 16095
rect 3695 16028 3721 16062
rect 3755 16028 3793 16062
rect 3827 16028 3855 16062
rect 4235 16061 4251 16095
rect 4316 16061 4320 16095
rect 4354 16061 4355 16095
rect 4423 16061 4428 16095
rect 4492 16061 4501 16095
rect 4561 16061 4574 16095
rect 4630 16061 4647 16095
rect 4699 16061 4720 16095
rect 4769 16061 4793 16095
rect 4839 16061 4866 16095
rect 4909 16061 4939 16095
rect 4979 16061 5012 16095
rect 5049 16061 5085 16095
rect 5119 16061 5155 16095
rect 5192 16061 5225 16095
rect 5265 16061 5295 16095
rect 5338 16061 5365 16095
rect 5411 16061 5435 16095
rect 5484 16061 5505 16095
rect 5557 16061 5575 16095
rect 5630 16061 5645 16095
rect 5703 16061 5715 16095
rect 5776 16061 5785 16095
rect 5819 16061 5835 16095
rect 6245 16081 6337 16104
rect 3076 15986 3122 15997
rect 3076 15929 3082 15986
rect 3116 15929 3122 15986
rect 3076 15913 3122 15929
rect 3076 15861 3082 15913
rect 3116 15861 3122 15913
rect 3076 15840 3122 15861
rect 3076 15793 3082 15840
rect 3116 15793 3122 15840
rect 3076 15767 3122 15793
rect 3076 15725 3082 15767
rect 3116 15725 3122 15767
rect 3076 15694 3122 15725
rect 3076 15657 3082 15694
rect 3116 15657 3122 15694
rect 3076 15623 3122 15657
rect 3076 15587 3082 15623
rect 3116 15587 3122 15623
rect 3076 15555 3122 15587
rect 3076 15514 3082 15555
rect 3116 15514 3122 15555
rect 3076 15487 3122 15514
rect 3076 15441 3082 15487
rect 3116 15441 3122 15487
rect 3076 15419 3122 15441
rect 3076 15368 3082 15419
rect 3116 15368 3122 15419
rect 3076 15351 3122 15368
rect 3076 15295 3082 15351
rect 3116 15295 3122 15351
rect 3076 15283 3122 15295
rect 3076 15222 3082 15283
rect 3116 15222 3122 15283
rect 3076 15215 3122 15222
rect 3076 15149 3082 15215
rect 3116 15149 3122 15215
rect 3076 15147 3122 15149
rect 3076 15113 3082 15147
rect 3116 15113 3122 15147
rect 3076 15110 3122 15113
rect 3076 15045 3082 15110
rect 3116 15045 3122 15110
rect 3076 15037 3122 15045
rect 3076 14977 3082 15037
rect 3116 14977 3122 15037
rect 3076 14964 3122 14977
rect 3076 14909 3082 14964
rect 3116 14909 3122 14964
rect 3076 14891 3122 14909
rect 3076 14841 3082 14891
rect 3116 14841 3122 14891
rect 3076 14819 3122 14841
rect 3076 14773 3082 14819
rect 3116 14773 3122 14819
rect 3076 14747 3122 14773
rect 3076 14705 3082 14747
rect 3116 14705 3122 14747
rect 3076 14675 3122 14705
rect 3076 14637 3082 14675
rect 3116 14637 3122 14675
rect 3076 14609 3122 14637
rect 3695 15989 3855 16028
rect 3695 15984 3721 15989
rect 3755 15955 3793 15989
rect 3827 15984 3855 15989
rect 3729 15950 3821 15955
rect 3695 15916 3855 15950
rect 3695 15882 3721 15916
rect 3755 15882 3793 15916
rect 3827 15882 3855 15916
rect 3695 15843 3855 15882
rect 3695 15839 3721 15843
rect 3755 15809 3793 15843
rect 3827 15839 3855 15843
rect 3729 15805 3821 15809
rect 3695 15770 3855 15805
rect 3695 15736 3721 15770
rect 3755 15736 3793 15770
rect 3827 15736 3855 15770
rect 3695 15697 3855 15736
rect 3695 15693 3721 15697
rect 3755 15663 3793 15697
rect 3827 15693 3855 15697
rect 3729 15659 3821 15663
rect 3695 15624 3855 15659
rect 3695 15590 3721 15624
rect 3755 15590 3793 15624
rect 3827 15590 3855 15624
rect 3695 15551 3855 15590
rect 3695 15547 3721 15551
rect 3755 15517 3793 15551
rect 3827 15547 3855 15551
rect 3729 15513 3821 15517
rect 3695 15478 3855 15513
rect 3695 15444 3721 15478
rect 3755 15444 3793 15478
rect 3827 15444 3855 15478
rect 3695 15405 3855 15444
rect 3695 15401 3721 15405
rect 3755 15371 3793 15405
rect 3827 15401 3855 15405
rect 3729 15367 3821 15371
rect 3695 15332 3855 15367
rect 6211 16047 6237 16070
rect 6271 16047 6309 16081
rect 6343 16047 6371 16070
rect 6211 16007 6371 16047
rect 6211 15973 6237 16007
rect 6271 15973 6309 16007
rect 6343 15973 6371 16007
rect 6211 15961 6371 15973
rect 6245 15933 6337 15961
rect 6211 15899 6237 15927
rect 6271 15899 6309 15933
rect 6343 15899 6371 15927
rect 6211 15859 6371 15899
rect 6211 15825 6237 15859
rect 6271 15825 6309 15859
rect 6343 15825 6371 15859
rect 6211 15818 6371 15825
rect 6245 15785 6337 15818
rect 6211 15751 6237 15784
rect 6271 15751 6309 15785
rect 6343 15751 6371 15784
rect 6211 15711 6371 15751
rect 6211 15677 6237 15711
rect 6271 15677 6309 15711
rect 6343 15677 6371 15711
rect 6211 15675 6371 15677
rect 6245 15641 6337 15675
rect 6211 15637 6371 15641
rect 6211 15603 6237 15637
rect 6271 15603 6309 15637
rect 6343 15603 6371 15637
rect 6211 15563 6371 15603
rect 6211 15532 6237 15563
rect 6271 15529 6309 15563
rect 6343 15532 6371 15563
rect 6245 15498 6337 15529
rect 6211 15489 6371 15498
rect 6211 15455 6237 15489
rect 6271 15455 6309 15489
rect 6343 15455 6371 15489
rect 6211 15415 6371 15455
rect 6211 15389 6237 15415
rect 6271 15381 6309 15415
rect 6343 15389 6371 15415
rect 3695 15298 3721 15332
rect 3755 15298 3793 15332
rect 3827 15298 3855 15332
rect 4235 15331 4251 15365
rect 4316 15331 4320 15365
rect 4354 15331 4355 15365
rect 4423 15331 4428 15365
rect 4492 15331 4501 15365
rect 4561 15331 4574 15365
rect 4630 15331 4647 15365
rect 4699 15331 4720 15365
rect 4769 15331 4793 15365
rect 4839 15331 4866 15365
rect 4909 15331 4939 15365
rect 4979 15331 5012 15365
rect 5049 15331 5085 15365
rect 5119 15331 5155 15365
rect 5192 15331 5225 15365
rect 5265 15331 5295 15365
rect 5338 15331 5365 15365
rect 5411 15331 5435 15365
rect 5484 15331 5505 15365
rect 5557 15331 5575 15365
rect 5630 15331 5645 15365
rect 5703 15331 5715 15365
rect 5776 15331 5785 15365
rect 5819 15331 5835 15365
rect 6245 15355 6337 15381
rect 6211 15341 6371 15355
rect 3695 15259 3855 15298
rect 3695 15255 3721 15259
rect 3755 15225 3793 15259
rect 3827 15255 3855 15259
rect 3729 15221 3821 15225
rect 3695 15186 3855 15221
rect 3695 15152 3721 15186
rect 3755 15152 3793 15186
rect 3827 15152 3855 15186
rect 3695 15113 3855 15152
rect 3695 15109 3721 15113
rect 3755 15079 3793 15113
rect 3827 15109 3855 15113
rect 3729 15075 3821 15079
rect 3695 15040 3855 15075
rect 3695 15006 3721 15040
rect 3755 15006 3793 15040
rect 3827 15006 3855 15040
rect 3695 14967 3855 15006
rect 3695 14963 3721 14967
rect 3755 14933 3793 14967
rect 3827 14963 3855 14967
rect 3729 14929 3821 14933
rect 3695 14894 3855 14929
rect 3695 14860 3721 14894
rect 3755 14860 3793 14894
rect 3827 14860 3855 14894
rect 3695 14821 3855 14860
rect 3695 14817 3721 14821
rect 3755 14787 3793 14821
rect 3827 14817 3855 14821
rect 3729 14783 3821 14787
rect 3695 14748 3855 14783
rect 3695 14714 3721 14748
rect 3755 14714 3793 14748
rect 3827 14714 3855 14748
rect 3695 14675 3855 14714
rect 3695 14671 3721 14675
rect 3755 14641 3793 14675
rect 3827 14671 3855 14675
rect 3729 14637 3821 14641
rect 3695 14609 3855 14637
rect 6211 15307 6237 15341
rect 6271 15307 6309 15341
rect 6343 15307 6371 15341
rect 6211 15267 6371 15307
rect 6211 15246 6237 15267
rect 6271 15233 6309 15267
rect 6343 15246 6371 15267
rect 6245 15212 6337 15233
rect 6211 15193 6371 15212
rect 6211 15159 6237 15193
rect 6271 15159 6309 15193
rect 6343 15159 6371 15193
rect 6211 15119 6371 15159
rect 6211 15103 6237 15119
rect 6271 15085 6309 15119
rect 6343 15103 6371 15119
rect 6245 15069 6337 15085
rect 6211 15045 6371 15069
rect 6211 15011 6237 15045
rect 6271 15011 6309 15045
rect 6343 15011 6371 15045
rect 6211 14971 6371 15011
rect 6211 14959 6237 14971
rect 6271 14937 6309 14971
rect 6343 14959 6371 14971
rect 6245 14925 6337 14937
rect 6211 14897 6371 14925
rect 6211 14863 6237 14897
rect 6271 14863 6309 14897
rect 6343 14863 6371 14897
rect 6211 14823 6371 14863
rect 6211 14815 6237 14823
rect 6271 14789 6309 14823
rect 6343 14815 6371 14823
rect 6245 14781 6337 14789
rect 6211 14749 6371 14781
rect 6211 14715 6237 14749
rect 6271 14715 6309 14749
rect 6343 14715 6371 14749
rect 6211 14675 6371 14715
rect 6211 14671 6237 14675
rect 6343 14671 6371 14675
rect 6211 14609 6237 14637
rect 3076 14603 6237 14609
rect 6343 14609 6371 14637
rect 6470 16975 6476 17011
rect 6510 16975 6516 17011
rect 6470 16941 6516 16975
rect 6470 16904 6476 16941
rect 6510 16904 6516 16941
rect 6470 16873 6516 16904
rect 6470 16831 6476 16873
rect 6510 16831 6516 16873
rect 6470 16805 6516 16831
rect 6470 16758 6476 16805
rect 6510 16758 6516 16805
rect 6470 16737 6516 16758
rect 6470 16685 6476 16737
rect 6510 16685 6516 16737
rect 6470 16669 6516 16685
rect 6470 16612 6476 16669
rect 6510 16612 6516 16669
rect 6470 16601 6516 16612
rect 6470 16539 6476 16601
rect 6510 16539 6516 16601
rect 6470 16533 6516 16539
rect 6470 16466 6476 16533
rect 6510 16466 6516 16533
rect 6470 16465 6516 16466
rect 6470 16431 6476 16465
rect 6510 16431 6516 16465
rect 6470 16427 6516 16431
rect 6470 16363 6476 16427
rect 6510 16363 6516 16427
rect 6470 16354 6516 16363
rect 6470 16295 6476 16354
rect 6510 16295 6516 16354
rect 6470 16281 6516 16295
rect 6470 16227 6476 16281
rect 6510 16227 6516 16281
rect 6470 16208 6516 16227
rect 6470 16159 6476 16208
rect 6510 16159 6516 16208
rect 6470 16135 6516 16159
rect 6470 16091 6476 16135
rect 6510 16091 6516 16135
rect 6470 16062 6516 16091
rect 6470 16023 6476 16062
rect 6510 16023 6516 16062
rect 6470 15989 6516 16023
rect 6470 15955 6476 15989
rect 6510 15955 6516 15989
rect 6470 15921 6516 15955
rect 6470 15882 6476 15921
rect 6510 15882 6516 15921
rect 6470 15853 6516 15882
rect 6470 15809 6476 15853
rect 6510 15809 6516 15853
rect 6470 15785 6516 15809
rect 6470 15736 6476 15785
rect 6510 15736 6516 15785
rect 6470 15717 6516 15736
rect 6470 15663 6476 15717
rect 6510 15663 6516 15717
rect 6470 15649 6516 15663
rect 6470 15590 6476 15649
rect 6510 15590 6516 15649
rect 6470 15581 6516 15590
rect 6470 15517 6476 15581
rect 6510 15517 6516 15581
rect 6470 15513 6516 15517
rect 6470 15479 6476 15513
rect 6510 15479 6516 15513
rect 6470 15478 6516 15479
rect 6470 15411 6476 15478
rect 6510 15411 6516 15478
rect 6470 15405 6516 15411
rect 6470 15343 6476 15405
rect 6510 15343 6516 15405
rect 6470 15332 6516 15343
rect 6470 15275 6476 15332
rect 6510 15275 6516 15332
rect 6470 15259 6516 15275
rect 6470 15207 6476 15259
rect 6510 15207 6516 15259
rect 6470 15186 6516 15207
rect 6470 15139 6476 15186
rect 6510 15139 6516 15186
rect 6470 15113 6516 15139
rect 6470 15071 6476 15113
rect 6510 15071 6516 15113
rect 6470 15040 6516 15071
rect 6470 15003 6476 15040
rect 6510 15003 6516 15040
rect 6470 14969 6516 15003
rect 6470 14933 6476 14969
rect 6510 14933 6516 14969
rect 6470 14901 6516 14933
rect 6470 14860 6476 14901
rect 6510 14860 6516 14901
rect 6470 14833 6516 14860
rect 6470 14787 6476 14833
rect 6510 14787 6516 14833
rect 6470 14765 6516 14787
rect 6470 14714 6476 14765
rect 6510 14714 6516 14765
rect 6470 14697 6516 14714
rect 6470 14641 6476 14697
rect 6510 14641 6516 14697
rect 6470 14609 6516 14641
rect 6343 14603 6516 14609
rect 3076 14569 3154 14603
rect 3188 14569 3212 14603
rect 3261 14569 3280 14603
rect 3334 14569 3348 14603
rect 3407 14569 3416 14603
rect 3480 14569 3484 14603
rect 3518 14569 3519 14603
rect 3586 14569 3592 14603
rect 3654 14569 3665 14603
rect 3722 14569 3738 14603
rect 3790 14569 3811 14603
rect 3858 14569 3884 14603
rect 3926 14569 3956 14603
rect 3994 14569 4028 14603
rect 4062 14569 4096 14603
rect 4134 14569 4164 14603
rect 4206 14569 4232 14603
rect 4278 14569 4300 14603
rect 4350 14569 4368 14603
rect 4422 14569 4436 14603
rect 4494 14569 4504 14603
rect 4566 14569 4572 14603
rect 4638 14569 4640 14603
rect 4674 14569 4676 14603
rect 4742 14569 4748 14603
rect 4810 14569 4820 14603
rect 4878 14569 4892 14603
rect 4946 14569 4964 14603
rect 5014 14569 5036 14603
rect 5082 14569 5108 14603
rect 5150 14569 5180 14603
rect 5218 14569 5252 14603
rect 5286 14569 5320 14603
rect 5358 14569 5388 14603
rect 5430 14569 5456 14603
rect 5502 14569 5524 14603
rect 5574 14569 5592 14603
rect 5646 14569 5660 14603
rect 5718 14569 5728 14603
rect 5790 14569 5796 14603
rect 5862 14569 5864 14603
rect 5898 14569 5900 14603
rect 5966 14569 5972 14603
rect 6034 14569 6044 14603
rect 6102 14569 6116 14603
rect 6170 14569 6188 14603
rect 6374 14569 6404 14603
rect 6442 14569 6516 14603
rect 3076 14563 6516 14569
rect 6744 18017 6790 18036
rect 6744 17963 6750 18017
rect 6784 17963 6790 18017
rect 6744 17949 6790 17963
rect 6744 17890 6750 17949
rect 6784 17890 6790 17949
rect 6744 17881 6790 17890
rect 6744 17817 6750 17881
rect 6784 17817 6790 17881
rect 6744 17813 6790 17817
rect 6744 17779 6750 17813
rect 6784 17779 6790 17813
rect 6744 17778 6790 17779
rect 6744 17711 6750 17778
rect 6784 17711 6790 17778
rect 6744 17705 6790 17711
rect 6744 17643 6750 17705
rect 6784 17643 6790 17705
rect 6744 17632 6790 17643
rect 6744 17575 6750 17632
rect 6784 17575 6790 17632
rect 6744 17559 6790 17575
rect 6744 17507 6750 17559
rect 6784 17507 6790 17559
rect 6744 17486 6790 17507
rect 6744 17439 6750 17486
rect 6784 17439 6790 17486
rect 6744 17413 6790 17439
rect 6744 17371 6750 17413
rect 6784 17371 6790 17413
rect 6744 17340 6790 17371
rect 6744 17303 6750 17340
rect 6784 17303 6790 17340
rect 6744 17269 6790 17303
rect 6744 17233 6750 17269
rect 6784 17233 6790 17269
rect 6744 17201 6790 17233
rect 6744 17160 6750 17201
rect 6784 17160 6790 17201
rect 6744 17133 6790 17160
rect 6744 17087 6750 17133
rect 6784 17087 6790 17133
rect 6744 17065 6790 17087
rect 6744 17014 6750 17065
rect 6784 17014 6790 17065
rect 6744 16997 6790 17014
rect 6744 16941 6750 16997
rect 6784 16941 6790 16997
rect 6744 16929 6790 16941
rect 6744 16868 6750 16929
rect 6784 16868 6790 16929
rect 6744 16861 6790 16868
rect 6744 16795 6750 16861
rect 6784 16795 6790 16861
rect 6744 16793 6790 16795
rect 6744 16759 6750 16793
rect 6784 16759 6790 16793
rect 6744 16756 6790 16759
rect 6744 16691 6750 16756
rect 6784 16691 6790 16756
rect 6744 16683 6790 16691
rect 6744 16623 6750 16683
rect 6784 16623 6790 16683
rect 6744 16610 6790 16623
rect 6744 16555 6750 16610
rect 6784 16555 6790 16610
rect 6744 16537 6790 16555
rect 6744 16487 6750 16537
rect 6784 16487 6790 16537
rect 6744 16464 6790 16487
rect 6744 16419 6750 16464
rect 6784 16419 6790 16464
rect 6744 16391 6790 16419
rect 6744 16351 6750 16391
rect 6784 16351 6790 16391
rect 6744 16318 6790 16351
rect 6744 16283 6750 16318
rect 6784 16283 6790 16318
rect 6744 16249 6790 16283
rect 6744 16211 6750 16249
rect 6784 16211 6790 16249
rect 6744 16181 6790 16211
rect 6744 16138 6750 16181
rect 6784 16138 6790 16181
rect 6744 16113 6790 16138
rect 6744 16065 6750 16113
rect 6784 16065 6790 16113
rect 6744 16045 6790 16065
rect 6744 15992 6750 16045
rect 6784 15992 6790 16045
rect 6744 15977 6790 15992
rect 6744 15919 6750 15977
rect 6784 15919 6790 15977
rect 6744 15909 6790 15919
rect 6744 15846 6750 15909
rect 6784 15846 6790 15909
rect 6744 15841 6790 15846
rect 6744 15739 6750 15841
rect 6784 15739 6790 15841
rect 6744 15734 6790 15739
rect 6744 15671 6750 15734
rect 6784 15671 6790 15734
rect 6744 15661 6790 15671
rect 6744 15603 6750 15661
rect 6784 15603 6790 15661
rect 6744 15588 6790 15603
rect 6744 15535 6750 15588
rect 6784 15535 6790 15588
rect 6744 15515 6790 15535
rect 6744 15467 6750 15515
rect 6784 15467 6790 15515
rect 6744 15442 6790 15467
rect 6744 15399 6750 15442
rect 6784 15399 6790 15442
rect 6744 15369 6790 15399
rect 6744 15331 6750 15369
rect 6784 15331 6790 15369
rect 6744 15297 6790 15331
rect 6744 15262 6750 15297
rect 6784 15262 6790 15297
rect 6744 15229 6790 15262
rect 6744 15189 6750 15229
rect 6784 15189 6790 15229
rect 6744 15161 6790 15189
rect 6744 15116 6750 15161
rect 6784 15116 6790 15161
rect 6744 15093 6790 15116
rect 6744 15043 6750 15093
rect 6784 15043 6790 15093
rect 6744 15025 6790 15043
rect 6744 14970 6750 15025
rect 6784 14970 6790 15025
rect 6744 14957 6790 14970
rect 6744 14897 6750 14957
rect 6784 14897 6790 14957
rect 6744 14889 6790 14897
rect 6744 14824 6750 14889
rect 6784 14824 6790 14889
rect 6744 14821 6790 14824
rect 6744 14787 6750 14821
rect 6784 14787 6790 14821
rect 6744 14785 6790 14787
rect 6744 14719 6750 14785
rect 6784 14719 6790 14785
rect 6744 14711 6790 14719
rect 6744 14651 6750 14711
rect 6784 14651 6790 14711
rect 6744 14637 6790 14651
rect 6744 14583 6750 14637
rect 6784 14583 6790 14637
rect 6744 14563 6790 14583
rect 2816 14513 2822 14562
rect 2856 14513 2862 14562
rect 2816 14489 2862 14513
rect 2816 14445 2822 14489
rect 2856 14445 2862 14489
rect 2816 14416 2862 14445
rect 2816 14377 2822 14416
rect 2856 14377 2862 14416
rect 2816 14349 2862 14377
rect 6744 14515 6750 14563
rect 6784 14515 6790 14563
rect 6744 14489 6790 14515
rect 6744 14447 6750 14489
rect 6784 14447 6790 14489
rect 6744 14415 6790 14447
rect 6744 14379 6750 14415
rect 6784 14379 6790 14415
rect 6744 14349 6790 14379
rect 2816 14343 6790 14349
rect 2816 14309 2894 14343
rect 2928 14309 2942 14343
rect 3001 14309 3010 14343
rect 3074 14309 3078 14343
rect 3112 14309 3113 14343
rect 3180 14309 3186 14343
rect 3248 14309 3259 14343
rect 3316 14309 3332 14343
rect 3384 14309 3405 14343
rect 3452 14309 3478 14343
rect 3520 14309 3551 14343
rect 3588 14309 3622 14343
rect 3658 14309 3690 14343
rect 3731 14309 3758 14343
rect 3804 14309 3826 14343
rect 3877 14309 3894 14343
rect 3950 14309 3962 14343
rect 4023 14309 4030 14343
rect 4096 14309 4098 14343
rect 4132 14309 4135 14343
rect 4200 14309 4208 14343
rect 4268 14309 4281 14343
rect 4336 14309 4354 14343
rect 4404 14309 4427 14343
rect 4472 14309 4500 14343
rect 4540 14309 4573 14343
rect 4608 14309 4642 14343
rect 4680 14309 4710 14343
rect 4753 14309 4778 14343
rect 4826 14309 4846 14343
rect 4899 14309 4914 14343
rect 4972 14309 4982 14343
rect 5045 14309 5050 14343
rect 5152 14309 5157 14343
rect 5220 14309 5230 14343
rect 5288 14309 5303 14343
rect 5356 14309 5376 14343
rect 5424 14309 5449 14343
rect 5492 14309 5522 14343
rect 5560 14309 5594 14343
rect 5629 14309 5662 14343
rect 5702 14309 5730 14343
rect 5775 14309 5798 14343
rect 5848 14309 5866 14343
rect 5920 14309 5934 14343
rect 5992 14309 6002 14343
rect 6064 14309 6070 14343
rect 6136 14309 6138 14343
rect 6172 14309 6174 14343
rect 6240 14309 6246 14343
rect 6308 14309 6318 14343
rect 6376 14309 6390 14343
rect 6444 14309 6462 14343
rect 6512 14309 6534 14343
rect 6580 14309 6606 14343
rect 6648 14309 6678 14343
rect 6716 14309 6790 14343
rect 2816 14303 6790 14309
<< viali >>
rect 2897 39840 2918 39874
rect 2918 39840 2931 39874
rect 2972 39840 2986 39874
rect 2986 39840 3006 39874
rect 3047 39840 3054 39874
rect 3054 39840 3081 39874
rect 3123 39840 3156 39874
rect 3156 39840 3157 39874
rect 3199 39840 3224 39874
rect 3224 39840 3233 39874
rect 3275 39840 3292 39874
rect 3292 39840 3309 39874
rect 3351 39840 3360 39874
rect 3360 39840 3385 39874
rect 3427 39840 3428 39874
rect 3428 39840 3461 39874
rect 3503 39840 3530 39874
rect 3530 39840 3537 39874
rect 3579 39840 3598 39874
rect 3598 39840 3613 39874
rect 3655 39840 3666 39874
rect 3666 39840 3689 39874
rect 3731 39840 3734 39874
rect 3734 39840 3765 39874
rect 3807 39840 3836 39874
rect 3836 39840 3841 39874
rect 3883 39840 3904 39874
rect 3904 39840 3917 39874
rect 3959 39840 3972 39874
rect 3972 39840 3993 39874
rect 4035 39840 4040 39874
rect 4040 39840 4069 39874
rect 4111 39840 4142 39874
rect 4142 39840 4145 39874
rect 4221 39840 4244 39874
rect 4244 39840 4255 39874
rect 4294 39840 4312 39874
rect 4312 39840 4328 39874
rect 4367 39840 4380 39874
rect 4380 39840 4401 39874
rect 4440 39840 4448 39874
rect 4448 39840 4474 39874
rect 4513 39840 4516 39874
rect 4516 39840 4547 39874
rect 4586 39840 4618 39874
rect 4618 39840 4620 39874
rect 4659 39840 4686 39874
rect 4686 39840 4693 39874
rect 4732 39840 4754 39874
rect 4754 39840 4766 39874
rect 4805 39840 4822 39874
rect 4822 39840 4839 39874
rect 4878 39840 4890 39874
rect 4890 39840 4912 39874
rect 4951 39840 4958 39874
rect 4958 39840 4985 39874
rect 5024 39840 5026 39874
rect 5026 39840 5058 39874
rect 5097 39840 5128 39874
rect 5128 39840 5131 39874
rect 5170 39840 5196 39874
rect 5196 39840 5204 39874
rect 5243 39840 5264 39874
rect 5264 39840 5277 39874
rect 5316 39840 5332 39874
rect 5332 39840 5350 39874
rect 5389 39840 5400 39874
rect 5400 39840 5423 39874
rect 5462 39840 5468 39874
rect 5468 39840 5496 39874
rect 5535 39840 5536 39874
rect 5536 39840 5569 39874
rect 5608 39840 5638 39874
rect 5638 39840 5642 39874
rect 5681 39840 5706 39874
rect 5706 39840 5715 39874
rect 5754 39840 5774 39874
rect 5774 39840 5788 39874
rect 5827 39840 5842 39874
rect 5842 39840 5861 39874
rect 5900 39840 5910 39874
rect 5910 39840 5934 39874
rect 5973 39840 5978 39874
rect 5978 39840 6007 39874
rect 6046 39840 6080 39874
rect 6120 39840 6148 39874
rect 6148 39840 6154 39874
rect 6194 39840 6216 39874
rect 6216 39840 6228 39874
rect 6268 39840 6284 39874
rect 6284 39840 6302 39874
rect 6342 39840 6352 39874
rect 6352 39840 6376 39874
rect 6416 39840 6420 39874
rect 6420 39840 6450 39874
rect 6490 39840 6522 39874
rect 6522 39840 6524 39874
rect 6564 39840 6590 39874
rect 6590 39840 6598 39874
rect 6638 39840 6658 39874
rect 6658 39840 6672 39874
rect 6712 39840 6726 39874
rect 6726 39840 6746 39874
rect 6786 39840 6794 39874
rect 6794 39840 6820 39874
rect 6860 39840 6862 39874
rect 6862 39840 6894 39874
rect 6934 39840 6964 39874
rect 6964 39840 6968 39874
rect 7008 39840 7032 39874
rect 7032 39840 7042 39874
rect 7082 39840 7100 39874
rect 7100 39840 7116 39874
rect 7156 39840 7168 39874
rect 7168 39840 7190 39874
rect 7230 39840 7236 39874
rect 7236 39840 7264 39874
rect 7304 39840 7338 39874
rect 7378 39840 7406 39874
rect 7406 39840 7412 39874
rect 7452 39840 7474 39874
rect 7474 39840 7486 39874
rect 7526 39840 7542 39874
rect 7542 39840 7560 39874
rect 7600 39840 7610 39874
rect 7610 39840 7634 39874
rect 7674 39840 7678 39874
rect 7678 39840 7708 39874
rect 2822 39772 2856 39802
rect 2822 39768 2856 39772
rect 2822 39704 2856 39729
rect 2822 39695 2856 39704
rect 2822 39636 2856 39656
rect 2822 39622 2856 39636
rect 7746 39768 7780 39802
rect 7746 39700 7780 39730
rect 7746 39696 7780 39700
rect 7746 39632 7780 39658
rect 7746 39624 7780 39632
rect 2822 39568 2856 39583
rect 2822 39549 2856 39568
rect 2822 39500 2856 39510
rect 2822 39476 2856 39500
rect 2822 39432 2856 39437
rect 2822 39403 2856 39432
rect 2822 39330 2856 39364
rect 2822 39262 2856 39291
rect 2822 39257 2856 39262
rect 2822 39194 2856 39218
rect 2822 39184 2856 39194
rect 2822 39126 2856 39145
rect 2822 39111 2856 39126
rect 2822 39058 2856 39072
rect 2822 39038 2856 39058
rect 2822 38990 2856 38999
rect 2822 38965 2856 38990
rect 2822 38922 2856 38926
rect 2822 38892 2856 38922
rect 2822 38820 2856 38853
rect 2822 38819 2856 38820
rect 2822 38752 2856 38780
rect 2822 38746 2856 38752
rect 2822 38684 2856 38707
rect 2822 38673 2856 38684
rect 2822 38616 2856 38634
rect 2822 38600 2856 38616
rect 2822 38548 2856 38561
rect 2822 38527 2856 38548
rect 2822 38480 2856 38488
rect 2822 38454 2856 38480
rect 2822 38412 2856 38415
rect 2822 38381 2856 38412
rect 2822 38310 2856 38342
rect 2822 38308 2856 38310
rect 2822 38242 2856 38269
rect 2822 38235 2856 38242
rect 2822 38174 2856 38196
rect 2822 38162 2856 38174
rect 2822 38106 2856 38123
rect 2822 38089 2856 38106
rect 2822 38038 2856 38050
rect 2822 38016 2856 38038
rect 2822 37970 2856 37977
rect 2822 37943 2856 37970
rect 2822 37902 2856 37904
rect 2822 37870 2856 37902
rect 2822 37800 2856 37831
rect 2822 37797 2856 37800
rect 2822 37732 2856 37758
rect 2822 37724 2856 37732
rect 2822 37664 2856 37685
rect 2822 37651 2856 37664
rect 2822 37596 2856 37612
rect 2822 37578 2856 37596
rect 2822 37528 2856 37539
rect 2822 37505 2856 37528
rect 2822 37460 2856 37466
rect 2822 37432 2856 37460
rect 2822 37392 2856 37393
rect 2822 37359 2856 37392
rect 2822 37290 2856 37320
rect 2822 37286 2856 37290
rect 2822 37222 2856 37247
rect 2822 37213 2856 37222
rect 2822 37154 2856 37174
rect 2822 37140 2856 37154
rect 2822 37086 2856 37102
rect 2822 37068 2856 37086
rect 2822 37018 2856 37030
rect 2822 36996 2856 37018
rect 2822 36950 2856 36958
rect 2822 36924 2856 36950
rect 2822 36882 2856 36886
rect 2822 36852 2856 36882
rect 2822 36780 2856 36814
rect 2822 36712 2856 36742
rect 2822 36708 2856 36712
rect 2822 36644 2856 36670
rect 2822 36636 2856 36644
rect 2822 36576 2856 36598
rect 2822 36564 2856 36576
rect 2822 36508 2856 36526
rect 2822 36492 2856 36508
rect 2822 36440 2856 36454
rect 2822 36420 2856 36440
rect 2822 36372 2856 36382
rect 2822 36348 2856 36372
rect 2822 36304 2856 36310
rect 2822 36276 2856 36304
rect 2822 36236 2856 36238
rect 2822 36204 2856 36236
rect 2822 36134 2856 36166
rect 2822 36132 2856 36134
rect 2822 36066 2856 36094
rect 2822 36060 2856 36066
rect 2822 35998 2856 36022
rect 2822 35988 2856 35998
rect 2822 35930 2856 35950
rect 2822 35916 2856 35930
rect 2822 35862 2856 35878
rect 2822 35844 2856 35862
rect 2822 35794 2856 35806
rect 2822 35772 2856 35794
rect 2822 35726 2856 35734
rect 2822 35700 2856 35726
rect 2822 35658 2856 35662
rect 2822 35628 2856 35658
rect 2822 35556 2856 35590
rect 2822 35488 2856 35518
rect 2822 35484 2856 35488
rect 2822 35420 2856 35446
rect 2822 35412 2856 35420
rect 2822 35352 2856 35374
rect 2822 35340 2856 35352
rect 2822 35284 2856 35302
rect 2822 35268 2856 35284
rect 2822 35216 2856 35230
rect 2822 35196 2856 35216
rect 2822 35148 2856 35158
rect 2822 35124 2856 35148
rect 2822 35080 2856 35086
rect 2822 35052 2856 35080
rect 2822 35012 2856 35014
rect 2822 34980 2856 35012
rect 2822 34910 2856 34942
rect 2822 34908 2856 34910
rect 2822 34842 2856 34870
rect 2822 34836 2856 34842
rect 2822 34774 2856 34798
rect 2822 34764 2856 34774
rect 2822 34706 2856 34726
rect 2822 34692 2856 34706
rect 2822 34638 2856 34654
rect 2822 34620 2856 34638
rect 2822 34570 2856 34582
rect 2822 34548 2856 34570
rect 2822 34502 2856 34510
rect 2822 34476 2856 34502
rect 2822 34434 2856 34438
rect 2822 34404 2856 34434
rect 2822 34332 2856 34366
rect 2822 34264 2856 34294
rect 2822 34260 2856 34264
rect 2822 34196 2856 34222
rect 2822 34188 2856 34196
rect 2822 34128 2856 34150
rect 2822 34116 2856 34128
rect 2822 34060 2856 34078
rect 2822 34044 2856 34060
rect 2822 33992 2856 34006
rect 2822 33972 2856 33992
rect 2822 33924 2856 33934
rect 2822 33900 2856 33924
rect 2822 33856 2856 33862
rect 2822 33828 2856 33856
rect 2822 33788 2856 33790
rect 2822 33756 2856 33788
rect 2822 33686 2856 33718
rect 2822 33684 2856 33686
rect 2822 33618 2856 33646
rect 2822 33612 2856 33618
rect 2822 33550 2856 33574
rect 2822 33540 2856 33550
rect 2822 33482 2856 33502
rect 2822 33468 2856 33482
rect 2822 33414 2856 33430
rect 2822 33396 2856 33414
rect 2822 33346 2856 33358
rect 2822 33324 2856 33346
rect 2822 33278 2856 33286
rect 2822 33252 2856 33278
rect 2822 33210 2856 33214
rect 2822 33180 2856 33210
rect 2822 33108 2856 33142
rect 2822 33040 2856 33070
rect 2822 33036 2856 33040
rect 2822 32972 2856 32998
rect 2822 32964 2856 32972
rect 2822 32904 2856 32926
rect 2822 32892 2856 32904
rect 2822 32836 2856 32854
rect 2822 32820 2856 32836
rect 2822 32768 2856 32782
rect 2822 32748 2856 32768
rect 2822 32700 2856 32710
rect 2822 32676 2856 32700
rect 2822 32632 2856 32638
rect 2822 32604 2856 32632
rect 2822 32564 2856 32566
rect 2822 32532 2856 32564
rect 2822 32462 2856 32494
rect 2822 32460 2856 32462
rect 2822 32394 2856 32422
rect 2822 32388 2856 32394
rect 2822 32326 2856 32350
rect 2822 32316 2856 32326
rect 2822 32258 2856 32278
rect 2822 32244 2856 32258
rect 2822 32190 2856 32206
rect 2822 32172 2856 32190
rect 2822 32122 2856 32134
rect 2822 32100 2856 32122
rect 2822 32054 2856 32062
rect 2822 32028 2856 32054
rect 2822 31986 2856 31990
rect 2822 31956 2856 31986
rect 2822 31884 2856 31918
rect 2822 31816 2856 31846
rect 2822 31812 2856 31816
rect 2822 31748 2856 31774
rect 2822 31740 2856 31748
rect 2822 31680 2856 31702
rect 2822 31668 2856 31680
rect 2822 31612 2856 31630
rect 2822 31596 2856 31612
rect 2822 31544 2856 31558
rect 2822 31524 2856 31544
rect 2822 31476 2856 31486
rect 2822 31452 2856 31476
rect 2822 31408 2856 31414
rect 2822 31380 2856 31408
rect 2822 31340 2856 31342
rect 2822 31308 2856 31340
rect 2822 31238 2856 31270
rect 2822 31236 2856 31238
rect 2822 31170 2856 31198
rect 2822 31164 2856 31170
rect 2822 31102 2856 31126
rect 2822 31092 2856 31102
rect 2822 31034 2856 31054
rect 2822 31020 2856 31034
rect 2822 30966 2856 30982
rect 2822 30948 2856 30966
rect 2822 30898 2856 30910
rect 2822 30876 2856 30898
rect 2822 30830 2856 30838
rect 2822 30804 2856 30830
rect 2822 30762 2856 30766
rect 2822 30732 2856 30762
rect 2822 30660 2856 30694
rect 2822 30592 2856 30622
rect 2822 30588 2856 30592
rect 2822 30524 2856 30550
rect 2822 30516 2856 30524
rect 2822 30456 2856 30478
rect 2822 30444 2856 30456
rect 2822 30388 2856 30406
rect 2822 30372 2856 30388
rect 2822 30320 2856 30334
rect 2822 30300 2856 30320
rect 2822 30252 2856 30262
rect 2822 30228 2856 30252
rect 2822 30184 2856 30190
rect 2822 30156 2856 30184
rect 2822 30116 2856 30118
rect 2822 30084 2856 30116
rect 2822 30014 2856 30046
rect 2822 30012 2856 30014
rect 2822 29946 2856 29974
rect 2822 29940 2856 29946
rect 2822 29878 2856 29902
rect 2822 29868 2856 29878
rect 2822 29810 2856 29830
rect 2822 29796 2856 29810
rect 2822 29742 2856 29758
rect 2822 29724 2856 29742
rect 2822 29674 2856 29686
rect 2822 29652 2856 29674
rect 2822 29606 2856 29614
rect 2822 29580 2856 29606
rect 2822 29538 2856 29542
rect 2822 29508 2856 29538
rect 2822 29436 2856 29470
rect 2822 29368 2856 29398
rect 2822 29364 2856 29368
rect 2822 29300 2856 29326
rect 2822 29292 2856 29300
rect 2822 29232 2856 29254
rect 2822 29220 2856 29232
rect 2822 29164 2856 29182
rect 2822 29148 2856 29164
rect 2822 29096 2856 29110
rect 2822 29076 2856 29096
rect 2822 29028 2856 29038
rect 2822 29004 2856 29028
rect 2822 28960 2856 28966
rect 2822 28932 2856 28960
rect 2822 28892 2856 28894
rect 2822 28860 2856 28892
rect 2822 28790 2856 28822
rect 2822 28788 2856 28790
rect 2822 28722 2856 28750
rect 2822 28716 2856 28722
rect 2822 28654 2856 28678
rect 2822 28644 2856 28654
rect 2822 28586 2856 28606
rect 2822 28572 2856 28586
rect 2822 28518 2856 28534
rect 2822 28500 2856 28518
rect 2822 28450 2856 28462
rect 2822 28428 2856 28450
rect 3157 39580 3188 39614
rect 3188 39580 3191 39614
rect 3232 39580 3256 39614
rect 3256 39580 3266 39614
rect 3307 39580 3324 39614
rect 3324 39580 3341 39614
rect 3382 39580 3392 39614
rect 3392 39580 3416 39614
rect 3457 39580 3460 39614
rect 3460 39580 3491 39614
rect 3532 39580 3562 39614
rect 3562 39580 3566 39614
rect 3607 39580 3630 39614
rect 3630 39580 3641 39614
rect 3682 39580 3698 39614
rect 3698 39580 3716 39614
rect 3757 39580 3766 39614
rect 3766 39580 3791 39614
rect 3832 39580 3834 39614
rect 3834 39580 3866 39614
rect 3907 39580 3936 39614
rect 3936 39580 3941 39614
rect 3982 39580 4004 39614
rect 4004 39580 4016 39614
rect 4057 39580 4072 39614
rect 4072 39580 4091 39614
rect 4132 39580 4140 39614
rect 4140 39580 4166 39614
rect 4207 39580 4208 39614
rect 4208 39580 4241 39614
rect 4282 39580 4310 39614
rect 4310 39580 4316 39614
rect 4357 39580 4378 39614
rect 4378 39580 4391 39614
rect 4433 39580 4446 39614
rect 4446 39580 4467 39614
rect 4509 39580 4514 39614
rect 4514 39580 4543 39614
rect 4619 39580 4650 39614
rect 4650 39580 4653 39614
rect 4698 39580 4718 39614
rect 4718 39580 4732 39614
rect 4778 39580 4786 39614
rect 4786 39580 4812 39614
rect 4858 39580 4888 39614
rect 4888 39580 4892 39614
rect 4938 39580 4956 39614
rect 4956 39580 4972 39614
rect 5018 39580 5024 39614
rect 5024 39580 5052 39614
rect 5098 39580 5126 39614
rect 5126 39580 5132 39614
rect 5178 39580 5194 39614
rect 5194 39580 5212 39614
rect 5258 39580 5262 39614
rect 5262 39580 5292 39614
rect 3082 39512 3116 39542
rect 3082 39508 3116 39512
rect 3082 39444 3116 39469
rect 3082 39435 3116 39444
rect 5330 39508 5364 39542
rect 3082 39376 3116 39396
rect 3082 39362 3116 39376
rect 3082 39308 3116 39323
rect 3082 39289 3116 39308
rect 3082 39240 3116 39250
rect 3082 39216 3116 39240
rect 3082 39172 3116 39177
rect 3082 39143 3116 39172
rect 3082 39070 3116 39104
rect 3082 39002 3116 39031
rect 3082 38997 3116 39002
rect 3082 38934 3116 38958
rect 3082 38924 3116 38934
rect 3082 38866 3116 38885
rect 3082 38851 3116 38866
rect 3082 38798 3116 38812
rect 3082 38778 3116 38798
rect 3082 38730 3116 38739
rect 3082 38705 3116 38730
rect 3082 38662 3116 38666
rect 3082 38632 3116 38662
rect 3082 38560 3116 38593
rect 3082 38559 3116 38560
rect 3082 38492 3116 38520
rect 3082 38486 3116 38492
rect 3082 38424 3116 38447
rect 3082 38413 3116 38424
rect 3082 38356 3116 38374
rect 3082 38340 3116 38356
rect 3082 38288 3116 38301
rect 3082 38267 3116 38288
rect 3082 38220 3116 38228
rect 3082 38194 3116 38220
rect 3082 38152 3116 38155
rect 3082 38121 3116 38152
rect 3082 38050 3116 38082
rect 3082 38048 3116 38050
rect 3082 37982 3116 38010
rect 3082 37976 3116 37982
rect 3082 37914 3116 37938
rect 3082 37904 3116 37914
rect 3082 37846 3116 37866
rect 3082 37832 3116 37846
rect 3082 37778 3116 37794
rect 3082 37760 3116 37778
rect 3082 37710 3116 37722
rect 3082 37688 3116 37710
rect 3082 37642 3116 37650
rect 3082 37616 3116 37642
rect 3082 37574 3116 37578
rect 3082 37544 3116 37574
rect 3082 37472 3116 37506
rect 3082 37404 3116 37434
rect 3082 37400 3116 37404
rect 3082 37336 3116 37362
rect 3082 37328 3116 37336
rect 3082 37268 3116 37290
rect 3082 37256 3116 37268
rect 3082 37200 3116 37218
rect 3082 37184 3116 37200
rect 3082 37132 3116 37146
rect 3082 37112 3116 37132
rect 3082 37064 3116 37074
rect 3082 37040 3116 37064
rect 3082 36996 3116 37002
rect 3082 36968 3116 36996
rect 3082 36928 3116 36930
rect 3082 36896 3116 36928
rect 3082 36826 3116 36858
rect 3082 36824 3116 36826
rect 3082 36758 3116 36786
rect 3082 36752 3116 36758
rect 3082 36690 3116 36714
rect 3082 36680 3116 36690
rect 3082 36622 3116 36642
rect 3082 36608 3116 36622
rect 3082 36554 3116 36570
rect 3082 36536 3116 36554
rect 3082 36486 3116 36498
rect 3082 36464 3116 36486
rect 3082 36418 3116 36426
rect 3082 36392 3116 36418
rect 3082 36350 3116 36354
rect 3082 36320 3116 36350
rect 3082 36248 3116 36282
rect 3082 36180 3116 36210
rect 3082 36176 3116 36180
rect 3082 36112 3116 36138
rect 3082 36104 3116 36112
rect 3082 36044 3116 36066
rect 3082 36032 3116 36044
rect 3082 35976 3116 35994
rect 3082 35960 3116 35976
rect 3082 35908 3116 35922
rect 3082 35888 3116 35908
rect 3082 35840 3116 35850
rect 3082 35816 3116 35840
rect 3082 35772 3116 35778
rect 3082 35744 3116 35772
rect 3082 35704 3116 35706
rect 3082 35672 3116 35704
rect 3082 35602 3116 35634
rect 3082 35600 3116 35602
rect 3082 35534 3116 35562
rect 3082 35528 3116 35534
rect 3082 35466 3116 35490
rect 3082 35456 3116 35466
rect 3082 35398 3116 35418
rect 3082 35384 3116 35398
rect 3082 35330 3116 35346
rect 3082 35312 3116 35330
rect 3082 35262 3116 35274
rect 3082 35240 3116 35262
rect 3082 35194 3116 35202
rect 3082 35168 3116 35194
rect 3082 35126 3116 35130
rect 3082 35096 3116 35126
rect 3082 35024 3116 35058
rect 3082 34956 3116 34986
rect 3082 34952 3116 34956
rect 3082 34888 3116 34914
rect 3082 34880 3116 34888
rect 3082 34820 3116 34842
rect 3082 34808 3116 34820
rect 3082 34752 3116 34770
rect 3082 34736 3116 34752
rect 3082 34684 3116 34698
rect 3082 34664 3116 34684
rect 3082 34616 3116 34626
rect 3082 34592 3116 34616
rect 3082 34548 3116 34554
rect 3082 34520 3116 34548
rect 3082 34480 3116 34482
rect 3082 34448 3116 34480
rect 3082 34378 3116 34410
rect 3082 34376 3116 34378
rect 3082 34310 3116 34338
rect 3082 34304 3116 34310
rect 3082 34242 3116 34266
rect 3082 34232 3116 34242
rect 3082 34174 3116 34194
rect 3082 34160 3116 34174
rect 3082 34106 3116 34122
rect 3082 34088 3116 34106
rect 3082 34038 3116 34050
rect 3082 34016 3116 34038
rect 3082 33970 3116 33978
rect 3082 33944 3116 33970
rect 3082 33902 3116 33906
rect 3082 33872 3116 33902
rect 3082 33800 3116 33834
rect 3082 33732 3116 33762
rect 3082 33728 3116 33732
rect 3082 33664 3116 33690
rect 3082 33656 3116 33664
rect 3082 33596 3116 33618
rect 3082 33584 3116 33596
rect 3082 33528 3116 33546
rect 3082 33512 3116 33528
rect 3082 33460 3116 33474
rect 3082 33440 3116 33460
rect 3082 33392 3116 33402
rect 3082 33368 3116 33392
rect 3082 33324 3116 33330
rect 3082 33296 3116 33324
rect 3082 33256 3116 33258
rect 3082 33224 3116 33256
rect 3082 33154 3116 33186
rect 3082 33152 3116 33154
rect 3082 33086 3116 33114
rect 3082 33080 3116 33086
rect 3082 33018 3116 33042
rect 3082 33008 3116 33018
rect 3082 32950 3116 32970
rect 3082 32936 3116 32950
rect 3082 32882 3116 32898
rect 3082 32864 3116 32882
rect 3082 32814 3116 32826
rect 3082 32792 3116 32814
rect 3082 32746 3116 32754
rect 3082 32720 3116 32746
rect 3082 32678 3116 32682
rect 3082 32648 3116 32678
rect 3082 32576 3116 32610
rect 3082 32508 3116 32538
rect 3082 32504 3116 32508
rect 3082 32440 3116 32466
rect 3082 32432 3116 32440
rect 3082 32372 3116 32394
rect 3082 32360 3116 32372
rect 3082 32304 3116 32322
rect 3082 32288 3116 32304
rect 3082 32236 3116 32250
rect 3082 32216 3116 32236
rect 3082 32168 3116 32178
rect 3082 32144 3116 32168
rect 3082 32100 3116 32106
rect 3082 32072 3116 32100
rect 3082 32032 3116 32034
rect 3082 32000 3116 32032
rect 3082 31930 3116 31962
rect 3082 31928 3116 31930
rect 3082 31862 3116 31890
rect 3082 31856 3116 31862
rect 3082 31794 3116 31818
rect 3082 31784 3116 31794
rect 3082 31726 3116 31746
rect 3082 31712 3116 31726
rect 3082 31658 3116 31674
rect 3082 31640 3116 31658
rect 3082 31590 3116 31602
rect 3082 31568 3116 31590
rect 3082 31522 3116 31530
rect 3082 31496 3116 31522
rect 3082 31454 3116 31458
rect 3082 31424 3116 31454
rect 3082 31352 3116 31386
rect 3082 31284 3116 31314
rect 3082 31280 3116 31284
rect 3082 31216 3116 31242
rect 3082 31208 3116 31216
rect 3082 31148 3116 31170
rect 3082 31136 3116 31148
rect 3082 31080 3116 31098
rect 3082 31064 3116 31080
rect 3082 31012 3116 31026
rect 3082 30992 3116 31012
rect 3082 30944 3116 30954
rect 3082 30920 3116 30944
rect 3082 30876 3116 30882
rect 3082 30848 3116 30876
rect 3082 30808 3116 30810
rect 3082 30776 3116 30808
rect 3082 30706 3116 30738
rect 3082 30704 3116 30706
rect 3082 30638 3116 30666
rect 3082 30632 3116 30638
rect 3082 30570 3116 30594
rect 3082 30560 3116 30570
rect 3082 30502 3116 30522
rect 3082 30488 3116 30502
rect 3082 30434 3116 30450
rect 3082 30416 3116 30434
rect 3174 39329 3208 39353
rect 3174 39319 3208 39329
rect 3174 39261 3208 39281
rect 3174 39247 3208 39261
rect 3174 39193 3208 39209
rect 3174 39175 3208 39193
rect 3174 39125 3208 39137
rect 3174 39103 3208 39125
rect 3174 39057 3208 39065
rect 3174 39031 3208 39057
rect 3174 38989 3208 38993
rect 3174 38959 3208 38989
rect 3174 38887 3208 38921
rect 3174 38819 3208 38849
rect 3174 38815 3208 38819
rect 3174 38751 3208 38777
rect 3174 38743 3208 38751
rect 3174 38683 3208 38705
rect 3174 38671 3208 38683
rect 3174 38615 3208 38633
rect 3174 38599 3208 38615
rect 3174 38547 3208 38561
rect 3174 38527 3208 38547
rect 3174 38479 3208 38489
rect 3174 38455 3208 38479
rect 3174 38411 3208 38417
rect 3174 38383 3208 38411
rect 3174 38343 3208 38345
rect 3174 38311 3208 38343
rect 3174 38241 3208 38273
rect 3174 38239 3208 38241
rect 3174 38173 3208 38201
rect 3174 38167 3208 38173
rect 3174 38105 3208 38129
rect 3174 38095 3208 38105
rect 3174 38037 3208 38057
rect 3174 38023 3208 38037
rect 3174 37969 3208 37985
rect 3174 37951 3208 37969
rect 3174 37901 3208 37913
rect 3174 37879 3208 37901
rect 3174 37833 3208 37841
rect 3174 37807 3208 37833
rect 3174 37765 3208 37769
rect 3174 37735 3208 37765
rect 3174 37663 3208 37697
rect 3174 37595 3208 37625
rect 3174 37591 3208 37595
rect 3174 37527 3208 37553
rect 3174 37519 3208 37527
rect 3174 37459 3208 37481
rect 3174 37447 3208 37459
rect 3174 37391 3208 37409
rect 3174 37375 3208 37391
rect 3174 37323 3208 37337
rect 3174 37303 3208 37323
rect 3174 37255 3208 37265
rect 3174 37231 3208 37255
rect 3174 37187 3208 37193
rect 3174 37159 3208 37187
rect 3174 37119 3208 37121
rect 3174 37087 3208 37119
rect 3174 37017 3208 37049
rect 3174 37015 3208 37017
rect 3174 36949 3208 36977
rect 3174 36943 3208 36949
rect 3174 36881 3208 36905
rect 3174 36871 3208 36881
rect 3174 36813 3208 36833
rect 3174 36799 3208 36813
rect 3174 36745 3208 36761
rect 3174 36727 3208 36745
rect 3174 36677 3208 36689
rect 3174 36655 3208 36677
rect 3174 36609 3208 36617
rect 3174 36583 3208 36609
rect 3174 36541 3208 36545
rect 3174 36511 3208 36541
rect 3174 36439 3208 36473
rect 3174 36371 3208 36401
rect 3174 36367 3208 36371
rect 3174 36303 3208 36329
rect 3174 36295 3208 36303
rect 3174 36235 3208 36257
rect 3174 36223 3208 36235
rect 3174 36167 3208 36185
rect 3174 36151 3208 36167
rect 3174 36099 3208 36113
rect 3174 36079 3208 36099
rect 3174 36031 3208 36041
rect 3174 36007 3208 36031
rect 3174 35963 3208 35969
rect 3174 35935 3208 35963
rect 3174 35895 3208 35897
rect 3174 35863 3208 35895
rect 3174 35793 3208 35825
rect 3174 35791 3208 35793
rect 3174 35725 3208 35753
rect 3174 35719 3208 35725
rect 3174 35657 3208 35681
rect 3174 35647 3208 35657
rect 3174 35589 3208 35609
rect 3174 35575 3208 35589
rect 3174 35521 3208 35537
rect 3174 35503 3208 35521
rect 3174 35453 3208 35465
rect 3174 35431 3208 35453
rect 3174 35385 3208 35393
rect 3174 35359 3208 35385
rect 3174 35317 3208 35321
rect 3174 35287 3208 35317
rect 3174 35215 3208 35249
rect 3174 35147 3208 35177
rect 3174 35143 3208 35147
rect 3174 35079 3208 35105
rect 3174 35071 3208 35079
rect 3174 35011 3208 35033
rect 3174 34999 3208 35011
rect 3174 34943 3208 34961
rect 3174 34927 3208 34943
rect 3174 34875 3208 34889
rect 3174 34855 3208 34875
rect 3174 34807 3208 34817
rect 3174 34783 3208 34807
rect 3174 34739 3208 34745
rect 3174 34711 3208 34739
rect 3174 34671 3208 34673
rect 3174 34639 3208 34671
rect 3174 34569 3208 34601
rect 3174 34567 3208 34569
rect 3174 34501 3208 34529
rect 3174 34495 3208 34501
rect 3174 34433 3208 34457
rect 3174 34423 3208 34433
rect 3174 34365 3208 34385
rect 3174 34351 3208 34365
rect 3174 34297 3208 34313
rect 3174 34279 3208 34297
rect 3174 34229 3208 34241
rect 3174 34207 3208 34229
rect 3174 34161 3208 34169
rect 3174 34135 3208 34161
rect 3174 34093 3208 34097
rect 3174 34063 3208 34093
rect 3174 33991 3208 34025
rect 3174 33923 3208 33953
rect 3174 33919 3208 33923
rect 3174 33855 3208 33881
rect 3174 33847 3208 33855
rect 3174 33787 3208 33809
rect 3174 33775 3208 33787
rect 3174 33719 3208 33737
rect 3174 33703 3208 33719
rect 3174 33651 3208 33665
rect 3174 33631 3208 33651
rect 3174 33583 3208 33593
rect 3174 33559 3208 33583
rect 3174 33515 3208 33521
rect 3174 33487 3208 33515
rect 3174 33447 3208 33449
rect 3174 33415 3208 33447
rect 3174 33345 3208 33377
rect 3174 33343 3208 33345
rect 3174 33277 3208 33305
rect 3174 33271 3208 33277
rect 3174 33209 3208 33233
rect 3174 33199 3208 33209
rect 3174 33141 3208 33161
rect 3174 33127 3208 33141
rect 3174 33073 3208 33089
rect 3174 33055 3208 33073
rect 3174 33005 3208 33017
rect 3174 32983 3208 33005
rect 3174 32937 3208 32945
rect 3174 32911 3208 32937
rect 3174 32869 3208 32873
rect 3174 32839 3208 32869
rect 3174 32767 3208 32801
rect 3174 32699 3208 32729
rect 3174 32695 3208 32699
rect 3174 32631 3208 32657
rect 3174 32623 3208 32631
rect 3174 32563 3208 32585
rect 3174 32551 3208 32563
rect 3174 32495 3208 32513
rect 3174 32479 3208 32495
rect 3174 32427 3208 32441
rect 3174 32407 3208 32427
rect 3174 32359 3208 32369
rect 3174 32335 3208 32359
rect 3174 32291 3208 32296
rect 3174 32262 3208 32291
rect 3174 32189 3208 32223
rect 3174 32121 3208 32150
rect 3174 32116 3208 32121
rect 3174 32053 3208 32077
rect 3174 32043 3208 32053
rect 3174 31985 3208 32004
rect 3174 31970 3208 31985
rect 3174 31917 3208 31931
rect 3174 31897 3208 31917
rect 3174 31848 3208 31858
rect 3174 31824 3208 31848
rect 3174 31779 3208 31785
rect 3174 31751 3208 31779
rect 3174 31710 3208 31712
rect 3174 31678 3208 31710
rect 3174 31606 3208 31639
rect 3174 31605 3208 31606
rect 3174 31537 3208 31566
rect 3174 31532 3208 31537
rect 3174 31468 3208 31493
rect 3174 31459 3208 31468
rect 3174 31399 3208 31420
rect 3174 31386 3208 31399
rect 3174 31330 3208 31347
rect 3174 31313 3208 31330
rect 3174 31261 3208 31274
rect 3174 31240 3208 31261
rect 3174 31192 3208 31201
rect 3174 31167 3208 31192
rect 3174 31123 3208 31128
rect 3174 31094 3208 31123
rect 3174 31054 3208 31055
rect 3174 31021 3208 31054
rect 3174 30951 3208 30982
rect 3174 30948 3208 30951
rect 3174 30882 3208 30909
rect 3174 30875 3208 30882
rect 3174 30813 3208 30836
rect 3174 30802 3208 30813
rect 3174 30744 3208 30763
rect 3174 30729 3208 30744
rect 3174 30675 3208 30690
rect 3174 30656 3208 30675
rect 3174 30606 3208 30617
rect 3174 30583 3208 30606
rect 3174 30537 3208 30544
rect 3174 30510 3208 30537
rect 3174 30468 3208 30471
rect 3174 30437 3208 30468
rect 5330 39440 5364 39470
rect 5330 39436 5364 39440
rect 5330 39372 5364 39398
rect 5330 39364 5364 39372
rect 5330 39304 5364 39326
rect 5330 39292 5364 39304
rect 5330 39236 5364 39254
rect 5330 39220 5364 39236
rect 5330 39168 5364 39182
rect 5330 39148 5364 39168
rect 5330 39100 5364 39110
rect 5330 39076 5364 39100
rect 5330 39032 5364 39038
rect 5330 39004 5364 39032
rect 5330 38964 5364 38966
rect 5330 38932 5364 38964
rect 5330 38862 5364 38894
rect 5330 38860 5364 38862
rect 5330 38794 5364 38822
rect 5330 38788 5364 38794
rect 5330 38726 5364 38750
rect 5330 38716 5364 38726
rect 5330 38658 5364 38678
rect 5330 38644 5364 38658
rect 5330 38590 5364 38606
rect 5330 38572 5364 38590
rect 5330 38522 5364 38534
rect 5330 38500 5364 38522
rect 5330 38454 5364 38462
rect 5330 38428 5364 38454
rect 5330 38386 5364 38390
rect 5330 38356 5364 38386
rect 5330 38284 5364 38318
rect 5330 38216 5364 38246
rect 5330 38212 5364 38216
rect 5330 38148 5364 38174
rect 5330 38140 5364 38148
rect 5330 38080 5364 38102
rect 5330 38068 5364 38080
rect 5330 38012 5364 38030
rect 5330 37996 5364 38012
rect 5330 37944 5364 37958
rect 5330 37924 5364 37944
rect 5330 37876 5364 37886
rect 5330 37852 5364 37876
rect 5330 37808 5364 37814
rect 5330 37780 5364 37808
rect 5330 37740 5364 37742
rect 5330 37708 5364 37740
rect 5330 37638 5364 37670
rect 5330 37636 5364 37638
rect 5330 37570 5364 37598
rect 5330 37564 5364 37570
rect 5330 37502 5364 37526
rect 5330 37492 5364 37502
rect 5330 37434 5364 37454
rect 5330 37420 5364 37434
rect 5330 37366 5364 37382
rect 5330 37348 5364 37366
rect 5330 37298 5364 37310
rect 5330 37276 5364 37298
rect 5330 37230 5364 37238
rect 5330 37204 5364 37230
rect 5330 37162 5364 37166
rect 5330 37132 5364 37162
rect 5330 37060 5364 37094
rect 5330 36992 5364 37022
rect 5330 36988 5364 36992
rect 5330 36924 5364 36950
rect 5330 36916 5364 36924
rect 5330 36856 5364 36878
rect 5330 36844 5364 36856
rect 5330 36788 5364 36806
rect 5330 36772 5364 36788
rect 5330 36720 5364 36734
rect 5330 36700 5364 36720
rect 5330 36652 5364 36662
rect 5330 36628 5364 36652
rect 5330 36584 5364 36590
rect 5330 36556 5364 36584
rect 5330 36516 5364 36518
rect 5330 36484 5364 36516
rect 5330 36414 5364 36446
rect 5330 36412 5364 36414
rect 5330 36346 5364 36374
rect 5330 36340 5364 36346
rect 5330 36278 5364 36302
rect 5330 36268 5364 36278
rect 5330 36210 5364 36230
rect 5330 36196 5364 36210
rect 5330 36142 5364 36158
rect 5330 36124 5364 36142
rect 5330 36074 5364 36086
rect 5330 36052 5364 36074
rect 5330 36006 5364 36014
rect 5330 35980 5364 36006
rect 5330 35938 5364 35942
rect 5330 35908 5364 35938
rect 5330 35836 5364 35870
rect 5330 35768 5364 35798
rect 5330 35764 5364 35768
rect 5330 35700 5364 35726
rect 5330 35692 5364 35700
rect 5330 35632 5364 35654
rect 5330 35620 5364 35632
rect 5330 35564 5364 35582
rect 5330 35548 5364 35564
rect 5330 35496 5364 35510
rect 5330 35476 5364 35496
rect 5330 35428 5364 35438
rect 5330 35404 5364 35428
rect 5330 35360 5364 35366
rect 5330 35332 5364 35360
rect 5330 35292 5364 35294
rect 5330 35260 5364 35292
rect 5330 35190 5364 35222
rect 5330 35188 5364 35190
rect 5330 35122 5364 35149
rect 5330 35115 5364 35122
rect 5330 35054 5364 35076
rect 5330 35042 5364 35054
rect 5330 34986 5364 35003
rect 5330 34969 5364 34986
rect 5330 34918 5364 34930
rect 5330 34896 5364 34918
rect 5330 34850 5364 34857
rect 5330 34823 5364 34850
rect 5330 34782 5364 34784
rect 5330 34750 5364 34782
rect 5330 34680 5364 34711
rect 5330 34677 5364 34680
rect 5330 34612 5364 34638
rect 5330 34604 5364 34612
rect 5330 34544 5364 34565
rect 5330 34531 5364 34544
rect 5330 34476 5364 34492
rect 5330 34458 5364 34476
rect 5330 34408 5364 34419
rect 5330 34385 5364 34408
rect 5330 34340 5364 34346
rect 5330 34312 5364 34340
rect 5330 34272 5364 34273
rect 5330 34239 5364 34272
rect 5330 34170 5364 34200
rect 5330 34166 5364 34170
rect 5330 34102 5364 34127
rect 5330 34093 5364 34102
rect 5330 34034 5364 34054
rect 5330 34020 5364 34034
rect 5330 33966 5364 33981
rect 5330 33947 5364 33966
rect 5330 33898 5364 33908
rect 5330 33874 5364 33898
rect 5330 33830 5364 33835
rect 5330 33801 5364 33830
rect 5330 33728 5364 33762
rect 5330 33660 5364 33689
rect 5330 33655 5364 33660
rect 5330 33592 5364 33616
rect 5330 33582 5364 33592
rect 5330 33524 5364 33543
rect 5330 33509 5364 33524
rect 5330 33456 5364 33470
rect 5330 33436 5364 33456
rect 5330 33388 5364 33397
rect 5330 33363 5364 33388
rect 5330 33320 5364 33324
rect 5330 33290 5364 33320
rect 5330 33218 5364 33251
rect 5330 33217 5364 33218
rect 5330 33150 5364 33178
rect 5330 33144 5364 33150
rect 5330 33082 5364 33105
rect 5330 33071 5364 33082
rect 5330 33014 5364 33032
rect 5330 32998 5364 33014
rect 5330 32946 5364 32959
rect 5330 32925 5364 32946
rect 5330 32878 5364 32886
rect 5330 32852 5364 32878
rect 5330 32810 5364 32813
rect 5330 32779 5364 32810
rect 5330 32708 5364 32740
rect 5330 32706 5364 32708
rect 5330 32640 5364 32667
rect 5330 32633 5364 32640
rect 5330 32572 5364 32594
rect 5330 32560 5364 32572
rect 5330 32504 5364 32521
rect 5330 32487 5364 32504
rect 5330 32436 5364 32448
rect 5330 32414 5364 32436
rect 5330 32368 5364 32375
rect 5330 32341 5364 32368
rect 5330 32300 5364 32302
rect 5330 32268 5364 32300
rect 5330 32198 5364 32229
rect 5330 32195 5364 32198
rect 5330 32130 5364 32156
rect 5330 32122 5364 32130
rect 5330 32062 5364 32083
rect 5330 32049 5364 32062
rect 5330 31994 5364 32010
rect 5330 31976 5364 31994
rect 5330 31926 5364 31937
rect 5330 31903 5364 31926
rect 5330 31858 5364 31864
rect 5330 31830 5364 31858
rect 5330 31790 5364 31791
rect 5330 31757 5364 31790
rect 5330 31688 5364 31718
rect 5330 31684 5364 31688
rect 5330 31620 5364 31645
rect 5330 31611 5364 31620
rect 5330 31552 5364 31572
rect 5330 31538 5364 31552
rect 5330 31484 5364 31499
rect 5330 31465 5364 31484
rect 5330 31416 5364 31426
rect 5330 31392 5364 31416
rect 5330 31348 5364 31353
rect 5330 31319 5364 31348
rect 5330 31246 5364 31280
rect 5330 31178 5364 31207
rect 5330 31173 5364 31178
rect 5330 31110 5364 31134
rect 5330 31100 5364 31110
rect 5330 31042 5364 31061
rect 5330 31027 5364 31042
rect 5330 30974 5364 30988
rect 5330 30954 5364 30974
rect 5330 30906 5364 30915
rect 5330 30881 5364 30906
rect 5330 30838 5364 30842
rect 5330 30808 5364 30838
rect 5330 30736 5364 30769
rect 5330 30735 5364 30736
rect 5330 30668 5364 30696
rect 5330 30662 5364 30668
rect 5330 30600 5364 30623
rect 5330 30589 5364 30600
rect 5330 30532 5364 30550
rect 5330 30516 5364 30532
rect 5330 30464 5364 30477
rect 5330 30443 5364 30464
rect 3082 30366 3116 30378
rect 3082 30344 3116 30366
rect 5330 30396 5364 30404
rect 5330 30370 5364 30396
rect 7746 39564 7780 39586
rect 7746 39552 7780 39564
rect 7746 39496 7780 39514
rect 7746 39480 7780 39496
rect 7746 39428 7780 39442
rect 7746 39408 7780 39428
rect 7746 39360 7780 39370
rect 7746 39336 7780 39360
rect 7746 39292 7780 39298
rect 7746 39264 7780 39292
rect 7746 39224 7780 39226
rect 7746 39192 7780 39224
rect 7746 39122 7780 39154
rect 7746 39120 7780 39122
rect 7746 39054 7780 39082
rect 7746 39048 7780 39054
rect 7746 38986 7780 39010
rect 7746 38976 7780 38986
rect 7746 38918 7780 38938
rect 7746 38904 7780 38918
rect 7746 38850 7780 38866
rect 7746 38832 7780 38850
rect 7746 38782 7780 38794
rect 7746 38760 7780 38782
rect 7746 38714 7780 38722
rect 7746 38688 7780 38714
rect 7746 38646 7780 38650
rect 7746 38616 7780 38646
rect 7746 38544 7780 38578
rect 7746 38476 7780 38506
rect 7746 38472 7780 38476
rect 7746 38408 7780 38434
rect 7746 38400 7780 38408
rect 7746 38340 7780 38362
rect 7746 38328 7780 38340
rect 7746 38272 7780 38290
rect 7746 38256 7780 38272
rect 7746 38204 7780 38218
rect 7746 38184 7780 38204
rect 7746 38136 7780 38146
rect 7746 38112 7780 38136
rect 7746 38068 7780 38074
rect 7746 38040 7780 38068
rect 7746 38000 7780 38002
rect 7746 37968 7780 38000
rect 7746 37898 7780 37930
rect 7746 37896 7780 37898
rect 7746 37830 7780 37858
rect 7746 37824 7780 37830
rect 7746 37762 7780 37786
rect 7746 37752 7780 37762
rect 7746 37694 7780 37714
rect 7746 37680 7780 37694
rect 7746 37626 7780 37642
rect 7746 37608 7780 37626
rect 7746 37558 7780 37570
rect 7746 37536 7780 37558
rect 7746 37490 7780 37498
rect 7746 37464 7780 37490
rect 7746 37422 7780 37426
rect 7746 37392 7780 37422
rect 7746 37320 7780 37354
rect 7746 37252 7780 37282
rect 7746 37248 7780 37252
rect 7746 37184 7780 37210
rect 7746 37176 7780 37184
rect 7746 37116 7780 37138
rect 7746 37104 7780 37116
rect 7746 37048 7780 37066
rect 7746 37032 7780 37048
rect 7746 36980 7780 36994
rect 7746 36960 7780 36980
rect 7746 36912 7780 36922
rect 7746 36888 7780 36912
rect 7746 36844 7780 36850
rect 7746 36816 7780 36844
rect 7746 36776 7780 36778
rect 7746 36744 7780 36776
rect 7746 36674 7780 36706
rect 7746 36672 7780 36674
rect 7746 36606 7780 36634
rect 7746 36600 7780 36606
rect 7746 36538 7780 36562
rect 7746 36528 7780 36538
rect 7746 36470 7780 36490
rect 7746 36456 7780 36470
rect 7746 36402 7780 36418
rect 7746 36384 7780 36402
rect 7746 36334 7780 36346
rect 7746 36312 7780 36334
rect 7746 36266 7780 36274
rect 7746 36240 7780 36266
rect 7746 36198 7780 36202
rect 7746 36168 7780 36198
rect 7746 36096 7780 36130
rect 7746 36028 7780 36058
rect 7746 36024 7780 36028
rect 7746 35960 7780 35986
rect 7746 35952 7780 35960
rect 7746 35892 7780 35914
rect 7746 35880 7780 35892
rect 7746 35824 7780 35842
rect 7746 35808 7780 35824
rect 7746 35756 7780 35770
rect 7746 35736 7780 35756
rect 7746 35688 7780 35698
rect 7746 35664 7780 35688
rect 7746 35620 7780 35626
rect 7746 35592 7780 35620
rect 7746 35552 7780 35554
rect 7746 35520 7780 35552
rect 7746 35450 7780 35482
rect 7746 35448 7780 35450
rect 7746 35382 7780 35410
rect 7746 35376 7780 35382
rect 7746 35314 7780 35338
rect 7746 35304 7780 35314
rect 7746 35246 7780 35266
rect 7746 35232 7780 35246
rect 7746 35178 7780 35194
rect 7746 35160 7780 35178
rect 7746 35110 7780 35122
rect 7746 35088 7780 35110
rect 7746 35042 7780 35050
rect 7746 35016 7780 35042
rect 7746 34974 7780 34978
rect 7746 34944 7780 34974
rect 7746 34872 7780 34906
rect 7746 34804 7780 34834
rect 7746 34800 7780 34804
rect 7746 34736 7780 34762
rect 7746 34728 7780 34736
rect 7746 34668 7780 34690
rect 7746 34656 7780 34668
rect 7746 34600 7780 34618
rect 7746 34584 7780 34600
rect 7746 34532 7780 34546
rect 7746 34512 7780 34532
rect 7746 34464 7780 34474
rect 7746 34440 7780 34464
rect 7746 34396 7780 34402
rect 7746 34368 7780 34396
rect 7746 34328 7780 34330
rect 7746 34296 7780 34328
rect 7746 34226 7780 34258
rect 7746 34224 7780 34226
rect 7746 34158 7780 34186
rect 7746 34152 7780 34158
rect 7746 34090 7780 34114
rect 7746 34080 7780 34090
rect 7746 34022 7780 34042
rect 7746 34008 7780 34022
rect 7746 33954 7780 33970
rect 7746 33936 7780 33954
rect 7746 33886 7780 33898
rect 7746 33864 7780 33886
rect 7746 33818 7780 33826
rect 7746 33792 7780 33818
rect 7746 33750 7780 33754
rect 7746 33720 7780 33750
rect 7746 33648 7780 33682
rect 7746 33580 7780 33610
rect 7746 33576 7780 33580
rect 7746 33512 7780 33538
rect 7746 33504 7780 33512
rect 7746 33444 7780 33466
rect 7746 33432 7780 33444
rect 7746 33376 7780 33394
rect 7746 33360 7780 33376
rect 7746 33308 7780 33322
rect 7746 33288 7780 33308
rect 7746 33240 7780 33250
rect 7746 33216 7780 33240
rect 7746 33172 7780 33178
rect 7746 33144 7780 33172
rect 7746 33104 7780 33106
rect 7746 33072 7780 33104
rect 7746 33002 7780 33034
rect 7746 33000 7780 33002
rect 7746 32934 7780 32962
rect 7746 32928 7780 32934
rect 7746 32866 7780 32890
rect 7746 32856 7780 32866
rect 7746 32798 7780 32818
rect 7746 32784 7780 32798
rect 7746 32730 7780 32746
rect 7746 32712 7780 32730
rect 7746 32662 7780 32674
rect 7746 32640 7780 32662
rect 7746 32594 7780 32602
rect 7746 32568 7780 32594
rect 7746 32526 7780 32530
rect 7746 32496 7780 32526
rect 7746 32424 7780 32458
rect 7746 32356 7780 32386
rect 7746 32352 7780 32356
rect 7746 32288 7780 32314
rect 7746 32280 7780 32288
rect 7746 32220 7780 32242
rect 7746 32208 7780 32220
rect 7746 32152 7780 32170
rect 7746 32136 7780 32152
rect 7746 32084 7780 32098
rect 7746 32064 7780 32084
rect 7746 32016 7780 32026
rect 7746 31992 7780 32016
rect 7746 31948 7780 31954
rect 7746 31920 7780 31948
rect 7746 31880 7780 31882
rect 7746 31848 7780 31880
rect 7746 31778 7780 31810
rect 7746 31776 7780 31778
rect 7746 31710 7780 31738
rect 7746 31704 7780 31710
rect 7746 31642 7780 31666
rect 7746 31632 7780 31642
rect 7746 31574 7780 31594
rect 7746 31560 7780 31574
rect 7746 31506 7780 31522
rect 7746 31488 7780 31506
rect 7746 31438 7780 31450
rect 7746 31416 7780 31438
rect 7746 31370 7780 31378
rect 7746 31344 7780 31370
rect 7746 31302 7780 31306
rect 7746 31272 7780 31302
rect 7746 31200 7780 31234
rect 7746 31132 7780 31162
rect 7746 31128 7780 31132
rect 7746 31064 7780 31090
rect 7746 31056 7780 31064
rect 7746 30996 7780 31018
rect 7746 30984 7780 30996
rect 7746 30928 7780 30946
rect 7746 30912 7780 30928
rect 7746 30860 7780 30874
rect 7746 30840 7780 30860
rect 7746 30792 7780 30801
rect 7746 30767 7780 30792
rect 7746 30724 7780 30728
rect 7746 30694 7780 30724
rect 7746 30622 7780 30655
rect 7746 30621 7780 30622
rect 7746 30554 7780 30582
rect 7746 30548 7780 30554
rect 7746 30486 7780 30509
rect 7746 30475 7780 30486
rect 7746 30418 7780 30436
rect 7746 30402 7780 30418
rect 3082 30298 3116 30306
rect 3082 30272 3116 30298
rect 3082 30230 3116 30234
rect 3082 30200 3116 30230
rect 7746 30350 7780 30363
rect 7746 30329 7780 30350
rect 7746 30282 7780 30290
rect 7746 30256 7780 30282
rect 5646 30163 5664 30197
rect 5664 30163 5680 30197
rect 5721 30163 5735 30197
rect 5735 30163 5755 30197
rect 5796 30163 5806 30197
rect 5806 30163 5830 30197
rect 5871 30163 5877 30197
rect 5877 30163 5905 30197
rect 5946 30163 5948 30197
rect 5948 30163 5980 30197
rect 6021 30163 6053 30197
rect 6053 30163 6055 30197
rect 6096 30163 6124 30197
rect 6124 30163 6130 30197
rect 6171 30163 6195 30197
rect 6195 30163 6205 30197
rect 6246 30163 6266 30197
rect 6266 30163 6280 30197
rect 6321 30163 6337 30197
rect 6337 30163 6355 30197
rect 6396 30163 6408 30197
rect 6408 30163 6430 30197
rect 6471 30163 6478 30197
rect 6478 30163 6505 30197
rect 6546 30163 6548 30197
rect 6548 30163 6580 30197
rect 6621 30163 6654 30197
rect 6654 30163 6655 30197
rect 6696 30163 6724 30197
rect 6724 30163 6730 30197
rect 6770 30163 6794 30197
rect 6794 30163 6804 30197
rect 6844 30163 6864 30197
rect 6864 30163 6878 30197
rect 6918 30163 6934 30197
rect 6934 30163 6952 30197
rect 6992 30163 7004 30197
rect 7004 30163 7026 30197
rect 7066 30163 7074 30197
rect 7074 30163 7100 30197
rect 7140 30163 7144 30197
rect 7144 30163 7174 30197
rect 7214 30163 7248 30197
rect 7288 30163 7318 30197
rect 7318 30163 7322 30197
rect 7362 30163 7388 30197
rect 7388 30163 7396 30197
rect 7436 30163 7458 30197
rect 7458 30163 7470 30197
rect 7746 30214 7780 30217
rect 7746 30183 7780 30214
rect 3082 30128 3116 30162
rect 3689 30123 3723 30125
rect 3764 30123 3798 30125
rect 3839 30123 3873 30125
rect 3914 30123 3948 30125
rect 3989 30123 4023 30125
rect 4064 30123 4098 30125
rect 4139 30123 4173 30125
rect 4214 30123 4248 30125
rect 4289 30123 4323 30125
rect 4364 30123 4398 30125
rect 4439 30123 4473 30125
rect 4514 30123 4548 30125
rect 4589 30123 4623 30125
rect 4664 30123 4698 30125
rect 4739 30123 4773 30125
rect 4814 30123 4848 30125
rect 4889 30123 4923 30125
rect 4964 30123 4998 30125
rect 3082 30060 3116 30090
rect 3082 30056 3116 30060
rect 3689 30091 3690 30123
rect 3690 30091 3723 30123
rect 3764 30091 3794 30123
rect 3794 30091 3798 30123
rect 3839 30091 3864 30123
rect 3864 30091 3873 30123
rect 3914 30091 3933 30123
rect 3933 30091 3948 30123
rect 3989 30091 4002 30123
rect 4002 30091 4023 30123
rect 4064 30091 4071 30123
rect 4071 30091 4098 30123
rect 4139 30091 4140 30123
rect 4140 30091 4173 30123
rect 4214 30091 4244 30123
rect 4244 30091 4248 30123
rect 4289 30091 4313 30123
rect 4313 30091 4323 30123
rect 4364 30091 4382 30123
rect 4382 30091 4398 30123
rect 4439 30091 4451 30123
rect 4451 30091 4473 30123
rect 4514 30091 4520 30123
rect 4520 30091 4548 30123
rect 4589 30091 4623 30123
rect 4664 30091 4692 30123
rect 4692 30091 4698 30123
rect 4739 30091 4761 30123
rect 4761 30091 4773 30123
rect 4814 30091 4830 30123
rect 4830 30091 4848 30123
rect 4889 30091 4899 30123
rect 4899 30091 4923 30123
rect 4964 30091 4968 30123
rect 4968 30091 4998 30123
rect 5038 30091 5072 30125
rect 5112 30123 5146 30125
rect 5186 30123 5220 30125
rect 5112 30091 5141 30123
rect 5141 30091 5146 30123
rect 5186 30091 5210 30123
rect 5210 30091 5220 30123
rect 7746 30112 7780 30144
rect 7746 30110 7780 30112
rect 3082 29992 3116 30018
rect 3082 29984 3116 29992
rect 3082 29924 3116 29946
rect 3082 29912 3116 29924
rect 3082 29856 3116 29874
rect 3082 29840 3116 29856
rect 3082 29788 3116 29802
rect 3082 29768 3116 29788
rect 3082 29720 3116 29730
rect 3082 29696 3116 29720
rect 3082 29652 3116 29658
rect 3082 29624 3116 29652
rect 3082 29584 3116 29586
rect 3082 29552 3116 29584
rect 3082 29482 3116 29514
rect 3082 29480 3116 29482
rect 3082 29414 3116 29442
rect 3082 29408 3116 29414
rect 3082 29346 3116 29370
rect 3082 29336 3116 29346
rect 3082 29278 3116 29298
rect 3082 29264 3116 29278
rect 5640 29998 5674 30002
rect 5640 29968 5674 29998
rect 5640 29896 5674 29928
rect 5640 29894 5674 29896
rect 7746 30044 7780 30071
rect 7746 30037 7780 30044
rect 7746 29976 7780 29998
rect 7746 29964 7780 29976
rect 7746 29908 7780 29925
rect 7746 29891 7780 29908
rect 5640 29828 5674 29854
rect 5640 29820 5674 29828
rect 6214 29854 6237 29888
rect 6237 29854 6248 29888
rect 6286 29854 6305 29888
rect 6305 29854 6320 29888
rect 6446 29854 6461 29888
rect 6461 29854 6480 29888
rect 6518 29854 6529 29888
rect 6529 29854 6552 29888
rect 5640 29760 5674 29780
rect 5640 29746 5674 29760
rect 5640 29692 5674 29706
rect 5640 29672 5674 29692
rect 5640 29624 5674 29631
rect 5640 29597 5674 29624
rect 5640 29522 5674 29556
rect 5640 29454 5674 29481
rect 5640 29447 5674 29454
rect 5640 29386 5674 29406
rect 5640 29372 5674 29386
rect 5640 29318 5674 29331
rect 5640 29297 5674 29318
rect 3715 29235 3724 29269
rect 3724 29235 3749 29269
rect 3789 29235 3794 29269
rect 3794 29235 3823 29269
rect 3863 29235 3864 29269
rect 3864 29235 3897 29269
rect 3937 29235 3968 29269
rect 3968 29235 3971 29269
rect 4011 29235 4037 29269
rect 4037 29235 4045 29269
rect 4085 29235 4106 29269
rect 4106 29235 4119 29269
rect 4159 29235 4175 29269
rect 4175 29235 4193 29269
rect 4232 29235 4244 29269
rect 4244 29235 4266 29269
rect 4305 29235 4313 29269
rect 4313 29235 4339 29269
rect 4378 29235 4382 29269
rect 4382 29235 4412 29269
rect 4451 29235 4485 29269
rect 4524 29235 4554 29269
rect 4554 29235 4558 29269
rect 4597 29235 4623 29269
rect 4623 29235 4631 29269
rect 4670 29235 4692 29269
rect 4692 29235 4704 29269
rect 4743 29235 4761 29269
rect 4761 29235 4777 29269
rect 4816 29235 4830 29269
rect 4830 29235 4850 29269
rect 4889 29235 4899 29269
rect 4899 29235 4923 29269
rect 4962 29235 4968 29269
rect 4968 29235 4996 29269
rect 5035 29235 5037 29269
rect 5037 29235 5069 29269
rect 5108 29235 5141 29269
rect 5141 29235 5142 29269
rect 5181 29235 5210 29269
rect 5210 29235 5215 29269
rect 3082 29210 3116 29226
rect 3082 29192 3116 29210
rect 3082 29142 3116 29154
rect 3082 29120 3116 29142
rect 5640 29250 5674 29256
rect 5640 29222 5674 29250
rect 5640 29148 5674 29181
rect 5640 29147 5674 29148
rect 3715 29105 3724 29139
rect 3724 29105 3749 29139
rect 3792 29105 3794 29139
rect 3794 29105 3826 29139
rect 3869 29105 3899 29139
rect 3899 29105 3903 29139
rect 3946 29105 3968 29139
rect 3968 29105 3980 29139
rect 4023 29105 4037 29139
rect 4037 29105 4057 29139
rect 4100 29105 4106 29139
rect 4106 29105 4134 29139
rect 4177 29105 4209 29139
rect 4209 29105 4211 29139
rect 4254 29105 4278 29139
rect 4278 29105 4288 29139
rect 4330 29105 4347 29139
rect 4347 29105 4364 29139
rect 4515 29105 4520 29139
rect 4520 29105 4549 29139
rect 4590 29105 4623 29139
rect 4623 29105 4624 29139
rect 4665 29105 4692 29139
rect 4692 29105 4699 29139
rect 4740 29105 4761 29139
rect 4761 29105 4774 29139
rect 4815 29105 4830 29139
rect 4830 29105 4849 29139
rect 4890 29105 4899 29139
rect 4899 29105 4924 29139
rect 4965 29105 4968 29139
rect 4968 29105 4999 29139
rect 5040 29105 5072 29139
rect 5072 29105 5074 29139
rect 5115 29105 5141 29139
rect 5141 29105 5149 29139
rect 5189 29105 5210 29139
rect 5210 29105 5223 29139
rect 3082 29074 3116 29082
rect 3082 29048 3116 29074
rect 3082 29006 3116 29010
rect 3082 28976 3116 29006
rect 3082 28904 3116 28938
rect 3082 28836 3116 28866
rect 3082 28832 3116 28836
rect 3082 28768 3116 28794
rect 3082 28760 3116 28768
rect 3082 28700 3116 28722
rect 3082 28688 3116 28700
rect 3082 28632 3116 28650
rect 3082 28616 3116 28632
rect 3082 28564 3116 28578
rect 3082 28544 3116 28564
rect 3082 28496 3116 28506
rect 3082 28472 3116 28496
rect 5640 29080 5674 29106
rect 5640 29072 5674 29080
rect 5640 29012 5674 29031
rect 5640 28997 5674 29012
rect 5640 28944 5674 28956
rect 5640 28922 5674 28944
rect 5640 28876 5674 28881
rect 5640 28847 5674 28876
rect 5640 28774 5674 28806
rect 5640 28772 5674 28774
rect 5640 28706 5674 28731
rect 5640 28697 5674 28706
rect 5640 28638 5674 28656
rect 5640 28622 5674 28638
rect 5640 28570 5674 28581
rect 5640 28547 5674 28570
rect 5640 28502 5674 28506
rect 5640 28472 5674 28502
rect 3154 28400 3184 28434
rect 3184 28400 3188 28434
rect 3228 28400 3252 28434
rect 3252 28400 3262 28434
rect 3302 28400 3320 28434
rect 3320 28400 3336 28434
rect 3376 28400 3388 28434
rect 3388 28400 3410 28434
rect 3450 28400 3456 28434
rect 3456 28400 3484 28434
rect 3523 28400 3524 28434
rect 3524 28400 3557 28434
rect 3596 28400 3626 28434
rect 3626 28400 3630 28434
rect 3669 28400 3694 28434
rect 3694 28400 3703 28434
rect 3742 28400 3762 28434
rect 3762 28400 3776 28434
rect 3815 28400 3830 28434
rect 3830 28400 3849 28434
rect 3888 28400 3898 28434
rect 3898 28400 3922 28434
rect 3961 28400 3966 28434
rect 3966 28400 3995 28434
rect 4034 28400 4068 28434
rect 4107 28400 4136 28434
rect 4136 28400 4141 28434
rect 4180 28400 4204 28434
rect 4204 28400 4214 28434
rect 4253 28400 4272 28434
rect 4272 28400 4287 28434
rect 4326 28400 4340 28434
rect 4340 28400 4360 28434
rect 4399 28400 4408 28434
rect 4408 28400 4433 28434
rect 4472 28400 4476 28434
rect 4476 28400 4506 28434
rect 4545 28400 4578 28434
rect 4578 28400 4579 28434
rect 4618 28400 4646 28434
rect 4646 28400 4652 28434
rect 4691 28400 4714 28434
rect 4714 28400 4725 28434
rect 4764 28400 4782 28434
rect 4782 28400 4798 28434
rect 4837 28400 4850 28434
rect 4850 28400 4871 28434
rect 4910 28400 4918 28434
rect 4918 28400 4944 28434
rect 4983 28400 4986 28434
rect 4986 28400 5017 28434
rect 5056 28400 5088 28434
rect 5088 28400 5090 28434
rect 5129 28400 5156 28434
rect 5156 28400 5163 28434
rect 5202 28400 5224 28434
rect 5224 28400 5236 28434
rect 5275 28400 5292 28434
rect 5292 28400 5309 28434
rect 5348 28400 5360 28434
rect 5360 28400 5382 28434
rect 5421 28400 5428 28434
rect 5428 28400 5455 28434
rect 5494 28400 5496 28434
rect 5496 28400 5528 28434
rect 5567 28400 5601 28434
rect 7746 29840 7780 29852
rect 7746 29818 7780 29840
rect 7746 29772 7780 29779
rect 7746 29745 7780 29772
rect 7746 29704 7780 29706
rect 7746 29672 7780 29704
rect 7746 29602 7780 29633
rect 7746 29599 7780 29602
rect 7746 29534 7780 29560
rect 7746 29526 7780 29534
rect 7746 29466 7780 29487
rect 7746 29453 7780 29466
rect 7746 29398 7780 29414
rect 7746 29380 7780 29398
rect 7746 29330 7780 29341
rect 7746 29307 7780 29330
rect 7746 29262 7780 29268
rect 7746 29234 7780 29262
rect 7746 29194 7780 29195
rect 7746 29161 7780 29194
rect 7746 29092 7780 29122
rect 7746 29088 7780 29092
rect 7746 29024 7780 29049
rect 7746 29015 7780 29024
rect 7746 28956 7780 28976
rect 7746 28942 7780 28956
rect 7746 28888 7780 28903
rect 7746 28869 7780 28888
rect 7746 28820 7780 28830
rect 7746 28796 7780 28820
rect 7746 28752 7780 28757
rect 7746 28723 7780 28752
rect 7746 28650 7780 28684
rect 7746 28582 7780 28611
rect 7746 28577 7780 28582
rect 7746 28514 7780 28538
rect 7746 28504 7780 28514
rect 7746 28446 7780 28465
rect 7746 28431 7780 28446
rect 2822 28382 2856 28390
rect 2822 28356 2856 28382
rect 2822 28284 2856 28318
rect 2822 28232 2856 28246
rect 2822 28212 2856 28232
rect 7746 28378 7780 28392
rect 7746 28358 7780 28378
rect 7746 28310 7780 28319
rect 7746 28285 7780 28310
rect 7746 28242 7780 28246
rect 7746 28212 7780 28242
rect 2894 28140 2924 28174
rect 2924 28140 2928 28174
rect 2967 28140 2992 28174
rect 2992 28140 3001 28174
rect 3040 28140 3060 28174
rect 3060 28140 3074 28174
rect 3113 28140 3128 28174
rect 3128 28140 3147 28174
rect 3186 28140 3196 28174
rect 3196 28140 3220 28174
rect 3259 28140 3264 28174
rect 3264 28140 3293 28174
rect 3332 28140 3366 28174
rect 3405 28140 3434 28174
rect 3434 28140 3439 28174
rect 3478 28140 3502 28174
rect 3502 28140 3512 28174
rect 3551 28140 3570 28174
rect 3570 28140 3585 28174
rect 3624 28140 3638 28174
rect 3638 28140 3658 28174
rect 3697 28140 3706 28174
rect 3706 28140 3731 28174
rect 3770 28140 3774 28174
rect 3774 28140 3804 28174
rect 3843 28140 3876 28174
rect 3876 28140 3877 28174
rect 3916 28140 3944 28174
rect 3944 28140 3950 28174
rect 3989 28140 4012 28174
rect 4012 28140 4023 28174
rect 4062 28140 4080 28174
rect 4080 28140 4096 28174
rect 4135 28140 4148 28174
rect 4148 28140 4169 28174
rect 4208 28140 4216 28174
rect 4216 28140 4242 28174
rect 4281 28140 4284 28174
rect 4284 28140 4315 28174
rect 4354 28140 4386 28174
rect 4386 28140 4388 28174
rect 4427 28140 4454 28174
rect 4454 28140 4461 28174
rect 4500 28140 4522 28174
rect 4522 28140 4534 28174
rect 4573 28140 4590 28174
rect 4590 28140 4607 28174
rect 4646 28140 4658 28174
rect 4658 28140 4680 28174
rect 4719 28140 4726 28174
rect 4726 28140 4753 28174
rect 4792 28140 4794 28174
rect 4794 28140 4826 28174
rect 4865 28140 4896 28174
rect 4896 28140 4899 28174
rect 4938 28140 4964 28174
rect 4964 28140 4972 28174
rect 5010 28140 5032 28174
rect 5032 28140 5044 28174
rect 5082 28140 5100 28174
rect 5100 28140 5116 28174
rect 5154 28140 5168 28174
rect 5168 28140 5188 28174
rect 5226 28140 5236 28174
rect 5236 28140 5260 28174
rect 5298 28140 5304 28174
rect 5304 28140 5332 28174
rect 5370 28140 5372 28174
rect 5372 28140 5404 28174
rect 5442 28140 5474 28174
rect 5474 28140 5476 28174
rect 5514 28140 5542 28174
rect 5542 28140 5548 28174
rect 5586 28140 5610 28174
rect 5610 28140 5620 28174
rect 5658 28140 5678 28174
rect 5678 28140 5692 28174
rect 5730 28140 5746 28174
rect 5746 28140 5764 28174
rect 5802 28140 5814 28174
rect 5814 28140 5836 28174
rect 5874 28140 5882 28174
rect 5882 28140 5908 28174
rect 5946 28140 5950 28174
rect 5950 28140 5980 28174
rect 6018 28140 6052 28174
rect 6090 28140 6120 28174
rect 6120 28140 6124 28174
rect 6162 28140 6188 28174
rect 6188 28140 6196 28174
rect 6234 28140 6256 28174
rect 6256 28140 6268 28174
rect 6306 28140 6324 28174
rect 6324 28140 6340 28174
rect 6378 28140 6392 28174
rect 6392 28140 6412 28174
rect 6450 28140 6460 28174
rect 6460 28140 6484 28174
rect 6522 28140 6528 28174
rect 6528 28140 6556 28174
rect 6594 28140 6596 28174
rect 6596 28140 6628 28174
rect 6666 28140 6698 28174
rect 6698 28140 6700 28174
rect 6738 28140 6766 28174
rect 6766 28140 6772 28174
rect 6810 28140 6834 28174
rect 6834 28140 6844 28174
rect 6882 28140 6902 28174
rect 6902 28140 6916 28174
rect 6954 28140 6970 28174
rect 6970 28140 6988 28174
rect 7026 28140 7038 28174
rect 7038 28140 7060 28174
rect 7098 28140 7106 28174
rect 7106 28140 7132 28174
rect 7170 28140 7174 28174
rect 7174 28140 7204 28174
rect 7242 28140 7276 28174
rect 7314 28140 7344 28174
rect 7344 28140 7348 28174
rect 7386 28140 7412 28174
rect 7412 28140 7420 28174
rect 7458 28140 7480 28174
rect 7480 28140 7492 28174
rect 7530 28140 7548 28174
rect 7548 28140 7564 28174
rect 7602 28140 7616 28174
rect 7616 28140 7636 28174
rect 7674 28140 7684 28174
rect 7684 28140 7708 28174
rect 4980 26165 5014 26199
rect 5059 26165 5084 26199
rect 5084 26165 5093 26199
rect 5138 26165 5154 26199
rect 5154 26165 5172 26199
rect 5217 26165 5224 26199
rect 5224 26165 5251 26199
rect 5295 26165 5329 26199
rect 5373 26165 5400 26199
rect 5400 26165 5407 26199
rect 5451 26165 5470 26199
rect 5470 26165 5485 26199
rect 5529 26165 5540 26199
rect 5540 26165 5563 26199
rect 4008 26082 4042 26116
rect 4008 26014 4042 26041
rect 4008 26007 4042 26014
rect 4008 25946 4042 25966
rect 4008 25932 4042 25946
rect 4008 25878 4042 25891
rect 4008 25857 4042 25878
rect 4008 25810 4042 25816
rect 4008 25782 4042 25810
rect 4008 25708 4042 25740
rect 4008 25706 4042 25708
rect 2850 25651 2882 25685
rect 2882 25651 2884 25685
rect 2928 25651 2950 25685
rect 2950 25651 2962 25685
rect 3005 25651 3018 25685
rect 3018 25651 3039 25685
rect 3082 25651 3086 25685
rect 3086 25651 3116 25685
rect 3159 25651 3188 25685
rect 3188 25651 3193 25685
rect 3236 25651 3256 25685
rect 3256 25651 3270 25685
rect 3313 25651 3324 25685
rect 3324 25651 3347 25685
rect 3390 25651 3392 25685
rect 3392 25651 3424 25685
rect 3467 25651 3494 25685
rect 3494 25651 3501 25685
rect 3544 25651 3562 25685
rect 3562 25651 3578 25685
rect 3621 25651 3630 25685
rect 3630 25651 3655 25685
rect 3698 25609 3732 25613
rect 3698 25579 3732 25609
rect 3698 25507 3732 25540
rect 3698 25506 3732 25507
rect 2832 25472 2866 25506
rect 2904 25472 2938 25506
rect 3536 25472 3570 25506
rect 3608 25472 3642 25506
rect 3698 25439 3732 25467
rect 3698 25433 3732 25439
rect 3698 25371 3732 25394
rect 3698 25360 3732 25371
rect 3698 25303 3732 25321
rect 3698 25287 3732 25303
rect 3698 25235 3732 25248
rect 3698 25214 3732 25235
rect 3698 25167 3732 25175
rect 3698 25141 3732 25167
rect 3698 25099 3732 25102
rect 3698 25068 3732 25099
rect 3698 24997 3732 25029
rect 3698 24995 3732 24997
rect 3698 24929 3732 24956
rect 3698 24922 3732 24929
rect 3698 24861 3732 24883
rect 3698 24849 3732 24861
rect 3698 24793 3732 24810
rect 3698 24776 3732 24793
rect 3698 24725 3732 24737
rect 3698 24703 3732 24725
rect 4008 25640 4042 25664
rect 4008 25630 4042 25640
rect 4008 25572 4042 25588
rect 4008 25554 4042 25572
rect 4008 25504 4042 25512
rect 4008 25478 4042 25504
rect 4008 25402 4042 25436
rect 4008 25334 4042 25360
rect 4008 25326 4042 25334
rect 4008 25266 4042 25284
rect 4008 25250 4042 25266
rect 4008 25198 4042 25208
rect 4008 25174 4042 25198
rect 4008 25130 4042 25132
rect 4008 25098 4042 25130
rect 4008 25028 4042 25056
rect 4008 25022 4042 25028
rect 4008 24960 4042 24980
rect 4008 24946 4042 24960
rect 4008 24892 4042 24904
rect 4008 24870 4042 24892
rect 4008 24824 4042 24828
rect 4008 24794 4042 24824
rect 4008 24718 4042 24752
rect 4353 26037 4387 26071
rect 4353 25964 4387 25998
rect 4353 25891 4387 25925
rect 4353 25818 4387 25852
rect 4353 25745 4387 25779
rect 4353 25672 4387 25706
rect 4353 25599 4387 25633
rect 4353 25526 4387 25560
rect 4353 25453 4387 25487
rect 4353 25379 4387 25413
rect 4353 25305 4387 25339
rect 4353 25231 4387 25265
rect 4353 25157 4387 25191
rect 4353 25083 4387 25117
rect 4353 25009 4387 25043
rect 4353 24935 4387 24969
rect 4353 24861 4387 24895
rect 4353 24787 4387 24821
rect 4353 24713 4387 24747
rect 4509 26037 4543 26071
rect 4509 25964 4543 25998
rect 4509 25891 4543 25925
rect 4509 25818 4543 25852
rect 4509 25745 4543 25779
rect 4509 25672 4543 25706
rect 4509 25599 4543 25633
rect 4509 25526 4543 25560
rect 4509 25453 4543 25487
rect 4509 25379 4543 25413
rect 4509 25305 4543 25339
rect 4509 25231 4543 25265
rect 4509 25157 4543 25191
rect 4509 25083 4543 25117
rect 4509 25009 4543 25043
rect 4509 24935 4543 24969
rect 4509 24861 4543 24895
rect 4509 24787 4543 24821
rect 4509 24713 4543 24747
rect 4665 26037 4699 26071
rect 4665 25964 4699 25998
rect 4665 25891 4699 25925
rect 4665 25818 4699 25852
rect 4665 25745 4699 25779
rect 4665 25672 4699 25706
rect 4665 25599 4699 25633
rect 4665 25526 4699 25560
rect 4665 25453 4699 25487
rect 4665 25379 4699 25413
rect 4665 25305 4699 25339
rect 4665 25231 4699 25265
rect 4665 25157 4699 25191
rect 4665 25083 4699 25117
rect 4665 25009 4699 25043
rect 4665 24935 4699 24969
rect 4665 24861 4699 24895
rect 4665 24787 4699 24821
rect 4665 24713 4699 24747
rect 4821 26037 4855 26071
rect 4821 25964 4855 25998
rect 4821 25891 4855 25925
rect 4821 25818 4855 25852
rect 4821 25745 4855 25779
rect 4821 25672 4855 25706
rect 4821 25599 4855 25633
rect 4821 25526 4855 25560
rect 4821 25453 4855 25487
rect 4821 25379 4855 25413
rect 4821 25305 4855 25339
rect 4821 25231 4855 25265
rect 4821 25157 4855 25191
rect 4821 25083 4855 25117
rect 4821 25009 4855 25043
rect 4821 24935 4855 24969
rect 4821 24861 4855 24895
rect 4821 24787 4855 24821
rect 4821 24713 4855 24747
rect 4977 26037 5011 26071
rect 4977 25964 5011 25998
rect 4977 25891 5011 25925
rect 4977 25818 5011 25852
rect 4977 25745 5011 25779
rect 4977 25672 5011 25706
rect 4977 25599 5011 25633
rect 4977 25526 5011 25560
rect 4977 25453 5011 25487
rect 4977 25379 5011 25413
rect 4977 25305 5011 25339
rect 4977 25231 5011 25265
rect 4977 25157 5011 25191
rect 4977 25083 5011 25117
rect 4977 25009 5011 25043
rect 4977 24935 5011 24969
rect 4977 24861 5011 24895
rect 4977 24787 5011 24821
rect 4977 24713 5011 24747
rect 5133 26037 5167 26071
rect 5133 25964 5167 25998
rect 5133 25891 5167 25925
rect 5133 25818 5167 25852
rect 5133 25745 5167 25779
rect 5133 25672 5167 25706
rect 5133 25599 5167 25633
rect 5133 25526 5167 25560
rect 5133 25453 5167 25487
rect 5133 25379 5167 25413
rect 5133 25305 5167 25339
rect 5133 25231 5167 25265
rect 5133 25157 5167 25191
rect 5133 25083 5167 25117
rect 5133 25009 5167 25043
rect 5133 24935 5167 24969
rect 5133 24861 5167 24895
rect 5133 24787 5167 24821
rect 5133 24713 5167 24747
rect 5289 26037 5323 26071
rect 5289 25964 5323 25998
rect 5289 25891 5323 25925
rect 5289 25818 5323 25852
rect 5289 25745 5323 25779
rect 5289 25672 5323 25706
rect 5289 25599 5323 25633
rect 5289 25526 5323 25560
rect 5289 25453 5323 25487
rect 5289 25379 5323 25413
rect 5289 25305 5323 25339
rect 5289 25231 5323 25265
rect 5289 25157 5323 25191
rect 5289 25083 5323 25117
rect 5289 25009 5323 25043
rect 5289 24935 5323 24969
rect 5289 24861 5323 24895
rect 5289 24787 5323 24821
rect 5289 24713 5323 24747
rect 5445 26037 5479 26071
rect 5445 25964 5479 25998
rect 5445 25891 5479 25925
rect 5445 25818 5479 25852
rect 5445 25745 5479 25779
rect 5445 25672 5479 25706
rect 5445 25599 5479 25633
rect 5445 25526 5479 25560
rect 5445 25453 5479 25487
rect 5445 25379 5479 25413
rect 5445 25305 5479 25339
rect 5445 25231 5479 25265
rect 5445 25157 5479 25191
rect 5445 25083 5479 25117
rect 5445 25009 5479 25043
rect 5445 24935 5479 24969
rect 5445 24861 5479 24895
rect 5445 24787 5479 24821
rect 5445 24713 5479 24747
rect 5601 26037 5635 26071
rect 5601 25964 5635 25998
rect 5601 25891 5635 25925
rect 5601 25818 5635 25852
rect 5601 25745 5635 25779
rect 5601 25672 5635 25706
rect 5601 25599 5635 25633
rect 5601 25526 5635 25560
rect 5601 25453 5635 25487
rect 5601 25379 5635 25413
rect 5601 25305 5635 25339
rect 5601 25231 5635 25265
rect 5601 25157 5635 25191
rect 5601 25083 5635 25117
rect 5601 25009 5635 25043
rect 5601 24935 5635 24969
rect 5601 24861 5635 24895
rect 5601 24787 5635 24821
rect 5601 24713 5635 24747
rect 5946 26048 5980 26071
rect 5946 26037 5980 26048
rect 5946 25980 5980 25998
rect 5946 25964 5980 25980
rect 5946 25912 5980 25925
rect 5946 25891 5980 25912
rect 5946 25844 5980 25852
rect 5946 25818 5980 25844
rect 5946 25776 5980 25779
rect 5946 25745 5980 25776
rect 5946 25674 5980 25706
rect 5946 25672 5980 25674
rect 5946 25606 5980 25633
rect 5946 25599 5980 25606
rect 5946 25538 5980 25560
rect 5946 25526 5980 25538
rect 5946 25470 5980 25487
rect 5946 25453 5980 25470
rect 5946 25402 5980 25413
rect 5946 25379 5980 25402
rect 5946 25334 5980 25339
rect 5946 25305 5980 25334
rect 5946 25232 5980 25265
rect 5946 25231 5980 25232
rect 5946 25164 5980 25191
rect 5946 25157 5980 25164
rect 5946 25096 5980 25117
rect 5946 25083 5980 25096
rect 5946 25028 5980 25043
rect 5946 25009 5980 25028
rect 5946 24960 5980 24969
rect 5946 24935 5980 24960
rect 5946 24892 5980 24895
rect 5946 24861 5980 24892
rect 5946 24790 5980 24821
rect 5946 24787 5980 24790
rect 5946 24713 5980 24747
rect 3698 24657 3732 24664
rect 3698 24630 3732 24657
rect 3698 24589 3732 24591
rect 3698 24557 3732 24589
rect 3698 24487 3732 24518
rect 3698 24484 3732 24487
rect 3698 24419 3732 24445
rect 3698 24411 3732 24419
rect 3698 24351 3732 24372
rect 3698 24338 3732 24351
rect 3698 24283 3732 24299
rect 3698 24265 3732 24283
rect 3698 24215 3732 24226
rect 3698 24192 3732 24215
rect 3698 24147 3732 24153
rect 3698 24119 3732 24147
rect 3698 24079 3732 24080
rect 3698 24046 3732 24079
rect 3698 23977 3732 24007
rect 3698 23973 3732 23977
rect 3698 23909 3732 23934
rect 3698 23900 3732 23909
rect 3698 23841 3732 23861
rect 3698 23827 3732 23841
rect 3698 23773 3732 23788
rect 3698 23754 3732 23773
rect 3698 23705 3732 23715
rect 3698 23681 3732 23705
rect 3698 23637 3732 23642
rect 3698 23608 3732 23637
rect 3698 23535 3732 23569
rect 3698 23467 3732 23496
rect 3698 23462 3732 23467
rect 3698 23399 3732 23423
rect 3698 23389 3732 23399
rect 3698 23331 3732 23350
rect 3698 23316 3732 23331
rect 3698 23263 3732 23277
rect 3698 23243 3732 23263
rect 3698 23195 3732 23204
rect 3698 23170 3732 23195
rect 3698 23127 3732 23131
rect 3698 23097 3732 23127
rect 3698 23025 3732 23058
rect 3698 23024 3732 23025
rect 3698 22957 3732 22985
rect 3698 22951 3732 22957
rect 3698 22889 3732 22912
rect 3698 22878 3732 22889
rect 3698 22821 3732 22839
rect 3698 22805 3732 22821
rect 3698 22753 3732 22766
rect 3698 22732 3732 22753
rect 3698 22685 3732 22693
rect 3698 22659 3732 22685
rect 3698 22617 3732 22621
rect 3698 22587 3732 22617
rect 3698 22515 3732 22549
rect 3698 22447 3732 22477
rect 3698 22443 3732 22447
rect 3698 22379 3732 22405
rect 3698 22371 3732 22379
rect 3698 22311 3732 22333
rect 3698 22299 3732 22311
rect 3698 22243 3732 22261
rect 3698 22227 3732 22243
rect 3698 22175 3732 22189
rect 3698 22155 3732 22175
rect 3698 22107 3732 22117
rect 3698 22083 3732 22107
rect 3698 22039 3732 22045
rect 3698 22011 3732 22039
rect 3698 21971 3732 21973
rect 3698 21939 3732 21971
rect 3698 21869 3732 21901
rect 3698 21867 3732 21869
rect 3698 21801 3732 21829
rect 3698 21795 3732 21801
rect 3698 21733 3732 21757
rect 3698 21723 3732 21733
rect 3698 21665 3732 21685
rect 3698 21651 3732 21665
rect 3698 21597 3732 21613
rect 3698 21579 3732 21597
rect 3698 21529 3732 21541
rect 3698 21507 3732 21529
rect 3698 21461 3732 21469
rect 3698 21435 3732 21461
rect 3698 21393 3732 21397
rect 3698 21363 3732 21393
rect 3698 21291 3732 21325
rect 3698 21223 3732 21253
rect 3698 21219 3732 21223
rect 3698 21155 3732 21181
rect 3698 21147 3732 21155
rect 3698 21087 3732 21109
rect 3698 21075 3732 21087
rect 3698 21019 3732 21037
rect 3698 21003 3732 21019
rect 3698 20951 3732 20965
rect 3698 20931 3732 20951
rect 3698 20883 3732 20893
rect 3698 20859 3732 20883
rect 3698 20815 3732 20821
rect 3698 20787 3732 20815
rect 3698 20747 3732 20749
rect 3698 20715 3732 20747
rect 3698 20645 3732 20677
rect 3698 20643 3732 20645
rect 3698 20577 3732 20605
rect 3698 20571 3732 20577
rect 3698 20509 3732 20533
rect 3698 20499 3732 20509
rect 3698 20441 3732 20461
rect 3698 20427 3732 20441
rect 3698 20373 3732 20389
rect 3698 20355 3732 20373
rect 3698 20305 3732 20317
rect 3698 20283 3732 20305
rect 3698 20237 3732 20245
rect 3698 20211 3732 20237
rect 3698 20169 3732 20173
rect 3698 20139 3732 20169
rect 3698 20067 3732 20101
rect 3698 19999 3732 20029
rect 3698 19995 3732 19999
rect 3698 19931 3732 19957
rect 3698 19923 3732 19931
rect 3698 19863 3732 19885
rect 3698 19851 3732 19863
rect 3698 19795 3732 19813
rect 3698 19779 3732 19795
rect 3698 19727 3732 19741
rect 3698 19707 3732 19727
rect 3698 19659 3732 19669
rect 3698 19635 3732 19659
rect 3698 19591 3732 19597
rect 3698 19563 3732 19591
rect 3698 19523 3732 19525
rect 3698 19491 3732 19523
rect 3698 19421 3732 19453
rect 3698 19419 3732 19421
rect 3698 19353 3732 19381
rect 3698 19347 3732 19353
rect 3698 19285 3732 19309
rect 3698 19275 3732 19285
rect 3698 19217 3732 19237
rect 3698 19203 3732 19217
rect 3698 19149 3732 19165
rect 3698 19131 3732 19149
rect 3698 19081 3732 19093
rect 3698 19059 3732 19081
rect 3698 19013 3732 19021
rect 3698 18987 3732 19013
rect 3698 18945 3732 18949
rect 3698 18915 3732 18945
rect 3698 18843 3732 18877
rect 3698 18775 3732 18805
rect 3698 18771 3732 18775
rect 3698 18707 3732 18733
rect 3698 18699 3732 18707
rect 3698 18639 3732 18661
rect 3698 18627 3732 18639
rect 3698 18571 3732 18589
rect 3698 18555 3732 18571
rect 4555 24150 4562 24184
rect 4562 24150 4589 24184
rect 4687 24150 4698 24184
rect 4698 24150 4721 24184
rect 4760 24150 4766 24184
rect 4766 24150 4794 24184
rect 4833 24150 4834 24184
rect 4834 24150 4867 24184
rect 4906 24150 4936 24184
rect 4936 24150 4940 24184
rect 4979 24150 5004 24184
rect 5004 24150 5013 24184
rect 5052 24150 5072 24184
rect 5072 24150 5086 24184
rect 5125 24150 5140 24184
rect 5140 24150 5159 24184
rect 5198 24150 5208 24184
rect 5208 24150 5232 24184
rect 5271 24150 5276 24184
rect 5276 24150 5305 24184
rect 5344 24150 5378 24184
rect 5417 24150 5446 24184
rect 5446 24150 5451 24184
rect 5490 24150 5514 24184
rect 5514 24150 5524 24184
rect 5564 24150 5582 24184
rect 5582 24150 5598 24184
rect 5638 24150 5650 24184
rect 5650 24150 5672 24184
rect 5712 24150 5718 24184
rect 5718 24150 5746 24184
rect 5786 24150 5820 24184
rect 4460 24110 4494 24112
rect 4460 24078 4494 24110
rect 4460 24005 4494 24039
rect 4460 23956 4494 23966
rect 4460 23932 4494 23956
rect 4460 23888 4494 23893
rect 4460 23859 4494 23888
rect 5858 24082 5892 24112
rect 5858 24078 5892 24082
rect 5858 24014 5892 24040
rect 5858 24006 5892 24014
rect 5858 23946 5892 23968
rect 5858 23934 5892 23946
rect 5858 23878 5892 23896
rect 5858 23862 5892 23878
rect 4460 23786 4494 23820
rect 4460 23718 4494 23747
rect 4460 23713 4494 23718
rect 4651 23800 4685 23834
rect 4731 23800 4765 23834
rect 4810 23800 4844 23834
rect 4651 23728 4685 23762
rect 4731 23728 4765 23762
rect 4810 23728 4844 23762
rect 5060 23830 5166 23854
rect 5060 23796 5102 23830
rect 5102 23796 5136 23830
rect 5136 23796 5166 23830
rect 5060 23748 5166 23796
rect 5315 23830 5421 23848
rect 5315 23796 5358 23830
rect 5358 23796 5392 23830
rect 5392 23796 5421 23830
rect 5315 23742 5421 23796
rect 5858 23810 5892 23824
rect 5858 23790 5892 23810
rect 5858 23742 5892 23752
rect 5858 23718 5892 23742
rect 4460 23650 4494 23674
rect 4460 23640 4494 23650
rect 4460 23582 4494 23601
rect 4460 23567 4494 23582
rect 4460 23514 4494 23528
rect 4460 23494 4494 23514
rect 4460 23446 4494 23455
rect 4460 23421 4494 23446
rect 4460 23378 4494 23382
rect 4460 23348 4494 23378
rect 4460 23276 4494 23309
rect 4460 23275 4494 23276
rect 4460 23208 4494 23236
rect 4460 23202 4494 23208
rect 4460 23140 4494 23163
rect 4460 23129 4494 23140
rect 4460 23072 4494 23090
rect 4460 23056 4494 23072
rect 4460 23004 4494 23017
rect 4460 22983 4494 23004
rect 4460 22936 4494 22944
rect 4460 22910 4494 22936
rect 4460 22868 4494 22871
rect 4460 22837 4494 22868
rect 4460 22766 4494 22798
rect 4460 22764 4494 22766
rect 4460 22698 4494 22725
rect 4460 22691 4494 22698
rect 4460 22630 4494 22652
rect 4460 22618 4494 22630
rect 4460 22562 4494 22579
rect 4460 22545 4494 22562
rect 4460 22494 4494 22506
rect 4460 22472 4494 22494
rect 4460 22426 4494 22433
rect 4460 22399 4494 22426
rect 4460 22358 4494 22360
rect 4460 22326 4494 22358
rect 4460 22256 4494 22287
rect 4460 22253 4494 22256
rect 4460 22188 4494 22214
rect 4460 22180 4494 22188
rect 4460 22120 4494 22141
rect 4460 22107 4494 22120
rect 4888 23631 4922 23660
rect 4888 23626 4922 23631
rect 4888 23561 4922 23587
rect 4888 23553 4922 23561
rect 4888 23491 4922 23514
rect 4888 23480 4922 23491
rect 4888 23421 4922 23441
rect 4888 23407 4922 23421
rect 4888 23351 4922 23368
rect 4888 23334 4922 23351
rect 4888 23281 4922 23295
rect 4888 23261 4922 23281
rect 4888 23211 4922 23222
rect 4888 23188 4922 23211
rect 4888 23141 4922 23149
rect 4888 23115 4922 23141
rect 4888 23071 4922 23076
rect 4888 23042 4922 23071
rect 4888 23001 4922 23003
rect 4888 22969 4922 23001
rect 4888 22897 4922 22930
rect 4888 22896 4922 22897
rect 4888 22827 4922 22857
rect 4888 22823 4922 22827
rect 4888 22757 4922 22784
rect 4888 22750 4922 22757
rect 4888 22687 4922 22711
rect 4888 22677 4922 22687
rect 4888 22617 4922 22638
rect 4888 22604 4922 22617
rect 4888 22547 4922 22565
rect 4888 22531 4922 22547
rect 4888 22478 4922 22492
rect 4888 22458 4922 22478
rect 4888 22409 4922 22419
rect 4888 22385 4922 22409
rect 4888 22340 4922 22346
rect 4888 22312 4922 22340
rect 4888 22271 4922 22273
rect 4888 22239 4922 22271
rect 4888 22167 4922 22200
rect 4888 22166 4922 22167
rect 4642 22072 4676 22106
rect 4715 22072 4749 22106
rect 4788 22072 4822 22106
rect 4888 22098 4922 22127
rect 4888 22093 4922 22098
rect 4460 22052 4494 22068
rect 4460 22034 4494 22052
rect 4460 21984 4494 21995
rect 4460 21961 4494 21984
rect 4460 21916 4494 21922
rect 4460 21888 4494 21916
rect 4460 21848 4494 21849
rect 4460 21815 4494 21848
rect 4460 21746 4494 21776
rect 4460 21742 4494 21746
rect 4460 21678 4494 21703
rect 4460 21669 4494 21678
rect 4460 21610 4494 21630
rect 4460 21596 4494 21610
rect 4460 21542 4494 21557
rect 4460 21523 4494 21542
rect 4460 21474 4494 21484
rect 4460 21450 4494 21474
rect 4460 21406 4494 21411
rect 4460 21377 4494 21406
rect 4460 21304 4494 21338
rect 4460 21236 4494 21265
rect 4460 21231 4494 21236
rect 4460 21168 4494 21192
rect 4460 21158 4494 21168
rect 4460 21100 4494 21119
rect 4460 21085 4494 21100
rect 4460 21032 4494 21046
rect 4460 21012 4494 21032
rect 4460 20964 4494 20973
rect 4460 20939 4494 20964
rect 4460 20896 4494 20900
rect 4460 20866 4494 20896
rect 4460 20794 4494 20827
rect 4460 20793 4494 20794
rect 4460 20726 4494 20754
rect 4460 20720 4494 20726
rect 4460 20658 4494 20681
rect 4460 20647 4494 20658
rect 4460 20590 4494 20608
rect 4460 20574 4494 20590
rect 4460 20522 4494 20535
rect 4460 20501 4494 20522
rect 4460 20454 4494 20462
rect 4460 20428 4494 20454
rect 4888 22029 4922 22054
rect 4888 22020 4922 22029
rect 4888 21960 4922 21981
rect 4888 21947 4922 21960
rect 4888 21891 4922 21908
rect 4888 21874 4922 21891
rect 4888 21822 4922 21835
rect 4888 21801 4922 21822
rect 4888 21753 4922 21762
rect 4888 21728 4922 21753
rect 4888 21684 4922 21689
rect 4888 21655 4922 21684
rect 4888 21615 4922 21616
rect 4888 21582 4922 21615
rect 4888 21512 4922 21543
rect 4888 21509 4922 21512
rect 4888 21443 4922 21470
rect 4888 21436 4922 21443
rect 4888 21374 4922 21397
rect 4888 21363 4922 21374
rect 4888 21305 4922 21324
rect 4888 21290 4922 21305
rect 4888 21236 4922 21251
rect 4888 21217 4922 21236
rect 4888 21167 4922 21178
rect 4888 21144 4922 21167
rect 4888 21098 4922 21105
rect 4888 21071 4922 21098
rect 4888 21029 4922 21032
rect 4888 20998 4922 21029
rect 4888 20925 4922 20959
rect 4888 20856 4922 20886
rect 4888 20852 4922 20856
rect 4888 20787 4922 20813
rect 4888 20779 4922 20787
rect 4888 20718 4922 20740
rect 4888 20706 4922 20718
rect 4888 20649 4922 20667
rect 4888 20633 4922 20649
rect 4888 20580 4922 20594
rect 4888 20560 4922 20580
rect 4888 20511 4922 20520
rect 4888 20486 4922 20511
rect 5196 23631 5230 23637
rect 5196 23603 5230 23631
rect 5196 23562 5230 23564
rect 5196 23530 5230 23562
rect 5196 23459 5230 23491
rect 5196 23457 5230 23459
rect 5196 23390 5230 23418
rect 5196 23384 5230 23390
rect 5196 23321 5230 23345
rect 5196 23311 5230 23321
rect 5196 23252 5230 23272
rect 5196 23238 5230 23252
rect 5196 23183 5230 23199
rect 5196 23165 5230 23183
rect 5196 23114 5230 23126
rect 5196 23092 5230 23114
rect 5196 23045 5230 23053
rect 5196 23019 5230 23045
rect 5196 22976 5230 22980
rect 5196 22946 5230 22976
rect 5196 22873 5230 22907
rect 5196 22803 5230 22834
rect 5196 22800 5230 22803
rect 5196 22734 5230 22761
rect 5196 22727 5230 22734
rect 5196 22665 5230 22688
rect 5196 22654 5230 22665
rect 5196 22596 5230 22615
rect 5196 22581 5230 22596
rect 5196 22527 5230 22542
rect 5196 22508 5230 22527
rect 5196 22458 5230 22469
rect 5196 22435 5230 22458
rect 5196 22389 5230 22396
rect 5196 22362 5230 22389
rect 5196 22320 5230 22323
rect 5196 22289 5230 22320
rect 5196 22217 5230 22250
rect 5196 22216 5230 22217
rect 5196 22148 5230 22177
rect 5196 22143 5230 22148
rect 5196 22079 5230 22104
rect 5196 22070 5230 22079
rect 5196 22010 5230 22031
rect 5196 21997 5230 22010
rect 5196 21941 5230 21958
rect 5196 21924 5230 21941
rect 5196 21872 5230 21885
rect 5196 21851 5230 21872
rect 5196 21803 5230 21812
rect 5196 21778 5230 21803
rect 5196 21734 5230 21739
rect 5196 21705 5230 21734
rect 5196 21665 5230 21666
rect 5196 21632 5230 21665
rect 5196 21561 5230 21593
rect 5196 21559 5230 21561
rect 5196 21492 5230 21520
rect 5196 21486 5230 21492
rect 5196 21423 5230 21447
rect 5196 21413 5230 21423
rect 5196 21354 5230 21374
rect 5196 21340 5230 21354
rect 5196 21285 5230 21301
rect 5196 21267 5230 21285
rect 5196 21216 5230 21228
rect 5196 21194 5230 21216
rect 5196 21147 5230 21155
rect 5196 21121 5230 21147
rect 5196 21078 5230 21082
rect 5196 21048 5230 21078
rect 5196 20975 5230 21009
rect 5196 20906 5230 20936
rect 5196 20902 5230 20906
rect 5196 20837 5230 20863
rect 5196 20829 5230 20837
rect 5196 20768 5230 20790
rect 5196 20756 5230 20768
rect 5196 20699 5230 20717
rect 5196 20683 5230 20699
rect 5196 20630 5230 20644
rect 5196 20610 5230 20630
rect 5196 20561 5230 20571
rect 5196 20537 5230 20561
rect 5196 20492 5230 20498
rect 5196 20464 5230 20492
rect 4460 20386 4494 20389
rect 4460 20355 4494 20386
rect 4642 20411 4676 20445
rect 4726 20411 4760 20445
rect 4810 20411 4844 20445
rect 4642 20339 4676 20373
rect 4726 20339 4760 20373
rect 4810 20339 4844 20373
rect 5196 20423 5230 20425
rect 5196 20391 5230 20423
rect 4460 20284 4494 20316
rect 4460 20282 4494 20284
rect 4460 20216 4494 20244
rect 4460 20210 4494 20216
rect 4460 20148 4494 20172
rect 4460 20138 4494 20148
rect 4460 20080 4494 20100
rect 4460 20066 4494 20080
rect 5196 20319 5230 20352
rect 5196 20318 5230 20319
rect 5196 20250 5230 20278
rect 5196 20244 5230 20250
rect 5196 20181 5230 20204
rect 5196 20170 5230 20181
rect 5196 20112 5230 20130
rect 5196 20096 5230 20112
rect 4585 20059 4619 20093
rect 4660 20059 4694 20093
rect 4735 20059 4769 20093
rect 4809 20059 4843 20093
rect 4460 20012 4494 20028
rect 4460 19994 4494 20012
rect 4460 19944 4494 19956
rect 4460 19922 4494 19944
rect 4899 20032 4933 20036
rect 4899 20002 4933 20032
rect 4899 19961 4933 19964
rect 4642 19903 4676 19937
rect 4726 19903 4760 19937
rect 4809 19903 4843 19937
rect 4899 19930 4933 19961
rect 4460 19876 4494 19884
rect 4460 19850 4494 19876
rect 4460 19808 4494 19812
rect 4460 19778 4494 19808
rect 4899 19890 4933 19891
rect 4899 19857 4933 19890
rect 4899 19784 4933 19818
rect 4585 19747 4619 19781
rect 4657 19747 4691 19781
rect 4729 19747 4763 19781
rect 4460 19706 4494 19740
rect 4460 19638 4494 19668
rect 4460 19634 4494 19638
rect 4899 19712 4933 19745
rect 5196 20043 5230 20056
rect 5196 20022 5230 20043
rect 5196 19974 5230 19982
rect 5196 19948 5230 19974
rect 5196 19905 5230 19908
rect 5196 19874 5230 19905
rect 5196 19802 5230 19834
rect 5196 19800 5230 19802
rect 5452 23631 5486 23637
rect 5452 23603 5486 23631
rect 5452 23562 5486 23564
rect 5452 23530 5486 23562
rect 5452 23459 5486 23491
rect 5452 23457 5486 23459
rect 5452 23390 5486 23418
rect 5452 23384 5486 23390
rect 5452 23321 5486 23345
rect 5452 23311 5486 23321
rect 5452 23252 5486 23272
rect 5452 23238 5486 23252
rect 5452 23183 5486 23199
rect 5452 23165 5486 23183
rect 5452 23114 5486 23126
rect 5452 23092 5486 23114
rect 5452 23045 5486 23053
rect 5452 23019 5486 23045
rect 5452 22976 5486 22980
rect 5452 22946 5486 22976
rect 5452 22873 5486 22907
rect 5452 22803 5486 22834
rect 5452 22800 5486 22803
rect 5452 22734 5486 22761
rect 5452 22727 5486 22734
rect 5452 22665 5486 22688
rect 5452 22654 5486 22665
rect 5452 22596 5486 22615
rect 5452 22581 5486 22596
rect 5452 22527 5486 22542
rect 5452 22508 5486 22527
rect 5452 22458 5486 22469
rect 5452 22435 5486 22458
rect 5452 22389 5486 22396
rect 5452 22362 5486 22389
rect 5452 22320 5486 22323
rect 5452 22289 5486 22320
rect 5452 22217 5486 22250
rect 5452 22216 5486 22217
rect 5452 22148 5486 22177
rect 5452 22143 5486 22148
rect 5452 22079 5486 22104
rect 5452 22070 5486 22079
rect 5452 22010 5486 22031
rect 5452 21997 5486 22010
rect 5452 21941 5486 21958
rect 5452 21924 5486 21941
rect 5452 21872 5486 21885
rect 5452 21851 5486 21872
rect 5452 21803 5486 21812
rect 5452 21778 5486 21803
rect 5452 21734 5486 21739
rect 5452 21705 5486 21734
rect 5452 21665 5486 21666
rect 5452 21632 5486 21665
rect 5452 21561 5486 21593
rect 5452 21559 5486 21561
rect 5452 21492 5486 21520
rect 5452 21486 5486 21492
rect 5452 21423 5486 21447
rect 5452 21413 5486 21423
rect 5452 21354 5486 21374
rect 5452 21340 5486 21354
rect 5452 21285 5486 21301
rect 5452 21267 5486 21285
rect 5452 21216 5486 21228
rect 5452 21194 5486 21216
rect 5452 21147 5486 21155
rect 5452 21121 5486 21147
rect 5452 21078 5486 21082
rect 5452 21048 5486 21078
rect 5452 20975 5486 21009
rect 5452 20906 5486 20936
rect 5452 20902 5486 20906
rect 5452 20837 5486 20863
rect 5452 20829 5486 20837
rect 5452 20768 5486 20790
rect 5452 20756 5486 20768
rect 5452 20699 5486 20717
rect 5452 20683 5486 20699
rect 5452 20630 5486 20644
rect 5452 20610 5486 20630
rect 5452 20561 5486 20571
rect 5452 20537 5486 20561
rect 5452 20492 5486 20498
rect 5452 20464 5486 20492
rect 5452 20423 5486 20425
rect 5452 20391 5486 20423
rect 5452 20319 5486 20352
rect 5452 20318 5486 20319
rect 5452 20250 5486 20278
rect 5452 20244 5486 20250
rect 5452 20181 5486 20204
rect 5452 20170 5486 20181
rect 5452 20112 5486 20130
rect 5452 20096 5486 20112
rect 5452 20043 5486 20056
rect 5452 20022 5486 20043
rect 5452 19974 5486 19982
rect 5452 19948 5486 19974
rect 5452 19905 5486 19908
rect 5452 19874 5486 19905
rect 5452 19802 5486 19834
rect 5452 19800 5486 19802
rect 5858 23674 5892 23680
rect 5858 23646 5892 23674
rect 5858 23606 5892 23608
rect 5858 23574 5892 23606
rect 5858 23504 5892 23536
rect 5858 23502 5892 23504
rect 5858 23436 5892 23464
rect 5858 23430 5892 23436
rect 5858 23368 5892 23392
rect 5858 23358 5892 23368
rect 5858 23300 5892 23320
rect 5858 23286 5892 23300
rect 5858 23232 5892 23248
rect 5858 23214 5892 23232
rect 5858 23164 5892 23176
rect 5858 23142 5892 23164
rect 5858 23096 5892 23104
rect 5858 23070 5892 23096
rect 5858 23028 5892 23032
rect 5858 22998 5892 23028
rect 5858 22926 5892 22960
rect 5858 22858 5892 22888
rect 5858 22854 5892 22858
rect 5858 22790 5892 22816
rect 5858 22782 5892 22790
rect 5858 22722 5892 22744
rect 5858 22710 5892 22722
rect 5858 22654 5892 22672
rect 5858 22638 5892 22654
rect 5858 22586 5892 22600
rect 5858 22566 5892 22586
rect 5858 22518 5892 22528
rect 5858 22494 5892 22518
rect 5858 22450 5892 22456
rect 5858 22422 5892 22450
rect 5858 22382 5892 22384
rect 5858 22350 5892 22382
rect 5858 22280 5892 22311
rect 5858 22277 5892 22280
rect 5858 22212 5892 22238
rect 5858 22204 5892 22212
rect 5858 22144 5892 22165
rect 5858 22131 5892 22144
rect 5858 22076 5892 22092
rect 5858 22058 5892 22076
rect 5858 22008 5892 22019
rect 5858 21985 5892 22008
rect 7340 22000 7363 22034
rect 7363 22000 7374 22034
rect 7412 22000 7431 22034
rect 7431 22000 7446 22034
rect 7572 22000 7587 22034
rect 7587 22000 7606 22034
rect 7644 22000 7655 22034
rect 7655 22000 7678 22034
rect 5858 21940 5892 21946
rect 5858 21912 5892 21940
rect 5858 21872 5892 21873
rect 5858 21839 5892 21872
rect 5858 21770 5892 21800
rect 5858 21766 5892 21770
rect 5858 21702 5892 21727
rect 5858 21693 5892 21702
rect 5858 21634 5892 21654
rect 5858 21620 5892 21634
rect 5858 21566 5892 21581
rect 5858 21547 5892 21566
rect 5858 21498 5892 21508
rect 5858 21474 5892 21498
rect 7342 21485 7376 21519
rect 7417 21485 7420 21519
rect 7420 21485 7451 21519
rect 7492 21485 7522 21519
rect 7522 21485 7526 21519
rect 7567 21485 7590 21519
rect 7590 21485 7601 21519
rect 7642 21485 7658 21519
rect 7658 21485 7676 21519
rect 5858 21430 5892 21435
rect 5858 21401 5892 21430
rect 5858 21328 5892 21362
rect 5858 21260 5892 21289
rect 5858 21255 5892 21260
rect 5858 21192 5892 21216
rect 5858 21182 5892 21192
rect 5858 21124 5892 21143
rect 5858 21109 5892 21124
rect 5858 21056 5892 21070
rect 5858 21036 5892 21056
rect 5858 20988 5892 20997
rect 5858 20963 5892 20988
rect 5858 20920 5892 20924
rect 5858 20890 5892 20920
rect 5858 20818 5892 20851
rect 5858 20817 5892 20818
rect 5858 20750 5892 20778
rect 5858 20744 5892 20750
rect 5858 20682 5892 20705
rect 5858 20671 5892 20682
rect 5858 20614 5892 20632
rect 5858 20598 5892 20614
rect 5858 20546 5892 20559
rect 5858 20525 5892 20546
rect 5858 20478 5892 20486
rect 5858 20452 5892 20478
rect 5858 20410 5892 20413
rect 5858 20379 5892 20410
rect 5858 20308 5892 20340
rect 5858 20306 5892 20308
rect 5858 20240 5892 20267
rect 5858 20233 5892 20240
rect 5858 20172 5892 20194
rect 5858 20160 5892 20172
rect 5858 20104 5892 20121
rect 5858 20087 5892 20104
rect 5858 20036 5892 20048
rect 5858 20014 5892 20036
rect 5858 19968 5892 19975
rect 5858 19941 5892 19968
rect 5858 19900 5892 19902
rect 5858 19868 5892 19900
rect 5858 19798 5892 19829
rect 5858 19795 5892 19798
rect 5858 19730 5892 19756
rect 5858 19722 5892 19730
rect 4899 19711 4933 19712
rect 4899 19640 4933 19672
rect 4899 19638 4933 19640
rect 4460 19570 4494 19596
rect 4460 19562 4494 19570
rect 4642 19591 4676 19625
rect 4726 19591 4760 19625
rect 4809 19591 4843 19625
rect 4460 19502 4494 19524
rect 4460 19490 4494 19502
rect 4899 19568 4933 19599
rect 5086 19666 5120 19700
rect 5086 19604 5102 19628
rect 5102 19604 5120 19628
rect 5362 19666 5396 19700
rect 5362 19604 5392 19628
rect 5392 19604 5396 19628
rect 5858 19662 5892 19683
rect 5858 19649 5892 19662
rect 5086 19594 5120 19604
rect 5362 19594 5396 19604
rect 4899 19565 4933 19568
rect 4899 19496 4933 19526
rect 4899 19492 4933 19496
rect 5858 19594 5892 19610
rect 5858 19576 5892 19594
rect 5858 19526 5892 19537
rect 5858 19503 5892 19526
rect 4460 19434 4494 19452
rect 4460 19418 4494 19434
rect 4585 19435 4619 19469
rect 4660 19435 4694 19469
rect 4735 19435 4769 19469
rect 4809 19435 4843 19469
rect 4460 19366 4494 19380
rect 4460 19346 4494 19366
rect 4460 19298 4494 19308
rect 4460 19274 4494 19298
rect 4460 19230 4494 19236
rect 4460 19202 4494 19230
rect 4460 19162 4494 19164
rect 4460 19130 4494 19162
rect 4460 19060 4494 19092
rect 4460 19058 4494 19060
rect 5858 19458 5892 19464
rect 5858 19430 5892 19458
rect 5858 19390 5892 19391
rect 5858 19357 5892 19390
rect 5858 19288 5892 19318
rect 5858 19284 5892 19288
rect 5858 19220 5892 19245
rect 5858 19211 5892 19220
rect 5858 19152 5892 19172
rect 5858 19138 5892 19152
rect 5080 19034 5092 19068
rect 5092 19034 5114 19068
rect 5152 19034 5186 19068
rect 5858 19084 5892 19099
rect 5858 19065 5892 19084
rect 4460 18992 4494 19020
rect 4460 18986 4494 18992
rect 4460 18924 4494 18948
rect 4460 18914 4494 18924
rect 4460 18856 4494 18876
rect 4460 18842 4494 18856
rect 4460 18788 4494 18804
rect 4460 18770 4494 18788
rect 4460 18720 4494 18732
rect 4460 18698 4494 18720
rect 4460 18652 4494 18660
rect 4460 18626 4494 18652
rect 4460 18584 4494 18588
rect 4460 18554 4494 18584
rect 5858 19016 5892 19026
rect 5858 18992 5892 19016
rect 5858 18948 5892 18953
rect 5858 18919 5892 18948
rect 5858 18846 5892 18880
rect 5858 18778 5892 18807
rect 5858 18773 5892 18778
rect 5858 18710 5892 18734
rect 5858 18700 5892 18710
rect 5858 18642 5892 18661
rect 5858 18627 5892 18642
rect 5858 18574 5892 18588
rect 5858 18554 5892 18574
rect 4532 18482 4566 18516
rect 4606 18482 4634 18516
rect 4634 18482 4640 18516
rect 4680 18482 4702 18516
rect 4702 18482 4714 18516
rect 4754 18482 4770 18516
rect 4770 18482 4788 18516
rect 4828 18482 4838 18516
rect 4838 18482 4862 18516
rect 4902 18482 4906 18516
rect 4906 18482 4936 18516
rect 4976 18482 5008 18516
rect 5008 18482 5010 18516
rect 5050 18482 5076 18516
rect 5076 18482 5084 18516
rect 5124 18482 5144 18516
rect 5144 18482 5158 18516
rect 5198 18482 5212 18516
rect 5212 18482 5232 18516
rect 5272 18482 5280 18516
rect 5280 18482 5306 18516
rect 5346 18482 5348 18516
rect 5348 18482 5380 18516
rect 5420 18482 5450 18516
rect 5450 18482 5454 18516
rect 5493 18482 5518 18516
rect 5518 18482 5527 18516
rect 5566 18482 5586 18516
rect 5586 18482 5600 18516
rect 5639 18482 5654 18516
rect 5654 18482 5673 18516
rect 5712 18482 5722 18516
rect 5722 18482 5746 18516
rect 5785 18482 5790 18516
rect 5790 18482 5819 18516
rect 2899 18255 2924 18289
rect 2924 18255 2933 18289
rect 2977 18255 2992 18289
rect 2992 18255 3011 18289
rect 3055 18255 3060 18289
rect 3060 18255 3089 18289
rect 3133 18255 3162 18289
rect 3162 18255 3167 18289
rect 3211 18255 3230 18289
rect 3230 18255 3245 18289
rect 3289 18255 3298 18289
rect 3298 18255 3323 18289
rect 3367 18255 3400 18289
rect 3400 18255 3401 18289
rect 3445 18255 3468 18289
rect 3468 18255 3479 18289
rect 3523 18255 3536 18289
rect 3536 18255 3557 18289
rect 3601 18255 3604 18289
rect 3604 18255 3635 18289
rect 3679 18255 3706 18289
rect 3706 18255 3713 18289
rect 3789 18255 3808 18289
rect 3808 18255 3823 18289
rect 3861 18255 3876 18289
rect 3876 18255 3895 18289
rect 3933 18255 3944 18289
rect 3944 18255 3967 18289
rect 4005 18255 4012 18289
rect 4012 18255 4039 18289
rect 4077 18255 4080 18289
rect 4080 18255 4111 18289
rect 4149 18255 4182 18289
rect 4182 18255 4183 18289
rect 4221 18255 4250 18289
rect 4250 18255 4255 18289
rect 4293 18255 4318 18289
rect 4318 18255 4327 18289
rect 4365 18255 4386 18289
rect 4386 18255 4399 18289
rect 4437 18255 4454 18289
rect 4454 18255 4471 18289
rect 4509 18255 4522 18289
rect 4522 18255 4543 18289
rect 4581 18255 4590 18289
rect 4590 18255 4615 18289
rect 4653 18255 4658 18289
rect 4658 18255 4687 18289
rect 4725 18255 4726 18289
rect 4726 18255 4759 18289
rect 4797 18255 4828 18289
rect 4828 18255 4831 18289
rect 4869 18255 4896 18289
rect 4896 18255 4903 18289
rect 4941 18255 4964 18289
rect 4964 18255 4975 18289
rect 5013 18255 5032 18289
rect 5032 18255 5047 18289
rect 5085 18255 5100 18289
rect 5100 18255 5119 18289
rect 5157 18255 5168 18289
rect 5168 18255 5191 18289
rect 5229 18255 5236 18289
rect 5236 18255 5263 18289
rect 5301 18255 5304 18289
rect 5304 18255 5335 18289
rect 5373 18255 5406 18289
rect 5406 18255 5407 18289
rect 5445 18255 5474 18289
rect 5474 18255 5479 18289
rect 5517 18255 5542 18289
rect 5542 18255 5551 18289
rect 5589 18255 5610 18289
rect 5610 18255 5623 18289
rect 5661 18255 5678 18289
rect 5678 18255 5695 18289
rect 5733 18255 5746 18289
rect 5746 18255 5767 18289
rect 5805 18255 5814 18289
rect 5814 18255 5839 18289
rect 5877 18255 5882 18289
rect 5882 18255 5911 18289
rect 5949 18255 5950 18289
rect 5950 18255 5983 18289
rect 6021 18255 6052 18289
rect 6052 18255 6055 18289
rect 6094 18255 6120 18289
rect 6120 18255 6128 18289
rect 6167 18255 6188 18289
rect 6188 18255 6201 18289
rect 6240 18255 6256 18289
rect 6256 18255 6274 18289
rect 6313 18255 6324 18289
rect 6324 18255 6347 18289
rect 6386 18255 6392 18289
rect 6392 18255 6420 18289
rect 6459 18255 6460 18289
rect 6460 18255 6493 18289
rect 6532 18255 6562 18289
rect 6562 18255 6566 18289
rect 6605 18255 6630 18289
rect 6630 18255 6639 18289
rect 6678 18255 6712 18289
rect 2822 18197 2856 18217
rect 2822 18183 2856 18197
rect 2822 18109 2856 18143
rect 2822 18049 2856 18069
rect 2822 18035 2856 18049
rect 6750 18187 6784 18216
rect 6750 18182 6784 18187
rect 6750 18119 6784 18143
rect 6750 18109 6784 18119
rect 6750 18051 6784 18070
rect 6750 18036 6784 18051
rect 2822 17981 2856 17995
rect 2822 17961 2856 17981
rect 2822 17913 2856 17921
rect 2822 17887 2856 17913
rect 2822 17845 2856 17847
rect 2822 17813 2856 17845
rect 2822 17743 2856 17774
rect 2822 17740 2856 17743
rect 2822 17675 2856 17701
rect 2822 17667 2856 17675
rect 2822 17607 2856 17628
rect 2822 17594 2856 17607
rect 2822 17539 2856 17555
rect 2822 17521 2856 17539
rect 2822 17471 2856 17482
rect 2822 17448 2856 17471
rect 2822 17403 2856 17409
rect 2822 17375 2856 17403
rect 2822 17335 2856 17336
rect 2822 17302 2856 17335
rect 2822 17233 2856 17263
rect 2822 17229 2856 17233
rect 2822 17165 2856 17190
rect 2822 17156 2856 17165
rect 2822 17097 2856 17117
rect 2822 17083 2856 17097
rect 2822 17029 2856 17044
rect 2822 17010 2856 17029
rect 2822 16961 2856 16971
rect 2822 16937 2856 16961
rect 2822 16893 2856 16898
rect 2822 16864 2856 16893
rect 2822 16791 2856 16825
rect 2822 16723 2856 16752
rect 2822 16718 2856 16723
rect 2822 16655 2856 16679
rect 2822 16645 2856 16655
rect 2822 16587 2856 16606
rect 2822 16572 2856 16587
rect 2822 16519 2856 16533
rect 2822 16499 2856 16519
rect 2822 16451 2856 16460
rect 2822 16426 2856 16451
rect 2822 16383 2856 16387
rect 2822 16353 2856 16383
rect 2822 16281 2856 16314
rect 2822 16280 2856 16281
rect 2822 16213 2856 16241
rect 2822 16207 2856 16213
rect 2822 16145 2856 16168
rect 2822 16134 2856 16145
rect 2822 16077 2856 16095
rect 2822 16061 2856 16077
rect 2822 16009 2856 16022
rect 2822 15988 2856 16009
rect 2822 15941 2856 15949
rect 2822 15915 2856 15941
rect 2822 15873 2856 15876
rect 2822 15842 2856 15873
rect 2822 15771 2856 15803
rect 2822 15769 2856 15771
rect 2822 15703 2856 15730
rect 2822 15696 2856 15703
rect 2822 15635 2856 15657
rect 2822 15623 2856 15635
rect 2822 15567 2856 15584
rect 2822 15550 2856 15567
rect 2822 15499 2856 15511
rect 2822 15477 2856 15499
rect 2822 15431 2856 15438
rect 2822 15404 2856 15431
rect 2822 15363 2856 15365
rect 2822 15331 2856 15363
rect 2822 15261 2856 15292
rect 2822 15258 2856 15261
rect 2822 15193 2856 15219
rect 2822 15185 2856 15193
rect 2822 15125 2856 15146
rect 2822 15112 2856 15125
rect 2822 15057 2856 15073
rect 2822 15039 2856 15057
rect 2822 14989 2856 15000
rect 2822 14966 2856 14989
rect 2822 14921 2856 14927
rect 2822 14893 2856 14921
rect 2822 14853 2856 14854
rect 2822 14820 2856 14853
rect 2822 14751 2856 14781
rect 2822 14747 2856 14751
rect 2822 14683 2856 14708
rect 2822 14674 2856 14683
rect 2822 14615 2856 14635
rect 2822 14601 2856 14615
rect 3161 17995 3184 18029
rect 3184 17995 3195 18029
rect 3240 17995 3252 18029
rect 3252 17995 3274 18029
rect 3319 17995 3320 18029
rect 3320 17995 3353 18029
rect 3398 17995 3422 18029
rect 3422 17995 3432 18029
rect 3478 17995 3490 18029
rect 3490 17995 3512 18029
rect 3558 17995 3592 18029
rect 3638 17995 3660 18029
rect 3660 17995 3672 18029
rect 3718 17995 3728 18029
rect 3728 17995 3752 18029
rect 3798 17995 3830 18029
rect 3830 17995 3832 18029
rect 3908 17995 3932 18029
rect 3932 17995 3942 18029
rect 3981 17995 4000 18029
rect 4000 17995 4015 18029
rect 4054 17995 4068 18029
rect 4068 17995 4088 18029
rect 4127 17995 4136 18029
rect 4136 17995 4161 18029
rect 4200 17995 4204 18029
rect 4204 17995 4234 18029
rect 4273 17995 4306 18029
rect 4306 17995 4307 18029
rect 4346 17995 4374 18029
rect 4374 17995 4380 18029
rect 4419 17995 4442 18029
rect 4442 17995 4453 18029
rect 4492 17995 4510 18029
rect 4510 17995 4526 18029
rect 4565 17995 4578 18029
rect 4578 17995 4599 18029
rect 4638 17995 4646 18029
rect 4646 17995 4672 18029
rect 4711 17995 4714 18029
rect 4714 17995 4745 18029
rect 4784 17995 4816 18029
rect 4816 17995 4818 18029
rect 4857 17995 4884 18029
rect 4884 17995 4891 18029
rect 4930 17995 4952 18029
rect 4952 17995 4964 18029
rect 5003 17995 5020 18029
rect 5020 17995 5037 18029
rect 5076 17995 5088 18029
rect 5088 17995 5110 18029
rect 5149 17995 5156 18029
rect 5156 17995 5183 18029
rect 5222 17995 5224 18029
rect 5224 17995 5256 18029
rect 5295 17995 5326 18029
rect 5326 17995 5329 18029
rect 5368 17995 5394 18029
rect 5394 17995 5402 18029
rect 5442 17995 5462 18029
rect 5462 17995 5476 18029
rect 5516 17995 5530 18029
rect 5530 17995 5550 18029
rect 5590 17995 5598 18029
rect 5598 17995 5624 18029
rect 5664 17995 5666 18029
rect 5666 17995 5698 18029
rect 5738 17995 5768 18029
rect 5768 17995 5772 18029
rect 5812 17995 5836 18029
rect 5836 17995 5846 18029
rect 5886 17995 5904 18029
rect 5904 17995 5920 18029
rect 5960 17995 5972 18029
rect 5972 17995 5994 18029
rect 6034 17995 6040 18029
rect 6040 17995 6068 18029
rect 6108 17995 6142 18029
rect 6182 17995 6210 18029
rect 6210 17995 6216 18029
rect 6256 17995 6278 18029
rect 6278 17995 6290 18029
rect 6330 17995 6346 18029
rect 6346 17995 6364 18029
rect 6404 17995 6438 18029
rect 3082 17935 3116 17957
rect 3082 17923 3116 17935
rect 3082 17867 3116 17884
rect 3082 17850 3116 17867
rect 3082 17799 3116 17811
rect 3082 17777 3116 17799
rect 6476 17927 6510 17957
rect 6476 17923 6510 17927
rect 6476 17859 6510 17885
rect 6476 17851 6510 17859
rect 6476 17791 6510 17813
rect 6476 17779 6510 17791
rect 3082 17731 3116 17738
rect 3082 17704 3116 17731
rect 3654 17711 3688 17745
rect 3745 17711 3779 17745
rect 3836 17711 3870 17745
rect 6476 17723 6510 17741
rect 6476 17707 6510 17723
rect 3082 17663 3116 17665
rect 3082 17631 3116 17663
rect 3552 17650 3586 17670
rect 3552 17636 3586 17650
rect 3082 17561 3116 17592
rect 3082 17558 3116 17561
rect 3082 17493 3116 17519
rect 3082 17485 3116 17493
rect 3082 17425 3116 17446
rect 3082 17412 3116 17425
rect 3082 17357 3116 17373
rect 3082 17339 3116 17357
rect 3082 17289 3116 17300
rect 3082 17266 3116 17289
rect 3082 17221 3116 17227
rect 3082 17193 3116 17221
rect 3082 17153 3116 17154
rect 3082 17120 3116 17153
rect 3082 17051 3116 17081
rect 3082 17047 3116 17051
rect 3082 16983 3116 17008
rect 3082 16974 3116 16983
rect 3082 16915 3116 16935
rect 3082 16901 3116 16915
rect 3082 16847 3116 16862
rect 3082 16828 3116 16847
rect 3082 16779 3116 16789
rect 3082 16755 3116 16779
rect 3082 16711 3116 16716
rect 3082 16682 3116 16711
rect 3082 16609 3116 16643
rect 3082 16541 3116 16570
rect 3082 16536 3116 16541
rect 3082 16473 3116 16497
rect 3082 16463 3116 16473
rect 3082 16405 3116 16424
rect 3082 16390 3116 16405
rect 3082 16337 3116 16351
rect 3082 16317 3116 16337
rect 3082 16269 3116 16278
rect 3082 16244 3116 16269
rect 3082 16201 3116 16205
rect 3082 16171 3116 16201
rect 3082 16099 3116 16132
rect 3082 16098 3116 16099
rect 3082 16031 3116 16059
rect 3082 16025 3116 16031
rect 3444 17599 3478 17603
rect 3444 17569 3478 17599
rect 3444 17496 3478 17529
rect 3444 17495 3478 17496
rect 3444 17427 3478 17455
rect 3444 17421 3478 17427
rect 3444 17358 3478 17381
rect 3444 17347 3478 17358
rect 3444 17289 3478 17306
rect 3444 17272 3478 17289
rect 3444 17220 3478 17231
rect 3444 17197 3478 17220
rect 3444 17151 3478 17156
rect 3444 17122 3478 17151
rect 6476 17655 6510 17668
rect 6476 17634 6510 17655
rect 3552 17579 3586 17589
rect 3552 17555 3586 17579
rect 3654 17555 3688 17589
rect 3728 17555 3762 17589
rect 6476 17587 6510 17595
rect 6476 17561 6510 17587
rect 3552 17474 3586 17508
rect 6476 17519 6510 17522
rect 6476 17488 6510 17519
rect 3552 17398 3586 17427
rect 3712 17399 3746 17433
rect 3786 17399 3820 17433
rect 3552 17393 3586 17398
rect 3552 17326 3586 17345
rect 3552 17311 3586 17326
rect 6476 17417 6510 17449
rect 6476 17415 6510 17417
rect 6476 17349 6510 17376
rect 6476 17342 6510 17349
rect 3552 17254 3586 17263
rect 3552 17229 3586 17254
rect 3654 17243 3688 17277
rect 3728 17243 3762 17277
rect 6476 17281 6510 17303
rect 6476 17269 6510 17281
rect 3552 17148 3586 17181
rect 3552 17147 3586 17148
rect 6476 17213 6510 17230
rect 6476 17196 6510 17213
rect 3654 17087 3688 17121
rect 3745 17087 3779 17121
rect 3836 17087 3870 17121
rect 6476 17145 6510 17157
rect 6476 17123 6510 17145
rect 3444 17047 3478 17081
rect 3444 16975 3478 17006
rect 6476 17077 6510 17084
rect 6476 17050 6510 17077
rect 3444 16972 3478 16975
rect 3444 16905 3478 16931
rect 3444 16897 3478 16905
rect 6237 16962 6271 16964
rect 6237 16930 6245 16962
rect 6245 16930 6271 16962
rect 6309 16962 6343 16964
rect 6309 16930 6337 16962
rect 6337 16930 6343 16962
rect 3444 16835 3478 16856
rect 3444 16822 3478 16835
rect 4314 16833 4319 16867
rect 4319 16833 4348 16867
rect 4387 16833 4391 16867
rect 4391 16833 4421 16867
rect 4460 16833 4463 16867
rect 4463 16833 4494 16867
rect 4533 16833 4535 16867
rect 4535 16833 4567 16867
rect 4606 16833 4607 16867
rect 4607 16833 4640 16867
rect 4679 16833 4713 16867
rect 4752 16833 4786 16867
rect 4958 16833 4981 16867
rect 4981 16833 4992 16867
rect 5041 16833 5053 16867
rect 5053 16833 5075 16867
rect 5124 16833 5125 16867
rect 5125 16833 5158 16867
rect 5207 16833 5231 16867
rect 5231 16833 5241 16867
rect 5289 16833 5303 16867
rect 5303 16833 5323 16867
rect 5371 16833 5374 16867
rect 5374 16833 5405 16867
rect 6237 16857 6271 16891
rect 6309 16857 6343 16891
rect 3444 16765 3478 16781
rect 3444 16747 3478 16765
rect 6237 16785 6245 16818
rect 6245 16785 6271 16818
rect 6237 16784 6271 16785
rect 6309 16785 6337 16818
rect 6337 16785 6343 16818
rect 6309 16784 6343 16785
rect 3444 16695 3478 16706
rect 3444 16672 3478 16695
rect 3444 16625 3478 16631
rect 3444 16597 3478 16625
rect 3444 16555 3478 16556
rect 3444 16522 3478 16555
rect 3444 16451 3478 16481
rect 3444 16447 3478 16451
rect 3444 16381 3478 16406
rect 3444 16372 3478 16381
rect 3444 16311 3478 16331
rect 3444 16297 3478 16311
rect 3444 16241 3478 16256
rect 3444 16222 3478 16241
rect 3444 16171 3478 16181
rect 3444 16147 3478 16171
rect 3444 16101 3478 16106
rect 3444 16072 3478 16101
rect 3721 16709 3827 16711
rect 3721 16675 3729 16709
rect 3729 16675 3821 16709
rect 3821 16675 3827 16709
rect 3721 16564 3827 16675
rect 3721 16530 3729 16564
rect 3729 16530 3821 16564
rect 3821 16530 3827 16564
rect 3721 16419 3827 16530
rect 3721 16385 3729 16419
rect 3729 16385 3821 16419
rect 3821 16385 3827 16419
rect 3721 16274 3827 16385
rect 3721 16240 3729 16274
rect 3729 16240 3821 16274
rect 3821 16240 3827 16274
rect 3721 16129 3827 16240
rect 3721 16101 3729 16129
rect 3729 16101 3821 16129
rect 3821 16101 3827 16129
rect 6237 16711 6271 16745
rect 6309 16711 6343 16745
rect 6237 16642 6245 16672
rect 6245 16642 6271 16672
rect 6237 16638 6271 16642
rect 6309 16642 6337 16672
rect 6337 16642 6343 16672
rect 6309 16638 6343 16642
rect 6237 16565 6271 16599
rect 6309 16565 6343 16599
rect 6237 16499 6245 16525
rect 6245 16499 6271 16525
rect 6237 16491 6271 16499
rect 6309 16499 6337 16525
rect 6337 16499 6343 16525
rect 6309 16491 6343 16499
rect 6237 16417 6271 16451
rect 6309 16417 6343 16451
rect 6237 16356 6245 16377
rect 6245 16356 6271 16377
rect 6237 16343 6271 16356
rect 6309 16356 6337 16377
rect 6337 16356 6343 16377
rect 6309 16343 6343 16356
rect 6237 16269 6271 16303
rect 6309 16269 6343 16303
rect 6237 16213 6245 16229
rect 6245 16213 6271 16229
rect 6237 16195 6271 16213
rect 6309 16213 6337 16229
rect 6337 16213 6343 16229
rect 6309 16195 6343 16213
rect 6237 16121 6271 16155
rect 6309 16121 6343 16155
rect 3721 16028 3755 16062
rect 3793 16028 3827 16062
rect 4282 16061 4285 16095
rect 4285 16061 4316 16095
rect 4355 16061 4389 16095
rect 4428 16061 4458 16095
rect 4458 16061 4462 16095
rect 4501 16061 4527 16095
rect 4527 16061 4535 16095
rect 4574 16061 4596 16095
rect 4596 16061 4608 16095
rect 4647 16061 4665 16095
rect 4665 16061 4681 16095
rect 4720 16061 4735 16095
rect 4735 16061 4754 16095
rect 4793 16061 4805 16095
rect 4805 16061 4827 16095
rect 4866 16061 4875 16095
rect 4875 16061 4900 16095
rect 4939 16061 4945 16095
rect 4945 16061 4973 16095
rect 5012 16061 5015 16095
rect 5015 16061 5046 16095
rect 5085 16061 5119 16095
rect 5158 16061 5189 16095
rect 5189 16061 5192 16095
rect 5231 16061 5259 16095
rect 5259 16061 5265 16095
rect 5304 16061 5329 16095
rect 5329 16061 5338 16095
rect 5377 16061 5399 16095
rect 5399 16061 5411 16095
rect 5450 16061 5469 16095
rect 5469 16061 5484 16095
rect 5523 16061 5539 16095
rect 5539 16061 5557 16095
rect 5596 16061 5609 16095
rect 5609 16061 5630 16095
rect 5669 16061 5679 16095
rect 5679 16061 5703 16095
rect 5742 16061 5749 16095
rect 5749 16061 5776 16095
rect 6237 16070 6245 16081
rect 6245 16070 6271 16081
rect 3082 15963 3116 15986
rect 3082 15952 3116 15963
rect 3082 15895 3116 15913
rect 3082 15879 3116 15895
rect 3082 15827 3116 15840
rect 3082 15806 3116 15827
rect 3082 15759 3116 15767
rect 3082 15733 3116 15759
rect 3082 15691 3116 15694
rect 3082 15660 3116 15691
rect 3082 15589 3116 15621
rect 3082 15587 3116 15589
rect 3082 15521 3116 15548
rect 3082 15514 3116 15521
rect 3082 15453 3116 15475
rect 3082 15441 3116 15453
rect 3082 15385 3116 15402
rect 3082 15368 3116 15385
rect 3082 15317 3116 15329
rect 3082 15295 3116 15317
rect 3082 15249 3116 15256
rect 3082 15222 3116 15249
rect 3082 15181 3116 15183
rect 3082 15149 3116 15181
rect 3082 15079 3116 15110
rect 3082 15076 3116 15079
rect 3082 15011 3116 15037
rect 3082 15003 3116 15011
rect 3082 14943 3116 14964
rect 3082 14930 3116 14943
rect 3082 14875 3116 14891
rect 3082 14857 3116 14875
rect 3082 14807 3116 14819
rect 3082 14785 3116 14807
rect 3082 14739 3116 14747
rect 3082 14713 3116 14739
rect 3082 14671 3116 14675
rect 3082 14641 3116 14671
rect 3721 15984 3755 15989
rect 3721 15955 3729 15984
rect 3729 15955 3755 15984
rect 3793 15984 3827 15989
rect 3793 15955 3821 15984
rect 3821 15955 3827 15984
rect 3721 15882 3755 15916
rect 3793 15882 3827 15916
rect 3721 15839 3755 15843
rect 3721 15809 3729 15839
rect 3729 15809 3755 15839
rect 3793 15839 3827 15843
rect 3793 15809 3821 15839
rect 3821 15809 3827 15839
rect 3721 15736 3755 15770
rect 3793 15736 3827 15770
rect 3721 15693 3755 15697
rect 3721 15663 3729 15693
rect 3729 15663 3755 15693
rect 3793 15693 3827 15697
rect 3793 15663 3821 15693
rect 3821 15663 3827 15693
rect 3721 15590 3755 15624
rect 3793 15590 3827 15624
rect 3721 15547 3755 15551
rect 3721 15517 3729 15547
rect 3729 15517 3755 15547
rect 3793 15547 3827 15551
rect 3793 15517 3821 15547
rect 3821 15517 3827 15547
rect 3721 15444 3755 15478
rect 3793 15444 3827 15478
rect 3721 15401 3755 15405
rect 3721 15371 3729 15401
rect 3729 15371 3755 15401
rect 3793 15401 3827 15405
rect 3793 15371 3821 15401
rect 3821 15371 3827 15401
rect 6237 16047 6271 16070
rect 6309 16070 6337 16081
rect 6337 16070 6343 16081
rect 6309 16047 6343 16070
rect 6237 15973 6271 16007
rect 6309 15973 6343 16007
rect 6237 15927 6245 15933
rect 6245 15927 6271 15933
rect 6237 15899 6271 15927
rect 6309 15927 6337 15933
rect 6337 15927 6343 15933
rect 6309 15899 6343 15927
rect 6237 15825 6271 15859
rect 6309 15825 6343 15859
rect 6237 15784 6245 15785
rect 6245 15784 6271 15785
rect 6237 15751 6271 15784
rect 6309 15784 6337 15785
rect 6337 15784 6343 15785
rect 6309 15751 6343 15784
rect 6237 15677 6271 15711
rect 6309 15677 6343 15711
rect 6237 15603 6271 15637
rect 6309 15603 6343 15637
rect 6237 15532 6271 15563
rect 6237 15529 6245 15532
rect 6245 15529 6271 15532
rect 6309 15532 6343 15563
rect 6309 15529 6337 15532
rect 6337 15529 6343 15532
rect 6237 15455 6271 15489
rect 6309 15455 6343 15489
rect 6237 15389 6271 15415
rect 6237 15381 6245 15389
rect 6245 15381 6271 15389
rect 6309 15389 6343 15415
rect 6309 15381 6337 15389
rect 6337 15381 6343 15389
rect 3721 15298 3755 15332
rect 3793 15298 3827 15332
rect 4282 15331 4285 15365
rect 4285 15331 4316 15365
rect 4355 15331 4389 15365
rect 4428 15331 4458 15365
rect 4458 15331 4462 15365
rect 4501 15331 4527 15365
rect 4527 15331 4535 15365
rect 4574 15331 4596 15365
rect 4596 15331 4608 15365
rect 4647 15331 4665 15365
rect 4665 15331 4681 15365
rect 4720 15331 4735 15365
rect 4735 15331 4754 15365
rect 4793 15331 4805 15365
rect 4805 15331 4827 15365
rect 4866 15331 4875 15365
rect 4875 15331 4900 15365
rect 4939 15331 4945 15365
rect 4945 15331 4973 15365
rect 5012 15331 5015 15365
rect 5015 15331 5046 15365
rect 5085 15331 5119 15365
rect 5158 15331 5189 15365
rect 5189 15331 5192 15365
rect 5231 15331 5259 15365
rect 5259 15331 5265 15365
rect 5304 15331 5329 15365
rect 5329 15331 5338 15365
rect 5377 15331 5399 15365
rect 5399 15331 5411 15365
rect 5450 15331 5469 15365
rect 5469 15331 5484 15365
rect 5523 15331 5539 15365
rect 5539 15331 5557 15365
rect 5596 15331 5609 15365
rect 5609 15331 5630 15365
rect 5669 15331 5679 15365
rect 5679 15331 5703 15365
rect 5742 15331 5749 15365
rect 5749 15331 5776 15365
rect 3721 15255 3755 15259
rect 3721 15225 3729 15255
rect 3729 15225 3755 15255
rect 3793 15255 3827 15259
rect 3793 15225 3821 15255
rect 3821 15225 3827 15255
rect 3721 15152 3755 15186
rect 3793 15152 3827 15186
rect 3721 15109 3755 15113
rect 3721 15079 3729 15109
rect 3729 15079 3755 15109
rect 3793 15109 3827 15113
rect 3793 15079 3821 15109
rect 3821 15079 3827 15109
rect 3721 15006 3755 15040
rect 3793 15006 3827 15040
rect 3721 14963 3755 14967
rect 3721 14933 3729 14963
rect 3729 14933 3755 14963
rect 3793 14963 3827 14967
rect 3793 14933 3821 14963
rect 3821 14933 3827 14963
rect 3721 14860 3755 14894
rect 3793 14860 3827 14894
rect 3721 14817 3755 14821
rect 3721 14787 3729 14817
rect 3729 14787 3755 14817
rect 3793 14817 3827 14821
rect 3793 14787 3821 14817
rect 3821 14787 3827 14817
rect 3721 14714 3755 14748
rect 3793 14714 3827 14748
rect 3721 14671 3755 14675
rect 3721 14641 3729 14671
rect 3729 14641 3755 14671
rect 3793 14671 3827 14675
rect 3793 14641 3821 14671
rect 3821 14641 3827 14671
rect 6237 15307 6271 15341
rect 6309 15307 6343 15341
rect 6237 15246 6271 15267
rect 6237 15233 6245 15246
rect 6245 15233 6271 15246
rect 6309 15246 6343 15267
rect 6309 15233 6337 15246
rect 6337 15233 6343 15246
rect 6237 15159 6271 15193
rect 6309 15159 6343 15193
rect 6237 15103 6271 15119
rect 6237 15085 6245 15103
rect 6245 15085 6271 15103
rect 6309 15103 6343 15119
rect 6309 15085 6337 15103
rect 6337 15085 6343 15103
rect 6237 15011 6271 15045
rect 6309 15011 6343 15045
rect 6237 14959 6271 14971
rect 6237 14937 6245 14959
rect 6245 14937 6271 14959
rect 6309 14959 6343 14971
rect 6309 14937 6337 14959
rect 6337 14937 6343 14959
rect 6237 14863 6271 14897
rect 6309 14863 6343 14897
rect 6237 14815 6271 14823
rect 6237 14789 6245 14815
rect 6245 14789 6271 14815
rect 6309 14815 6343 14823
rect 6309 14789 6337 14815
rect 6337 14789 6343 14815
rect 6237 14715 6271 14749
rect 6309 14715 6343 14749
rect 6237 14671 6343 14675
rect 6237 14637 6245 14671
rect 6245 14637 6337 14671
rect 6337 14637 6343 14671
rect 6237 14603 6343 14637
rect 6476 17009 6510 17011
rect 6476 16977 6510 17009
rect 6476 16907 6510 16938
rect 6476 16904 6510 16907
rect 6476 16839 6510 16865
rect 6476 16831 6510 16839
rect 6476 16771 6510 16792
rect 6476 16758 6510 16771
rect 6476 16703 6510 16719
rect 6476 16685 6510 16703
rect 6476 16635 6510 16646
rect 6476 16612 6510 16635
rect 6476 16567 6510 16573
rect 6476 16539 6510 16567
rect 6476 16499 6510 16500
rect 6476 16466 6510 16499
rect 6476 16397 6510 16427
rect 6476 16393 6510 16397
rect 6476 16329 6510 16354
rect 6476 16320 6510 16329
rect 6476 16261 6510 16281
rect 6476 16247 6510 16261
rect 6476 16193 6510 16208
rect 6476 16174 6510 16193
rect 6476 16125 6510 16135
rect 6476 16101 6510 16125
rect 6476 16057 6510 16062
rect 6476 16028 6510 16057
rect 6476 15955 6510 15989
rect 6476 15887 6510 15916
rect 6476 15882 6510 15887
rect 6476 15819 6510 15843
rect 6476 15809 6510 15819
rect 6476 15751 6510 15770
rect 6476 15736 6510 15751
rect 6476 15683 6510 15697
rect 6476 15663 6510 15683
rect 6476 15615 6510 15624
rect 6476 15590 6510 15615
rect 6476 15547 6510 15551
rect 6476 15517 6510 15547
rect 6476 15445 6510 15478
rect 6476 15444 6510 15445
rect 6476 15377 6510 15405
rect 6476 15371 6510 15377
rect 6476 15309 6510 15332
rect 6476 15298 6510 15309
rect 6476 15241 6510 15259
rect 6476 15225 6510 15241
rect 6476 15173 6510 15186
rect 6476 15152 6510 15173
rect 6476 15105 6510 15113
rect 6476 15079 6510 15105
rect 6476 15037 6510 15040
rect 6476 15006 6510 15037
rect 6476 14935 6510 14967
rect 6476 14933 6510 14935
rect 6476 14867 6510 14894
rect 6476 14860 6510 14867
rect 6476 14799 6510 14821
rect 6476 14787 6510 14799
rect 6476 14731 6510 14748
rect 6476 14714 6510 14731
rect 6476 14663 6510 14675
rect 6476 14641 6510 14663
rect 3154 14569 3188 14603
rect 3227 14569 3246 14603
rect 3246 14569 3261 14603
rect 3300 14569 3314 14603
rect 3314 14569 3334 14603
rect 3373 14569 3382 14603
rect 3382 14569 3407 14603
rect 3446 14569 3450 14603
rect 3450 14569 3480 14603
rect 3519 14569 3552 14603
rect 3552 14569 3553 14603
rect 3592 14569 3620 14603
rect 3620 14569 3626 14603
rect 3665 14569 3688 14603
rect 3688 14569 3699 14603
rect 3738 14569 3756 14603
rect 3756 14569 3772 14603
rect 3811 14569 3824 14603
rect 3824 14569 3845 14603
rect 3884 14569 3892 14603
rect 3892 14569 3918 14603
rect 3956 14569 3960 14603
rect 3960 14569 3990 14603
rect 4028 14569 4062 14603
rect 4100 14569 4130 14603
rect 4130 14569 4134 14603
rect 4172 14569 4198 14603
rect 4198 14569 4206 14603
rect 4244 14569 4266 14603
rect 4266 14569 4278 14603
rect 4316 14569 4334 14603
rect 4334 14569 4350 14603
rect 4388 14569 4402 14603
rect 4402 14569 4422 14603
rect 4460 14569 4470 14603
rect 4470 14569 4494 14603
rect 4532 14569 4538 14603
rect 4538 14569 4566 14603
rect 4604 14569 4606 14603
rect 4606 14569 4638 14603
rect 4676 14569 4708 14603
rect 4708 14569 4710 14603
rect 4748 14569 4776 14603
rect 4776 14569 4782 14603
rect 4820 14569 4844 14603
rect 4844 14569 4854 14603
rect 4892 14569 4912 14603
rect 4912 14569 4926 14603
rect 4964 14569 4980 14603
rect 4980 14569 4998 14603
rect 5036 14569 5048 14603
rect 5048 14569 5070 14603
rect 5108 14569 5116 14603
rect 5116 14569 5142 14603
rect 5180 14569 5184 14603
rect 5184 14569 5214 14603
rect 5252 14569 5286 14603
rect 5324 14569 5354 14603
rect 5354 14569 5358 14603
rect 5396 14569 5422 14603
rect 5422 14569 5430 14603
rect 5468 14569 5490 14603
rect 5490 14569 5502 14603
rect 5540 14569 5558 14603
rect 5558 14569 5574 14603
rect 5612 14569 5626 14603
rect 5626 14569 5646 14603
rect 5684 14569 5694 14603
rect 5694 14569 5718 14603
rect 5756 14569 5762 14603
rect 5762 14569 5790 14603
rect 5828 14569 5830 14603
rect 5830 14569 5862 14603
rect 5900 14569 5932 14603
rect 5932 14569 5934 14603
rect 5972 14569 6000 14603
rect 6000 14569 6006 14603
rect 6044 14569 6068 14603
rect 6068 14569 6078 14603
rect 6116 14569 6136 14603
rect 6136 14569 6150 14603
rect 6188 14569 6204 14603
rect 6204 14569 6222 14603
rect 6237 14569 6238 14603
rect 6238 14569 6272 14603
rect 6272 14569 6306 14603
rect 6306 14569 6340 14603
rect 6340 14569 6366 14603
rect 6404 14569 6408 14603
rect 6408 14569 6438 14603
rect 6750 17983 6784 17997
rect 6750 17963 6784 17983
rect 6750 17915 6784 17924
rect 6750 17890 6784 17915
rect 6750 17847 6784 17851
rect 6750 17817 6784 17847
rect 6750 17745 6784 17778
rect 6750 17744 6784 17745
rect 6750 17677 6784 17705
rect 6750 17671 6784 17677
rect 6750 17609 6784 17632
rect 6750 17598 6784 17609
rect 6750 17541 6784 17559
rect 6750 17525 6784 17541
rect 6750 17473 6784 17486
rect 6750 17452 6784 17473
rect 6750 17405 6784 17413
rect 6750 17379 6784 17405
rect 6750 17337 6784 17340
rect 6750 17306 6784 17337
rect 6750 17235 6784 17267
rect 6750 17233 6784 17235
rect 6750 17167 6784 17194
rect 6750 17160 6784 17167
rect 6750 17099 6784 17121
rect 6750 17087 6784 17099
rect 6750 17031 6784 17048
rect 6750 17014 6784 17031
rect 6750 16963 6784 16975
rect 6750 16941 6784 16963
rect 6750 16895 6784 16902
rect 6750 16868 6784 16895
rect 6750 16827 6784 16829
rect 6750 16795 6784 16827
rect 6750 16725 6784 16756
rect 6750 16722 6784 16725
rect 6750 16657 6784 16683
rect 6750 16649 6784 16657
rect 6750 16589 6784 16610
rect 6750 16576 6784 16589
rect 6750 16521 6784 16537
rect 6750 16503 6784 16521
rect 6750 16453 6784 16464
rect 6750 16430 6784 16453
rect 6750 16385 6784 16391
rect 6750 16357 6784 16385
rect 6750 16317 6784 16318
rect 6750 16284 6784 16317
rect 6750 16215 6784 16245
rect 6750 16211 6784 16215
rect 6750 16147 6784 16172
rect 6750 16138 6784 16147
rect 6750 16079 6784 16099
rect 6750 16065 6784 16079
rect 6750 16011 6784 16026
rect 6750 15992 6784 16011
rect 6750 15943 6784 15953
rect 6750 15919 6784 15943
rect 6750 15875 6784 15880
rect 6750 15846 6784 15875
rect 6750 15773 6784 15807
rect 6750 15705 6784 15734
rect 6750 15700 6784 15705
rect 6750 15637 6784 15661
rect 6750 15627 6784 15637
rect 6750 15569 6784 15588
rect 6750 15554 6784 15569
rect 6750 15501 6784 15515
rect 6750 15481 6784 15501
rect 6750 15433 6784 15442
rect 6750 15408 6784 15433
rect 6750 15365 6784 15369
rect 6750 15335 6784 15365
rect 6750 15263 6784 15296
rect 6750 15262 6784 15263
rect 6750 15195 6784 15223
rect 6750 15189 6784 15195
rect 6750 15127 6784 15150
rect 6750 15116 6784 15127
rect 6750 15059 6784 15077
rect 6750 15043 6784 15059
rect 6750 14991 6784 15004
rect 6750 14970 6784 14991
rect 6750 14923 6784 14931
rect 6750 14897 6784 14923
rect 6750 14855 6784 14858
rect 6750 14824 6784 14855
rect 6750 14753 6784 14785
rect 6750 14751 6784 14753
rect 6750 14685 6784 14711
rect 6750 14677 6784 14685
rect 6750 14617 6784 14637
rect 6750 14603 6784 14617
rect 2822 14547 2856 14562
rect 2822 14528 2856 14547
rect 2822 14479 2856 14489
rect 2822 14455 2856 14479
rect 2822 14411 2856 14416
rect 2822 14382 2856 14411
rect 6750 14549 6784 14563
rect 6750 14529 6784 14549
rect 6750 14481 6784 14489
rect 6750 14455 6784 14481
rect 6750 14413 6784 14415
rect 6750 14381 6784 14413
rect 2894 14309 2928 14343
rect 2967 14309 2976 14343
rect 2976 14309 3001 14343
rect 3040 14309 3044 14343
rect 3044 14309 3074 14343
rect 3113 14309 3146 14343
rect 3146 14309 3147 14343
rect 3186 14309 3214 14343
rect 3214 14309 3220 14343
rect 3259 14309 3282 14343
rect 3282 14309 3293 14343
rect 3332 14309 3350 14343
rect 3350 14309 3366 14343
rect 3405 14309 3418 14343
rect 3418 14309 3439 14343
rect 3478 14309 3486 14343
rect 3486 14309 3512 14343
rect 3551 14309 3554 14343
rect 3554 14309 3585 14343
rect 3624 14309 3656 14343
rect 3656 14309 3658 14343
rect 3697 14309 3724 14343
rect 3724 14309 3731 14343
rect 3770 14309 3792 14343
rect 3792 14309 3804 14343
rect 3843 14309 3860 14343
rect 3860 14309 3877 14343
rect 3916 14309 3928 14343
rect 3928 14309 3950 14343
rect 3989 14309 3996 14343
rect 3996 14309 4023 14343
rect 4062 14309 4064 14343
rect 4064 14309 4096 14343
rect 4135 14309 4166 14343
rect 4166 14309 4169 14343
rect 4208 14309 4234 14343
rect 4234 14309 4242 14343
rect 4281 14309 4302 14343
rect 4302 14309 4315 14343
rect 4354 14309 4370 14343
rect 4370 14309 4388 14343
rect 4427 14309 4438 14343
rect 4438 14309 4461 14343
rect 4500 14309 4506 14343
rect 4506 14309 4534 14343
rect 4573 14309 4574 14343
rect 4574 14309 4607 14343
rect 4646 14309 4676 14343
rect 4676 14309 4680 14343
rect 4719 14309 4744 14343
rect 4744 14309 4753 14343
rect 4792 14309 4812 14343
rect 4812 14309 4826 14343
rect 4865 14309 4880 14343
rect 4880 14309 4899 14343
rect 4938 14309 4948 14343
rect 4948 14309 4972 14343
rect 5011 14309 5016 14343
rect 5016 14309 5045 14343
rect 5084 14309 5118 14343
rect 5157 14309 5186 14343
rect 5186 14309 5191 14343
rect 5230 14309 5254 14343
rect 5254 14309 5264 14343
rect 5303 14309 5322 14343
rect 5322 14309 5337 14343
rect 5376 14309 5390 14343
rect 5390 14309 5410 14343
rect 5449 14309 5458 14343
rect 5458 14309 5483 14343
rect 5522 14309 5526 14343
rect 5526 14309 5556 14343
rect 5595 14309 5628 14343
rect 5628 14309 5629 14343
rect 5668 14309 5696 14343
rect 5696 14309 5702 14343
rect 5741 14309 5764 14343
rect 5764 14309 5775 14343
rect 5814 14309 5832 14343
rect 5832 14309 5848 14343
rect 5886 14309 5900 14343
rect 5900 14309 5920 14343
rect 5958 14309 5968 14343
rect 5968 14309 5992 14343
rect 6030 14309 6036 14343
rect 6036 14309 6064 14343
rect 6102 14309 6104 14343
rect 6104 14309 6136 14343
rect 6174 14309 6206 14343
rect 6206 14309 6208 14343
rect 6246 14309 6274 14343
rect 6274 14309 6280 14343
rect 6318 14309 6342 14343
rect 6342 14309 6352 14343
rect 6390 14309 6410 14343
rect 6410 14309 6424 14343
rect 6462 14309 6478 14343
rect 6478 14309 6496 14343
rect 6534 14309 6546 14343
rect 6546 14309 6568 14343
rect 6606 14309 6614 14343
rect 6614 14309 6640 14343
rect 6678 14309 6682 14343
rect 6682 14309 6712 14343
<< metal1 >>
rect 2816 39874 7786 39880
rect 2816 39840 2897 39874
rect 2931 39840 2972 39874
rect 3006 39840 3047 39874
rect 3081 39840 3123 39874
rect 3157 39840 3199 39874
rect 3233 39840 3275 39874
rect 3309 39840 3351 39874
rect 3385 39840 3427 39874
rect 3461 39840 3503 39874
rect 3537 39840 3579 39874
rect 3613 39840 3655 39874
rect 3689 39840 3731 39874
rect 3765 39840 3807 39874
rect 3841 39840 3883 39874
rect 3917 39840 3959 39874
rect 3993 39840 4035 39874
rect 4069 39840 4111 39874
rect 4145 39840 4221 39874
rect 4255 39840 4294 39874
rect 4328 39840 4367 39874
rect 4401 39840 4440 39874
rect 4474 39840 4513 39874
rect 4547 39840 4586 39874
rect 4620 39840 4659 39874
rect 4693 39840 4732 39874
rect 4766 39840 4805 39874
rect 4839 39840 4878 39874
rect 4912 39840 4951 39874
rect 4985 39840 5024 39874
rect 5058 39840 5097 39874
rect 5131 39840 5170 39874
rect 5204 39840 5243 39874
rect 5277 39840 5316 39874
rect 5350 39840 5389 39874
rect 5423 39840 5462 39874
rect 5496 39840 5535 39874
rect 5569 39840 5608 39874
rect 5642 39840 5681 39874
rect 5715 39840 5754 39874
rect 5788 39840 5827 39874
rect 5861 39840 5900 39874
rect 5934 39840 5973 39874
rect 6007 39840 6046 39874
rect 6080 39840 6120 39874
rect 6154 39840 6194 39874
rect 6228 39840 6268 39874
rect 6302 39840 6342 39874
rect 6376 39840 6416 39874
rect 6450 39840 6490 39874
rect 6524 39840 6564 39874
rect 6598 39840 6638 39874
rect 6672 39840 6712 39874
rect 6746 39840 6786 39874
rect 6820 39840 6860 39874
rect 6894 39840 6934 39874
rect 6968 39840 7008 39874
rect 7042 39840 7082 39874
rect 7116 39840 7156 39874
rect 7190 39840 7230 39874
rect 7264 39840 7304 39874
rect 7338 39840 7378 39874
rect 7412 39840 7452 39874
rect 7486 39840 7526 39874
rect 7560 39840 7600 39874
rect 7634 39840 7674 39874
rect 7708 39840 7786 39874
rect 2816 39834 7786 39840
rect 2816 39802 2862 39834
rect 2816 39768 2822 39802
rect 2856 39768 2862 39802
rect 2816 39729 2862 39768
rect 2816 39695 2822 39729
rect 2856 39695 2862 39729
rect 2816 39656 2862 39695
rect 2816 39622 2822 39656
rect 2856 39622 2862 39656
rect 2816 39583 2862 39622
rect 7740 39802 7786 39834
rect 7740 39768 7746 39802
rect 7780 39768 7786 39802
rect 7740 39730 7786 39768
rect 7740 39696 7746 39730
rect 7780 39696 7786 39730
rect 7740 39658 7786 39696
rect 7740 39624 7746 39658
rect 7780 39624 7786 39658
rect 2816 39549 2822 39583
rect 2856 39549 2862 39583
rect 2816 39510 2862 39549
rect 2816 39476 2822 39510
rect 2856 39476 2862 39510
rect 2816 39437 2862 39476
rect 2816 39403 2822 39437
rect 2856 39403 2862 39437
rect 2816 39364 2862 39403
rect 2816 39330 2822 39364
rect 2856 39330 2862 39364
rect 2816 39291 2862 39330
rect 2816 39257 2822 39291
rect 2856 39257 2862 39291
rect 2816 39218 2862 39257
rect 2816 39184 2822 39218
rect 2856 39184 2862 39218
rect 2816 39145 2862 39184
rect 2816 39111 2822 39145
rect 2856 39111 2862 39145
rect 2816 39072 2862 39111
rect 2816 39038 2822 39072
rect 2856 39038 2862 39072
rect 2816 38999 2862 39038
rect 2816 38965 2822 38999
rect 2856 38965 2862 38999
rect 2816 38926 2862 38965
rect 2816 38892 2822 38926
rect 2856 38892 2862 38926
rect 2816 38853 2862 38892
rect 2816 38819 2822 38853
rect 2856 38819 2862 38853
rect 2816 38780 2862 38819
rect 2816 38746 2822 38780
rect 2856 38746 2862 38780
rect 2816 38707 2862 38746
rect 2816 38673 2822 38707
rect 2856 38673 2862 38707
rect 2816 38634 2862 38673
rect 2816 38600 2822 38634
rect 2856 38600 2862 38634
rect 2816 38561 2862 38600
rect 2816 38527 2822 38561
rect 2856 38527 2862 38561
rect 2816 38488 2862 38527
rect 2816 38454 2822 38488
rect 2856 38454 2862 38488
rect 2816 38415 2862 38454
rect 2816 38381 2822 38415
rect 2856 38381 2862 38415
rect 2816 38342 2862 38381
rect 2816 38308 2822 38342
rect 2856 38308 2862 38342
rect 2816 38269 2862 38308
rect 2816 38235 2822 38269
rect 2856 38235 2862 38269
rect 2816 38196 2862 38235
rect 2816 38162 2822 38196
rect 2856 38162 2862 38196
rect 2816 38123 2862 38162
rect 2816 38089 2822 38123
rect 2856 38089 2862 38123
rect 2816 38050 2862 38089
rect 2816 38016 2822 38050
rect 2856 38016 2862 38050
rect 2816 37977 2862 38016
rect 2816 37943 2822 37977
rect 2856 37943 2862 37977
rect 2816 37904 2862 37943
rect 2816 37870 2822 37904
rect 2856 37870 2862 37904
rect 2816 37831 2862 37870
rect 2816 37797 2822 37831
rect 2856 37797 2862 37831
rect 2816 37758 2862 37797
rect 2816 37724 2822 37758
rect 2856 37724 2862 37758
rect 2816 37685 2862 37724
rect 2816 37651 2822 37685
rect 2856 37651 2862 37685
rect 2816 37612 2862 37651
rect 2816 37578 2822 37612
rect 2856 37578 2862 37612
rect 2816 37539 2862 37578
rect 2816 37505 2822 37539
rect 2856 37505 2862 37539
rect 2816 37466 2862 37505
rect 2816 37432 2822 37466
rect 2856 37432 2862 37466
rect 2816 37393 2862 37432
rect 2816 37359 2822 37393
rect 2856 37359 2862 37393
rect 2816 37320 2862 37359
rect 2816 37286 2822 37320
rect 2856 37286 2862 37320
rect 2816 37247 2862 37286
rect 2816 37213 2822 37247
rect 2856 37213 2862 37247
rect 2816 37174 2862 37213
rect 2816 37140 2822 37174
rect 2856 37140 2862 37174
rect 2816 37102 2862 37140
rect 2816 37068 2822 37102
rect 2856 37068 2862 37102
rect 2816 37030 2862 37068
rect 2816 36996 2822 37030
rect 2856 36996 2862 37030
rect 2816 36958 2862 36996
rect 2816 36924 2822 36958
rect 2856 36924 2862 36958
rect 2816 36886 2862 36924
rect 2816 36852 2822 36886
rect 2856 36852 2862 36886
rect 2816 36814 2862 36852
rect 2816 36780 2822 36814
rect 2856 36780 2862 36814
rect 2816 36742 2862 36780
rect 2816 36708 2822 36742
rect 2856 36708 2862 36742
rect 2816 36670 2862 36708
rect 2816 36636 2822 36670
rect 2856 36636 2862 36670
rect 2816 36598 2862 36636
rect 2816 36564 2822 36598
rect 2856 36564 2862 36598
rect 2816 36526 2862 36564
rect 2816 36492 2822 36526
rect 2856 36492 2862 36526
rect 2816 36454 2862 36492
rect 2816 36420 2822 36454
rect 2856 36420 2862 36454
rect 2816 36382 2862 36420
rect 2816 36348 2822 36382
rect 2856 36348 2862 36382
rect 2816 36310 2862 36348
rect 2816 36276 2822 36310
rect 2856 36276 2862 36310
rect 2816 36238 2862 36276
rect 2816 36204 2822 36238
rect 2856 36204 2862 36238
rect 2816 36166 2862 36204
rect 2816 36132 2822 36166
rect 2856 36132 2862 36166
rect 2816 36094 2862 36132
rect 2816 36060 2822 36094
rect 2856 36060 2862 36094
rect 2816 36022 2862 36060
rect 2816 35988 2822 36022
rect 2856 35988 2862 36022
rect 2816 35950 2862 35988
rect 2816 35916 2822 35950
rect 2856 35916 2862 35950
rect 2816 35878 2862 35916
rect 2816 35844 2822 35878
rect 2856 35844 2862 35878
rect 2816 35806 2862 35844
rect 2816 35772 2822 35806
rect 2856 35772 2862 35806
rect 2816 35734 2862 35772
rect 2816 35700 2822 35734
rect 2856 35700 2862 35734
rect 2816 35662 2862 35700
rect 1187 35643 1287 35649
rect 1187 35591 1211 35643
rect 1263 35591 1287 35643
rect 1187 35579 1287 35591
rect 1187 35527 1211 35579
rect 1263 35527 1287 35579
rect 1187 26202 1287 35527
rect 2816 35628 2822 35662
rect 2856 35628 2862 35662
rect 2816 35590 2862 35628
rect 2816 35556 2822 35590
rect 2856 35556 2862 35590
rect 2816 35518 2862 35556
rect 2816 35484 2822 35518
rect 2856 35484 2862 35518
rect 2816 35446 2862 35484
rect 2816 35412 2822 35446
rect 2856 35412 2862 35446
rect 2816 35374 2862 35412
rect 2816 35340 2822 35374
rect 2856 35340 2862 35374
rect 2816 35302 2862 35340
rect 2816 35268 2822 35302
rect 2856 35268 2862 35302
rect 2816 35230 2862 35268
rect 2816 35196 2822 35230
rect 2856 35196 2862 35230
rect 2816 35158 2862 35196
rect 2816 35124 2822 35158
rect 2856 35124 2862 35158
rect 2816 35086 2862 35124
rect 2816 35052 2822 35086
rect 2856 35052 2862 35086
rect 2816 35014 2862 35052
rect 2816 34980 2822 35014
rect 2856 34980 2862 35014
rect 2816 34942 2862 34980
rect 2816 34908 2822 34942
rect 2856 34908 2862 34942
rect 2816 34870 2862 34908
rect 2816 34836 2822 34870
rect 2856 34836 2862 34870
rect 2816 34798 2862 34836
rect 2816 34764 2822 34798
rect 2856 34764 2862 34798
rect 2816 34726 2862 34764
rect 2816 34692 2822 34726
rect 2856 34692 2862 34726
rect 2816 34654 2862 34692
rect 2816 34620 2822 34654
rect 2856 34620 2862 34654
rect 2816 34582 2862 34620
rect 2816 34548 2822 34582
rect 2856 34548 2862 34582
rect 2816 34510 2862 34548
rect 2816 34476 2822 34510
rect 2856 34476 2862 34510
rect 2816 34438 2862 34476
rect 2816 34404 2822 34438
rect 2856 34404 2862 34438
rect 2816 34366 2862 34404
rect 2816 34332 2822 34366
rect 2856 34332 2862 34366
rect 2816 34294 2862 34332
rect 2816 34260 2822 34294
rect 2856 34260 2862 34294
rect 2816 34222 2862 34260
rect 2816 34188 2822 34222
rect 2856 34188 2862 34222
rect 2816 34150 2862 34188
rect 2816 34116 2822 34150
rect 2856 34116 2862 34150
rect 2816 34078 2862 34116
rect 2816 34044 2822 34078
rect 2856 34044 2862 34078
rect 2816 34006 2862 34044
rect 2816 33972 2822 34006
rect 2856 33972 2862 34006
rect 2816 33934 2862 33972
rect 2816 33900 2822 33934
rect 2856 33900 2862 33934
rect 2816 33862 2862 33900
rect 2816 33828 2822 33862
rect 2856 33828 2862 33862
rect 2816 33790 2862 33828
rect 2816 33756 2822 33790
rect 2856 33756 2862 33790
rect 2816 33718 2862 33756
rect 2816 33684 2822 33718
rect 2856 33684 2862 33718
rect 2816 33646 2862 33684
rect 2816 33612 2822 33646
rect 2856 33612 2862 33646
rect 2816 33574 2862 33612
rect 2816 33540 2822 33574
rect 2856 33540 2862 33574
rect 2816 33502 2862 33540
rect 2816 33468 2822 33502
rect 2856 33468 2862 33502
rect 2816 33430 2862 33468
rect 2816 33396 2822 33430
rect 2856 33396 2862 33430
rect 2816 33358 2862 33396
rect 2816 33324 2822 33358
rect 2856 33324 2862 33358
rect 2816 33286 2862 33324
rect 2816 33252 2822 33286
rect 2856 33252 2862 33286
rect 2816 33214 2862 33252
rect 2816 33180 2822 33214
rect 2856 33180 2862 33214
rect 2816 33142 2862 33180
rect 2816 33108 2822 33142
rect 2856 33108 2862 33142
rect 2816 33070 2862 33108
rect 2816 33036 2822 33070
rect 2856 33036 2862 33070
rect 2816 32998 2862 33036
rect 2816 32964 2822 32998
rect 2856 32964 2862 32998
rect 2816 32926 2862 32964
rect 2816 32892 2822 32926
rect 2856 32892 2862 32926
rect 2816 32854 2862 32892
rect 2816 32820 2822 32854
rect 2856 32820 2862 32854
rect 2816 32782 2862 32820
rect 2816 32748 2822 32782
rect 2856 32748 2862 32782
rect 2816 32710 2862 32748
rect 2816 32676 2822 32710
rect 2856 32676 2862 32710
rect 2816 32638 2862 32676
rect 2816 32604 2822 32638
rect 2856 32604 2862 32638
rect 2816 32566 2862 32604
rect 2816 32532 2822 32566
rect 2856 32532 2862 32566
rect 2816 32494 2862 32532
rect 2816 32460 2822 32494
rect 2856 32460 2862 32494
rect 2816 32422 2862 32460
rect 2816 32388 2822 32422
rect 2856 32388 2862 32422
rect 2816 32350 2862 32388
rect 2816 32316 2822 32350
rect 2856 32316 2862 32350
rect 2816 32278 2862 32316
rect 2816 32244 2822 32278
rect 2856 32244 2862 32278
rect 2816 32206 2862 32244
rect 2816 32172 2822 32206
rect 2856 32172 2862 32206
rect 2816 32134 2862 32172
rect 2816 32100 2822 32134
rect 2856 32100 2862 32134
rect 2816 32062 2862 32100
rect 2816 32028 2822 32062
rect 2856 32028 2862 32062
rect 2816 31990 2862 32028
rect 2816 31956 2822 31990
rect 2856 31956 2862 31990
rect 2816 31918 2862 31956
rect 2816 31884 2822 31918
rect 2856 31884 2862 31918
rect 2816 31846 2862 31884
rect 2816 31812 2822 31846
rect 2856 31812 2862 31846
rect 2816 31774 2862 31812
rect 2816 31740 2822 31774
rect 2856 31740 2862 31774
rect 2816 31702 2862 31740
rect 2816 31668 2822 31702
rect 2856 31668 2862 31702
rect 2816 31630 2862 31668
rect 2816 31596 2822 31630
rect 2856 31596 2862 31630
rect 2816 31558 2862 31596
rect 2816 31524 2822 31558
rect 2856 31524 2862 31558
rect 2816 31486 2862 31524
rect 2816 31452 2822 31486
rect 2856 31452 2862 31486
rect 2816 31414 2862 31452
rect 2816 31380 2822 31414
rect 2856 31380 2862 31414
rect 2816 31342 2862 31380
rect 2816 31308 2822 31342
rect 2856 31308 2862 31342
rect 2816 31270 2862 31308
rect 2816 31236 2822 31270
rect 2856 31236 2862 31270
rect 2816 31198 2862 31236
rect 2816 31164 2822 31198
rect 2856 31164 2862 31198
rect 2816 31126 2862 31164
rect 2816 31092 2822 31126
rect 2856 31092 2862 31126
rect 2816 31054 2862 31092
rect 2816 31020 2822 31054
rect 2856 31020 2862 31054
rect 2816 30982 2862 31020
rect 2816 30948 2822 30982
rect 2856 30948 2862 30982
rect 2816 30910 2862 30948
rect 2816 30876 2822 30910
rect 2856 30876 2862 30910
rect 2816 30838 2862 30876
rect 2816 30804 2822 30838
rect 2856 30804 2862 30838
rect 2816 30766 2862 30804
rect 2816 30732 2822 30766
rect 2856 30732 2862 30766
rect 2816 30694 2862 30732
rect 2816 30660 2822 30694
rect 2856 30660 2862 30694
rect 2816 30622 2862 30660
rect 2816 30588 2822 30622
rect 2856 30588 2862 30622
rect 2816 30550 2862 30588
rect 2816 30516 2822 30550
rect 2856 30516 2862 30550
rect 2816 30478 2862 30516
rect 2816 30444 2822 30478
rect 2856 30444 2862 30478
rect 2816 30406 2862 30444
rect 2816 30372 2822 30406
rect 2856 30372 2862 30406
rect 2816 30334 2862 30372
rect 2816 30300 2822 30334
rect 2856 30300 2862 30334
rect 2816 30262 2862 30300
rect 2816 30228 2822 30262
rect 2856 30228 2862 30262
rect 2816 30190 2862 30228
rect 2816 30156 2822 30190
rect 2856 30156 2862 30190
rect 2816 30118 2862 30156
rect 2816 30084 2822 30118
rect 2856 30084 2862 30118
rect 2816 30046 2862 30084
rect 2816 30012 2822 30046
rect 2856 30012 2862 30046
rect 2816 29974 2862 30012
rect 2816 29940 2822 29974
rect 2856 29940 2862 29974
rect 2816 29902 2862 29940
rect 2816 29868 2822 29902
rect 2856 29868 2862 29902
rect 2816 29830 2862 29868
rect 2816 29796 2822 29830
rect 2856 29796 2862 29830
rect 2816 29758 2862 29796
rect 2816 29724 2822 29758
rect 2856 29724 2862 29758
rect 2816 29686 2862 29724
rect 2816 29652 2822 29686
rect 2856 29652 2862 29686
rect 2816 29614 2862 29652
rect 2816 29580 2822 29614
rect 2856 29580 2862 29614
rect 2816 29542 2862 29580
rect 2816 29508 2822 29542
rect 2856 29508 2862 29542
rect 2627 29435 2633 29487
rect 2685 29435 2730 29487
rect 2782 29435 2788 29487
rect 2627 29411 2788 29435
rect 2627 29359 2633 29411
rect 2685 29359 2730 29411
rect 2782 29359 2788 29411
rect 1239 26150 1287 26202
rect 1187 26138 1287 26150
rect 1239 26086 1287 26138
rect 908 25807 1008 25813
rect 908 25755 932 25807
rect 984 25755 1008 25807
rect 908 25743 1008 25755
rect 908 25691 932 25743
rect 984 25691 1008 25743
rect 908 16786 1008 25691
rect 960 16734 1008 16786
rect 908 16720 1008 16734
rect 960 16668 1008 16720
rect 908 16654 1008 16668
rect 960 16602 1008 16654
rect 908 16588 1008 16602
rect 960 16536 1008 16588
rect 908 16530 1008 16536
rect 1187 25601 1287 26086
rect 1239 25549 1287 25601
rect 1187 25537 1287 25549
rect 1239 25485 1287 25537
rect 1187 16901 1287 25485
rect 2288 28957 2294 29009
rect 2346 28957 2391 29009
rect 2443 28957 2449 29009
rect 2288 22530 2449 28957
rect 2288 22478 2294 22530
rect 2346 22478 2391 22530
rect 2443 22478 2449 22530
rect 2288 22454 2449 22478
rect 2288 22402 2294 22454
rect 2346 22402 2391 22454
rect 2443 22402 2449 22454
rect 2288 19271 2449 22402
rect 2288 19219 2294 19271
rect 2346 19219 2391 19271
rect 2443 19219 2449 19271
rect 2288 19207 2449 19219
rect 2288 19155 2294 19207
rect 2346 19155 2391 19207
rect 2443 19155 2449 19207
rect 2288 17619 2449 19155
rect 2627 21692 2788 29359
rect 2816 29470 2862 29508
rect 2816 29436 2822 29470
rect 2856 29436 2862 29470
rect 2816 29398 2862 29436
rect 2816 29364 2822 29398
rect 2856 29364 2862 29398
rect 2816 29326 2862 29364
rect 2816 29292 2822 29326
rect 2856 29292 2862 29326
rect 2816 29254 2862 29292
rect 2816 29220 2822 29254
rect 2856 29220 2862 29254
rect 2816 29182 2862 29220
rect 2816 29148 2822 29182
rect 2856 29148 2862 29182
rect 2816 29110 2862 29148
rect 2816 29076 2822 29110
rect 2856 29076 2862 29110
rect 2816 29038 2862 29076
rect 2816 29004 2822 29038
rect 2856 29004 2862 29038
rect 2816 28966 2862 29004
rect 2816 28932 2822 28966
rect 2856 28932 2862 28966
rect 2816 28894 2862 28932
rect 2816 28860 2822 28894
rect 2856 28860 2862 28894
rect 2816 28822 2862 28860
rect 2816 28788 2822 28822
rect 2856 28788 2862 28822
rect 2816 28750 2862 28788
rect 2816 28716 2822 28750
rect 2856 28716 2862 28750
rect 2816 28678 2862 28716
rect 2816 28644 2822 28678
rect 2856 28644 2862 28678
rect 2816 28606 2862 28644
rect 2816 28572 2822 28606
rect 2856 28572 2862 28606
rect 2816 28534 2862 28572
rect 2816 28500 2822 28534
rect 2856 28500 2862 28534
rect 2816 28462 2862 28500
rect 2816 28428 2822 28462
rect 2856 28428 2862 28462
rect 2816 28390 2862 28428
rect 3076 39614 5370 39620
rect 3076 39580 3157 39614
rect 3191 39580 3232 39614
rect 3266 39580 3307 39614
rect 3341 39580 3382 39614
rect 3416 39580 3457 39614
rect 3491 39580 3532 39614
rect 3566 39580 3607 39614
rect 3641 39580 3682 39614
rect 3716 39580 3757 39614
rect 3791 39580 3832 39614
rect 3866 39580 3907 39614
rect 3941 39580 3982 39614
rect 4016 39580 4057 39614
rect 4091 39580 4132 39614
rect 4166 39580 4207 39614
rect 4241 39580 4282 39614
rect 4316 39580 4357 39614
rect 4391 39580 4433 39614
rect 4467 39580 4509 39614
rect 4543 39580 4619 39614
rect 4653 39580 4698 39614
rect 4732 39580 4778 39614
rect 4812 39580 4858 39614
rect 4892 39580 4938 39614
rect 4972 39580 5018 39614
rect 5052 39580 5098 39614
rect 5132 39580 5178 39614
rect 5212 39580 5258 39614
rect 5292 39580 5370 39614
rect 3076 39574 5370 39580
rect 3076 39542 3122 39574
rect 3076 39508 3082 39542
rect 3116 39508 3122 39542
rect 3076 39469 3122 39508
rect 3076 39435 3082 39469
rect 3116 39435 3122 39469
rect 3076 39396 3122 39435
rect 3076 39362 3082 39396
rect 3116 39362 3122 39396
rect 3076 39323 3122 39362
rect 3076 39289 3082 39323
rect 3116 39289 3122 39323
rect 3076 39250 3122 39289
rect 3076 39216 3082 39250
rect 3116 39216 3122 39250
rect 3076 39177 3122 39216
rect 3076 39143 3082 39177
rect 3116 39143 3122 39177
rect 3076 39104 3122 39143
rect 3076 39070 3082 39104
rect 3116 39070 3122 39104
rect 3076 39031 3122 39070
rect 3076 38997 3082 39031
rect 3116 38997 3122 39031
rect 3076 38958 3122 38997
rect 3076 38924 3082 38958
rect 3116 38924 3122 38958
rect 3076 38885 3122 38924
rect 3076 38851 3082 38885
rect 3116 38851 3122 38885
rect 3076 38812 3122 38851
rect 3076 38778 3082 38812
rect 3116 38778 3122 38812
rect 3076 38739 3122 38778
rect 3076 38705 3082 38739
rect 3116 38705 3122 38739
rect 3076 38666 3122 38705
rect 3076 38632 3082 38666
rect 3116 38632 3122 38666
rect 3076 38593 3122 38632
rect 3076 38559 3082 38593
rect 3116 38559 3122 38593
rect 3076 38520 3122 38559
rect 3076 38486 3082 38520
rect 3116 38486 3122 38520
rect 3076 38447 3122 38486
rect 3076 38413 3082 38447
rect 3116 38413 3122 38447
rect 3076 38374 3122 38413
rect 3076 38340 3082 38374
rect 3116 38340 3122 38374
rect 3076 38301 3122 38340
rect 3076 38267 3082 38301
rect 3116 38267 3122 38301
rect 3076 38228 3122 38267
rect 3076 38194 3082 38228
rect 3116 38194 3122 38228
rect 3076 38155 3122 38194
rect 3076 38121 3082 38155
rect 3116 38121 3122 38155
rect 3076 38082 3122 38121
rect 3076 38048 3082 38082
rect 3116 38048 3122 38082
rect 3076 38010 3122 38048
rect 3076 37976 3082 38010
rect 3116 37976 3122 38010
rect 3076 37938 3122 37976
rect 3076 37904 3082 37938
rect 3116 37904 3122 37938
rect 3076 37866 3122 37904
rect 3076 37832 3082 37866
rect 3116 37832 3122 37866
rect 3076 37794 3122 37832
rect 3076 37760 3082 37794
rect 3116 37760 3122 37794
rect 3076 37722 3122 37760
rect 3076 37688 3082 37722
rect 3116 37688 3122 37722
rect 3076 37650 3122 37688
rect 3076 37616 3082 37650
rect 3116 37616 3122 37650
rect 3076 37578 3122 37616
rect 3076 37544 3082 37578
rect 3116 37544 3122 37578
rect 3076 37506 3122 37544
rect 3076 37472 3082 37506
rect 3116 37472 3122 37506
rect 3076 37434 3122 37472
rect 3076 37400 3082 37434
rect 3116 37400 3122 37434
rect 3076 37362 3122 37400
rect 3076 37328 3082 37362
rect 3116 37328 3122 37362
rect 3076 37290 3122 37328
rect 3076 37256 3082 37290
rect 3116 37256 3122 37290
rect 3076 37218 3122 37256
rect 3076 37184 3082 37218
rect 3116 37184 3122 37218
rect 3076 37146 3122 37184
rect 3076 37112 3082 37146
rect 3116 37112 3122 37146
rect 3076 37074 3122 37112
rect 3076 37040 3082 37074
rect 3116 37040 3122 37074
rect 3076 37002 3122 37040
rect 3076 36968 3082 37002
rect 3116 36968 3122 37002
rect 3076 36930 3122 36968
rect 3076 36896 3082 36930
rect 3116 36896 3122 36930
rect 3076 36858 3122 36896
rect 3076 36824 3082 36858
rect 3116 36824 3122 36858
rect 3076 36786 3122 36824
rect 3076 36752 3082 36786
rect 3116 36752 3122 36786
rect 3076 36714 3122 36752
rect 3076 36680 3082 36714
rect 3116 36680 3122 36714
rect 3076 36642 3122 36680
rect 3076 36608 3082 36642
rect 3116 36608 3122 36642
rect 3076 36570 3122 36608
rect 3076 36536 3082 36570
rect 3116 36536 3122 36570
rect 3076 36498 3122 36536
rect 3076 36464 3082 36498
rect 3116 36464 3122 36498
rect 3076 36426 3122 36464
rect 3076 36392 3082 36426
rect 3116 36392 3122 36426
rect 3076 36354 3122 36392
rect 3076 36320 3082 36354
rect 3116 36320 3122 36354
rect 3076 36282 3122 36320
rect 3076 36248 3082 36282
rect 3116 36248 3122 36282
rect 3076 36210 3122 36248
rect 3076 36176 3082 36210
rect 3116 36176 3122 36210
rect 3076 36138 3122 36176
rect 3076 36104 3082 36138
rect 3116 36104 3122 36138
rect 3076 36066 3122 36104
rect 3076 36032 3082 36066
rect 3116 36032 3122 36066
rect 3076 35994 3122 36032
rect 3076 35960 3082 35994
rect 3116 35960 3122 35994
rect 3076 35922 3122 35960
rect 3076 35888 3082 35922
rect 3116 35888 3122 35922
rect 3076 35850 3122 35888
rect 3076 35816 3082 35850
rect 3116 35816 3122 35850
rect 3076 35778 3122 35816
rect 3076 35744 3082 35778
rect 3116 35744 3122 35778
rect 3076 35706 3122 35744
rect 3076 35672 3082 35706
rect 3116 35672 3122 35706
rect 3076 35634 3122 35672
rect 3168 39353 3214 39365
rect 3168 39319 3174 39353
rect 3208 39319 3214 39353
rect 3168 39281 3214 39319
rect 3168 39247 3174 39281
rect 3208 39247 3214 39281
rect 3168 39209 3214 39247
rect 3168 39175 3174 39209
rect 3208 39175 3214 39209
rect 3168 39137 3214 39175
rect 3168 39103 3174 39137
rect 3208 39103 3214 39137
rect 3168 39065 3214 39103
rect 3168 39031 3174 39065
rect 3208 39031 3214 39065
rect 3168 38993 3214 39031
rect 3168 38959 3174 38993
rect 3208 38959 3214 38993
rect 3168 38921 3214 38959
rect 3168 38887 3174 38921
rect 3208 38887 3214 38921
rect 3168 38849 3214 38887
rect 3168 38815 3174 38849
rect 3208 38815 3214 38849
rect 3168 38777 3214 38815
rect 3168 38743 3174 38777
rect 3208 38743 3214 38777
rect 3168 38705 3214 38743
rect 3168 38671 3174 38705
rect 3208 38671 3214 38705
rect 3168 38633 3214 38671
rect 3168 38599 3174 38633
rect 3208 38599 3214 38633
rect 3168 38561 3214 38599
rect 3168 38527 3174 38561
rect 3208 38527 3214 38561
rect 3168 38489 3214 38527
rect 3168 38455 3174 38489
rect 3208 38455 3214 38489
rect 3168 38417 3214 38455
rect 3168 38383 3174 38417
rect 3208 38383 3214 38417
rect 3168 38345 3214 38383
rect 3168 38311 3174 38345
rect 3208 38311 3214 38345
rect 3168 38273 3214 38311
rect 3168 38239 3174 38273
rect 3208 38239 3214 38273
rect 3168 38201 3214 38239
rect 3168 38167 3174 38201
rect 3208 38167 3214 38201
rect 3168 38129 3214 38167
rect 3168 38095 3174 38129
rect 3208 38095 3214 38129
rect 3168 38057 3214 38095
rect 3168 38023 3174 38057
rect 3208 38023 3214 38057
rect 3168 37985 3214 38023
rect 3168 37951 3174 37985
rect 3208 37951 3214 37985
rect 3168 37913 3214 37951
rect 3168 37879 3174 37913
rect 3208 37879 3214 37913
rect 3168 37841 3214 37879
rect 3168 37807 3174 37841
rect 3208 37807 3214 37841
rect 3168 37769 3214 37807
rect 3168 37735 3174 37769
rect 3208 37735 3214 37769
rect 3168 37697 3214 37735
rect 3168 37663 3174 37697
rect 3208 37663 3214 37697
rect 3168 37625 3214 37663
rect 3168 37591 3174 37625
rect 3208 37591 3214 37625
rect 3168 37553 3214 37591
rect 3168 37519 3174 37553
rect 3208 37519 3214 37553
rect 3168 37481 3214 37519
rect 3168 37447 3174 37481
rect 3208 37447 3214 37481
rect 3168 37409 3214 37447
rect 3168 37375 3174 37409
rect 3208 37375 3214 37409
rect 3168 37337 3214 37375
rect 3168 37303 3174 37337
rect 3208 37303 3214 37337
rect 3168 37265 3214 37303
rect 3168 37231 3174 37265
rect 3208 37231 3214 37265
rect 3168 37193 3214 37231
rect 3168 37159 3174 37193
rect 3208 37159 3214 37193
rect 3168 37121 3214 37159
rect 3168 37087 3174 37121
rect 3208 37087 3214 37121
rect 3168 37049 3214 37087
rect 3168 37015 3174 37049
rect 3208 37015 3214 37049
rect 3168 36977 3214 37015
rect 3168 36943 3174 36977
rect 3208 36943 3214 36977
rect 3168 36905 3214 36943
rect 3168 36871 3174 36905
rect 3208 36871 3214 36905
rect 3168 36833 3214 36871
rect 3168 36799 3174 36833
rect 3208 36799 3214 36833
rect 3168 36761 3214 36799
rect 3168 36727 3174 36761
rect 3208 36727 3214 36761
rect 3168 36689 3214 36727
rect 3168 36655 3174 36689
rect 3208 36655 3214 36689
rect 3168 36617 3214 36655
rect 3168 36583 3174 36617
rect 3208 36583 3214 36617
rect 3168 36545 3214 36583
rect 3168 36511 3174 36545
rect 3208 36511 3214 36545
rect 3168 36473 3214 36511
rect 3168 36439 3174 36473
rect 3208 36439 3214 36473
rect 3168 36401 3214 36439
rect 3168 36367 3174 36401
rect 3208 36367 3214 36401
rect 3168 36329 3214 36367
rect 3168 36295 3174 36329
rect 3208 36295 3214 36329
rect 3168 36257 3214 36295
rect 3168 36223 3174 36257
rect 3208 36223 3214 36257
rect 3168 36185 3214 36223
rect 3168 36151 3174 36185
rect 3208 36151 3214 36185
rect 3168 36113 3214 36151
rect 3168 36079 3174 36113
rect 3208 36079 3214 36113
rect 3168 36041 3214 36079
rect 3168 36007 3174 36041
rect 3208 36007 3214 36041
rect 3168 35969 3214 36007
rect 3168 35935 3174 35969
rect 3208 35935 3214 35969
rect 3168 35897 3214 35935
rect 3168 35863 3174 35897
rect 3208 35863 3214 35897
rect 3168 35825 3214 35863
rect 3168 35791 3174 35825
rect 3208 35791 3214 35825
rect 3168 35753 3214 35791
rect 3168 35719 3174 35753
rect 3208 35719 3214 35753
rect 3168 35681 3214 35719
rect 3168 35649 3174 35681
rect 3076 35600 3082 35634
rect 3116 35600 3122 35634
rect 3076 35562 3122 35600
rect 3076 35528 3082 35562
rect 3116 35528 3122 35562
rect 3076 35490 3122 35528
rect 3165 35647 3174 35649
rect 3208 35649 3214 35681
rect 4489 39201 5273 39574
rect 5324 39542 5370 39574
rect 5324 39508 5330 39542
rect 5364 39508 5370 39542
rect 5324 39470 5370 39508
rect 5324 39436 5330 39470
rect 5364 39436 5370 39470
rect 5324 39398 5370 39436
rect 5324 39364 5330 39398
rect 5364 39364 5370 39398
rect 5324 39326 5370 39364
rect 5324 39292 5330 39326
rect 5364 39292 5370 39326
rect 5324 39254 5370 39292
rect 5324 39220 5330 39254
rect 5364 39220 5370 39254
rect 5324 39201 5370 39220
rect 7740 39586 7786 39624
rect 7740 39552 7746 39586
rect 7780 39552 7786 39586
rect 7740 39514 7786 39552
rect 7740 39480 7746 39514
rect 7780 39480 7786 39514
rect 7740 39442 7786 39480
rect 7740 39408 7746 39442
rect 7780 39408 7786 39442
rect 7740 39370 7786 39408
rect 7740 39336 7746 39370
rect 7780 39336 7786 39370
rect 7740 39298 7786 39336
rect 7740 39264 7746 39298
rect 7780 39264 7786 39298
rect 7740 39226 7786 39264
rect 4489 39195 5447 39201
rect 4489 39143 4666 39195
rect 4718 39143 4732 39195
rect 4784 39143 4798 39195
rect 4850 39143 4864 39195
rect 4916 39143 4930 39195
rect 4982 39143 4996 39195
rect 5048 39143 5062 39195
rect 5114 39143 5128 39195
rect 5180 39143 5194 39195
rect 5246 39143 5260 39195
rect 5312 39143 5326 39195
rect 5378 39143 5392 39195
rect 5444 39143 5447 39195
rect 4489 39131 5447 39143
rect 4489 39079 4666 39131
rect 4718 39079 4732 39131
rect 4784 39079 4798 39131
rect 4850 39079 4864 39131
rect 4916 39079 4930 39131
rect 4982 39079 4996 39131
rect 5048 39079 5062 39131
rect 5114 39079 5128 39131
rect 5180 39079 5194 39131
rect 5246 39079 5260 39131
rect 5312 39079 5326 39131
rect 5378 39079 5392 39131
rect 5444 39079 5447 39131
rect 4489 39076 5330 39079
rect 5364 39076 5447 39079
rect 4489 39067 5447 39076
rect 4489 39015 4666 39067
rect 4718 39015 4732 39067
rect 4784 39015 4798 39067
rect 4850 39015 4864 39067
rect 4916 39015 4930 39067
rect 4982 39015 4996 39067
rect 5048 39015 5062 39067
rect 5114 39015 5128 39067
rect 5180 39015 5194 39067
rect 5246 39015 5260 39067
rect 5312 39015 5326 39067
rect 5378 39015 5392 39067
rect 5444 39015 5447 39067
rect 4489 39004 5330 39015
rect 5364 39004 5447 39015
rect 4489 39003 5447 39004
rect 4489 38951 4666 39003
rect 4718 38951 4732 39003
rect 4784 38951 4798 39003
rect 4850 38951 4864 39003
rect 4916 38951 4930 39003
rect 4982 38951 4996 39003
rect 5048 38951 5062 39003
rect 5114 38951 5128 39003
rect 5180 38951 5194 39003
rect 5246 38951 5260 39003
rect 5312 38951 5326 39003
rect 5378 38951 5392 39003
rect 5444 38951 5447 39003
rect 4489 38939 5330 38951
rect 5364 38939 5447 38951
rect 4489 38887 4666 38939
rect 4718 38887 4732 38939
rect 4784 38887 4798 38939
rect 4850 38887 4864 38939
rect 4916 38887 4930 38939
rect 4982 38887 4996 38939
rect 5048 38887 5062 38939
rect 5114 38887 5128 38939
rect 5180 38887 5194 38939
rect 5246 38887 5260 38939
rect 5312 38887 5326 38939
rect 5378 38887 5392 38939
rect 5444 38887 5447 38939
rect 4489 38875 5330 38887
rect 5364 38875 5447 38887
rect 4489 38823 4666 38875
rect 4718 38823 4732 38875
rect 4784 38823 4798 38875
rect 4850 38823 4864 38875
rect 4916 38823 4930 38875
rect 4982 38823 4996 38875
rect 5048 38823 5062 38875
rect 5114 38823 5128 38875
rect 5180 38823 5194 38875
rect 5246 38823 5260 38875
rect 5312 38823 5326 38875
rect 5378 38823 5392 38875
rect 5444 38823 5447 38875
rect 4489 38822 5447 38823
rect 4489 38811 5330 38822
rect 5364 38811 5447 38822
rect 4489 38759 4666 38811
rect 4718 38759 4732 38811
rect 4784 38759 4798 38811
rect 4850 38759 4864 38811
rect 4916 38759 4930 38811
rect 4982 38759 4996 38811
rect 5048 38759 5062 38811
rect 5114 38759 5128 38811
rect 5180 38759 5194 38811
rect 5246 38759 5260 38811
rect 5312 38759 5326 38811
rect 5378 38759 5392 38811
rect 5444 38759 5447 38811
rect 4489 38750 5447 38759
rect 4489 38747 5330 38750
rect 5364 38747 5447 38750
rect 4489 38695 4666 38747
rect 4718 38695 4732 38747
rect 4784 38695 4798 38747
rect 4850 38695 4864 38747
rect 4916 38695 4930 38747
rect 4982 38695 4996 38747
rect 5048 38695 5062 38747
rect 5114 38695 5128 38747
rect 5180 38695 5194 38747
rect 5246 38695 5260 38747
rect 5312 38695 5326 38747
rect 5378 38695 5392 38747
rect 5444 38695 5447 38747
rect 4489 38683 5447 38695
rect 4489 38631 4666 38683
rect 4718 38631 4732 38683
rect 4784 38631 4798 38683
rect 4850 38631 4864 38683
rect 4916 38631 4930 38683
rect 4982 38631 4996 38683
rect 5048 38631 5062 38683
rect 5114 38631 5128 38683
rect 5180 38631 5194 38683
rect 5246 38631 5260 38683
rect 5312 38631 5326 38683
rect 5378 38631 5392 38683
rect 5444 38631 5447 38683
rect 4489 38619 5447 38631
rect 4489 38567 4666 38619
rect 4718 38567 4732 38619
rect 4784 38567 4798 38619
rect 4850 38567 4864 38619
rect 4916 38567 4930 38619
rect 4982 38567 4996 38619
rect 5048 38567 5062 38619
rect 5114 38567 5128 38619
rect 5180 38567 5194 38619
rect 5246 38567 5260 38619
rect 5312 38567 5326 38619
rect 5378 38567 5392 38619
rect 5444 38567 5447 38619
rect 4489 38555 5447 38567
rect 4489 38503 4666 38555
rect 4718 38503 4732 38555
rect 4784 38503 4798 38555
rect 4850 38503 4864 38555
rect 4916 38503 4930 38555
rect 4982 38503 4996 38555
rect 5048 38503 5062 38555
rect 5114 38503 5128 38555
rect 5180 38503 5194 38555
rect 5246 38503 5260 38555
rect 5312 38503 5326 38555
rect 5378 38503 5392 38555
rect 5444 38503 5447 38555
rect 4489 38500 5330 38503
rect 5364 38500 5447 38503
rect 4489 38491 5447 38500
rect 4489 38439 4666 38491
rect 4718 38439 4732 38491
rect 4784 38439 4798 38491
rect 4850 38439 4864 38491
rect 4916 38439 4930 38491
rect 4982 38439 4996 38491
rect 5048 38439 5062 38491
rect 5114 38439 5128 38491
rect 5180 38439 5194 38491
rect 5246 38439 5260 38491
rect 5312 38439 5326 38491
rect 5378 38439 5392 38491
rect 5444 38439 5447 38491
rect 4489 38428 5330 38439
rect 5364 38428 5447 38439
rect 4489 38427 5447 38428
rect 4489 38375 4666 38427
rect 4718 38375 4732 38427
rect 4784 38375 4798 38427
rect 4850 38375 4864 38427
rect 4916 38375 4930 38427
rect 4982 38375 4996 38427
rect 5048 38375 5062 38427
rect 5114 38375 5128 38427
rect 5180 38375 5194 38427
rect 5246 38375 5260 38427
rect 5312 38375 5326 38427
rect 5378 38375 5392 38427
rect 5444 38375 5447 38427
rect 4489 38363 5330 38375
rect 5364 38363 5447 38375
rect 4489 38311 4666 38363
rect 4718 38311 4732 38363
rect 4784 38311 4798 38363
rect 4850 38311 4864 38363
rect 4916 38311 4930 38363
rect 4982 38311 4996 38363
rect 5048 38311 5062 38363
rect 5114 38311 5128 38363
rect 5180 38311 5194 38363
rect 5246 38311 5260 38363
rect 5312 38311 5326 38363
rect 5378 38311 5392 38363
rect 5444 38311 5447 38363
rect 4489 38299 5330 38311
rect 5364 38299 5447 38311
rect 4489 38247 4666 38299
rect 4718 38247 4732 38299
rect 4784 38247 4798 38299
rect 4850 38247 4864 38299
rect 4916 38247 4930 38299
rect 4982 38247 4996 38299
rect 5048 38247 5062 38299
rect 5114 38247 5128 38299
rect 5180 38247 5194 38299
rect 5246 38247 5260 38299
rect 5312 38247 5326 38299
rect 5378 38247 5392 38299
rect 5444 38247 5447 38299
rect 4489 38246 5447 38247
rect 4489 38235 5330 38246
rect 5364 38235 5447 38246
rect 4489 38183 4666 38235
rect 4718 38183 4732 38235
rect 4784 38183 4798 38235
rect 4850 38183 4864 38235
rect 4916 38183 4930 38235
rect 4982 38183 4996 38235
rect 5048 38183 5062 38235
rect 5114 38183 5128 38235
rect 5180 38183 5194 38235
rect 5246 38183 5260 38235
rect 5312 38183 5326 38235
rect 5378 38183 5392 38235
rect 5444 38183 5447 38235
rect 4489 38174 5447 38183
rect 4489 38171 5330 38174
rect 5364 38171 5447 38174
rect 4489 38119 4666 38171
rect 4718 38119 4732 38171
rect 4784 38119 4798 38171
rect 4850 38119 4864 38171
rect 4916 38119 4930 38171
rect 4982 38119 4996 38171
rect 5048 38119 5062 38171
rect 5114 38119 5128 38171
rect 5180 38119 5194 38171
rect 5246 38119 5260 38171
rect 5312 38119 5326 38171
rect 5378 38119 5392 38171
rect 5444 38119 5447 38171
rect 4489 38107 5447 38119
rect 4489 38055 4666 38107
rect 4718 38055 4732 38107
rect 4784 38055 4798 38107
rect 4850 38055 4864 38107
rect 4916 38055 4930 38107
rect 4982 38055 4996 38107
rect 5048 38055 5062 38107
rect 5114 38055 5128 38107
rect 5180 38055 5194 38107
rect 5246 38055 5260 38107
rect 5312 38055 5326 38107
rect 5378 38055 5392 38107
rect 5444 38055 5447 38107
rect 4489 38043 5447 38055
rect 4489 37991 4666 38043
rect 4718 37991 4732 38043
rect 4784 37991 4798 38043
rect 4850 37991 4864 38043
rect 4916 37991 4930 38043
rect 4982 37991 4996 38043
rect 5048 37991 5062 38043
rect 5114 37991 5128 38043
rect 5180 37991 5194 38043
rect 5246 37991 5260 38043
rect 5312 37991 5326 38043
rect 5378 37991 5392 38043
rect 5444 37991 5447 38043
rect 4489 37979 5447 37991
rect 4489 37927 4666 37979
rect 4718 37927 4732 37979
rect 4784 37927 4798 37979
rect 4850 37927 4864 37979
rect 4916 37927 4930 37979
rect 4982 37927 4996 37979
rect 5048 37927 5062 37979
rect 5114 37927 5128 37979
rect 5180 37927 5194 37979
rect 5246 37927 5260 37979
rect 5312 37927 5326 37979
rect 5378 37927 5392 37979
rect 5444 37927 5447 37979
rect 4489 37924 5330 37927
rect 5364 37924 5447 37927
rect 4489 37915 5447 37924
rect 4489 37863 4666 37915
rect 4718 37863 4732 37915
rect 4784 37863 4798 37915
rect 4850 37863 4864 37915
rect 4916 37863 4930 37915
rect 4982 37863 4996 37915
rect 5048 37863 5062 37915
rect 5114 37863 5128 37915
rect 5180 37863 5194 37915
rect 5246 37863 5260 37915
rect 5312 37863 5326 37915
rect 5378 37863 5392 37915
rect 5444 37863 5447 37915
rect 4489 37852 5330 37863
rect 5364 37852 5447 37863
rect 4489 37851 5447 37852
rect 4489 37799 4666 37851
rect 4718 37799 4732 37851
rect 4784 37799 4798 37851
rect 4850 37799 4864 37851
rect 4916 37799 4930 37851
rect 4982 37799 4996 37851
rect 5048 37799 5062 37851
rect 5114 37799 5128 37851
rect 5180 37799 5194 37851
rect 5246 37799 5260 37851
rect 5312 37799 5326 37851
rect 5378 37799 5392 37851
rect 5444 37799 5447 37851
rect 4489 37787 5330 37799
rect 5364 37787 5447 37799
rect 4489 37735 4666 37787
rect 4718 37735 4732 37787
rect 4784 37735 4798 37787
rect 4850 37735 4864 37787
rect 4916 37735 4930 37787
rect 4982 37735 4996 37787
rect 5048 37735 5062 37787
rect 5114 37735 5128 37787
rect 5180 37735 5194 37787
rect 5246 37735 5260 37787
rect 5312 37735 5326 37787
rect 5378 37735 5392 37787
rect 5444 37735 5447 37787
rect 4489 37723 5330 37735
rect 5364 37723 5447 37735
rect 4489 37671 4666 37723
rect 4718 37671 4732 37723
rect 4784 37671 4798 37723
rect 4850 37671 4864 37723
rect 4916 37671 4930 37723
rect 4982 37671 4996 37723
rect 5048 37671 5062 37723
rect 5114 37671 5128 37723
rect 5180 37671 5194 37723
rect 5246 37671 5260 37723
rect 5312 37671 5326 37723
rect 5378 37671 5392 37723
rect 5444 37671 5447 37723
rect 4489 37670 5447 37671
rect 4489 37659 5330 37670
rect 5364 37659 5447 37670
rect 4489 37607 4666 37659
rect 4718 37607 4732 37659
rect 4784 37607 4798 37659
rect 4850 37607 4864 37659
rect 4916 37607 4930 37659
rect 4982 37607 4996 37659
rect 5048 37607 5062 37659
rect 5114 37607 5128 37659
rect 5180 37607 5194 37659
rect 5246 37607 5260 37659
rect 5312 37607 5326 37659
rect 5378 37607 5392 37659
rect 5444 37607 5447 37659
rect 4489 37598 5447 37607
rect 4489 37595 5330 37598
rect 5364 37595 5447 37598
rect 4489 37543 4666 37595
rect 4718 37543 4732 37595
rect 4784 37543 4798 37595
rect 4850 37543 4864 37595
rect 4916 37543 4930 37595
rect 4982 37543 4996 37595
rect 5048 37543 5062 37595
rect 5114 37543 5128 37595
rect 5180 37543 5194 37595
rect 5246 37543 5260 37595
rect 5312 37543 5326 37595
rect 5378 37543 5392 37595
rect 5444 37543 5447 37595
rect 4489 37531 5447 37543
rect 4489 37479 4666 37531
rect 4718 37479 4732 37531
rect 4784 37479 4798 37531
rect 4850 37479 4864 37531
rect 4916 37479 4930 37531
rect 4982 37479 4996 37531
rect 5048 37479 5062 37531
rect 5114 37479 5128 37531
rect 5180 37479 5194 37531
rect 5246 37479 5260 37531
rect 5312 37479 5326 37531
rect 5378 37479 5392 37531
rect 5444 37479 5447 37531
rect 4489 37467 5447 37479
rect 4489 37415 4666 37467
rect 4718 37415 4732 37467
rect 4784 37415 4798 37467
rect 4850 37415 4864 37467
rect 4916 37415 4930 37467
rect 4982 37415 4996 37467
rect 5048 37415 5062 37467
rect 5114 37415 5128 37467
rect 5180 37415 5194 37467
rect 5246 37415 5260 37467
rect 5312 37415 5326 37467
rect 5378 37415 5392 37467
rect 5444 37415 5447 37467
rect 4489 37403 5447 37415
rect 4489 37351 4666 37403
rect 4718 37351 4732 37403
rect 4784 37351 4798 37403
rect 4850 37351 4864 37403
rect 4916 37351 4930 37403
rect 4982 37351 4996 37403
rect 5048 37351 5062 37403
rect 5114 37351 5128 37403
rect 5180 37351 5194 37403
rect 5246 37351 5260 37403
rect 5312 37351 5326 37403
rect 5378 37351 5392 37403
rect 5444 37351 5447 37403
rect 4489 37348 5330 37351
rect 5364 37348 5447 37351
rect 4489 37339 5447 37348
rect 4489 37287 4666 37339
rect 4718 37287 4732 37339
rect 4784 37287 4798 37339
rect 4850 37287 4864 37339
rect 4916 37287 4930 37339
rect 4982 37287 4996 37339
rect 5048 37287 5062 37339
rect 5114 37287 5128 37339
rect 5180 37287 5194 37339
rect 5246 37287 5260 37339
rect 5312 37287 5326 37339
rect 5378 37287 5392 37339
rect 5444 37287 5447 37339
rect 4489 37276 5330 37287
rect 5364 37276 5447 37287
rect 4489 37275 5447 37276
rect 4489 37223 4666 37275
rect 4718 37223 4732 37275
rect 4784 37223 4798 37275
rect 4850 37223 4864 37275
rect 4916 37223 4930 37275
rect 4982 37223 4996 37275
rect 5048 37223 5062 37275
rect 5114 37223 5128 37275
rect 5180 37223 5194 37275
rect 5246 37223 5260 37275
rect 5312 37223 5326 37275
rect 5378 37223 5392 37275
rect 5444 37223 5447 37275
rect 4489 37211 5330 37223
rect 5364 37211 5447 37223
rect 4489 37159 4666 37211
rect 4718 37159 4732 37211
rect 4784 37159 4798 37211
rect 4850 37159 4864 37211
rect 4916 37159 4930 37211
rect 4982 37159 4996 37211
rect 5048 37159 5062 37211
rect 5114 37159 5128 37211
rect 5180 37159 5194 37211
rect 5246 37159 5260 37211
rect 5312 37159 5326 37211
rect 5378 37159 5392 37211
rect 5444 37159 5447 37211
rect 4489 37147 5330 37159
rect 5364 37147 5447 37159
rect 4489 37095 4666 37147
rect 4718 37095 4732 37147
rect 4784 37095 4798 37147
rect 4850 37095 4864 37147
rect 4916 37095 4930 37147
rect 4982 37095 4996 37147
rect 5048 37095 5062 37147
rect 5114 37095 5128 37147
rect 5180 37095 5194 37147
rect 5246 37095 5260 37147
rect 5312 37095 5326 37147
rect 5378 37095 5392 37147
rect 5444 37095 5447 37147
rect 4489 37094 5447 37095
rect 4489 37083 5330 37094
rect 5364 37083 5447 37094
rect 4489 37031 4666 37083
rect 4718 37031 4732 37083
rect 4784 37031 4798 37083
rect 4850 37031 4864 37083
rect 4916 37031 4930 37083
rect 4982 37031 4996 37083
rect 5048 37031 5062 37083
rect 5114 37031 5128 37083
rect 5180 37031 5194 37083
rect 5246 37031 5260 37083
rect 5312 37031 5326 37083
rect 5378 37031 5392 37083
rect 5444 37031 5447 37083
rect 4489 37022 5447 37031
rect 4489 37019 5330 37022
rect 5364 37019 5447 37022
rect 4489 36967 4666 37019
rect 4718 36967 4732 37019
rect 4784 36967 4798 37019
rect 4850 36967 4864 37019
rect 4916 36967 4930 37019
rect 4982 36967 4996 37019
rect 5048 36967 5062 37019
rect 5114 36967 5128 37019
rect 5180 36967 5194 37019
rect 5246 36967 5260 37019
rect 5312 36967 5326 37019
rect 5378 36967 5392 37019
rect 5444 36967 5447 37019
rect 4489 36955 5447 36967
rect 4489 36903 4666 36955
rect 4718 36903 4732 36955
rect 4784 36903 4798 36955
rect 4850 36903 4864 36955
rect 4916 36903 4930 36955
rect 4982 36903 4996 36955
rect 5048 36903 5062 36955
rect 5114 36903 5128 36955
rect 5180 36903 5194 36955
rect 5246 36903 5260 36955
rect 5312 36903 5326 36955
rect 5378 36903 5392 36955
rect 5444 36903 5447 36955
rect 4489 36891 5447 36903
rect 4489 36839 4666 36891
rect 4718 36839 4732 36891
rect 4784 36839 4798 36891
rect 4850 36839 4864 36891
rect 4916 36839 4930 36891
rect 4982 36839 4996 36891
rect 5048 36839 5062 36891
rect 5114 36839 5128 36891
rect 5180 36839 5194 36891
rect 5246 36839 5260 36891
rect 5312 36839 5326 36891
rect 5378 36839 5392 36891
rect 5444 36839 5447 36891
rect 4489 36827 5447 36839
rect 4489 36775 4666 36827
rect 4718 36775 4732 36827
rect 4784 36775 4798 36827
rect 4850 36775 4864 36827
rect 4916 36775 4930 36827
rect 4982 36775 4996 36827
rect 5048 36775 5062 36827
rect 5114 36775 5128 36827
rect 5180 36775 5194 36827
rect 5246 36775 5260 36827
rect 5312 36775 5326 36827
rect 5378 36775 5392 36827
rect 5444 36775 5447 36827
rect 4489 36772 5330 36775
rect 5364 36772 5447 36775
rect 4489 36763 5447 36772
rect 4489 36711 4666 36763
rect 4718 36711 4732 36763
rect 4784 36711 4798 36763
rect 4850 36711 4864 36763
rect 4916 36711 4930 36763
rect 4982 36711 4996 36763
rect 5048 36711 5062 36763
rect 5114 36711 5128 36763
rect 5180 36711 5194 36763
rect 5246 36711 5260 36763
rect 5312 36711 5326 36763
rect 5378 36711 5392 36763
rect 5444 36711 5447 36763
rect 4489 36700 5330 36711
rect 5364 36700 5447 36711
rect 4489 36699 5447 36700
rect 4489 36647 4666 36699
rect 4718 36647 4732 36699
rect 4784 36647 4798 36699
rect 4850 36647 4864 36699
rect 4916 36647 4930 36699
rect 4982 36647 4996 36699
rect 5048 36647 5062 36699
rect 5114 36647 5128 36699
rect 5180 36647 5194 36699
rect 5246 36647 5260 36699
rect 5312 36647 5326 36699
rect 5378 36647 5392 36699
rect 5444 36647 5447 36699
rect 4489 36635 5330 36647
rect 5364 36635 5447 36647
rect 4489 36583 4666 36635
rect 4718 36583 4732 36635
rect 4784 36583 4798 36635
rect 4850 36583 4864 36635
rect 4916 36583 4930 36635
rect 4982 36583 4996 36635
rect 5048 36583 5062 36635
rect 5114 36583 5128 36635
rect 5180 36583 5194 36635
rect 5246 36583 5260 36635
rect 5312 36583 5326 36635
rect 5378 36583 5392 36635
rect 5444 36583 5447 36635
rect 4489 36571 5330 36583
rect 5364 36571 5447 36583
rect 4489 36519 4666 36571
rect 4718 36519 4732 36571
rect 4784 36519 4798 36571
rect 4850 36519 4864 36571
rect 4916 36519 4930 36571
rect 4982 36519 4996 36571
rect 5048 36519 5062 36571
rect 5114 36519 5128 36571
rect 5180 36519 5194 36571
rect 5246 36519 5260 36571
rect 5312 36519 5326 36571
rect 5378 36519 5392 36571
rect 5444 36519 5447 36571
rect 4489 36518 5447 36519
rect 4489 36507 5330 36518
rect 5364 36507 5447 36518
rect 4489 36455 4666 36507
rect 4718 36455 4732 36507
rect 4784 36455 4798 36507
rect 4850 36455 4864 36507
rect 4916 36455 4930 36507
rect 4982 36455 4996 36507
rect 5048 36455 5062 36507
rect 5114 36455 5128 36507
rect 5180 36455 5194 36507
rect 5246 36455 5260 36507
rect 5312 36455 5326 36507
rect 5378 36455 5392 36507
rect 5444 36455 5447 36507
rect 4489 36446 5447 36455
rect 4489 36443 5330 36446
rect 5364 36443 5447 36446
rect 4489 36391 4666 36443
rect 4718 36391 4732 36443
rect 4784 36391 4798 36443
rect 4850 36391 4864 36443
rect 4916 36391 4930 36443
rect 4982 36391 4996 36443
rect 5048 36391 5062 36443
rect 5114 36391 5128 36443
rect 5180 36391 5194 36443
rect 5246 36391 5260 36443
rect 5312 36391 5326 36443
rect 5378 36391 5392 36443
rect 5444 36391 5447 36443
rect 4489 36379 5447 36391
rect 4489 36327 4666 36379
rect 4718 36327 4732 36379
rect 4784 36327 4798 36379
rect 4850 36327 4864 36379
rect 4916 36327 4930 36379
rect 4982 36327 4996 36379
rect 5048 36327 5062 36379
rect 5114 36327 5128 36379
rect 5180 36327 5194 36379
rect 5246 36327 5260 36379
rect 5312 36327 5326 36379
rect 5378 36327 5392 36379
rect 5444 36327 5447 36379
rect 4489 36315 5447 36327
rect 4489 36263 4666 36315
rect 4718 36263 4732 36315
rect 4784 36263 4798 36315
rect 4850 36263 4864 36315
rect 4916 36263 4930 36315
rect 4982 36263 4996 36315
rect 5048 36263 5062 36315
rect 5114 36263 5128 36315
rect 5180 36263 5194 36315
rect 5246 36263 5260 36315
rect 5312 36263 5326 36315
rect 5378 36263 5392 36315
rect 5444 36263 5447 36315
rect 4489 36251 5447 36263
rect 4489 36199 4666 36251
rect 4718 36199 4732 36251
rect 4784 36199 4798 36251
rect 4850 36199 4864 36251
rect 4916 36199 4930 36251
rect 4982 36199 4996 36251
rect 5048 36199 5062 36251
rect 5114 36199 5128 36251
rect 5180 36199 5194 36251
rect 5246 36199 5260 36251
rect 5312 36199 5326 36251
rect 5378 36199 5392 36251
rect 5444 36199 5447 36251
rect 4489 36196 5330 36199
rect 5364 36196 5447 36199
rect 4489 36187 5447 36196
rect 4489 36135 4666 36187
rect 4718 36135 4732 36187
rect 4784 36135 4798 36187
rect 4850 36135 4864 36187
rect 4916 36135 4930 36187
rect 4982 36135 4996 36187
rect 5048 36135 5062 36187
rect 5114 36135 5128 36187
rect 5180 36135 5194 36187
rect 5246 36135 5260 36187
rect 5312 36135 5326 36187
rect 5378 36135 5392 36187
rect 5444 36135 5447 36187
rect 4489 36124 5330 36135
rect 5364 36124 5447 36135
rect 4489 36123 5447 36124
rect 4489 36071 4666 36123
rect 4718 36071 4732 36123
rect 4784 36071 4798 36123
rect 4850 36071 4864 36123
rect 4916 36071 4930 36123
rect 4982 36071 4996 36123
rect 5048 36071 5062 36123
rect 5114 36071 5128 36123
rect 5180 36071 5194 36123
rect 5246 36071 5260 36123
rect 5312 36071 5326 36123
rect 5378 36071 5392 36123
rect 5444 36071 5447 36123
rect 4489 36059 5330 36071
rect 5364 36059 5447 36071
rect 4489 36007 4666 36059
rect 4718 36007 4732 36059
rect 4784 36007 4798 36059
rect 4850 36007 4864 36059
rect 4916 36007 4930 36059
rect 4982 36007 4996 36059
rect 5048 36007 5062 36059
rect 5114 36007 5128 36059
rect 5180 36007 5194 36059
rect 5246 36007 5260 36059
rect 5312 36007 5326 36059
rect 5378 36007 5392 36059
rect 5444 36007 5447 36059
rect 4489 35995 5330 36007
rect 5364 35995 5447 36007
rect 4489 35943 4666 35995
rect 4718 35943 4732 35995
rect 4784 35943 4798 35995
rect 4850 35943 4864 35995
rect 4916 35943 4930 35995
rect 4982 35943 4996 35995
rect 5048 35943 5062 35995
rect 5114 35943 5128 35995
rect 5180 35943 5194 35995
rect 5246 35943 5260 35995
rect 5312 35943 5326 35995
rect 5378 35943 5392 35995
rect 5444 35943 5447 35995
rect 4489 35942 5447 35943
rect 4489 35931 5330 35942
rect 5364 35931 5447 35942
rect 4489 35879 4666 35931
rect 4718 35879 4732 35931
rect 4784 35879 4798 35931
rect 4850 35879 4864 35931
rect 4916 35879 4930 35931
rect 4982 35879 4996 35931
rect 5048 35879 5062 35931
rect 5114 35879 5128 35931
rect 5180 35879 5194 35931
rect 5246 35879 5260 35931
rect 5312 35879 5326 35931
rect 5378 35879 5392 35931
rect 5444 35879 5447 35931
rect 4489 35870 5447 35879
rect 4489 35867 5330 35870
rect 5364 35867 5447 35870
rect 4489 35815 4666 35867
rect 4718 35815 4732 35867
rect 4784 35815 4798 35867
rect 4850 35815 4864 35867
rect 4916 35815 4930 35867
rect 4982 35815 4996 35867
rect 5048 35815 5062 35867
rect 5114 35815 5128 35867
rect 5180 35815 5194 35867
rect 5246 35815 5260 35867
rect 5312 35815 5326 35867
rect 5378 35815 5392 35867
rect 5444 35815 5447 35867
rect 4489 35803 5447 35815
rect 4489 35751 4666 35803
rect 4718 35751 4732 35803
rect 4784 35751 4798 35803
rect 4850 35751 4864 35803
rect 4916 35751 4930 35803
rect 4982 35751 4996 35803
rect 5048 35751 5062 35803
rect 5114 35751 5128 35803
rect 5180 35751 5194 35803
rect 5246 35751 5260 35803
rect 5312 35751 5326 35803
rect 5378 35751 5392 35803
rect 5444 35751 5447 35803
rect 4489 35739 5447 35751
rect 4489 35687 4666 35739
rect 4718 35687 4732 35739
rect 4784 35687 4798 35739
rect 4850 35687 4864 35739
rect 4916 35687 4930 35739
rect 4982 35687 4996 35739
rect 5048 35687 5062 35739
rect 5114 35687 5128 35739
rect 5180 35687 5194 35739
rect 5246 35687 5260 35739
rect 5312 35687 5326 35739
rect 5378 35687 5392 35739
rect 5444 35687 5447 35739
rect 4489 35675 5447 35687
rect 3208 35647 3217 35649
rect 3165 35643 3217 35647
rect 3165 35579 3174 35591
rect 3208 35579 3217 35591
rect 3165 35521 3174 35527
rect 3076 35456 3082 35490
rect 3116 35456 3122 35490
rect 3076 35418 3122 35456
rect 3076 35384 3082 35418
rect 3116 35384 3122 35418
rect 3076 35346 3122 35384
rect 3076 35312 3082 35346
rect 3116 35312 3122 35346
rect 3076 35274 3122 35312
rect 3076 35240 3082 35274
rect 3116 35240 3122 35274
rect 3076 35202 3122 35240
rect 3076 35168 3082 35202
rect 3116 35168 3122 35202
rect 3076 35130 3122 35168
rect 3076 35096 3082 35130
rect 3116 35096 3122 35130
rect 3076 35058 3122 35096
rect 3076 35024 3082 35058
rect 3116 35024 3122 35058
rect 3076 34986 3122 35024
rect 3076 34952 3082 34986
rect 3116 34952 3122 34986
rect 3076 34914 3122 34952
rect 3076 34880 3082 34914
rect 3116 34880 3122 34914
rect 3076 34842 3122 34880
rect 3076 34808 3082 34842
rect 3116 34808 3122 34842
rect 3076 34770 3122 34808
rect 3076 34736 3082 34770
rect 3116 34736 3122 34770
rect 3076 34698 3122 34736
rect 3076 34664 3082 34698
rect 3116 34664 3122 34698
rect 3076 34626 3122 34664
rect 3076 34592 3082 34626
rect 3116 34592 3122 34626
rect 3076 34554 3122 34592
rect 3076 34520 3082 34554
rect 3116 34520 3122 34554
rect 3076 34482 3122 34520
rect 3076 34448 3082 34482
rect 3116 34448 3122 34482
rect 3076 34410 3122 34448
rect 3076 34376 3082 34410
rect 3116 34376 3122 34410
rect 3076 34338 3122 34376
rect 3076 34304 3082 34338
rect 3116 34304 3122 34338
rect 3076 34266 3122 34304
rect 3076 34232 3082 34266
rect 3116 34232 3122 34266
rect 3076 34194 3122 34232
rect 3076 34160 3082 34194
rect 3116 34160 3122 34194
rect 3076 34122 3122 34160
rect 3076 34088 3082 34122
rect 3116 34088 3122 34122
rect 3076 34050 3122 34088
rect 3076 34016 3082 34050
rect 3116 34016 3122 34050
rect 3076 33978 3122 34016
rect 3076 33944 3082 33978
rect 3116 33944 3122 33978
rect 3076 33906 3122 33944
rect 3076 33872 3082 33906
rect 3116 33872 3122 33906
rect 3076 33834 3122 33872
rect 3076 33800 3082 33834
rect 3116 33800 3122 33834
rect 3076 33762 3122 33800
rect 3076 33728 3082 33762
rect 3116 33728 3122 33762
rect 3076 33690 3122 33728
rect 3076 33656 3082 33690
rect 3116 33656 3122 33690
rect 3076 33618 3122 33656
rect 3076 33584 3082 33618
rect 3116 33584 3122 33618
rect 3076 33546 3122 33584
rect 3076 33512 3082 33546
rect 3116 33512 3122 33546
rect 3076 33474 3122 33512
rect 3076 33440 3082 33474
rect 3116 33440 3122 33474
rect 3076 33402 3122 33440
rect 3076 33368 3082 33402
rect 3116 33368 3122 33402
rect 3076 33330 3122 33368
rect 3076 33296 3082 33330
rect 3116 33296 3122 33330
rect 3076 33258 3122 33296
rect 3076 33224 3082 33258
rect 3116 33224 3122 33258
rect 3076 33186 3122 33224
rect 3076 33152 3082 33186
rect 3116 33152 3122 33186
rect 3076 33114 3122 33152
rect 3076 33080 3082 33114
rect 3116 33080 3122 33114
rect 3076 33042 3122 33080
rect 3076 33008 3082 33042
rect 3116 33008 3122 33042
rect 3076 32970 3122 33008
rect 3076 32936 3082 32970
rect 3116 32936 3122 32970
rect 3076 32898 3122 32936
rect 3076 32864 3082 32898
rect 3116 32864 3122 32898
rect 3076 32826 3122 32864
rect 3076 32792 3082 32826
rect 3116 32792 3122 32826
rect 3076 32754 3122 32792
rect 3076 32720 3082 32754
rect 3116 32720 3122 32754
rect 3076 32682 3122 32720
rect 3076 32648 3082 32682
rect 3116 32648 3122 32682
rect 3076 32610 3122 32648
rect 3076 32576 3082 32610
rect 3116 32576 3122 32610
rect 3076 32538 3122 32576
rect 3076 32504 3082 32538
rect 3116 32504 3122 32538
rect 3076 32466 3122 32504
rect 3076 32432 3082 32466
rect 3116 32432 3122 32466
rect 3076 32394 3122 32432
rect 3076 32360 3082 32394
rect 3116 32360 3122 32394
rect 3076 32322 3122 32360
rect 3076 32288 3082 32322
rect 3116 32288 3122 32322
rect 3076 32250 3122 32288
rect 3076 32216 3082 32250
rect 3116 32216 3122 32250
rect 3076 32178 3122 32216
rect 3076 32144 3082 32178
rect 3116 32144 3122 32178
rect 3076 32106 3122 32144
rect 3076 32072 3082 32106
rect 3116 32072 3122 32106
rect 3076 32034 3122 32072
rect 3076 32000 3082 32034
rect 3116 32000 3122 32034
rect 3076 31962 3122 32000
rect 3076 31928 3082 31962
rect 3116 31928 3122 31962
rect 3076 31890 3122 31928
rect 3076 31856 3082 31890
rect 3116 31856 3122 31890
rect 3076 31818 3122 31856
rect 3076 31784 3082 31818
rect 3116 31784 3122 31818
rect 3076 31746 3122 31784
rect 3076 31712 3082 31746
rect 3116 31712 3122 31746
rect 3076 31674 3122 31712
rect 3076 31640 3082 31674
rect 3116 31640 3122 31674
rect 3076 31602 3122 31640
rect 3076 31568 3082 31602
rect 3116 31568 3122 31602
rect 3076 31530 3122 31568
rect 3076 31496 3082 31530
rect 3116 31496 3122 31530
rect 3076 31458 3122 31496
rect 3076 31424 3082 31458
rect 3116 31424 3122 31458
rect 3076 31386 3122 31424
rect 3076 31352 3082 31386
rect 3116 31352 3122 31386
rect 3076 31314 3122 31352
rect 3076 31280 3082 31314
rect 3116 31280 3122 31314
rect 3076 31242 3122 31280
rect 3076 31208 3082 31242
rect 3116 31208 3122 31242
rect 3076 31170 3122 31208
rect 3076 31136 3082 31170
rect 3116 31136 3122 31170
rect 3076 31098 3122 31136
rect 3076 31064 3082 31098
rect 3116 31064 3122 31098
rect 3076 31026 3122 31064
rect 3076 30992 3082 31026
rect 3116 30992 3122 31026
rect 3076 30954 3122 30992
rect 3076 30920 3082 30954
rect 3116 30920 3122 30954
rect 3076 30882 3122 30920
rect 3076 30848 3082 30882
rect 3116 30848 3122 30882
rect 3076 30810 3122 30848
rect 3076 30776 3082 30810
rect 3116 30776 3122 30810
rect 3076 30738 3122 30776
rect 3076 30704 3082 30738
rect 3116 30704 3122 30738
rect 3076 30666 3122 30704
rect 3076 30632 3082 30666
rect 3116 30632 3122 30666
rect 3076 30594 3122 30632
rect 3076 30560 3082 30594
rect 3116 30560 3122 30594
rect 3076 30522 3122 30560
rect 3076 30488 3082 30522
rect 3116 30488 3122 30522
rect 3076 30450 3122 30488
rect 3076 30416 3082 30450
rect 3116 30416 3122 30450
rect 3168 35503 3174 35521
rect 3208 35521 3217 35527
rect 4489 35623 4666 35675
rect 4718 35623 4732 35675
rect 4784 35623 4798 35675
rect 4850 35623 4864 35675
rect 4916 35623 4930 35675
rect 4982 35623 4996 35675
rect 5048 35623 5062 35675
rect 5114 35623 5128 35675
rect 5180 35623 5194 35675
rect 5246 35623 5260 35675
rect 5312 35623 5326 35675
rect 5378 35623 5392 35675
rect 5444 35623 5447 35675
rect 4489 35620 5330 35623
rect 5364 35620 5447 35623
rect 4489 35611 5447 35620
rect 4489 35559 4666 35611
rect 4718 35559 4732 35611
rect 4784 35559 4798 35611
rect 4850 35559 4864 35611
rect 4916 35559 4930 35611
rect 4982 35559 4996 35611
rect 5048 35559 5062 35611
rect 5114 35559 5128 35611
rect 5180 35559 5194 35611
rect 5246 35559 5260 35611
rect 5312 35559 5326 35611
rect 5378 35559 5392 35611
rect 5444 35559 5447 35611
rect 4489 35548 5330 35559
rect 5364 35548 5447 35559
rect 4489 35547 5447 35548
rect 3208 35503 3214 35521
rect 3168 35465 3214 35503
rect 3168 35431 3174 35465
rect 3208 35431 3214 35465
rect 3168 35393 3214 35431
rect 3168 35359 3174 35393
rect 3208 35359 3214 35393
rect 3168 35321 3214 35359
rect 3168 35287 3174 35321
rect 3208 35287 3214 35321
rect 3168 35249 3214 35287
rect 3168 35215 3174 35249
rect 3208 35215 3214 35249
rect 3168 35177 3214 35215
rect 3168 35143 3174 35177
rect 3208 35143 3214 35177
rect 3168 35105 3214 35143
rect 3168 35071 3174 35105
rect 3208 35071 3214 35105
rect 3168 35033 3214 35071
rect 3168 34999 3174 35033
rect 3208 34999 3214 35033
rect 3168 34961 3214 34999
rect 3168 34927 3174 34961
rect 3208 34927 3214 34961
rect 3168 34889 3214 34927
rect 3168 34855 3174 34889
rect 3208 34855 3214 34889
rect 3168 34817 3214 34855
rect 3168 34783 3174 34817
rect 3208 34783 3214 34817
rect 3168 34745 3214 34783
rect 3168 34711 3174 34745
rect 3208 34711 3214 34745
rect 3168 34673 3214 34711
rect 3168 34639 3174 34673
rect 3208 34639 3214 34673
rect 3168 34601 3214 34639
rect 3168 34567 3174 34601
rect 3208 34567 3214 34601
rect 3168 34529 3214 34567
rect 3168 34495 3174 34529
rect 3208 34495 3214 34529
rect 3168 34457 3214 34495
rect 3168 34423 3174 34457
rect 3208 34423 3214 34457
rect 3168 34385 3214 34423
rect 3168 34351 3174 34385
rect 3208 34351 3214 34385
rect 3168 34313 3214 34351
rect 3168 34279 3174 34313
rect 3208 34279 3214 34313
rect 3168 34241 3214 34279
rect 3168 34207 3174 34241
rect 3208 34207 3214 34241
rect 3168 34169 3214 34207
rect 3168 34135 3174 34169
rect 3208 34135 3214 34169
rect 3168 34097 3214 34135
rect 3168 34063 3174 34097
rect 3208 34063 3214 34097
rect 3168 34025 3214 34063
rect 3168 33991 3174 34025
rect 3208 33991 3214 34025
rect 3168 33953 3214 33991
rect 3168 33919 3174 33953
rect 3208 33919 3214 33953
rect 3168 33881 3214 33919
rect 3168 33847 3174 33881
rect 3208 33847 3214 33881
rect 3168 33809 3214 33847
rect 3168 33775 3174 33809
rect 3208 33775 3214 33809
rect 3168 33737 3214 33775
rect 3168 33703 3174 33737
rect 3208 33703 3214 33737
rect 3168 33665 3214 33703
rect 3168 33631 3174 33665
rect 3208 33631 3214 33665
rect 3168 33593 3214 33631
rect 3168 33559 3174 33593
rect 3208 33559 3214 33593
rect 3168 33521 3214 33559
rect 3168 33487 3174 33521
rect 3208 33487 3214 33521
rect 3168 33449 3214 33487
rect 3168 33415 3174 33449
rect 3208 33415 3214 33449
rect 3168 33377 3214 33415
rect 3168 33343 3174 33377
rect 3208 33343 3214 33377
rect 3168 33305 3214 33343
rect 3168 33271 3174 33305
rect 3208 33271 3214 33305
rect 3168 33233 3214 33271
rect 3168 33199 3174 33233
rect 3208 33199 3214 33233
rect 3168 33161 3214 33199
rect 3168 33127 3174 33161
rect 3208 33127 3214 33161
rect 3168 33089 3214 33127
rect 3168 33055 3174 33089
rect 3208 33055 3214 33089
rect 3168 33017 3214 33055
rect 3168 32983 3174 33017
rect 3208 32983 3214 33017
rect 3168 32945 3214 32983
rect 3168 32911 3174 32945
rect 3208 32911 3214 32945
rect 3168 32873 3214 32911
rect 3168 32839 3174 32873
rect 3208 32839 3214 32873
rect 3168 32801 3214 32839
rect 3168 32767 3174 32801
rect 3208 32767 3214 32801
rect 3168 32729 3214 32767
rect 3168 32695 3174 32729
rect 3208 32695 3214 32729
rect 3168 32657 3214 32695
rect 3168 32623 3174 32657
rect 3208 32623 3214 32657
rect 3168 32585 3214 32623
rect 3168 32551 3174 32585
rect 3208 32551 3214 32585
rect 3168 32513 3214 32551
rect 3168 32479 3174 32513
rect 3208 32479 3214 32513
rect 3168 32441 3214 32479
rect 3168 32407 3174 32441
rect 3208 32407 3214 32441
rect 3168 32369 3214 32407
rect 3168 32335 3174 32369
rect 3208 32335 3214 32369
rect 3168 32296 3214 32335
rect 3168 32262 3174 32296
rect 3208 32262 3214 32296
rect 3168 32223 3214 32262
rect 3168 32189 3174 32223
rect 3208 32189 3214 32223
rect 3168 32150 3214 32189
rect 3168 32116 3174 32150
rect 3208 32116 3214 32150
rect 3168 32077 3214 32116
rect 3168 32043 3174 32077
rect 3208 32043 3214 32077
rect 3168 32004 3214 32043
rect 3168 31970 3174 32004
rect 3208 31970 3214 32004
rect 3168 31931 3214 31970
rect 3168 31897 3174 31931
rect 3208 31897 3214 31931
rect 3168 31858 3214 31897
rect 3168 31824 3174 31858
rect 3208 31824 3214 31858
rect 3168 31785 3214 31824
rect 3168 31751 3174 31785
rect 3208 31751 3214 31785
rect 3168 31712 3214 31751
rect 3168 31678 3174 31712
rect 3208 31678 3214 31712
rect 3168 31639 3214 31678
rect 3168 31605 3174 31639
rect 3208 31605 3214 31639
rect 3168 31566 3214 31605
rect 3168 31532 3174 31566
rect 3208 31532 3214 31566
rect 3168 31493 3214 31532
rect 3168 31459 3174 31493
rect 3208 31459 3214 31493
rect 3168 31420 3214 31459
rect 3168 31386 3174 31420
rect 3208 31386 3214 31420
rect 3168 31347 3214 31386
rect 3168 31313 3174 31347
rect 3208 31313 3214 31347
rect 3168 31274 3214 31313
rect 3168 31240 3174 31274
rect 3208 31240 3214 31274
rect 3168 31201 3214 31240
rect 3168 31167 3174 31201
rect 3208 31167 3214 31201
rect 3168 31128 3214 31167
rect 3168 31094 3174 31128
rect 3208 31094 3214 31128
rect 3168 31055 3214 31094
rect 3168 31021 3174 31055
rect 3208 31021 3214 31055
rect 3168 30982 3214 31021
rect 3168 30948 3174 30982
rect 3208 30948 3214 30982
rect 3168 30909 3214 30948
rect 3168 30875 3174 30909
rect 3208 30875 3214 30909
rect 3168 30836 3214 30875
rect 3168 30802 3174 30836
rect 3208 30802 3214 30836
rect 3168 30763 3214 30802
rect 3168 30729 3174 30763
rect 3208 30729 3214 30763
rect 3168 30690 3214 30729
rect 3168 30656 3174 30690
rect 3208 30656 3214 30690
rect 3168 30617 3214 30656
rect 3168 30583 3174 30617
rect 3208 30583 3214 30617
rect 3168 30544 3214 30583
rect 3168 30510 3174 30544
rect 3208 30510 3214 30544
rect 3168 30471 3214 30510
rect 3168 30437 3174 30471
rect 3208 30437 3214 30471
rect 3168 30425 3214 30437
rect 4489 35495 4666 35547
rect 4718 35495 4732 35547
rect 4784 35495 4798 35547
rect 4850 35495 4864 35547
rect 4916 35495 4930 35547
rect 4982 35495 4996 35547
rect 5048 35495 5062 35547
rect 5114 35495 5128 35547
rect 5180 35495 5194 35547
rect 5246 35495 5260 35547
rect 5312 35495 5326 35547
rect 5378 35495 5392 35547
rect 5444 35495 5447 35547
rect 4489 35483 5330 35495
rect 5364 35483 5447 35495
rect 4489 35431 4666 35483
rect 4718 35431 4732 35483
rect 4784 35431 4798 35483
rect 4850 35431 4864 35483
rect 4916 35431 4930 35483
rect 4982 35431 4996 35483
rect 5048 35431 5062 35483
rect 5114 35431 5128 35483
rect 5180 35431 5194 35483
rect 5246 35431 5260 35483
rect 5312 35431 5326 35483
rect 5378 35431 5392 35483
rect 5444 35431 5447 35483
rect 4489 35419 5330 35431
rect 5364 35419 5447 35431
rect 4489 35367 4666 35419
rect 4718 35367 4732 35419
rect 4784 35367 4798 35419
rect 4850 35367 4864 35419
rect 4916 35367 4930 35419
rect 4982 35367 4996 35419
rect 5048 35367 5062 35419
rect 5114 35367 5128 35419
rect 5180 35367 5194 35419
rect 5246 35367 5260 35419
rect 5312 35367 5326 35419
rect 5378 35367 5392 35419
rect 5444 35367 5447 35419
rect 4489 35366 5447 35367
rect 4489 35355 5330 35366
rect 5364 35355 5447 35366
rect 4489 35303 4666 35355
rect 4718 35303 4732 35355
rect 4784 35303 4798 35355
rect 4850 35303 4864 35355
rect 4916 35303 4930 35355
rect 4982 35303 4996 35355
rect 5048 35303 5062 35355
rect 5114 35303 5128 35355
rect 5180 35303 5194 35355
rect 5246 35303 5260 35355
rect 5312 35303 5326 35355
rect 5378 35303 5392 35355
rect 5444 35303 5447 35355
rect 4489 35294 5447 35303
rect 4489 35291 5330 35294
rect 5364 35291 5447 35294
rect 4489 35239 4666 35291
rect 4718 35239 4732 35291
rect 4784 35239 4798 35291
rect 4850 35239 4864 35291
rect 4916 35239 4930 35291
rect 4982 35239 4996 35291
rect 5048 35239 5062 35291
rect 5114 35239 5128 35291
rect 5180 35239 5194 35291
rect 5246 35239 5260 35291
rect 5312 35239 5326 35291
rect 5378 35239 5392 35291
rect 5444 35239 5447 35291
rect 4489 35227 5447 35239
rect 4489 35175 4666 35227
rect 4718 35175 4732 35227
rect 4784 35175 4798 35227
rect 4850 35175 4864 35227
rect 4916 35175 4930 35227
rect 4982 35175 4996 35227
rect 5048 35175 5062 35227
rect 5114 35175 5128 35227
rect 5180 35175 5194 35227
rect 5246 35175 5260 35227
rect 5312 35175 5326 35227
rect 5378 35175 5392 35227
rect 5444 35175 5447 35227
rect 4489 35163 5447 35175
rect 4489 35111 4666 35163
rect 4718 35111 4732 35163
rect 4784 35111 4798 35163
rect 4850 35111 4864 35163
rect 4916 35111 4930 35163
rect 4982 35111 4996 35163
rect 5048 35111 5062 35163
rect 5114 35111 5128 35163
rect 5180 35111 5194 35163
rect 5246 35111 5260 35163
rect 5312 35111 5326 35163
rect 5378 35111 5392 35163
rect 5444 35111 5447 35163
rect 4489 35099 5447 35111
rect 4489 35047 4666 35099
rect 4718 35047 4732 35099
rect 4784 35047 4798 35099
rect 4850 35047 4864 35099
rect 4916 35047 4930 35099
rect 4982 35047 4996 35099
rect 5048 35047 5062 35099
rect 5114 35047 5128 35099
rect 5180 35047 5194 35099
rect 5246 35047 5260 35099
rect 5312 35047 5326 35099
rect 5378 35047 5392 35099
rect 5444 35047 5447 35099
rect 4489 35042 5330 35047
rect 5364 35042 5447 35047
rect 4489 35035 5447 35042
rect 4489 34983 4666 35035
rect 4718 34983 4732 35035
rect 4784 34983 4798 35035
rect 4850 34983 4864 35035
rect 4916 34983 4930 35035
rect 4982 34983 4996 35035
rect 5048 34983 5062 35035
rect 5114 34983 5128 35035
rect 5180 34983 5194 35035
rect 5246 34983 5260 35035
rect 5312 34983 5326 35035
rect 5378 34983 5392 35035
rect 5444 34983 5447 35035
rect 4489 34971 5330 34983
rect 5364 34971 5447 34983
rect 4489 34919 4666 34971
rect 4718 34919 4732 34971
rect 4784 34919 4798 34971
rect 4850 34919 4864 34971
rect 4916 34919 4930 34971
rect 4982 34919 4996 34971
rect 5048 34919 5062 34971
rect 5114 34919 5128 34971
rect 5180 34919 5194 34971
rect 5246 34919 5260 34971
rect 5312 34919 5326 34971
rect 5378 34919 5392 34971
rect 5444 34919 5447 34971
rect 4489 34907 5330 34919
rect 5364 34907 5447 34919
rect 4489 34855 4666 34907
rect 4718 34855 4732 34907
rect 4784 34855 4798 34907
rect 4850 34855 4864 34907
rect 4916 34855 4930 34907
rect 4982 34855 4996 34907
rect 5048 34855 5062 34907
rect 5114 34855 5128 34907
rect 5180 34855 5194 34907
rect 5246 34855 5260 34907
rect 5312 34855 5326 34907
rect 5378 34855 5392 34907
rect 5444 34855 5447 34907
rect 4489 34843 5330 34855
rect 5364 34843 5447 34855
rect 4489 34791 4666 34843
rect 4718 34791 4732 34843
rect 4784 34791 4798 34843
rect 4850 34791 4864 34843
rect 4916 34791 4930 34843
rect 4982 34791 4996 34843
rect 5048 34791 5062 34843
rect 5114 34791 5128 34843
rect 5180 34791 5194 34843
rect 5246 34791 5260 34843
rect 5312 34791 5326 34843
rect 5378 34791 5392 34843
rect 5444 34791 5447 34843
rect 4489 34784 5447 34791
rect 4489 34779 5330 34784
rect 5364 34779 5447 34784
rect 4489 34727 4666 34779
rect 4718 34727 4732 34779
rect 4784 34727 4798 34779
rect 4850 34727 4864 34779
rect 4916 34727 4930 34779
rect 4982 34727 4996 34779
rect 5048 34727 5062 34779
rect 5114 34727 5128 34779
rect 5180 34727 5194 34779
rect 5246 34727 5260 34779
rect 5312 34727 5326 34779
rect 5378 34727 5392 34779
rect 5444 34727 5447 34779
rect 4489 34715 5447 34727
rect 4489 34663 4666 34715
rect 4718 34663 4732 34715
rect 4784 34663 4798 34715
rect 4850 34663 4864 34715
rect 4916 34663 4930 34715
rect 4982 34663 4996 34715
rect 5048 34663 5062 34715
rect 5114 34663 5128 34715
rect 5180 34663 5194 34715
rect 5246 34663 5260 34715
rect 5312 34663 5326 34715
rect 5378 34663 5392 34715
rect 5444 34663 5447 34715
rect 4489 34651 5447 34663
rect 4489 34599 4666 34651
rect 4718 34599 4732 34651
rect 4784 34599 4798 34651
rect 4850 34599 4864 34651
rect 4916 34599 4930 34651
rect 4982 34599 4996 34651
rect 5048 34599 5062 34651
rect 5114 34599 5128 34651
rect 5180 34599 5194 34651
rect 5246 34599 5260 34651
rect 5312 34599 5326 34651
rect 5378 34599 5392 34651
rect 5444 34599 5447 34651
rect 4489 34587 5447 34599
rect 4489 34535 4666 34587
rect 4718 34535 4732 34587
rect 4784 34535 4798 34587
rect 4850 34535 4864 34587
rect 4916 34535 4930 34587
rect 4982 34535 4996 34587
rect 5048 34535 5062 34587
rect 5114 34535 5128 34587
rect 5180 34535 5194 34587
rect 5246 34535 5260 34587
rect 5312 34535 5326 34587
rect 5378 34535 5392 34587
rect 5444 34535 5447 34587
rect 4489 34531 5330 34535
rect 5364 34531 5447 34535
rect 4489 34523 5447 34531
rect 4489 34471 4666 34523
rect 4718 34471 4732 34523
rect 4784 34471 4798 34523
rect 4850 34471 4864 34523
rect 4916 34471 4930 34523
rect 4982 34471 4996 34523
rect 5048 34471 5062 34523
rect 5114 34471 5128 34523
rect 5180 34471 5194 34523
rect 5246 34471 5260 34523
rect 5312 34471 5326 34523
rect 5378 34471 5392 34523
rect 5444 34471 5447 34523
rect 4489 34459 5330 34471
rect 5364 34459 5447 34471
rect 4489 34407 4666 34459
rect 4718 34407 4732 34459
rect 4784 34407 4798 34459
rect 4850 34407 4864 34459
rect 4916 34407 4930 34459
rect 4982 34407 4996 34459
rect 5048 34407 5062 34459
rect 5114 34407 5128 34459
rect 5180 34407 5194 34459
rect 5246 34407 5260 34459
rect 5312 34407 5326 34459
rect 5378 34407 5392 34459
rect 5444 34407 5447 34459
rect 4489 34395 5330 34407
rect 5364 34395 5447 34407
rect 4489 34343 4666 34395
rect 4718 34343 4732 34395
rect 4784 34343 4798 34395
rect 4850 34343 4864 34395
rect 4916 34343 4930 34395
rect 4982 34343 4996 34395
rect 5048 34343 5062 34395
rect 5114 34343 5128 34395
rect 5180 34343 5194 34395
rect 5246 34343 5260 34395
rect 5312 34343 5326 34395
rect 5378 34343 5392 34395
rect 5444 34343 5447 34395
rect 4489 34331 5330 34343
rect 5364 34331 5447 34343
rect 4489 34279 4666 34331
rect 4718 34279 4732 34331
rect 4784 34279 4798 34331
rect 4850 34279 4864 34331
rect 4916 34279 4930 34331
rect 4982 34279 4996 34331
rect 5048 34279 5062 34331
rect 5114 34279 5128 34331
rect 5180 34279 5194 34331
rect 5246 34279 5260 34331
rect 5312 34279 5326 34331
rect 5378 34279 5392 34331
rect 5444 34279 5447 34331
rect 4489 34273 5447 34279
rect 4489 34267 5330 34273
rect 5364 34267 5447 34273
rect 4489 34215 4666 34267
rect 4718 34215 4732 34267
rect 4784 34215 4798 34267
rect 4850 34215 4864 34267
rect 4916 34215 4930 34267
rect 4982 34215 4996 34267
rect 5048 34215 5062 34267
rect 5114 34215 5128 34267
rect 5180 34215 5194 34267
rect 5246 34215 5260 34267
rect 5312 34215 5326 34267
rect 5378 34215 5392 34267
rect 5444 34215 5447 34267
rect 4489 34203 5447 34215
rect 4489 34151 4666 34203
rect 4718 34151 4732 34203
rect 4784 34151 4798 34203
rect 4850 34151 4864 34203
rect 4916 34151 4930 34203
rect 4982 34151 4996 34203
rect 5048 34151 5062 34203
rect 5114 34151 5128 34203
rect 5180 34151 5194 34203
rect 5246 34151 5260 34203
rect 5312 34151 5326 34203
rect 5378 34151 5392 34203
rect 5444 34151 5447 34203
rect 4489 34139 5447 34151
rect 4489 34087 4666 34139
rect 4718 34087 4732 34139
rect 4784 34087 4798 34139
rect 4850 34087 4864 34139
rect 4916 34087 4930 34139
rect 4982 34087 4996 34139
rect 5048 34087 5062 34139
rect 5114 34087 5128 34139
rect 5180 34087 5194 34139
rect 5246 34087 5260 34139
rect 5312 34087 5326 34139
rect 5378 34087 5392 34139
rect 5444 34087 5447 34139
rect 4489 34075 5447 34087
rect 4489 34023 4666 34075
rect 4718 34023 4732 34075
rect 4784 34023 4798 34075
rect 4850 34023 4864 34075
rect 4916 34023 4930 34075
rect 4982 34023 4996 34075
rect 5048 34023 5062 34075
rect 5114 34023 5128 34075
rect 5180 34023 5194 34075
rect 5246 34023 5260 34075
rect 5312 34023 5326 34075
rect 5378 34023 5392 34075
rect 5444 34023 5447 34075
rect 4489 34020 5330 34023
rect 5364 34020 5447 34023
rect 4489 34011 5447 34020
rect 4489 33959 4666 34011
rect 4718 33959 4732 34011
rect 4784 33959 4798 34011
rect 4850 33959 4864 34011
rect 4916 33959 4930 34011
rect 4982 33959 4996 34011
rect 5048 33959 5062 34011
rect 5114 33959 5128 34011
rect 5180 33959 5194 34011
rect 5246 33959 5260 34011
rect 5312 33959 5326 34011
rect 5378 33959 5392 34011
rect 5444 33959 5447 34011
rect 4489 33947 5330 33959
rect 5364 33947 5447 33959
rect 4489 33895 4666 33947
rect 4718 33895 4732 33947
rect 4784 33895 4798 33947
rect 4850 33895 4864 33947
rect 4916 33895 4930 33947
rect 4982 33895 4996 33947
rect 5048 33895 5062 33947
rect 5114 33895 5128 33947
rect 5180 33895 5194 33947
rect 5246 33895 5260 33947
rect 5312 33895 5326 33947
rect 5378 33895 5392 33947
rect 5444 33895 5447 33947
rect 4489 33883 5330 33895
rect 5364 33883 5447 33895
rect 4489 33831 4666 33883
rect 4718 33831 4732 33883
rect 4784 33831 4798 33883
rect 4850 33831 4864 33883
rect 4916 33831 4930 33883
rect 4982 33831 4996 33883
rect 5048 33831 5062 33883
rect 5114 33831 5128 33883
rect 5180 33831 5194 33883
rect 5246 33831 5260 33883
rect 5312 33831 5326 33883
rect 5378 33831 5392 33883
rect 5444 33831 5447 33883
rect 4489 33819 5330 33831
rect 5364 33819 5447 33831
rect 4489 33767 4666 33819
rect 4718 33767 4732 33819
rect 4784 33767 4798 33819
rect 4850 33767 4864 33819
rect 4916 33767 4930 33819
rect 4982 33767 4996 33819
rect 5048 33767 5062 33819
rect 5114 33767 5128 33819
rect 5180 33767 5194 33819
rect 5246 33767 5260 33819
rect 5312 33767 5326 33819
rect 5378 33767 5392 33819
rect 5444 33767 5447 33819
rect 4489 33762 5447 33767
rect 4489 33755 5330 33762
rect 5364 33755 5447 33762
rect 4489 33703 4666 33755
rect 4718 33703 4732 33755
rect 4784 33703 4798 33755
rect 4850 33703 4864 33755
rect 4916 33703 4930 33755
rect 4982 33703 4996 33755
rect 5048 33703 5062 33755
rect 5114 33703 5128 33755
rect 5180 33703 5194 33755
rect 5246 33703 5260 33755
rect 5312 33703 5326 33755
rect 5378 33703 5392 33755
rect 5444 33703 5447 33755
rect 4489 33691 5447 33703
rect 4489 33639 4666 33691
rect 4718 33639 4732 33691
rect 4784 33639 4798 33691
rect 4850 33639 4864 33691
rect 4916 33639 4930 33691
rect 4982 33639 4996 33691
rect 5048 33639 5062 33691
rect 5114 33639 5128 33691
rect 5180 33639 5194 33691
rect 5246 33639 5260 33691
rect 5312 33639 5326 33691
rect 5378 33639 5392 33691
rect 5444 33639 5447 33691
rect 4489 33627 5447 33639
rect 4489 33575 4666 33627
rect 4718 33575 4732 33627
rect 4784 33575 4798 33627
rect 4850 33575 4864 33627
rect 4916 33575 4930 33627
rect 4982 33575 4996 33627
rect 5048 33575 5062 33627
rect 5114 33575 5128 33627
rect 5180 33575 5194 33627
rect 5246 33575 5260 33627
rect 5312 33575 5326 33627
rect 5378 33575 5392 33627
rect 5444 33575 5447 33627
rect 4489 33563 5447 33575
rect 4489 33511 4666 33563
rect 4718 33511 4732 33563
rect 4784 33511 4798 33563
rect 4850 33511 4864 33563
rect 4916 33511 4930 33563
rect 4982 33511 4996 33563
rect 5048 33511 5062 33563
rect 5114 33511 5128 33563
rect 5180 33511 5194 33563
rect 5246 33511 5260 33563
rect 5312 33511 5326 33563
rect 5378 33511 5392 33563
rect 5444 33511 5447 33563
rect 4489 33509 5330 33511
rect 5364 33509 5447 33511
rect 4489 33499 5447 33509
rect 4489 33447 4666 33499
rect 4718 33447 4732 33499
rect 4784 33447 4798 33499
rect 4850 33447 4864 33499
rect 4916 33447 4930 33499
rect 4982 33447 4996 33499
rect 5048 33447 5062 33499
rect 5114 33447 5128 33499
rect 5180 33447 5194 33499
rect 5246 33447 5260 33499
rect 5312 33447 5326 33499
rect 5378 33447 5392 33499
rect 5444 33447 5447 33499
rect 4489 33436 5330 33447
rect 5364 33436 5447 33447
rect 4489 33435 5447 33436
rect 4489 33383 4666 33435
rect 4718 33383 4732 33435
rect 4784 33383 4798 33435
rect 4850 33383 4864 33435
rect 4916 33383 4930 33435
rect 4982 33383 4996 33435
rect 5048 33383 5062 33435
rect 5114 33383 5128 33435
rect 5180 33383 5194 33435
rect 5246 33383 5260 33435
rect 5312 33383 5326 33435
rect 5378 33383 5392 33435
rect 5444 33383 5447 33435
rect 4489 33371 5330 33383
rect 5364 33371 5447 33383
rect 4489 33319 4666 33371
rect 4718 33319 4732 33371
rect 4784 33319 4798 33371
rect 4850 33319 4864 33371
rect 4916 33319 4930 33371
rect 4982 33319 4996 33371
rect 5048 33319 5062 33371
rect 5114 33319 5128 33371
rect 5180 33319 5194 33371
rect 5246 33319 5260 33371
rect 5312 33319 5326 33371
rect 5378 33319 5392 33371
rect 5444 33319 5447 33371
rect 4489 33307 5330 33319
rect 5364 33307 5447 33319
rect 4489 33255 4666 33307
rect 4718 33255 4732 33307
rect 4784 33255 4798 33307
rect 4850 33255 4864 33307
rect 4916 33255 4930 33307
rect 4982 33255 4996 33307
rect 5048 33255 5062 33307
rect 5114 33255 5128 33307
rect 5180 33255 5194 33307
rect 5246 33255 5260 33307
rect 5312 33255 5326 33307
rect 5378 33255 5392 33307
rect 5444 33255 5447 33307
rect 4489 33251 5447 33255
rect 4489 33243 5330 33251
rect 5364 33243 5447 33251
rect 4489 33191 4666 33243
rect 4718 33191 4732 33243
rect 4784 33191 4798 33243
rect 4850 33191 4864 33243
rect 4916 33191 4930 33243
rect 4982 33191 4996 33243
rect 5048 33191 5062 33243
rect 5114 33191 5128 33243
rect 5180 33191 5194 33243
rect 5246 33191 5260 33243
rect 5312 33191 5326 33243
rect 5378 33191 5392 33243
rect 5444 33191 5447 33243
rect 4489 33179 5447 33191
rect 4489 33127 4666 33179
rect 4718 33127 4732 33179
rect 4784 33127 4798 33179
rect 4850 33127 4864 33179
rect 4916 33127 4930 33179
rect 4982 33127 4996 33179
rect 5048 33127 5062 33179
rect 5114 33127 5128 33179
rect 5180 33127 5194 33179
rect 5246 33127 5260 33179
rect 5312 33127 5326 33179
rect 5378 33127 5392 33179
rect 5444 33127 5447 33179
rect 4489 33115 5447 33127
rect 4489 33063 4666 33115
rect 4718 33063 4732 33115
rect 4784 33063 4798 33115
rect 4850 33063 4864 33115
rect 4916 33063 4930 33115
rect 4982 33063 4996 33115
rect 5048 33063 5062 33115
rect 5114 33063 5128 33115
rect 5180 33063 5194 33115
rect 5246 33063 5260 33115
rect 5312 33063 5326 33115
rect 5378 33063 5392 33115
rect 5444 33063 5447 33115
rect 4489 33051 5447 33063
rect 4489 32999 4666 33051
rect 4718 32999 4732 33051
rect 4784 32999 4798 33051
rect 4850 32999 4864 33051
rect 4916 32999 4930 33051
rect 4982 32999 4996 33051
rect 5048 32999 5062 33051
rect 5114 32999 5128 33051
rect 5180 32999 5194 33051
rect 5246 32999 5260 33051
rect 5312 32999 5326 33051
rect 5378 32999 5392 33051
rect 5444 32999 5447 33051
rect 4489 32998 5330 32999
rect 5364 32998 5447 32999
rect 4489 32987 5447 32998
rect 4489 32935 4666 32987
rect 4718 32935 4732 32987
rect 4784 32935 4798 32987
rect 4850 32935 4864 32987
rect 4916 32935 4930 32987
rect 4982 32935 4996 32987
rect 5048 32935 5062 32987
rect 5114 32935 5128 32987
rect 5180 32935 5194 32987
rect 5246 32935 5260 32987
rect 5312 32935 5326 32987
rect 5378 32935 5392 32987
rect 5444 32935 5447 32987
rect 4489 32925 5330 32935
rect 5364 32925 5447 32935
rect 4489 32923 5447 32925
rect 4489 32871 4666 32923
rect 4718 32871 4732 32923
rect 4784 32871 4798 32923
rect 4850 32871 4864 32923
rect 4916 32871 4930 32923
rect 4982 32871 4996 32923
rect 5048 32871 5062 32923
rect 5114 32871 5128 32923
rect 5180 32871 5194 32923
rect 5246 32871 5260 32923
rect 5312 32871 5326 32923
rect 5378 32871 5392 32923
rect 5444 32871 5447 32923
rect 4489 32859 5330 32871
rect 5364 32859 5447 32871
rect 4489 32807 4666 32859
rect 4718 32807 4732 32859
rect 4784 32807 4798 32859
rect 4850 32807 4864 32859
rect 4916 32807 4930 32859
rect 4982 32807 4996 32859
rect 5048 32807 5062 32859
rect 5114 32807 5128 32859
rect 5180 32807 5194 32859
rect 5246 32807 5260 32859
rect 5312 32807 5326 32859
rect 5378 32807 5392 32859
rect 5444 32807 5447 32859
rect 4489 32795 5330 32807
rect 5364 32795 5447 32807
rect 4489 32743 4666 32795
rect 4718 32743 4732 32795
rect 4784 32743 4798 32795
rect 4850 32743 4864 32795
rect 4916 32743 4930 32795
rect 4982 32743 4996 32795
rect 5048 32743 5062 32795
rect 5114 32743 5128 32795
rect 5180 32743 5194 32795
rect 5246 32743 5260 32795
rect 5312 32743 5326 32795
rect 5378 32743 5392 32795
rect 5444 32743 5447 32795
rect 4489 32740 5447 32743
rect 4489 32730 5330 32740
rect 5364 32730 5447 32740
rect 4489 32678 4666 32730
rect 4718 32678 4732 32730
rect 4784 32678 4798 32730
rect 4850 32678 4864 32730
rect 4916 32678 4930 32730
rect 4982 32678 4996 32730
rect 5048 32678 5062 32730
rect 5114 32678 5128 32730
rect 5180 32678 5194 32730
rect 5246 32678 5260 32730
rect 5312 32678 5326 32730
rect 5378 32678 5392 32730
rect 5444 32678 5447 32730
rect 4489 32667 5447 32678
rect 4489 32665 5330 32667
rect 5364 32665 5447 32667
rect 4489 32613 4666 32665
rect 4718 32613 4732 32665
rect 4784 32613 4798 32665
rect 4850 32613 4864 32665
rect 4916 32613 4930 32665
rect 4982 32613 4996 32665
rect 5048 32613 5062 32665
rect 5114 32613 5128 32665
rect 5180 32613 5194 32665
rect 5246 32613 5260 32665
rect 5312 32613 5326 32665
rect 5378 32613 5392 32665
rect 5444 32613 5447 32665
rect 4489 32600 5447 32613
rect 4489 32548 4666 32600
rect 4718 32548 4732 32600
rect 4784 32548 4798 32600
rect 4850 32548 4864 32600
rect 4916 32548 4930 32600
rect 4982 32548 4996 32600
rect 5048 32548 5062 32600
rect 5114 32548 5128 32600
rect 5180 32548 5194 32600
rect 5246 32548 5260 32600
rect 5312 32548 5326 32600
rect 5378 32548 5392 32600
rect 5444 32548 5447 32600
rect 4489 32535 5447 32548
rect 4489 32483 4666 32535
rect 4718 32483 4732 32535
rect 4784 32483 4798 32535
rect 4850 32483 4864 32535
rect 4916 32483 4930 32535
rect 4982 32483 4996 32535
rect 5048 32483 5062 32535
rect 5114 32483 5128 32535
rect 5180 32483 5194 32535
rect 5246 32483 5260 32535
rect 5312 32483 5326 32535
rect 5378 32483 5392 32535
rect 5444 32483 5447 32535
rect 4489 32470 5447 32483
rect 4489 32418 4666 32470
rect 4718 32418 4732 32470
rect 4784 32418 4798 32470
rect 4850 32418 4864 32470
rect 4916 32418 4930 32470
rect 4982 32418 4996 32470
rect 5048 32418 5062 32470
rect 5114 32418 5128 32470
rect 5180 32418 5194 32470
rect 5246 32418 5260 32470
rect 5312 32418 5326 32470
rect 5378 32418 5392 32470
rect 5444 32418 5447 32470
rect 4489 32414 5330 32418
rect 5364 32414 5447 32418
rect 4489 32405 5447 32414
rect 4489 32353 4666 32405
rect 4718 32353 4732 32405
rect 4784 32353 4798 32405
rect 4850 32353 4864 32405
rect 4916 32353 4930 32405
rect 4982 32353 4996 32405
rect 5048 32353 5062 32405
rect 5114 32353 5128 32405
rect 5180 32353 5194 32405
rect 5246 32353 5260 32405
rect 5312 32353 5326 32405
rect 5378 32353 5392 32405
rect 5444 32353 5447 32405
rect 4489 32341 5330 32353
rect 5364 32341 5447 32353
rect 4489 32340 5447 32341
rect 4489 32288 4666 32340
rect 4718 32288 4732 32340
rect 4784 32288 4798 32340
rect 4850 32288 4864 32340
rect 4916 32288 4930 32340
rect 4982 32288 4996 32340
rect 5048 32288 5062 32340
rect 5114 32288 5128 32340
rect 5180 32288 5194 32340
rect 5246 32288 5260 32340
rect 5312 32288 5326 32340
rect 5378 32288 5392 32340
rect 5444 32288 5447 32340
rect 4489 32275 5330 32288
rect 5364 32275 5447 32288
rect 4489 32223 4666 32275
rect 4718 32223 4732 32275
rect 4784 32223 4798 32275
rect 4850 32223 4864 32275
rect 4916 32223 4930 32275
rect 4982 32223 4996 32275
rect 5048 32223 5062 32275
rect 5114 32223 5128 32275
rect 5180 32223 5194 32275
rect 5246 32223 5260 32275
rect 5312 32223 5326 32275
rect 5378 32223 5392 32275
rect 5444 32223 5447 32275
rect 4489 32210 5330 32223
rect 5364 32210 5447 32223
rect 4489 32158 4666 32210
rect 4718 32158 4732 32210
rect 4784 32158 4798 32210
rect 4850 32158 4864 32210
rect 4916 32158 4930 32210
rect 4982 32158 4996 32210
rect 5048 32158 5062 32210
rect 5114 32158 5128 32210
rect 5180 32158 5194 32210
rect 5246 32158 5260 32210
rect 5312 32158 5326 32210
rect 5378 32158 5392 32210
rect 5444 32158 5447 32210
rect 4489 32156 5447 32158
rect 4489 32145 5330 32156
rect 5364 32145 5447 32156
rect 4489 32093 4666 32145
rect 4718 32093 4732 32145
rect 4784 32093 4798 32145
rect 4850 32093 4864 32145
rect 4916 32093 4930 32145
rect 4982 32093 4996 32145
rect 5048 32093 5062 32145
rect 5114 32093 5128 32145
rect 5180 32093 5194 32145
rect 5246 32093 5260 32145
rect 5312 32093 5326 32145
rect 5378 32093 5392 32145
rect 5444 32093 5447 32145
rect 4489 32083 5447 32093
rect 4489 32080 5330 32083
rect 5364 32080 5447 32083
rect 4489 32028 4666 32080
rect 4718 32028 4732 32080
rect 4784 32028 4798 32080
rect 4850 32028 4864 32080
rect 4916 32028 4930 32080
rect 4982 32028 4996 32080
rect 5048 32028 5062 32080
rect 5114 32028 5128 32080
rect 5180 32028 5194 32080
rect 5246 32028 5260 32080
rect 5312 32028 5326 32080
rect 5378 32028 5392 32080
rect 5444 32028 5447 32080
rect 4489 32015 5447 32028
rect 4489 31963 4666 32015
rect 4718 31963 4732 32015
rect 4784 31963 4798 32015
rect 4850 31963 4864 32015
rect 4916 31963 4930 32015
rect 4982 31963 4996 32015
rect 5048 31963 5062 32015
rect 5114 31963 5128 32015
rect 5180 31963 5194 32015
rect 5246 31963 5260 32015
rect 5312 31963 5326 32015
rect 5378 31963 5392 32015
rect 5444 31963 5447 32015
rect 4489 31950 5447 31963
rect 4489 31898 4666 31950
rect 4718 31898 4732 31950
rect 4784 31898 4798 31950
rect 4850 31898 4864 31950
rect 4916 31898 4930 31950
rect 4982 31898 4996 31950
rect 5048 31898 5062 31950
rect 5114 31898 5128 31950
rect 5180 31898 5194 31950
rect 5246 31898 5260 31950
rect 5312 31898 5326 31950
rect 5378 31898 5392 31950
rect 5444 31898 5447 31950
rect 4489 31885 5447 31898
rect 4489 31833 4666 31885
rect 4718 31833 4732 31885
rect 4784 31833 4798 31885
rect 4850 31833 4864 31885
rect 4916 31833 4930 31885
rect 4982 31833 4996 31885
rect 5048 31833 5062 31885
rect 5114 31833 5128 31885
rect 5180 31833 5194 31885
rect 5246 31833 5260 31885
rect 5312 31833 5326 31885
rect 5378 31833 5392 31885
rect 5444 31833 5447 31885
rect 4489 31830 5330 31833
rect 5364 31830 5447 31833
rect 4489 31820 5447 31830
rect 4489 31768 4666 31820
rect 4718 31768 4732 31820
rect 4784 31768 4798 31820
rect 4850 31768 4864 31820
rect 4916 31768 4930 31820
rect 4982 31768 4996 31820
rect 5048 31768 5062 31820
rect 5114 31768 5128 31820
rect 5180 31768 5194 31820
rect 5246 31768 5260 31820
rect 5312 31768 5326 31820
rect 5378 31768 5392 31820
rect 5444 31768 5447 31820
rect 4489 31757 5330 31768
rect 5364 31757 5447 31768
rect 4489 31755 5447 31757
rect 4489 31703 4666 31755
rect 4718 31703 4732 31755
rect 4784 31703 4798 31755
rect 4850 31703 4864 31755
rect 4916 31703 4930 31755
rect 4982 31703 4996 31755
rect 5048 31703 5062 31755
rect 5114 31703 5128 31755
rect 5180 31703 5194 31755
rect 5246 31703 5260 31755
rect 5312 31703 5326 31755
rect 5378 31703 5392 31755
rect 5444 31703 5447 31755
rect 4489 31690 5330 31703
rect 5364 31690 5447 31703
rect 4489 31638 4666 31690
rect 4718 31638 4732 31690
rect 4784 31638 4798 31690
rect 4850 31638 4864 31690
rect 4916 31638 4930 31690
rect 4982 31638 4996 31690
rect 5048 31638 5062 31690
rect 5114 31638 5128 31690
rect 5180 31638 5194 31690
rect 5246 31638 5260 31690
rect 5312 31638 5326 31690
rect 5378 31638 5392 31690
rect 5444 31638 5447 31690
rect 4489 31625 5330 31638
rect 5364 31625 5447 31638
rect 4489 31573 4666 31625
rect 4718 31573 4732 31625
rect 4784 31573 4798 31625
rect 4850 31573 4864 31625
rect 4916 31573 4930 31625
rect 4982 31573 4996 31625
rect 5048 31573 5062 31625
rect 5114 31573 5128 31625
rect 5180 31573 5194 31625
rect 5246 31573 5260 31625
rect 5312 31573 5326 31625
rect 5378 31573 5392 31625
rect 5444 31573 5447 31625
rect 4489 31572 5447 31573
rect 4489 31560 5330 31572
rect 5364 31560 5447 31572
rect 4489 31508 4666 31560
rect 4718 31508 4732 31560
rect 4784 31508 4798 31560
rect 4850 31508 4864 31560
rect 4916 31508 4930 31560
rect 4982 31508 4996 31560
rect 5048 31508 5062 31560
rect 5114 31508 5128 31560
rect 5180 31508 5194 31560
rect 5246 31508 5260 31560
rect 5312 31508 5326 31560
rect 5378 31508 5392 31560
rect 5444 31508 5447 31560
rect 4489 31499 5447 31508
rect 4489 31495 5330 31499
rect 5364 31495 5447 31499
rect 4489 31443 4666 31495
rect 4718 31443 4732 31495
rect 4784 31443 4798 31495
rect 4850 31443 4864 31495
rect 4916 31443 4930 31495
rect 4982 31443 4996 31495
rect 5048 31443 5062 31495
rect 5114 31443 5128 31495
rect 5180 31443 5194 31495
rect 5246 31443 5260 31495
rect 5312 31443 5326 31495
rect 5378 31443 5392 31495
rect 5444 31443 5447 31495
rect 4489 31430 5447 31443
rect 4489 31378 4666 31430
rect 4718 31378 4732 31430
rect 4784 31378 4798 31430
rect 4850 31378 4864 31430
rect 4916 31378 4930 31430
rect 4982 31378 4996 31430
rect 5048 31378 5062 31430
rect 5114 31378 5128 31430
rect 5180 31378 5194 31430
rect 5246 31378 5260 31430
rect 5312 31378 5326 31430
rect 5378 31378 5392 31430
rect 5444 31378 5447 31430
rect 4489 31365 5447 31378
rect 4489 31313 4666 31365
rect 4718 31313 4732 31365
rect 4784 31313 4798 31365
rect 4850 31313 4864 31365
rect 4916 31313 4930 31365
rect 4982 31313 4996 31365
rect 5048 31313 5062 31365
rect 5114 31313 5128 31365
rect 5180 31313 5194 31365
rect 5246 31313 5260 31365
rect 5312 31313 5326 31365
rect 5378 31313 5392 31365
rect 5444 31313 5447 31365
rect 4489 31300 5447 31313
rect 4489 31248 4666 31300
rect 4718 31248 4732 31300
rect 4784 31248 4798 31300
rect 4850 31248 4864 31300
rect 4916 31248 4930 31300
rect 4982 31248 4996 31300
rect 5048 31248 5062 31300
rect 5114 31248 5128 31300
rect 5180 31248 5194 31300
rect 5246 31248 5260 31300
rect 5312 31248 5326 31300
rect 5378 31248 5392 31300
rect 5444 31248 5447 31300
rect 4489 31246 5330 31248
rect 5364 31246 5447 31248
rect 4489 31235 5447 31246
rect 4489 31183 4666 31235
rect 4718 31183 4732 31235
rect 4784 31183 4798 31235
rect 4850 31183 4864 31235
rect 4916 31183 4930 31235
rect 4982 31183 4996 31235
rect 5048 31183 5062 31235
rect 5114 31183 5128 31235
rect 5180 31183 5194 31235
rect 5246 31183 5260 31235
rect 5312 31183 5326 31235
rect 5378 31183 5392 31235
rect 5444 31183 5447 31235
rect 4489 31173 5330 31183
rect 5364 31173 5447 31183
rect 4489 31170 5447 31173
rect 4489 31118 4666 31170
rect 4718 31118 4732 31170
rect 4784 31118 4798 31170
rect 4850 31118 4864 31170
rect 4916 31118 4930 31170
rect 4982 31118 4996 31170
rect 5048 31118 5062 31170
rect 5114 31118 5128 31170
rect 5180 31118 5194 31170
rect 5246 31118 5260 31170
rect 5312 31118 5326 31170
rect 5378 31118 5392 31170
rect 5444 31118 5447 31170
rect 4489 31105 5330 31118
rect 5364 31105 5447 31118
rect 4489 31053 4666 31105
rect 4718 31053 4732 31105
rect 4784 31053 4798 31105
rect 4850 31053 4864 31105
rect 4916 31053 4930 31105
rect 4982 31053 4996 31105
rect 5048 31053 5062 31105
rect 5114 31053 5128 31105
rect 5180 31053 5194 31105
rect 5246 31053 5260 31105
rect 5312 31053 5326 31105
rect 5378 31053 5392 31105
rect 5444 31053 5447 31105
rect 4489 31040 5330 31053
rect 5364 31040 5447 31053
rect 4489 30988 4666 31040
rect 4718 30988 4732 31040
rect 4784 30988 4798 31040
rect 4850 30988 4864 31040
rect 4916 30988 4930 31040
rect 4982 30988 4996 31040
rect 5048 30988 5062 31040
rect 5114 30988 5128 31040
rect 5180 30988 5194 31040
rect 5246 30988 5260 31040
rect 5312 30988 5326 31040
rect 5378 30988 5392 31040
rect 5444 30988 5447 31040
rect 4489 30975 5330 30988
rect 5364 30975 5447 30988
rect 4489 30923 4666 30975
rect 4718 30923 4732 30975
rect 4784 30923 4798 30975
rect 4850 30923 4864 30975
rect 4916 30923 4930 30975
rect 4982 30923 4996 30975
rect 5048 30923 5062 30975
rect 5114 30923 5128 30975
rect 5180 30923 5194 30975
rect 5246 30923 5260 30975
rect 5312 30923 5326 30975
rect 5378 30923 5392 30975
rect 5444 30923 5447 30975
rect 4489 30915 5447 30923
rect 4489 30910 5330 30915
rect 5364 30910 5447 30915
rect 4489 30858 4666 30910
rect 4718 30858 4732 30910
rect 4784 30858 4798 30910
rect 4850 30858 4864 30910
rect 4916 30858 4930 30910
rect 4982 30858 4996 30910
rect 5048 30858 5062 30910
rect 5114 30858 5128 30910
rect 5180 30858 5194 30910
rect 5246 30858 5260 30910
rect 5312 30858 5326 30910
rect 5378 30858 5392 30910
rect 5444 30858 5447 30910
rect 4489 30845 5447 30858
rect 4489 30793 4666 30845
rect 4718 30793 4732 30845
rect 4784 30793 4798 30845
rect 4850 30793 4864 30845
rect 4916 30793 4930 30845
rect 4982 30793 4996 30845
rect 5048 30793 5062 30845
rect 5114 30793 5128 30845
rect 5180 30793 5194 30845
rect 5246 30793 5260 30845
rect 5312 30793 5326 30845
rect 5378 30793 5392 30845
rect 5444 30793 5447 30845
rect 4489 30780 5447 30793
rect 4489 30728 4666 30780
rect 4718 30728 4732 30780
rect 4784 30728 4798 30780
rect 4850 30728 4864 30780
rect 4916 30728 4930 30780
rect 4982 30728 4996 30780
rect 5048 30728 5062 30780
rect 5114 30728 5128 30780
rect 5180 30728 5194 30780
rect 5246 30728 5260 30780
rect 5312 30728 5326 30780
rect 5378 30728 5392 30780
rect 5444 30728 5447 30780
rect 4489 30715 5447 30728
rect 4489 30663 4666 30715
rect 4718 30663 4732 30715
rect 4784 30663 4798 30715
rect 4850 30663 4864 30715
rect 4916 30663 4930 30715
rect 4982 30663 4996 30715
rect 5048 30663 5062 30715
rect 5114 30663 5128 30715
rect 5180 30663 5194 30715
rect 5246 30663 5260 30715
rect 5312 30663 5326 30715
rect 5378 30663 5392 30715
rect 5444 30663 5447 30715
rect 4489 30662 5330 30663
rect 5364 30662 5447 30663
rect 4489 30650 5447 30662
rect 4489 30598 4666 30650
rect 4718 30598 4732 30650
rect 4784 30598 4798 30650
rect 4850 30598 4864 30650
rect 4916 30598 4930 30650
rect 4982 30598 4996 30650
rect 5048 30598 5062 30650
rect 5114 30598 5128 30650
rect 5180 30598 5194 30650
rect 5246 30598 5260 30650
rect 5312 30598 5326 30650
rect 5378 30598 5392 30650
rect 5444 30598 5447 30650
rect 4489 30589 5330 30598
rect 5364 30589 5447 30598
rect 4489 30585 5447 30589
rect 4489 30533 4666 30585
rect 4718 30533 4732 30585
rect 4784 30533 4798 30585
rect 4850 30533 4864 30585
rect 4916 30533 4930 30585
rect 4982 30533 4996 30585
rect 5048 30533 5062 30585
rect 5114 30533 5128 30585
rect 5180 30533 5194 30585
rect 5246 30533 5260 30585
rect 5312 30533 5326 30585
rect 5378 30533 5392 30585
rect 5444 30533 5447 30585
rect 4489 30520 5330 30533
rect 5364 30520 5447 30533
rect 4489 30468 4666 30520
rect 4718 30468 4732 30520
rect 4784 30468 4798 30520
rect 4850 30468 4864 30520
rect 4916 30468 4930 30520
rect 4982 30468 4996 30520
rect 5048 30468 5062 30520
rect 5114 30468 5128 30520
rect 5180 30468 5194 30520
rect 5246 30468 5260 30520
rect 5312 30468 5326 30520
rect 5378 30468 5392 30520
rect 5444 30468 5447 30520
rect 4489 30455 5330 30468
rect 5364 30455 5447 30468
rect 3076 30378 3122 30416
rect 3076 30344 3082 30378
rect 3116 30344 3122 30378
rect 3076 30306 3122 30344
rect 4489 30403 4666 30455
rect 4718 30403 4732 30455
rect 4784 30403 4798 30455
rect 4850 30403 4864 30455
rect 4916 30403 4930 30455
rect 4982 30403 4996 30455
rect 5048 30403 5062 30455
rect 5114 30403 5128 30455
rect 5180 30403 5194 30455
rect 5246 30403 5260 30455
rect 5312 30403 5326 30455
rect 5378 30403 5392 30455
rect 5444 30403 5447 30455
rect 4489 30390 5330 30403
rect 5364 30390 5447 30403
rect 4489 30338 4666 30390
rect 4718 30338 4732 30390
rect 4784 30338 4798 30390
rect 4850 30338 4864 30390
rect 4916 30338 4930 30390
rect 4982 30338 4996 30390
rect 5048 30338 5062 30390
rect 5114 30338 5128 30390
rect 5180 30338 5194 30390
rect 5246 30338 5260 30390
rect 5312 30338 5326 30390
rect 5378 30338 5392 30390
rect 5444 30338 5447 30390
rect 4489 30332 5447 30338
rect 7740 39192 7746 39226
rect 7780 39192 7786 39226
rect 7740 39154 7786 39192
rect 7740 39120 7746 39154
rect 7780 39120 7786 39154
rect 7740 39082 7786 39120
rect 7740 39048 7746 39082
rect 7780 39048 7786 39082
rect 7740 39010 7786 39048
rect 7740 38976 7746 39010
rect 7780 38976 7786 39010
rect 7740 38938 7786 38976
rect 7740 38904 7746 38938
rect 7780 38904 7786 38938
rect 7740 38866 7786 38904
rect 7740 38832 7746 38866
rect 7780 38832 7786 38866
rect 7740 38794 7786 38832
rect 7740 38760 7746 38794
rect 7780 38760 7786 38794
rect 7740 38722 7786 38760
rect 7740 38688 7746 38722
rect 7780 38688 7786 38722
rect 7740 38650 7786 38688
rect 7740 38616 7746 38650
rect 7780 38616 7786 38650
rect 7740 38578 7786 38616
rect 7740 38544 7746 38578
rect 7780 38544 7786 38578
rect 7740 38506 7786 38544
rect 7740 38472 7746 38506
rect 7780 38472 7786 38506
rect 7740 38434 7786 38472
rect 7740 38400 7746 38434
rect 7780 38400 7786 38434
rect 7740 38362 7786 38400
rect 7740 38328 7746 38362
rect 7780 38328 7786 38362
rect 7740 38290 7786 38328
rect 7740 38256 7746 38290
rect 7780 38256 7786 38290
rect 7740 38218 7786 38256
rect 7740 38184 7746 38218
rect 7780 38184 7786 38218
rect 7740 38146 7786 38184
rect 7740 38112 7746 38146
rect 7780 38112 7786 38146
rect 7740 38074 7786 38112
rect 7740 38040 7746 38074
rect 7780 38040 7786 38074
rect 7740 38002 7786 38040
rect 7740 37968 7746 38002
rect 7780 37968 7786 38002
rect 7740 37930 7786 37968
rect 7740 37896 7746 37930
rect 7780 37896 7786 37930
rect 7740 37858 7786 37896
rect 7740 37824 7746 37858
rect 7780 37824 7786 37858
rect 7740 37786 7786 37824
rect 7740 37752 7746 37786
rect 7780 37752 7786 37786
rect 7740 37714 7786 37752
rect 7740 37680 7746 37714
rect 7780 37680 7786 37714
rect 7740 37642 7786 37680
rect 7740 37608 7746 37642
rect 7780 37608 7786 37642
rect 7740 37570 7786 37608
rect 7740 37536 7746 37570
rect 7780 37536 7786 37570
rect 7740 37498 7786 37536
rect 7740 37464 7746 37498
rect 7780 37464 7786 37498
rect 7740 37426 7786 37464
rect 7740 37392 7746 37426
rect 7780 37392 7786 37426
rect 7740 37354 7786 37392
rect 7740 37320 7746 37354
rect 7780 37320 7786 37354
rect 7740 37282 7786 37320
rect 7740 37248 7746 37282
rect 7780 37248 7786 37282
rect 7740 37210 7786 37248
rect 7740 37176 7746 37210
rect 7780 37176 7786 37210
rect 7740 37138 7786 37176
rect 7740 37104 7746 37138
rect 7780 37104 7786 37138
rect 7740 37066 7786 37104
rect 7740 37032 7746 37066
rect 7780 37032 7786 37066
rect 7740 36994 7786 37032
rect 7740 36960 7746 36994
rect 7780 36960 7786 36994
rect 7740 36922 7786 36960
rect 7740 36888 7746 36922
rect 7780 36888 7786 36922
rect 7740 36850 7786 36888
rect 7740 36816 7746 36850
rect 7780 36816 7786 36850
rect 7740 36778 7786 36816
rect 7740 36744 7746 36778
rect 7780 36744 7786 36778
rect 7740 36706 7786 36744
rect 7740 36672 7746 36706
rect 7780 36672 7786 36706
rect 7740 36634 7786 36672
rect 7740 36600 7746 36634
rect 7780 36600 7786 36634
rect 7740 36562 7786 36600
rect 7740 36528 7746 36562
rect 7780 36528 7786 36562
rect 7740 36490 7786 36528
rect 7740 36456 7746 36490
rect 7780 36456 7786 36490
rect 7740 36418 7786 36456
rect 7740 36384 7746 36418
rect 7780 36384 7786 36418
rect 7740 36346 7786 36384
rect 7740 36312 7746 36346
rect 7780 36312 7786 36346
rect 7740 36274 7786 36312
rect 7740 36240 7746 36274
rect 7780 36240 7786 36274
rect 7740 36202 7786 36240
rect 7740 36168 7746 36202
rect 7780 36168 7786 36202
rect 7740 36130 7786 36168
rect 7740 36096 7746 36130
rect 7780 36096 7786 36130
rect 7740 36058 7786 36096
rect 7740 36024 7746 36058
rect 7780 36024 7786 36058
rect 7740 35986 7786 36024
rect 7740 35952 7746 35986
rect 7780 35952 7786 35986
rect 7740 35914 7786 35952
rect 7740 35880 7746 35914
rect 7780 35880 7786 35914
rect 7740 35842 7786 35880
rect 7740 35808 7746 35842
rect 7780 35808 7786 35842
rect 7740 35770 7786 35808
rect 7740 35736 7746 35770
rect 7780 35736 7786 35770
rect 7740 35698 7786 35736
rect 7740 35664 7746 35698
rect 7780 35664 7786 35698
rect 7740 35626 7786 35664
rect 7740 35592 7746 35626
rect 7780 35592 7786 35626
rect 7740 35554 7786 35592
rect 7740 35520 7746 35554
rect 7780 35520 7786 35554
rect 7740 35482 7786 35520
rect 7740 35448 7746 35482
rect 7780 35448 7786 35482
rect 7740 35410 7786 35448
rect 7740 35376 7746 35410
rect 7780 35376 7786 35410
rect 7740 35338 7786 35376
rect 7740 35304 7746 35338
rect 7780 35304 7786 35338
rect 7740 35266 7786 35304
rect 7740 35232 7746 35266
rect 7780 35232 7786 35266
rect 7740 35194 7786 35232
rect 7740 35160 7746 35194
rect 7780 35160 7786 35194
rect 7740 35122 7786 35160
rect 7740 35088 7746 35122
rect 7780 35088 7786 35122
rect 7740 35050 7786 35088
rect 7740 35016 7746 35050
rect 7780 35016 7786 35050
rect 7740 34978 7786 35016
rect 7740 34944 7746 34978
rect 7780 34944 7786 34978
rect 7740 34906 7786 34944
rect 7740 34872 7746 34906
rect 7780 34872 7786 34906
rect 7740 34834 7786 34872
rect 7740 34800 7746 34834
rect 7780 34800 7786 34834
rect 7740 34762 7786 34800
rect 7740 34728 7746 34762
rect 7780 34728 7786 34762
rect 7740 34690 7786 34728
rect 7740 34656 7746 34690
rect 7780 34656 7786 34690
rect 7740 34618 7786 34656
rect 7740 34584 7746 34618
rect 7780 34584 7786 34618
rect 7740 34546 7786 34584
rect 7740 34512 7746 34546
rect 7780 34512 7786 34546
rect 7740 34474 7786 34512
rect 7740 34440 7746 34474
rect 7780 34440 7786 34474
rect 7740 34402 7786 34440
rect 7740 34368 7746 34402
rect 7780 34368 7786 34402
rect 7740 34330 7786 34368
rect 7740 34296 7746 34330
rect 7780 34296 7786 34330
rect 7740 34258 7786 34296
rect 7740 34224 7746 34258
rect 7780 34224 7786 34258
rect 7740 34186 7786 34224
rect 7740 34152 7746 34186
rect 7780 34152 7786 34186
rect 7740 34114 7786 34152
rect 7740 34080 7746 34114
rect 7780 34080 7786 34114
rect 7740 34042 7786 34080
rect 7740 34008 7746 34042
rect 7780 34008 7786 34042
rect 7740 33970 7786 34008
rect 7740 33936 7746 33970
rect 7780 33936 7786 33970
rect 7740 33898 7786 33936
rect 7740 33864 7746 33898
rect 7780 33864 7786 33898
rect 7740 33826 7786 33864
rect 7740 33792 7746 33826
rect 7780 33792 7786 33826
rect 7740 33754 7786 33792
rect 7740 33720 7746 33754
rect 7780 33720 7786 33754
rect 7740 33682 7786 33720
rect 7740 33648 7746 33682
rect 7780 33648 7786 33682
rect 7740 33610 7786 33648
rect 7740 33576 7746 33610
rect 7780 33576 7786 33610
rect 7740 33538 7786 33576
rect 7740 33504 7746 33538
rect 7780 33504 7786 33538
rect 7740 33466 7786 33504
rect 7740 33432 7746 33466
rect 7780 33432 7786 33466
rect 7740 33394 7786 33432
rect 7740 33360 7746 33394
rect 7780 33360 7786 33394
rect 7740 33322 7786 33360
rect 7740 33288 7746 33322
rect 7780 33288 7786 33322
rect 7740 33250 7786 33288
rect 7740 33216 7746 33250
rect 7780 33216 7786 33250
rect 7740 33178 7786 33216
rect 7740 33144 7746 33178
rect 7780 33144 7786 33178
rect 7740 33106 7786 33144
rect 7740 33072 7746 33106
rect 7780 33072 7786 33106
rect 7740 33034 7786 33072
rect 7740 33000 7746 33034
rect 7780 33000 7786 33034
rect 7740 32962 7786 33000
rect 7740 32928 7746 32962
rect 7780 32928 7786 32962
rect 7740 32890 7786 32928
rect 7740 32856 7746 32890
rect 7780 32856 7786 32890
rect 7740 32818 7786 32856
rect 7740 32784 7746 32818
rect 7780 32784 7786 32818
rect 7740 32746 7786 32784
rect 7740 32712 7746 32746
rect 7780 32712 7786 32746
rect 7740 32674 7786 32712
rect 7740 32640 7746 32674
rect 7780 32640 7786 32674
rect 7740 32602 7786 32640
rect 7740 32568 7746 32602
rect 7780 32568 7786 32602
rect 7740 32530 7786 32568
rect 7740 32496 7746 32530
rect 7780 32496 7786 32530
rect 7740 32458 7786 32496
rect 7740 32424 7746 32458
rect 7780 32424 7786 32458
rect 7740 32386 7786 32424
rect 7740 32352 7746 32386
rect 7780 32352 7786 32386
rect 7740 32314 7786 32352
rect 7740 32280 7746 32314
rect 7780 32280 7786 32314
rect 7740 32242 7786 32280
rect 7740 32208 7746 32242
rect 7780 32208 7786 32242
rect 7740 32170 7786 32208
rect 7740 32136 7746 32170
rect 7780 32136 7786 32170
rect 7740 32098 7786 32136
rect 7740 32064 7746 32098
rect 7780 32064 7786 32098
rect 7740 32026 7786 32064
rect 7740 31992 7746 32026
rect 7780 31992 7786 32026
rect 7740 31954 7786 31992
rect 7740 31920 7746 31954
rect 7780 31920 7786 31954
rect 7740 31882 7786 31920
rect 7740 31848 7746 31882
rect 7780 31848 7786 31882
rect 7740 31810 7786 31848
rect 7740 31776 7746 31810
rect 7780 31776 7786 31810
rect 7740 31738 7786 31776
rect 7740 31704 7746 31738
rect 7780 31704 7786 31738
rect 7740 31666 7786 31704
rect 7740 31632 7746 31666
rect 7780 31632 7786 31666
rect 7740 31594 7786 31632
rect 7740 31560 7746 31594
rect 7780 31560 7786 31594
rect 7740 31522 7786 31560
rect 7740 31488 7746 31522
rect 7780 31488 7786 31522
rect 7740 31450 7786 31488
rect 7740 31416 7746 31450
rect 7780 31416 7786 31450
rect 7740 31378 7786 31416
rect 7740 31344 7746 31378
rect 7780 31344 7786 31378
rect 7740 31306 7786 31344
rect 7740 31272 7746 31306
rect 7780 31272 7786 31306
rect 7740 31234 7786 31272
rect 7740 31200 7746 31234
rect 7780 31200 7786 31234
rect 7740 31162 7786 31200
rect 7740 31128 7746 31162
rect 7780 31128 7786 31162
rect 7740 31090 7786 31128
rect 7740 31056 7746 31090
rect 7780 31056 7786 31090
rect 7740 31018 7786 31056
rect 7740 30984 7746 31018
rect 7780 30984 7786 31018
rect 7740 30946 7786 30984
rect 7740 30912 7746 30946
rect 7780 30912 7786 30946
rect 7740 30874 7786 30912
rect 7740 30840 7746 30874
rect 7780 30840 7786 30874
rect 7740 30801 7786 30840
rect 7740 30767 7746 30801
rect 7780 30767 7786 30801
rect 7740 30728 7786 30767
rect 7740 30694 7746 30728
rect 7780 30694 7786 30728
rect 7740 30655 7786 30694
rect 7740 30621 7746 30655
rect 7780 30621 7786 30655
rect 7740 30582 7786 30621
rect 7740 30548 7746 30582
rect 7780 30548 7786 30582
rect 7740 30509 7786 30548
rect 7740 30475 7746 30509
rect 7780 30475 7786 30509
rect 7740 30436 7786 30475
rect 7740 30402 7746 30436
rect 7780 30402 7786 30436
rect 7740 30363 7786 30402
rect 3076 30272 3082 30306
rect 3116 30272 3122 30306
rect 3076 30234 3122 30272
rect 3076 30200 3082 30234
rect 3116 30200 3122 30234
rect 7740 30329 7746 30363
rect 7780 30329 7786 30363
rect 7740 30290 7786 30329
rect 7740 30256 7746 30290
rect 7780 30256 7786 30290
rect 7740 30217 7786 30256
rect 3076 30162 3122 30200
rect 3076 30128 3082 30162
rect 3116 30128 3122 30162
rect 5634 30197 7482 30203
rect 5634 30163 5646 30197
rect 5680 30163 5721 30197
rect 5755 30163 5796 30197
rect 5830 30163 5871 30197
rect 5905 30163 5946 30197
rect 5980 30163 6021 30197
rect 6055 30163 6096 30197
rect 6130 30163 6171 30197
rect 6205 30163 6246 30197
rect 6280 30163 6321 30197
rect 6355 30163 6396 30197
rect 6430 30163 6471 30197
rect 6505 30163 6546 30197
rect 6580 30163 6621 30197
rect 6655 30163 6696 30197
rect 6730 30163 6770 30197
rect 6804 30163 6844 30197
rect 6878 30163 6918 30197
rect 6952 30163 6992 30197
rect 7026 30163 7066 30197
rect 7100 30163 7140 30197
rect 7174 30163 7214 30197
rect 7248 30163 7288 30197
rect 7322 30163 7362 30197
rect 7396 30163 7436 30197
rect 7470 30163 7482 30197
rect 5634 30157 7482 30163
rect 7740 30183 7746 30217
rect 7780 30183 7786 30217
rect 5634 30144 5701 30157
tri 5701 30144 5714 30157 nw
rect 7740 30144 7786 30183
rect 4863 30131 4869 30134
rect 3076 30090 3122 30128
rect 3076 30056 3082 30090
rect 3116 30056 3122 30090
rect 3677 30125 4869 30131
rect 4921 30125 4946 30134
rect 3677 30091 3689 30125
rect 3723 30091 3764 30125
rect 3798 30091 3839 30125
rect 3873 30091 3914 30125
rect 3948 30091 3989 30125
rect 4023 30091 4064 30125
rect 4098 30091 4139 30125
rect 4173 30091 4214 30125
rect 4248 30091 4289 30125
rect 4323 30091 4364 30125
rect 4398 30091 4439 30125
rect 4473 30091 4514 30125
rect 4548 30091 4589 30125
rect 4623 30091 4664 30125
rect 4698 30091 4739 30125
rect 4773 30091 4814 30125
rect 4848 30091 4869 30125
rect 4923 30091 4946 30125
rect 3677 30085 4869 30091
rect 4863 30082 4869 30085
rect 4921 30082 4946 30091
rect 4998 30082 5022 30134
rect 5074 30082 5098 30134
rect 5150 30082 5174 30134
rect 5226 30082 5232 30134
rect 3076 30018 3122 30056
rect 3076 29984 3082 30018
rect 3116 29984 3122 30018
rect 3076 29946 3122 29984
rect 3076 29912 3082 29946
rect 3116 29912 3122 29946
rect 3076 29874 3122 29912
rect 5634 30002 5680 30144
tri 5680 30123 5701 30144 nw
rect 7740 30110 7746 30144
rect 7780 30110 7786 30144
rect 5634 29968 5640 30002
rect 5674 29968 5680 30002
rect 6188 30099 6240 30105
rect 7740 30071 7786 30110
rect 6188 30035 6240 30047
rect 6348 30002 6354 30054
rect 6406 30002 6418 30054
rect 6470 30002 6476 30054
rect 7740 30037 7746 30071
rect 7780 30037 7786 30071
rect 6188 29977 6240 29983
rect 7740 29998 7786 30037
rect 5634 29928 5680 29968
rect 3076 29840 3082 29874
rect 3116 29840 3122 29874
rect 3076 29802 3122 29840
rect 3076 29768 3082 29802
rect 3116 29768 3122 29802
rect 3550 29905 3602 29911
rect 3550 29841 3602 29853
rect 5261 29905 5313 29911
rect 5261 29841 5313 29853
rect 3550 29783 3602 29789
rect 3076 29730 3122 29768
rect 3076 29696 3082 29730
rect 3116 29696 3122 29730
rect 3076 29658 3122 29696
rect 3076 29624 3082 29658
rect 3116 29624 3122 29658
rect 3076 29586 3122 29624
rect 4409 29617 4455 29789
rect 5261 29783 5313 29789
rect 5634 29894 5640 29928
rect 5674 29894 5680 29928
rect 6483 29922 6489 29974
rect 6541 29922 6553 29974
rect 6605 29922 6611 29974
rect 7740 29964 7746 29998
rect 7780 29964 7786 29998
rect 7740 29925 7786 29964
rect 5634 29854 5680 29894
rect 5634 29820 5640 29854
rect 5674 29820 5680 29854
rect 5634 29780 5680 29820
rect 5634 29746 5640 29780
rect 5674 29746 5680 29780
rect 5634 29706 5680 29746
rect 5634 29672 5640 29706
rect 5674 29672 5680 29706
rect 6202 29888 6564 29894
rect 6202 29854 6214 29888
rect 6248 29854 6286 29888
rect 6320 29854 6446 29888
rect 6480 29854 6518 29888
rect 6552 29854 6564 29888
rect 6202 29848 6564 29854
rect 6202 29818 6254 29848
tri 6254 29818 6284 29848 nw
tri 6326 29818 6356 29848 ne
rect 6356 29818 6410 29848
tri 6410 29818 6440 29848 nw
tri 6482 29818 6512 29848 ne
rect 6512 29818 6564 29848
rect 6202 29692 6250 29818
tri 6250 29814 6254 29818 nw
tri 6356 29814 6360 29818 ne
rect 6360 29746 6406 29818
tri 6406 29814 6410 29818 nw
tri 6512 29814 6516 29818 ne
rect 6516 29692 6564 29818
rect 7740 29891 7746 29925
rect 7780 29891 7786 29925
rect 7740 29852 7786 29891
rect 7740 29818 7746 29852
rect 7780 29818 7786 29852
rect 7740 29779 7786 29818
rect 7740 29745 7746 29779
rect 7780 29745 7786 29779
rect 7740 29706 7786 29745
rect 5634 29631 5680 29672
rect 3076 29552 3082 29586
rect 3116 29552 3122 29586
rect 3076 29514 3122 29552
rect 3076 29480 3082 29514
rect 3116 29480 3122 29514
rect 5634 29597 5640 29631
rect 5674 29597 5680 29631
rect 5634 29556 5680 29597
rect 5634 29522 5640 29556
rect 5674 29522 5680 29556
rect 3076 29442 3122 29480
rect 3076 29408 3082 29442
rect 3116 29408 3122 29442
rect 3076 29370 3122 29408
rect 3076 29336 3082 29370
rect 3116 29336 3122 29370
rect 3550 29481 3602 29487
rect 3550 29417 3602 29429
rect 3550 29359 3602 29365
rect 5261 29481 5313 29487
rect 5261 29417 5313 29429
rect 5261 29359 5313 29365
rect 5634 29481 5680 29522
rect 5634 29447 5640 29481
rect 5674 29447 5680 29481
rect 5634 29406 5680 29447
rect 5634 29372 5640 29406
rect 5674 29372 5680 29406
rect 3076 29298 3122 29336
rect 3076 29264 3082 29298
rect 3116 29264 3122 29298
rect 5634 29331 5680 29372
rect 5634 29297 5640 29331
rect 5674 29297 5680 29331
rect 3076 29226 3122 29264
rect 3703 29269 5227 29275
rect 3703 29235 3715 29269
rect 3749 29235 3789 29269
rect 3823 29235 3863 29269
rect 3897 29235 3937 29269
rect 3971 29235 4011 29269
rect 4045 29235 4085 29269
rect 4119 29235 4159 29269
rect 4193 29235 4232 29269
rect 4266 29235 4305 29269
rect 4339 29235 4378 29269
rect 4412 29235 4451 29269
rect 4485 29235 4524 29269
rect 4558 29235 4597 29269
rect 4631 29235 4670 29269
rect 4704 29235 4743 29269
rect 4777 29235 4816 29269
rect 4850 29235 4889 29269
rect 4923 29235 4962 29269
rect 4996 29235 5035 29269
rect 5069 29235 5108 29269
rect 5142 29235 5181 29269
rect 5215 29235 5227 29269
rect 3703 29229 5227 29235
rect 5634 29256 5680 29297
rect 3076 29192 3082 29226
rect 3116 29192 3122 29226
rect 3076 29154 3122 29192
rect 3076 29120 3082 29154
rect 3116 29120 3122 29154
rect 4201 29145 4207 29147
rect 3076 29082 3122 29120
rect 3703 29139 4207 29145
rect 4259 29139 4271 29147
rect 4323 29145 4329 29147
rect 4323 29139 4376 29145
rect 3703 29105 3715 29139
rect 3749 29105 3792 29139
rect 3826 29105 3869 29139
rect 3903 29105 3946 29139
rect 3980 29105 4023 29139
rect 4057 29105 4100 29139
rect 4134 29105 4177 29139
rect 4323 29105 4330 29139
rect 4364 29105 4376 29139
rect 3703 29099 4207 29105
rect 4201 29095 4207 29099
rect 4259 29095 4271 29105
rect 4323 29099 4376 29105
rect 4323 29095 4329 29099
rect 3076 29048 3082 29082
rect 3116 29048 3122 29082
rect 3076 29010 3122 29048
rect 4409 29016 4455 29229
rect 5634 29222 5640 29256
rect 5674 29222 5680 29256
rect 5634 29181 5680 29222
rect 5634 29147 5640 29181
rect 5674 29147 5680 29181
rect 4738 29145 4744 29147
rect 4503 29139 4744 29145
rect 4503 29105 4515 29139
rect 4549 29105 4590 29139
rect 4624 29105 4665 29139
rect 4699 29105 4740 29139
rect 4503 29099 4744 29105
rect 4738 29095 4744 29099
rect 4796 29095 4808 29147
rect 4860 29145 4866 29147
rect 4860 29139 5235 29145
rect 4860 29105 4890 29139
rect 4924 29105 4965 29139
rect 4999 29105 5040 29139
rect 5074 29105 5115 29139
rect 5149 29105 5189 29139
rect 5223 29105 5235 29139
rect 4860 29099 5235 29105
rect 5634 29106 5680 29147
rect 4860 29095 4866 29099
rect 5634 29072 5640 29106
rect 5674 29072 5680 29106
rect 5634 29031 5680 29072
rect 3076 28976 3082 29010
rect 3116 28976 3122 29010
rect 3076 28938 3122 28976
rect 4374 28957 4380 29009
rect 4432 28957 4444 29009
rect 4496 28957 4502 29009
rect 5634 28997 5640 29031
rect 5674 28997 5680 29031
rect 3076 28904 3082 28938
rect 3116 28904 3122 28938
rect 5634 28956 5680 28997
rect 3076 28866 3122 28904
rect 3076 28832 3082 28866
rect 3116 28832 3122 28866
rect 3076 28794 3122 28832
rect 3550 28921 3602 28927
rect 3550 28857 3602 28869
rect 3550 28799 3602 28805
rect 5261 28921 5313 28927
rect 5261 28857 5313 28869
rect 5261 28799 5313 28805
rect 5634 28922 5640 28956
rect 5674 28922 5680 28956
rect 5634 28881 5680 28922
rect 5634 28847 5640 28881
rect 5674 28847 5680 28881
rect 5634 28806 5680 28847
rect 3076 28760 3082 28794
rect 3116 28760 3122 28794
rect 3076 28722 3122 28760
rect 3076 28688 3082 28722
rect 3116 28688 3122 28722
rect 3076 28650 3122 28688
rect 3076 28616 3082 28650
rect 3116 28616 3122 28650
rect 3076 28578 3122 28616
rect 3076 28544 3082 28578
rect 3116 28544 3122 28578
rect 3076 28506 3122 28544
rect 3076 28472 3082 28506
rect 3116 28472 3122 28506
rect 3076 28440 3122 28472
rect 5634 28772 5640 28806
rect 5674 28772 5680 28806
rect 5634 28731 5680 28772
rect 5634 28697 5640 28731
rect 5674 28697 5680 28731
rect 5634 28656 5680 28697
rect 5634 28622 5640 28656
rect 5674 28622 5680 28656
rect 5634 28581 5680 28622
rect 5634 28547 5640 28581
rect 5674 28547 5680 28581
rect 5634 28506 5680 28547
rect 5634 28472 5640 28506
rect 5674 28472 5680 28506
rect 5634 28443 5680 28472
rect 4663 28440 4669 28443
rect 3076 28434 4669 28440
rect 4721 28434 4736 28443
rect 4788 28434 4803 28443
rect 4855 28434 4870 28443
rect 4922 28434 4937 28443
rect 4989 28434 5004 28443
rect 5056 28434 5071 28443
rect 5123 28434 5138 28443
rect 5190 28434 5205 28443
rect 3076 28400 3154 28434
rect 3188 28400 3228 28434
rect 3262 28400 3302 28434
rect 3336 28400 3376 28434
rect 3410 28400 3450 28434
rect 3484 28400 3523 28434
rect 3557 28400 3596 28434
rect 3630 28400 3669 28434
rect 3703 28400 3742 28434
rect 3776 28400 3815 28434
rect 3849 28400 3888 28434
rect 3922 28400 3961 28434
rect 3995 28400 4034 28434
rect 4068 28400 4107 28434
rect 4141 28400 4180 28434
rect 4214 28400 4253 28434
rect 4287 28400 4326 28434
rect 4360 28400 4399 28434
rect 4433 28400 4472 28434
rect 4506 28400 4545 28434
rect 4579 28400 4618 28434
rect 4652 28400 4669 28434
rect 4725 28400 4736 28434
rect 4798 28400 4803 28434
rect 5123 28400 5129 28434
rect 5190 28400 5202 28434
rect 3076 28394 4669 28400
rect 4663 28391 4669 28394
rect 4721 28391 4736 28400
rect 4788 28391 4803 28400
rect 4855 28391 4870 28400
rect 4922 28391 4937 28400
rect 4989 28391 5004 28400
rect 5056 28391 5071 28400
rect 5123 28391 5138 28400
rect 5190 28391 5205 28400
rect 5257 28391 5272 28443
rect 5324 28391 5339 28443
rect 5391 28391 5406 28443
rect 5458 28391 5473 28443
rect 5525 28434 5539 28443
rect 5591 28434 5605 28443
rect 5528 28400 5539 28434
rect 5601 28400 5605 28434
rect 5525 28391 5539 28400
rect 5591 28391 5605 28400
rect 5657 28394 5680 28443
rect 7740 29672 7746 29706
rect 7780 29672 7786 29706
rect 7740 29633 7786 29672
rect 7740 29599 7746 29633
rect 7780 29599 7786 29633
rect 7740 29560 7786 29599
rect 7740 29526 7746 29560
rect 7780 29526 7786 29560
rect 7740 29487 7786 29526
rect 7740 29453 7746 29487
rect 7780 29453 7786 29487
rect 7740 29414 7786 29453
rect 7740 29380 7746 29414
rect 7780 29380 7786 29414
rect 7740 29341 7786 29380
rect 7740 29307 7746 29341
rect 7780 29307 7786 29341
rect 7740 29268 7786 29307
rect 7740 29234 7746 29268
rect 7780 29234 7786 29268
rect 7740 29195 7786 29234
rect 7740 29161 7746 29195
rect 7780 29161 7786 29195
rect 7740 29122 7786 29161
rect 7740 29088 7746 29122
rect 7780 29088 7786 29122
rect 7740 29049 7786 29088
rect 7740 29015 7746 29049
rect 7780 29015 7786 29049
rect 7740 28976 7786 29015
rect 7740 28942 7746 28976
rect 7780 28942 7786 28976
rect 7740 28903 7786 28942
rect 7740 28869 7746 28903
rect 7780 28869 7786 28903
rect 7740 28830 7786 28869
rect 7740 28796 7746 28830
rect 7780 28796 7786 28830
rect 7740 28757 7786 28796
rect 7740 28723 7746 28757
rect 7780 28723 7786 28757
rect 7740 28684 7786 28723
rect 7740 28650 7746 28684
rect 7780 28650 7786 28684
rect 7740 28611 7786 28650
rect 7740 28577 7746 28611
rect 7780 28577 7786 28611
rect 7740 28538 7786 28577
rect 7740 28504 7746 28538
rect 7780 28504 7786 28538
rect 7740 28465 7786 28504
rect 7740 28431 7746 28465
rect 7780 28431 7786 28465
rect 5657 28391 5663 28394
rect 7740 28392 7786 28431
rect 2816 28356 2822 28390
rect 2856 28356 2862 28390
rect 2816 28318 2862 28356
rect 2816 28284 2822 28318
rect 2856 28284 2862 28318
rect 2816 28246 2862 28284
rect 2816 28212 2822 28246
rect 2856 28212 2862 28246
rect 7740 28358 7746 28392
rect 7780 28358 7786 28392
rect 7740 28319 7786 28358
rect 7740 28285 7746 28319
rect 7780 28285 7786 28319
rect 7740 28246 7786 28285
tri 7735 28212 7740 28217 se
rect 7740 28212 7746 28246
rect 7780 28212 7786 28246
rect 2816 28180 2862 28212
tri 7706 28183 7735 28212 se
rect 7735 28183 7786 28212
rect 3703 28180 3709 28183
rect 2816 28174 3709 28180
rect 3761 28174 3776 28183
rect 2816 28140 2894 28174
rect 2928 28140 2967 28174
rect 3001 28140 3040 28174
rect 3074 28140 3113 28174
rect 3147 28140 3186 28174
rect 3220 28140 3259 28174
rect 3293 28140 3332 28174
rect 3366 28140 3405 28174
rect 3439 28140 3478 28174
rect 3512 28140 3551 28174
rect 3585 28140 3624 28174
rect 3658 28140 3697 28174
rect 3761 28140 3770 28174
rect 2816 28134 3709 28140
rect 3703 28131 3709 28134
rect 3761 28131 3776 28140
rect 3828 28131 3843 28183
rect 3895 28131 3910 28183
rect 3962 28131 3977 28183
rect 4029 28131 4044 28183
rect 4096 28131 4111 28183
rect 4163 28174 4178 28183
rect 4230 28174 4245 28183
rect 4297 28174 4312 28183
rect 4364 28174 4379 28183
rect 4431 28174 4445 28183
rect 4497 28180 4503 28183
rect 5926 28180 7786 28183
rect 4497 28174 7786 28180
rect 4169 28140 4178 28174
rect 4242 28140 4245 28174
rect 4497 28140 4500 28174
rect 4534 28140 4573 28174
rect 4607 28140 4646 28174
rect 4680 28140 4719 28174
rect 4753 28140 4792 28174
rect 4826 28140 4865 28174
rect 4899 28140 4938 28174
rect 4972 28140 5010 28174
rect 5044 28140 5082 28174
rect 5116 28140 5154 28174
rect 5188 28140 5226 28174
rect 5260 28140 5298 28174
rect 5332 28140 5370 28174
rect 5404 28140 5442 28174
rect 5476 28140 5514 28174
rect 5548 28140 5586 28174
rect 5620 28140 5658 28174
rect 5692 28140 5730 28174
rect 5764 28140 5802 28174
rect 5836 28140 5874 28174
rect 5908 28140 5946 28174
rect 5980 28140 6018 28174
rect 6052 28140 6090 28174
rect 6124 28140 6162 28174
rect 6196 28140 6234 28174
rect 6268 28140 6306 28174
rect 6340 28140 6378 28174
rect 6412 28140 6450 28174
rect 6484 28140 6522 28174
rect 6556 28140 6594 28174
rect 6628 28140 6666 28174
rect 6700 28140 6738 28174
rect 6772 28140 6810 28174
rect 6844 28140 6882 28174
rect 6916 28140 6954 28174
rect 6988 28140 7026 28174
rect 7060 28140 7098 28174
rect 7132 28140 7170 28174
rect 7204 28140 7242 28174
rect 7276 28140 7314 28174
rect 7348 28140 7386 28174
rect 7420 28140 7458 28174
rect 7492 28140 7530 28174
rect 7564 28140 7602 28174
rect 7636 28140 7674 28174
rect 7708 28140 7786 28174
rect 4163 28131 4178 28140
rect 4230 28131 4245 28140
rect 4297 28131 4312 28140
rect 4364 28131 4379 28140
rect 4431 28131 4445 28140
rect 4497 28134 7786 28140
rect 4497 28131 4503 28134
rect 5926 28131 7786 28134
rect 8223 30469 8229 30521
rect 8281 30469 8293 30521
rect 8345 30469 8351 30521
rect 4435 26156 4441 26208
rect 4493 26156 4508 26208
rect 4560 26156 4575 26208
rect 4627 26156 4642 26208
rect 4694 26156 4709 26208
rect 4761 26156 4776 26208
rect 4828 26156 4843 26208
rect 4895 26156 4910 26208
rect 4962 26156 4977 26208
rect 5029 26156 5044 26208
rect 5096 26205 5102 26208
rect 5096 26199 5575 26205
rect 5096 26165 5138 26199
rect 5172 26165 5217 26199
rect 5251 26165 5295 26199
rect 5329 26165 5373 26199
rect 5407 26165 5451 26199
rect 5485 26165 5529 26199
rect 5563 26165 5575 26199
rect 5096 26159 5575 26165
rect 5096 26156 5102 26159
rect 4002 26116 4048 26128
rect 4002 26082 4008 26116
rect 4042 26082 4048 26116
rect 4002 26041 4048 26082
rect 4002 26007 4008 26041
rect 4042 26007 4048 26041
rect 4002 25966 4048 26007
rect 4002 25932 4008 25966
rect 4042 25932 4048 25966
rect 4002 25891 4048 25932
rect 4002 25857 4008 25891
rect 4042 25857 4048 25891
rect 4002 25816 4048 25857
rect 4002 25782 4008 25816
rect 4042 25782 4048 25816
rect 4002 25740 4048 25782
rect 4002 25706 4008 25740
rect 4042 25706 4048 25740
rect 2838 25685 3738 25691
rect 2838 25651 2850 25685
rect 2884 25651 2928 25685
rect 2962 25651 3005 25685
rect 3039 25651 3082 25685
rect 3116 25651 3159 25685
rect 3193 25651 3236 25685
rect 3270 25651 3313 25685
rect 3347 25651 3390 25685
rect 3424 25651 3467 25685
rect 3501 25651 3544 25685
rect 3578 25651 3621 25685
rect 3655 25651 3738 25685
rect 2838 25645 3738 25651
tri 3658 25630 3673 25645 ne
rect 3673 25630 3738 25645
tri 3673 25613 3690 25630 ne
rect 3690 25613 3738 25630
tri 3690 25611 3692 25613 ne
rect 3692 25579 3698 25613
rect 3732 25579 3738 25613
rect 2820 25479 2826 25531
rect 2878 25479 2890 25531
rect 2942 25512 2948 25531
rect 2942 25479 2950 25512
rect 2820 25472 2832 25479
rect 2866 25472 2904 25479
rect 2938 25472 2950 25479
rect 2820 25466 2950 25472
rect 3524 25507 3530 25559
rect 3582 25507 3596 25559
rect 3648 25507 3654 25559
rect 3524 25506 3654 25507
rect 3524 25472 3536 25506
rect 3570 25472 3608 25506
rect 3642 25472 3654 25506
rect 3524 25466 3654 25472
rect 3692 25540 3738 25579
rect 4002 25664 4048 25706
rect 4002 25630 4008 25664
rect 4042 25630 4048 25664
rect 4002 25588 4048 25630
rect 3692 25506 3698 25540
rect 3732 25506 3738 25540
rect 3692 25467 3738 25506
rect 3692 25433 3698 25467
rect 3732 25433 3738 25467
rect 3692 25394 3738 25433
rect 3692 25360 3698 25394
rect 3732 25360 3738 25394
rect 3692 25321 3738 25360
rect 3692 25287 3698 25321
rect 3732 25287 3738 25321
rect 3692 25248 3738 25287
rect 3692 25214 3698 25248
rect 3732 25214 3738 25248
rect 3692 25175 3738 25214
rect 3692 25141 3698 25175
rect 3732 25141 3738 25175
rect 3692 25102 3738 25141
rect 3692 25068 3698 25102
rect 3732 25068 3738 25102
rect 3692 25029 3738 25068
rect 3692 24995 3698 25029
rect 3732 24995 3738 25029
rect 3692 24956 3738 24995
rect 3692 24922 3698 24956
rect 3732 24922 3738 24956
rect 3692 24883 3738 24922
rect 3692 24849 3698 24883
rect 3732 24849 3738 24883
rect 3692 24810 3738 24849
rect 3692 24776 3698 24810
rect 3732 24776 3738 24810
rect 3692 24737 3738 24776
rect 3692 24703 3698 24737
rect 3732 24703 3738 24737
rect 3692 24664 3738 24703
rect 3692 24630 3698 24664
rect 3732 24630 3738 24664
rect 3692 24591 3738 24630
rect 3692 24557 3698 24591
rect 3732 24557 3738 24591
rect 3692 24518 3738 24557
rect 3692 24484 3698 24518
rect 3732 24484 3738 24518
rect 3692 24445 3738 24484
rect 3692 24411 3698 24445
rect 3732 24411 3738 24445
rect 3692 24372 3738 24411
rect 3692 24338 3698 24372
rect 3732 24338 3738 24372
rect 3692 24299 3738 24338
rect 3692 24265 3698 24299
rect 3732 24265 3738 24299
rect 3692 24226 3738 24265
rect 3692 24192 3698 24226
rect 3732 24192 3738 24226
rect 3692 24153 3738 24192
rect 3692 24119 3698 24153
rect 3732 24119 3738 24153
rect 3692 24080 3738 24119
rect 3692 24046 3698 24080
rect 3732 24046 3738 24080
rect 3692 24007 3738 24046
rect 3692 23973 3698 24007
rect 3732 23973 3738 24007
rect 3692 23934 3738 23973
rect 3692 23900 3698 23934
rect 3732 23900 3738 23934
rect 3692 23861 3738 23900
rect 3692 23827 3698 23861
rect 3732 23827 3738 23861
rect 3692 23788 3738 23827
rect 3692 23754 3698 23788
rect 3732 23754 3738 23788
rect 3692 23715 3738 23754
rect 3692 23681 3698 23715
rect 3732 23681 3738 23715
rect 3692 23642 3738 23681
rect 3692 23608 3698 23642
rect 3732 23608 3738 23642
rect 3692 23569 3738 23608
rect 3692 23535 3698 23569
rect 3732 23535 3738 23569
rect 3692 23496 3738 23535
rect 3692 23462 3698 23496
rect 3732 23462 3738 23496
rect 3692 23423 3738 23462
rect 3692 23389 3698 23423
rect 3732 23389 3738 23423
rect 3692 23350 3738 23389
rect 3692 23316 3698 23350
rect 3732 23316 3738 23350
rect 3692 23277 3738 23316
rect 3692 23243 3698 23277
rect 3732 23243 3738 23277
rect 3692 23204 3738 23243
rect 3692 23170 3698 23204
rect 3732 23170 3738 23204
rect 3692 23131 3738 23170
rect 3692 23097 3698 23131
rect 3732 23097 3738 23131
rect 3692 23058 3738 23097
rect 3692 23024 3698 23058
rect 3732 23024 3738 23058
rect 3692 22985 3738 23024
rect 3692 22951 3698 22985
rect 3732 22951 3738 22985
rect 3692 22912 3738 22951
rect 3692 22878 3698 22912
rect 3732 22878 3738 22912
rect 3692 22839 3738 22878
rect 3692 22805 3698 22839
rect 3732 22805 3738 22839
rect 3692 22766 3738 22805
rect 3692 22732 3698 22766
rect 3732 22732 3738 22766
rect 3692 22693 3738 22732
rect 3692 22659 3698 22693
rect 3732 22659 3738 22693
rect 3692 22621 3738 22659
rect 3692 22587 3698 22621
rect 3732 22587 3738 22621
rect 3692 22549 3738 22587
rect 3692 22515 3698 22549
rect 3732 22515 3738 22549
rect 3692 22477 3738 22515
rect 3692 22443 3698 22477
rect 3732 22443 3738 22477
rect 3692 22405 3738 22443
rect 3692 22371 3698 22405
rect 3732 22371 3738 22405
rect 3692 22333 3738 22371
rect 3692 22299 3698 22333
rect 3732 22299 3738 22333
rect 3692 22261 3738 22299
rect 3692 22227 3698 22261
rect 3732 22227 3738 22261
rect 2627 21640 2633 21692
rect 2685 21640 2730 21692
rect 2782 21640 2788 21692
rect 2627 21616 2788 21640
rect 2627 21564 2633 21616
rect 2685 21564 2730 21616
rect 2782 21564 2788 21616
rect 2627 19706 2788 21564
rect 2627 19654 2633 19706
rect 2685 19654 2730 19706
rect 2782 19654 2788 19706
rect 2627 19630 2788 19654
rect 2627 19578 2633 19630
rect 2685 19578 2730 19630
rect 2782 19578 2788 19630
rect 2627 18746 2788 19578
rect 2627 18694 2633 18746
rect 2685 18694 2730 18746
rect 2782 18694 2788 18746
rect 2627 17775 2788 18694
rect 2996 22185 3048 22194
rect 2996 22121 3048 22133
rect 2996 19834 3048 22069
rect 3692 22189 3738 22227
rect 3692 22155 3698 22189
rect 3732 22155 3738 22189
rect 3692 22117 3738 22155
rect 3692 22083 3698 22117
rect 3732 22083 3738 22117
rect 3692 22045 3738 22083
rect 3692 22011 3698 22045
rect 3732 22011 3738 22045
rect 3692 21973 3738 22011
rect 3692 21939 3698 21973
rect 3732 21939 3738 21973
rect 3692 21901 3738 21939
rect 3692 21867 3698 21901
rect 3732 21867 3738 21901
rect 3692 21829 3738 21867
rect 3692 21795 3698 21829
rect 3732 21795 3738 21829
rect 3692 21757 3738 21795
rect 3692 21723 3698 21757
rect 3732 21723 3738 21757
rect 3692 21685 3738 21723
rect 3692 21651 3698 21685
rect 3732 21651 3738 21685
rect 3692 21613 3738 21651
rect 3692 21579 3698 21613
rect 3732 21579 3738 21613
rect 3692 21541 3738 21579
rect 3692 21507 3698 21541
rect 3732 21507 3738 21541
rect 3692 21469 3738 21507
rect 3692 21435 3698 21469
rect 3732 21435 3738 21469
rect 3692 21397 3738 21435
rect 3692 21363 3698 21397
rect 3732 21363 3738 21397
rect 3770 25506 3776 25558
rect 3828 25506 3844 25558
rect 3896 25506 3912 25558
rect 3964 25506 3970 25558
rect 3770 21450 3970 25506
rect 4002 25554 4008 25588
rect 4042 25554 4048 25588
rect 4002 25512 4048 25554
rect 4002 25478 4008 25512
rect 4042 25478 4048 25512
rect 4002 25451 4048 25478
rect 4347 26071 4393 26083
rect 4347 26037 4353 26071
rect 4387 26037 4393 26071
rect 4347 25998 4393 26037
rect 4347 25964 4353 25998
rect 4387 25964 4393 25998
rect 4347 25925 4393 25964
rect 4347 25891 4353 25925
rect 4387 25891 4393 25925
rect 4347 25852 4393 25891
rect 4347 25818 4353 25852
rect 4387 25818 4393 25852
rect 4347 25779 4393 25818
rect 4503 26071 4549 26083
rect 4503 26037 4509 26071
rect 4543 26037 4549 26071
rect 4503 25998 4549 26037
rect 4503 25964 4509 25998
rect 4543 25964 4549 25998
rect 4503 25925 4549 25964
rect 4503 25891 4509 25925
rect 4543 25891 4549 25925
rect 4503 25852 4549 25891
rect 4503 25818 4509 25852
rect 4543 25818 4549 25852
rect 4503 25813 4549 25818
rect 4659 26071 4705 26083
rect 4659 26037 4665 26071
rect 4699 26037 4705 26071
rect 4659 25998 4705 26037
rect 4659 25964 4665 25998
rect 4699 25964 4705 25998
rect 4659 25925 4705 25964
rect 4659 25891 4665 25925
rect 4699 25891 4705 25925
rect 4659 25852 4705 25891
rect 4659 25818 4665 25852
rect 4699 25818 4705 25852
rect 4347 25745 4353 25779
rect 4387 25745 4393 25779
rect 4347 25706 4393 25745
rect 4347 25672 4353 25706
rect 4387 25672 4393 25706
rect 4500 25807 4552 25813
rect 4500 25745 4509 25755
rect 4543 25745 4552 25755
rect 4500 25743 4552 25745
rect 4500 25685 4509 25691
rect 4347 25633 4393 25672
rect 4347 25599 4353 25633
rect 4387 25599 4393 25633
rect 4347 25560 4393 25599
rect 4347 25526 4353 25560
rect 4387 25526 4393 25560
rect 4347 25487 4393 25526
rect 4347 25453 4353 25487
rect 4387 25453 4393 25487
rect 4347 25451 4393 25453
rect 4503 25672 4509 25685
rect 4543 25685 4552 25691
rect 4659 25779 4705 25818
rect 4815 26071 4861 26083
rect 4815 26037 4821 26071
rect 4855 26037 4861 26071
rect 4815 25998 4861 26037
rect 4815 25964 4821 25998
rect 4855 25964 4861 25998
rect 4815 25925 4861 25964
rect 4815 25891 4821 25925
rect 4855 25891 4861 25925
rect 4815 25852 4861 25891
rect 4815 25818 4821 25852
rect 4855 25818 4861 25852
rect 4815 25813 4861 25818
rect 4971 26071 5017 26083
rect 4971 26037 4977 26071
rect 5011 26037 5017 26071
rect 4971 25998 5017 26037
rect 4971 25964 4977 25998
rect 5011 25964 5017 25998
rect 4971 25925 5017 25964
rect 4971 25891 4977 25925
rect 5011 25891 5017 25925
rect 4971 25852 5017 25891
rect 4971 25818 4977 25852
rect 5011 25818 5017 25852
rect 4659 25745 4665 25779
rect 4699 25745 4705 25779
rect 4659 25706 4705 25745
rect 4543 25672 4549 25685
rect 4503 25633 4549 25672
rect 4503 25599 4509 25633
rect 4543 25599 4549 25633
rect 4503 25560 4549 25599
rect 4503 25526 4509 25560
rect 4543 25526 4549 25560
rect 4503 25487 4549 25526
rect 4503 25453 4509 25487
rect 4543 25453 4549 25487
rect 3999 25445 4051 25451
rect 3999 25367 4051 25393
rect 3999 25288 4051 25315
rect 3999 25209 4051 25236
rect 3999 25151 4051 25157
rect 4344 25445 4396 25451
rect 4344 25379 4353 25393
rect 4387 25379 4396 25393
rect 4344 25367 4396 25379
rect 4344 25305 4353 25315
rect 4387 25305 4396 25315
rect 4344 25288 4396 25305
rect 4344 25231 4353 25236
rect 4387 25231 4396 25236
rect 4344 25209 4396 25231
rect 4344 25151 4396 25157
rect 4503 25413 4549 25453
rect 4659 25672 4665 25706
rect 4699 25672 4705 25706
rect 4812 25807 4864 25813
rect 4812 25745 4821 25755
rect 4855 25745 4864 25755
rect 4812 25743 4864 25745
rect 4812 25685 4821 25691
rect 4659 25633 4705 25672
rect 4659 25599 4665 25633
rect 4699 25599 4705 25633
rect 4659 25560 4705 25599
rect 4659 25526 4665 25560
rect 4699 25526 4705 25560
rect 4659 25487 4705 25526
rect 4659 25453 4665 25487
rect 4699 25453 4705 25487
rect 4659 25451 4705 25453
rect 4815 25672 4821 25685
rect 4855 25685 4864 25691
rect 4971 25779 5017 25818
rect 5127 26071 5173 26083
rect 5127 26037 5133 26071
rect 5167 26037 5173 26071
rect 5127 25998 5173 26037
rect 5127 25964 5133 25998
rect 5167 25964 5173 25998
rect 5127 25925 5173 25964
rect 5127 25891 5133 25925
rect 5167 25891 5173 25925
rect 5127 25852 5173 25891
rect 5127 25818 5133 25852
rect 5167 25818 5173 25852
rect 5127 25813 5173 25818
rect 5283 26071 5329 26083
rect 5283 26037 5289 26071
rect 5323 26037 5329 26071
rect 5283 25998 5329 26037
rect 5283 25964 5289 25998
rect 5323 25964 5329 25998
rect 5283 25925 5329 25964
rect 5283 25891 5289 25925
rect 5323 25891 5329 25925
rect 5283 25852 5329 25891
rect 5283 25818 5289 25852
rect 5323 25818 5329 25852
rect 4971 25745 4977 25779
rect 5011 25745 5017 25779
rect 4971 25706 5017 25745
rect 4855 25672 4861 25685
rect 4815 25633 4861 25672
rect 4815 25599 4821 25633
rect 4855 25599 4861 25633
rect 4815 25560 4861 25599
rect 4815 25526 4821 25560
rect 4855 25526 4861 25560
rect 4815 25487 4861 25526
rect 4815 25453 4821 25487
rect 4855 25453 4861 25487
rect 4503 25379 4509 25413
rect 4543 25379 4549 25413
rect 4503 25339 4549 25379
rect 4503 25305 4509 25339
rect 4543 25305 4549 25339
rect 4503 25265 4549 25305
rect 4503 25231 4509 25265
rect 4543 25231 4549 25265
rect 4503 25191 4549 25231
rect 4503 25157 4509 25191
rect 4543 25157 4549 25191
rect 4002 25132 4048 25151
rect 4002 25098 4008 25132
rect 4042 25098 4048 25132
rect 4002 25056 4048 25098
rect 4002 25022 4008 25056
rect 4042 25022 4048 25056
rect 4002 24980 4048 25022
rect 4002 24946 4008 24980
rect 4042 24946 4048 24980
rect 4002 24904 4048 24946
rect 4002 24870 4008 24904
rect 4042 24870 4048 24904
rect 4002 24828 4048 24870
rect 4002 24794 4008 24828
rect 4042 24794 4048 24828
rect 4002 24752 4048 24794
rect 4002 24718 4008 24752
rect 4042 24718 4048 24752
rect 4002 24706 4048 24718
rect 4347 25117 4393 25151
rect 4347 25083 4353 25117
rect 4387 25083 4393 25117
rect 4347 25043 4393 25083
rect 4347 25009 4353 25043
rect 4387 25009 4393 25043
rect 4347 24969 4393 25009
rect 4347 24935 4353 24969
rect 4387 24935 4393 24969
rect 4347 24895 4393 24935
rect 4347 24861 4353 24895
rect 4387 24861 4393 24895
rect 4347 24821 4393 24861
rect 4347 24787 4353 24821
rect 4387 24787 4393 24821
rect 4347 24747 4393 24787
rect 4347 24713 4353 24747
rect 4387 24713 4393 24747
rect 4347 24701 4393 24713
rect 4503 25117 4549 25157
rect 4656 25445 4708 25451
rect 4656 25379 4665 25393
rect 4699 25379 4708 25393
rect 4656 25367 4708 25379
rect 4656 25305 4665 25315
rect 4699 25305 4708 25315
rect 4656 25288 4708 25305
rect 4656 25231 4665 25236
rect 4699 25231 4708 25236
rect 4656 25209 4708 25231
rect 4656 25151 4708 25157
rect 4815 25413 4861 25453
rect 4971 25672 4977 25706
rect 5011 25672 5017 25706
rect 5124 25807 5176 25813
rect 5124 25745 5133 25755
rect 5167 25745 5176 25755
rect 5124 25743 5176 25745
rect 5124 25685 5133 25691
rect 4971 25633 5017 25672
rect 4971 25599 4977 25633
rect 5011 25599 5017 25633
rect 4971 25560 5017 25599
rect 4971 25526 4977 25560
rect 5011 25526 5017 25560
rect 4971 25487 5017 25526
rect 4971 25453 4977 25487
rect 5011 25453 5017 25487
rect 4971 25451 5017 25453
rect 5127 25672 5133 25685
rect 5167 25685 5176 25691
rect 5283 25779 5329 25818
rect 5439 26071 5485 26083
rect 5439 26037 5445 26071
rect 5479 26037 5485 26071
rect 5439 25998 5485 26037
rect 5439 25964 5445 25998
rect 5479 25964 5485 25998
rect 5439 25925 5485 25964
rect 5439 25891 5445 25925
rect 5479 25891 5485 25925
rect 5439 25852 5485 25891
rect 5439 25818 5445 25852
rect 5479 25818 5485 25852
rect 5439 25813 5485 25818
rect 5595 26071 5641 26083
rect 5595 26037 5601 26071
rect 5635 26037 5641 26071
rect 5595 25998 5641 26037
rect 5595 25964 5601 25998
rect 5635 25964 5641 25998
rect 5595 25925 5641 25964
rect 5595 25891 5601 25925
rect 5635 25891 5641 25925
rect 5595 25852 5641 25891
rect 5595 25818 5601 25852
rect 5635 25818 5641 25852
rect 5283 25745 5289 25779
rect 5323 25745 5329 25779
rect 5283 25706 5329 25745
rect 5167 25672 5173 25685
rect 5127 25633 5173 25672
rect 5127 25599 5133 25633
rect 5167 25599 5173 25633
rect 5127 25560 5173 25599
rect 5127 25526 5133 25560
rect 5167 25526 5173 25560
rect 5127 25487 5173 25526
rect 5127 25453 5133 25487
rect 5167 25453 5173 25487
rect 4815 25379 4821 25413
rect 4855 25379 4861 25413
rect 4815 25339 4861 25379
rect 4815 25305 4821 25339
rect 4855 25305 4861 25339
rect 4815 25265 4861 25305
rect 4815 25231 4821 25265
rect 4855 25231 4861 25265
rect 4815 25191 4861 25231
rect 4815 25157 4821 25191
rect 4855 25157 4861 25191
rect 4503 25083 4509 25117
rect 4543 25083 4549 25117
rect 4503 25043 4549 25083
rect 4503 25009 4509 25043
rect 4543 25009 4549 25043
rect 4503 24969 4549 25009
rect 4503 24935 4509 24969
rect 4543 24935 4549 24969
rect 4503 24895 4549 24935
rect 4503 24861 4509 24895
rect 4543 24861 4549 24895
rect 4503 24821 4549 24861
rect 4503 24787 4509 24821
rect 4543 24787 4549 24821
rect 4503 24747 4549 24787
rect 4503 24713 4509 24747
rect 4543 24713 4549 24747
rect 4503 24701 4549 24713
rect 4659 25117 4705 25151
rect 4659 25083 4665 25117
rect 4699 25083 4705 25117
rect 4659 25043 4705 25083
rect 4659 25009 4665 25043
rect 4699 25009 4705 25043
rect 4659 24969 4705 25009
rect 4659 24935 4665 24969
rect 4699 24935 4705 24969
rect 4659 24895 4705 24935
rect 4659 24861 4665 24895
rect 4699 24861 4705 24895
rect 4659 24821 4705 24861
rect 4659 24787 4665 24821
rect 4699 24787 4705 24821
rect 4659 24747 4705 24787
rect 4659 24713 4665 24747
rect 4699 24713 4705 24747
rect 4659 24701 4705 24713
rect 4815 25117 4861 25157
rect 4968 25445 5020 25451
rect 4968 25379 4977 25393
rect 5011 25379 5020 25393
rect 4968 25367 5020 25379
rect 4968 25305 4977 25315
rect 5011 25305 5020 25315
rect 4968 25288 5020 25305
rect 4968 25231 4977 25236
rect 5011 25231 5020 25236
rect 4968 25209 5020 25231
rect 4968 25151 5020 25157
rect 5127 25413 5173 25453
rect 5283 25672 5289 25706
rect 5323 25672 5329 25706
rect 5436 25807 5488 25813
rect 5436 25745 5445 25755
rect 5479 25745 5488 25755
rect 5436 25743 5488 25745
rect 5436 25685 5445 25691
rect 5283 25633 5329 25672
rect 5283 25599 5289 25633
rect 5323 25599 5329 25633
rect 5283 25560 5329 25599
rect 5283 25526 5289 25560
rect 5323 25526 5329 25560
rect 5283 25487 5329 25526
rect 5283 25453 5289 25487
rect 5323 25453 5329 25487
rect 5283 25451 5329 25453
rect 5439 25672 5445 25685
rect 5479 25685 5488 25691
rect 5595 25779 5641 25818
rect 5595 25745 5601 25779
rect 5635 25745 5641 25779
rect 5595 25706 5641 25745
rect 5479 25672 5485 25685
rect 5439 25633 5485 25672
rect 5439 25599 5445 25633
rect 5479 25599 5485 25633
rect 5439 25560 5485 25599
rect 5439 25526 5445 25560
rect 5479 25526 5485 25560
rect 5439 25487 5485 25526
rect 5439 25453 5445 25487
rect 5479 25453 5485 25487
rect 5127 25379 5133 25413
rect 5167 25379 5173 25413
rect 5127 25339 5173 25379
rect 5127 25305 5133 25339
rect 5167 25305 5173 25339
rect 5127 25265 5173 25305
rect 5127 25231 5133 25265
rect 5167 25231 5173 25265
rect 5127 25191 5173 25231
rect 5127 25157 5133 25191
rect 5167 25157 5173 25191
rect 4815 25083 4821 25117
rect 4855 25083 4861 25117
rect 4815 25043 4861 25083
rect 4815 25009 4821 25043
rect 4855 25009 4861 25043
rect 4815 24969 4861 25009
rect 4815 24935 4821 24969
rect 4855 24935 4861 24969
rect 4815 24895 4861 24935
rect 4815 24861 4821 24895
rect 4855 24861 4861 24895
rect 4815 24821 4861 24861
rect 4815 24787 4821 24821
rect 4855 24787 4861 24821
rect 4815 24747 4861 24787
rect 4815 24713 4821 24747
rect 4855 24713 4861 24747
rect 4815 24701 4861 24713
rect 4971 25117 5017 25151
rect 4971 25083 4977 25117
rect 5011 25083 5017 25117
rect 4971 25043 5017 25083
rect 4971 25009 4977 25043
rect 5011 25009 5017 25043
rect 4971 24969 5017 25009
rect 4971 24935 4977 24969
rect 5011 24935 5017 24969
rect 4971 24895 5017 24935
rect 4971 24861 4977 24895
rect 5011 24861 5017 24895
rect 4971 24821 5017 24861
rect 4971 24787 4977 24821
rect 5011 24787 5017 24821
rect 4971 24747 5017 24787
rect 4971 24713 4977 24747
rect 5011 24713 5017 24747
rect 4971 24701 5017 24713
rect 5127 25117 5173 25157
rect 5280 25445 5332 25451
rect 5280 25379 5289 25393
rect 5323 25379 5332 25393
rect 5280 25367 5332 25379
rect 5280 25305 5289 25315
rect 5323 25305 5332 25315
rect 5280 25288 5332 25305
rect 5280 25231 5289 25236
rect 5323 25231 5332 25236
rect 5280 25209 5332 25231
rect 5280 25151 5332 25157
rect 5439 25413 5485 25453
rect 5595 25672 5601 25706
rect 5635 25672 5641 25706
rect 5595 25633 5641 25672
rect 5595 25599 5601 25633
rect 5635 25599 5641 25633
rect 5595 25560 5641 25599
rect 5595 25526 5601 25560
rect 5635 25526 5641 25560
rect 5595 25487 5641 25526
rect 5595 25453 5601 25487
rect 5635 25453 5641 25487
rect 5595 25451 5641 25453
rect 5940 26071 5986 26083
rect 5940 26037 5946 26071
rect 5980 26037 5986 26071
rect 5940 25998 5986 26037
rect 5940 25964 5946 25998
rect 5980 25964 5986 25998
rect 5940 25925 5986 25964
rect 5940 25891 5946 25925
rect 5980 25891 5986 25925
rect 5940 25852 5986 25891
rect 5940 25818 5946 25852
rect 5980 25818 5986 25852
rect 5940 25779 5986 25818
rect 5940 25745 5946 25779
rect 5980 25745 5986 25779
rect 5940 25706 5986 25745
rect 5940 25672 5946 25706
rect 5980 25672 5986 25706
rect 5940 25633 5986 25672
rect 5940 25599 5946 25633
rect 5980 25599 5986 25633
rect 5940 25560 5986 25599
rect 5940 25526 5946 25560
rect 5980 25526 5986 25560
rect 5940 25487 5986 25526
rect 5940 25453 5946 25487
rect 5980 25453 5986 25487
rect 5940 25451 5986 25453
rect 5439 25379 5445 25413
rect 5479 25379 5485 25413
rect 5439 25339 5485 25379
rect 5439 25305 5445 25339
rect 5479 25305 5485 25339
rect 5439 25265 5485 25305
rect 5439 25231 5445 25265
rect 5479 25231 5485 25265
rect 5439 25191 5485 25231
rect 5439 25157 5445 25191
rect 5479 25157 5485 25191
rect 5127 25083 5133 25117
rect 5167 25083 5173 25117
rect 5127 25043 5173 25083
rect 5127 25009 5133 25043
rect 5167 25009 5173 25043
rect 5127 24969 5173 25009
rect 5127 24935 5133 24969
rect 5167 24935 5173 24969
rect 5127 24895 5173 24935
rect 5127 24861 5133 24895
rect 5167 24861 5173 24895
rect 5127 24821 5173 24861
rect 5127 24787 5133 24821
rect 5167 24787 5173 24821
rect 5127 24747 5173 24787
rect 5127 24713 5133 24747
rect 5167 24713 5173 24747
rect 5127 24701 5173 24713
rect 5283 25117 5329 25151
rect 5283 25083 5289 25117
rect 5323 25083 5329 25117
rect 5283 25043 5329 25083
rect 5283 25009 5289 25043
rect 5323 25009 5329 25043
rect 5283 24969 5329 25009
rect 5283 24935 5289 24969
rect 5323 24935 5329 24969
rect 5283 24895 5329 24935
rect 5283 24861 5289 24895
rect 5323 24861 5329 24895
rect 5283 24821 5329 24861
rect 5283 24787 5289 24821
rect 5323 24787 5329 24821
rect 5283 24747 5329 24787
rect 5283 24713 5289 24747
rect 5323 24713 5329 24747
rect 5283 24701 5329 24713
rect 5439 25117 5485 25157
rect 5592 25445 5644 25451
rect 5592 25379 5601 25393
rect 5635 25379 5644 25393
rect 5592 25367 5644 25379
rect 5592 25305 5601 25315
rect 5635 25305 5644 25315
rect 5592 25288 5644 25305
rect 5592 25231 5601 25236
rect 5635 25231 5644 25236
rect 5592 25209 5644 25231
rect 5592 25151 5644 25157
rect 5937 25445 5989 25451
rect 5937 25379 5946 25393
rect 5980 25379 5989 25393
rect 5937 25367 5989 25379
rect 5937 25305 5946 25315
rect 5980 25305 5989 25315
rect 5937 25288 5989 25305
rect 5937 25231 5946 25236
rect 5980 25231 5989 25236
rect 5937 25209 5989 25231
rect 5937 25151 5989 25157
rect 5439 25083 5445 25117
rect 5479 25083 5485 25117
rect 5439 25043 5485 25083
rect 5439 25009 5445 25043
rect 5479 25009 5485 25043
rect 5439 24969 5485 25009
rect 5439 24935 5445 24969
rect 5479 24935 5485 24969
rect 5439 24895 5485 24935
rect 5439 24861 5445 24895
rect 5479 24861 5485 24895
rect 5439 24821 5485 24861
rect 5439 24787 5445 24821
rect 5479 24787 5485 24821
rect 5439 24747 5485 24787
rect 5439 24713 5445 24747
rect 5479 24713 5485 24747
rect 5439 24701 5485 24713
rect 5595 25117 5641 25151
rect 5595 25083 5601 25117
rect 5635 25083 5641 25117
rect 5595 25043 5641 25083
rect 5595 25009 5601 25043
rect 5635 25009 5641 25043
rect 5595 24969 5641 25009
rect 5595 24935 5601 24969
rect 5635 24935 5641 24969
rect 5595 24895 5641 24935
rect 5595 24861 5601 24895
rect 5635 24861 5641 24895
rect 5595 24821 5641 24861
rect 5595 24787 5601 24821
rect 5635 24787 5641 24821
rect 5595 24747 5641 24787
rect 5595 24713 5601 24747
rect 5635 24713 5641 24747
rect 5595 24701 5641 24713
rect 5940 25117 5986 25151
rect 5940 25083 5946 25117
rect 5980 25083 5986 25117
rect 5940 25043 5986 25083
rect 5940 25009 5946 25043
rect 5980 25009 5986 25043
rect 5940 24969 5986 25009
rect 5940 24935 5946 24969
rect 5980 24935 5986 24969
rect 5940 24895 5986 24935
rect 5940 24861 5946 24895
rect 5980 24861 5986 24895
rect 5940 24821 5986 24861
rect 5940 24787 5946 24821
rect 5980 24787 5986 24821
rect 5940 24747 5986 24787
rect 5940 24713 5946 24747
rect 5980 24713 5986 24747
rect 5940 24701 5986 24713
rect 4451 24184 5901 24190
rect 4451 24150 4555 24184
rect 4589 24150 4687 24184
rect 4721 24150 4760 24184
rect 4794 24150 4833 24184
rect 4867 24150 4906 24184
rect 4940 24150 4979 24184
rect 5013 24150 5052 24184
rect 5086 24150 5125 24184
rect 5159 24150 5198 24184
rect 5232 24150 5271 24184
rect 5305 24150 5344 24184
rect 5378 24150 5417 24184
rect 5451 24150 5490 24184
rect 5524 24150 5564 24184
rect 5598 24150 5638 24184
rect 5672 24150 5712 24184
rect 5746 24150 5786 24184
rect 5820 24150 5901 24184
rect 4451 24144 5901 24150
rect 4451 24112 4505 24144
tri 4505 24112 4537 24144 nw
tri 5815 24112 5847 24144 ne
rect 5847 24112 5901 24144
rect 4451 24078 4460 24112
rect 4494 24078 4503 24112
tri 4503 24110 4505 24112 nw
tri 5847 24110 5849 24112 ne
rect 4451 24039 4503 24078
rect 4451 24005 4460 24039
rect 4494 24005 4503 24039
rect 4451 23966 4503 24005
rect 4451 23932 4460 23966
rect 4494 23932 4503 23966
rect 4451 23893 4503 23932
rect 4451 23859 4460 23893
rect 4494 23859 4503 23893
rect 5849 24078 5858 24112
rect 5892 24078 5901 24112
rect 5849 24040 5901 24078
rect 5849 24006 5858 24040
rect 5892 24006 5901 24040
rect 5849 23968 5901 24006
rect 5849 23934 5858 23968
rect 5892 23934 5901 23968
rect 5849 23896 5901 23934
rect 5849 23862 5858 23896
rect 5892 23862 5901 23896
rect 4451 23844 4503 23859
rect 5048 23854 5178 23860
rect 4451 23786 4460 23792
rect 4494 23786 4503 23792
rect 4451 23780 4503 23786
rect 4451 23713 4460 23728
rect 4494 23713 4503 23728
rect 4639 23838 4856 23840
rect 4639 23786 4646 23838
rect 4698 23786 4722 23838
rect 4774 23786 4797 23838
rect 4849 23786 4856 23838
rect 4639 23774 4856 23786
rect 4639 23722 4646 23774
rect 4698 23722 4722 23774
rect 4774 23722 4797 23774
rect 4849 23722 4856 23774
rect 5048 23838 5060 23854
rect 5166 23838 5178 23854
rect 5048 23722 5055 23838
rect 5171 23722 5178 23838
rect 5303 23848 5433 23854
rect 5303 23838 5315 23848
rect 5421 23838 5433 23848
rect 5303 23722 5310 23838
rect 5426 23722 5433 23838
rect 5849 23844 5901 23862
rect 5849 23790 5858 23792
rect 5892 23790 5901 23792
rect 5849 23780 5901 23790
rect 4451 23674 4503 23713
rect 4451 23640 4460 23674
rect 4494 23640 4503 23674
rect 5849 23718 5858 23728
rect 5892 23718 5901 23728
rect 5849 23680 5901 23718
rect 4451 23601 4503 23640
rect 4451 23567 4460 23601
rect 4494 23567 4503 23601
rect 4451 23528 4503 23567
rect 4451 23494 4460 23528
rect 4494 23494 4503 23528
rect 4451 23455 4503 23494
rect 4451 23421 4460 23455
rect 4494 23421 4503 23455
rect 4451 23382 4503 23421
rect 4451 23348 4460 23382
rect 4494 23348 4503 23382
rect 4451 23309 4503 23348
rect 4451 23275 4460 23309
rect 4494 23275 4503 23309
rect 4451 23236 4503 23275
rect 4451 23202 4460 23236
rect 4494 23202 4503 23236
rect 4451 23163 4503 23202
rect 4451 23129 4460 23163
rect 4494 23129 4503 23163
rect 4451 23090 4503 23129
rect 4451 23056 4460 23090
rect 4494 23056 4503 23090
rect 4451 23017 4503 23056
rect 4451 22983 4460 23017
rect 4494 22983 4503 23017
rect 4451 22944 4503 22983
rect 4451 22910 4460 22944
rect 4494 22910 4503 22944
rect 4451 22871 4503 22910
rect 4451 22837 4460 22871
rect 4494 22837 4503 22871
rect 4451 22798 4503 22837
rect 4451 22764 4460 22798
rect 4494 22764 4503 22798
rect 4451 22725 4503 22764
rect 4451 22691 4460 22725
rect 4494 22691 4503 22725
rect 4451 22652 4503 22691
rect 4451 22618 4460 22652
rect 4494 22618 4503 22652
rect 4451 22579 4503 22618
rect 4451 22545 4460 22579
rect 4494 22545 4503 22579
rect 4451 22506 4503 22545
rect 4451 22472 4460 22506
rect 4494 22472 4503 22506
rect 4451 22433 4503 22472
rect 4451 22399 4460 22433
rect 4494 22399 4503 22433
rect 4451 22360 4503 22399
rect 4451 22326 4460 22360
rect 4494 22326 4503 22360
rect 4451 22287 4503 22326
rect 4451 22253 4460 22287
rect 4494 22253 4503 22287
rect 4451 22214 4503 22253
rect 4451 22180 4460 22214
rect 4494 22180 4503 22214
rect 4451 22141 4503 22180
rect 4451 22107 4460 22141
rect 4494 22107 4503 22141
rect 4879 23660 4931 23672
rect 4879 23626 4888 23660
rect 4922 23626 4931 23660
rect 4879 23587 4931 23626
rect 4879 23553 4888 23587
rect 4922 23553 4931 23587
rect 4879 23514 4931 23553
rect 4879 23480 4888 23514
rect 4922 23480 4931 23514
rect 4879 23441 4931 23480
rect 4879 23407 4888 23441
rect 4922 23407 4931 23441
rect 4879 23368 4931 23407
rect 4879 23334 4888 23368
rect 4922 23334 4931 23368
rect 4879 23295 4931 23334
rect 4879 23261 4888 23295
rect 4922 23261 4931 23295
rect 4879 23222 4931 23261
rect 4879 23188 4888 23222
rect 4922 23188 4931 23222
rect 4879 23149 4931 23188
rect 4879 23115 4888 23149
rect 4922 23115 4931 23149
rect 4879 23076 4931 23115
rect 4879 23042 4888 23076
rect 4922 23042 4931 23076
rect 4879 23003 4931 23042
rect 4879 22969 4888 23003
rect 4922 22969 4931 23003
rect 4879 22930 4931 22969
rect 4879 22896 4888 22930
rect 4922 22896 4931 22930
rect 4879 22857 4931 22896
rect 4879 22823 4888 22857
rect 4922 22823 4931 22857
rect 4879 22784 4931 22823
rect 4879 22750 4888 22784
rect 4922 22750 4931 22784
rect 4879 22711 4931 22750
rect 4879 22677 4888 22711
rect 4922 22677 4931 22711
rect 4879 22638 4931 22677
rect 4879 22604 4888 22638
rect 4922 22604 4931 22638
rect 4879 22565 4931 22604
rect 4879 22531 4888 22565
rect 4922 22531 4931 22565
rect 4879 22524 4931 22531
rect 4879 22460 4888 22472
rect 4922 22460 4931 22472
rect 4879 22385 4888 22408
rect 4922 22385 4931 22408
rect 4879 22346 4931 22385
rect 4879 22312 4888 22346
rect 4922 22312 4931 22346
rect 4879 22273 4931 22312
rect 4879 22239 4888 22273
rect 4922 22239 4931 22273
rect 4879 22200 4931 22239
rect 4879 22166 4888 22200
rect 4922 22166 4931 22200
rect 4879 22127 4931 22166
rect 4451 22068 4503 22107
rect 4451 22034 4460 22068
rect 4494 22034 4503 22068
rect 4630 22106 4686 22115
rect 4738 22106 4750 22115
rect 4802 22106 4834 22115
rect 4630 22072 4642 22106
rect 4676 22072 4686 22106
rect 4749 22072 4750 22106
rect 4822 22072 4834 22106
rect 4630 22063 4686 22072
rect 4738 22063 4750 22072
rect 4802 22063 4834 22072
rect 4879 22093 4888 22127
rect 4922 22093 4931 22127
rect 4451 21995 4503 22034
rect 4451 21961 4460 21995
rect 4494 21961 4503 21995
rect 4451 21922 4503 21961
rect 4451 21888 4460 21922
rect 4494 21888 4503 21922
rect 4451 21849 4503 21888
rect 4451 21815 4460 21849
rect 4494 21815 4503 21849
rect 4451 21776 4503 21815
rect 4451 21742 4460 21776
rect 4494 21742 4503 21776
rect 4451 21703 4503 21742
rect 4451 21669 4460 21703
rect 4494 21669 4503 21703
rect 4451 21630 4503 21669
rect 4451 21596 4460 21630
rect 4494 21596 4503 21630
rect 4451 21557 4503 21596
rect 4451 21523 4460 21557
rect 4494 21523 4503 21557
rect 4451 21484 4503 21523
tri 3970 21450 3972 21452 sw
rect 4451 21450 4460 21484
rect 4494 21450 4503 21484
rect 3770 21436 3972 21450
tri 3972 21436 3986 21450 sw
rect 3770 21413 3986 21436
tri 3986 21413 4009 21436 sw
rect 3770 21411 4009 21413
tri 4009 21411 4011 21413 sw
rect 4451 21411 4503 21450
rect 3770 21377 4011 21411
tri 4011 21377 4045 21411 sw
rect 4451 21377 4460 21411
rect 4494 21377 4503 21411
rect 3770 21370 4045 21377
tri 4045 21370 4052 21377 sw
tri 3770 21363 3777 21370 ne
rect 3777 21363 4052 21370
tri 4052 21363 4059 21370 sw
rect 3692 21325 3738 21363
tri 3777 21340 3800 21363 ne
rect 3800 21340 4059 21363
tri 4059 21340 4082 21363 sw
tri 3800 21338 3802 21340 ne
rect 3802 21338 4082 21340
tri 4082 21338 4084 21340 sw
rect 4451 21338 4503 21377
rect 3692 21291 3698 21325
rect 3732 21291 3738 21325
tri 3802 21304 3836 21338 ne
rect 3836 21304 4084 21338
tri 4084 21304 4118 21338 sw
rect 4451 21304 4460 21338
rect 4494 21304 4503 21338
rect 3692 21253 3738 21291
tri 3836 21290 3850 21304 ne
rect 3850 21290 4118 21304
tri 4118 21290 4132 21304 sw
tri 3850 21267 3873 21290 ne
rect 3873 21274 4132 21290
tri 4132 21274 4148 21290 sw
rect 3873 21267 4148 21274
tri 3873 21265 3875 21267 ne
rect 3875 21265 4148 21267
rect 3692 21219 3698 21253
rect 3732 21219 3738 21253
tri 3875 21231 3909 21265 ne
rect 3909 21231 4148 21265
rect 3692 21181 3738 21219
tri 3909 21217 3923 21231 ne
rect 3923 21217 4148 21231
tri 3923 21194 3946 21217 ne
rect 3946 21194 4148 21217
tri 3946 21192 3948 21194 ne
rect 3692 21147 3698 21181
rect 3732 21147 3738 21181
rect 3692 21109 3738 21147
rect 3692 21075 3698 21109
rect 3732 21075 3738 21109
rect 3692 21037 3738 21075
rect 3692 21003 3698 21037
rect 3732 21003 3738 21037
rect 3692 20965 3738 21003
rect 3692 20931 3698 20965
rect 3732 20931 3738 20965
rect 3692 20893 3738 20931
rect 3692 20859 3698 20893
rect 3732 20859 3738 20893
rect 3692 20821 3738 20859
rect 3692 20787 3698 20821
rect 3732 20787 3738 20821
rect 3692 20749 3738 20787
tri 3932 20756 3948 20772 se
rect 3948 20756 4148 21194
rect 4451 21265 4503 21304
rect 4451 21231 4460 21265
rect 4494 21231 4503 21265
rect 4451 21192 4503 21231
rect 4451 21158 4460 21192
rect 4494 21158 4503 21192
rect 4451 21119 4503 21158
rect 4451 21085 4460 21119
rect 4494 21085 4503 21119
rect 4451 21046 4503 21085
rect 4451 21012 4460 21046
rect 4494 21012 4503 21046
rect 4451 20973 4503 21012
rect 4451 20939 4460 20973
rect 4494 20939 4503 20973
rect 4451 20900 4503 20939
rect 4451 20866 4460 20900
rect 4494 20866 4503 20900
rect 4451 20827 4503 20866
rect 4451 20793 4460 20827
rect 4494 20793 4503 20827
tri 4148 20756 4164 20772 sw
tri 3930 20754 3932 20756 se
rect 3932 20754 4164 20756
tri 4164 20754 4166 20756 sw
rect 4451 20754 4503 20793
rect 3692 20715 3698 20749
rect 3732 20715 3738 20749
tri 3914 20738 3930 20754 se
rect 3930 20738 4166 20754
tri 4166 20738 4182 20754 sw
rect 3692 20677 3738 20715
rect 3692 20643 3698 20677
rect 3732 20643 3738 20677
rect 3692 20605 3738 20643
rect 3692 20571 3698 20605
rect 3732 20571 3738 20605
rect 3692 20533 3738 20571
rect 3692 20499 3698 20533
rect 3732 20499 3738 20533
rect 3692 20461 3738 20499
rect 3692 20427 3698 20461
rect 3732 20427 3738 20461
rect 3692 20389 3738 20427
rect 3692 20355 3698 20389
rect 3732 20355 3738 20389
rect 3692 20317 3738 20355
rect 3692 20283 3698 20317
rect 3732 20283 3738 20317
rect 3692 20245 3738 20283
rect 3692 20211 3698 20245
rect 3732 20211 3738 20245
rect 3692 20173 3738 20211
rect 3692 20139 3698 20173
rect 3732 20139 3738 20173
rect 3692 20101 3738 20139
rect 3692 20067 3698 20101
rect 3732 20067 3738 20101
rect 3692 20029 3738 20067
rect 3692 19995 3698 20029
rect 3732 19995 3738 20029
rect 3692 19957 3738 19995
rect 3692 19923 3698 19957
rect 3732 19923 3738 19957
rect 3692 19885 3738 19923
rect 3692 19851 3698 19885
rect 3732 19851 3738 19885
tri 3048 19834 3064 19850 sw
rect 2996 19818 3064 19834
tri 3064 19818 3080 19834 sw
rect 2996 19816 3080 19818
tri 3080 19816 3082 19818 sw
rect 2996 19764 3002 19816
rect 3054 19764 3066 19816
rect 3118 19764 3124 19816
rect 3692 19813 3738 19851
rect 3692 19779 3698 19813
rect 3732 19779 3738 19813
rect 2996 19747 3065 19764
tri 3065 19747 3082 19764 nw
rect 2996 19745 3063 19747
tri 3063 19745 3065 19747 nw
rect 2996 19741 3059 19745
tri 3059 19741 3063 19745 nw
rect 3692 19741 3738 19779
rect 2996 18473 3048 19741
tri 3048 19730 3059 19741 nw
rect 3692 19707 3698 19741
rect 3732 19707 3738 19741
rect 3692 19669 3738 19707
rect 3692 19635 3698 19669
rect 3732 19635 3738 19669
rect 3692 19597 3738 19635
rect 3692 19563 3698 19597
rect 3732 19563 3738 19597
rect 3692 19525 3738 19563
rect 3692 19491 3698 19525
rect 3732 19491 3738 19525
rect 3692 19453 3738 19491
rect 3692 19419 3698 19453
rect 3732 19419 3738 19453
rect 3692 19381 3738 19419
rect 3692 19347 3698 19381
rect 3732 19347 3738 19381
rect 3692 19309 3738 19347
rect 3692 19275 3698 19309
rect 3732 19275 3738 19309
rect 3692 19237 3738 19275
rect 3692 19203 3698 19237
rect 3732 19203 3738 19237
rect 3692 19165 3738 19203
rect 3692 19131 3698 19165
rect 3732 19131 3738 19165
rect 3692 19093 3738 19131
rect 3692 19059 3698 19093
rect 3732 19059 3738 19093
rect 3692 19021 3738 19059
rect 3692 18987 3698 19021
rect 3732 18987 3738 19021
rect 3692 18949 3738 18987
rect 3692 18915 3698 18949
rect 3732 18915 3738 18949
rect 3692 18877 3738 18915
rect 3692 18843 3698 18877
rect 3732 18843 3738 18877
rect 3692 18805 3738 18843
rect 3692 18771 3698 18805
rect 3732 18771 3738 18805
rect 3692 18733 3738 18771
rect 3692 18699 3698 18733
rect 3732 18699 3738 18733
rect 3692 18661 3738 18699
rect 3692 18627 3698 18661
rect 3732 18627 3738 18661
rect 3692 18589 3738 18627
rect 3692 18555 3698 18589
rect 3732 18555 3738 18589
rect 3692 18543 3738 18555
rect 4451 20720 4460 20754
rect 4494 20720 4503 20754
rect 4451 20681 4503 20720
rect 4451 20647 4460 20681
rect 4494 20647 4503 20681
rect 4451 20608 4503 20647
rect 4451 20574 4460 20608
rect 4494 20574 4503 20608
rect 4451 20535 4503 20574
rect 4451 20501 4460 20535
rect 4494 20501 4503 20535
rect 4451 20462 4503 20501
rect 4879 22054 4931 22093
rect 4879 22020 4888 22054
rect 4922 22020 4931 22054
rect 4879 21981 4931 22020
rect 4879 21947 4888 21981
rect 4922 21947 4931 21981
rect 4879 21908 4931 21947
rect 4879 21874 4888 21908
rect 4922 21874 4931 21908
rect 4879 21835 4931 21874
rect 4879 21801 4888 21835
rect 4922 21801 4931 21835
rect 4879 21762 4931 21801
rect 4879 21728 4888 21762
rect 4922 21728 4931 21762
rect 4879 21689 4931 21728
rect 4879 21655 4888 21689
rect 4922 21655 4931 21689
rect 4879 21616 4931 21655
rect 4879 21582 4888 21616
rect 4922 21582 4931 21616
rect 4879 21543 4931 21582
rect 4879 21509 4888 21543
rect 4922 21509 4931 21543
rect 4879 21470 4931 21509
rect 4879 21436 4888 21470
rect 4922 21436 4931 21470
rect 4879 21397 4931 21436
rect 4879 21363 4888 21397
rect 4922 21363 4931 21397
rect 4879 21324 4931 21363
rect 4879 21290 4888 21324
rect 4922 21290 4931 21324
rect 4879 21251 4931 21290
rect 4879 21217 4888 21251
rect 4922 21217 4931 21251
rect 4879 21178 4931 21217
rect 4879 21144 4888 21178
rect 4922 21144 4931 21178
rect 4879 21105 4931 21144
rect 4879 21071 4888 21105
rect 4922 21071 4931 21105
rect 4879 21032 4931 21071
rect 4879 20998 4888 21032
rect 4922 20998 4931 21032
rect 4879 20959 4931 20998
rect 4879 20925 4888 20959
rect 4922 20925 4931 20959
rect 4879 20886 4931 20925
rect 4879 20852 4888 20886
rect 4922 20852 4931 20886
rect 4879 20813 4931 20852
rect 4879 20779 4888 20813
rect 4922 20779 4931 20813
rect 4879 20740 4931 20779
rect 4879 20706 4888 20740
rect 4922 20706 4931 20740
rect 4879 20667 4931 20706
rect 4879 20633 4888 20667
rect 4922 20633 4931 20667
rect 4879 20594 4931 20633
rect 4879 20560 4888 20594
rect 4922 20560 4931 20594
rect 4879 20520 4931 20560
rect 4879 20486 4888 20520
rect 4922 20486 4931 20520
rect 4879 20474 4931 20486
rect 5187 23637 5239 23649
rect 5187 23603 5196 23637
rect 5230 23603 5239 23637
rect 5187 23564 5239 23603
rect 5187 23530 5196 23564
rect 5230 23530 5239 23564
rect 5187 23491 5239 23530
rect 5187 23457 5196 23491
rect 5230 23457 5239 23491
rect 5187 23418 5239 23457
rect 5187 23384 5196 23418
rect 5230 23384 5239 23418
rect 5187 23345 5239 23384
rect 5187 23311 5196 23345
rect 5230 23311 5239 23345
rect 5187 23272 5239 23311
rect 5187 23238 5196 23272
rect 5230 23238 5239 23272
rect 5187 23199 5239 23238
rect 5187 23165 5196 23199
rect 5230 23165 5239 23199
rect 5187 23126 5239 23165
rect 5187 23092 5196 23126
rect 5230 23092 5239 23126
rect 5187 23053 5239 23092
rect 5187 23019 5196 23053
rect 5230 23019 5239 23053
rect 5187 22980 5239 23019
rect 5187 22946 5196 22980
rect 5230 22946 5239 22980
rect 5187 22907 5239 22946
rect 5187 22873 5196 22907
rect 5230 22873 5239 22907
rect 5187 22834 5239 22873
rect 5187 22800 5196 22834
rect 5230 22800 5239 22834
rect 5187 22761 5239 22800
rect 5187 22727 5196 22761
rect 5230 22727 5239 22761
rect 5187 22688 5239 22727
rect 5187 22654 5196 22688
rect 5230 22654 5239 22688
rect 5187 22615 5239 22654
rect 5187 22581 5196 22615
rect 5230 22581 5239 22615
rect 5187 22542 5239 22581
rect 5187 22508 5196 22542
rect 5230 22508 5239 22542
rect 5187 22469 5239 22508
rect 5187 22435 5196 22469
rect 5230 22435 5239 22469
rect 5187 22396 5239 22435
rect 5187 22362 5196 22396
rect 5230 22362 5239 22396
rect 5187 22323 5239 22362
rect 5187 22289 5196 22323
rect 5230 22289 5239 22323
rect 5187 22250 5239 22289
rect 5187 22216 5196 22250
rect 5230 22216 5239 22250
rect 5187 22177 5239 22216
rect 5187 22143 5196 22177
rect 5230 22143 5239 22177
rect 5187 22104 5239 22143
rect 5187 22070 5196 22104
rect 5230 22070 5239 22104
rect 5187 22031 5239 22070
rect 5187 21997 5196 22031
rect 5230 21997 5239 22031
rect 5187 21958 5239 21997
rect 5187 21924 5196 21958
rect 5230 21924 5239 21958
rect 5187 21885 5239 21924
rect 5187 21851 5196 21885
rect 5230 21851 5239 21885
rect 5187 21812 5239 21851
rect 5187 21778 5196 21812
rect 5230 21778 5239 21812
rect 5187 21739 5239 21778
rect 5187 21705 5196 21739
rect 5230 21705 5239 21739
rect 5187 21686 5239 21705
rect 5187 21632 5196 21634
rect 5230 21632 5239 21634
rect 5187 21622 5239 21632
rect 5187 21559 5196 21570
rect 5230 21559 5239 21570
rect 5187 21520 5239 21559
rect 5187 21486 5196 21520
rect 5230 21486 5239 21520
rect 5187 21447 5239 21486
rect 5187 21413 5196 21447
rect 5230 21413 5239 21447
rect 5187 21374 5239 21413
rect 5187 21340 5196 21374
rect 5230 21340 5239 21374
rect 5187 21301 5239 21340
rect 5187 21267 5196 21301
rect 5230 21267 5239 21301
rect 5187 21228 5239 21267
rect 5187 21194 5196 21228
rect 5230 21194 5239 21228
rect 5187 21155 5239 21194
rect 5187 21121 5196 21155
rect 5230 21121 5239 21155
rect 5187 21082 5239 21121
rect 5187 21048 5196 21082
rect 5230 21048 5239 21082
rect 5187 21009 5239 21048
rect 5187 20975 5196 21009
rect 5230 20975 5239 21009
rect 5187 20936 5239 20975
rect 5187 20902 5196 20936
rect 5230 20902 5239 20936
rect 5187 20863 5239 20902
rect 5187 20829 5196 20863
rect 5230 20829 5239 20863
rect 5187 20790 5239 20829
rect 5187 20756 5196 20790
rect 5230 20756 5239 20790
rect 5187 20717 5239 20756
rect 5187 20683 5196 20717
rect 5230 20683 5239 20717
rect 5187 20644 5239 20683
rect 5187 20610 5196 20644
rect 5230 20610 5239 20644
rect 5187 20571 5239 20610
rect 5187 20537 5196 20571
rect 5230 20537 5239 20571
rect 5187 20498 5239 20537
rect 4451 20428 4460 20462
rect 4494 20428 4503 20462
rect 5187 20464 5196 20498
rect 5230 20464 5239 20498
rect 4451 20389 4503 20428
rect 4451 20355 4460 20389
rect 4494 20355 4503 20389
rect 4451 20316 4503 20355
rect 4630 20449 4856 20451
rect 4630 20445 4646 20449
rect 4630 20411 4642 20445
rect 4630 20397 4646 20411
rect 4698 20397 4722 20449
rect 4774 20397 4797 20449
rect 4849 20397 4856 20449
rect 4630 20385 4856 20397
rect 4630 20373 4646 20385
rect 4630 20339 4642 20373
rect 4630 20333 4646 20339
rect 4698 20333 4722 20385
rect 4774 20333 4797 20385
rect 4849 20333 4856 20385
rect 5187 20425 5239 20464
rect 5187 20391 5196 20425
rect 5230 20391 5239 20425
rect 5187 20352 5239 20391
rect 4451 20282 4460 20316
rect 4494 20282 4503 20316
rect 4451 20244 4503 20282
rect 4451 20210 4460 20244
rect 4494 20210 4503 20244
rect 4451 20172 4503 20210
rect 4451 20138 4460 20172
rect 4494 20138 4503 20172
rect 4451 20130 4503 20138
rect 5187 20318 5196 20352
rect 5230 20318 5239 20352
rect 5187 20278 5239 20318
rect 5187 20244 5196 20278
rect 5230 20244 5239 20278
rect 5187 20204 5239 20244
rect 5187 20170 5196 20204
rect 5230 20170 5239 20204
tri 4503 20130 4506 20133 sw
rect 5187 20130 5239 20170
rect 4451 20100 4506 20130
rect 4451 20066 4460 20100
rect 4494 20099 4506 20100
tri 4506 20099 4537 20130 sw
rect 4494 20093 4855 20099
rect 4494 20066 4585 20093
rect 4451 20059 4585 20066
rect 4619 20059 4660 20093
rect 4694 20059 4735 20093
rect 4769 20059 4809 20093
rect 4843 20059 4855 20093
rect 4451 20054 4855 20059
rect 4451 20028 4472 20054
rect 4588 20053 4855 20054
rect 5187 20096 5196 20130
rect 5230 20096 5239 20130
rect 5187 20056 5239 20096
rect 4588 20036 4611 20053
tri 4611 20036 4628 20053 nw
rect 4893 20036 4945 20048
rect 4451 19994 4460 20028
rect 4451 19956 4472 19994
rect 4451 19922 4460 19956
rect 4588 19938 4594 20036
tri 4594 20019 4611 20036 nw
tri 4714 19964 4727 19977 se
rect 4727 19971 4733 20023
rect 4785 19971 4797 20023
rect 4849 19971 4855 20023
rect 4727 19964 4855 19971
tri 4693 19943 4714 19964 se
rect 4714 19943 4855 19964
rect 4494 19922 4594 19938
rect 4451 19884 4594 19922
rect 4630 19937 4855 19943
rect 4630 19903 4642 19937
rect 4676 19903 4726 19937
rect 4760 19903 4809 19937
rect 4843 19903 4855 19937
rect 4630 19897 4855 19903
tri 4769 19891 4775 19897 ne
rect 4775 19891 4855 19897
rect 4451 19850 4460 19884
rect 4494 19850 4594 19884
tri 4775 19863 4803 19891 ne
rect 4451 19818 4594 19850
tri 4594 19818 4597 19821 sw
rect 4451 19812 4597 19818
rect 4451 19778 4460 19812
rect 4494 19787 4597 19812
tri 4597 19787 4628 19818 sw
rect 4494 19781 4775 19787
rect 4494 19778 4585 19781
rect 4451 19747 4585 19778
rect 4619 19747 4657 19781
rect 4691 19747 4729 19781
rect 4763 19747 4775 19781
rect 4451 19741 4775 19747
rect 4451 19740 4598 19741
rect 4451 19706 4460 19740
rect 4494 19711 4598 19740
tri 4598 19711 4628 19741 nw
rect 4494 19706 4594 19711
tri 4594 19707 4598 19711 nw
rect 4451 19668 4594 19706
rect 4451 19634 4460 19668
rect 4494 19634 4594 19668
tri 4776 19638 4803 19665 se
rect 4803 19638 4855 19891
rect 4451 19596 4594 19634
tri 4769 19631 4776 19638 se
rect 4776 19631 4855 19638
rect 4451 19562 4460 19596
rect 4494 19562 4594 19596
rect 4630 19625 4855 19631
rect 4630 19591 4642 19625
rect 4676 19591 4726 19625
rect 4760 19591 4809 19625
rect 4843 19591 4855 19625
rect 4630 19585 4855 19591
rect 4893 20002 4899 20036
rect 4933 20002 4945 20036
rect 4893 19964 4945 20002
rect 4893 19930 4899 19964
rect 4933 19930 4945 19964
rect 4893 19891 4945 19930
rect 4893 19886 4899 19891
rect 4933 19886 4945 19891
rect 4893 19822 4945 19834
rect 5187 20022 5196 20056
rect 5230 20022 5239 20056
rect 5187 19982 5239 20022
rect 5187 19948 5196 19982
rect 5230 19948 5239 19982
rect 5187 19908 5239 19948
rect 5187 19874 5196 19908
rect 5230 19874 5239 19908
rect 5187 19834 5239 19874
rect 5187 19800 5196 19834
rect 5230 19800 5239 19834
rect 5187 19788 5239 19800
rect 5443 23637 5495 23649
rect 5443 23603 5452 23637
rect 5486 23603 5495 23637
rect 5443 23564 5495 23603
rect 5443 23530 5452 23564
rect 5486 23530 5495 23564
rect 5443 23491 5495 23530
rect 5443 23457 5452 23491
rect 5486 23457 5495 23491
rect 5443 23418 5495 23457
rect 5443 23384 5452 23418
rect 5486 23384 5495 23418
rect 5443 23345 5495 23384
rect 5443 23311 5452 23345
rect 5486 23311 5495 23345
rect 5443 23272 5495 23311
rect 5443 23238 5452 23272
rect 5486 23238 5495 23272
rect 5443 23199 5495 23238
rect 5443 23165 5452 23199
rect 5486 23165 5495 23199
rect 5443 23126 5495 23165
rect 5443 23092 5452 23126
rect 5486 23092 5495 23126
rect 5443 23053 5495 23092
rect 5443 23019 5452 23053
rect 5486 23019 5495 23053
rect 5443 22980 5495 23019
rect 5443 22946 5452 22980
rect 5486 22946 5495 22980
rect 5443 22907 5495 22946
rect 5443 22873 5452 22907
rect 5486 22873 5495 22907
rect 5443 22834 5495 22873
rect 5443 22800 5452 22834
rect 5486 22800 5495 22834
rect 5443 22761 5495 22800
rect 5443 22727 5452 22761
rect 5486 22727 5495 22761
rect 5443 22688 5495 22727
rect 5443 22654 5452 22688
rect 5486 22654 5495 22688
rect 5443 22615 5495 22654
rect 5443 22581 5452 22615
rect 5486 22581 5495 22615
rect 5443 22542 5495 22581
rect 5443 22524 5452 22542
rect 5486 22524 5495 22542
rect 5443 22469 5495 22472
rect 5443 22460 5452 22469
rect 5486 22460 5495 22469
rect 5443 22396 5495 22408
rect 5443 22362 5452 22396
rect 5486 22362 5495 22396
rect 5443 22323 5495 22362
rect 5443 22289 5452 22323
rect 5486 22289 5495 22323
rect 5443 22250 5495 22289
rect 5443 22216 5452 22250
rect 5486 22216 5495 22250
rect 5443 22177 5495 22216
rect 5443 22143 5452 22177
rect 5486 22143 5495 22177
rect 5443 22104 5495 22143
rect 5443 22070 5452 22104
rect 5486 22070 5495 22104
rect 5443 22031 5495 22070
rect 5443 21997 5452 22031
rect 5486 21997 5495 22031
rect 5443 21958 5495 21997
rect 5443 21924 5452 21958
rect 5486 21924 5495 21958
rect 5443 21885 5495 21924
rect 5443 21851 5452 21885
rect 5486 21851 5495 21885
rect 5443 21812 5495 21851
rect 5443 21778 5452 21812
rect 5486 21778 5495 21812
rect 5443 21739 5495 21778
rect 5443 21705 5452 21739
rect 5486 21705 5495 21739
rect 5443 21666 5495 21705
rect 5443 21632 5452 21666
rect 5486 21632 5495 21666
rect 5443 21593 5495 21632
rect 5443 21559 5452 21593
rect 5486 21559 5495 21593
rect 5443 21520 5495 21559
rect 5443 21486 5452 21520
rect 5486 21486 5495 21520
rect 5443 21447 5495 21486
rect 5443 21413 5452 21447
rect 5486 21413 5495 21447
rect 5443 21374 5495 21413
rect 5443 21340 5452 21374
rect 5486 21340 5495 21374
rect 5443 21301 5495 21340
rect 5443 21267 5452 21301
rect 5486 21267 5495 21301
rect 5443 21228 5495 21267
rect 5443 21194 5452 21228
rect 5486 21194 5495 21228
rect 5443 21155 5495 21194
rect 5443 21121 5452 21155
rect 5486 21121 5495 21155
rect 5443 21082 5495 21121
rect 5443 21048 5452 21082
rect 5486 21048 5495 21082
rect 5443 21009 5495 21048
rect 5443 20975 5452 21009
rect 5486 20975 5495 21009
rect 5443 20936 5495 20975
rect 5443 20902 5452 20936
rect 5486 20902 5495 20936
rect 5443 20863 5495 20902
rect 5443 20829 5452 20863
rect 5486 20829 5495 20863
rect 5443 20790 5495 20829
rect 5443 20756 5452 20790
rect 5486 20756 5495 20790
rect 5443 20717 5495 20756
rect 5443 20683 5452 20717
rect 5486 20683 5495 20717
rect 5443 20644 5495 20683
rect 5443 20610 5452 20644
rect 5486 20610 5495 20644
rect 5443 20571 5495 20610
rect 5443 20537 5452 20571
rect 5486 20537 5495 20571
rect 5443 20498 5495 20537
rect 5443 20464 5452 20498
rect 5486 20464 5495 20498
rect 5443 20425 5495 20464
rect 5443 20391 5452 20425
rect 5486 20391 5495 20425
rect 5443 20352 5495 20391
rect 5443 20318 5452 20352
rect 5486 20318 5495 20352
rect 5443 20278 5495 20318
rect 5443 20244 5452 20278
rect 5486 20244 5495 20278
rect 5849 23646 5858 23680
rect 5892 23646 5901 23680
rect 5849 23608 5901 23646
rect 5849 23574 5858 23608
rect 5892 23574 5901 23608
rect 5849 23536 5901 23574
rect 5849 23502 5858 23536
rect 5892 23502 5901 23536
rect 5849 23464 5901 23502
rect 5849 23430 5858 23464
rect 5892 23430 5901 23464
rect 5849 23392 5901 23430
rect 5849 23358 5858 23392
rect 5892 23358 5901 23392
rect 5849 23320 5901 23358
rect 5849 23286 5858 23320
rect 5892 23286 5901 23320
rect 5849 23248 5901 23286
rect 5849 23214 5858 23248
rect 5892 23214 5901 23248
rect 5849 23176 5901 23214
rect 5849 23142 5858 23176
rect 5892 23142 5901 23176
rect 5849 23104 5901 23142
rect 5849 23070 5858 23104
rect 5892 23070 5901 23104
rect 5849 23032 5901 23070
rect 5849 22998 5858 23032
rect 5892 22998 5901 23032
rect 5849 22960 5901 22998
rect 5849 22926 5858 22960
rect 5892 22926 5901 22960
rect 5849 22888 5901 22926
rect 5849 22854 5858 22888
rect 5892 22854 5901 22888
rect 5849 22816 5901 22854
rect 5849 22782 5858 22816
rect 5892 22782 5901 22816
rect 5849 22744 5901 22782
rect 5849 22710 5858 22744
rect 5892 22710 5901 22744
rect 5849 22672 5901 22710
rect 5849 22638 5858 22672
rect 5892 22638 5901 22672
rect 5849 22600 5901 22638
rect 5849 22566 5858 22600
rect 5892 22566 5901 22600
rect 5849 22528 5901 22566
rect 5849 22494 5858 22528
rect 5892 22494 5901 22528
rect 5849 22456 5901 22494
rect 5849 22422 5858 22456
rect 5892 22422 5901 22456
rect 5849 22384 5901 22422
rect 5849 22350 5858 22384
rect 5892 22350 5901 22384
rect 5849 22311 5901 22350
rect 5849 22277 5858 22311
rect 5892 22277 5901 22311
rect 7618 22285 7624 22337
rect 7676 22285 7688 22337
rect 7740 22285 7746 22337
rect 5849 22238 5901 22277
rect 5849 22204 5858 22238
rect 5892 22204 5901 22238
rect 7486 22205 7492 22257
rect 7544 22205 7556 22257
rect 7608 22205 7614 22257
rect 5849 22165 5901 22204
rect 5849 22131 5858 22165
rect 5892 22131 5901 22165
rect 5849 22092 5901 22131
rect 7306 22125 7312 22177
rect 7364 22125 7376 22177
rect 7428 22125 7434 22177
rect 5849 22058 5858 22092
rect 5892 22058 5901 22092
rect 5849 22019 5901 22058
rect 5849 21985 5858 22019
rect 5892 21985 5901 22019
rect 5849 21946 5901 21985
rect 5849 21912 5858 21946
rect 5892 21912 5901 21946
rect 5849 21873 5901 21912
rect 5849 21839 5858 21873
rect 5892 21839 5901 21873
rect 5849 21800 5901 21839
rect 5849 21766 5858 21800
rect 5892 21766 5901 21800
rect 5849 21727 5901 21766
rect 5849 21693 5858 21727
rect 5892 21693 5901 21727
rect 5849 21654 5901 21693
rect 5849 21620 5858 21654
rect 5892 21620 5901 21654
rect 5849 21581 5901 21620
rect 5849 21547 5858 21581
rect 5892 21547 5901 21581
rect 5849 21519 5901 21547
rect 7328 22034 7690 22040
rect 7328 22000 7340 22034
rect 7374 22000 7412 22034
rect 7446 22000 7572 22034
rect 7606 22000 7644 22034
rect 7678 22000 7690 22034
rect 7328 21994 7690 22000
tri 5901 21519 5926 21544 sw
tri 7303 21519 7328 21544 se
rect 7328 21525 7376 21994
tri 7376 21960 7410 21994 nw
tri 7452 21960 7486 21994 ne
rect 7486 21886 7532 21994
tri 7532 21960 7566 21994 nw
tri 7608 21960 7642 21994 ne
tri 7376 21525 7410 21559 sw
tri 7452 21525 7486 21559 se
rect 7486 21525 7532 21644
tri 7532 21525 7566 21559 sw
tri 7608 21525 7642 21559 se
rect 7642 21525 7690 21994
rect 7328 21519 7690 21525
rect 5849 21510 5926 21519
tri 5926 21510 5935 21519 sw
tri 7294 21510 7303 21519 se
rect 7303 21510 7342 21519
rect 5849 21508 7342 21510
rect 5849 21474 5858 21508
rect 5892 21485 7342 21508
rect 7376 21485 7417 21519
rect 7451 21485 7492 21519
rect 7526 21485 7567 21519
rect 7601 21485 7642 21519
rect 7676 21485 7690 21519
rect 5892 21474 7690 21485
rect 5849 21454 7690 21474
rect 5849 21435 5901 21454
rect 5849 21401 5858 21435
rect 5892 21401 5901 21435
tri 5901 21420 5935 21454 nw
rect 5849 21362 5901 21401
rect 5849 21328 5858 21362
rect 5892 21328 5901 21362
rect 5849 21289 5901 21328
rect 5849 21255 5858 21289
rect 5892 21255 5901 21289
rect 5849 21216 5901 21255
rect 5849 21182 5858 21216
rect 5892 21182 5901 21216
rect 5849 21143 5901 21182
rect 5849 21109 5858 21143
rect 5892 21109 5901 21143
rect 5849 21070 5901 21109
rect 5849 21036 5858 21070
rect 5892 21036 5901 21070
rect 5849 20997 5901 21036
rect 5849 20963 5858 20997
rect 5892 20963 5901 20997
rect 5849 20924 5901 20963
rect 5849 20890 5858 20924
rect 5892 20890 5901 20924
rect 5849 20851 5901 20890
rect 5849 20817 5858 20851
rect 5892 20817 5901 20851
rect 5849 20778 5901 20817
rect 5849 20744 5858 20778
rect 5892 20744 5901 20778
rect 5849 20705 5901 20744
rect 5849 20671 5858 20705
rect 5892 20671 5901 20705
rect 5849 20632 5901 20671
rect 5849 20598 5858 20632
rect 5892 20598 5901 20632
rect 5849 20559 5901 20598
rect 5849 20525 5858 20559
rect 5892 20525 5901 20559
rect 5849 20486 5901 20525
rect 5849 20452 5858 20486
rect 5892 20452 5901 20486
rect 5849 20413 5901 20452
rect 5849 20379 5858 20413
rect 5892 20379 5901 20413
rect 5849 20340 5901 20379
rect 5849 20306 5858 20340
rect 5892 20306 5901 20340
rect 5849 20267 5901 20306
rect 5443 20204 5495 20244
rect 5443 20170 5452 20204
rect 5486 20170 5495 20204
rect 5443 20130 5495 20170
rect 5443 20096 5452 20130
rect 5486 20096 5495 20130
rect 5443 20056 5495 20096
rect 5443 20022 5452 20056
rect 5486 20022 5495 20056
rect 5443 19982 5495 20022
rect 5443 19948 5452 19982
rect 5486 19948 5495 19982
rect 5443 19908 5495 19948
rect 5443 19874 5452 19908
rect 5486 19874 5495 19908
rect 5443 19834 5495 19874
rect 5443 19800 5452 19834
rect 5486 19800 5495 19834
rect 5443 19788 5495 19800
rect 5699 20253 5751 20259
rect 5699 20189 5751 20201
rect 4893 19745 4945 19770
rect 4893 19711 4899 19745
rect 4933 19711 4945 19745
rect 4893 19672 4945 19711
rect 4893 19638 4899 19672
rect 4933 19638 4945 19672
rect 4893 19599 4945 19638
rect 4451 19524 4594 19562
rect 4451 19490 4460 19524
rect 4494 19492 4594 19524
rect 4893 19565 4899 19599
rect 4933 19565 4945 19599
rect 4893 19526 4945 19565
tri 4594 19492 4611 19509 sw
rect 4893 19492 4899 19526
rect 4933 19492 4945 19526
rect 4494 19490 4611 19492
rect 4451 19480 4611 19490
tri 4611 19480 4623 19492 sw
rect 4893 19480 4945 19492
rect 5074 19700 5152 19706
rect 5074 19666 5086 19700
rect 5120 19666 5152 19700
rect 5074 19628 5152 19666
rect 5074 19594 5086 19628
rect 5120 19594 5152 19628
rect 4451 19475 4623 19480
tri 4623 19475 4628 19480 sw
rect 4451 19469 4855 19475
rect 4451 19452 4585 19469
rect 4451 19418 4460 19452
rect 4494 19435 4585 19452
rect 4619 19435 4660 19469
rect 4694 19435 4735 19469
rect 4769 19435 4809 19469
rect 4843 19435 4855 19469
rect 4494 19429 4855 19435
rect 4494 19418 4503 19429
rect 4451 19380 4503 19418
tri 4503 19395 4537 19429 nw
rect 4451 19346 4460 19380
rect 4494 19346 4503 19380
rect 4451 19308 4503 19346
rect 4451 19274 4460 19308
rect 4494 19274 4503 19308
rect 4451 19236 4503 19274
rect 4451 19202 4460 19236
rect 4494 19202 4503 19236
rect 4451 19164 4503 19202
rect 4451 19130 4460 19164
rect 4494 19130 4503 19164
rect 5074 19271 5152 19594
rect 5350 19700 5514 19706
rect 5350 19666 5362 19700
rect 5396 19666 5461 19700
rect 5350 19648 5461 19666
rect 5513 19648 5514 19700
rect 5350 19636 5514 19648
rect 5350 19628 5461 19636
rect 5350 19594 5362 19628
rect 5396 19594 5461 19628
rect 5350 19584 5461 19594
rect 5513 19584 5514 19636
rect 5350 19578 5514 19584
rect 5074 19219 5080 19271
rect 5132 19219 5152 19271
rect 5074 19207 5152 19219
rect 5074 19155 5080 19207
rect 5132 19155 5152 19207
rect 4451 19092 4503 19130
tri 5690 19099 5699 19108 se
rect 5699 19099 5751 20137
rect 4451 19058 4460 19092
rect 4494 19058 4503 19092
tri 5665 19074 5690 19099 se
rect 5690 19074 5751 19099
rect 4451 19020 4503 19058
rect 5068 19068 5751 19074
rect 5068 19034 5080 19068
rect 5114 19034 5152 19068
rect 5186 19034 5751 19068
rect 5068 19028 5751 19034
rect 5849 20233 5858 20267
rect 5892 20233 5901 20267
rect 5849 20194 5901 20233
rect 5849 20160 5858 20194
rect 5892 20160 5901 20194
rect 5849 20121 5901 20160
rect 8223 20253 8351 30469
rect 9567 30128 9619 30134
rect 9567 30064 9619 30076
rect 9456 30048 9508 30054
rect 9456 29984 9508 29996
rect 9300 29968 9352 29974
rect 9300 29904 9352 29916
tri 9266 22337 9300 22371 se
rect 9300 22337 9352 29852
rect 9224 22285 9230 22337
rect 9282 22285 9294 22337
rect 9346 22285 9352 22337
tri 9450 22285 9456 22291 se
rect 9456 22285 9508 29932
tri 9422 22257 9450 22285 se
rect 9450 22257 9508 22285
rect 9380 22205 9386 22257
rect 9438 22205 9450 22257
rect 9502 22205 9508 22257
rect 9567 22171 9619 30012
rect 9567 22107 9619 22119
rect 9567 22049 9619 22055
rect 8275 20201 8299 20253
rect 8223 20189 8351 20201
rect 8275 20137 8299 20189
rect 8223 20131 8351 20137
rect 5849 20087 5858 20121
rect 5892 20087 5901 20121
rect 5849 20048 5901 20087
rect 5849 20014 5858 20048
rect 5892 20014 5901 20048
rect 5849 19975 5901 20014
rect 5849 19941 5858 19975
rect 5892 19941 5901 19975
rect 5849 19902 5901 19941
rect 5849 19868 5858 19902
rect 5892 19868 5901 19902
rect 5849 19829 5901 19868
rect 5849 19795 5858 19829
rect 5892 19795 5901 19829
rect 5849 19756 5901 19795
rect 5849 19722 5858 19756
rect 5892 19722 5901 19756
rect 5849 19683 5901 19722
rect 5849 19649 5858 19683
rect 5892 19649 5901 19683
rect 5849 19610 5901 19649
rect 5849 19576 5858 19610
rect 5892 19576 5901 19610
rect 5849 19537 5901 19576
rect 5849 19503 5858 19537
rect 5892 19503 5901 19537
rect 5849 19464 5901 19503
rect 5849 19430 5858 19464
rect 5892 19430 5901 19464
rect 5849 19391 5901 19430
rect 5849 19357 5858 19391
rect 5892 19357 5901 19391
rect 5849 19318 5901 19357
rect 5849 19284 5858 19318
rect 5892 19284 5901 19318
rect 5849 19245 5901 19284
rect 5849 19211 5858 19245
rect 5892 19211 5901 19245
rect 5849 19172 5901 19211
rect 5849 19138 5858 19172
rect 5892 19138 5901 19172
rect 5849 19099 5901 19138
rect 5849 19065 5858 19099
rect 5892 19065 5901 19099
rect 4451 18986 4460 19020
rect 4494 18986 4503 19020
rect 5849 19026 5901 19065
rect 4451 18948 4503 18986
rect 4451 18914 4460 18948
rect 4494 18914 4503 18948
rect 4451 18876 4503 18914
rect 4451 18842 4460 18876
rect 4494 18842 4503 18876
rect 4451 18804 4503 18842
rect 4451 18770 4460 18804
rect 4494 18770 4503 18804
rect 4987 18996 5039 19002
rect 5849 18992 5858 19026
rect 5892 18992 5901 19026
rect 4987 18932 5039 18944
rect 4987 18770 5039 18880
rect 5247 18816 5299 18972
rect 4451 18732 4503 18770
rect 4451 18698 4460 18732
rect 4494 18698 4503 18732
rect 4451 18660 4503 18698
rect 5247 18752 5299 18764
rect 5247 18694 5299 18700
rect 5849 18953 5901 18992
rect 5849 18919 5858 18953
rect 5892 18919 5901 18953
rect 5849 18880 5901 18919
rect 5849 18846 5858 18880
rect 5892 18846 5901 18880
rect 5849 18807 5901 18846
rect 5849 18773 5858 18807
rect 5892 18773 5901 18807
rect 5849 18734 5901 18773
rect 5849 18700 5858 18734
rect 5892 18700 5901 18734
rect 4451 18626 4460 18660
rect 4494 18626 4503 18660
rect 4451 18588 4503 18626
rect 4451 18554 4460 18588
rect 4494 18554 4503 18588
rect 5849 18661 5901 18700
rect 5849 18627 5858 18661
rect 5892 18627 5901 18661
rect 5849 18588 5901 18627
tri 4503 18554 4505 18556 sw
tri 5847 18554 5849 18556 se
rect 5849 18554 5858 18588
rect 5892 18554 5901 18588
rect 3926 18476 4192 18528
rect 4451 18522 4505 18554
tri 4505 18522 4537 18554 sw
tri 5815 18522 5847 18554 se
rect 5847 18522 5901 18554
rect 4451 18516 5901 18522
rect 4451 18482 4532 18516
rect 4566 18482 4606 18516
rect 4640 18482 4680 18516
rect 4714 18482 4754 18516
rect 4788 18482 4828 18516
rect 4862 18482 4902 18516
rect 4936 18482 4976 18516
rect 5010 18482 5050 18516
rect 5084 18482 5124 18516
rect 5158 18482 5198 18516
rect 5232 18482 5272 18516
rect 5306 18482 5346 18516
rect 5380 18482 5420 18516
rect 5454 18482 5493 18516
rect 5527 18482 5566 18516
rect 5600 18482 5639 18516
rect 5673 18482 5712 18516
rect 5746 18482 5785 18516
rect 5819 18482 5901 18516
rect 4451 18476 5901 18482
rect 8793 19971 8799 20023
rect 8851 19971 8863 20023
rect 8915 19971 8921 20023
rect 2996 18409 3048 18421
rect 2996 18351 3048 18357
rect 2627 17723 2633 17775
rect 2685 17723 2730 17775
rect 2782 17723 2788 17775
rect 2627 17699 2788 17723
rect 2627 17647 2633 17699
rect 2685 17647 2730 17699
rect 2782 17647 2788 17699
rect 2816 18289 3709 18298
rect 2816 18255 2899 18289
rect 2933 18255 2977 18289
rect 3011 18255 3055 18289
rect 3089 18255 3133 18289
rect 3167 18255 3211 18289
rect 3245 18255 3289 18289
rect 3323 18255 3367 18289
rect 3401 18255 3445 18289
rect 3479 18255 3523 18289
rect 3557 18255 3601 18289
rect 3635 18255 3679 18289
rect 2816 18246 3709 18255
rect 3761 18246 3776 18298
rect 3828 18246 3843 18298
rect 3895 18246 3910 18298
rect 3962 18289 3977 18298
rect 4029 18289 4044 18298
rect 4096 18289 4111 18298
rect 4163 18289 4178 18298
rect 4230 18289 4245 18298
rect 4297 18289 4312 18298
rect 4364 18289 4379 18298
rect 4431 18289 4445 18298
rect 4497 18289 6790 18298
rect 3967 18255 3977 18289
rect 4039 18255 4044 18289
rect 4364 18255 4365 18289
rect 4431 18255 4437 18289
rect 4497 18255 4509 18289
rect 4543 18255 4581 18289
rect 4615 18255 4653 18289
rect 4687 18255 4725 18289
rect 4759 18255 4797 18289
rect 4831 18255 4869 18289
rect 4903 18255 4941 18289
rect 4975 18255 5013 18289
rect 5047 18255 5085 18289
rect 5119 18255 5157 18289
rect 5191 18255 5229 18289
rect 5263 18255 5301 18289
rect 5335 18255 5373 18289
rect 5407 18255 5445 18289
rect 5479 18255 5517 18289
rect 5551 18255 5589 18289
rect 5623 18255 5661 18289
rect 5695 18255 5733 18289
rect 5767 18255 5805 18289
rect 5839 18255 5877 18289
rect 5911 18255 5949 18289
rect 5983 18255 6021 18289
rect 6055 18255 6094 18289
rect 6128 18255 6167 18289
rect 6201 18255 6240 18289
rect 6274 18255 6313 18289
rect 6347 18255 6386 18289
rect 6420 18255 6459 18289
rect 6493 18255 6532 18289
rect 6566 18255 6605 18289
rect 6639 18255 6678 18289
rect 6712 18255 6790 18289
rect 3962 18246 3977 18255
rect 4029 18246 4044 18255
rect 4096 18246 4111 18255
rect 4163 18246 4178 18255
rect 4230 18246 4245 18255
rect 4297 18246 4312 18255
rect 4364 18246 4379 18255
rect 4431 18246 4445 18255
rect 4497 18246 6790 18255
rect 2816 18217 2866 18246
rect 2816 18183 2822 18217
rect 2856 18216 2866 18217
tri 2866 18216 2896 18246 nw
tri 6710 18216 6740 18246 ne
rect 6740 18216 6790 18246
rect 2856 18183 2862 18216
tri 2862 18212 2866 18216 nw
tri 6740 18212 6744 18216 ne
rect 2816 18143 2862 18183
rect 2816 18109 2822 18143
rect 2856 18109 2862 18143
rect 2816 18069 2862 18109
rect 2816 18035 2822 18069
rect 2856 18035 2862 18069
rect 2816 17995 2862 18035
rect 2816 17961 2822 17995
rect 2856 17961 2862 17995
rect 2816 17921 2862 17961
rect 2816 17887 2822 17921
rect 2856 17887 2862 17921
rect 2816 17847 2862 17887
rect 2816 17813 2822 17847
rect 2856 17813 2862 17847
rect 2816 17774 2862 17813
rect 2816 17740 2822 17774
rect 2856 17740 2862 17774
rect 2816 17701 2862 17740
rect 2816 17667 2822 17701
rect 2856 17667 2862 17701
rect 2288 17567 2294 17619
rect 2346 17567 2391 17619
rect 2443 17567 2449 17619
rect 2288 17543 2449 17567
rect 2288 17491 2294 17543
rect 2346 17491 2391 17543
rect 2443 17491 2449 17543
rect 2816 17628 2862 17667
rect 2816 17594 2822 17628
rect 2856 17594 2862 17628
rect 2816 17555 2862 17594
rect 2816 17521 2822 17555
rect 2856 17521 2862 17555
rect 2816 17482 2862 17521
rect 2816 17448 2822 17482
rect 2856 17448 2862 17482
rect 2816 17409 2862 17448
rect 2816 17375 2822 17409
rect 2856 17375 2862 17409
rect 2816 17336 2862 17375
rect 2816 17302 2822 17336
rect 2856 17302 2862 17336
rect 2816 17263 2862 17302
rect 2816 17229 2822 17263
rect 2856 17229 2862 17263
rect 2816 17190 2862 17229
rect 2816 17156 2822 17190
rect 2856 17156 2862 17190
rect 2816 17117 2862 17156
rect 2816 17083 2822 17117
rect 2856 17083 2862 17117
rect 2816 17044 2862 17083
rect 2816 17010 2822 17044
rect 2856 17010 2862 17044
rect 2816 16971 2862 17010
rect 2816 16937 2822 16971
rect 2856 16937 2862 16971
tri 1287 16901 1290 16904 sw
rect 1187 16898 1290 16901
tri 1290 16898 1293 16901 sw
rect 2816 16898 2862 16937
rect 1187 16876 1293 16898
tri 1293 16876 1315 16898 sw
rect 1187 16824 1193 16876
rect 1245 16824 1257 16876
rect 1309 16824 1315 16876
rect 1187 16426 1287 16824
tri 1287 16796 1315 16824 nw
rect 2816 16864 2822 16898
rect 2856 16864 2862 16898
rect 2816 16825 2862 16864
rect 2816 16791 2822 16825
rect 2856 16791 2862 16825
rect 2816 16752 2862 16791
rect 2816 16718 2822 16752
rect 2856 16718 2862 16752
rect 2816 16679 2862 16718
rect 2816 16645 2822 16679
rect 2856 16645 2862 16679
rect 2816 16606 2862 16645
rect 2816 16572 2822 16606
rect 2856 16572 2862 16606
rect 2816 16533 2862 16572
rect 2816 16499 2822 16533
rect 2856 16499 2862 16533
rect 2816 16460 2862 16499
tri 1287 16426 1309 16448 sw
rect 2816 16426 2822 16460
rect 2856 16426 2862 16460
rect 1187 16424 1309 16426
tri 1309 16424 1311 16426 sw
rect 1187 16420 1311 16424
tri 1311 16420 1315 16424 sw
rect 1187 16368 1193 16420
rect 1245 16368 1257 16420
rect 1309 16368 1315 16420
rect 2816 16387 2862 16426
rect 2816 16353 2822 16387
rect 2856 16353 2862 16387
rect 2816 16314 2862 16353
rect 2816 16280 2822 16314
rect 2856 16280 2862 16314
rect 2816 16241 2862 16280
rect 2816 16207 2822 16241
rect 2856 16207 2862 16241
rect 2816 16168 2862 16207
rect 2816 16134 2822 16168
rect 2856 16134 2862 16168
rect 2816 16095 2862 16134
rect 2816 16061 2822 16095
rect 2856 16061 2862 16095
rect 2816 16022 2862 16061
rect 2816 15988 2822 16022
rect 2856 15988 2862 16022
rect 2816 15949 2862 15988
rect 2816 15915 2822 15949
rect 2856 15915 2862 15949
rect 2816 15876 2862 15915
rect 2996 18202 3048 18208
rect 2996 18138 3048 18150
rect 2996 17453 3048 18086
rect 6744 18182 6750 18216
rect 6784 18182 6790 18216
rect 6744 18143 6790 18182
rect 6744 18109 6750 18143
rect 6784 18109 6790 18143
rect 6744 18070 6790 18109
rect 6744 18036 6750 18070
rect 6784 18036 6790 18070
rect 2996 17389 3048 17401
rect 2996 16006 3048 17337
rect 2996 15942 3048 15954
rect 2996 15884 3048 15890
rect 3076 18029 6516 18035
rect 3076 17995 3161 18029
rect 3195 17995 3240 18029
rect 3274 17995 3319 18029
rect 3353 17995 3398 18029
rect 3432 17995 3478 18029
rect 3512 17995 3558 18029
rect 3592 17995 3638 18029
rect 3672 17995 3718 18029
rect 3752 17995 3798 18029
rect 3832 17995 3908 18029
rect 3942 17995 3981 18029
rect 4015 17995 4054 18029
rect 4088 17995 4127 18029
rect 4161 17995 4200 18029
rect 4234 17995 4273 18029
rect 4307 17995 4346 18029
rect 4380 17995 4419 18029
rect 4453 17995 4492 18029
rect 4526 17995 4565 18029
rect 4599 17995 4638 18029
rect 4672 17995 4711 18029
rect 4745 17995 4784 18029
rect 4818 17995 4857 18029
rect 4891 17995 4930 18029
rect 4964 17995 5003 18029
rect 5037 17995 5076 18029
rect 5110 17995 5149 18029
rect 5183 17995 5222 18029
rect 5256 17995 5295 18029
rect 5329 17995 5368 18029
rect 5402 17995 5442 18029
rect 5476 17995 5516 18029
rect 5550 17995 5590 18029
rect 5624 17995 5664 18029
rect 5698 17995 5738 18029
rect 5772 17995 5812 18029
rect 5846 17995 5886 18029
rect 5920 17995 5960 18029
rect 5994 17995 6034 18029
rect 6068 17995 6108 18029
rect 6142 17995 6182 18029
rect 6216 17995 6256 18029
rect 6290 17995 6330 18029
rect 6364 17995 6404 18029
rect 6438 17995 6516 18029
rect 3076 17989 6516 17995
rect 3076 17963 3136 17989
tri 3136 17963 3162 17989 nw
tri 6436 17963 6462 17989 ne
rect 6462 17963 6516 17989
rect 3076 17957 3130 17963
tri 3130 17957 3136 17963 nw
tri 6462 17957 6468 17963 ne
rect 6468 17957 6516 17963
rect 3076 17925 3082 17957
rect 3116 17925 3128 17957
tri 3128 17955 3130 17957 nw
tri 6468 17955 6470 17957 ne
rect 3076 17861 3082 17873
rect 3116 17861 3128 17873
rect 3076 17777 3082 17809
rect 3116 17777 3128 17809
rect 3076 17738 3128 17777
rect 3076 17704 3082 17738
rect 3116 17704 3128 17738
rect 3076 17665 3128 17704
rect 3076 17631 3082 17665
rect 3116 17631 3128 17665
rect 3076 17592 3128 17631
rect 3177 17879 3183 17931
rect 3235 17879 3254 17931
rect 3306 17879 3324 17931
rect 3376 17879 3382 17931
rect 3177 17855 3382 17879
rect 3177 17803 3183 17855
rect 3235 17803 3254 17855
rect 3306 17803 3324 17855
rect 3376 17803 3382 17855
rect 3177 17620 3382 17803
rect 3921 17925 4022 17935
rect 3921 17873 3946 17925
rect 3998 17873 4022 17925
rect 3921 17861 4022 17873
rect 3921 17809 3946 17861
rect 3998 17809 4022 17861
tri 3915 17779 3921 17785 se
rect 3921 17779 4022 17809
tri 3914 17778 3915 17779 se
rect 3915 17778 4022 17779
tri 3887 17751 3914 17778 se
rect 3914 17751 4022 17778
rect 3642 17745 4022 17751
rect 3642 17711 3654 17745
rect 3688 17711 3745 17745
rect 3779 17711 3836 17745
rect 3870 17711 4022 17745
rect 3642 17705 4022 17711
tri 3887 17682 3910 17705 ne
rect 3910 17682 4022 17705
rect 3540 17670 3592 17682
tri 3910 17671 3921 17682 ne
rect 3540 17636 3552 17670
rect 3586 17636 3592 17670
rect 3076 17558 3082 17592
rect 3116 17558 3128 17592
rect 3076 17519 3128 17558
rect 3076 17485 3082 17519
rect 3116 17485 3128 17519
rect 3076 17446 3128 17485
rect 3076 17412 3082 17446
rect 3116 17412 3128 17446
rect 3076 17373 3128 17412
rect 3076 17339 3082 17373
rect 3116 17339 3128 17373
rect 3076 17300 3128 17339
rect 3076 17266 3082 17300
rect 3116 17266 3128 17300
rect 3076 17227 3128 17266
rect 3076 17193 3082 17227
rect 3116 17193 3128 17227
rect 3076 17154 3128 17193
rect 3076 17120 3082 17154
rect 3116 17120 3128 17154
rect 3076 17081 3128 17120
rect 3076 17047 3082 17081
rect 3116 17047 3128 17081
rect 3076 17008 3128 17047
rect 3076 16974 3082 17008
rect 3116 16974 3128 17008
rect 3076 16935 3128 16974
rect 3076 16901 3082 16935
rect 3116 16901 3128 16935
rect 3076 16862 3128 16901
rect 3076 16828 3082 16862
rect 3116 16828 3128 16862
rect 3076 16789 3128 16828
rect 3076 16755 3082 16789
rect 3116 16755 3128 16789
rect 3076 16716 3128 16755
rect 3076 16682 3082 16716
rect 3116 16682 3128 16716
rect 3076 16643 3128 16682
rect 3076 16609 3082 16643
rect 3116 16609 3128 16643
rect 3076 16570 3128 16609
rect 3076 16536 3082 16570
rect 3116 16536 3128 16570
rect 3076 16497 3128 16536
rect 3076 16463 3082 16497
rect 3116 16463 3128 16497
rect 3076 16424 3128 16463
rect 3076 16390 3082 16424
rect 3116 16390 3128 16424
rect 3076 16351 3128 16390
rect 3076 16317 3082 16351
rect 3116 16317 3128 16351
rect 3076 16278 3128 16317
rect 3076 16244 3082 16278
rect 3116 16244 3128 16278
rect 3076 16205 3128 16244
rect 3076 16171 3082 16205
rect 3116 16171 3128 16205
rect 3076 16132 3128 16171
rect 3076 16098 3082 16132
rect 3116 16098 3128 16132
rect 3076 16059 3128 16098
rect 3435 17613 3487 17619
rect 3435 17549 3487 17561
rect 3435 17495 3444 17497
rect 3478 17495 3487 17497
rect 3435 17455 3487 17495
rect 3435 17421 3444 17455
rect 3478 17421 3487 17455
rect 3435 17381 3487 17421
rect 3435 17347 3444 17381
rect 3478 17347 3487 17381
rect 3435 17306 3487 17347
rect 3435 17272 3444 17306
rect 3478 17272 3487 17306
rect 3435 17231 3487 17272
rect 3435 17197 3444 17231
rect 3478 17197 3487 17231
rect 3435 17156 3487 17197
rect 3435 17122 3444 17156
rect 3478 17122 3487 17156
rect 3540 17589 3592 17636
rect 3540 17555 3552 17589
rect 3586 17555 3592 17589
rect 3540 17508 3592 17555
rect 3540 17474 3552 17508
rect 3586 17474 3592 17508
rect 3540 17453 3592 17474
rect 3540 17393 3552 17401
rect 3586 17393 3592 17401
rect 3540 17389 3592 17393
rect 3540 17311 3552 17337
rect 3586 17311 3592 17337
rect 3540 17263 3592 17311
rect 3540 17229 3552 17263
rect 3586 17229 3592 17263
rect 3620 17589 3774 17595
rect 3620 17555 3654 17589
rect 3688 17555 3728 17589
rect 3762 17555 3774 17589
rect 3620 17549 3774 17555
rect 3620 17525 3682 17549
tri 3682 17525 3706 17549 nw
rect 3620 17522 3679 17525
tri 3679 17522 3682 17525 nw
rect 3620 17457 3672 17522
tri 3672 17515 3679 17522 nw
tri 3900 17452 3921 17473 se
rect 3921 17452 4022 17682
tri 3897 17449 3900 17452 se
rect 3900 17449 4022 17452
tri 3887 17439 3897 17449 se
rect 3897 17439 4022 17449
rect 3620 17393 3672 17405
rect 3700 17433 4022 17439
rect 3700 17399 3712 17433
rect 3746 17399 3786 17433
rect 3820 17399 4022 17433
rect 3700 17393 4022 17399
tri 3887 17379 3901 17393 ne
rect 3901 17379 4022 17393
tri 3901 17376 3904 17379 ne
rect 3904 17376 4022 17379
tri 3904 17359 3921 17376 ne
rect 3620 17306 3672 17341
tri 3672 17306 3683 17317 sw
rect 3620 17303 3683 17306
tri 3683 17303 3686 17306 sw
rect 3620 17283 3686 17303
tri 3686 17283 3706 17303 sw
rect 3620 17277 3774 17283
rect 3620 17243 3654 17277
rect 3688 17243 3728 17277
rect 3762 17243 3774 17277
rect 3620 17237 3774 17243
rect 3540 17181 3592 17229
rect 3540 17147 3552 17181
rect 3586 17147 3592 17181
tri 3920 17160 3921 17161 se
rect 3921 17160 4022 17376
tri 3917 17157 3920 17160 se
rect 3920 17157 4022 17160
rect 3540 17135 3592 17147
tri 3895 17135 3917 17157 se
rect 3917 17135 4022 17157
tri 3887 17127 3895 17135 se
rect 3895 17127 4022 17135
rect 3435 17081 3487 17122
rect 3642 17121 4022 17127
rect 3642 17087 3654 17121
rect 3688 17087 3745 17121
rect 3779 17087 3836 17121
rect 3870 17087 4022 17121
rect 3642 17081 4022 17087
rect 4215 17925 4267 17931
rect 4215 17861 4267 17873
rect 3435 17047 3444 17081
rect 3478 17047 3487 17081
rect 3435 17006 3487 17047
rect 3435 16972 3444 17006
rect 3478 16972 3487 17006
rect 3435 16931 3487 16972
rect 4215 16937 4267 17809
rect 4371 17769 4423 17931
rect 4371 17705 4423 17717
rect 4371 16937 4423 17653
rect 4527 17925 4579 17931
rect 4527 17861 4579 17873
rect 4527 16937 4579 17809
rect 4682 17769 4734 17931
rect 4682 17705 4734 17717
rect 4682 16937 4734 17653
rect 4839 17925 4891 17931
rect 4839 17861 4891 17873
rect 4839 16937 4891 17809
rect 4995 17613 5047 17931
rect 4995 17549 5047 17561
rect 4995 16937 5047 17497
rect 5151 17925 5203 17931
rect 5151 17861 5203 17873
rect 5151 16937 5203 17809
rect 5307 17613 5359 17931
rect 5307 17549 5359 17561
rect 5307 16937 5359 17497
rect 5462 17925 5514 17931
rect 5462 17861 5514 17873
rect 5462 16937 5514 17809
rect 5832 17925 5884 17931
rect 5832 17861 5884 17873
rect 5832 17803 5884 17809
rect 6470 17923 6476 17957
rect 6510 17923 6516 17957
rect 6470 17885 6516 17923
rect 6470 17851 6476 17885
rect 6510 17851 6516 17885
rect 6470 17813 6516 17851
rect 6470 17779 6476 17813
rect 6510 17779 6516 17813
rect 6470 17741 6516 17779
rect 6470 17707 6476 17741
rect 6510 17707 6516 17741
rect 6470 17668 6516 17707
rect 6470 17634 6476 17668
rect 6510 17634 6516 17668
rect 6470 17595 6516 17634
rect 6470 17561 6476 17595
rect 6510 17561 6516 17595
rect 6470 17522 6516 17561
rect 6470 17488 6476 17522
rect 6510 17488 6516 17522
rect 6470 17449 6516 17488
rect 6470 17415 6476 17449
rect 6510 17415 6516 17449
rect 6470 17376 6516 17415
rect 6470 17342 6476 17376
rect 6510 17342 6516 17376
rect 6470 17303 6516 17342
rect 6470 17269 6476 17303
rect 6510 17269 6516 17303
rect 6470 17230 6516 17269
rect 6470 17196 6476 17230
rect 6510 17196 6516 17230
rect 6470 17157 6516 17196
rect 6470 17123 6476 17157
rect 6510 17123 6516 17157
rect 6470 17084 6516 17123
rect 6470 17050 6476 17084
rect 6510 17050 6516 17084
tri 6454 17014 6470 17030 se
rect 6470 17014 6516 17050
tri 6451 17011 6454 17014 se
rect 6454 17011 6516 17014
tri 6436 16996 6451 17011 se
rect 6451 16996 6476 17011
rect 6211 16977 6476 16996
rect 6510 16977 6516 17011
rect 6211 16964 6516 16977
rect 3435 16897 3444 16931
rect 3478 16897 3487 16931
rect 3435 16856 3487 16897
rect 6211 16930 6237 16964
rect 6271 16930 6309 16964
rect 6343 16938 6516 16964
rect 6343 16930 6476 16938
rect 6211 16904 6476 16930
rect 6510 16904 6516 16938
rect 6211 16891 6516 16904
rect 3435 16822 3444 16856
rect 3478 16822 3487 16856
rect 4302 16867 4383 16876
rect 4302 16833 4314 16867
rect 4348 16833 4383 16867
rect 4302 16824 4383 16833
rect 4435 16824 4447 16876
rect 4499 16867 4798 16876
rect 4499 16833 4533 16867
rect 4567 16833 4606 16867
rect 4640 16833 4679 16867
rect 4713 16833 4752 16867
rect 4786 16833 4798 16867
rect 4499 16824 4798 16833
rect 4946 16867 5417 16873
rect 4946 16833 4958 16867
rect 4992 16833 5041 16867
rect 5075 16833 5124 16867
rect 5158 16833 5207 16867
rect 5241 16833 5289 16867
rect 5323 16833 5371 16867
rect 5405 16833 5417 16867
rect 4946 16827 5417 16833
rect 6211 16857 6237 16891
rect 6271 16857 6309 16891
rect 6343 16865 6516 16891
rect 6343 16857 6476 16865
rect 6211 16831 6476 16857
rect 6510 16831 6516 16865
tri 5016 16824 5019 16827 ne
rect 5019 16824 5203 16827
rect 3435 16781 3487 16822
tri 5019 16818 5025 16824 ne
rect 5025 16818 5203 16824
tri 5203 16818 5212 16827 nw
rect 6211 16818 6516 16831
tri 5025 16793 5050 16818 ne
rect 3435 16747 3444 16781
rect 3478 16747 3487 16781
rect 3435 16706 3487 16747
rect 5050 16792 5178 16818
tri 5178 16793 5203 16818 nw
rect 3435 16672 3444 16706
rect 3478 16672 3487 16706
rect 3435 16631 3487 16672
rect 3435 16597 3444 16631
rect 3478 16597 3487 16631
rect 3435 16556 3487 16597
rect 3435 16522 3444 16556
rect 3478 16522 3487 16556
rect 3435 16481 3487 16522
rect 3435 16447 3444 16481
rect 3478 16447 3487 16481
rect 3435 16406 3487 16447
rect 3435 16372 3444 16406
rect 3478 16372 3487 16406
rect 3435 16331 3487 16372
rect 3435 16297 3444 16331
rect 3478 16297 3487 16331
rect 3435 16256 3487 16297
rect 3435 16222 3444 16256
rect 3478 16222 3487 16256
rect 3435 16181 3487 16222
rect 3435 16147 3444 16181
rect 3478 16147 3487 16181
rect 3435 16106 3487 16147
rect 3435 16072 3444 16106
rect 3478 16072 3487 16106
rect 3435 16060 3487 16072
rect 3715 16711 3833 16743
rect 5050 16740 5056 16792
rect 5108 16740 5120 16792
rect 5172 16740 5178 16792
rect 6211 16784 6237 16818
rect 6271 16784 6309 16818
rect 6343 16792 6516 16818
rect 6343 16784 6476 16792
rect 6211 16758 6476 16784
rect 6510 16758 6516 16792
rect 6211 16745 6516 16758
rect 3715 16101 3721 16711
rect 3827 16101 3833 16711
rect 6211 16711 6237 16745
rect 6271 16711 6309 16745
rect 6343 16719 6516 16745
rect 6343 16711 6476 16719
rect 4180 16652 4232 16689
rect 4180 16588 4232 16600
rect 4180 16127 4232 16536
rect 4878 16368 4884 16420
rect 4936 16368 4948 16420
rect 5000 16368 5006 16420
tri 4870 16127 4878 16135 se
rect 4878 16127 5006 16368
tri 4864 16121 4870 16127 se
rect 4870 16121 5006 16127
tri 5006 16121 5020 16135 sw
tri 4844 16101 4864 16121 se
rect 4864 16101 5020 16121
tri 5020 16101 5040 16121 sw
rect 3715 16062 3833 16101
rect 3076 16025 3082 16059
rect 3116 16025 3128 16059
rect 3076 15986 3128 16025
rect 3715 16028 3721 16062
rect 3755 16028 3793 16062
rect 3827 16028 3833 16062
rect 4270 16095 5788 16101
rect 4270 16061 4282 16095
rect 4316 16061 4355 16095
rect 4389 16061 4428 16095
rect 4462 16061 4501 16095
rect 4535 16061 4574 16095
rect 4608 16061 4647 16095
rect 4681 16061 4720 16095
rect 4754 16061 4793 16095
rect 4827 16061 4866 16095
rect 4900 16061 4939 16095
rect 4973 16061 5012 16095
rect 5046 16061 5085 16095
rect 5119 16061 5158 16095
rect 5192 16061 5231 16095
rect 5265 16061 5304 16095
rect 5338 16061 5377 16095
rect 5411 16061 5450 16095
rect 5484 16061 5523 16095
rect 5557 16061 5596 16095
rect 5630 16061 5669 16095
rect 5703 16061 5742 16095
rect 5776 16061 5788 16095
rect 4270 16055 5788 16061
tri 4844 16047 4852 16055 ne
rect 4852 16047 5032 16055
tri 5032 16047 5040 16055 nw
tri 4852 16028 4871 16047 ne
rect 4871 16028 5013 16047
tri 5013 16028 5032 16047 nw
rect 3076 15952 3082 15986
rect 3116 15952 3128 15986
rect 3180 15960 3234 16012
rect 3286 15960 3298 16012
rect 3350 15960 3382 16012
rect 3715 15989 3833 16028
tri 4871 16026 4873 16028 ne
rect 4873 16026 5011 16028
tri 5011 16026 5013 16028 nw
tri 4873 16021 4878 16026 ne
rect 3076 15913 3128 15952
rect 2816 15842 2822 15876
rect 2856 15842 2862 15876
rect 2816 15803 2862 15842
rect 2816 15769 2822 15803
rect 2856 15769 2862 15803
rect 2816 15730 2862 15769
rect 2816 15696 2822 15730
rect 2856 15696 2862 15730
rect 2816 15657 2862 15696
rect 2816 15623 2822 15657
rect 2856 15623 2862 15657
rect 2816 15584 2862 15623
rect 2816 15550 2822 15584
rect 2856 15550 2862 15584
rect 2816 15511 2862 15550
rect 2816 15477 2822 15511
rect 2856 15477 2862 15511
rect 2816 15438 2862 15477
rect 2816 15404 2822 15438
rect 2856 15404 2862 15438
rect 2816 15365 2862 15404
rect 2816 15331 2822 15365
rect 2856 15331 2862 15365
rect 2816 15292 2862 15331
rect 2816 15258 2822 15292
rect 2856 15258 2862 15292
rect 2816 15219 2862 15258
rect 2816 15185 2822 15219
rect 2856 15185 2862 15219
rect 2816 15146 2862 15185
rect 2816 15112 2822 15146
rect 2856 15112 2862 15146
rect 2816 15073 2862 15112
rect 2816 15039 2822 15073
rect 2856 15039 2862 15073
rect 2816 15000 2862 15039
rect 2816 14966 2822 15000
rect 2856 14966 2862 15000
rect 2816 14927 2862 14966
rect 2816 14893 2822 14927
rect 2856 14893 2862 14927
rect 2816 14854 2862 14893
rect 2816 14820 2822 14854
rect 2856 14820 2862 14854
rect 2816 14781 2862 14820
rect 2816 14747 2822 14781
rect 2856 14747 2862 14781
rect 2816 14708 2862 14747
rect 2816 14674 2822 14708
rect 2856 14674 2862 14708
rect 2816 14635 2862 14674
rect 2816 14601 2822 14635
rect 2856 14601 2862 14635
rect 2816 14562 2862 14601
rect 3076 15879 3082 15913
rect 3116 15879 3128 15913
rect 3076 15872 3128 15879
rect 3076 15808 3082 15820
rect 3116 15808 3128 15820
rect 3076 15733 3082 15756
rect 3116 15733 3128 15756
rect 3076 15694 3128 15733
rect 3076 15660 3082 15694
rect 3116 15660 3128 15694
rect 3076 15621 3128 15660
rect 3076 15587 3082 15621
rect 3116 15587 3128 15621
rect 3076 15548 3128 15587
rect 3076 15514 3082 15548
rect 3116 15514 3128 15548
rect 3076 15475 3128 15514
rect 3076 15441 3082 15475
rect 3116 15441 3128 15475
rect 3076 15402 3128 15441
rect 3076 15368 3082 15402
rect 3116 15368 3128 15402
rect 3076 15329 3128 15368
rect 3076 15295 3082 15329
rect 3116 15295 3128 15329
rect 3076 15256 3128 15295
rect 3076 15222 3082 15256
rect 3116 15222 3128 15256
rect 3076 15183 3128 15222
rect 3076 15149 3082 15183
rect 3116 15149 3128 15183
rect 3076 15110 3128 15149
rect 3076 15076 3082 15110
rect 3116 15076 3128 15110
rect 3076 15037 3128 15076
rect 3076 15003 3082 15037
rect 3116 15003 3128 15037
rect 3076 14964 3128 15003
rect 3076 14930 3082 14964
rect 3116 14930 3128 14964
rect 3076 14891 3128 14930
rect 3076 14857 3082 14891
rect 3116 14857 3128 14891
rect 3076 14819 3128 14857
rect 3076 14785 3082 14819
rect 3116 14785 3128 14819
rect 3076 14747 3128 14785
rect 3076 14713 3082 14747
rect 3116 14713 3128 14747
rect 3076 14675 3128 14713
rect 3076 14641 3082 14675
rect 3116 14641 3128 14675
rect 3715 15955 3721 15989
rect 3755 15955 3793 15989
rect 3827 15955 3833 15989
rect 3715 15916 3833 15955
rect 3715 15882 3721 15916
rect 3755 15882 3793 15916
rect 3827 15882 3833 15916
rect 3715 15843 3833 15882
rect 3715 15809 3721 15843
rect 3755 15809 3793 15843
rect 3827 15809 3833 15843
rect 3715 15770 3833 15809
rect 3715 15736 3721 15770
rect 3755 15736 3793 15770
rect 3827 15736 3833 15770
rect 3715 15697 3833 15736
rect 3715 15663 3721 15697
rect 3755 15663 3793 15697
rect 3827 15663 3833 15697
rect 3715 15624 3833 15663
rect 3715 15590 3721 15624
rect 3755 15590 3793 15624
rect 3827 15590 3833 15624
rect 3715 15551 3833 15590
rect 3715 15517 3721 15551
rect 3755 15517 3793 15551
rect 3827 15517 3833 15551
rect 3715 15478 3833 15517
rect 3715 15444 3721 15478
rect 3755 15444 3793 15478
rect 3827 15444 3833 15478
rect 3715 15405 3833 15444
rect 3715 15371 3721 15405
rect 3755 15371 3793 15405
rect 3827 15371 3833 15405
rect 3715 15332 3833 15371
rect 3715 15298 3721 15332
rect 3755 15298 3793 15332
rect 3827 15298 3833 15332
rect 3715 15259 3833 15298
rect 3715 15225 3721 15259
rect 3755 15225 3793 15259
rect 3827 15225 3833 15259
rect 3715 15186 3833 15225
rect 3715 15152 3721 15186
rect 3755 15152 3793 15186
rect 3827 15152 3833 15186
rect 3715 15113 3833 15152
rect 3715 15079 3721 15113
rect 3755 15079 3793 15113
rect 3827 15079 3833 15113
rect 3715 15040 3833 15079
rect 3715 15006 3721 15040
rect 3755 15006 3793 15040
rect 3827 15006 3833 15040
rect 3715 14967 3833 15006
rect 3715 14933 3721 14967
rect 3755 14933 3793 14967
rect 3827 14933 3833 14967
rect 3715 14894 3833 14933
rect 3715 14860 3721 14894
rect 3755 14860 3793 14894
rect 3827 14860 3833 14894
rect 3715 14821 3833 14860
rect 3715 14787 3721 14821
rect 3755 14787 3793 14821
rect 3827 14787 3833 14821
rect 3715 14748 3833 14787
rect 3715 14714 3721 14748
rect 3755 14714 3793 14748
rect 3827 14714 3833 14748
rect 3715 14675 3833 14714
tri 3128 14641 3130 14643 sw
tri 3713 14641 3715 14643 se
rect 3715 14641 3721 14675
rect 3755 14641 3793 14675
rect 3827 14641 3833 14675
rect 4130 14667 4230 15959
tri 4854 15381 4878 15405 se
rect 4878 15381 5006 16026
tri 5006 16021 5011 16026 nw
tri 5006 15381 5030 15405 sw
rect 5840 15397 5940 16689
rect 6211 16685 6476 16711
rect 6510 16685 6516 16719
rect 6211 16672 6516 16685
rect 6211 16638 6237 16672
rect 6271 16638 6309 16672
rect 6343 16646 6516 16672
rect 6343 16638 6476 16646
rect 6211 16612 6476 16638
rect 6510 16612 6516 16646
rect 6211 16599 6516 16612
rect 6211 16565 6237 16599
rect 6271 16565 6309 16599
rect 6343 16573 6516 16599
rect 6343 16565 6476 16573
rect 6211 16539 6476 16565
rect 6510 16539 6516 16573
rect 6211 16525 6516 16539
rect 6211 16491 6237 16525
rect 6271 16491 6309 16525
rect 6343 16500 6516 16525
rect 6343 16491 6476 16500
rect 6211 16466 6476 16491
rect 6510 16466 6516 16500
rect 6211 16451 6516 16466
rect 6211 16417 6237 16451
rect 6271 16417 6309 16451
rect 6343 16427 6516 16451
rect 6343 16417 6476 16427
rect 6211 16393 6476 16417
rect 6510 16393 6516 16427
rect 6211 16377 6516 16393
rect 6211 16343 6237 16377
rect 6271 16343 6309 16377
rect 6343 16354 6516 16377
rect 6343 16343 6476 16354
rect 6211 16320 6476 16343
rect 6510 16320 6516 16354
rect 6211 16303 6516 16320
rect 6211 16269 6237 16303
rect 6271 16269 6309 16303
rect 6343 16281 6516 16303
rect 6343 16269 6476 16281
rect 6211 16247 6476 16269
rect 6510 16247 6516 16281
rect 6211 16229 6516 16247
rect 6211 16195 6237 16229
rect 6271 16195 6309 16229
rect 6343 16208 6516 16229
rect 6343 16195 6476 16208
rect 6211 16174 6476 16195
rect 6510 16174 6516 16208
rect 6211 16155 6516 16174
rect 6211 16121 6237 16155
rect 6271 16121 6309 16155
rect 6343 16135 6516 16155
rect 6343 16121 6476 16135
rect 6211 16101 6476 16121
rect 6510 16101 6516 16135
rect 6211 16081 6516 16101
rect 6211 16047 6237 16081
rect 6271 16047 6309 16081
rect 6343 16062 6516 16081
rect 6343 16047 6476 16062
rect 6211 16028 6476 16047
rect 6510 16028 6516 16062
rect 6211 16007 6516 16028
rect 6211 15973 6237 16007
rect 6271 15973 6309 16007
rect 6343 15989 6516 16007
rect 6343 15973 6476 15989
rect 6211 15955 6476 15973
rect 6510 15955 6516 15989
rect 6211 15933 6516 15955
rect 6211 15899 6237 15933
rect 6271 15899 6309 15933
rect 6343 15916 6516 15933
rect 6343 15899 6476 15916
rect 6211 15882 6476 15899
rect 6510 15882 6516 15916
rect 6211 15872 6516 15882
rect 6211 15859 6464 15872
rect 6211 15825 6237 15859
rect 6271 15825 6309 15859
rect 6343 15825 6464 15859
rect 6211 15820 6464 15825
rect 6211 15809 6476 15820
rect 6510 15809 6516 15820
rect 6211 15808 6516 15809
rect 6211 15785 6464 15808
rect 6211 15751 6237 15785
rect 6271 15751 6309 15785
rect 6343 15756 6464 15785
rect 6343 15751 6476 15756
rect 6211 15736 6476 15751
rect 6510 15736 6516 15756
rect 6211 15711 6516 15736
rect 6211 15677 6237 15711
rect 6271 15677 6309 15711
rect 6343 15697 6516 15711
rect 6343 15677 6476 15697
rect 6211 15663 6476 15677
rect 6510 15663 6516 15697
rect 6211 15637 6516 15663
rect 6211 15603 6237 15637
rect 6271 15603 6309 15637
rect 6343 15624 6516 15637
rect 6343 15603 6476 15624
rect 6211 15590 6476 15603
rect 6510 15590 6516 15624
rect 6211 15563 6516 15590
rect 6211 15529 6237 15563
rect 6271 15529 6309 15563
rect 6343 15551 6516 15563
rect 6343 15529 6476 15551
rect 6211 15517 6476 15529
rect 6510 15517 6516 15551
rect 6211 15489 6516 15517
rect 6211 15455 6237 15489
rect 6271 15455 6309 15489
rect 6343 15478 6516 15489
rect 6343 15455 6476 15478
rect 6211 15444 6476 15455
rect 6510 15444 6516 15478
rect 6211 15415 6516 15444
rect 6211 15381 6237 15415
rect 6271 15381 6309 15415
rect 6343 15405 6516 15415
rect 6343 15381 6476 15405
tri 4844 15371 4854 15381 se
rect 4854 15371 5030 15381
tri 5030 15371 5040 15381 sw
rect 6211 15371 6476 15381
rect 6510 15371 6516 15405
rect 4270 15365 5788 15371
rect 4270 15331 4282 15365
rect 4316 15331 4355 15365
rect 4389 15331 4428 15365
rect 4462 15331 4501 15365
rect 4535 15331 4574 15365
rect 4608 15331 4647 15365
rect 4681 15331 4720 15365
rect 4754 15331 4793 15365
rect 4827 15331 4866 15365
rect 4900 15331 4939 15365
rect 4973 15331 5012 15365
rect 5046 15331 5085 15365
rect 5119 15331 5158 15365
rect 5192 15331 5231 15365
rect 5265 15331 5304 15365
rect 5338 15331 5377 15365
rect 5411 15331 5450 15365
rect 5484 15331 5523 15365
rect 5557 15331 5596 15365
rect 5630 15331 5669 15365
rect 5703 15331 5742 15365
rect 5776 15331 5788 15365
rect 4270 15325 5788 15331
rect 6211 15341 6516 15371
rect 6211 15307 6237 15341
rect 6271 15307 6309 15341
rect 6343 15332 6516 15341
rect 6343 15307 6476 15332
rect 6211 15298 6476 15307
rect 6510 15298 6516 15332
rect 6211 15267 6516 15298
rect 6211 15233 6237 15267
rect 6271 15233 6309 15267
rect 6343 15259 6516 15267
rect 6343 15233 6476 15259
rect 6211 15225 6476 15233
rect 6510 15225 6516 15259
rect 6211 15193 6516 15225
rect 6211 15159 6237 15193
rect 6271 15159 6309 15193
rect 6343 15186 6516 15193
rect 6343 15159 6476 15186
rect 6211 15152 6476 15159
rect 6510 15152 6516 15186
rect 6211 15119 6516 15152
rect 6211 15085 6237 15119
rect 6271 15085 6309 15119
rect 6343 15113 6516 15119
rect 6343 15085 6476 15113
rect 6211 15079 6476 15085
rect 6510 15079 6516 15113
rect 6211 15045 6516 15079
rect 6211 15011 6237 15045
rect 6271 15011 6309 15045
rect 6343 15040 6516 15045
rect 6343 15011 6476 15040
rect 6211 15006 6476 15011
rect 6510 15006 6516 15040
rect 6211 14971 6516 15006
rect 6211 14937 6237 14971
rect 6271 14937 6309 14971
rect 6343 14967 6516 14971
rect 6343 14937 6476 14967
rect 6211 14933 6476 14937
rect 6510 14933 6516 14967
rect 6211 14897 6516 14933
rect 5837 14861 5889 14867
rect 5837 14793 5889 14809
rect 5837 14725 5889 14741
rect 5837 14667 5889 14673
rect 6211 14863 6237 14897
rect 6271 14863 6309 14897
rect 6343 14894 6516 14897
rect 6343 14863 6476 14894
rect 6211 14861 6476 14863
rect 6510 14861 6516 14894
rect 6263 14823 6295 14861
rect 6271 14809 6295 14823
rect 6347 14809 6379 14861
rect 6431 14809 6463 14861
rect 6515 14809 6516 14861
rect 6211 14793 6237 14809
rect 6271 14793 6309 14809
rect 6343 14793 6476 14809
rect 6510 14793 6516 14809
rect 6271 14789 6295 14793
rect 6263 14749 6295 14789
rect 6271 14741 6295 14749
rect 6347 14741 6379 14793
rect 6431 14741 6463 14793
rect 6515 14741 6516 14793
rect 6211 14725 6237 14741
rect 6271 14725 6309 14741
rect 6343 14725 6476 14741
rect 6510 14725 6516 14741
rect 6271 14715 6295 14725
rect 6263 14675 6295 14715
rect 6347 14673 6379 14725
rect 6431 14673 6463 14725
rect 6515 14673 6516 14725
rect 3076 14609 3130 14641
tri 3130 14609 3162 14641 sw
tri 3681 14609 3713 14641 se
rect 3713 14609 3833 14641
tri 3833 14609 3867 14643 sw
tri 6177 14609 6211 14643 se
rect 6211 14609 6237 14673
rect 3076 14603 6237 14609
rect 6343 14641 6476 14673
rect 6510 14641 6516 14673
rect 6343 14603 6516 14641
rect 3076 14569 3154 14603
rect 3188 14569 3227 14603
rect 3261 14569 3300 14603
rect 3334 14569 3373 14603
rect 3407 14569 3446 14603
rect 3480 14569 3519 14603
rect 3553 14569 3592 14603
rect 3626 14569 3665 14603
rect 3699 14569 3738 14603
rect 3772 14569 3811 14603
rect 3845 14569 3884 14603
rect 3918 14569 3956 14603
rect 3990 14569 4028 14603
rect 4062 14569 4100 14603
rect 4134 14569 4172 14603
rect 4206 14569 4244 14603
rect 4278 14569 4316 14603
rect 4350 14569 4388 14603
rect 4422 14569 4460 14603
rect 4494 14569 4532 14603
rect 4566 14569 4604 14603
rect 4638 14569 4676 14603
rect 4710 14569 4748 14603
rect 4782 14569 4820 14603
rect 4854 14569 4892 14603
rect 4926 14569 4964 14603
rect 4998 14569 5036 14603
rect 5070 14569 5108 14603
rect 5142 14569 5180 14603
rect 5214 14569 5252 14603
rect 5286 14569 5324 14603
rect 5358 14569 5396 14603
rect 5430 14569 5468 14603
rect 5502 14569 5540 14603
rect 5574 14569 5612 14603
rect 5646 14569 5684 14603
rect 5718 14569 5756 14603
rect 5790 14569 5828 14603
rect 5862 14569 5900 14603
rect 5934 14569 5972 14603
rect 6006 14569 6044 14603
rect 6078 14569 6116 14603
rect 6150 14569 6188 14603
rect 6222 14569 6237 14603
rect 6366 14569 6404 14603
rect 6438 14569 6516 14603
rect 3076 14563 6516 14569
rect 6744 17997 6790 18036
rect 6744 17963 6750 17997
rect 6784 17963 6790 17997
rect 6744 17924 6790 17963
rect 6744 17890 6750 17924
rect 6784 17890 6790 17924
rect 6744 17851 6790 17890
rect 6744 17817 6750 17851
rect 6784 17817 6790 17851
rect 6744 17778 6790 17817
rect 6744 17744 6750 17778
rect 6784 17744 6790 17778
rect 6744 17705 6790 17744
rect 6744 17671 6750 17705
rect 6784 17671 6790 17705
rect 6744 17632 6790 17671
rect 6744 17598 6750 17632
rect 6784 17598 6790 17632
rect 6744 17559 6790 17598
rect 6744 17525 6750 17559
rect 6784 17525 6790 17559
rect 6744 17486 6790 17525
rect 6744 17452 6750 17486
rect 6784 17452 6790 17486
rect 6744 17413 6790 17452
rect 6744 17379 6750 17413
rect 6784 17379 6790 17413
rect 8793 17461 8921 19971
rect 8793 17409 8799 17461
rect 8851 17409 8863 17461
rect 8915 17409 8921 17461
rect 8793 17403 8921 17409
rect 6744 17340 6790 17379
rect 6744 17306 6750 17340
rect 6784 17306 6790 17340
rect 6744 17267 6790 17306
rect 6744 17233 6750 17267
rect 6784 17233 6790 17267
rect 6744 17194 6790 17233
rect 6744 17160 6750 17194
rect 6784 17160 6790 17194
rect 6744 17121 6790 17160
rect 6744 17087 6750 17121
rect 6784 17087 6790 17121
rect 6744 17048 6790 17087
rect 6744 17014 6750 17048
rect 6784 17014 6790 17048
rect 6744 16975 6790 17014
rect 6744 16941 6750 16975
rect 6784 16941 6790 16975
rect 6744 16902 6790 16941
rect 6744 16868 6750 16902
rect 6784 16868 6790 16902
rect 6744 16829 6790 16868
rect 6744 16795 6750 16829
rect 6784 16795 6790 16829
rect 6744 16756 6790 16795
rect 6744 16722 6750 16756
rect 6784 16722 6790 16756
rect 6744 16683 6790 16722
rect 6744 16649 6750 16683
rect 6784 16649 6790 16683
rect 6744 16610 6790 16649
rect 6744 16576 6750 16610
rect 6784 16576 6790 16610
rect 6744 16537 6790 16576
rect 6744 16503 6750 16537
rect 6784 16503 6790 16537
rect 6744 16464 6790 16503
rect 6744 16430 6750 16464
rect 6784 16430 6790 16464
rect 6744 16391 6790 16430
rect 6744 16357 6750 16391
rect 6784 16357 6790 16391
rect 6744 16318 6790 16357
rect 6744 16284 6750 16318
rect 6784 16284 6790 16318
rect 6744 16245 6790 16284
rect 6744 16211 6750 16245
rect 6784 16211 6790 16245
rect 6744 16172 6790 16211
rect 6744 16138 6750 16172
rect 6784 16138 6790 16172
rect 6744 16099 6790 16138
rect 6744 16065 6750 16099
rect 6784 16065 6790 16099
rect 6744 16026 6790 16065
rect 6744 15992 6750 16026
rect 6784 15992 6790 16026
rect 6744 15953 6790 15992
rect 6744 15919 6750 15953
rect 6784 15919 6790 15953
rect 6744 15880 6790 15919
rect 6744 15846 6750 15880
rect 6784 15846 6790 15880
rect 6744 15807 6790 15846
rect 6744 15773 6750 15807
rect 6784 15773 6790 15807
rect 6744 15734 6790 15773
rect 6744 15700 6750 15734
rect 6784 15700 6790 15734
rect 6744 15661 6790 15700
rect 6744 15627 6750 15661
rect 6784 15627 6790 15661
rect 6744 15588 6790 15627
rect 6744 15554 6750 15588
rect 6784 15554 6790 15588
rect 6744 15515 6790 15554
rect 6744 15481 6750 15515
rect 6784 15481 6790 15515
rect 6744 15442 6790 15481
rect 6744 15408 6750 15442
rect 6784 15408 6790 15442
rect 6744 15369 6790 15408
rect 6744 15335 6750 15369
rect 6784 15335 6790 15369
rect 6744 15296 6790 15335
rect 6744 15262 6750 15296
rect 6784 15262 6790 15296
rect 6744 15223 6790 15262
rect 6744 15189 6750 15223
rect 6784 15189 6790 15223
rect 6744 15150 6790 15189
rect 6744 15116 6750 15150
rect 6784 15116 6790 15150
rect 6744 15077 6790 15116
rect 6744 15043 6750 15077
rect 6784 15043 6790 15077
rect 6744 15004 6790 15043
rect 6744 14970 6750 15004
rect 6784 14970 6790 15004
rect 6744 14931 6790 14970
rect 6744 14897 6750 14931
rect 6784 14897 6790 14931
rect 6744 14858 6790 14897
rect 6744 14824 6750 14858
rect 6784 14824 6790 14858
rect 6744 14785 6790 14824
rect 6744 14751 6750 14785
rect 6784 14751 6790 14785
rect 6744 14711 6790 14751
rect 6744 14677 6750 14711
rect 6784 14677 6790 14711
rect 6744 14637 6790 14677
rect 6744 14603 6750 14637
rect 6784 14603 6790 14637
rect 6744 14563 6790 14603
rect 2816 14528 2822 14562
rect 2856 14528 2862 14562
rect 2816 14489 2862 14528
rect 2816 14455 2822 14489
rect 2856 14455 2862 14489
rect 2816 14416 2862 14455
rect 2816 14382 2822 14416
rect 2856 14382 2862 14416
rect 6744 14529 6750 14563
rect 6784 14529 6790 14563
rect 6744 14489 6790 14529
rect 6744 14455 6750 14489
rect 6784 14455 6790 14489
rect 6744 14415 6790 14455
rect 2816 14381 2862 14382
tri 2862 14381 2867 14386 sw
tri 6739 14381 6744 14386 se
rect 6744 14381 6750 14415
rect 6784 14381 6790 14415
rect 2816 14352 2867 14381
tri 2867 14352 2896 14381 sw
tri 6710 14352 6739 14381 se
rect 6739 14352 6790 14381
rect 2816 14343 6790 14352
rect 2816 14309 2894 14343
rect 2928 14309 2967 14343
rect 3001 14309 3040 14343
rect 3074 14309 3113 14343
rect 3147 14309 3186 14343
rect 3220 14309 3259 14343
rect 3293 14309 3332 14343
rect 3366 14309 3405 14343
rect 3439 14309 3478 14343
rect 3512 14309 3551 14343
rect 3585 14309 3624 14343
rect 3658 14309 3697 14343
rect 3731 14309 3770 14343
rect 3804 14309 3843 14343
rect 3877 14309 3916 14343
rect 3950 14309 3989 14343
rect 4023 14309 4062 14343
rect 4096 14309 4135 14343
rect 4169 14309 4208 14343
rect 4242 14309 4281 14343
rect 4315 14309 4354 14343
rect 4388 14309 4427 14343
rect 4461 14309 4500 14343
rect 4534 14309 4573 14343
rect 4607 14309 4646 14343
rect 4680 14309 4719 14343
rect 4753 14309 4792 14343
rect 4826 14309 4865 14343
rect 4899 14309 4938 14343
rect 4972 14309 5011 14343
rect 5045 14309 5084 14343
rect 5118 14309 5157 14343
rect 5191 14309 5230 14343
rect 5264 14309 5303 14343
rect 5337 14309 5376 14343
rect 5410 14309 5449 14343
rect 5483 14309 5522 14343
rect 5556 14309 5595 14343
rect 5629 14309 5668 14343
rect 5702 14309 5741 14343
rect 5775 14309 5814 14343
rect 5848 14309 5886 14343
rect 5920 14309 5958 14343
rect 5992 14309 6030 14343
rect 6064 14309 6102 14343
rect 6136 14309 6174 14343
rect 6208 14309 6246 14343
rect 6280 14309 6318 14343
rect 6352 14309 6390 14343
rect 6424 14309 6462 14343
rect 6496 14309 6534 14343
rect 6568 14309 6606 14343
rect 6640 14309 6678 14343
rect 6712 14309 6790 14343
rect 2816 14300 6790 14309
<< via1 >>
rect 1211 35591 1263 35643
rect 1211 35527 1263 35579
rect 2633 29435 2685 29487
rect 2730 29435 2782 29487
rect 2633 29359 2685 29411
rect 2730 29359 2782 29411
rect 1187 26150 1239 26202
rect 1187 26086 1239 26138
rect 932 25755 984 25807
rect 932 25691 984 25743
rect 908 16734 960 16786
rect 908 16668 960 16720
rect 908 16602 960 16654
rect 908 16536 960 16588
rect 1187 25549 1239 25601
rect 1187 25485 1239 25537
rect 2294 28957 2346 29009
rect 2391 28957 2443 29009
rect 2294 22478 2346 22530
rect 2391 22478 2443 22530
rect 2294 22402 2346 22454
rect 2391 22402 2443 22454
rect 2294 19219 2346 19271
rect 2391 19219 2443 19271
rect 2294 19155 2346 19207
rect 2391 19155 2443 19207
rect 4666 39143 4718 39195
rect 4732 39143 4784 39195
rect 4798 39143 4850 39195
rect 4864 39143 4916 39195
rect 4930 39143 4982 39195
rect 4996 39143 5048 39195
rect 5062 39143 5114 39195
rect 5128 39143 5180 39195
rect 5194 39143 5246 39195
rect 5260 39143 5312 39195
rect 5326 39182 5378 39195
rect 5326 39148 5330 39182
rect 5330 39148 5364 39182
rect 5364 39148 5378 39182
rect 5326 39143 5378 39148
rect 5392 39143 5444 39195
rect 4666 39079 4718 39131
rect 4732 39079 4784 39131
rect 4798 39079 4850 39131
rect 4864 39079 4916 39131
rect 4930 39079 4982 39131
rect 4996 39079 5048 39131
rect 5062 39079 5114 39131
rect 5128 39079 5180 39131
rect 5194 39079 5246 39131
rect 5260 39079 5312 39131
rect 5326 39110 5378 39131
rect 5326 39079 5330 39110
rect 5330 39079 5364 39110
rect 5364 39079 5378 39110
rect 5392 39079 5444 39131
rect 4666 39015 4718 39067
rect 4732 39015 4784 39067
rect 4798 39015 4850 39067
rect 4864 39015 4916 39067
rect 4930 39015 4982 39067
rect 4996 39015 5048 39067
rect 5062 39015 5114 39067
rect 5128 39015 5180 39067
rect 5194 39015 5246 39067
rect 5260 39015 5312 39067
rect 5326 39038 5378 39067
rect 5326 39015 5330 39038
rect 5330 39015 5364 39038
rect 5364 39015 5378 39038
rect 5392 39015 5444 39067
rect 4666 38951 4718 39003
rect 4732 38951 4784 39003
rect 4798 38951 4850 39003
rect 4864 38951 4916 39003
rect 4930 38951 4982 39003
rect 4996 38951 5048 39003
rect 5062 38951 5114 39003
rect 5128 38951 5180 39003
rect 5194 38951 5246 39003
rect 5260 38951 5312 39003
rect 5326 38966 5378 39003
rect 5326 38951 5330 38966
rect 5330 38951 5364 38966
rect 5364 38951 5378 38966
rect 5392 38951 5444 39003
rect 4666 38887 4718 38939
rect 4732 38887 4784 38939
rect 4798 38887 4850 38939
rect 4864 38887 4916 38939
rect 4930 38887 4982 38939
rect 4996 38887 5048 38939
rect 5062 38887 5114 38939
rect 5128 38887 5180 38939
rect 5194 38887 5246 38939
rect 5260 38887 5312 38939
rect 5326 38932 5330 38939
rect 5330 38932 5364 38939
rect 5364 38932 5378 38939
rect 5326 38894 5378 38932
rect 5326 38887 5330 38894
rect 5330 38887 5364 38894
rect 5364 38887 5378 38894
rect 5392 38887 5444 38939
rect 4666 38823 4718 38875
rect 4732 38823 4784 38875
rect 4798 38823 4850 38875
rect 4864 38823 4916 38875
rect 4930 38823 4982 38875
rect 4996 38823 5048 38875
rect 5062 38823 5114 38875
rect 5128 38823 5180 38875
rect 5194 38823 5246 38875
rect 5260 38823 5312 38875
rect 5326 38860 5330 38875
rect 5330 38860 5364 38875
rect 5364 38860 5378 38875
rect 5326 38823 5378 38860
rect 5392 38823 5444 38875
rect 4666 38759 4718 38811
rect 4732 38759 4784 38811
rect 4798 38759 4850 38811
rect 4864 38759 4916 38811
rect 4930 38759 4982 38811
rect 4996 38759 5048 38811
rect 5062 38759 5114 38811
rect 5128 38759 5180 38811
rect 5194 38759 5246 38811
rect 5260 38759 5312 38811
rect 5326 38788 5330 38811
rect 5330 38788 5364 38811
rect 5364 38788 5378 38811
rect 5326 38759 5378 38788
rect 5392 38759 5444 38811
rect 4666 38695 4718 38747
rect 4732 38695 4784 38747
rect 4798 38695 4850 38747
rect 4864 38695 4916 38747
rect 4930 38695 4982 38747
rect 4996 38695 5048 38747
rect 5062 38695 5114 38747
rect 5128 38695 5180 38747
rect 5194 38695 5246 38747
rect 5260 38695 5312 38747
rect 5326 38716 5330 38747
rect 5330 38716 5364 38747
rect 5364 38716 5378 38747
rect 5326 38695 5378 38716
rect 5392 38695 5444 38747
rect 4666 38631 4718 38683
rect 4732 38631 4784 38683
rect 4798 38631 4850 38683
rect 4864 38631 4916 38683
rect 4930 38631 4982 38683
rect 4996 38631 5048 38683
rect 5062 38631 5114 38683
rect 5128 38631 5180 38683
rect 5194 38631 5246 38683
rect 5260 38631 5312 38683
rect 5326 38678 5378 38683
rect 5326 38644 5330 38678
rect 5330 38644 5364 38678
rect 5364 38644 5378 38678
rect 5326 38631 5378 38644
rect 5392 38631 5444 38683
rect 4666 38567 4718 38619
rect 4732 38567 4784 38619
rect 4798 38567 4850 38619
rect 4864 38567 4916 38619
rect 4930 38567 4982 38619
rect 4996 38567 5048 38619
rect 5062 38567 5114 38619
rect 5128 38567 5180 38619
rect 5194 38567 5246 38619
rect 5260 38567 5312 38619
rect 5326 38606 5378 38619
rect 5326 38572 5330 38606
rect 5330 38572 5364 38606
rect 5364 38572 5378 38606
rect 5326 38567 5378 38572
rect 5392 38567 5444 38619
rect 4666 38503 4718 38555
rect 4732 38503 4784 38555
rect 4798 38503 4850 38555
rect 4864 38503 4916 38555
rect 4930 38503 4982 38555
rect 4996 38503 5048 38555
rect 5062 38503 5114 38555
rect 5128 38503 5180 38555
rect 5194 38503 5246 38555
rect 5260 38503 5312 38555
rect 5326 38534 5378 38555
rect 5326 38503 5330 38534
rect 5330 38503 5364 38534
rect 5364 38503 5378 38534
rect 5392 38503 5444 38555
rect 4666 38439 4718 38491
rect 4732 38439 4784 38491
rect 4798 38439 4850 38491
rect 4864 38439 4916 38491
rect 4930 38439 4982 38491
rect 4996 38439 5048 38491
rect 5062 38439 5114 38491
rect 5128 38439 5180 38491
rect 5194 38439 5246 38491
rect 5260 38439 5312 38491
rect 5326 38462 5378 38491
rect 5326 38439 5330 38462
rect 5330 38439 5364 38462
rect 5364 38439 5378 38462
rect 5392 38439 5444 38491
rect 4666 38375 4718 38427
rect 4732 38375 4784 38427
rect 4798 38375 4850 38427
rect 4864 38375 4916 38427
rect 4930 38375 4982 38427
rect 4996 38375 5048 38427
rect 5062 38375 5114 38427
rect 5128 38375 5180 38427
rect 5194 38375 5246 38427
rect 5260 38375 5312 38427
rect 5326 38390 5378 38427
rect 5326 38375 5330 38390
rect 5330 38375 5364 38390
rect 5364 38375 5378 38390
rect 5392 38375 5444 38427
rect 4666 38311 4718 38363
rect 4732 38311 4784 38363
rect 4798 38311 4850 38363
rect 4864 38311 4916 38363
rect 4930 38311 4982 38363
rect 4996 38311 5048 38363
rect 5062 38311 5114 38363
rect 5128 38311 5180 38363
rect 5194 38311 5246 38363
rect 5260 38311 5312 38363
rect 5326 38356 5330 38363
rect 5330 38356 5364 38363
rect 5364 38356 5378 38363
rect 5326 38318 5378 38356
rect 5326 38311 5330 38318
rect 5330 38311 5364 38318
rect 5364 38311 5378 38318
rect 5392 38311 5444 38363
rect 4666 38247 4718 38299
rect 4732 38247 4784 38299
rect 4798 38247 4850 38299
rect 4864 38247 4916 38299
rect 4930 38247 4982 38299
rect 4996 38247 5048 38299
rect 5062 38247 5114 38299
rect 5128 38247 5180 38299
rect 5194 38247 5246 38299
rect 5260 38247 5312 38299
rect 5326 38284 5330 38299
rect 5330 38284 5364 38299
rect 5364 38284 5378 38299
rect 5326 38247 5378 38284
rect 5392 38247 5444 38299
rect 4666 38183 4718 38235
rect 4732 38183 4784 38235
rect 4798 38183 4850 38235
rect 4864 38183 4916 38235
rect 4930 38183 4982 38235
rect 4996 38183 5048 38235
rect 5062 38183 5114 38235
rect 5128 38183 5180 38235
rect 5194 38183 5246 38235
rect 5260 38183 5312 38235
rect 5326 38212 5330 38235
rect 5330 38212 5364 38235
rect 5364 38212 5378 38235
rect 5326 38183 5378 38212
rect 5392 38183 5444 38235
rect 4666 38119 4718 38171
rect 4732 38119 4784 38171
rect 4798 38119 4850 38171
rect 4864 38119 4916 38171
rect 4930 38119 4982 38171
rect 4996 38119 5048 38171
rect 5062 38119 5114 38171
rect 5128 38119 5180 38171
rect 5194 38119 5246 38171
rect 5260 38119 5312 38171
rect 5326 38140 5330 38171
rect 5330 38140 5364 38171
rect 5364 38140 5378 38171
rect 5326 38119 5378 38140
rect 5392 38119 5444 38171
rect 4666 38055 4718 38107
rect 4732 38055 4784 38107
rect 4798 38055 4850 38107
rect 4864 38055 4916 38107
rect 4930 38055 4982 38107
rect 4996 38055 5048 38107
rect 5062 38055 5114 38107
rect 5128 38055 5180 38107
rect 5194 38055 5246 38107
rect 5260 38055 5312 38107
rect 5326 38102 5378 38107
rect 5326 38068 5330 38102
rect 5330 38068 5364 38102
rect 5364 38068 5378 38102
rect 5326 38055 5378 38068
rect 5392 38055 5444 38107
rect 4666 37991 4718 38043
rect 4732 37991 4784 38043
rect 4798 37991 4850 38043
rect 4864 37991 4916 38043
rect 4930 37991 4982 38043
rect 4996 37991 5048 38043
rect 5062 37991 5114 38043
rect 5128 37991 5180 38043
rect 5194 37991 5246 38043
rect 5260 37991 5312 38043
rect 5326 38030 5378 38043
rect 5326 37996 5330 38030
rect 5330 37996 5364 38030
rect 5364 37996 5378 38030
rect 5326 37991 5378 37996
rect 5392 37991 5444 38043
rect 4666 37927 4718 37979
rect 4732 37927 4784 37979
rect 4798 37927 4850 37979
rect 4864 37927 4916 37979
rect 4930 37927 4982 37979
rect 4996 37927 5048 37979
rect 5062 37927 5114 37979
rect 5128 37927 5180 37979
rect 5194 37927 5246 37979
rect 5260 37927 5312 37979
rect 5326 37958 5378 37979
rect 5326 37927 5330 37958
rect 5330 37927 5364 37958
rect 5364 37927 5378 37958
rect 5392 37927 5444 37979
rect 4666 37863 4718 37915
rect 4732 37863 4784 37915
rect 4798 37863 4850 37915
rect 4864 37863 4916 37915
rect 4930 37863 4982 37915
rect 4996 37863 5048 37915
rect 5062 37863 5114 37915
rect 5128 37863 5180 37915
rect 5194 37863 5246 37915
rect 5260 37863 5312 37915
rect 5326 37886 5378 37915
rect 5326 37863 5330 37886
rect 5330 37863 5364 37886
rect 5364 37863 5378 37886
rect 5392 37863 5444 37915
rect 4666 37799 4718 37851
rect 4732 37799 4784 37851
rect 4798 37799 4850 37851
rect 4864 37799 4916 37851
rect 4930 37799 4982 37851
rect 4996 37799 5048 37851
rect 5062 37799 5114 37851
rect 5128 37799 5180 37851
rect 5194 37799 5246 37851
rect 5260 37799 5312 37851
rect 5326 37814 5378 37851
rect 5326 37799 5330 37814
rect 5330 37799 5364 37814
rect 5364 37799 5378 37814
rect 5392 37799 5444 37851
rect 4666 37735 4718 37787
rect 4732 37735 4784 37787
rect 4798 37735 4850 37787
rect 4864 37735 4916 37787
rect 4930 37735 4982 37787
rect 4996 37735 5048 37787
rect 5062 37735 5114 37787
rect 5128 37735 5180 37787
rect 5194 37735 5246 37787
rect 5260 37735 5312 37787
rect 5326 37780 5330 37787
rect 5330 37780 5364 37787
rect 5364 37780 5378 37787
rect 5326 37742 5378 37780
rect 5326 37735 5330 37742
rect 5330 37735 5364 37742
rect 5364 37735 5378 37742
rect 5392 37735 5444 37787
rect 4666 37671 4718 37723
rect 4732 37671 4784 37723
rect 4798 37671 4850 37723
rect 4864 37671 4916 37723
rect 4930 37671 4982 37723
rect 4996 37671 5048 37723
rect 5062 37671 5114 37723
rect 5128 37671 5180 37723
rect 5194 37671 5246 37723
rect 5260 37671 5312 37723
rect 5326 37708 5330 37723
rect 5330 37708 5364 37723
rect 5364 37708 5378 37723
rect 5326 37671 5378 37708
rect 5392 37671 5444 37723
rect 4666 37607 4718 37659
rect 4732 37607 4784 37659
rect 4798 37607 4850 37659
rect 4864 37607 4916 37659
rect 4930 37607 4982 37659
rect 4996 37607 5048 37659
rect 5062 37607 5114 37659
rect 5128 37607 5180 37659
rect 5194 37607 5246 37659
rect 5260 37607 5312 37659
rect 5326 37636 5330 37659
rect 5330 37636 5364 37659
rect 5364 37636 5378 37659
rect 5326 37607 5378 37636
rect 5392 37607 5444 37659
rect 4666 37543 4718 37595
rect 4732 37543 4784 37595
rect 4798 37543 4850 37595
rect 4864 37543 4916 37595
rect 4930 37543 4982 37595
rect 4996 37543 5048 37595
rect 5062 37543 5114 37595
rect 5128 37543 5180 37595
rect 5194 37543 5246 37595
rect 5260 37543 5312 37595
rect 5326 37564 5330 37595
rect 5330 37564 5364 37595
rect 5364 37564 5378 37595
rect 5326 37543 5378 37564
rect 5392 37543 5444 37595
rect 4666 37479 4718 37531
rect 4732 37479 4784 37531
rect 4798 37479 4850 37531
rect 4864 37479 4916 37531
rect 4930 37479 4982 37531
rect 4996 37479 5048 37531
rect 5062 37479 5114 37531
rect 5128 37479 5180 37531
rect 5194 37479 5246 37531
rect 5260 37479 5312 37531
rect 5326 37526 5378 37531
rect 5326 37492 5330 37526
rect 5330 37492 5364 37526
rect 5364 37492 5378 37526
rect 5326 37479 5378 37492
rect 5392 37479 5444 37531
rect 4666 37415 4718 37467
rect 4732 37415 4784 37467
rect 4798 37415 4850 37467
rect 4864 37415 4916 37467
rect 4930 37415 4982 37467
rect 4996 37415 5048 37467
rect 5062 37415 5114 37467
rect 5128 37415 5180 37467
rect 5194 37415 5246 37467
rect 5260 37415 5312 37467
rect 5326 37454 5378 37467
rect 5326 37420 5330 37454
rect 5330 37420 5364 37454
rect 5364 37420 5378 37454
rect 5326 37415 5378 37420
rect 5392 37415 5444 37467
rect 4666 37351 4718 37403
rect 4732 37351 4784 37403
rect 4798 37351 4850 37403
rect 4864 37351 4916 37403
rect 4930 37351 4982 37403
rect 4996 37351 5048 37403
rect 5062 37351 5114 37403
rect 5128 37351 5180 37403
rect 5194 37351 5246 37403
rect 5260 37351 5312 37403
rect 5326 37382 5378 37403
rect 5326 37351 5330 37382
rect 5330 37351 5364 37382
rect 5364 37351 5378 37382
rect 5392 37351 5444 37403
rect 4666 37287 4718 37339
rect 4732 37287 4784 37339
rect 4798 37287 4850 37339
rect 4864 37287 4916 37339
rect 4930 37287 4982 37339
rect 4996 37287 5048 37339
rect 5062 37287 5114 37339
rect 5128 37287 5180 37339
rect 5194 37287 5246 37339
rect 5260 37287 5312 37339
rect 5326 37310 5378 37339
rect 5326 37287 5330 37310
rect 5330 37287 5364 37310
rect 5364 37287 5378 37310
rect 5392 37287 5444 37339
rect 4666 37223 4718 37275
rect 4732 37223 4784 37275
rect 4798 37223 4850 37275
rect 4864 37223 4916 37275
rect 4930 37223 4982 37275
rect 4996 37223 5048 37275
rect 5062 37223 5114 37275
rect 5128 37223 5180 37275
rect 5194 37223 5246 37275
rect 5260 37223 5312 37275
rect 5326 37238 5378 37275
rect 5326 37223 5330 37238
rect 5330 37223 5364 37238
rect 5364 37223 5378 37238
rect 5392 37223 5444 37275
rect 4666 37159 4718 37211
rect 4732 37159 4784 37211
rect 4798 37159 4850 37211
rect 4864 37159 4916 37211
rect 4930 37159 4982 37211
rect 4996 37159 5048 37211
rect 5062 37159 5114 37211
rect 5128 37159 5180 37211
rect 5194 37159 5246 37211
rect 5260 37159 5312 37211
rect 5326 37204 5330 37211
rect 5330 37204 5364 37211
rect 5364 37204 5378 37211
rect 5326 37166 5378 37204
rect 5326 37159 5330 37166
rect 5330 37159 5364 37166
rect 5364 37159 5378 37166
rect 5392 37159 5444 37211
rect 4666 37095 4718 37147
rect 4732 37095 4784 37147
rect 4798 37095 4850 37147
rect 4864 37095 4916 37147
rect 4930 37095 4982 37147
rect 4996 37095 5048 37147
rect 5062 37095 5114 37147
rect 5128 37095 5180 37147
rect 5194 37095 5246 37147
rect 5260 37095 5312 37147
rect 5326 37132 5330 37147
rect 5330 37132 5364 37147
rect 5364 37132 5378 37147
rect 5326 37095 5378 37132
rect 5392 37095 5444 37147
rect 4666 37031 4718 37083
rect 4732 37031 4784 37083
rect 4798 37031 4850 37083
rect 4864 37031 4916 37083
rect 4930 37031 4982 37083
rect 4996 37031 5048 37083
rect 5062 37031 5114 37083
rect 5128 37031 5180 37083
rect 5194 37031 5246 37083
rect 5260 37031 5312 37083
rect 5326 37060 5330 37083
rect 5330 37060 5364 37083
rect 5364 37060 5378 37083
rect 5326 37031 5378 37060
rect 5392 37031 5444 37083
rect 4666 36967 4718 37019
rect 4732 36967 4784 37019
rect 4798 36967 4850 37019
rect 4864 36967 4916 37019
rect 4930 36967 4982 37019
rect 4996 36967 5048 37019
rect 5062 36967 5114 37019
rect 5128 36967 5180 37019
rect 5194 36967 5246 37019
rect 5260 36967 5312 37019
rect 5326 36988 5330 37019
rect 5330 36988 5364 37019
rect 5364 36988 5378 37019
rect 5326 36967 5378 36988
rect 5392 36967 5444 37019
rect 4666 36903 4718 36955
rect 4732 36903 4784 36955
rect 4798 36903 4850 36955
rect 4864 36903 4916 36955
rect 4930 36903 4982 36955
rect 4996 36903 5048 36955
rect 5062 36903 5114 36955
rect 5128 36903 5180 36955
rect 5194 36903 5246 36955
rect 5260 36903 5312 36955
rect 5326 36950 5378 36955
rect 5326 36916 5330 36950
rect 5330 36916 5364 36950
rect 5364 36916 5378 36950
rect 5326 36903 5378 36916
rect 5392 36903 5444 36955
rect 4666 36839 4718 36891
rect 4732 36839 4784 36891
rect 4798 36839 4850 36891
rect 4864 36839 4916 36891
rect 4930 36839 4982 36891
rect 4996 36839 5048 36891
rect 5062 36839 5114 36891
rect 5128 36839 5180 36891
rect 5194 36839 5246 36891
rect 5260 36839 5312 36891
rect 5326 36878 5378 36891
rect 5326 36844 5330 36878
rect 5330 36844 5364 36878
rect 5364 36844 5378 36878
rect 5326 36839 5378 36844
rect 5392 36839 5444 36891
rect 4666 36775 4718 36827
rect 4732 36775 4784 36827
rect 4798 36775 4850 36827
rect 4864 36775 4916 36827
rect 4930 36775 4982 36827
rect 4996 36775 5048 36827
rect 5062 36775 5114 36827
rect 5128 36775 5180 36827
rect 5194 36775 5246 36827
rect 5260 36775 5312 36827
rect 5326 36806 5378 36827
rect 5326 36775 5330 36806
rect 5330 36775 5364 36806
rect 5364 36775 5378 36806
rect 5392 36775 5444 36827
rect 4666 36711 4718 36763
rect 4732 36711 4784 36763
rect 4798 36711 4850 36763
rect 4864 36711 4916 36763
rect 4930 36711 4982 36763
rect 4996 36711 5048 36763
rect 5062 36711 5114 36763
rect 5128 36711 5180 36763
rect 5194 36711 5246 36763
rect 5260 36711 5312 36763
rect 5326 36734 5378 36763
rect 5326 36711 5330 36734
rect 5330 36711 5364 36734
rect 5364 36711 5378 36734
rect 5392 36711 5444 36763
rect 4666 36647 4718 36699
rect 4732 36647 4784 36699
rect 4798 36647 4850 36699
rect 4864 36647 4916 36699
rect 4930 36647 4982 36699
rect 4996 36647 5048 36699
rect 5062 36647 5114 36699
rect 5128 36647 5180 36699
rect 5194 36647 5246 36699
rect 5260 36647 5312 36699
rect 5326 36662 5378 36699
rect 5326 36647 5330 36662
rect 5330 36647 5364 36662
rect 5364 36647 5378 36662
rect 5392 36647 5444 36699
rect 4666 36583 4718 36635
rect 4732 36583 4784 36635
rect 4798 36583 4850 36635
rect 4864 36583 4916 36635
rect 4930 36583 4982 36635
rect 4996 36583 5048 36635
rect 5062 36583 5114 36635
rect 5128 36583 5180 36635
rect 5194 36583 5246 36635
rect 5260 36583 5312 36635
rect 5326 36628 5330 36635
rect 5330 36628 5364 36635
rect 5364 36628 5378 36635
rect 5326 36590 5378 36628
rect 5326 36583 5330 36590
rect 5330 36583 5364 36590
rect 5364 36583 5378 36590
rect 5392 36583 5444 36635
rect 4666 36519 4718 36571
rect 4732 36519 4784 36571
rect 4798 36519 4850 36571
rect 4864 36519 4916 36571
rect 4930 36519 4982 36571
rect 4996 36519 5048 36571
rect 5062 36519 5114 36571
rect 5128 36519 5180 36571
rect 5194 36519 5246 36571
rect 5260 36519 5312 36571
rect 5326 36556 5330 36571
rect 5330 36556 5364 36571
rect 5364 36556 5378 36571
rect 5326 36519 5378 36556
rect 5392 36519 5444 36571
rect 4666 36455 4718 36507
rect 4732 36455 4784 36507
rect 4798 36455 4850 36507
rect 4864 36455 4916 36507
rect 4930 36455 4982 36507
rect 4996 36455 5048 36507
rect 5062 36455 5114 36507
rect 5128 36455 5180 36507
rect 5194 36455 5246 36507
rect 5260 36455 5312 36507
rect 5326 36484 5330 36507
rect 5330 36484 5364 36507
rect 5364 36484 5378 36507
rect 5326 36455 5378 36484
rect 5392 36455 5444 36507
rect 4666 36391 4718 36443
rect 4732 36391 4784 36443
rect 4798 36391 4850 36443
rect 4864 36391 4916 36443
rect 4930 36391 4982 36443
rect 4996 36391 5048 36443
rect 5062 36391 5114 36443
rect 5128 36391 5180 36443
rect 5194 36391 5246 36443
rect 5260 36391 5312 36443
rect 5326 36412 5330 36443
rect 5330 36412 5364 36443
rect 5364 36412 5378 36443
rect 5326 36391 5378 36412
rect 5392 36391 5444 36443
rect 4666 36327 4718 36379
rect 4732 36327 4784 36379
rect 4798 36327 4850 36379
rect 4864 36327 4916 36379
rect 4930 36327 4982 36379
rect 4996 36327 5048 36379
rect 5062 36327 5114 36379
rect 5128 36327 5180 36379
rect 5194 36327 5246 36379
rect 5260 36327 5312 36379
rect 5326 36374 5378 36379
rect 5326 36340 5330 36374
rect 5330 36340 5364 36374
rect 5364 36340 5378 36374
rect 5326 36327 5378 36340
rect 5392 36327 5444 36379
rect 4666 36263 4718 36315
rect 4732 36263 4784 36315
rect 4798 36263 4850 36315
rect 4864 36263 4916 36315
rect 4930 36263 4982 36315
rect 4996 36263 5048 36315
rect 5062 36263 5114 36315
rect 5128 36263 5180 36315
rect 5194 36263 5246 36315
rect 5260 36263 5312 36315
rect 5326 36302 5378 36315
rect 5326 36268 5330 36302
rect 5330 36268 5364 36302
rect 5364 36268 5378 36302
rect 5326 36263 5378 36268
rect 5392 36263 5444 36315
rect 4666 36199 4718 36251
rect 4732 36199 4784 36251
rect 4798 36199 4850 36251
rect 4864 36199 4916 36251
rect 4930 36199 4982 36251
rect 4996 36199 5048 36251
rect 5062 36199 5114 36251
rect 5128 36199 5180 36251
rect 5194 36199 5246 36251
rect 5260 36199 5312 36251
rect 5326 36230 5378 36251
rect 5326 36199 5330 36230
rect 5330 36199 5364 36230
rect 5364 36199 5378 36230
rect 5392 36199 5444 36251
rect 4666 36135 4718 36187
rect 4732 36135 4784 36187
rect 4798 36135 4850 36187
rect 4864 36135 4916 36187
rect 4930 36135 4982 36187
rect 4996 36135 5048 36187
rect 5062 36135 5114 36187
rect 5128 36135 5180 36187
rect 5194 36135 5246 36187
rect 5260 36135 5312 36187
rect 5326 36158 5378 36187
rect 5326 36135 5330 36158
rect 5330 36135 5364 36158
rect 5364 36135 5378 36158
rect 5392 36135 5444 36187
rect 4666 36071 4718 36123
rect 4732 36071 4784 36123
rect 4798 36071 4850 36123
rect 4864 36071 4916 36123
rect 4930 36071 4982 36123
rect 4996 36071 5048 36123
rect 5062 36071 5114 36123
rect 5128 36071 5180 36123
rect 5194 36071 5246 36123
rect 5260 36071 5312 36123
rect 5326 36086 5378 36123
rect 5326 36071 5330 36086
rect 5330 36071 5364 36086
rect 5364 36071 5378 36086
rect 5392 36071 5444 36123
rect 4666 36007 4718 36059
rect 4732 36007 4784 36059
rect 4798 36007 4850 36059
rect 4864 36007 4916 36059
rect 4930 36007 4982 36059
rect 4996 36007 5048 36059
rect 5062 36007 5114 36059
rect 5128 36007 5180 36059
rect 5194 36007 5246 36059
rect 5260 36007 5312 36059
rect 5326 36052 5330 36059
rect 5330 36052 5364 36059
rect 5364 36052 5378 36059
rect 5326 36014 5378 36052
rect 5326 36007 5330 36014
rect 5330 36007 5364 36014
rect 5364 36007 5378 36014
rect 5392 36007 5444 36059
rect 4666 35943 4718 35995
rect 4732 35943 4784 35995
rect 4798 35943 4850 35995
rect 4864 35943 4916 35995
rect 4930 35943 4982 35995
rect 4996 35943 5048 35995
rect 5062 35943 5114 35995
rect 5128 35943 5180 35995
rect 5194 35943 5246 35995
rect 5260 35943 5312 35995
rect 5326 35980 5330 35995
rect 5330 35980 5364 35995
rect 5364 35980 5378 35995
rect 5326 35943 5378 35980
rect 5392 35943 5444 35995
rect 4666 35879 4718 35931
rect 4732 35879 4784 35931
rect 4798 35879 4850 35931
rect 4864 35879 4916 35931
rect 4930 35879 4982 35931
rect 4996 35879 5048 35931
rect 5062 35879 5114 35931
rect 5128 35879 5180 35931
rect 5194 35879 5246 35931
rect 5260 35879 5312 35931
rect 5326 35908 5330 35931
rect 5330 35908 5364 35931
rect 5364 35908 5378 35931
rect 5326 35879 5378 35908
rect 5392 35879 5444 35931
rect 4666 35815 4718 35867
rect 4732 35815 4784 35867
rect 4798 35815 4850 35867
rect 4864 35815 4916 35867
rect 4930 35815 4982 35867
rect 4996 35815 5048 35867
rect 5062 35815 5114 35867
rect 5128 35815 5180 35867
rect 5194 35815 5246 35867
rect 5260 35815 5312 35867
rect 5326 35836 5330 35867
rect 5330 35836 5364 35867
rect 5364 35836 5378 35867
rect 5326 35815 5378 35836
rect 5392 35815 5444 35867
rect 4666 35751 4718 35803
rect 4732 35751 4784 35803
rect 4798 35751 4850 35803
rect 4864 35751 4916 35803
rect 4930 35751 4982 35803
rect 4996 35751 5048 35803
rect 5062 35751 5114 35803
rect 5128 35751 5180 35803
rect 5194 35751 5246 35803
rect 5260 35751 5312 35803
rect 5326 35798 5378 35803
rect 5326 35764 5330 35798
rect 5330 35764 5364 35798
rect 5364 35764 5378 35798
rect 5326 35751 5378 35764
rect 5392 35751 5444 35803
rect 4666 35687 4718 35739
rect 4732 35687 4784 35739
rect 4798 35687 4850 35739
rect 4864 35687 4916 35739
rect 4930 35687 4982 35739
rect 4996 35687 5048 35739
rect 5062 35687 5114 35739
rect 5128 35687 5180 35739
rect 5194 35687 5246 35739
rect 5260 35687 5312 35739
rect 5326 35726 5378 35739
rect 5326 35692 5330 35726
rect 5330 35692 5364 35726
rect 5364 35692 5378 35726
rect 5326 35687 5378 35692
rect 5392 35687 5444 35739
rect 3165 35609 3217 35643
rect 3165 35591 3174 35609
rect 3174 35591 3208 35609
rect 3208 35591 3217 35609
rect 3165 35575 3174 35579
rect 3174 35575 3208 35579
rect 3208 35575 3217 35579
rect 3165 35537 3217 35575
rect 3165 35527 3174 35537
rect 3174 35527 3208 35537
rect 3208 35527 3217 35537
rect 4666 35623 4718 35675
rect 4732 35623 4784 35675
rect 4798 35623 4850 35675
rect 4864 35623 4916 35675
rect 4930 35623 4982 35675
rect 4996 35623 5048 35675
rect 5062 35623 5114 35675
rect 5128 35623 5180 35675
rect 5194 35623 5246 35675
rect 5260 35623 5312 35675
rect 5326 35654 5378 35675
rect 5326 35623 5330 35654
rect 5330 35623 5364 35654
rect 5364 35623 5378 35654
rect 5392 35623 5444 35675
rect 4666 35559 4718 35611
rect 4732 35559 4784 35611
rect 4798 35559 4850 35611
rect 4864 35559 4916 35611
rect 4930 35559 4982 35611
rect 4996 35559 5048 35611
rect 5062 35559 5114 35611
rect 5128 35559 5180 35611
rect 5194 35559 5246 35611
rect 5260 35559 5312 35611
rect 5326 35582 5378 35611
rect 5326 35559 5330 35582
rect 5330 35559 5364 35582
rect 5364 35559 5378 35582
rect 5392 35559 5444 35611
rect 4666 35495 4718 35547
rect 4732 35495 4784 35547
rect 4798 35495 4850 35547
rect 4864 35495 4916 35547
rect 4930 35495 4982 35547
rect 4996 35495 5048 35547
rect 5062 35495 5114 35547
rect 5128 35495 5180 35547
rect 5194 35495 5246 35547
rect 5260 35495 5312 35547
rect 5326 35510 5378 35547
rect 5326 35495 5330 35510
rect 5330 35495 5364 35510
rect 5364 35495 5378 35510
rect 5392 35495 5444 35547
rect 4666 35431 4718 35483
rect 4732 35431 4784 35483
rect 4798 35431 4850 35483
rect 4864 35431 4916 35483
rect 4930 35431 4982 35483
rect 4996 35431 5048 35483
rect 5062 35431 5114 35483
rect 5128 35431 5180 35483
rect 5194 35431 5246 35483
rect 5260 35431 5312 35483
rect 5326 35476 5330 35483
rect 5330 35476 5364 35483
rect 5364 35476 5378 35483
rect 5326 35438 5378 35476
rect 5326 35431 5330 35438
rect 5330 35431 5364 35438
rect 5364 35431 5378 35438
rect 5392 35431 5444 35483
rect 4666 35367 4718 35419
rect 4732 35367 4784 35419
rect 4798 35367 4850 35419
rect 4864 35367 4916 35419
rect 4930 35367 4982 35419
rect 4996 35367 5048 35419
rect 5062 35367 5114 35419
rect 5128 35367 5180 35419
rect 5194 35367 5246 35419
rect 5260 35367 5312 35419
rect 5326 35404 5330 35419
rect 5330 35404 5364 35419
rect 5364 35404 5378 35419
rect 5326 35367 5378 35404
rect 5392 35367 5444 35419
rect 4666 35303 4718 35355
rect 4732 35303 4784 35355
rect 4798 35303 4850 35355
rect 4864 35303 4916 35355
rect 4930 35303 4982 35355
rect 4996 35303 5048 35355
rect 5062 35303 5114 35355
rect 5128 35303 5180 35355
rect 5194 35303 5246 35355
rect 5260 35303 5312 35355
rect 5326 35332 5330 35355
rect 5330 35332 5364 35355
rect 5364 35332 5378 35355
rect 5326 35303 5378 35332
rect 5392 35303 5444 35355
rect 4666 35239 4718 35291
rect 4732 35239 4784 35291
rect 4798 35239 4850 35291
rect 4864 35239 4916 35291
rect 4930 35239 4982 35291
rect 4996 35239 5048 35291
rect 5062 35239 5114 35291
rect 5128 35239 5180 35291
rect 5194 35239 5246 35291
rect 5260 35239 5312 35291
rect 5326 35260 5330 35291
rect 5330 35260 5364 35291
rect 5364 35260 5378 35291
rect 5326 35239 5378 35260
rect 5392 35239 5444 35291
rect 4666 35175 4718 35227
rect 4732 35175 4784 35227
rect 4798 35175 4850 35227
rect 4864 35175 4916 35227
rect 4930 35175 4982 35227
rect 4996 35175 5048 35227
rect 5062 35175 5114 35227
rect 5128 35175 5180 35227
rect 5194 35175 5246 35227
rect 5260 35175 5312 35227
rect 5326 35222 5378 35227
rect 5326 35188 5330 35222
rect 5330 35188 5364 35222
rect 5364 35188 5378 35222
rect 5326 35175 5378 35188
rect 5392 35175 5444 35227
rect 4666 35111 4718 35163
rect 4732 35111 4784 35163
rect 4798 35111 4850 35163
rect 4864 35111 4916 35163
rect 4930 35111 4982 35163
rect 4996 35111 5048 35163
rect 5062 35111 5114 35163
rect 5128 35111 5180 35163
rect 5194 35111 5246 35163
rect 5260 35111 5312 35163
rect 5326 35149 5378 35163
rect 5326 35115 5330 35149
rect 5330 35115 5364 35149
rect 5364 35115 5378 35149
rect 5326 35111 5378 35115
rect 5392 35111 5444 35163
rect 4666 35047 4718 35099
rect 4732 35047 4784 35099
rect 4798 35047 4850 35099
rect 4864 35047 4916 35099
rect 4930 35047 4982 35099
rect 4996 35047 5048 35099
rect 5062 35047 5114 35099
rect 5128 35047 5180 35099
rect 5194 35047 5246 35099
rect 5260 35047 5312 35099
rect 5326 35076 5378 35099
rect 5326 35047 5330 35076
rect 5330 35047 5364 35076
rect 5364 35047 5378 35076
rect 5392 35047 5444 35099
rect 4666 34983 4718 35035
rect 4732 34983 4784 35035
rect 4798 34983 4850 35035
rect 4864 34983 4916 35035
rect 4930 34983 4982 35035
rect 4996 34983 5048 35035
rect 5062 34983 5114 35035
rect 5128 34983 5180 35035
rect 5194 34983 5246 35035
rect 5260 34983 5312 35035
rect 5326 35003 5378 35035
rect 5326 34983 5330 35003
rect 5330 34983 5364 35003
rect 5364 34983 5378 35003
rect 5392 34983 5444 35035
rect 4666 34919 4718 34971
rect 4732 34919 4784 34971
rect 4798 34919 4850 34971
rect 4864 34919 4916 34971
rect 4930 34919 4982 34971
rect 4996 34919 5048 34971
rect 5062 34919 5114 34971
rect 5128 34919 5180 34971
rect 5194 34919 5246 34971
rect 5260 34919 5312 34971
rect 5326 34969 5330 34971
rect 5330 34969 5364 34971
rect 5364 34969 5378 34971
rect 5326 34930 5378 34969
rect 5326 34919 5330 34930
rect 5330 34919 5364 34930
rect 5364 34919 5378 34930
rect 5392 34919 5444 34971
rect 4666 34855 4718 34907
rect 4732 34855 4784 34907
rect 4798 34855 4850 34907
rect 4864 34855 4916 34907
rect 4930 34855 4982 34907
rect 4996 34855 5048 34907
rect 5062 34855 5114 34907
rect 5128 34855 5180 34907
rect 5194 34855 5246 34907
rect 5260 34855 5312 34907
rect 5326 34896 5330 34907
rect 5330 34896 5364 34907
rect 5364 34896 5378 34907
rect 5326 34857 5378 34896
rect 5326 34855 5330 34857
rect 5330 34855 5364 34857
rect 5364 34855 5378 34857
rect 5392 34855 5444 34907
rect 4666 34791 4718 34843
rect 4732 34791 4784 34843
rect 4798 34791 4850 34843
rect 4864 34791 4916 34843
rect 4930 34791 4982 34843
rect 4996 34791 5048 34843
rect 5062 34791 5114 34843
rect 5128 34791 5180 34843
rect 5194 34791 5246 34843
rect 5260 34791 5312 34843
rect 5326 34823 5330 34843
rect 5330 34823 5364 34843
rect 5364 34823 5378 34843
rect 5326 34791 5378 34823
rect 5392 34791 5444 34843
rect 4666 34727 4718 34779
rect 4732 34727 4784 34779
rect 4798 34727 4850 34779
rect 4864 34727 4916 34779
rect 4930 34727 4982 34779
rect 4996 34727 5048 34779
rect 5062 34727 5114 34779
rect 5128 34727 5180 34779
rect 5194 34727 5246 34779
rect 5260 34727 5312 34779
rect 5326 34750 5330 34779
rect 5330 34750 5364 34779
rect 5364 34750 5378 34779
rect 5326 34727 5378 34750
rect 5392 34727 5444 34779
rect 4666 34663 4718 34715
rect 4732 34663 4784 34715
rect 4798 34663 4850 34715
rect 4864 34663 4916 34715
rect 4930 34663 4982 34715
rect 4996 34663 5048 34715
rect 5062 34663 5114 34715
rect 5128 34663 5180 34715
rect 5194 34663 5246 34715
rect 5260 34663 5312 34715
rect 5326 34711 5378 34715
rect 5326 34677 5330 34711
rect 5330 34677 5364 34711
rect 5364 34677 5378 34711
rect 5326 34663 5378 34677
rect 5392 34663 5444 34715
rect 4666 34599 4718 34651
rect 4732 34599 4784 34651
rect 4798 34599 4850 34651
rect 4864 34599 4916 34651
rect 4930 34599 4982 34651
rect 4996 34599 5048 34651
rect 5062 34599 5114 34651
rect 5128 34599 5180 34651
rect 5194 34599 5246 34651
rect 5260 34599 5312 34651
rect 5326 34638 5378 34651
rect 5326 34604 5330 34638
rect 5330 34604 5364 34638
rect 5364 34604 5378 34638
rect 5326 34599 5378 34604
rect 5392 34599 5444 34651
rect 4666 34535 4718 34587
rect 4732 34535 4784 34587
rect 4798 34535 4850 34587
rect 4864 34535 4916 34587
rect 4930 34535 4982 34587
rect 4996 34535 5048 34587
rect 5062 34535 5114 34587
rect 5128 34535 5180 34587
rect 5194 34535 5246 34587
rect 5260 34535 5312 34587
rect 5326 34565 5378 34587
rect 5326 34535 5330 34565
rect 5330 34535 5364 34565
rect 5364 34535 5378 34565
rect 5392 34535 5444 34587
rect 4666 34471 4718 34523
rect 4732 34471 4784 34523
rect 4798 34471 4850 34523
rect 4864 34471 4916 34523
rect 4930 34471 4982 34523
rect 4996 34471 5048 34523
rect 5062 34471 5114 34523
rect 5128 34471 5180 34523
rect 5194 34471 5246 34523
rect 5260 34471 5312 34523
rect 5326 34492 5378 34523
rect 5326 34471 5330 34492
rect 5330 34471 5364 34492
rect 5364 34471 5378 34492
rect 5392 34471 5444 34523
rect 4666 34407 4718 34459
rect 4732 34407 4784 34459
rect 4798 34407 4850 34459
rect 4864 34407 4916 34459
rect 4930 34407 4982 34459
rect 4996 34407 5048 34459
rect 5062 34407 5114 34459
rect 5128 34407 5180 34459
rect 5194 34407 5246 34459
rect 5260 34407 5312 34459
rect 5326 34458 5330 34459
rect 5330 34458 5364 34459
rect 5364 34458 5378 34459
rect 5326 34419 5378 34458
rect 5326 34407 5330 34419
rect 5330 34407 5364 34419
rect 5364 34407 5378 34419
rect 5392 34407 5444 34459
rect 4666 34343 4718 34395
rect 4732 34343 4784 34395
rect 4798 34343 4850 34395
rect 4864 34343 4916 34395
rect 4930 34343 4982 34395
rect 4996 34343 5048 34395
rect 5062 34343 5114 34395
rect 5128 34343 5180 34395
rect 5194 34343 5246 34395
rect 5260 34343 5312 34395
rect 5326 34385 5330 34395
rect 5330 34385 5364 34395
rect 5364 34385 5378 34395
rect 5326 34346 5378 34385
rect 5326 34343 5330 34346
rect 5330 34343 5364 34346
rect 5364 34343 5378 34346
rect 5392 34343 5444 34395
rect 4666 34279 4718 34331
rect 4732 34279 4784 34331
rect 4798 34279 4850 34331
rect 4864 34279 4916 34331
rect 4930 34279 4982 34331
rect 4996 34279 5048 34331
rect 5062 34279 5114 34331
rect 5128 34279 5180 34331
rect 5194 34279 5246 34331
rect 5260 34279 5312 34331
rect 5326 34312 5330 34331
rect 5330 34312 5364 34331
rect 5364 34312 5378 34331
rect 5326 34279 5378 34312
rect 5392 34279 5444 34331
rect 4666 34215 4718 34267
rect 4732 34215 4784 34267
rect 4798 34215 4850 34267
rect 4864 34215 4916 34267
rect 4930 34215 4982 34267
rect 4996 34215 5048 34267
rect 5062 34215 5114 34267
rect 5128 34215 5180 34267
rect 5194 34215 5246 34267
rect 5260 34215 5312 34267
rect 5326 34239 5330 34267
rect 5330 34239 5364 34267
rect 5364 34239 5378 34267
rect 5326 34215 5378 34239
rect 5392 34215 5444 34267
rect 4666 34151 4718 34203
rect 4732 34151 4784 34203
rect 4798 34151 4850 34203
rect 4864 34151 4916 34203
rect 4930 34151 4982 34203
rect 4996 34151 5048 34203
rect 5062 34151 5114 34203
rect 5128 34151 5180 34203
rect 5194 34151 5246 34203
rect 5260 34151 5312 34203
rect 5326 34200 5378 34203
rect 5326 34166 5330 34200
rect 5330 34166 5364 34200
rect 5364 34166 5378 34200
rect 5326 34151 5378 34166
rect 5392 34151 5444 34203
rect 4666 34087 4718 34139
rect 4732 34087 4784 34139
rect 4798 34087 4850 34139
rect 4864 34087 4916 34139
rect 4930 34087 4982 34139
rect 4996 34087 5048 34139
rect 5062 34087 5114 34139
rect 5128 34087 5180 34139
rect 5194 34087 5246 34139
rect 5260 34087 5312 34139
rect 5326 34127 5378 34139
rect 5326 34093 5330 34127
rect 5330 34093 5364 34127
rect 5364 34093 5378 34127
rect 5326 34087 5378 34093
rect 5392 34087 5444 34139
rect 4666 34023 4718 34075
rect 4732 34023 4784 34075
rect 4798 34023 4850 34075
rect 4864 34023 4916 34075
rect 4930 34023 4982 34075
rect 4996 34023 5048 34075
rect 5062 34023 5114 34075
rect 5128 34023 5180 34075
rect 5194 34023 5246 34075
rect 5260 34023 5312 34075
rect 5326 34054 5378 34075
rect 5326 34023 5330 34054
rect 5330 34023 5364 34054
rect 5364 34023 5378 34054
rect 5392 34023 5444 34075
rect 4666 33959 4718 34011
rect 4732 33959 4784 34011
rect 4798 33959 4850 34011
rect 4864 33959 4916 34011
rect 4930 33959 4982 34011
rect 4996 33959 5048 34011
rect 5062 33959 5114 34011
rect 5128 33959 5180 34011
rect 5194 33959 5246 34011
rect 5260 33959 5312 34011
rect 5326 33981 5378 34011
rect 5326 33959 5330 33981
rect 5330 33959 5364 33981
rect 5364 33959 5378 33981
rect 5392 33959 5444 34011
rect 4666 33895 4718 33947
rect 4732 33895 4784 33947
rect 4798 33895 4850 33947
rect 4864 33895 4916 33947
rect 4930 33895 4982 33947
rect 4996 33895 5048 33947
rect 5062 33895 5114 33947
rect 5128 33895 5180 33947
rect 5194 33895 5246 33947
rect 5260 33895 5312 33947
rect 5326 33908 5378 33947
rect 5326 33895 5330 33908
rect 5330 33895 5364 33908
rect 5364 33895 5378 33908
rect 5392 33895 5444 33947
rect 4666 33831 4718 33883
rect 4732 33831 4784 33883
rect 4798 33831 4850 33883
rect 4864 33831 4916 33883
rect 4930 33831 4982 33883
rect 4996 33831 5048 33883
rect 5062 33831 5114 33883
rect 5128 33831 5180 33883
rect 5194 33831 5246 33883
rect 5260 33831 5312 33883
rect 5326 33874 5330 33883
rect 5330 33874 5364 33883
rect 5364 33874 5378 33883
rect 5326 33835 5378 33874
rect 5326 33831 5330 33835
rect 5330 33831 5364 33835
rect 5364 33831 5378 33835
rect 5392 33831 5444 33883
rect 4666 33767 4718 33819
rect 4732 33767 4784 33819
rect 4798 33767 4850 33819
rect 4864 33767 4916 33819
rect 4930 33767 4982 33819
rect 4996 33767 5048 33819
rect 5062 33767 5114 33819
rect 5128 33767 5180 33819
rect 5194 33767 5246 33819
rect 5260 33767 5312 33819
rect 5326 33801 5330 33819
rect 5330 33801 5364 33819
rect 5364 33801 5378 33819
rect 5326 33767 5378 33801
rect 5392 33767 5444 33819
rect 4666 33703 4718 33755
rect 4732 33703 4784 33755
rect 4798 33703 4850 33755
rect 4864 33703 4916 33755
rect 4930 33703 4982 33755
rect 4996 33703 5048 33755
rect 5062 33703 5114 33755
rect 5128 33703 5180 33755
rect 5194 33703 5246 33755
rect 5260 33703 5312 33755
rect 5326 33728 5330 33755
rect 5330 33728 5364 33755
rect 5364 33728 5378 33755
rect 5326 33703 5378 33728
rect 5392 33703 5444 33755
rect 4666 33639 4718 33691
rect 4732 33639 4784 33691
rect 4798 33639 4850 33691
rect 4864 33639 4916 33691
rect 4930 33639 4982 33691
rect 4996 33639 5048 33691
rect 5062 33639 5114 33691
rect 5128 33639 5180 33691
rect 5194 33639 5246 33691
rect 5260 33639 5312 33691
rect 5326 33689 5378 33691
rect 5326 33655 5330 33689
rect 5330 33655 5364 33689
rect 5364 33655 5378 33689
rect 5326 33639 5378 33655
rect 5392 33639 5444 33691
rect 4666 33575 4718 33627
rect 4732 33575 4784 33627
rect 4798 33575 4850 33627
rect 4864 33575 4916 33627
rect 4930 33575 4982 33627
rect 4996 33575 5048 33627
rect 5062 33575 5114 33627
rect 5128 33575 5180 33627
rect 5194 33575 5246 33627
rect 5260 33575 5312 33627
rect 5326 33616 5378 33627
rect 5326 33582 5330 33616
rect 5330 33582 5364 33616
rect 5364 33582 5378 33616
rect 5326 33575 5378 33582
rect 5392 33575 5444 33627
rect 4666 33511 4718 33563
rect 4732 33511 4784 33563
rect 4798 33511 4850 33563
rect 4864 33511 4916 33563
rect 4930 33511 4982 33563
rect 4996 33511 5048 33563
rect 5062 33511 5114 33563
rect 5128 33511 5180 33563
rect 5194 33511 5246 33563
rect 5260 33511 5312 33563
rect 5326 33543 5378 33563
rect 5326 33511 5330 33543
rect 5330 33511 5364 33543
rect 5364 33511 5378 33543
rect 5392 33511 5444 33563
rect 4666 33447 4718 33499
rect 4732 33447 4784 33499
rect 4798 33447 4850 33499
rect 4864 33447 4916 33499
rect 4930 33447 4982 33499
rect 4996 33447 5048 33499
rect 5062 33447 5114 33499
rect 5128 33447 5180 33499
rect 5194 33447 5246 33499
rect 5260 33447 5312 33499
rect 5326 33470 5378 33499
rect 5326 33447 5330 33470
rect 5330 33447 5364 33470
rect 5364 33447 5378 33470
rect 5392 33447 5444 33499
rect 4666 33383 4718 33435
rect 4732 33383 4784 33435
rect 4798 33383 4850 33435
rect 4864 33383 4916 33435
rect 4930 33383 4982 33435
rect 4996 33383 5048 33435
rect 5062 33383 5114 33435
rect 5128 33383 5180 33435
rect 5194 33383 5246 33435
rect 5260 33383 5312 33435
rect 5326 33397 5378 33435
rect 5326 33383 5330 33397
rect 5330 33383 5364 33397
rect 5364 33383 5378 33397
rect 5392 33383 5444 33435
rect 4666 33319 4718 33371
rect 4732 33319 4784 33371
rect 4798 33319 4850 33371
rect 4864 33319 4916 33371
rect 4930 33319 4982 33371
rect 4996 33319 5048 33371
rect 5062 33319 5114 33371
rect 5128 33319 5180 33371
rect 5194 33319 5246 33371
rect 5260 33319 5312 33371
rect 5326 33363 5330 33371
rect 5330 33363 5364 33371
rect 5364 33363 5378 33371
rect 5326 33324 5378 33363
rect 5326 33319 5330 33324
rect 5330 33319 5364 33324
rect 5364 33319 5378 33324
rect 5392 33319 5444 33371
rect 4666 33255 4718 33307
rect 4732 33255 4784 33307
rect 4798 33255 4850 33307
rect 4864 33255 4916 33307
rect 4930 33255 4982 33307
rect 4996 33255 5048 33307
rect 5062 33255 5114 33307
rect 5128 33255 5180 33307
rect 5194 33255 5246 33307
rect 5260 33255 5312 33307
rect 5326 33290 5330 33307
rect 5330 33290 5364 33307
rect 5364 33290 5378 33307
rect 5326 33255 5378 33290
rect 5392 33255 5444 33307
rect 4666 33191 4718 33243
rect 4732 33191 4784 33243
rect 4798 33191 4850 33243
rect 4864 33191 4916 33243
rect 4930 33191 4982 33243
rect 4996 33191 5048 33243
rect 5062 33191 5114 33243
rect 5128 33191 5180 33243
rect 5194 33191 5246 33243
rect 5260 33191 5312 33243
rect 5326 33217 5330 33243
rect 5330 33217 5364 33243
rect 5364 33217 5378 33243
rect 5326 33191 5378 33217
rect 5392 33191 5444 33243
rect 4666 33127 4718 33179
rect 4732 33127 4784 33179
rect 4798 33127 4850 33179
rect 4864 33127 4916 33179
rect 4930 33127 4982 33179
rect 4996 33127 5048 33179
rect 5062 33127 5114 33179
rect 5128 33127 5180 33179
rect 5194 33127 5246 33179
rect 5260 33127 5312 33179
rect 5326 33178 5378 33179
rect 5326 33144 5330 33178
rect 5330 33144 5364 33178
rect 5364 33144 5378 33178
rect 5326 33127 5378 33144
rect 5392 33127 5444 33179
rect 4666 33063 4718 33115
rect 4732 33063 4784 33115
rect 4798 33063 4850 33115
rect 4864 33063 4916 33115
rect 4930 33063 4982 33115
rect 4996 33063 5048 33115
rect 5062 33063 5114 33115
rect 5128 33063 5180 33115
rect 5194 33063 5246 33115
rect 5260 33063 5312 33115
rect 5326 33105 5378 33115
rect 5326 33071 5330 33105
rect 5330 33071 5364 33105
rect 5364 33071 5378 33105
rect 5326 33063 5378 33071
rect 5392 33063 5444 33115
rect 4666 32999 4718 33051
rect 4732 32999 4784 33051
rect 4798 32999 4850 33051
rect 4864 32999 4916 33051
rect 4930 32999 4982 33051
rect 4996 32999 5048 33051
rect 5062 32999 5114 33051
rect 5128 32999 5180 33051
rect 5194 32999 5246 33051
rect 5260 32999 5312 33051
rect 5326 33032 5378 33051
rect 5326 32999 5330 33032
rect 5330 32999 5364 33032
rect 5364 32999 5378 33032
rect 5392 32999 5444 33051
rect 4666 32935 4718 32987
rect 4732 32935 4784 32987
rect 4798 32935 4850 32987
rect 4864 32935 4916 32987
rect 4930 32935 4982 32987
rect 4996 32935 5048 32987
rect 5062 32935 5114 32987
rect 5128 32935 5180 32987
rect 5194 32935 5246 32987
rect 5260 32935 5312 32987
rect 5326 32959 5378 32987
rect 5326 32935 5330 32959
rect 5330 32935 5364 32959
rect 5364 32935 5378 32959
rect 5392 32935 5444 32987
rect 4666 32871 4718 32923
rect 4732 32871 4784 32923
rect 4798 32871 4850 32923
rect 4864 32871 4916 32923
rect 4930 32871 4982 32923
rect 4996 32871 5048 32923
rect 5062 32871 5114 32923
rect 5128 32871 5180 32923
rect 5194 32871 5246 32923
rect 5260 32871 5312 32923
rect 5326 32886 5378 32923
rect 5326 32871 5330 32886
rect 5330 32871 5364 32886
rect 5364 32871 5378 32886
rect 5392 32871 5444 32923
rect 4666 32807 4718 32859
rect 4732 32807 4784 32859
rect 4798 32807 4850 32859
rect 4864 32807 4916 32859
rect 4930 32807 4982 32859
rect 4996 32807 5048 32859
rect 5062 32807 5114 32859
rect 5128 32807 5180 32859
rect 5194 32807 5246 32859
rect 5260 32807 5312 32859
rect 5326 32852 5330 32859
rect 5330 32852 5364 32859
rect 5364 32852 5378 32859
rect 5326 32813 5378 32852
rect 5326 32807 5330 32813
rect 5330 32807 5364 32813
rect 5364 32807 5378 32813
rect 5392 32807 5444 32859
rect 4666 32743 4718 32795
rect 4732 32743 4784 32795
rect 4798 32743 4850 32795
rect 4864 32743 4916 32795
rect 4930 32743 4982 32795
rect 4996 32743 5048 32795
rect 5062 32743 5114 32795
rect 5128 32743 5180 32795
rect 5194 32743 5246 32795
rect 5260 32743 5312 32795
rect 5326 32779 5330 32795
rect 5330 32779 5364 32795
rect 5364 32779 5378 32795
rect 5326 32743 5378 32779
rect 5392 32743 5444 32795
rect 4666 32678 4718 32730
rect 4732 32678 4784 32730
rect 4798 32678 4850 32730
rect 4864 32678 4916 32730
rect 4930 32678 4982 32730
rect 4996 32678 5048 32730
rect 5062 32678 5114 32730
rect 5128 32678 5180 32730
rect 5194 32678 5246 32730
rect 5260 32678 5312 32730
rect 5326 32706 5330 32730
rect 5330 32706 5364 32730
rect 5364 32706 5378 32730
rect 5326 32678 5378 32706
rect 5392 32678 5444 32730
rect 4666 32613 4718 32665
rect 4732 32613 4784 32665
rect 4798 32613 4850 32665
rect 4864 32613 4916 32665
rect 4930 32613 4982 32665
rect 4996 32613 5048 32665
rect 5062 32613 5114 32665
rect 5128 32613 5180 32665
rect 5194 32613 5246 32665
rect 5260 32613 5312 32665
rect 5326 32633 5330 32665
rect 5330 32633 5364 32665
rect 5364 32633 5378 32665
rect 5326 32613 5378 32633
rect 5392 32613 5444 32665
rect 4666 32548 4718 32600
rect 4732 32548 4784 32600
rect 4798 32548 4850 32600
rect 4864 32548 4916 32600
rect 4930 32548 4982 32600
rect 4996 32548 5048 32600
rect 5062 32548 5114 32600
rect 5128 32548 5180 32600
rect 5194 32548 5246 32600
rect 5260 32548 5312 32600
rect 5326 32594 5378 32600
rect 5326 32560 5330 32594
rect 5330 32560 5364 32594
rect 5364 32560 5378 32594
rect 5326 32548 5378 32560
rect 5392 32548 5444 32600
rect 4666 32483 4718 32535
rect 4732 32483 4784 32535
rect 4798 32483 4850 32535
rect 4864 32483 4916 32535
rect 4930 32483 4982 32535
rect 4996 32483 5048 32535
rect 5062 32483 5114 32535
rect 5128 32483 5180 32535
rect 5194 32483 5246 32535
rect 5260 32483 5312 32535
rect 5326 32521 5378 32535
rect 5326 32487 5330 32521
rect 5330 32487 5364 32521
rect 5364 32487 5378 32521
rect 5326 32483 5378 32487
rect 5392 32483 5444 32535
rect 4666 32418 4718 32470
rect 4732 32418 4784 32470
rect 4798 32418 4850 32470
rect 4864 32418 4916 32470
rect 4930 32418 4982 32470
rect 4996 32418 5048 32470
rect 5062 32418 5114 32470
rect 5128 32418 5180 32470
rect 5194 32418 5246 32470
rect 5260 32418 5312 32470
rect 5326 32448 5378 32470
rect 5326 32418 5330 32448
rect 5330 32418 5364 32448
rect 5364 32418 5378 32448
rect 5392 32418 5444 32470
rect 4666 32353 4718 32405
rect 4732 32353 4784 32405
rect 4798 32353 4850 32405
rect 4864 32353 4916 32405
rect 4930 32353 4982 32405
rect 4996 32353 5048 32405
rect 5062 32353 5114 32405
rect 5128 32353 5180 32405
rect 5194 32353 5246 32405
rect 5260 32353 5312 32405
rect 5326 32375 5378 32405
rect 5326 32353 5330 32375
rect 5330 32353 5364 32375
rect 5364 32353 5378 32375
rect 5392 32353 5444 32405
rect 4666 32288 4718 32340
rect 4732 32288 4784 32340
rect 4798 32288 4850 32340
rect 4864 32288 4916 32340
rect 4930 32288 4982 32340
rect 4996 32288 5048 32340
rect 5062 32288 5114 32340
rect 5128 32288 5180 32340
rect 5194 32288 5246 32340
rect 5260 32288 5312 32340
rect 5326 32302 5378 32340
rect 5326 32288 5330 32302
rect 5330 32288 5364 32302
rect 5364 32288 5378 32302
rect 5392 32288 5444 32340
rect 4666 32223 4718 32275
rect 4732 32223 4784 32275
rect 4798 32223 4850 32275
rect 4864 32223 4916 32275
rect 4930 32223 4982 32275
rect 4996 32223 5048 32275
rect 5062 32223 5114 32275
rect 5128 32223 5180 32275
rect 5194 32223 5246 32275
rect 5260 32223 5312 32275
rect 5326 32268 5330 32275
rect 5330 32268 5364 32275
rect 5364 32268 5378 32275
rect 5326 32229 5378 32268
rect 5326 32223 5330 32229
rect 5330 32223 5364 32229
rect 5364 32223 5378 32229
rect 5392 32223 5444 32275
rect 4666 32158 4718 32210
rect 4732 32158 4784 32210
rect 4798 32158 4850 32210
rect 4864 32158 4916 32210
rect 4930 32158 4982 32210
rect 4996 32158 5048 32210
rect 5062 32158 5114 32210
rect 5128 32158 5180 32210
rect 5194 32158 5246 32210
rect 5260 32158 5312 32210
rect 5326 32195 5330 32210
rect 5330 32195 5364 32210
rect 5364 32195 5378 32210
rect 5326 32158 5378 32195
rect 5392 32158 5444 32210
rect 4666 32093 4718 32145
rect 4732 32093 4784 32145
rect 4798 32093 4850 32145
rect 4864 32093 4916 32145
rect 4930 32093 4982 32145
rect 4996 32093 5048 32145
rect 5062 32093 5114 32145
rect 5128 32093 5180 32145
rect 5194 32093 5246 32145
rect 5260 32093 5312 32145
rect 5326 32122 5330 32145
rect 5330 32122 5364 32145
rect 5364 32122 5378 32145
rect 5326 32093 5378 32122
rect 5392 32093 5444 32145
rect 4666 32028 4718 32080
rect 4732 32028 4784 32080
rect 4798 32028 4850 32080
rect 4864 32028 4916 32080
rect 4930 32028 4982 32080
rect 4996 32028 5048 32080
rect 5062 32028 5114 32080
rect 5128 32028 5180 32080
rect 5194 32028 5246 32080
rect 5260 32028 5312 32080
rect 5326 32049 5330 32080
rect 5330 32049 5364 32080
rect 5364 32049 5378 32080
rect 5326 32028 5378 32049
rect 5392 32028 5444 32080
rect 4666 31963 4718 32015
rect 4732 31963 4784 32015
rect 4798 31963 4850 32015
rect 4864 31963 4916 32015
rect 4930 31963 4982 32015
rect 4996 31963 5048 32015
rect 5062 31963 5114 32015
rect 5128 31963 5180 32015
rect 5194 31963 5246 32015
rect 5260 31963 5312 32015
rect 5326 32010 5378 32015
rect 5326 31976 5330 32010
rect 5330 31976 5364 32010
rect 5364 31976 5378 32010
rect 5326 31963 5378 31976
rect 5392 31963 5444 32015
rect 4666 31898 4718 31950
rect 4732 31898 4784 31950
rect 4798 31898 4850 31950
rect 4864 31898 4916 31950
rect 4930 31898 4982 31950
rect 4996 31898 5048 31950
rect 5062 31898 5114 31950
rect 5128 31898 5180 31950
rect 5194 31898 5246 31950
rect 5260 31898 5312 31950
rect 5326 31937 5378 31950
rect 5326 31903 5330 31937
rect 5330 31903 5364 31937
rect 5364 31903 5378 31937
rect 5326 31898 5378 31903
rect 5392 31898 5444 31950
rect 4666 31833 4718 31885
rect 4732 31833 4784 31885
rect 4798 31833 4850 31885
rect 4864 31833 4916 31885
rect 4930 31833 4982 31885
rect 4996 31833 5048 31885
rect 5062 31833 5114 31885
rect 5128 31833 5180 31885
rect 5194 31833 5246 31885
rect 5260 31833 5312 31885
rect 5326 31864 5378 31885
rect 5326 31833 5330 31864
rect 5330 31833 5364 31864
rect 5364 31833 5378 31864
rect 5392 31833 5444 31885
rect 4666 31768 4718 31820
rect 4732 31768 4784 31820
rect 4798 31768 4850 31820
rect 4864 31768 4916 31820
rect 4930 31768 4982 31820
rect 4996 31768 5048 31820
rect 5062 31768 5114 31820
rect 5128 31768 5180 31820
rect 5194 31768 5246 31820
rect 5260 31768 5312 31820
rect 5326 31791 5378 31820
rect 5326 31768 5330 31791
rect 5330 31768 5364 31791
rect 5364 31768 5378 31791
rect 5392 31768 5444 31820
rect 4666 31703 4718 31755
rect 4732 31703 4784 31755
rect 4798 31703 4850 31755
rect 4864 31703 4916 31755
rect 4930 31703 4982 31755
rect 4996 31703 5048 31755
rect 5062 31703 5114 31755
rect 5128 31703 5180 31755
rect 5194 31703 5246 31755
rect 5260 31703 5312 31755
rect 5326 31718 5378 31755
rect 5326 31703 5330 31718
rect 5330 31703 5364 31718
rect 5364 31703 5378 31718
rect 5392 31703 5444 31755
rect 4666 31638 4718 31690
rect 4732 31638 4784 31690
rect 4798 31638 4850 31690
rect 4864 31638 4916 31690
rect 4930 31638 4982 31690
rect 4996 31638 5048 31690
rect 5062 31638 5114 31690
rect 5128 31638 5180 31690
rect 5194 31638 5246 31690
rect 5260 31638 5312 31690
rect 5326 31684 5330 31690
rect 5330 31684 5364 31690
rect 5364 31684 5378 31690
rect 5326 31645 5378 31684
rect 5326 31638 5330 31645
rect 5330 31638 5364 31645
rect 5364 31638 5378 31645
rect 5392 31638 5444 31690
rect 4666 31573 4718 31625
rect 4732 31573 4784 31625
rect 4798 31573 4850 31625
rect 4864 31573 4916 31625
rect 4930 31573 4982 31625
rect 4996 31573 5048 31625
rect 5062 31573 5114 31625
rect 5128 31573 5180 31625
rect 5194 31573 5246 31625
rect 5260 31573 5312 31625
rect 5326 31611 5330 31625
rect 5330 31611 5364 31625
rect 5364 31611 5378 31625
rect 5326 31573 5378 31611
rect 5392 31573 5444 31625
rect 4666 31508 4718 31560
rect 4732 31508 4784 31560
rect 4798 31508 4850 31560
rect 4864 31508 4916 31560
rect 4930 31508 4982 31560
rect 4996 31508 5048 31560
rect 5062 31508 5114 31560
rect 5128 31508 5180 31560
rect 5194 31508 5246 31560
rect 5260 31508 5312 31560
rect 5326 31538 5330 31560
rect 5330 31538 5364 31560
rect 5364 31538 5378 31560
rect 5326 31508 5378 31538
rect 5392 31508 5444 31560
rect 4666 31443 4718 31495
rect 4732 31443 4784 31495
rect 4798 31443 4850 31495
rect 4864 31443 4916 31495
rect 4930 31443 4982 31495
rect 4996 31443 5048 31495
rect 5062 31443 5114 31495
rect 5128 31443 5180 31495
rect 5194 31443 5246 31495
rect 5260 31443 5312 31495
rect 5326 31465 5330 31495
rect 5330 31465 5364 31495
rect 5364 31465 5378 31495
rect 5326 31443 5378 31465
rect 5392 31443 5444 31495
rect 4666 31378 4718 31430
rect 4732 31378 4784 31430
rect 4798 31378 4850 31430
rect 4864 31378 4916 31430
rect 4930 31378 4982 31430
rect 4996 31378 5048 31430
rect 5062 31378 5114 31430
rect 5128 31378 5180 31430
rect 5194 31378 5246 31430
rect 5260 31378 5312 31430
rect 5326 31426 5378 31430
rect 5326 31392 5330 31426
rect 5330 31392 5364 31426
rect 5364 31392 5378 31426
rect 5326 31378 5378 31392
rect 5392 31378 5444 31430
rect 4666 31313 4718 31365
rect 4732 31313 4784 31365
rect 4798 31313 4850 31365
rect 4864 31313 4916 31365
rect 4930 31313 4982 31365
rect 4996 31313 5048 31365
rect 5062 31313 5114 31365
rect 5128 31313 5180 31365
rect 5194 31313 5246 31365
rect 5260 31313 5312 31365
rect 5326 31353 5378 31365
rect 5326 31319 5330 31353
rect 5330 31319 5364 31353
rect 5364 31319 5378 31353
rect 5326 31313 5378 31319
rect 5392 31313 5444 31365
rect 4666 31248 4718 31300
rect 4732 31248 4784 31300
rect 4798 31248 4850 31300
rect 4864 31248 4916 31300
rect 4930 31248 4982 31300
rect 4996 31248 5048 31300
rect 5062 31248 5114 31300
rect 5128 31248 5180 31300
rect 5194 31248 5246 31300
rect 5260 31248 5312 31300
rect 5326 31280 5378 31300
rect 5326 31248 5330 31280
rect 5330 31248 5364 31280
rect 5364 31248 5378 31280
rect 5392 31248 5444 31300
rect 4666 31183 4718 31235
rect 4732 31183 4784 31235
rect 4798 31183 4850 31235
rect 4864 31183 4916 31235
rect 4930 31183 4982 31235
rect 4996 31183 5048 31235
rect 5062 31183 5114 31235
rect 5128 31183 5180 31235
rect 5194 31183 5246 31235
rect 5260 31183 5312 31235
rect 5326 31207 5378 31235
rect 5326 31183 5330 31207
rect 5330 31183 5364 31207
rect 5364 31183 5378 31207
rect 5392 31183 5444 31235
rect 4666 31118 4718 31170
rect 4732 31118 4784 31170
rect 4798 31118 4850 31170
rect 4864 31118 4916 31170
rect 4930 31118 4982 31170
rect 4996 31118 5048 31170
rect 5062 31118 5114 31170
rect 5128 31118 5180 31170
rect 5194 31118 5246 31170
rect 5260 31118 5312 31170
rect 5326 31134 5378 31170
rect 5326 31118 5330 31134
rect 5330 31118 5364 31134
rect 5364 31118 5378 31134
rect 5392 31118 5444 31170
rect 4666 31053 4718 31105
rect 4732 31053 4784 31105
rect 4798 31053 4850 31105
rect 4864 31053 4916 31105
rect 4930 31053 4982 31105
rect 4996 31053 5048 31105
rect 5062 31053 5114 31105
rect 5128 31053 5180 31105
rect 5194 31053 5246 31105
rect 5260 31053 5312 31105
rect 5326 31100 5330 31105
rect 5330 31100 5364 31105
rect 5364 31100 5378 31105
rect 5326 31061 5378 31100
rect 5326 31053 5330 31061
rect 5330 31053 5364 31061
rect 5364 31053 5378 31061
rect 5392 31053 5444 31105
rect 4666 30988 4718 31040
rect 4732 30988 4784 31040
rect 4798 30988 4850 31040
rect 4864 30988 4916 31040
rect 4930 30988 4982 31040
rect 4996 30988 5048 31040
rect 5062 30988 5114 31040
rect 5128 30988 5180 31040
rect 5194 30988 5246 31040
rect 5260 30988 5312 31040
rect 5326 31027 5330 31040
rect 5330 31027 5364 31040
rect 5364 31027 5378 31040
rect 5326 30988 5378 31027
rect 5392 30988 5444 31040
rect 4666 30923 4718 30975
rect 4732 30923 4784 30975
rect 4798 30923 4850 30975
rect 4864 30923 4916 30975
rect 4930 30923 4982 30975
rect 4996 30923 5048 30975
rect 5062 30923 5114 30975
rect 5128 30923 5180 30975
rect 5194 30923 5246 30975
rect 5260 30923 5312 30975
rect 5326 30954 5330 30975
rect 5330 30954 5364 30975
rect 5364 30954 5378 30975
rect 5326 30923 5378 30954
rect 5392 30923 5444 30975
rect 4666 30858 4718 30910
rect 4732 30858 4784 30910
rect 4798 30858 4850 30910
rect 4864 30858 4916 30910
rect 4930 30858 4982 30910
rect 4996 30858 5048 30910
rect 5062 30858 5114 30910
rect 5128 30858 5180 30910
rect 5194 30858 5246 30910
rect 5260 30858 5312 30910
rect 5326 30881 5330 30910
rect 5330 30881 5364 30910
rect 5364 30881 5378 30910
rect 5326 30858 5378 30881
rect 5392 30858 5444 30910
rect 4666 30793 4718 30845
rect 4732 30793 4784 30845
rect 4798 30793 4850 30845
rect 4864 30793 4916 30845
rect 4930 30793 4982 30845
rect 4996 30793 5048 30845
rect 5062 30793 5114 30845
rect 5128 30793 5180 30845
rect 5194 30793 5246 30845
rect 5260 30793 5312 30845
rect 5326 30842 5378 30845
rect 5326 30808 5330 30842
rect 5330 30808 5364 30842
rect 5364 30808 5378 30842
rect 5326 30793 5378 30808
rect 5392 30793 5444 30845
rect 4666 30728 4718 30780
rect 4732 30728 4784 30780
rect 4798 30728 4850 30780
rect 4864 30728 4916 30780
rect 4930 30728 4982 30780
rect 4996 30728 5048 30780
rect 5062 30728 5114 30780
rect 5128 30728 5180 30780
rect 5194 30728 5246 30780
rect 5260 30728 5312 30780
rect 5326 30769 5378 30780
rect 5326 30735 5330 30769
rect 5330 30735 5364 30769
rect 5364 30735 5378 30769
rect 5326 30728 5378 30735
rect 5392 30728 5444 30780
rect 4666 30663 4718 30715
rect 4732 30663 4784 30715
rect 4798 30663 4850 30715
rect 4864 30663 4916 30715
rect 4930 30663 4982 30715
rect 4996 30663 5048 30715
rect 5062 30663 5114 30715
rect 5128 30663 5180 30715
rect 5194 30663 5246 30715
rect 5260 30663 5312 30715
rect 5326 30696 5378 30715
rect 5326 30663 5330 30696
rect 5330 30663 5364 30696
rect 5364 30663 5378 30696
rect 5392 30663 5444 30715
rect 4666 30598 4718 30650
rect 4732 30598 4784 30650
rect 4798 30598 4850 30650
rect 4864 30598 4916 30650
rect 4930 30598 4982 30650
rect 4996 30598 5048 30650
rect 5062 30598 5114 30650
rect 5128 30598 5180 30650
rect 5194 30598 5246 30650
rect 5260 30598 5312 30650
rect 5326 30623 5378 30650
rect 5326 30598 5330 30623
rect 5330 30598 5364 30623
rect 5364 30598 5378 30623
rect 5392 30598 5444 30650
rect 4666 30533 4718 30585
rect 4732 30533 4784 30585
rect 4798 30533 4850 30585
rect 4864 30533 4916 30585
rect 4930 30533 4982 30585
rect 4996 30533 5048 30585
rect 5062 30533 5114 30585
rect 5128 30533 5180 30585
rect 5194 30533 5246 30585
rect 5260 30533 5312 30585
rect 5326 30550 5378 30585
rect 5326 30533 5330 30550
rect 5330 30533 5364 30550
rect 5364 30533 5378 30550
rect 5392 30533 5444 30585
rect 4666 30468 4718 30520
rect 4732 30468 4784 30520
rect 4798 30468 4850 30520
rect 4864 30468 4916 30520
rect 4930 30468 4982 30520
rect 4996 30468 5048 30520
rect 5062 30468 5114 30520
rect 5128 30468 5180 30520
rect 5194 30468 5246 30520
rect 5260 30468 5312 30520
rect 5326 30516 5330 30520
rect 5330 30516 5364 30520
rect 5364 30516 5378 30520
rect 5326 30477 5378 30516
rect 5326 30468 5330 30477
rect 5330 30468 5364 30477
rect 5364 30468 5378 30477
rect 5392 30468 5444 30520
rect 4666 30403 4718 30455
rect 4732 30403 4784 30455
rect 4798 30403 4850 30455
rect 4864 30403 4916 30455
rect 4930 30403 4982 30455
rect 4996 30403 5048 30455
rect 5062 30403 5114 30455
rect 5128 30403 5180 30455
rect 5194 30403 5246 30455
rect 5260 30403 5312 30455
rect 5326 30443 5330 30455
rect 5330 30443 5364 30455
rect 5364 30443 5378 30455
rect 5326 30404 5378 30443
rect 5326 30403 5330 30404
rect 5330 30403 5364 30404
rect 5364 30403 5378 30404
rect 5392 30403 5444 30455
rect 4666 30338 4718 30390
rect 4732 30338 4784 30390
rect 4798 30338 4850 30390
rect 4864 30338 4916 30390
rect 4930 30338 4982 30390
rect 4996 30338 5048 30390
rect 5062 30338 5114 30390
rect 5128 30338 5180 30390
rect 5194 30338 5246 30390
rect 5260 30338 5312 30390
rect 5326 30370 5330 30390
rect 5330 30370 5364 30390
rect 5364 30370 5378 30390
rect 5326 30338 5378 30370
rect 5392 30338 5444 30390
rect 4869 30125 4921 30134
rect 4946 30125 4998 30134
rect 4869 30091 4889 30125
rect 4889 30091 4921 30125
rect 4946 30091 4964 30125
rect 4964 30091 4998 30125
rect 4869 30082 4921 30091
rect 4946 30082 4998 30091
rect 5022 30125 5074 30134
rect 5022 30091 5038 30125
rect 5038 30091 5072 30125
rect 5072 30091 5074 30125
rect 5022 30082 5074 30091
rect 5098 30125 5150 30134
rect 5098 30091 5112 30125
rect 5112 30091 5146 30125
rect 5146 30091 5150 30125
rect 5098 30082 5150 30091
rect 5174 30125 5226 30134
rect 5174 30091 5186 30125
rect 5186 30091 5220 30125
rect 5220 30091 5226 30125
rect 5174 30082 5226 30091
rect 6188 30047 6240 30099
rect 6188 29983 6240 30035
rect 6354 30002 6406 30054
rect 6418 30002 6470 30054
rect 3550 29853 3602 29905
rect 3550 29789 3602 29841
rect 5261 29853 5313 29905
rect 5261 29789 5313 29841
rect 6489 29922 6541 29974
rect 6553 29922 6605 29974
rect 3550 29429 3602 29481
rect 3550 29365 3602 29417
rect 5261 29429 5313 29481
rect 5261 29365 5313 29417
rect 4207 29139 4259 29147
rect 4271 29139 4323 29147
rect 4207 29105 4211 29139
rect 4211 29105 4254 29139
rect 4254 29105 4259 29139
rect 4271 29105 4288 29139
rect 4288 29105 4323 29139
rect 4207 29095 4259 29105
rect 4271 29095 4323 29105
rect 4744 29139 4796 29147
rect 4744 29105 4774 29139
rect 4774 29105 4796 29139
rect 4744 29095 4796 29105
rect 4808 29139 4860 29147
rect 4808 29105 4815 29139
rect 4815 29105 4849 29139
rect 4849 29105 4860 29139
rect 4808 29095 4860 29105
rect 4380 28957 4432 29009
rect 4444 28957 4496 29009
rect 3550 28869 3602 28921
rect 3550 28805 3602 28857
rect 5261 28869 5313 28921
rect 5261 28805 5313 28857
rect 4669 28434 4721 28443
rect 4736 28434 4788 28443
rect 4803 28434 4855 28443
rect 4870 28434 4922 28443
rect 4937 28434 4989 28443
rect 5004 28434 5056 28443
rect 5071 28434 5123 28443
rect 5138 28434 5190 28443
rect 5205 28434 5257 28443
rect 4669 28400 4691 28434
rect 4691 28400 4721 28434
rect 4736 28400 4764 28434
rect 4764 28400 4788 28434
rect 4803 28400 4837 28434
rect 4837 28400 4855 28434
rect 4870 28400 4871 28434
rect 4871 28400 4910 28434
rect 4910 28400 4922 28434
rect 4937 28400 4944 28434
rect 4944 28400 4983 28434
rect 4983 28400 4989 28434
rect 5004 28400 5017 28434
rect 5017 28400 5056 28434
rect 5071 28400 5090 28434
rect 5090 28400 5123 28434
rect 5138 28400 5163 28434
rect 5163 28400 5190 28434
rect 5205 28400 5236 28434
rect 5236 28400 5257 28434
rect 4669 28391 4721 28400
rect 4736 28391 4788 28400
rect 4803 28391 4855 28400
rect 4870 28391 4922 28400
rect 4937 28391 4989 28400
rect 5004 28391 5056 28400
rect 5071 28391 5123 28400
rect 5138 28391 5190 28400
rect 5205 28391 5257 28400
rect 5272 28434 5324 28443
rect 5272 28400 5275 28434
rect 5275 28400 5309 28434
rect 5309 28400 5324 28434
rect 5272 28391 5324 28400
rect 5339 28434 5391 28443
rect 5339 28400 5348 28434
rect 5348 28400 5382 28434
rect 5382 28400 5391 28434
rect 5339 28391 5391 28400
rect 5406 28434 5458 28443
rect 5406 28400 5421 28434
rect 5421 28400 5455 28434
rect 5455 28400 5458 28434
rect 5406 28391 5458 28400
rect 5473 28434 5525 28443
rect 5539 28434 5591 28443
rect 5473 28400 5494 28434
rect 5494 28400 5525 28434
rect 5539 28400 5567 28434
rect 5567 28400 5591 28434
rect 5473 28391 5525 28400
rect 5539 28391 5591 28400
rect 5605 28391 5657 28443
rect 3709 28174 3761 28183
rect 3776 28174 3828 28183
rect 3709 28140 3731 28174
rect 3731 28140 3761 28174
rect 3776 28140 3804 28174
rect 3804 28140 3828 28174
rect 3709 28131 3761 28140
rect 3776 28131 3828 28140
rect 3843 28174 3895 28183
rect 3843 28140 3877 28174
rect 3877 28140 3895 28174
rect 3843 28131 3895 28140
rect 3910 28174 3962 28183
rect 3910 28140 3916 28174
rect 3916 28140 3950 28174
rect 3950 28140 3962 28174
rect 3910 28131 3962 28140
rect 3977 28174 4029 28183
rect 3977 28140 3989 28174
rect 3989 28140 4023 28174
rect 4023 28140 4029 28174
rect 3977 28131 4029 28140
rect 4044 28174 4096 28183
rect 4044 28140 4062 28174
rect 4062 28140 4096 28174
rect 4044 28131 4096 28140
rect 4111 28174 4163 28183
rect 4178 28174 4230 28183
rect 4245 28174 4297 28183
rect 4312 28174 4364 28183
rect 4379 28174 4431 28183
rect 4445 28174 4497 28183
rect 4111 28140 4135 28174
rect 4135 28140 4163 28174
rect 4178 28140 4208 28174
rect 4208 28140 4230 28174
rect 4245 28140 4281 28174
rect 4281 28140 4297 28174
rect 4312 28140 4315 28174
rect 4315 28140 4354 28174
rect 4354 28140 4364 28174
rect 4379 28140 4388 28174
rect 4388 28140 4427 28174
rect 4427 28140 4431 28174
rect 4445 28140 4461 28174
rect 4461 28140 4497 28174
rect 4111 28131 4163 28140
rect 4178 28131 4230 28140
rect 4245 28131 4297 28140
rect 4312 28131 4364 28140
rect 4379 28131 4431 28140
rect 4445 28131 4497 28140
rect 8229 30469 8281 30521
rect 8293 30469 8345 30521
rect 4441 26156 4493 26208
rect 4508 26156 4560 26208
rect 4575 26156 4627 26208
rect 4642 26156 4694 26208
rect 4709 26156 4761 26208
rect 4776 26156 4828 26208
rect 4843 26156 4895 26208
rect 4910 26156 4962 26208
rect 4977 26199 5029 26208
rect 4977 26165 4980 26199
rect 4980 26165 5014 26199
rect 5014 26165 5029 26199
rect 4977 26156 5029 26165
rect 5044 26199 5096 26208
rect 5044 26165 5059 26199
rect 5059 26165 5093 26199
rect 5093 26165 5096 26199
rect 5044 26156 5096 26165
rect 2826 25506 2878 25531
rect 2826 25479 2832 25506
rect 2832 25479 2866 25506
rect 2866 25479 2878 25506
rect 2890 25506 2942 25531
rect 2890 25479 2904 25506
rect 2904 25479 2938 25506
rect 2938 25479 2942 25506
rect 3530 25507 3582 25559
rect 3596 25507 3648 25559
rect 2633 21640 2685 21692
rect 2730 21640 2782 21692
rect 2633 21564 2685 21616
rect 2730 21564 2782 21616
rect 2633 19654 2685 19706
rect 2730 19654 2782 19706
rect 2633 19578 2685 19630
rect 2730 19578 2782 19630
rect 2633 18694 2685 18746
rect 2730 18694 2782 18746
rect 2996 22133 3048 22185
rect 2996 22069 3048 22121
rect 3776 25506 3828 25558
rect 3844 25506 3896 25558
rect 3912 25506 3964 25558
rect 4500 25779 4552 25807
rect 4500 25755 4509 25779
rect 4509 25755 4543 25779
rect 4543 25755 4552 25779
rect 4500 25706 4552 25743
rect 4500 25691 4509 25706
rect 4509 25691 4543 25706
rect 4543 25691 4552 25706
rect 3999 25436 4051 25445
rect 3999 25402 4008 25436
rect 4008 25402 4042 25436
rect 4042 25402 4051 25436
rect 3999 25393 4051 25402
rect 3999 25360 4051 25367
rect 3999 25326 4008 25360
rect 4008 25326 4042 25360
rect 4042 25326 4051 25360
rect 3999 25315 4051 25326
rect 3999 25284 4051 25288
rect 3999 25250 4008 25284
rect 4008 25250 4042 25284
rect 4042 25250 4051 25284
rect 3999 25236 4051 25250
rect 3999 25208 4051 25209
rect 3999 25174 4008 25208
rect 4008 25174 4042 25208
rect 4042 25174 4051 25208
rect 3999 25157 4051 25174
rect 4344 25413 4396 25445
rect 4344 25393 4353 25413
rect 4353 25393 4387 25413
rect 4387 25393 4396 25413
rect 4344 25339 4396 25367
rect 4344 25315 4353 25339
rect 4353 25315 4387 25339
rect 4387 25315 4396 25339
rect 4344 25265 4396 25288
rect 4344 25236 4353 25265
rect 4353 25236 4387 25265
rect 4387 25236 4396 25265
rect 4344 25191 4396 25209
rect 4344 25157 4353 25191
rect 4353 25157 4387 25191
rect 4387 25157 4396 25191
rect 4812 25779 4864 25807
rect 4812 25755 4821 25779
rect 4821 25755 4855 25779
rect 4855 25755 4864 25779
rect 4812 25706 4864 25743
rect 4812 25691 4821 25706
rect 4821 25691 4855 25706
rect 4855 25691 4864 25706
rect 4656 25413 4708 25445
rect 4656 25393 4665 25413
rect 4665 25393 4699 25413
rect 4699 25393 4708 25413
rect 4656 25339 4708 25367
rect 4656 25315 4665 25339
rect 4665 25315 4699 25339
rect 4699 25315 4708 25339
rect 4656 25265 4708 25288
rect 4656 25236 4665 25265
rect 4665 25236 4699 25265
rect 4699 25236 4708 25265
rect 4656 25191 4708 25209
rect 4656 25157 4665 25191
rect 4665 25157 4699 25191
rect 4699 25157 4708 25191
rect 5124 25779 5176 25807
rect 5124 25755 5133 25779
rect 5133 25755 5167 25779
rect 5167 25755 5176 25779
rect 5124 25706 5176 25743
rect 5124 25691 5133 25706
rect 5133 25691 5167 25706
rect 5167 25691 5176 25706
rect 4968 25413 5020 25445
rect 4968 25393 4977 25413
rect 4977 25393 5011 25413
rect 5011 25393 5020 25413
rect 4968 25339 5020 25367
rect 4968 25315 4977 25339
rect 4977 25315 5011 25339
rect 5011 25315 5020 25339
rect 4968 25265 5020 25288
rect 4968 25236 4977 25265
rect 4977 25236 5011 25265
rect 5011 25236 5020 25265
rect 4968 25191 5020 25209
rect 4968 25157 4977 25191
rect 4977 25157 5011 25191
rect 5011 25157 5020 25191
rect 5436 25779 5488 25807
rect 5436 25755 5445 25779
rect 5445 25755 5479 25779
rect 5479 25755 5488 25779
rect 5436 25706 5488 25743
rect 5436 25691 5445 25706
rect 5445 25691 5479 25706
rect 5479 25691 5488 25706
rect 5280 25413 5332 25445
rect 5280 25393 5289 25413
rect 5289 25393 5323 25413
rect 5323 25393 5332 25413
rect 5280 25339 5332 25367
rect 5280 25315 5289 25339
rect 5289 25315 5323 25339
rect 5323 25315 5332 25339
rect 5280 25265 5332 25288
rect 5280 25236 5289 25265
rect 5289 25236 5323 25265
rect 5323 25236 5332 25265
rect 5280 25191 5332 25209
rect 5280 25157 5289 25191
rect 5289 25157 5323 25191
rect 5323 25157 5332 25191
rect 5592 25413 5644 25445
rect 5592 25393 5601 25413
rect 5601 25393 5635 25413
rect 5635 25393 5644 25413
rect 5592 25339 5644 25367
rect 5592 25315 5601 25339
rect 5601 25315 5635 25339
rect 5635 25315 5644 25339
rect 5592 25265 5644 25288
rect 5592 25236 5601 25265
rect 5601 25236 5635 25265
rect 5635 25236 5644 25265
rect 5592 25191 5644 25209
rect 5592 25157 5601 25191
rect 5601 25157 5635 25191
rect 5635 25157 5644 25191
rect 5937 25413 5989 25445
rect 5937 25393 5946 25413
rect 5946 25393 5980 25413
rect 5980 25393 5989 25413
rect 5937 25339 5989 25367
rect 5937 25315 5946 25339
rect 5946 25315 5980 25339
rect 5980 25315 5989 25339
rect 5937 25265 5989 25288
rect 5937 25236 5946 25265
rect 5946 25236 5980 25265
rect 5980 25236 5989 25265
rect 5937 25191 5989 25209
rect 5937 25157 5946 25191
rect 5946 25157 5980 25191
rect 5980 25157 5989 25191
rect 4451 23820 4503 23844
rect 4451 23792 4460 23820
rect 4460 23792 4494 23820
rect 4494 23792 4503 23820
rect 4451 23747 4503 23780
rect 4451 23728 4460 23747
rect 4460 23728 4494 23747
rect 4494 23728 4503 23747
rect 4646 23834 4698 23838
rect 4646 23800 4651 23834
rect 4651 23800 4685 23834
rect 4685 23800 4698 23834
rect 4646 23786 4698 23800
rect 4722 23834 4774 23838
rect 4722 23800 4731 23834
rect 4731 23800 4765 23834
rect 4765 23800 4774 23834
rect 4722 23786 4774 23800
rect 4797 23834 4849 23838
rect 4797 23800 4810 23834
rect 4810 23800 4844 23834
rect 4844 23800 4849 23834
rect 4797 23786 4849 23800
rect 4646 23762 4698 23774
rect 4646 23728 4651 23762
rect 4651 23728 4685 23762
rect 4685 23728 4698 23762
rect 4646 23722 4698 23728
rect 4722 23762 4774 23774
rect 4722 23728 4731 23762
rect 4731 23728 4765 23762
rect 4765 23728 4774 23762
rect 4722 23722 4774 23728
rect 4797 23762 4849 23774
rect 4797 23728 4810 23762
rect 4810 23728 4844 23762
rect 4844 23728 4849 23762
rect 4797 23722 4849 23728
rect 5055 23748 5060 23838
rect 5060 23748 5166 23838
rect 5166 23748 5171 23838
rect 5055 23722 5171 23748
rect 5310 23742 5315 23838
rect 5315 23742 5421 23838
rect 5421 23742 5426 23838
rect 5310 23722 5426 23742
rect 5849 23824 5901 23844
rect 5849 23792 5858 23824
rect 5858 23792 5892 23824
rect 5892 23792 5901 23824
rect 5849 23752 5901 23780
rect 5849 23728 5858 23752
rect 5858 23728 5892 23752
rect 5892 23728 5901 23752
rect 4879 22492 4931 22524
rect 4879 22472 4888 22492
rect 4888 22472 4922 22492
rect 4922 22472 4931 22492
rect 4879 22458 4888 22460
rect 4888 22458 4922 22460
rect 4922 22458 4931 22460
rect 4879 22419 4931 22458
rect 4879 22408 4888 22419
rect 4888 22408 4922 22419
rect 4922 22408 4931 22419
rect 4686 22106 4738 22115
rect 4750 22106 4802 22115
rect 4686 22072 4715 22106
rect 4715 22072 4738 22106
rect 4750 22072 4788 22106
rect 4788 22072 4802 22106
rect 4686 22063 4738 22072
rect 4750 22063 4802 22072
rect 3002 19764 3054 19816
rect 3066 19764 3118 19816
rect 5187 21666 5239 21686
rect 5187 21634 5196 21666
rect 5196 21634 5230 21666
rect 5230 21634 5239 21666
rect 5187 21593 5239 21622
rect 5187 21570 5196 21593
rect 5196 21570 5230 21593
rect 5230 21570 5239 21593
rect 4646 20445 4698 20449
rect 4646 20411 4676 20445
rect 4676 20411 4698 20445
rect 4646 20397 4698 20411
rect 4722 20445 4774 20449
rect 4722 20411 4726 20445
rect 4726 20411 4760 20445
rect 4760 20411 4774 20445
rect 4722 20397 4774 20411
rect 4797 20445 4849 20449
rect 4797 20411 4810 20445
rect 4810 20411 4844 20445
rect 4844 20411 4849 20445
rect 4797 20397 4849 20411
rect 4646 20373 4698 20385
rect 4646 20339 4676 20373
rect 4676 20339 4698 20373
rect 4646 20333 4698 20339
rect 4722 20373 4774 20385
rect 4722 20339 4726 20373
rect 4726 20339 4760 20373
rect 4760 20339 4774 20373
rect 4722 20333 4774 20339
rect 4797 20373 4849 20385
rect 4797 20339 4810 20373
rect 4810 20339 4844 20373
rect 4844 20339 4849 20373
rect 4797 20333 4849 20339
rect 4472 20028 4588 20054
rect 4472 19994 4494 20028
rect 4494 19994 4588 20028
rect 4472 19956 4588 19994
rect 4472 19938 4494 19956
rect 4494 19938 4588 19956
rect 4733 19971 4785 20023
rect 4797 19971 4849 20023
rect 4893 19857 4899 19886
rect 4899 19857 4933 19886
rect 4933 19857 4945 19886
rect 4893 19834 4945 19857
rect 4893 19818 4945 19822
rect 4893 19784 4899 19818
rect 4899 19784 4933 19818
rect 4933 19784 4945 19818
rect 5443 22508 5452 22524
rect 5452 22508 5486 22524
rect 5486 22508 5495 22524
rect 5443 22472 5495 22508
rect 5443 22435 5452 22460
rect 5452 22435 5486 22460
rect 5486 22435 5495 22460
rect 5443 22408 5495 22435
rect 7624 22285 7676 22337
rect 7688 22285 7740 22337
rect 7492 22205 7544 22257
rect 7556 22205 7608 22257
rect 7312 22125 7364 22177
rect 7376 22125 7428 22177
rect 5699 20201 5751 20253
rect 5699 20137 5751 20189
rect 4893 19770 4945 19784
rect 5461 19648 5513 19700
rect 5461 19584 5513 19636
rect 5080 19219 5132 19271
rect 5080 19155 5132 19207
rect 9567 30076 9619 30128
rect 9456 29996 9508 30048
rect 9300 29916 9352 29968
rect 9300 29852 9352 29904
rect 9230 22285 9282 22337
rect 9294 22285 9346 22337
rect 9456 29932 9508 29984
rect 9386 22205 9438 22257
rect 9450 22205 9502 22257
rect 9567 30012 9619 30064
rect 9567 22119 9619 22171
rect 9567 22055 9619 22107
rect 8223 20201 8275 20253
rect 8299 20201 8351 20253
rect 8223 20137 8275 20189
rect 8299 20137 8351 20189
rect 4987 18944 5039 18996
rect 4987 18880 5039 18932
rect 5247 18764 5299 18816
rect 5247 18700 5299 18752
rect 8799 19971 8851 20023
rect 8863 19971 8915 20023
rect 2996 18421 3048 18473
rect 2996 18357 3048 18409
rect 2633 17723 2685 17775
rect 2730 17723 2782 17775
rect 2633 17647 2685 17699
rect 2730 17647 2782 17699
rect 3709 18289 3761 18298
rect 3709 18255 3713 18289
rect 3713 18255 3761 18289
rect 3709 18246 3761 18255
rect 3776 18289 3828 18298
rect 3776 18255 3789 18289
rect 3789 18255 3823 18289
rect 3823 18255 3828 18289
rect 3776 18246 3828 18255
rect 3843 18289 3895 18298
rect 3843 18255 3861 18289
rect 3861 18255 3895 18289
rect 3843 18246 3895 18255
rect 3910 18289 3962 18298
rect 3977 18289 4029 18298
rect 4044 18289 4096 18298
rect 4111 18289 4163 18298
rect 4178 18289 4230 18298
rect 4245 18289 4297 18298
rect 4312 18289 4364 18298
rect 4379 18289 4431 18298
rect 4445 18289 4497 18298
rect 3910 18255 3933 18289
rect 3933 18255 3962 18289
rect 3977 18255 4005 18289
rect 4005 18255 4029 18289
rect 4044 18255 4077 18289
rect 4077 18255 4096 18289
rect 4111 18255 4149 18289
rect 4149 18255 4163 18289
rect 4178 18255 4183 18289
rect 4183 18255 4221 18289
rect 4221 18255 4230 18289
rect 4245 18255 4255 18289
rect 4255 18255 4293 18289
rect 4293 18255 4297 18289
rect 4312 18255 4327 18289
rect 4327 18255 4364 18289
rect 4379 18255 4399 18289
rect 4399 18255 4431 18289
rect 4445 18255 4471 18289
rect 4471 18255 4497 18289
rect 3910 18246 3962 18255
rect 3977 18246 4029 18255
rect 4044 18246 4096 18255
rect 4111 18246 4163 18255
rect 4178 18246 4230 18255
rect 4245 18246 4297 18255
rect 4312 18246 4364 18255
rect 4379 18246 4431 18255
rect 4445 18246 4497 18255
rect 2294 17567 2346 17619
rect 2391 17567 2443 17619
rect 2294 17491 2346 17543
rect 2391 17491 2443 17543
rect 1193 16824 1245 16876
rect 1257 16824 1309 16876
rect 1193 16368 1245 16420
rect 1257 16368 1309 16420
rect 2996 18150 3048 18202
rect 2996 18086 3048 18138
rect 2996 17401 3048 17453
rect 2996 17337 3048 17389
rect 2996 15954 3048 16006
rect 2996 15890 3048 15942
rect 3076 17923 3082 17925
rect 3082 17923 3116 17925
rect 3116 17923 3128 17925
rect 3076 17884 3128 17923
rect 3076 17873 3082 17884
rect 3082 17873 3116 17884
rect 3116 17873 3128 17884
rect 3076 17850 3082 17861
rect 3082 17850 3116 17861
rect 3116 17850 3128 17861
rect 3076 17811 3128 17850
rect 3076 17809 3082 17811
rect 3082 17809 3116 17811
rect 3116 17809 3128 17811
rect 3183 17879 3235 17931
rect 3254 17879 3306 17931
rect 3324 17879 3376 17931
rect 3183 17803 3235 17855
rect 3254 17803 3306 17855
rect 3324 17803 3376 17855
rect 3946 17873 3998 17925
rect 3946 17809 3998 17861
rect 3435 17603 3487 17613
rect 3435 17569 3444 17603
rect 3444 17569 3478 17603
rect 3478 17569 3487 17603
rect 3435 17561 3487 17569
rect 3435 17529 3487 17549
rect 3435 17497 3444 17529
rect 3444 17497 3478 17529
rect 3478 17497 3487 17529
rect 3540 17427 3592 17453
rect 3540 17401 3552 17427
rect 3552 17401 3586 17427
rect 3586 17401 3592 17427
rect 3540 17345 3592 17389
rect 3540 17337 3552 17345
rect 3552 17337 3586 17345
rect 3586 17337 3592 17345
rect 3620 17405 3672 17457
rect 3620 17341 3672 17393
rect 4215 17873 4267 17925
rect 4215 17809 4267 17861
rect 4371 17717 4423 17769
rect 4371 17653 4423 17705
rect 4527 17873 4579 17925
rect 4527 17809 4579 17861
rect 4682 17717 4734 17769
rect 4682 17653 4734 17705
rect 4839 17873 4891 17925
rect 4839 17809 4891 17861
rect 4995 17561 5047 17613
rect 4995 17497 5047 17549
rect 5151 17873 5203 17925
rect 5151 17809 5203 17861
rect 5307 17561 5359 17613
rect 5307 17497 5359 17549
rect 5462 17873 5514 17925
rect 5462 17809 5514 17861
rect 5832 17873 5884 17925
rect 5832 17809 5884 17861
rect 4383 16867 4435 16876
rect 4383 16833 4387 16867
rect 4387 16833 4421 16867
rect 4421 16833 4435 16867
rect 4383 16824 4435 16833
rect 4447 16867 4499 16876
rect 4447 16833 4460 16867
rect 4460 16833 4494 16867
rect 4494 16833 4499 16867
rect 4447 16824 4499 16833
rect 5056 16740 5108 16792
rect 5120 16740 5172 16792
rect 4180 16600 4232 16652
rect 4180 16536 4232 16588
rect 4884 16368 4936 16420
rect 4948 16368 5000 16420
rect 3234 15960 3286 16012
rect 3298 15960 3350 16012
rect 3076 15840 3128 15872
rect 3076 15820 3082 15840
rect 3082 15820 3116 15840
rect 3116 15820 3128 15840
rect 3076 15806 3082 15808
rect 3082 15806 3116 15808
rect 3116 15806 3128 15808
rect 3076 15767 3128 15806
rect 3076 15756 3082 15767
rect 3082 15756 3116 15767
rect 3116 15756 3128 15767
rect 6464 15843 6516 15872
rect 6464 15820 6476 15843
rect 6476 15820 6510 15843
rect 6510 15820 6516 15843
rect 6464 15770 6516 15808
rect 6464 15756 6476 15770
rect 6476 15756 6510 15770
rect 6510 15756 6516 15770
rect 5837 14809 5889 14861
rect 5837 14741 5889 14793
rect 5837 14673 5889 14725
rect 6211 14823 6263 14861
rect 6295 14823 6347 14861
rect 6211 14809 6237 14823
rect 6237 14809 6263 14823
rect 6295 14809 6309 14823
rect 6309 14809 6343 14823
rect 6343 14809 6347 14823
rect 6379 14809 6431 14861
rect 6463 14860 6476 14861
rect 6476 14860 6510 14861
rect 6510 14860 6515 14861
rect 6463 14821 6515 14860
rect 6463 14809 6476 14821
rect 6476 14809 6510 14821
rect 6510 14809 6515 14821
rect 6211 14789 6237 14793
rect 6237 14789 6263 14793
rect 6295 14789 6309 14793
rect 6309 14789 6343 14793
rect 6343 14789 6347 14793
rect 6211 14749 6263 14789
rect 6295 14749 6347 14789
rect 6211 14741 6237 14749
rect 6237 14741 6263 14749
rect 6295 14741 6309 14749
rect 6309 14741 6343 14749
rect 6343 14741 6347 14749
rect 6379 14741 6431 14793
rect 6463 14787 6476 14793
rect 6476 14787 6510 14793
rect 6510 14787 6515 14793
rect 6463 14748 6515 14787
rect 6463 14741 6476 14748
rect 6476 14741 6510 14748
rect 6510 14741 6515 14748
rect 6211 14715 6237 14725
rect 6237 14715 6263 14725
rect 6295 14715 6309 14725
rect 6309 14715 6343 14725
rect 6343 14715 6347 14725
rect 6211 14675 6263 14715
rect 6295 14675 6347 14715
rect 6211 14673 6237 14675
rect 6237 14673 6263 14675
rect 6295 14673 6343 14675
rect 6343 14673 6347 14675
rect 6379 14673 6431 14725
rect 6463 14714 6476 14725
rect 6476 14714 6510 14725
rect 6510 14714 6515 14725
rect 6463 14675 6515 14714
rect 6463 14673 6476 14675
rect 6476 14673 6510 14675
rect 6510 14673 6515 14675
rect 8799 17409 8851 17461
rect 8863 17409 8915 17461
<< metal2 >>
rect 4663 39195 5663 39276
rect 4663 39143 4666 39195
rect 4718 39143 4732 39195
rect 4784 39192 4798 39195
rect 4850 39192 4864 39195
rect 4916 39192 4930 39195
rect 4982 39192 4996 39195
rect 5048 39192 5062 39195
rect 5114 39192 5128 39195
rect 5180 39192 5194 39195
rect 5246 39192 5260 39195
rect 5312 39192 5326 39195
rect 5378 39192 5392 39195
rect 5444 39192 5663 39195
rect 4663 39131 4775 39143
rect 4663 39079 4666 39131
rect 4718 39079 4732 39131
rect 4663 39067 4775 39079
rect 4663 39015 4666 39067
rect 4718 39015 4732 39067
rect 4663 39003 4775 39015
rect 4663 38951 4666 39003
rect 4718 38951 4732 39003
rect 4663 38939 4775 38951
rect 4663 38887 4666 38939
rect 4718 38887 4732 38939
rect 4663 38875 4775 38887
rect 4663 38823 4666 38875
rect 4718 38823 4732 38875
rect 4663 38811 4775 38823
rect 4663 38759 4666 38811
rect 4718 38759 4732 38811
rect 4663 38747 4775 38759
rect 4663 38695 4666 38747
rect 4718 38695 4732 38747
rect 4663 38683 4775 38695
rect 4663 38631 4666 38683
rect 4718 38631 4732 38683
rect 4663 38619 4775 38631
rect 4663 38567 4666 38619
rect 4718 38567 4732 38619
rect 4663 38555 4775 38567
rect 4663 38503 4666 38555
rect 4718 38503 4732 38555
rect 4663 38491 4775 38503
rect 4663 38439 4666 38491
rect 4718 38439 4732 38491
rect 4663 38427 4775 38439
rect 4663 38375 4666 38427
rect 4718 38375 4732 38427
rect 4663 38363 4775 38375
rect 4663 38311 4666 38363
rect 4718 38311 4732 38363
rect 4663 38299 4775 38311
rect 4663 38247 4666 38299
rect 4718 38247 4732 38299
rect 4663 38235 4775 38247
rect 4663 38183 4666 38235
rect 4718 38183 4732 38235
rect 4663 38171 4775 38183
rect 4663 38119 4666 38171
rect 4718 38119 4732 38171
rect 4663 38107 4775 38119
rect 4663 38055 4666 38107
rect 4718 38055 4732 38107
rect 4663 38043 4775 38055
rect 4663 37991 4666 38043
rect 4718 37991 4732 38043
rect 4663 37979 4775 37991
rect 4663 37927 4666 37979
rect 4718 37927 4732 37979
rect 4663 37915 4775 37927
rect 4663 37863 4666 37915
rect 4718 37863 4732 37915
rect 4663 37851 4775 37863
rect 4663 37799 4666 37851
rect 4718 37799 4732 37851
rect 4663 37787 4775 37799
rect 4663 37735 4666 37787
rect 4718 37735 4732 37787
rect 4663 37723 4775 37735
rect 4663 37671 4666 37723
rect 4718 37671 4732 37723
rect 4663 37659 4775 37671
rect 4663 37607 4666 37659
rect 4718 37607 4732 37659
rect 4663 37595 4775 37607
rect 4663 37543 4666 37595
rect 4718 37543 4732 37595
rect 4663 37531 4775 37543
rect 4663 37479 4666 37531
rect 4718 37479 4732 37531
rect 4663 37467 4775 37479
rect 4663 37415 4666 37467
rect 4718 37415 4732 37467
rect 4663 37403 4775 37415
rect 4663 37351 4666 37403
rect 4718 37351 4732 37403
rect 4663 37339 4775 37351
rect 4663 37287 4666 37339
rect 4718 37287 4732 37339
rect 4663 37275 4775 37287
rect 4663 37223 4666 37275
rect 4718 37223 4732 37275
rect 4663 37211 4775 37223
rect 4663 37159 4666 37211
rect 4718 37159 4732 37211
rect 4663 37147 4775 37159
rect 4663 37095 4666 37147
rect 4718 37095 4732 37147
rect 4663 37083 4775 37095
rect 4663 37031 4666 37083
rect 4718 37031 4732 37083
rect 4663 37019 4775 37031
rect 4663 36967 4666 37019
rect 4718 36967 4732 37019
rect 4663 36955 4775 36967
rect 4663 36903 4666 36955
rect 4718 36903 4732 36955
rect 4663 36891 4775 36903
rect 4663 36839 4666 36891
rect 4718 36839 4732 36891
rect 4663 36827 4775 36839
rect 4663 36775 4666 36827
rect 4718 36775 4732 36827
rect 4663 36763 4775 36775
rect 4663 36711 4666 36763
rect 4718 36711 4732 36763
rect 4663 36699 4775 36711
rect 4663 36647 4666 36699
rect 4718 36647 4732 36699
rect 4663 36635 4775 36647
rect 4663 36583 4666 36635
rect 4718 36583 4732 36635
rect 4663 36571 4775 36583
rect 4663 36519 4666 36571
rect 4718 36519 4732 36571
rect 4663 36507 4775 36519
rect 4663 36455 4666 36507
rect 4718 36455 4732 36507
rect 4663 36443 4775 36455
rect 4663 36391 4666 36443
rect 4718 36391 4732 36443
rect 5551 36416 5663 39192
rect 4784 36391 4798 36416
rect 4850 36391 4864 36416
rect 4916 36391 4930 36416
rect 4982 36391 4996 36416
rect 5048 36391 5062 36416
rect 5114 36391 5128 36416
rect 5180 36391 5194 36416
rect 5246 36391 5260 36416
rect 5312 36391 5326 36416
rect 5378 36391 5392 36416
rect 5444 36391 5663 36416
rect 4663 36379 4775 36391
rect 4831 36379 4855 36391
rect 4911 36379 4935 36391
rect 4991 36379 5015 36391
rect 5071 36379 5095 36391
rect 5151 36379 5175 36391
rect 5231 36379 5255 36391
rect 5311 36379 5335 36391
rect 5391 36379 5415 36391
rect 4663 36327 4666 36379
rect 4718 36327 4732 36379
rect 4850 36335 4855 36379
rect 4784 36327 4798 36335
rect 4850 36327 4864 36335
rect 4916 36327 4930 36379
rect 4991 36335 4996 36379
rect 5246 36335 5255 36379
rect 4982 36327 4996 36335
rect 5048 36327 5062 36335
rect 5114 36327 5128 36335
rect 5180 36327 5194 36335
rect 5246 36327 5260 36335
rect 5312 36327 5326 36379
rect 5391 36335 5392 36379
rect 5471 36335 5495 36391
rect 5551 36335 5663 36391
rect 5378 36327 5392 36335
rect 5444 36327 5663 36335
rect 4663 36315 5663 36327
rect 4663 36263 4666 36315
rect 4718 36263 4732 36315
rect 4784 36310 4798 36315
rect 4850 36310 4864 36315
rect 4850 36263 4855 36310
rect 4916 36263 4930 36315
rect 4982 36310 4996 36315
rect 5048 36310 5062 36315
rect 5114 36310 5128 36315
rect 5180 36310 5194 36315
rect 5246 36310 5260 36315
rect 4991 36263 4996 36310
rect 5246 36263 5255 36310
rect 5312 36263 5326 36315
rect 5378 36310 5392 36315
rect 5444 36310 5663 36315
rect 5391 36263 5392 36310
rect 4663 36254 4775 36263
rect 4831 36254 4855 36263
rect 4911 36254 4935 36263
rect 4991 36254 5015 36263
rect 5071 36254 5095 36263
rect 5151 36254 5175 36263
rect 5231 36254 5255 36263
rect 5311 36254 5335 36263
rect 5391 36254 5415 36263
rect 5471 36254 5495 36310
rect 5551 36254 5663 36310
rect 4663 36251 5663 36254
rect 4663 36199 4666 36251
rect 4718 36199 4732 36251
rect 4784 36229 4798 36251
rect 4850 36229 4864 36251
rect 4850 36199 4855 36229
rect 4916 36199 4930 36251
rect 4982 36229 4996 36251
rect 5048 36229 5062 36251
rect 5114 36229 5128 36251
rect 5180 36229 5194 36251
rect 5246 36229 5260 36251
rect 4991 36199 4996 36229
rect 5246 36199 5255 36229
rect 5312 36199 5326 36251
rect 5378 36229 5392 36251
rect 5444 36229 5663 36251
rect 5391 36199 5392 36229
rect 4663 36187 4775 36199
rect 4831 36187 4855 36199
rect 4911 36187 4935 36199
rect 4991 36187 5015 36199
rect 5071 36187 5095 36199
rect 5151 36187 5175 36199
rect 5231 36187 5255 36199
rect 5311 36187 5335 36199
rect 5391 36187 5415 36199
rect 4663 36135 4666 36187
rect 4718 36135 4732 36187
rect 4850 36173 4855 36187
rect 4784 36148 4798 36173
rect 4850 36148 4864 36173
rect 4850 36135 4855 36148
rect 4916 36135 4930 36187
rect 4991 36173 4996 36187
rect 5246 36173 5255 36187
rect 4982 36148 4996 36173
rect 5048 36148 5062 36173
rect 5114 36148 5128 36173
rect 5180 36148 5194 36173
rect 5246 36148 5260 36173
rect 4991 36135 4996 36148
rect 5246 36135 5255 36148
rect 5312 36135 5326 36187
rect 5391 36173 5392 36187
rect 5471 36173 5495 36229
rect 5551 36173 5663 36229
rect 5378 36148 5392 36173
rect 5444 36148 5663 36173
rect 5391 36135 5392 36148
rect 4663 36123 4775 36135
rect 4831 36123 4855 36135
rect 4911 36123 4935 36135
rect 4991 36123 5015 36135
rect 5071 36123 5095 36135
rect 5151 36123 5175 36135
rect 5231 36123 5255 36135
rect 5311 36123 5335 36135
rect 5391 36123 5415 36135
rect 4663 36071 4666 36123
rect 4718 36071 4732 36123
rect 4850 36092 4855 36123
rect 4784 36071 4798 36092
rect 4850 36071 4864 36092
rect 4916 36071 4930 36123
rect 4991 36092 4996 36123
rect 5246 36092 5255 36123
rect 4982 36071 4996 36092
rect 5048 36071 5062 36092
rect 5114 36071 5128 36092
rect 5180 36071 5194 36092
rect 5246 36071 5260 36092
rect 5312 36071 5326 36123
rect 5391 36092 5392 36123
rect 5471 36092 5495 36148
rect 5551 36092 5663 36148
rect 5378 36071 5392 36092
rect 5444 36071 5663 36092
rect 4663 36067 5663 36071
rect 4663 36059 4775 36067
rect 4831 36059 4855 36067
rect 4911 36059 4935 36067
rect 4991 36059 5015 36067
rect 5071 36059 5095 36067
rect 5151 36059 5175 36067
rect 5231 36059 5255 36067
rect 5311 36059 5335 36067
rect 5391 36059 5415 36067
rect 4663 36007 4666 36059
rect 4718 36007 4732 36059
rect 4850 36011 4855 36059
rect 4784 36007 4798 36011
rect 4850 36007 4864 36011
rect 4916 36007 4930 36059
rect 4991 36011 4996 36059
rect 5246 36011 5255 36059
rect 4982 36007 4996 36011
rect 5048 36007 5062 36011
rect 5114 36007 5128 36011
rect 5180 36007 5194 36011
rect 5246 36007 5260 36011
rect 5312 36007 5326 36059
rect 5391 36011 5392 36059
rect 5471 36011 5495 36067
rect 5551 36011 5663 36067
rect 5378 36007 5392 36011
rect 5444 36007 5663 36011
rect 4663 35995 5663 36007
rect 4663 35943 4666 35995
rect 4718 35943 4732 35995
rect 4784 35986 4798 35995
rect 4850 35986 4864 35995
rect 4850 35943 4855 35986
rect 4916 35943 4930 35995
rect 4982 35986 4996 35995
rect 5048 35986 5062 35995
rect 5114 35986 5128 35995
rect 5180 35986 5194 35995
rect 5246 35986 5260 35995
rect 4991 35943 4996 35986
rect 5246 35943 5255 35986
rect 5312 35943 5326 35995
rect 5378 35986 5392 35995
rect 5444 35986 5663 35995
rect 5391 35943 5392 35986
rect 4663 35931 4775 35943
rect 4831 35931 4855 35943
rect 4911 35931 4935 35943
rect 4991 35931 5015 35943
rect 5071 35931 5095 35943
rect 5151 35931 5175 35943
rect 5231 35931 5255 35943
rect 5311 35931 5335 35943
rect 5391 35931 5415 35943
rect 4663 35879 4666 35931
rect 4718 35879 4732 35931
rect 4850 35930 4855 35931
rect 4784 35905 4798 35930
rect 4850 35905 4864 35930
rect 4850 35879 4855 35905
rect 4916 35879 4930 35931
rect 4991 35930 4996 35931
rect 5246 35930 5255 35931
rect 4982 35905 4996 35930
rect 5048 35905 5062 35930
rect 5114 35905 5128 35930
rect 5180 35905 5194 35930
rect 5246 35905 5260 35930
rect 4991 35879 4996 35905
rect 5246 35879 5255 35905
rect 5312 35879 5326 35931
rect 5391 35930 5392 35931
rect 5471 35930 5495 35986
rect 5551 35930 5663 35986
rect 5378 35905 5392 35930
rect 5444 35905 5663 35930
rect 5391 35879 5392 35905
rect 4663 35867 4775 35879
rect 4831 35867 4855 35879
rect 4911 35867 4935 35879
rect 4991 35867 5015 35879
rect 5071 35867 5095 35879
rect 5151 35867 5175 35879
rect 5231 35867 5255 35879
rect 5311 35867 5335 35879
rect 5391 35867 5415 35879
rect 4663 35815 4666 35867
rect 4718 35815 4732 35867
rect 4850 35849 4855 35867
rect 4784 35824 4798 35849
rect 4850 35824 4864 35849
rect 4850 35815 4855 35824
rect 4916 35815 4930 35867
rect 4991 35849 4996 35867
rect 5246 35849 5255 35867
rect 4982 35824 4996 35849
rect 5048 35824 5062 35849
rect 5114 35824 5128 35849
rect 5180 35824 5194 35849
rect 5246 35824 5260 35849
rect 4991 35815 4996 35824
rect 5246 35815 5255 35824
rect 5312 35815 5326 35867
rect 5391 35849 5392 35867
rect 5471 35849 5495 35905
rect 5551 35849 5663 35905
rect 5378 35824 5392 35849
rect 5444 35824 5663 35849
rect 5391 35815 5392 35824
rect 4663 35803 4775 35815
rect 4831 35803 4855 35815
rect 4911 35803 4935 35815
rect 4991 35803 5015 35815
rect 5071 35803 5095 35815
rect 5151 35803 5175 35815
rect 5231 35803 5255 35815
rect 5311 35803 5335 35815
rect 5391 35803 5415 35815
rect 4663 35751 4666 35803
rect 4718 35751 4732 35803
rect 4850 35768 4855 35803
rect 4784 35751 4798 35768
rect 4850 35751 4864 35768
rect 4916 35751 4930 35803
rect 4991 35768 4996 35803
rect 5246 35768 5255 35803
rect 4982 35751 4996 35768
rect 5048 35751 5062 35768
rect 5114 35751 5128 35768
rect 5180 35751 5194 35768
rect 5246 35751 5260 35768
rect 5312 35751 5326 35803
rect 5391 35768 5392 35803
rect 5471 35768 5495 35824
rect 5551 35768 5663 35824
rect 5378 35751 5392 35768
rect 5444 35751 5663 35768
rect 4663 35743 5663 35751
rect 4663 35739 4775 35743
rect 4831 35739 4855 35743
rect 4911 35739 4935 35743
rect 4991 35739 5015 35743
rect 5071 35739 5095 35743
rect 5151 35739 5175 35743
rect 5231 35739 5255 35743
rect 5311 35739 5335 35743
rect 5391 35739 5415 35743
rect 4663 35687 4666 35739
rect 4718 35687 4732 35739
rect 4850 35687 4855 35739
rect 4916 35687 4930 35739
rect 4991 35687 4996 35739
rect 5246 35687 5255 35739
rect 5312 35687 5326 35739
rect 5391 35687 5392 35739
rect 5471 35687 5495 35743
rect 5551 35687 5663 35743
rect 4663 35675 5663 35687
rect 1187 35643 3217 35649
rect 1187 35591 1211 35643
rect 1263 35591 3165 35643
rect 1187 35579 3217 35591
rect 1187 35527 1211 35579
rect 1263 35527 3165 35579
rect 1187 35521 3217 35527
rect 4663 35623 4666 35675
rect 4718 35623 4732 35675
rect 4784 35662 4798 35675
rect 4850 35662 4864 35675
rect 4850 35623 4855 35662
rect 4916 35623 4930 35675
rect 4982 35662 4996 35675
rect 5048 35662 5062 35675
rect 5114 35662 5128 35675
rect 5180 35662 5194 35675
rect 5246 35662 5260 35675
rect 4991 35623 4996 35662
rect 5246 35623 5255 35662
rect 5312 35623 5326 35675
rect 5378 35662 5392 35675
rect 5444 35662 5663 35675
rect 5391 35623 5392 35662
rect 4663 35611 4775 35623
rect 4831 35611 4855 35623
rect 4911 35611 4935 35623
rect 4991 35611 5015 35623
rect 5071 35611 5095 35623
rect 5151 35611 5175 35623
rect 5231 35611 5255 35623
rect 5311 35611 5335 35623
rect 5391 35611 5415 35623
rect 4663 35559 4666 35611
rect 4718 35559 4732 35611
rect 4850 35606 4855 35611
rect 4784 35581 4798 35606
rect 4850 35581 4864 35606
rect 4850 35559 4855 35581
rect 4916 35559 4930 35611
rect 4991 35606 4996 35611
rect 5246 35606 5255 35611
rect 4982 35581 4996 35606
rect 5048 35581 5062 35606
rect 5114 35581 5128 35606
rect 5180 35581 5194 35606
rect 5246 35581 5260 35606
rect 4991 35559 4996 35581
rect 5246 35559 5255 35581
rect 5312 35559 5326 35611
rect 5391 35606 5392 35611
rect 5471 35606 5495 35662
rect 5551 35606 5663 35662
rect 5378 35581 5392 35606
rect 5444 35581 5663 35606
rect 5391 35559 5392 35581
rect 4663 35547 4775 35559
rect 4831 35547 4855 35559
rect 4911 35547 4935 35559
rect 4991 35547 5015 35559
rect 5071 35547 5095 35559
rect 5151 35547 5175 35559
rect 5231 35547 5255 35559
rect 5311 35547 5335 35559
rect 5391 35547 5415 35559
rect 4663 35495 4666 35547
rect 4718 35495 4732 35547
rect 4850 35525 4855 35547
rect 4784 35500 4798 35525
rect 4850 35500 4864 35525
rect 4850 35495 4855 35500
rect 4916 35495 4930 35547
rect 4991 35525 4996 35547
rect 5246 35525 5255 35547
rect 4982 35500 4996 35525
rect 5048 35500 5062 35525
rect 5114 35500 5128 35525
rect 5180 35500 5194 35525
rect 5246 35500 5260 35525
rect 4991 35495 4996 35500
rect 5246 35495 5255 35500
rect 5312 35495 5326 35547
rect 5391 35525 5392 35547
rect 5471 35525 5495 35581
rect 5551 35525 5663 35581
rect 5378 35500 5392 35525
rect 5444 35500 5663 35525
rect 5391 35495 5392 35500
rect 4663 35483 4775 35495
rect 4831 35483 4855 35495
rect 4911 35483 4935 35495
rect 4991 35483 5015 35495
rect 5071 35483 5095 35495
rect 5151 35483 5175 35495
rect 5231 35483 5255 35495
rect 5311 35483 5335 35495
rect 5391 35483 5415 35495
rect 4663 35431 4666 35483
rect 4718 35431 4732 35483
rect 4850 35444 4855 35483
rect 4784 35431 4798 35444
rect 4850 35431 4864 35444
rect 4916 35431 4930 35483
rect 4991 35444 4996 35483
rect 5246 35444 5255 35483
rect 4982 35431 4996 35444
rect 5048 35431 5062 35444
rect 5114 35431 5128 35444
rect 5180 35431 5194 35444
rect 5246 35431 5260 35444
rect 5312 35431 5326 35483
rect 5391 35444 5392 35483
rect 5471 35444 5495 35500
rect 5551 35444 5663 35500
rect 5378 35431 5392 35444
rect 5444 35431 5663 35444
rect 4663 35419 5663 35431
rect 4663 35367 4666 35419
rect 4718 35367 4732 35419
rect 4850 35367 4855 35419
rect 4916 35367 4930 35419
rect 4991 35367 4996 35419
rect 5246 35367 5255 35419
rect 5312 35367 5326 35419
rect 5391 35367 5392 35419
rect 4663 35363 4775 35367
rect 4831 35363 4855 35367
rect 4911 35363 4935 35367
rect 4991 35363 5015 35367
rect 5071 35363 5095 35367
rect 5151 35363 5175 35367
rect 5231 35363 5255 35367
rect 5311 35363 5335 35367
rect 5391 35363 5415 35367
rect 5471 35363 5495 35419
rect 5551 35363 5663 35419
rect 4663 35355 5663 35363
rect 4663 35303 4666 35355
rect 4718 35303 4732 35355
rect 4784 35338 4798 35355
rect 4850 35338 4864 35355
rect 4850 35303 4855 35338
rect 4916 35303 4930 35355
rect 4982 35338 4996 35355
rect 5048 35338 5062 35355
rect 5114 35338 5128 35355
rect 5180 35338 5194 35355
rect 5246 35338 5260 35355
rect 4991 35303 4996 35338
rect 5246 35303 5255 35338
rect 5312 35303 5326 35355
rect 5378 35338 5392 35355
rect 5444 35338 5663 35355
rect 5391 35303 5392 35338
rect 4663 35291 4775 35303
rect 4831 35291 4855 35303
rect 4911 35291 4935 35303
rect 4991 35291 5015 35303
rect 5071 35291 5095 35303
rect 5151 35291 5175 35303
rect 5231 35291 5255 35303
rect 5311 35291 5335 35303
rect 5391 35291 5415 35303
rect 4663 35239 4666 35291
rect 4718 35239 4732 35291
rect 4850 35282 4855 35291
rect 4784 35257 4798 35282
rect 4850 35257 4864 35282
rect 4850 35239 4855 35257
rect 4916 35239 4930 35291
rect 4991 35282 4996 35291
rect 5246 35282 5255 35291
rect 4982 35257 4996 35282
rect 5048 35257 5062 35282
rect 5114 35257 5128 35282
rect 5180 35257 5194 35282
rect 5246 35257 5260 35282
rect 4991 35239 4996 35257
rect 5246 35239 5255 35257
rect 5312 35239 5326 35291
rect 5391 35282 5392 35291
rect 5471 35282 5495 35338
rect 5551 35282 5663 35338
rect 5378 35257 5392 35282
rect 5444 35257 5663 35282
rect 5391 35239 5392 35257
rect 4663 35227 4775 35239
rect 4831 35227 4855 35239
rect 4911 35227 4935 35239
rect 4991 35227 5015 35239
rect 5071 35227 5095 35239
rect 5151 35227 5175 35239
rect 5231 35227 5255 35239
rect 5311 35227 5335 35239
rect 5391 35227 5415 35239
rect 4663 35175 4666 35227
rect 4718 35175 4732 35227
rect 4850 35201 4855 35227
rect 4784 35176 4798 35201
rect 4850 35176 4864 35201
rect 4850 35175 4855 35176
rect 4916 35175 4930 35227
rect 4991 35201 4996 35227
rect 5246 35201 5255 35227
rect 4982 35176 4996 35201
rect 5048 35176 5062 35201
rect 5114 35176 5128 35201
rect 5180 35176 5194 35201
rect 5246 35176 5260 35201
rect 4991 35175 4996 35176
rect 5246 35175 5255 35176
rect 5312 35175 5326 35227
rect 5391 35201 5392 35227
rect 5471 35201 5495 35257
rect 5551 35201 5663 35257
rect 5378 35176 5392 35201
rect 5444 35176 5663 35201
rect 5391 35175 5392 35176
rect 4663 35163 4775 35175
rect 4831 35163 4855 35175
rect 4911 35163 4935 35175
rect 4991 35163 5015 35175
rect 5071 35163 5095 35175
rect 5151 35163 5175 35175
rect 5231 35163 5255 35175
rect 5311 35163 5335 35175
rect 5391 35163 5415 35175
rect 4663 35111 4666 35163
rect 4718 35111 4732 35163
rect 4850 35120 4855 35163
rect 4784 35111 4798 35120
rect 4850 35111 4864 35120
rect 4916 35111 4930 35163
rect 4991 35120 4996 35163
rect 5246 35120 5255 35163
rect 4982 35111 4996 35120
rect 5048 35111 5062 35120
rect 5114 35111 5128 35120
rect 5180 35111 5194 35120
rect 5246 35111 5260 35120
rect 5312 35111 5326 35163
rect 5391 35120 5392 35163
rect 5471 35120 5495 35176
rect 5551 35120 5663 35176
rect 5378 35111 5392 35120
rect 5444 35111 5663 35120
rect 4663 35099 5663 35111
rect 4663 35047 4666 35099
rect 4718 35047 4732 35099
rect 4784 35095 4798 35099
rect 4850 35095 4864 35099
rect 4850 35047 4855 35095
rect 4916 35047 4930 35099
rect 4982 35095 4996 35099
rect 5048 35095 5062 35099
rect 5114 35095 5128 35099
rect 5180 35095 5194 35099
rect 5246 35095 5260 35099
rect 4991 35047 4996 35095
rect 5246 35047 5255 35095
rect 5312 35047 5326 35099
rect 5378 35095 5392 35099
rect 5444 35095 5663 35099
rect 5391 35047 5392 35095
rect 4663 35039 4775 35047
rect 4831 35039 4855 35047
rect 4911 35039 4935 35047
rect 4991 35039 5015 35047
rect 5071 35039 5095 35047
rect 5151 35039 5175 35047
rect 5231 35039 5255 35047
rect 5311 35039 5335 35047
rect 5391 35039 5415 35047
rect 5471 35039 5495 35095
rect 5551 35039 5663 35095
rect 4663 35035 5663 35039
rect 4663 34983 4666 35035
rect 4718 34983 4732 35035
rect 4784 35014 4798 35035
rect 4850 35014 4864 35035
rect 4850 34983 4855 35014
rect 4916 34983 4930 35035
rect 4982 35014 4996 35035
rect 5048 35014 5062 35035
rect 5114 35014 5128 35035
rect 5180 35014 5194 35035
rect 5246 35014 5260 35035
rect 4991 34983 4996 35014
rect 5246 34983 5255 35014
rect 5312 34983 5326 35035
rect 5378 35014 5392 35035
rect 5444 35014 5663 35035
rect 5391 34983 5392 35014
rect 4663 34971 4775 34983
rect 4831 34971 4855 34983
rect 4911 34971 4935 34983
rect 4991 34971 5015 34983
rect 5071 34971 5095 34983
rect 5151 34971 5175 34983
rect 5231 34971 5255 34983
rect 5311 34971 5335 34983
rect 5391 34971 5415 34983
rect 4663 34919 4666 34971
rect 4718 34919 4732 34971
rect 4850 34958 4855 34971
rect 4784 34933 4798 34958
rect 4850 34933 4864 34958
rect 4850 34919 4855 34933
rect 4916 34919 4930 34971
rect 4991 34958 4996 34971
rect 5246 34958 5255 34971
rect 4982 34933 4996 34958
rect 5048 34933 5062 34958
rect 5114 34933 5128 34958
rect 5180 34933 5194 34958
rect 5246 34933 5260 34958
rect 4991 34919 4996 34933
rect 5246 34919 5255 34933
rect 5312 34919 5326 34971
rect 5391 34958 5392 34971
rect 5471 34958 5495 35014
rect 5551 34958 5663 35014
rect 5378 34933 5392 34958
rect 5444 34933 5663 34958
rect 5391 34919 5392 34933
rect 4663 34907 4775 34919
rect 4831 34907 4855 34919
rect 4911 34907 4935 34919
rect 4991 34907 5015 34919
rect 5071 34907 5095 34919
rect 5151 34907 5175 34919
rect 5231 34907 5255 34919
rect 5311 34907 5335 34919
rect 5391 34907 5415 34919
rect 4663 34855 4666 34907
rect 4718 34855 4732 34907
rect 4850 34877 4855 34907
rect 4784 34855 4798 34877
rect 4850 34855 4864 34877
rect 4916 34855 4930 34907
rect 4991 34877 4996 34907
rect 5246 34877 5255 34907
rect 4982 34855 4996 34877
rect 5048 34855 5062 34877
rect 5114 34855 5128 34877
rect 5180 34855 5194 34877
rect 5246 34855 5260 34877
rect 5312 34855 5326 34907
rect 5391 34877 5392 34907
rect 5471 34877 5495 34933
rect 5551 34877 5663 34933
rect 5378 34855 5392 34877
rect 5444 34855 5663 34877
rect 4663 34852 5663 34855
rect 4663 34843 4775 34852
rect 4831 34843 4855 34852
rect 4911 34843 4935 34852
rect 4991 34843 5015 34852
rect 5071 34843 5095 34852
rect 5151 34843 5175 34852
rect 5231 34843 5255 34852
rect 5311 34843 5335 34852
rect 5391 34843 5415 34852
rect 4663 34791 4666 34843
rect 4718 34791 4732 34843
rect 4850 34796 4855 34843
rect 4784 34791 4798 34796
rect 4850 34791 4864 34796
rect 4916 34791 4930 34843
rect 4991 34796 4996 34843
rect 5246 34796 5255 34843
rect 4982 34791 4996 34796
rect 5048 34791 5062 34796
rect 5114 34791 5128 34796
rect 5180 34791 5194 34796
rect 5246 34791 5260 34796
rect 5312 34791 5326 34843
rect 5391 34796 5392 34843
rect 5471 34796 5495 34852
rect 5551 34796 5663 34852
rect 5378 34791 5392 34796
rect 5444 34791 5663 34796
rect 4663 34779 5663 34791
rect 4663 34727 4666 34779
rect 4718 34727 4732 34779
rect 4784 34771 4798 34779
rect 4850 34771 4864 34779
rect 4850 34727 4855 34771
rect 4916 34727 4930 34779
rect 4982 34771 4996 34779
rect 5048 34771 5062 34779
rect 5114 34771 5128 34779
rect 5180 34771 5194 34779
rect 5246 34771 5260 34779
rect 4991 34727 4996 34771
rect 5246 34727 5255 34771
rect 5312 34727 5326 34779
rect 5378 34771 5392 34779
rect 5444 34771 5663 34779
rect 5391 34727 5392 34771
rect 4663 34715 4775 34727
rect 4831 34715 4855 34727
rect 4911 34715 4935 34727
rect 4991 34715 5015 34727
rect 5071 34715 5095 34727
rect 5151 34715 5175 34727
rect 5231 34715 5255 34727
rect 5311 34715 5335 34727
rect 5391 34715 5415 34727
rect 5471 34715 5495 34771
rect 5551 34715 5663 34771
rect 4663 34663 4666 34715
rect 4718 34663 4732 34715
rect 4784 34690 4798 34715
rect 4850 34690 4864 34715
rect 4850 34663 4855 34690
rect 4916 34663 4930 34715
rect 4982 34690 4996 34715
rect 5048 34690 5062 34715
rect 5114 34690 5128 34715
rect 5180 34690 5194 34715
rect 5246 34690 5260 34715
rect 4991 34663 4996 34690
rect 5246 34663 5255 34690
rect 5312 34663 5326 34715
rect 5378 34690 5392 34715
rect 5444 34690 5663 34715
rect 5391 34663 5392 34690
rect 4663 34651 4775 34663
rect 4831 34651 4855 34663
rect 4911 34651 4935 34663
rect 4991 34651 5015 34663
rect 5071 34651 5095 34663
rect 5151 34651 5175 34663
rect 5231 34651 5255 34663
rect 5311 34651 5335 34663
rect 5391 34651 5415 34663
rect 4663 34599 4666 34651
rect 4718 34599 4732 34651
rect 4850 34634 4855 34651
rect 4784 34609 4798 34634
rect 4850 34609 4864 34634
rect 4850 34599 4855 34609
rect 4916 34599 4930 34651
rect 4991 34634 4996 34651
rect 5246 34634 5255 34651
rect 4982 34609 4996 34634
rect 5048 34609 5062 34634
rect 5114 34609 5128 34634
rect 5180 34609 5194 34634
rect 5246 34609 5260 34634
rect 4991 34599 4996 34609
rect 5246 34599 5255 34609
rect 5312 34599 5326 34651
rect 5391 34634 5392 34651
rect 5471 34634 5495 34690
rect 5551 34634 5663 34690
rect 5378 34609 5392 34634
rect 5444 34609 5663 34634
rect 5391 34599 5392 34609
rect 4663 34587 4775 34599
rect 4831 34587 4855 34599
rect 4911 34587 4935 34599
rect 4991 34587 5015 34599
rect 5071 34587 5095 34599
rect 5151 34587 5175 34599
rect 5231 34587 5255 34599
rect 5311 34587 5335 34599
rect 5391 34587 5415 34599
rect 4663 34535 4666 34587
rect 4718 34535 4732 34587
rect 4850 34553 4855 34587
rect 4784 34535 4798 34553
rect 4850 34535 4864 34553
rect 4916 34535 4930 34587
rect 4991 34553 4996 34587
rect 5246 34553 5255 34587
rect 4982 34535 4996 34553
rect 5048 34535 5062 34553
rect 5114 34535 5128 34553
rect 5180 34535 5194 34553
rect 5246 34535 5260 34553
rect 5312 34535 5326 34587
rect 5391 34553 5392 34587
rect 5471 34553 5495 34609
rect 5551 34553 5663 34609
rect 5378 34535 5392 34553
rect 5444 34535 5663 34553
rect 4663 34528 5663 34535
rect 4663 34523 4775 34528
rect 4831 34523 4855 34528
rect 4911 34523 4935 34528
rect 4991 34523 5015 34528
rect 5071 34523 5095 34528
rect 5151 34523 5175 34528
rect 5231 34523 5255 34528
rect 5311 34523 5335 34528
rect 5391 34523 5415 34528
rect 4663 34471 4666 34523
rect 4718 34471 4732 34523
rect 4850 34472 4855 34523
rect 4784 34471 4798 34472
rect 4850 34471 4864 34472
rect 4916 34471 4930 34523
rect 4991 34472 4996 34523
rect 5246 34472 5255 34523
rect 4982 34471 4996 34472
rect 5048 34471 5062 34472
rect 5114 34471 5128 34472
rect 5180 34471 5194 34472
rect 5246 34471 5260 34472
rect 5312 34471 5326 34523
rect 5391 34472 5392 34523
rect 5471 34472 5495 34528
rect 5551 34472 5663 34528
rect 5378 34471 5392 34472
rect 5444 34471 5663 34472
rect 4663 34459 5663 34471
rect 4663 34407 4666 34459
rect 4718 34407 4732 34459
rect 4784 34447 4798 34459
rect 4850 34447 4864 34459
rect 4850 34407 4855 34447
rect 4916 34407 4930 34459
rect 4982 34447 4996 34459
rect 5048 34447 5062 34459
rect 5114 34447 5128 34459
rect 5180 34447 5194 34459
rect 5246 34447 5260 34459
rect 4991 34407 4996 34447
rect 5246 34407 5255 34447
rect 5312 34407 5326 34459
rect 5378 34447 5392 34459
rect 5444 34447 5663 34459
rect 5391 34407 5392 34447
rect 4663 34395 4775 34407
rect 4831 34395 4855 34407
rect 4911 34395 4935 34407
rect 4991 34395 5015 34407
rect 5071 34395 5095 34407
rect 5151 34395 5175 34407
rect 5231 34395 5255 34407
rect 5311 34395 5335 34407
rect 5391 34395 5415 34407
rect 4663 34343 4666 34395
rect 4718 34343 4732 34395
rect 4850 34391 4855 34395
rect 4784 34366 4798 34391
rect 4850 34366 4864 34391
rect 4850 34343 4855 34366
rect 4916 34343 4930 34395
rect 4991 34391 4996 34395
rect 5246 34391 5255 34395
rect 4982 34366 4996 34391
rect 5048 34366 5062 34391
rect 5114 34366 5128 34391
rect 5180 34366 5194 34391
rect 5246 34366 5260 34391
rect 4991 34343 4996 34366
rect 5246 34343 5255 34366
rect 5312 34343 5326 34395
rect 5391 34391 5392 34395
rect 5471 34391 5495 34447
rect 5551 34391 5663 34447
rect 5378 34366 5392 34391
rect 5444 34366 5663 34391
rect 5391 34343 5392 34366
rect 4663 34331 4775 34343
rect 4831 34331 4855 34343
rect 4911 34331 4935 34343
rect 4991 34331 5015 34343
rect 5071 34331 5095 34343
rect 5151 34331 5175 34343
rect 5231 34331 5255 34343
rect 5311 34331 5335 34343
rect 5391 34331 5415 34343
rect 4663 34279 4666 34331
rect 4718 34279 4732 34331
rect 4850 34310 4855 34331
rect 4784 34285 4798 34310
rect 4850 34285 4864 34310
rect 4850 34279 4855 34285
rect 4916 34279 4930 34331
rect 4991 34310 4996 34331
rect 5246 34310 5255 34331
rect 4982 34285 4996 34310
rect 5048 34285 5062 34310
rect 5114 34285 5128 34310
rect 5180 34285 5194 34310
rect 5246 34285 5260 34310
rect 4991 34279 4996 34285
rect 5246 34279 5255 34285
rect 5312 34279 5326 34331
rect 5391 34310 5392 34331
rect 5471 34310 5495 34366
rect 5551 34310 5663 34366
rect 5378 34285 5392 34310
rect 5444 34285 5663 34310
rect 5391 34279 5392 34285
rect 4663 34267 4775 34279
rect 4831 34267 4855 34279
rect 4911 34267 4935 34279
rect 4991 34267 5015 34279
rect 5071 34267 5095 34279
rect 5151 34267 5175 34279
rect 5231 34267 5255 34279
rect 5311 34267 5335 34279
rect 5391 34267 5415 34279
rect 4663 34215 4666 34267
rect 4718 34215 4732 34267
rect 4850 34229 4855 34267
rect 4784 34215 4798 34229
rect 4850 34215 4864 34229
rect 4916 34215 4930 34267
rect 4991 34229 4996 34267
rect 5246 34229 5255 34267
rect 4982 34215 4996 34229
rect 5048 34215 5062 34229
rect 5114 34215 5128 34229
rect 5180 34215 5194 34229
rect 5246 34215 5260 34229
rect 5312 34215 5326 34267
rect 5391 34229 5392 34267
rect 5471 34229 5495 34285
rect 5551 34229 5663 34285
rect 5378 34215 5392 34229
rect 5444 34215 5663 34229
rect 4663 34204 5663 34215
rect 4663 34203 4775 34204
rect 4831 34203 4855 34204
rect 4911 34203 4935 34204
rect 4991 34203 5015 34204
rect 5071 34203 5095 34204
rect 5151 34203 5175 34204
rect 5231 34203 5255 34204
rect 5311 34203 5335 34204
rect 5391 34203 5415 34204
rect 4663 34151 4666 34203
rect 4718 34151 4732 34203
rect 4850 34151 4855 34203
rect 4916 34151 4930 34203
rect 4991 34151 4996 34203
rect 5246 34151 5255 34203
rect 5312 34151 5326 34203
rect 5391 34151 5392 34203
rect 4663 34148 4775 34151
rect 4831 34148 4855 34151
rect 4911 34148 4935 34151
rect 4991 34148 5015 34151
rect 5071 34148 5095 34151
rect 5151 34148 5175 34151
rect 5231 34148 5255 34151
rect 5311 34148 5335 34151
rect 5391 34148 5415 34151
rect 5471 34148 5495 34204
rect 5551 34148 5663 34204
rect 4663 34139 5663 34148
rect 4663 34087 4666 34139
rect 4718 34087 4732 34139
rect 4784 34123 4798 34139
rect 4850 34123 4864 34139
rect 4850 34087 4855 34123
rect 4916 34087 4930 34139
rect 4982 34123 4996 34139
rect 5048 34123 5062 34139
rect 5114 34123 5128 34139
rect 5180 34123 5194 34139
rect 5246 34123 5260 34139
rect 4991 34087 4996 34123
rect 5246 34087 5255 34123
rect 5312 34087 5326 34139
rect 5378 34123 5392 34139
rect 5444 34123 5663 34139
rect 5391 34087 5392 34123
rect 4663 34075 4775 34087
rect 4831 34075 4855 34087
rect 4911 34075 4935 34087
rect 4991 34075 5015 34087
rect 5071 34075 5095 34087
rect 5151 34075 5175 34087
rect 5231 34075 5255 34087
rect 5311 34075 5335 34087
rect 5391 34075 5415 34087
rect 4663 34023 4666 34075
rect 4718 34023 4732 34075
rect 4850 34067 4855 34075
rect 4784 34042 4798 34067
rect 4850 34042 4864 34067
rect 4850 34023 4855 34042
rect 4916 34023 4930 34075
rect 4991 34067 4996 34075
rect 5246 34067 5255 34075
rect 4982 34042 4996 34067
rect 5048 34042 5062 34067
rect 5114 34042 5128 34067
rect 5180 34042 5194 34067
rect 5246 34042 5260 34067
rect 4991 34023 4996 34042
rect 5246 34023 5255 34042
rect 5312 34023 5326 34075
rect 5391 34067 5392 34075
rect 5471 34067 5495 34123
rect 5551 34067 5663 34123
rect 5378 34042 5392 34067
rect 5444 34042 5663 34067
rect 5391 34023 5392 34042
rect 4663 34011 4775 34023
rect 4831 34011 4855 34023
rect 4911 34011 4935 34023
rect 4991 34011 5015 34023
rect 5071 34011 5095 34023
rect 5151 34011 5175 34023
rect 5231 34011 5255 34023
rect 5311 34011 5335 34023
rect 5391 34011 5415 34023
rect 4663 33959 4666 34011
rect 4718 33959 4732 34011
rect 4850 33986 4855 34011
rect 4784 33961 4798 33986
rect 4850 33961 4864 33986
rect 4850 33959 4855 33961
rect 4916 33959 4930 34011
rect 4991 33986 4996 34011
rect 5246 33986 5255 34011
rect 4982 33961 4996 33986
rect 5048 33961 5062 33986
rect 5114 33961 5128 33986
rect 5180 33961 5194 33986
rect 5246 33961 5260 33986
rect 4991 33959 4996 33961
rect 5246 33959 5255 33961
rect 5312 33959 5326 34011
rect 5391 33986 5392 34011
rect 5471 33986 5495 34042
rect 5551 33986 5663 34042
rect 5378 33961 5392 33986
rect 5444 33961 5663 33986
rect 5391 33959 5392 33961
rect 4663 33947 4775 33959
rect 4831 33947 4855 33959
rect 4911 33947 4935 33959
rect 4991 33947 5015 33959
rect 5071 33947 5095 33959
rect 5151 33947 5175 33959
rect 5231 33947 5255 33959
rect 5311 33947 5335 33959
rect 5391 33947 5415 33959
rect 4663 33895 4666 33947
rect 4718 33895 4732 33947
rect 4850 33905 4855 33947
rect 4784 33895 4798 33905
rect 4850 33895 4864 33905
rect 4916 33895 4930 33947
rect 4991 33905 4996 33947
rect 5246 33905 5255 33947
rect 4982 33895 4996 33905
rect 5048 33895 5062 33905
rect 5114 33895 5128 33905
rect 5180 33895 5194 33905
rect 5246 33895 5260 33905
rect 5312 33895 5326 33947
rect 5391 33905 5392 33947
rect 5471 33905 5495 33961
rect 5551 33905 5663 33961
rect 5378 33895 5392 33905
rect 5444 33895 5663 33905
rect 4663 33883 5663 33895
rect 4663 33831 4666 33883
rect 4718 33831 4732 33883
rect 4784 33880 4798 33883
rect 4850 33880 4864 33883
rect 4850 33831 4855 33880
rect 4916 33831 4930 33883
rect 4982 33880 4996 33883
rect 5048 33880 5062 33883
rect 5114 33880 5128 33883
rect 5180 33880 5194 33883
rect 5246 33880 5260 33883
rect 4991 33831 4996 33880
rect 5246 33831 5255 33880
rect 5312 33831 5326 33883
rect 5378 33880 5392 33883
rect 5444 33880 5663 33883
rect 5391 33831 5392 33880
rect 4663 33824 4775 33831
rect 4831 33824 4855 33831
rect 4911 33824 4935 33831
rect 4991 33824 5015 33831
rect 5071 33824 5095 33831
rect 5151 33824 5175 33831
rect 5231 33824 5255 33831
rect 5311 33824 5335 33831
rect 5391 33824 5415 33831
rect 5471 33824 5495 33880
rect 5551 33824 5663 33880
rect 4663 33819 5663 33824
rect 4663 33767 4666 33819
rect 4718 33767 4732 33819
rect 4784 33799 4798 33819
rect 4850 33799 4864 33819
rect 4850 33767 4855 33799
rect 4916 33767 4930 33819
rect 4982 33799 4996 33819
rect 5048 33799 5062 33819
rect 5114 33799 5128 33819
rect 5180 33799 5194 33819
rect 5246 33799 5260 33819
rect 4991 33767 4996 33799
rect 5246 33767 5255 33799
rect 5312 33767 5326 33819
rect 5378 33799 5392 33819
rect 5444 33799 5663 33819
rect 5391 33767 5392 33799
rect 4663 33755 4775 33767
rect 4831 33755 4855 33767
rect 4911 33755 4935 33767
rect 4991 33755 5015 33767
rect 5071 33755 5095 33767
rect 5151 33755 5175 33767
rect 5231 33755 5255 33767
rect 5311 33755 5335 33767
rect 5391 33755 5415 33767
rect 4663 33703 4666 33755
rect 4718 33703 4732 33755
rect 4850 33743 4855 33755
rect 4784 33718 4798 33743
rect 4850 33718 4864 33743
rect 4850 33703 4855 33718
rect 4916 33703 4930 33755
rect 4991 33743 4996 33755
rect 5246 33743 5255 33755
rect 4982 33718 4996 33743
rect 5048 33718 5062 33743
rect 5114 33718 5128 33743
rect 5180 33718 5194 33743
rect 5246 33718 5260 33743
rect 4991 33703 4996 33718
rect 5246 33703 5255 33718
rect 5312 33703 5326 33755
rect 5391 33743 5392 33755
rect 5471 33743 5495 33799
rect 5551 33743 5663 33799
rect 5378 33718 5392 33743
rect 5444 33718 5663 33743
rect 5391 33703 5392 33718
rect 4663 33691 4775 33703
rect 4831 33691 4855 33703
rect 4911 33691 4935 33703
rect 4991 33691 5015 33703
rect 5071 33691 5095 33703
rect 5151 33691 5175 33703
rect 5231 33691 5255 33703
rect 5311 33691 5335 33703
rect 5391 33691 5415 33703
rect 4663 33639 4666 33691
rect 4718 33639 4732 33691
rect 4850 33662 4855 33691
rect 4784 33639 4798 33662
rect 4850 33639 4864 33662
rect 4916 33639 4930 33691
rect 4991 33662 4996 33691
rect 5246 33662 5255 33691
rect 4982 33639 4996 33662
rect 5048 33639 5062 33662
rect 5114 33639 5128 33662
rect 5180 33639 5194 33662
rect 5246 33639 5260 33662
rect 5312 33639 5326 33691
rect 5391 33662 5392 33691
rect 5471 33662 5495 33718
rect 5551 33662 5663 33718
rect 5378 33639 5392 33662
rect 5444 33639 5663 33662
rect 4663 33637 5663 33639
rect 4663 33627 4775 33637
rect 4831 33627 4855 33637
rect 4911 33627 4935 33637
rect 4991 33627 5015 33637
rect 5071 33627 5095 33637
rect 5151 33627 5175 33637
rect 5231 33627 5255 33637
rect 5311 33627 5335 33637
rect 5391 33627 5415 33637
rect 4663 33575 4666 33627
rect 4718 33575 4732 33627
rect 4850 33581 4855 33627
rect 4784 33575 4798 33581
rect 4850 33575 4864 33581
rect 4916 33575 4930 33627
rect 4991 33581 4996 33627
rect 5246 33581 5255 33627
rect 4982 33575 4996 33581
rect 5048 33575 5062 33581
rect 5114 33575 5128 33581
rect 5180 33575 5194 33581
rect 5246 33575 5260 33581
rect 5312 33575 5326 33627
rect 5391 33581 5392 33627
rect 5471 33581 5495 33637
rect 5551 33581 5663 33637
rect 5378 33575 5392 33581
rect 5444 33575 5663 33581
rect 4663 33563 5663 33575
rect 4663 33511 4666 33563
rect 4718 33511 4732 33563
rect 4784 33556 4798 33563
rect 4850 33556 4864 33563
rect 4850 33511 4855 33556
rect 4916 33511 4930 33563
rect 4982 33556 4996 33563
rect 5048 33556 5062 33563
rect 5114 33556 5128 33563
rect 5180 33556 5194 33563
rect 5246 33556 5260 33563
rect 4991 33511 4996 33556
rect 5246 33511 5255 33556
rect 5312 33511 5326 33563
rect 5378 33556 5392 33563
rect 5444 33556 5663 33563
rect 5391 33511 5392 33556
rect 4663 33500 4775 33511
rect 4831 33500 4855 33511
rect 4911 33500 4935 33511
rect 4991 33500 5015 33511
rect 5071 33500 5095 33511
rect 5151 33500 5175 33511
rect 5231 33500 5255 33511
rect 5311 33500 5335 33511
rect 5391 33500 5415 33511
rect 5471 33500 5495 33556
rect 5551 33500 5663 33556
rect 4663 33499 5663 33500
rect 4663 33447 4666 33499
rect 4718 33447 4732 33499
rect 4784 33475 4798 33499
rect 4850 33475 4864 33499
rect 4850 33447 4855 33475
rect 4916 33447 4930 33499
rect 4982 33475 4996 33499
rect 5048 33475 5062 33499
rect 5114 33475 5128 33499
rect 5180 33475 5194 33499
rect 5246 33475 5260 33499
rect 4991 33447 4996 33475
rect 5246 33447 5255 33475
rect 5312 33447 5326 33499
rect 5378 33475 5392 33499
rect 5444 33475 5663 33499
rect 5391 33447 5392 33475
rect 4663 33435 4775 33447
rect 4831 33435 4855 33447
rect 4911 33435 4935 33447
rect 4991 33435 5015 33447
rect 5071 33435 5095 33447
rect 5151 33435 5175 33447
rect 5231 33435 5255 33447
rect 5311 33435 5335 33447
rect 5391 33435 5415 33447
rect 4663 33383 4666 33435
rect 4718 33383 4732 33435
rect 4850 33419 4855 33435
rect 4784 33394 4798 33419
rect 4850 33394 4864 33419
rect 4850 33383 4855 33394
rect 4916 33383 4930 33435
rect 4991 33419 4996 33435
rect 5246 33419 5255 33435
rect 4982 33394 4996 33419
rect 5048 33394 5062 33419
rect 5114 33394 5128 33419
rect 5180 33394 5194 33419
rect 5246 33394 5260 33419
rect 4991 33383 4996 33394
rect 5246 33383 5255 33394
rect 5312 33383 5326 33435
rect 5391 33419 5392 33435
rect 5471 33419 5495 33475
rect 5551 33419 5663 33475
rect 5378 33394 5392 33419
rect 5444 33394 5663 33419
rect 5391 33383 5392 33394
rect 4663 33371 4775 33383
rect 4831 33371 4855 33383
rect 4911 33371 4935 33383
rect 4991 33371 5015 33383
rect 5071 33371 5095 33383
rect 5151 33371 5175 33383
rect 5231 33371 5255 33383
rect 5311 33371 5335 33383
rect 5391 33371 5415 33383
rect 4663 33319 4666 33371
rect 4718 33319 4732 33371
rect 4850 33338 4855 33371
rect 4784 33319 4798 33338
rect 4850 33319 4864 33338
rect 4916 33319 4930 33371
rect 4991 33338 4996 33371
rect 5246 33338 5255 33371
rect 4982 33319 4996 33338
rect 5048 33319 5062 33338
rect 5114 33319 5128 33338
rect 5180 33319 5194 33338
rect 5246 33319 5260 33338
rect 5312 33319 5326 33371
rect 5391 33338 5392 33371
rect 5471 33338 5495 33394
rect 5551 33338 5663 33394
rect 5378 33319 5392 33338
rect 5444 33319 5663 33338
rect 4663 33313 5663 33319
rect 4663 33307 4775 33313
rect 4831 33307 4855 33313
rect 4911 33307 4935 33313
rect 4991 33307 5015 33313
rect 5071 33307 5095 33313
rect 5151 33307 5175 33313
rect 5231 33307 5255 33313
rect 5311 33307 5335 33313
rect 5391 33307 5415 33313
rect 4663 33255 4666 33307
rect 4718 33255 4732 33307
rect 4850 33257 4855 33307
rect 4784 33255 4798 33257
rect 4850 33255 4864 33257
rect 4916 33255 4930 33307
rect 4991 33257 4996 33307
rect 5246 33257 5255 33307
rect 4982 33255 4996 33257
rect 5048 33255 5062 33257
rect 5114 33255 5128 33257
rect 5180 33255 5194 33257
rect 5246 33255 5260 33257
rect 5312 33255 5326 33307
rect 5391 33257 5392 33307
rect 5471 33257 5495 33313
rect 5551 33257 5663 33313
rect 5378 33255 5392 33257
rect 5444 33255 5663 33257
rect 4663 33243 5663 33255
rect 4663 33191 4666 33243
rect 4718 33191 4732 33243
rect 4784 33232 4798 33243
rect 4850 33232 4864 33243
rect 4850 33191 4855 33232
rect 4916 33191 4930 33243
rect 4982 33232 4996 33243
rect 5048 33232 5062 33243
rect 5114 33232 5128 33243
rect 5180 33232 5194 33243
rect 5246 33232 5260 33243
rect 4991 33191 4996 33232
rect 5246 33191 5255 33232
rect 5312 33191 5326 33243
rect 5378 33232 5392 33243
rect 5444 33232 5663 33243
rect 5391 33191 5392 33232
rect 4663 33179 4775 33191
rect 4831 33179 4855 33191
rect 4911 33179 4935 33191
rect 4991 33179 5015 33191
rect 5071 33179 5095 33191
rect 5151 33179 5175 33191
rect 5231 33179 5255 33191
rect 5311 33179 5335 33191
rect 5391 33179 5415 33191
rect 4663 33127 4666 33179
rect 4718 33127 4732 33179
rect 4850 33176 4855 33179
rect 4784 33151 4798 33176
rect 4850 33151 4864 33176
rect 4850 33127 4855 33151
rect 4916 33127 4930 33179
rect 4991 33176 4996 33179
rect 5246 33176 5255 33179
rect 4982 33151 4996 33176
rect 5048 33151 5062 33176
rect 5114 33151 5128 33176
rect 5180 33151 5194 33176
rect 5246 33151 5260 33176
rect 4991 33127 4996 33151
rect 5246 33127 5255 33151
rect 5312 33127 5326 33179
rect 5391 33176 5392 33179
rect 5471 33176 5495 33232
rect 5551 33176 5663 33232
rect 5378 33151 5392 33176
rect 5444 33151 5663 33176
rect 5391 33127 5392 33151
rect 4663 33115 4775 33127
rect 4831 33115 4855 33127
rect 4911 33115 4935 33127
rect 4991 33115 5015 33127
rect 5071 33115 5095 33127
rect 5151 33115 5175 33127
rect 5231 33115 5255 33127
rect 5311 33115 5335 33127
rect 5391 33115 5415 33127
rect 4663 33063 4666 33115
rect 4718 33063 4732 33115
rect 4850 33095 4855 33115
rect 4784 33070 4798 33095
rect 4850 33070 4864 33095
rect 4850 33063 4855 33070
rect 4916 33063 4930 33115
rect 4991 33095 4996 33115
rect 5246 33095 5255 33115
rect 4982 33070 4996 33095
rect 5048 33070 5062 33095
rect 5114 33070 5128 33095
rect 5180 33070 5194 33095
rect 5246 33070 5260 33095
rect 4991 33063 4996 33070
rect 5246 33063 5255 33070
rect 5312 33063 5326 33115
rect 5391 33095 5392 33115
rect 5471 33095 5495 33151
rect 5551 33095 5663 33151
rect 5378 33070 5392 33095
rect 5444 33070 5663 33095
rect 5391 33063 5392 33070
rect 4663 33051 4775 33063
rect 4831 33051 4855 33063
rect 4911 33051 4935 33063
rect 4991 33051 5015 33063
rect 5071 33051 5095 33063
rect 5151 33051 5175 33063
rect 5231 33051 5255 33063
rect 5311 33051 5335 33063
rect 5391 33051 5415 33063
rect 4663 32999 4666 33051
rect 4718 32999 4732 33051
rect 4850 33014 4855 33051
rect 4784 32999 4798 33014
rect 4850 32999 4864 33014
rect 4916 32999 4930 33051
rect 4991 33014 4996 33051
rect 5246 33014 5255 33051
rect 4982 32999 4996 33014
rect 5048 32999 5062 33014
rect 5114 32999 5128 33014
rect 5180 32999 5194 33014
rect 5246 32999 5260 33014
rect 5312 32999 5326 33051
rect 5391 33014 5392 33051
rect 5471 33014 5495 33070
rect 5551 33014 5663 33070
rect 5378 32999 5392 33014
rect 5444 32999 5663 33014
rect 4663 32989 5663 32999
rect 4663 32987 4775 32989
rect 4831 32987 4855 32989
rect 4911 32987 4935 32989
rect 4991 32987 5015 32989
rect 5071 32987 5095 32989
rect 5151 32987 5175 32989
rect 5231 32987 5255 32989
rect 5311 32987 5335 32989
rect 5391 32987 5415 32989
rect 4663 32935 4666 32987
rect 4718 32935 4732 32987
rect 4850 32935 4855 32987
rect 4916 32935 4930 32987
rect 4991 32935 4996 32987
rect 5246 32935 5255 32987
rect 5312 32935 5326 32987
rect 5391 32935 5392 32987
rect 4663 32933 4775 32935
rect 4831 32933 4855 32935
rect 4911 32933 4935 32935
rect 4991 32933 5015 32935
rect 5071 32933 5095 32935
rect 5151 32933 5175 32935
rect 5231 32933 5255 32935
rect 5311 32933 5335 32935
rect 5391 32933 5415 32935
rect 5471 32933 5495 32989
rect 5551 32933 5663 32989
rect 4663 32923 5663 32933
rect 4663 32871 4666 32923
rect 4718 32871 4732 32923
rect 4784 32908 4798 32923
rect 4850 32908 4864 32923
rect 4850 32871 4855 32908
rect 4916 32871 4930 32923
rect 4982 32908 4996 32923
rect 5048 32908 5062 32923
rect 5114 32908 5128 32923
rect 5180 32908 5194 32923
rect 5246 32908 5260 32923
rect 4991 32871 4996 32908
rect 5246 32871 5255 32908
rect 5312 32871 5326 32923
rect 5378 32908 5392 32923
rect 5444 32908 5663 32923
rect 5391 32871 5392 32908
rect 4663 32859 4775 32871
rect 4831 32859 4855 32871
rect 4911 32859 4935 32871
rect 4991 32859 5015 32871
rect 5071 32859 5095 32871
rect 5151 32859 5175 32871
rect 5231 32859 5255 32871
rect 5311 32859 5335 32871
rect 5391 32859 5415 32871
rect 4663 32807 4666 32859
rect 4718 32807 4732 32859
rect 4850 32852 4855 32859
rect 4784 32827 4798 32852
rect 4850 32827 4864 32852
rect 4850 32807 4855 32827
rect 4916 32807 4930 32859
rect 4991 32852 4996 32859
rect 5246 32852 5255 32859
rect 4982 32827 4996 32852
rect 5048 32827 5062 32852
rect 5114 32827 5128 32852
rect 5180 32827 5194 32852
rect 5246 32827 5260 32852
rect 4991 32807 4996 32827
rect 5246 32807 5255 32827
rect 5312 32807 5326 32859
rect 5391 32852 5392 32859
rect 5471 32852 5495 32908
rect 5551 32852 5663 32908
rect 5378 32827 5392 32852
rect 5444 32827 5663 32852
rect 5391 32807 5392 32827
rect 4663 32795 4775 32807
rect 4831 32795 4855 32807
rect 4911 32795 4935 32807
rect 4991 32795 5015 32807
rect 5071 32795 5095 32807
rect 5151 32795 5175 32807
rect 5231 32795 5255 32807
rect 5311 32795 5335 32807
rect 5391 32795 5415 32807
rect 4663 32743 4666 32795
rect 4718 32743 4732 32795
rect 4850 32771 4855 32795
rect 4784 32746 4798 32771
rect 4850 32746 4864 32771
rect 4850 32743 4855 32746
rect 4916 32743 4930 32795
rect 4991 32771 4996 32795
rect 5246 32771 5255 32795
rect 4982 32746 4996 32771
rect 5048 32746 5062 32771
rect 5114 32746 5128 32771
rect 5180 32746 5194 32771
rect 5246 32746 5260 32771
rect 4991 32743 4996 32746
rect 5246 32743 5255 32746
rect 5312 32743 5326 32795
rect 5391 32771 5392 32795
rect 5471 32771 5495 32827
rect 5551 32771 5663 32827
rect 5378 32746 5392 32771
rect 5444 32746 5663 32771
rect 5391 32743 5392 32746
rect 4663 32730 4775 32743
rect 4831 32730 4855 32743
rect 4911 32730 4935 32743
rect 4991 32730 5015 32743
rect 5071 32730 5095 32743
rect 5151 32730 5175 32743
rect 5231 32730 5255 32743
rect 5311 32730 5335 32743
rect 5391 32730 5415 32743
rect 4663 32678 4666 32730
rect 4718 32678 4732 32730
rect 4850 32690 4855 32730
rect 4784 32678 4798 32690
rect 4850 32678 4864 32690
rect 4916 32678 4930 32730
rect 4991 32690 4996 32730
rect 5246 32690 5255 32730
rect 4982 32678 4996 32690
rect 5048 32678 5062 32690
rect 5114 32678 5128 32690
rect 5180 32678 5194 32690
rect 5246 32678 5260 32690
rect 5312 32678 5326 32730
rect 5391 32690 5392 32730
rect 5471 32690 5495 32746
rect 5551 32690 5663 32746
rect 5378 32678 5392 32690
rect 5444 32678 5663 32690
rect 4663 32665 5663 32678
rect 4663 32613 4666 32665
rect 4718 32613 4732 32665
rect 4850 32613 4855 32665
rect 4916 32613 4930 32665
rect 4991 32613 4996 32665
rect 5246 32613 5255 32665
rect 5312 32613 5326 32665
rect 5391 32613 5392 32665
rect 4663 32609 4775 32613
rect 4831 32609 4855 32613
rect 4911 32609 4935 32613
rect 4991 32609 5015 32613
rect 5071 32609 5095 32613
rect 5151 32609 5175 32613
rect 5231 32609 5255 32613
rect 5311 32609 5335 32613
rect 5391 32609 5415 32613
rect 5471 32609 5495 32665
rect 5551 32609 5663 32665
rect 4663 32600 5663 32609
rect 4663 32548 4666 32600
rect 4718 32548 4732 32600
rect 4784 32584 4798 32600
rect 4850 32584 4864 32600
rect 4850 32548 4855 32584
rect 4916 32548 4930 32600
rect 4982 32584 4996 32600
rect 5048 32584 5062 32600
rect 5114 32584 5128 32600
rect 5180 32584 5194 32600
rect 5246 32584 5260 32600
rect 4991 32548 4996 32584
rect 5246 32548 5255 32584
rect 5312 32548 5326 32600
rect 5378 32584 5392 32600
rect 5444 32584 5663 32600
rect 5391 32548 5392 32584
rect 4663 32535 4775 32548
rect 4831 32535 4855 32548
rect 4911 32535 4935 32548
rect 4991 32535 5015 32548
rect 5071 32535 5095 32548
rect 5151 32535 5175 32548
rect 5231 32535 5255 32548
rect 5311 32535 5335 32548
rect 5391 32535 5415 32548
rect 4663 32483 4666 32535
rect 4718 32483 4732 32535
rect 4850 32528 4855 32535
rect 4784 32503 4798 32528
rect 4850 32503 4864 32528
rect 4850 32483 4855 32503
rect 4916 32483 4930 32535
rect 4991 32528 4996 32535
rect 5246 32528 5255 32535
rect 4982 32503 4996 32528
rect 5048 32503 5062 32528
rect 5114 32503 5128 32528
rect 5180 32503 5194 32528
rect 5246 32503 5260 32528
rect 4991 32483 4996 32503
rect 5246 32483 5255 32503
rect 5312 32483 5326 32535
rect 5391 32528 5392 32535
rect 5471 32528 5495 32584
rect 5551 32528 5663 32584
rect 5378 32503 5392 32528
rect 5444 32503 5663 32528
rect 5391 32483 5392 32503
rect 4663 32470 4775 32483
rect 4831 32470 4855 32483
rect 4911 32470 4935 32483
rect 4991 32470 5015 32483
rect 5071 32470 5095 32483
rect 5151 32470 5175 32483
rect 5231 32470 5255 32483
rect 5311 32470 5335 32483
rect 5391 32470 5415 32483
rect 4663 32418 4666 32470
rect 4718 32418 4732 32470
rect 4850 32447 4855 32470
rect 4784 32422 4798 32447
rect 4850 32422 4864 32447
rect 4850 32418 4855 32422
rect 4916 32418 4930 32470
rect 4991 32447 4996 32470
rect 5246 32447 5255 32470
rect 4982 32422 4996 32447
rect 5048 32422 5062 32447
rect 5114 32422 5128 32447
rect 5180 32422 5194 32447
rect 5246 32422 5260 32447
rect 4991 32418 4996 32422
rect 5246 32418 5255 32422
rect 5312 32418 5326 32470
rect 5391 32447 5392 32470
rect 5471 32447 5495 32503
rect 5551 32447 5663 32503
rect 5378 32422 5392 32447
rect 5444 32422 5663 32447
rect 5391 32418 5392 32422
rect 4663 32405 4775 32418
rect 4831 32405 4855 32418
rect 4911 32405 4935 32418
rect 4991 32405 5015 32418
rect 5071 32405 5095 32418
rect 5151 32405 5175 32418
rect 5231 32405 5255 32418
rect 5311 32405 5335 32418
rect 5391 32405 5415 32418
rect 4663 32353 4666 32405
rect 4718 32353 4732 32405
rect 4850 32366 4855 32405
rect 4784 32353 4798 32366
rect 4850 32353 4864 32366
rect 4916 32353 4930 32405
rect 4991 32366 4996 32405
rect 5246 32366 5255 32405
rect 4982 32353 4996 32366
rect 5048 32353 5062 32366
rect 5114 32353 5128 32366
rect 5180 32353 5194 32366
rect 5246 32353 5260 32366
rect 5312 32353 5326 32405
rect 5391 32366 5392 32405
rect 5471 32366 5495 32422
rect 5551 32366 5663 32422
rect 5378 32353 5392 32366
rect 5444 32353 5663 32366
rect 4663 32341 5663 32353
rect 4663 32340 4775 32341
rect 4831 32340 4855 32341
rect 4911 32340 4935 32341
rect 4991 32340 5015 32341
rect 5071 32340 5095 32341
rect 5151 32340 5175 32341
rect 5231 32340 5255 32341
rect 5311 32340 5335 32341
rect 5391 32340 5415 32341
rect 4663 32288 4666 32340
rect 4718 32288 4732 32340
rect 4850 32288 4855 32340
rect 4916 32288 4930 32340
rect 4991 32288 4996 32340
rect 5246 32288 5255 32340
rect 5312 32288 5326 32340
rect 5391 32288 5392 32340
rect 4663 32285 4775 32288
rect 4831 32285 4855 32288
rect 4911 32285 4935 32288
rect 4991 32285 5015 32288
rect 5071 32285 5095 32288
rect 5151 32285 5175 32288
rect 5231 32285 5255 32288
rect 5311 32285 5335 32288
rect 5391 32285 5415 32288
rect 5471 32285 5495 32341
rect 5551 32285 5663 32341
rect 4663 32275 5663 32285
rect 4663 32223 4666 32275
rect 4718 32223 4732 32275
rect 4784 32260 4798 32275
rect 4850 32260 4864 32275
rect 4850 32223 4855 32260
rect 4916 32223 4930 32275
rect 4982 32260 4996 32275
rect 5048 32260 5062 32275
rect 5114 32260 5128 32275
rect 5180 32260 5194 32275
rect 5246 32260 5260 32275
rect 4991 32223 4996 32260
rect 5246 32223 5255 32260
rect 5312 32223 5326 32275
rect 5378 32260 5392 32275
rect 5444 32260 5663 32275
rect 5391 32223 5392 32260
rect 4663 32210 4775 32223
rect 4831 32210 4855 32223
rect 4911 32210 4935 32223
rect 4991 32210 5015 32223
rect 5071 32210 5095 32223
rect 5151 32210 5175 32223
rect 5231 32210 5255 32223
rect 5311 32210 5335 32223
rect 5391 32210 5415 32223
rect 4663 32158 4666 32210
rect 4718 32158 4732 32210
rect 4850 32204 4855 32210
rect 4784 32179 4798 32204
rect 4850 32179 4864 32204
rect 4850 32158 4855 32179
rect 4916 32158 4930 32210
rect 4991 32204 4996 32210
rect 5246 32204 5255 32210
rect 4982 32179 4996 32204
rect 5048 32179 5062 32204
rect 5114 32179 5128 32204
rect 5180 32179 5194 32204
rect 5246 32179 5260 32204
rect 4991 32158 4996 32179
rect 5246 32158 5255 32179
rect 5312 32158 5326 32210
rect 5391 32204 5392 32210
rect 5471 32204 5495 32260
rect 5551 32204 5663 32260
rect 5378 32179 5392 32204
rect 5444 32179 5663 32204
rect 5391 32158 5392 32179
rect 4663 32145 4775 32158
rect 4831 32145 4855 32158
rect 4911 32145 4935 32158
rect 4991 32145 5015 32158
rect 5071 32145 5095 32158
rect 5151 32145 5175 32158
rect 5231 32145 5255 32158
rect 5311 32145 5335 32158
rect 5391 32145 5415 32158
rect 4663 32093 4666 32145
rect 4718 32093 4732 32145
rect 4850 32123 4855 32145
rect 4784 32098 4798 32123
rect 4850 32098 4864 32123
rect 4850 32093 4855 32098
rect 4916 32093 4930 32145
rect 4991 32123 4996 32145
rect 5246 32123 5255 32145
rect 4982 32098 4996 32123
rect 5048 32098 5062 32123
rect 5114 32098 5128 32123
rect 5180 32098 5194 32123
rect 5246 32098 5260 32123
rect 4991 32093 4996 32098
rect 5246 32093 5255 32098
rect 5312 32093 5326 32145
rect 5391 32123 5392 32145
rect 5471 32123 5495 32179
rect 5551 32123 5663 32179
rect 5378 32098 5392 32123
rect 5444 32098 5663 32123
rect 5391 32093 5392 32098
rect 4663 32080 4775 32093
rect 4831 32080 4855 32093
rect 4911 32080 4935 32093
rect 4991 32080 5015 32093
rect 5071 32080 5095 32093
rect 5151 32080 5175 32093
rect 5231 32080 5255 32093
rect 5311 32080 5335 32093
rect 5391 32080 5415 32093
rect 4663 32028 4666 32080
rect 4718 32028 4732 32080
rect 4850 32042 4855 32080
rect 4784 32028 4798 32042
rect 4850 32028 4864 32042
rect 4916 32028 4930 32080
rect 4991 32042 4996 32080
rect 5246 32042 5255 32080
rect 4982 32028 4996 32042
rect 5048 32028 5062 32042
rect 5114 32028 5128 32042
rect 5180 32028 5194 32042
rect 5246 32028 5260 32042
rect 5312 32028 5326 32080
rect 5391 32042 5392 32080
rect 5471 32042 5495 32098
rect 5551 32042 5663 32098
rect 5378 32028 5392 32042
rect 5444 32028 5663 32042
rect 4663 32017 5663 32028
rect 4663 32015 4775 32017
rect 4831 32015 4855 32017
rect 4911 32015 4935 32017
rect 4991 32015 5015 32017
rect 5071 32015 5095 32017
rect 5151 32015 5175 32017
rect 5231 32015 5255 32017
rect 5311 32015 5335 32017
rect 5391 32015 5415 32017
rect 4663 31963 4666 32015
rect 4718 31963 4732 32015
rect 4850 31963 4855 32015
rect 4916 31963 4930 32015
rect 4991 31963 4996 32015
rect 5246 31963 5255 32015
rect 5312 31963 5326 32015
rect 5391 31963 5392 32015
rect 4663 31961 4775 31963
rect 4831 31961 4855 31963
rect 4911 31961 4935 31963
rect 4991 31961 5015 31963
rect 5071 31961 5095 31963
rect 5151 31961 5175 31963
rect 5231 31961 5255 31963
rect 5311 31961 5335 31963
rect 5391 31961 5415 31963
rect 5471 31961 5495 32017
rect 5551 31961 5663 32017
rect 4663 31950 5663 31961
rect 4663 31898 4666 31950
rect 4718 31898 4732 31950
rect 4784 31936 4798 31950
rect 4850 31936 4864 31950
rect 4850 31898 4855 31936
rect 4916 31898 4930 31950
rect 4982 31936 4996 31950
rect 5048 31936 5062 31950
rect 5114 31936 5128 31950
rect 5180 31936 5194 31950
rect 5246 31936 5260 31950
rect 4991 31898 4996 31936
rect 5246 31898 5255 31936
rect 5312 31898 5326 31950
rect 5378 31936 5392 31950
rect 5444 31936 5663 31950
rect 5391 31898 5392 31936
rect 4663 31885 4775 31898
rect 4831 31885 4855 31898
rect 4911 31885 4935 31898
rect 4991 31885 5015 31898
rect 5071 31885 5095 31898
rect 5151 31885 5175 31898
rect 5231 31885 5255 31898
rect 5311 31885 5335 31898
rect 5391 31885 5415 31898
rect 4663 31833 4666 31885
rect 4718 31833 4732 31885
rect 4850 31880 4855 31885
rect 4784 31855 4798 31880
rect 4850 31855 4864 31880
rect 4850 31833 4855 31855
rect 4916 31833 4930 31885
rect 4991 31880 4996 31885
rect 5246 31880 5255 31885
rect 4982 31855 4996 31880
rect 5048 31855 5062 31880
rect 5114 31855 5128 31880
rect 5180 31855 5194 31880
rect 5246 31855 5260 31880
rect 4991 31833 4996 31855
rect 5246 31833 5255 31855
rect 5312 31833 5326 31885
rect 5391 31880 5392 31885
rect 5471 31880 5495 31936
rect 5551 31880 5663 31936
rect 5378 31855 5392 31880
rect 5444 31855 5663 31880
rect 5391 31833 5392 31855
rect 4663 31820 4775 31833
rect 4831 31820 4855 31833
rect 4911 31820 4935 31833
rect 4991 31820 5015 31833
rect 5071 31820 5095 31833
rect 5151 31820 5175 31833
rect 5231 31820 5255 31833
rect 5311 31820 5335 31833
rect 5391 31820 5415 31833
rect 4663 31768 4666 31820
rect 4718 31768 4732 31820
rect 4850 31799 4855 31820
rect 4784 31774 4798 31799
rect 4850 31774 4864 31799
rect 4850 31768 4855 31774
rect 4916 31768 4930 31820
rect 4991 31799 4996 31820
rect 5246 31799 5255 31820
rect 4982 31774 4996 31799
rect 5048 31774 5062 31799
rect 5114 31774 5128 31799
rect 5180 31774 5194 31799
rect 5246 31774 5260 31799
rect 4991 31768 4996 31774
rect 5246 31768 5255 31774
rect 5312 31768 5326 31820
rect 5391 31799 5392 31820
rect 5471 31799 5495 31855
rect 5551 31799 5663 31855
rect 5378 31774 5392 31799
rect 5444 31774 5663 31799
rect 5391 31768 5392 31774
rect 4663 31755 4775 31768
rect 4831 31755 4855 31768
rect 4911 31755 4935 31768
rect 4991 31755 5015 31768
rect 5071 31755 5095 31768
rect 5151 31755 5175 31768
rect 5231 31755 5255 31768
rect 5311 31755 5335 31768
rect 5391 31755 5415 31768
rect 4663 31703 4666 31755
rect 4718 31703 4732 31755
rect 4850 31718 4855 31755
rect 4784 31703 4798 31718
rect 4850 31703 4864 31718
rect 4916 31703 4930 31755
rect 4991 31718 4996 31755
rect 5246 31718 5255 31755
rect 4982 31703 4996 31718
rect 5048 31703 5062 31718
rect 5114 31703 5128 31718
rect 5180 31703 5194 31718
rect 5246 31703 5260 31718
rect 5312 31703 5326 31755
rect 5391 31718 5392 31755
rect 5471 31718 5495 31774
rect 5551 31718 5663 31774
rect 5378 31703 5392 31718
rect 5444 31703 5663 31718
rect 4663 31693 5663 31703
rect 4663 31690 4775 31693
rect 4831 31690 4855 31693
rect 4911 31690 4935 31693
rect 4991 31690 5015 31693
rect 5071 31690 5095 31693
rect 5151 31690 5175 31693
rect 5231 31690 5255 31693
rect 5311 31690 5335 31693
rect 5391 31690 5415 31693
rect 4663 31638 4666 31690
rect 4718 31638 4732 31690
rect 4850 31638 4855 31690
rect 4916 31638 4930 31690
rect 4991 31638 4996 31690
rect 5246 31638 5255 31690
rect 5312 31638 5326 31690
rect 5391 31638 5392 31690
rect 4663 31637 4775 31638
rect 4831 31637 4855 31638
rect 4911 31637 4935 31638
rect 4991 31637 5015 31638
rect 5071 31637 5095 31638
rect 5151 31637 5175 31638
rect 5231 31637 5255 31638
rect 5311 31637 5335 31638
rect 5391 31637 5415 31638
rect 5471 31637 5495 31693
rect 5551 31637 5663 31693
rect 4663 31625 5663 31637
rect 4663 31573 4666 31625
rect 4718 31573 4732 31625
rect 4784 31612 4798 31625
rect 4850 31612 4864 31625
rect 4850 31573 4855 31612
rect 4916 31573 4930 31625
rect 4982 31612 4996 31625
rect 5048 31612 5062 31625
rect 5114 31612 5128 31625
rect 5180 31612 5194 31625
rect 5246 31612 5260 31625
rect 4991 31573 4996 31612
rect 5246 31573 5255 31612
rect 5312 31573 5326 31625
rect 5378 31612 5392 31625
rect 5444 31612 5663 31625
rect 5391 31573 5392 31612
rect 4663 31560 4775 31573
rect 4831 31560 4855 31573
rect 4911 31560 4935 31573
rect 4991 31560 5015 31573
rect 5071 31560 5095 31573
rect 5151 31560 5175 31573
rect 5231 31560 5255 31573
rect 5311 31560 5335 31573
rect 5391 31560 5415 31573
rect 4663 31508 4666 31560
rect 4718 31508 4732 31560
rect 4850 31556 4855 31560
rect 4784 31531 4798 31556
rect 4850 31531 4864 31556
rect 4850 31508 4855 31531
rect 4916 31508 4930 31560
rect 4991 31556 4996 31560
rect 5246 31556 5255 31560
rect 4982 31531 4996 31556
rect 5048 31531 5062 31556
rect 5114 31531 5128 31556
rect 5180 31531 5194 31556
rect 5246 31531 5260 31556
rect 4991 31508 4996 31531
rect 5246 31508 5255 31531
rect 5312 31508 5326 31560
rect 5391 31556 5392 31560
rect 5471 31556 5495 31612
rect 5551 31556 5663 31612
rect 5378 31531 5392 31556
rect 5444 31531 5663 31556
rect 5391 31508 5392 31531
rect 4663 31495 4775 31508
rect 4831 31495 4855 31508
rect 4911 31495 4935 31508
rect 4991 31495 5015 31508
rect 5071 31495 5095 31508
rect 5151 31495 5175 31508
rect 5231 31495 5255 31508
rect 5311 31495 5335 31508
rect 5391 31495 5415 31508
rect 4663 31443 4666 31495
rect 4718 31443 4732 31495
rect 4850 31475 4855 31495
rect 4784 31450 4798 31475
rect 4850 31450 4864 31475
rect 4850 31443 4855 31450
rect 4916 31443 4930 31495
rect 4991 31475 4996 31495
rect 5246 31475 5255 31495
rect 4982 31450 4996 31475
rect 5048 31450 5062 31475
rect 5114 31450 5128 31475
rect 5180 31450 5194 31475
rect 5246 31450 5260 31475
rect 4991 31443 4996 31450
rect 5246 31443 5255 31450
rect 5312 31443 5326 31495
rect 5391 31475 5392 31495
rect 5471 31475 5495 31531
rect 5551 31475 5663 31531
rect 5378 31450 5392 31475
rect 5444 31450 5663 31475
rect 5391 31443 5392 31450
rect 4663 31430 4775 31443
rect 4831 31430 4855 31443
rect 4911 31430 4935 31443
rect 4991 31430 5015 31443
rect 5071 31430 5095 31443
rect 5151 31430 5175 31443
rect 5231 31430 5255 31443
rect 5311 31430 5335 31443
rect 5391 31430 5415 31443
rect 4663 31378 4666 31430
rect 4718 31378 4732 31430
rect 4850 31394 4855 31430
rect 4784 31378 4798 31394
rect 4850 31378 4864 31394
rect 4916 31378 4930 31430
rect 4991 31394 4996 31430
rect 5246 31394 5255 31430
rect 4982 31378 4996 31394
rect 5048 31378 5062 31394
rect 5114 31378 5128 31394
rect 5180 31378 5194 31394
rect 5246 31378 5260 31394
rect 5312 31378 5326 31430
rect 5391 31394 5392 31430
rect 5471 31394 5495 31450
rect 5551 31394 5663 31450
rect 5378 31378 5392 31394
rect 5444 31378 5663 31394
rect 4663 31369 5663 31378
rect 4663 31365 4775 31369
rect 4831 31365 4855 31369
rect 4911 31365 4935 31369
rect 4991 31365 5015 31369
rect 5071 31365 5095 31369
rect 5151 31365 5175 31369
rect 5231 31365 5255 31369
rect 5311 31365 5335 31369
rect 5391 31365 5415 31369
rect 4663 31313 4666 31365
rect 4718 31313 4732 31365
rect 4850 31313 4855 31365
rect 4916 31313 4930 31365
rect 4991 31313 4996 31365
rect 5246 31313 5255 31365
rect 5312 31313 5326 31365
rect 5391 31313 5392 31365
rect 5471 31313 5495 31369
rect 5551 31313 5663 31369
rect 4663 31300 5663 31313
rect 4663 31248 4666 31300
rect 4718 31248 4732 31300
rect 4784 31288 4798 31300
rect 4850 31288 4864 31300
rect 4850 31248 4855 31288
rect 4916 31248 4930 31300
rect 4982 31288 4996 31300
rect 5048 31288 5062 31300
rect 5114 31288 5128 31300
rect 5180 31288 5194 31300
rect 5246 31288 5260 31300
rect 4991 31248 4996 31288
rect 5246 31248 5255 31288
rect 5312 31248 5326 31300
rect 5378 31288 5392 31300
rect 5444 31288 5663 31300
rect 5391 31248 5392 31288
rect 4663 31235 4775 31248
rect 4831 31235 4855 31248
rect 4911 31235 4935 31248
rect 4991 31235 5015 31248
rect 5071 31235 5095 31248
rect 5151 31235 5175 31248
rect 5231 31235 5255 31248
rect 5311 31235 5335 31248
rect 5391 31235 5415 31248
rect 4663 31183 4666 31235
rect 4718 31183 4732 31235
rect 4850 31232 4855 31235
rect 4784 31207 4798 31232
rect 4850 31207 4864 31232
rect 4850 31183 4855 31207
rect 4916 31183 4930 31235
rect 4991 31232 4996 31235
rect 5246 31232 5255 31235
rect 4982 31207 4996 31232
rect 5048 31207 5062 31232
rect 5114 31207 5128 31232
rect 5180 31207 5194 31232
rect 5246 31207 5260 31232
rect 4991 31183 4996 31207
rect 5246 31183 5255 31207
rect 5312 31183 5326 31235
rect 5391 31232 5392 31235
rect 5471 31232 5495 31288
rect 5551 31232 5663 31288
rect 5378 31207 5392 31232
rect 5444 31207 5663 31232
rect 5391 31183 5392 31207
rect 4663 31170 4775 31183
rect 4831 31170 4855 31183
rect 4911 31170 4935 31183
rect 4991 31170 5015 31183
rect 5071 31170 5095 31183
rect 5151 31170 5175 31183
rect 5231 31170 5255 31183
rect 5311 31170 5335 31183
rect 5391 31170 5415 31183
rect 4663 31118 4666 31170
rect 4718 31118 4732 31170
rect 4850 31151 4855 31170
rect 4784 31126 4798 31151
rect 4850 31126 4864 31151
rect 4850 31118 4855 31126
rect 4916 31118 4930 31170
rect 4991 31151 4996 31170
rect 5246 31151 5255 31170
rect 4982 31126 4996 31151
rect 5048 31126 5062 31151
rect 5114 31126 5128 31151
rect 5180 31126 5194 31151
rect 5246 31126 5260 31151
rect 4991 31118 4996 31126
rect 5246 31118 5255 31126
rect 5312 31118 5326 31170
rect 5391 31151 5392 31170
rect 5471 31151 5495 31207
rect 5551 31151 5663 31207
rect 5378 31126 5392 31151
rect 5444 31126 5663 31151
rect 5391 31118 5392 31126
rect 4663 31105 4775 31118
rect 4831 31105 4855 31118
rect 4911 31105 4935 31118
rect 4991 31105 5015 31118
rect 5071 31105 5095 31118
rect 5151 31105 5175 31118
rect 5231 31105 5255 31118
rect 5311 31105 5335 31118
rect 5391 31105 5415 31118
rect 4663 31053 4666 31105
rect 4718 31053 4732 31105
rect 4850 31070 4855 31105
rect 4784 31053 4798 31070
rect 4850 31053 4864 31070
rect 4916 31053 4930 31105
rect 4991 31070 4996 31105
rect 5246 31070 5255 31105
rect 4982 31053 4996 31070
rect 5048 31053 5062 31070
rect 5114 31053 5128 31070
rect 5180 31053 5194 31070
rect 5246 31053 5260 31070
rect 5312 31053 5326 31105
rect 5391 31070 5392 31105
rect 5471 31070 5495 31126
rect 5551 31070 5663 31126
rect 5378 31053 5392 31070
rect 5444 31053 5663 31070
rect 4663 31045 5663 31053
rect 4663 31040 4775 31045
rect 4831 31040 4855 31045
rect 4911 31040 4935 31045
rect 4991 31040 5015 31045
rect 5071 31040 5095 31045
rect 5151 31040 5175 31045
rect 5231 31040 5255 31045
rect 5311 31040 5335 31045
rect 5391 31040 5415 31045
rect 4663 30988 4666 31040
rect 4718 30988 4732 31040
rect 4850 30989 4855 31040
rect 4784 30988 4798 30989
rect 4850 30988 4864 30989
rect 4916 30988 4930 31040
rect 4991 30989 4996 31040
rect 5246 30989 5255 31040
rect 4982 30988 4996 30989
rect 5048 30988 5062 30989
rect 5114 30988 5128 30989
rect 5180 30988 5194 30989
rect 5246 30988 5260 30989
rect 5312 30988 5326 31040
rect 5391 30989 5392 31040
rect 5471 30989 5495 31045
rect 5551 30989 5663 31045
rect 5378 30988 5392 30989
rect 5444 30988 5663 30989
rect 4663 30975 5663 30988
rect 4663 30923 4666 30975
rect 4718 30923 4732 30975
rect 4784 30964 4798 30975
rect 4850 30964 4864 30975
rect 4850 30923 4855 30964
rect 4916 30923 4930 30975
rect 4982 30964 4996 30975
rect 5048 30964 5062 30975
rect 5114 30964 5128 30975
rect 5180 30964 5194 30975
rect 5246 30964 5260 30975
rect 4991 30923 4996 30964
rect 5246 30923 5255 30964
rect 5312 30923 5326 30975
rect 5378 30964 5392 30975
rect 5444 30964 5663 30975
rect 5391 30923 5392 30964
rect 4663 30910 4775 30923
rect 4831 30910 4855 30923
rect 4911 30910 4935 30923
rect 4991 30910 5015 30923
rect 5071 30910 5095 30923
rect 5151 30910 5175 30923
rect 5231 30910 5255 30923
rect 5311 30910 5335 30923
rect 5391 30910 5415 30923
rect 4663 30858 4666 30910
rect 4718 30858 4732 30910
rect 4850 30908 4855 30910
rect 4784 30883 4798 30908
rect 4850 30883 4864 30908
rect 4850 30858 4855 30883
rect 4916 30858 4930 30910
rect 4991 30908 4996 30910
rect 5246 30908 5255 30910
rect 4982 30883 4996 30908
rect 5048 30883 5062 30908
rect 5114 30883 5128 30908
rect 5180 30883 5194 30908
rect 5246 30883 5260 30908
rect 4991 30858 4996 30883
rect 5246 30858 5255 30883
rect 5312 30858 5326 30910
rect 5391 30908 5392 30910
rect 5471 30908 5495 30964
rect 5551 30908 5663 30964
rect 5378 30883 5392 30908
rect 5444 30883 5663 30908
rect 5391 30858 5392 30883
rect 4663 30845 4775 30858
rect 4831 30845 4855 30858
rect 4911 30845 4935 30858
rect 4991 30845 5015 30858
rect 5071 30845 5095 30858
rect 5151 30845 5175 30858
rect 5231 30845 5255 30858
rect 5311 30845 5335 30858
rect 5391 30845 5415 30858
rect 4663 30793 4666 30845
rect 4718 30793 4732 30845
rect 4850 30827 4855 30845
rect 4784 30802 4798 30827
rect 4850 30802 4864 30827
rect 4850 30793 4855 30802
rect 4916 30793 4930 30845
rect 4991 30827 4996 30845
rect 5246 30827 5255 30845
rect 4982 30802 4996 30827
rect 5048 30802 5062 30827
rect 5114 30802 5128 30827
rect 5180 30802 5194 30827
rect 5246 30802 5260 30827
rect 4991 30793 4996 30802
rect 5246 30793 5255 30802
rect 5312 30793 5326 30845
rect 5391 30827 5392 30845
rect 5471 30827 5495 30883
rect 5551 30827 5663 30883
rect 5378 30802 5392 30827
rect 5444 30802 5663 30827
rect 5391 30793 5392 30802
rect 4663 30780 4775 30793
rect 4831 30780 4855 30793
rect 4911 30780 4935 30793
rect 4991 30780 5015 30793
rect 5071 30780 5095 30793
rect 5151 30780 5175 30793
rect 5231 30780 5255 30793
rect 5311 30780 5335 30793
rect 5391 30780 5415 30793
rect 4663 30728 4666 30780
rect 4718 30728 4732 30780
rect 4850 30746 4855 30780
rect 4784 30728 4798 30746
rect 4850 30728 4864 30746
rect 4916 30728 4930 30780
rect 4991 30746 4996 30780
rect 5246 30746 5255 30780
rect 4982 30728 4996 30746
rect 5048 30728 5062 30746
rect 5114 30728 5128 30746
rect 5180 30728 5194 30746
rect 5246 30728 5260 30746
rect 5312 30728 5326 30780
rect 5391 30746 5392 30780
rect 5471 30746 5495 30802
rect 5551 30746 5663 30802
rect 5378 30728 5392 30746
rect 5444 30728 5663 30746
rect 4663 30721 5663 30728
rect 4663 30715 4775 30721
rect 4831 30715 4855 30721
rect 4911 30715 4935 30721
rect 4991 30715 5015 30721
rect 5071 30715 5095 30721
rect 5151 30715 5175 30721
rect 5231 30715 5255 30721
rect 5311 30715 5335 30721
rect 5391 30715 5415 30721
rect 4663 30663 4666 30715
rect 4718 30663 4732 30715
rect 4850 30665 4855 30715
rect 4784 30663 4798 30665
rect 4850 30663 4864 30665
rect 4916 30663 4930 30715
rect 4991 30665 4996 30715
rect 5246 30665 5255 30715
rect 4982 30663 4996 30665
rect 5048 30663 5062 30665
rect 5114 30663 5128 30665
rect 5180 30663 5194 30665
rect 5246 30663 5260 30665
rect 5312 30663 5326 30715
rect 5391 30665 5392 30715
rect 5471 30665 5495 30721
rect 5551 30665 5663 30721
rect 5378 30663 5392 30665
rect 5444 30663 5663 30665
rect 4663 30650 5663 30663
rect 4663 30598 4666 30650
rect 4718 30598 4732 30650
rect 4784 30640 4798 30650
rect 4850 30640 4864 30650
rect 4850 30598 4855 30640
rect 4916 30598 4930 30650
rect 4982 30640 4996 30650
rect 5048 30640 5062 30650
rect 5114 30640 5128 30650
rect 5180 30640 5194 30650
rect 5246 30640 5260 30650
rect 4991 30598 4996 30640
rect 5246 30598 5255 30640
rect 5312 30598 5326 30650
rect 5378 30640 5392 30650
rect 5444 30640 5663 30650
rect 5391 30598 5392 30640
rect 4663 30585 4775 30598
rect 4831 30585 4855 30598
rect 4911 30585 4935 30598
rect 4991 30585 5015 30598
rect 5071 30585 5095 30598
rect 5151 30585 5175 30598
rect 5231 30585 5255 30598
rect 5311 30585 5335 30598
rect 5391 30585 5415 30598
rect 4663 30533 4666 30585
rect 4718 30533 4732 30585
rect 4850 30584 4855 30585
rect 4784 30559 4798 30584
rect 4850 30559 4864 30584
rect 4850 30533 4855 30559
rect 4916 30533 4930 30585
rect 4991 30584 4996 30585
rect 5246 30584 5255 30585
rect 4982 30559 4996 30584
rect 5048 30559 5062 30584
rect 5114 30559 5128 30584
rect 5180 30559 5194 30584
rect 5246 30559 5260 30584
rect 4991 30533 4996 30559
rect 5246 30533 5255 30559
rect 5312 30533 5326 30585
rect 5391 30584 5392 30585
rect 5471 30584 5495 30640
rect 5551 30584 5663 30640
rect 5378 30559 5392 30584
rect 5444 30559 5663 30584
rect 5391 30533 5392 30559
rect 4663 30520 4775 30533
rect 4831 30520 4855 30533
rect 4911 30520 4935 30533
rect 4991 30520 5015 30533
rect 5071 30520 5095 30533
rect 5151 30520 5175 30533
rect 5231 30520 5255 30533
rect 5311 30520 5335 30533
rect 5391 30520 5415 30533
rect 4663 30468 4666 30520
rect 4718 30468 4732 30520
rect 4850 30503 4855 30520
rect 4784 30478 4798 30503
rect 4850 30478 4864 30503
rect 4850 30468 4855 30478
rect 4916 30468 4930 30520
rect 4991 30503 4996 30520
rect 5246 30503 5255 30520
rect 4982 30478 4996 30503
rect 5048 30478 5062 30503
rect 5114 30478 5128 30503
rect 5180 30478 5194 30503
rect 5246 30478 5260 30503
rect 4991 30468 4996 30478
rect 5246 30468 5255 30478
rect 5312 30468 5326 30520
rect 5391 30503 5392 30520
rect 5471 30503 5495 30559
rect 5551 30503 5663 30559
rect 5378 30478 5392 30503
rect 5444 30478 5663 30503
rect 5391 30468 5392 30478
rect 4663 30455 4775 30468
rect 4831 30455 4855 30468
rect 4911 30455 4935 30468
rect 4991 30455 5015 30468
rect 5071 30455 5095 30468
rect 5151 30455 5175 30468
rect 5231 30455 5255 30468
rect 5311 30455 5335 30468
rect 5391 30455 5415 30468
rect 4663 30403 4666 30455
rect 4718 30403 4732 30455
rect 4850 30422 4855 30455
rect 4784 30403 4798 30422
rect 4850 30403 4864 30422
rect 4916 30403 4930 30455
rect 4991 30422 4996 30455
rect 5246 30422 5255 30455
rect 4982 30403 4996 30422
rect 5048 30403 5062 30422
rect 5114 30403 5128 30422
rect 5180 30403 5194 30422
rect 5246 30403 5260 30422
rect 5312 30403 5326 30455
rect 5391 30422 5392 30455
rect 5471 30422 5495 30478
rect 5551 30422 5663 30478
rect 5378 30403 5392 30422
rect 5444 30403 5663 30422
rect 4663 30397 5663 30403
rect 4663 30390 4775 30397
rect 4831 30390 4855 30397
rect 4911 30390 4935 30397
rect 4991 30390 5015 30397
rect 5071 30390 5095 30397
rect 5151 30390 5175 30397
rect 5231 30390 5255 30397
rect 5311 30390 5335 30397
rect 5391 30390 5415 30397
rect 4663 30338 4666 30390
rect 4718 30338 4732 30390
rect 4850 30341 4855 30390
rect 4784 30338 4798 30341
rect 4850 30338 4864 30341
rect 4916 30338 4930 30390
rect 4991 30341 4996 30390
rect 5246 30341 5255 30390
rect 4982 30338 4996 30341
rect 5048 30338 5062 30341
rect 5114 30338 5128 30341
rect 5180 30338 5194 30341
rect 5246 30338 5260 30341
rect 5312 30338 5326 30390
rect 5391 30341 5392 30390
rect 5471 30341 5495 30397
rect 5551 30341 5663 30397
rect 5378 30338 5392 30341
rect 5444 30338 5663 30341
rect 4663 30332 5663 30338
rect 5864 30469 8229 30521
rect 8281 30469 8293 30521
rect 8345 30469 8351 30521
tri 5830 30134 5864 30168 se
rect 5864 30134 5916 30469
tri 5916 30435 5950 30469 nw
rect 4863 30082 4869 30134
rect 4921 30082 4946 30134
rect 4998 30082 5022 30134
rect 5074 30082 5098 30134
rect 5150 30082 5174 30134
rect 5226 30082 5916 30134
rect 6188 30128 9619 30134
rect 6188 30099 9567 30128
rect 6240 30082 9567 30099
rect 6240 30076 6268 30082
tri 6268 30076 6274 30082 nw
tri 9533 30076 9539 30082 ne
rect 9539 30076 9567 30082
rect 6240 30064 6256 30076
tri 6256 30064 6268 30076 nw
tri 9539 30064 9551 30076 ne
rect 9551 30064 9619 30076
rect 6240 30054 6246 30064
tri 6246 30054 6256 30064 nw
tri 9551 30054 9561 30064 ne
rect 9561 30054 9567 30064
tri 6240 30048 6246 30054 nw
rect 6188 30035 6240 30047
rect 6348 30002 6354 30054
rect 6406 30002 6418 30054
rect 6470 30048 9508 30054
tri 9561 30048 9567 30054 ne
rect 6470 30002 9456 30048
tri 9422 29996 9428 30002 ne
rect 9428 29996 9456 30002
rect 9567 30006 9619 30012
tri 9428 29984 9440 29996 ne
rect 9440 29984 9508 29996
rect 6188 29977 6240 29983
tri 9440 29977 9447 29984 ne
rect 9447 29977 9456 29984
tri 9447 29974 9450 29977 ne
rect 9450 29974 9456 29977
rect 6483 29922 6489 29974
rect 6541 29922 6553 29974
rect 6605 29968 9352 29974
tri 9450 29968 9456 29974 ne
rect 6605 29922 9300 29968
tri 9266 29916 9272 29922 ne
rect 9272 29916 9300 29922
rect 9456 29926 9508 29932
tri 9272 29911 9277 29916 ne
rect 9277 29911 9352 29916
rect 3550 29905 5663 29911
rect 3602 29875 5261 29905
rect 5313 29875 5663 29905
tri 9277 29904 9284 29911 ne
rect 9284 29904 9352 29911
tri 9284 29888 9300 29904 ne
rect 3602 29853 4672 29875
rect 3550 29841 4672 29853
rect 3602 29819 4672 29841
rect 4728 29819 4757 29875
rect 4813 29819 4842 29875
rect 4898 29819 4926 29875
rect 4982 29819 5010 29875
rect 5066 29819 5094 29875
rect 5150 29819 5178 29875
rect 5234 29853 5261 29875
rect 5234 29841 5262 29853
rect 5234 29819 5261 29841
rect 5318 29819 5346 29875
rect 5402 29819 5430 29875
rect 5486 29819 5514 29875
rect 5570 29819 5598 29875
rect 5654 29819 5663 29875
rect 9300 29846 9352 29852
rect 3602 29789 5261 29819
rect 5313 29789 5663 29819
rect 3550 29783 5663 29789
tri 8894 29613 8928 29647 ne
rect 2627 29435 2633 29487
rect 2685 29435 2730 29487
rect 2782 29481 5313 29487
rect 2782 29435 3550 29481
rect 2627 29429 3550 29435
rect 3602 29429 5261 29481
rect 2627 29417 5313 29429
rect 2627 29411 3550 29417
rect 2627 29359 2633 29411
rect 2685 29359 2730 29411
rect 2782 29365 3550 29411
rect 3602 29365 5261 29417
rect 2782 29359 5313 29365
tri 4167 29325 4201 29359 ne
rect 4201 29147 4329 29359
tri 4329 29325 4363 29359 nw
tri 4704 29325 4738 29359 ne
rect 4201 29095 4207 29147
rect 4259 29095 4271 29147
rect 4323 29095 4329 29147
rect 4738 29147 4866 29359
tri 4866 29325 4900 29359 nw
rect 4738 29095 4744 29147
rect 4796 29095 4808 29147
rect 4860 29095 4866 29147
rect 2288 28957 2294 29009
rect 2346 28957 2391 29009
rect 2443 28957 4380 29009
rect 4432 28957 4444 29009
rect 4496 28957 4502 29009
rect 3550 28921 5663 28927
rect 3602 28891 5261 28921
rect 5313 28891 5663 28921
rect 3602 28869 4672 28891
rect 3550 28857 4672 28869
rect 3602 28835 4672 28857
rect 4728 28835 4757 28891
rect 4813 28835 4842 28891
rect 4898 28835 4926 28891
rect 4982 28835 5010 28891
rect 5066 28835 5094 28891
rect 5150 28835 5178 28891
rect 5234 28869 5261 28891
rect 5234 28857 5262 28869
rect 5234 28835 5261 28857
rect 5318 28835 5346 28891
rect 5402 28835 5430 28891
rect 5486 28835 5514 28891
rect 5570 28835 5598 28891
rect 5654 28835 5663 28891
rect 3602 28805 5261 28835
rect 5313 28805 5663 28835
rect 3550 28799 5663 28805
rect 4663 28443 4672 28445
rect 4728 28443 4757 28445
rect 4813 28443 4842 28445
rect 4898 28443 4926 28445
rect 4982 28443 5010 28445
rect 5066 28443 5094 28445
rect 5150 28443 5178 28445
rect 5234 28443 5262 28445
rect 5318 28443 5346 28445
rect 5402 28443 5430 28445
rect 5486 28443 5514 28445
rect 5570 28443 5598 28445
rect 5654 28443 5663 28445
rect 4663 28391 4669 28443
rect 4728 28391 4736 28443
rect 4922 28391 4926 28443
rect 4989 28391 5004 28443
rect 5066 28391 5071 28443
rect 5257 28391 5262 28443
rect 5324 28391 5339 28443
rect 5402 28391 5406 28443
rect 5591 28391 5598 28443
rect 5657 28391 5663 28443
rect 4663 28389 4672 28391
rect 4728 28389 4757 28391
rect 4813 28389 4842 28391
rect 4898 28389 4926 28391
rect 4982 28389 5010 28391
rect 5066 28389 5094 28391
rect 5150 28389 5178 28391
rect 5234 28389 5262 28391
rect 5318 28389 5346 28391
rect 5402 28389 5430 28391
rect 5486 28389 5514 28391
rect 5570 28389 5598 28391
rect 5654 28389 5663 28391
rect 3703 28183 3712 28185
rect 3768 28183 3793 28185
rect 3849 28183 3874 28185
rect 3930 28183 3955 28185
rect 4011 28183 4036 28185
rect 4092 28183 4117 28185
rect 4173 28183 4198 28185
rect 4254 28183 4278 28185
rect 4334 28183 4358 28185
rect 4414 28183 4438 28185
rect 4494 28183 4503 28185
rect 3703 28131 3709 28183
rect 3768 28131 3776 28183
rect 4029 28131 4036 28183
rect 4096 28131 4111 28183
rect 4173 28131 4178 28183
rect 4431 28131 4438 28183
rect 4497 28131 4503 28183
rect 3703 28129 3712 28131
rect 3768 28129 3793 28131
rect 3849 28129 3874 28131
rect 3930 28129 3955 28131
rect 4011 28129 4036 28131
rect 4092 28129 4117 28131
rect 4173 28129 4198 28131
rect 4254 28129 4278 28131
rect 4334 28129 4358 28131
rect 4414 28129 4438 28131
rect 4494 28129 4503 28131
rect 1187 26202 4441 26208
rect 1239 26156 4441 26202
rect 4493 26156 4508 26208
rect 4560 26156 4575 26208
rect 4627 26156 4642 26208
rect 4694 26156 4709 26208
rect 4761 26156 4776 26208
rect 4828 26156 4843 26208
rect 4895 26156 4910 26208
rect 4962 26156 4977 26208
rect 5029 26156 5044 26208
rect 5096 26156 5102 26208
rect 1187 26138 1239 26150
tri 1239 26122 1273 26156 nw
rect 1187 26080 1239 26086
rect 908 25807 5488 25813
rect 908 25755 932 25807
rect 984 25755 4500 25807
rect 4552 25755 4812 25807
rect 4864 25755 5124 25807
rect 5176 25755 5436 25807
rect 908 25743 5488 25755
rect 908 25691 932 25743
rect 984 25691 4500 25743
rect 4552 25691 4812 25743
rect 4864 25691 5124 25743
rect 5176 25691 5436 25743
rect 908 25685 5488 25691
rect 1187 25601 1239 25607
tri 1239 25559 1245 25565 sw
rect 1239 25549 1245 25559
rect 1187 25537 1245 25549
rect 1239 25531 1245 25537
tri 1245 25531 1273 25559 sw
rect 1239 25485 2826 25531
rect 1187 25479 2826 25485
rect 2878 25479 2890 25531
rect 2942 25479 2948 25531
rect 3524 25507 3530 25559
rect 3582 25507 3596 25559
rect 3648 25558 3970 25559
rect 3648 25507 3776 25558
rect 3524 25506 3776 25507
rect 3828 25506 3844 25558
rect 3896 25506 3912 25558
rect 3964 25506 3970 25558
rect 1583 25449 5989 25451
rect 1583 25393 1592 25449
rect 1648 25393 1673 25449
rect 1729 25393 1754 25449
rect 1810 25393 1835 25449
rect 1891 25393 1916 25449
rect 1972 25393 1997 25449
rect 2053 25393 2078 25449
rect 1583 25369 2078 25393
rect 1583 25313 1592 25369
rect 1648 25313 1673 25369
rect 1729 25313 1754 25369
rect 1810 25313 1835 25369
rect 1891 25313 1916 25369
rect 1972 25313 1997 25369
rect 2053 25313 2078 25369
rect 1583 25289 2078 25313
rect 1583 25233 1592 25289
rect 1648 25233 1673 25289
rect 1729 25233 1754 25289
rect 1810 25233 1835 25289
rect 1891 25233 1916 25289
rect 1972 25233 1997 25289
rect 2053 25233 2078 25289
rect 1583 25209 2078 25233
rect 1583 25153 1592 25209
rect 1648 25153 1673 25209
rect 1729 25153 1754 25209
rect 1810 25153 1835 25209
rect 1891 25153 1916 25209
rect 1972 25153 1997 25209
rect 2053 25153 2078 25209
rect 2374 25445 5989 25449
rect 2374 25393 3999 25445
rect 4051 25393 4344 25445
rect 4396 25393 4656 25445
rect 4708 25393 4968 25445
rect 5020 25393 5280 25445
rect 5332 25393 5592 25445
rect 5644 25393 5937 25445
rect 2374 25367 5989 25393
rect 2374 25315 3999 25367
rect 4051 25315 4344 25367
rect 4396 25315 4656 25367
rect 4708 25315 4968 25367
rect 5020 25315 5280 25367
rect 5332 25315 5592 25367
rect 5644 25315 5937 25367
rect 2374 25288 5989 25315
rect 2374 25236 3999 25288
rect 4051 25236 4344 25288
rect 4396 25236 4656 25288
rect 4708 25236 4968 25288
rect 5020 25236 5280 25288
rect 5332 25236 5592 25288
rect 5644 25236 5937 25288
rect 2374 25209 5989 25236
rect 2374 25157 3999 25209
rect 4051 25157 4344 25209
rect 4396 25157 4656 25209
rect 4708 25157 4968 25209
rect 5020 25157 5280 25209
rect 5332 25157 5592 25209
rect 5644 25157 5937 25209
rect 2374 25153 5989 25157
rect 1583 25151 5989 25153
rect 3703 23844 5901 23850
rect 3703 23814 4451 23844
rect 4503 23838 5849 23844
rect 3703 23758 3712 23814
rect 3768 23758 3793 23814
rect 3849 23758 3874 23814
rect 3930 23758 3955 23814
rect 4011 23758 4036 23814
rect 4092 23758 4117 23814
rect 4173 23758 4198 23814
rect 4254 23758 4278 23814
rect 4334 23758 4358 23814
rect 4414 23758 4438 23814
rect 4503 23792 4646 23838
rect 4494 23786 4646 23792
rect 4698 23786 4722 23838
rect 4774 23786 4797 23838
rect 4849 23786 5055 23838
rect 4494 23780 5055 23786
rect 4503 23774 5055 23780
rect 3703 23728 4451 23758
rect 4503 23728 4646 23774
rect 3703 23722 4646 23728
rect 4698 23722 4722 23774
rect 4774 23722 4797 23774
rect 4849 23722 5055 23774
rect 5171 23722 5310 23838
rect 5426 23792 5849 23838
rect 5426 23780 5901 23792
rect 5426 23728 5849 23780
rect 5426 23722 5901 23728
rect 2288 22478 2294 22530
rect 2346 22478 2391 22530
rect 2443 22524 5495 22530
rect 2443 22478 4879 22524
rect 2288 22472 4879 22478
rect 4931 22472 5443 22524
rect 2288 22460 5495 22472
rect 2288 22454 4879 22460
rect 2288 22402 2294 22454
rect 2346 22402 2391 22454
rect 2443 22408 4879 22454
rect 4931 22408 5443 22460
rect 2443 22402 5495 22408
rect 7499 22285 7624 22337
rect 7676 22285 7688 22337
rect 7740 22285 9230 22337
rect 9282 22285 9294 22337
rect 9346 22285 9352 22337
rect 7346 22205 7492 22257
rect 7544 22205 7556 22257
rect 7608 22205 9386 22257
rect 9438 22205 9450 22257
rect 9502 22205 9508 22257
rect 2996 22185 3048 22191
rect 2996 22125 3048 22133
tri 3048 22125 3072 22149 sw
rect 7306 22125 7312 22177
rect 7364 22125 7376 22177
rect 7428 22171 9619 22177
rect 7428 22125 9567 22171
rect 2996 22121 3072 22125
rect 3048 22119 3072 22121
tri 3072 22119 3078 22125 sw
tri 9533 22119 9539 22125 ne
rect 9539 22119 9567 22125
rect 3048 22115 3078 22119
tri 3078 22115 3082 22119 sw
tri 9539 22115 9543 22119 ne
rect 9543 22115 9619 22119
rect 3048 22069 4686 22115
rect 2996 22063 4686 22069
rect 4738 22063 4750 22115
rect 4802 22063 4808 22115
tri 9543 22107 9551 22115 ne
rect 9551 22107 9619 22115
tri 9551 22091 9567 22107 ne
rect 9567 22049 9619 22055
rect 2627 21640 2633 21692
rect 2685 21640 2730 21692
rect 2782 21686 5239 21692
rect 2782 21640 5187 21686
rect 2627 21634 5187 21640
rect 2627 21622 5239 21634
rect 2627 21616 5187 21622
rect 2627 21564 2633 21616
rect 2685 21564 2730 21616
rect 2782 21570 5187 21616
rect 2782 21564 5239 21570
rect 3703 20419 4646 20449
rect 3703 20363 3712 20419
rect 3768 20363 3793 20419
rect 3849 20363 3874 20419
rect 3930 20363 3955 20419
rect 4011 20363 4036 20419
rect 4092 20363 4117 20419
rect 4173 20363 4198 20419
rect 4254 20363 4278 20419
rect 4334 20363 4358 20419
rect 4414 20363 4438 20419
rect 4494 20397 4646 20419
rect 4698 20397 4722 20449
rect 4774 20397 4797 20449
rect 4849 20397 4855 20449
rect 4494 20385 4855 20397
rect 4494 20363 4646 20385
rect 3703 20333 4646 20363
rect 4698 20333 4722 20385
rect 4774 20333 4797 20385
rect 4849 20333 4855 20385
rect 5699 20253 8351 20259
rect 5751 20201 8223 20253
rect 8275 20201 8299 20253
rect 5699 20189 8351 20201
rect 5751 20137 8223 20189
rect 8275 20137 8299 20189
rect 5699 20131 8351 20137
rect 3703 20024 4472 20054
rect 3703 19968 3712 20024
rect 3768 19968 3793 20024
rect 3849 19968 3874 20024
rect 3930 19968 3955 20024
rect 4011 19968 4036 20024
rect 4092 19968 4117 20024
rect 4173 19968 4198 20024
rect 4254 19968 4278 20024
rect 4334 19968 4358 20024
rect 4414 19968 4438 20024
rect 3703 19938 4472 19968
rect 4588 19938 4594 20054
rect 4727 19971 4733 20023
rect 4785 19971 4797 20023
rect 4849 19971 8799 20023
rect 8851 19971 8863 20023
rect 8915 19971 8921 20023
rect 4893 19886 4945 19892
tri 4877 19834 4893 19850 se
tri 4865 19822 4877 19834 se
rect 4877 19822 4945 19834
tri 4859 19816 4865 19822 se
rect 4865 19816 4893 19822
rect 2996 19764 3002 19816
rect 3054 19764 3066 19816
rect 3118 19770 4893 19816
rect 3118 19764 4945 19770
rect 2627 19654 2633 19706
rect 2685 19654 2730 19706
rect 2782 19700 5513 19706
rect 2782 19654 5461 19700
rect 2627 19648 5461 19654
rect 2627 19636 5513 19648
rect 2627 19630 5461 19636
rect 2627 19578 2633 19630
rect 2685 19578 2730 19630
rect 2782 19584 5461 19630
rect 2782 19578 5513 19584
rect 2288 19219 2294 19271
rect 2346 19219 2391 19271
rect 2443 19219 5080 19271
rect 5132 19219 5152 19271
rect 2288 19207 5152 19219
rect 2288 19155 2294 19207
rect 2346 19155 2391 19207
rect 2443 19155 5080 19207
rect 5132 19155 5152 19207
rect 4987 18996 5039 19002
rect 4987 18932 5039 18944
rect 4987 18874 5039 18880
rect 5247 18816 5299 18822
rect 5247 18752 5299 18764
rect 2627 18694 2633 18746
rect 2685 18694 2730 18746
rect 2782 18700 5247 18746
rect 2782 18694 5299 18700
rect 2996 18473 3048 18479
rect 2996 18409 3048 18421
rect 2996 18202 3048 18357
rect 3703 18298 3712 18300
rect 3768 18298 3793 18300
rect 3849 18298 3874 18300
rect 3930 18298 3955 18300
rect 4011 18298 4036 18300
rect 4092 18298 4117 18300
rect 4173 18298 4198 18300
rect 4254 18298 4278 18300
rect 4334 18298 4358 18300
rect 4414 18298 4438 18300
rect 4494 18298 4503 18300
rect 3703 18246 3709 18298
rect 3768 18246 3776 18298
rect 4029 18246 4036 18298
rect 4096 18246 4111 18298
rect 4173 18246 4178 18298
rect 4431 18246 4438 18298
rect 4497 18246 4503 18298
rect 3703 18244 3712 18246
rect 3768 18244 3793 18246
rect 3849 18244 3874 18246
rect 3930 18244 3955 18246
rect 4011 18244 4036 18246
rect 4092 18244 4117 18246
rect 4173 18244 4198 18246
rect 4254 18244 4278 18246
rect 4334 18244 4358 18246
rect 4414 18244 4438 18246
rect 4494 18244 4503 18246
rect 2996 18138 3048 18150
rect 2996 18080 3048 18086
rect 2993 17925 3183 17931
rect 2993 17873 3076 17925
rect 3128 17879 3183 17925
rect 3235 17879 3254 17931
rect 3306 17879 3324 17931
rect 3376 17925 6037 17931
rect 3376 17879 3946 17925
rect 3128 17873 3946 17879
rect 3998 17873 4215 17925
rect 4267 17873 4527 17925
rect 4579 17895 4839 17925
rect 4891 17895 5151 17925
rect 5203 17895 5462 17925
rect 5514 17895 5832 17925
rect 4579 17873 4672 17895
rect 2993 17861 4672 17873
rect 2993 17809 3076 17861
rect 3128 17855 3946 17861
rect 3128 17809 3183 17855
rect 2993 17803 3183 17809
rect 3235 17803 3254 17855
rect 3306 17803 3324 17855
rect 3376 17809 3946 17855
rect 3998 17809 4215 17861
rect 4267 17809 4527 17861
rect 4579 17839 4672 17861
rect 4728 17839 4757 17895
rect 4813 17873 4839 17895
rect 4813 17861 4842 17873
rect 4813 17839 4839 17861
rect 4898 17839 4926 17895
rect 4982 17839 5010 17895
rect 5066 17839 5094 17895
rect 5150 17873 5151 17895
rect 5150 17861 5178 17873
rect 5150 17839 5151 17861
rect 5234 17839 5262 17895
rect 5318 17839 5346 17895
rect 5402 17839 5430 17895
rect 5486 17861 5514 17873
rect 5570 17839 5598 17895
rect 5654 17873 5832 17895
rect 5884 17873 6037 17925
rect 5654 17861 6037 17873
rect 5654 17839 5832 17861
rect 4579 17809 4839 17839
rect 4891 17809 5151 17839
rect 5203 17809 5462 17839
rect 5514 17809 5832 17839
rect 5884 17809 6037 17861
rect 3376 17803 6037 17809
rect 2627 17723 2633 17775
rect 2685 17723 2730 17775
rect 2782 17769 4734 17775
rect 2782 17723 4371 17769
rect 2627 17717 4371 17723
rect 4423 17717 4682 17769
rect 2627 17705 4734 17717
rect 2627 17699 4371 17705
rect 2627 17647 2633 17699
rect 2685 17647 2730 17699
rect 2782 17653 4371 17699
rect 4423 17653 4682 17705
rect 2782 17647 4734 17653
rect 2288 17567 2294 17619
rect 2346 17567 2391 17619
rect 2443 17613 5359 17619
rect 2443 17567 3435 17613
rect 2288 17561 3435 17567
rect 3487 17561 4995 17613
rect 5047 17561 5307 17613
rect 2288 17549 5359 17561
rect 2288 17543 3435 17549
rect 2288 17491 2294 17543
rect 2346 17491 2391 17543
rect 2443 17497 3435 17543
rect 3487 17497 4995 17549
rect 5047 17497 5307 17549
rect 2443 17491 5359 17497
rect 3620 17461 8918 17463
rect 2996 17453 3592 17459
rect 3048 17407 3540 17453
rect 3048 17403 3078 17407
tri 3078 17403 3082 17407 nw
tri 3506 17403 3510 17407 ne
rect 3510 17403 3540 17407
rect 3048 17401 3076 17403
tri 3076 17401 3078 17403 nw
tri 3510 17401 3512 17403 ne
rect 3512 17401 3540 17403
rect 2996 17393 3068 17401
tri 3068 17393 3076 17401 nw
tri 3512 17393 3520 17401 ne
rect 3520 17393 3592 17401
rect 2996 17389 3064 17393
tri 3064 17389 3068 17393 nw
tri 3520 17389 3524 17393 ne
rect 3524 17389 3592 17393
tri 3048 17373 3064 17389 nw
tri 3524 17373 3540 17389 ne
rect 2996 17331 3048 17337
rect 3540 17331 3592 17337
rect 3620 17457 8799 17461
rect 3672 17409 8799 17457
rect 8851 17409 8863 17461
rect 8915 17409 8921 17461
rect 3672 17405 8918 17409
rect 3620 17403 8918 17405
rect 3620 17393 3672 17403
tri 3672 17369 3706 17403 nw
rect 3620 17335 3672 17341
rect 1187 16824 1193 16876
rect 1245 16824 1257 16876
rect 1309 16824 4383 16876
rect 4435 16824 4447 16876
rect 4499 16824 4505 16876
rect 908 16786 5056 16792
rect 960 16740 5056 16786
rect 5108 16740 5120 16792
rect 5172 16740 5178 16792
rect 908 16720 960 16734
tri 960 16706 994 16740 nw
rect 908 16654 960 16668
rect 4180 16652 4232 16658
rect 908 16600 960 16602
tri 960 16600 976 16616 sw
tri 4164 16600 4180 16616 se
rect 908 16588 976 16600
tri 976 16588 988 16600 sw
tri 4152 16588 4164 16600 se
rect 4164 16588 4232 16600
rect 960 16582 988 16588
tri 988 16582 994 16588 sw
tri 4146 16582 4152 16588 se
rect 4152 16582 4180 16588
rect 960 16536 4180 16582
rect 908 16530 4232 16536
rect 1187 16368 1193 16420
rect 1245 16368 1257 16420
rect 1309 16368 4884 16420
rect 4936 16368 4948 16420
rect 5000 16368 5007 16420
rect 2996 16006 3234 16012
rect 3048 15960 3234 16006
rect 3286 15960 3298 16012
rect 3350 15960 3356 16012
rect 2996 15942 3048 15954
tri 3048 15926 3082 15960 nw
rect 2996 15884 3048 15890
rect 3076 15872 6519 15878
rect 3128 15820 6464 15872
rect 6516 15820 6519 15872
rect 3076 15808 6519 15820
rect 3128 15756 6464 15808
rect 6516 15756 6519 15808
rect 3076 15750 6519 15756
rect 4663 14811 4672 14867
rect 4728 14811 4757 14867
rect 4813 14811 4842 14867
rect 4898 14811 4926 14867
rect 4982 14811 5010 14867
rect 5066 14811 5094 14867
rect 5150 14811 5178 14867
rect 5234 14811 5262 14867
rect 5318 14811 5346 14867
rect 5402 14811 5430 14867
rect 5486 14811 5514 14867
rect 5570 14811 5598 14867
rect 5654 14861 6516 14867
rect 5654 14811 5837 14861
rect 4663 14809 5837 14811
rect 5889 14809 6211 14861
rect 6263 14809 6295 14861
rect 6347 14809 6379 14861
rect 6431 14809 6463 14861
rect 6515 14809 6516 14861
rect 4663 14793 6516 14809
rect 4663 14741 5837 14793
rect 5889 14741 6211 14793
rect 6263 14741 6295 14793
rect 6347 14741 6379 14793
rect 6431 14741 6463 14793
rect 6515 14741 6516 14793
rect 4663 14725 6516 14741
rect 4663 14723 5837 14725
rect 4663 14667 4672 14723
rect 4728 14667 4757 14723
rect 4813 14667 4842 14723
rect 4898 14667 4926 14723
rect 4982 14667 5010 14723
rect 5066 14667 5094 14723
rect 5150 14667 5178 14723
rect 5234 14667 5262 14723
rect 5318 14667 5346 14723
rect 5402 14667 5430 14723
rect 5486 14667 5514 14723
rect 5570 14667 5598 14723
rect 5654 14673 5837 14723
rect 5889 14673 6211 14725
rect 6263 14673 6295 14725
rect 6347 14673 6379 14725
rect 6431 14673 6463 14725
rect 6515 14673 6516 14725
rect 5654 14667 6516 14673
<< via2 >>
rect 4775 39143 4784 39192
rect 4784 39143 4798 39192
rect 4798 39143 4850 39192
rect 4850 39143 4864 39192
rect 4864 39143 4916 39192
rect 4916 39143 4930 39192
rect 4930 39143 4982 39192
rect 4982 39143 4996 39192
rect 4996 39143 5048 39192
rect 5048 39143 5062 39192
rect 5062 39143 5114 39192
rect 5114 39143 5128 39192
rect 5128 39143 5180 39192
rect 5180 39143 5194 39192
rect 5194 39143 5246 39192
rect 5246 39143 5260 39192
rect 5260 39143 5312 39192
rect 5312 39143 5326 39192
rect 5326 39143 5378 39192
rect 5378 39143 5392 39192
rect 5392 39143 5444 39192
rect 5444 39143 5551 39192
rect 4775 39131 5551 39143
rect 4775 39079 4784 39131
rect 4784 39079 4798 39131
rect 4798 39079 4850 39131
rect 4850 39079 4864 39131
rect 4864 39079 4916 39131
rect 4916 39079 4930 39131
rect 4930 39079 4982 39131
rect 4982 39079 4996 39131
rect 4996 39079 5048 39131
rect 5048 39079 5062 39131
rect 5062 39079 5114 39131
rect 5114 39079 5128 39131
rect 5128 39079 5180 39131
rect 5180 39079 5194 39131
rect 5194 39079 5246 39131
rect 5246 39079 5260 39131
rect 5260 39079 5312 39131
rect 5312 39079 5326 39131
rect 5326 39079 5378 39131
rect 5378 39079 5392 39131
rect 5392 39079 5444 39131
rect 5444 39079 5551 39131
rect 4775 39067 5551 39079
rect 4775 39015 4784 39067
rect 4784 39015 4798 39067
rect 4798 39015 4850 39067
rect 4850 39015 4864 39067
rect 4864 39015 4916 39067
rect 4916 39015 4930 39067
rect 4930 39015 4982 39067
rect 4982 39015 4996 39067
rect 4996 39015 5048 39067
rect 5048 39015 5062 39067
rect 5062 39015 5114 39067
rect 5114 39015 5128 39067
rect 5128 39015 5180 39067
rect 5180 39015 5194 39067
rect 5194 39015 5246 39067
rect 5246 39015 5260 39067
rect 5260 39015 5312 39067
rect 5312 39015 5326 39067
rect 5326 39015 5378 39067
rect 5378 39015 5392 39067
rect 5392 39015 5444 39067
rect 5444 39015 5551 39067
rect 4775 39003 5551 39015
rect 4775 38951 4784 39003
rect 4784 38951 4798 39003
rect 4798 38951 4850 39003
rect 4850 38951 4864 39003
rect 4864 38951 4916 39003
rect 4916 38951 4930 39003
rect 4930 38951 4982 39003
rect 4982 38951 4996 39003
rect 4996 38951 5048 39003
rect 5048 38951 5062 39003
rect 5062 38951 5114 39003
rect 5114 38951 5128 39003
rect 5128 38951 5180 39003
rect 5180 38951 5194 39003
rect 5194 38951 5246 39003
rect 5246 38951 5260 39003
rect 5260 38951 5312 39003
rect 5312 38951 5326 39003
rect 5326 38951 5378 39003
rect 5378 38951 5392 39003
rect 5392 38951 5444 39003
rect 5444 38951 5551 39003
rect 4775 38939 5551 38951
rect 4775 38887 4784 38939
rect 4784 38887 4798 38939
rect 4798 38887 4850 38939
rect 4850 38887 4864 38939
rect 4864 38887 4916 38939
rect 4916 38887 4930 38939
rect 4930 38887 4982 38939
rect 4982 38887 4996 38939
rect 4996 38887 5048 38939
rect 5048 38887 5062 38939
rect 5062 38887 5114 38939
rect 5114 38887 5128 38939
rect 5128 38887 5180 38939
rect 5180 38887 5194 38939
rect 5194 38887 5246 38939
rect 5246 38887 5260 38939
rect 5260 38887 5312 38939
rect 5312 38887 5326 38939
rect 5326 38887 5378 38939
rect 5378 38887 5392 38939
rect 5392 38887 5444 38939
rect 5444 38887 5551 38939
rect 4775 38875 5551 38887
rect 4775 38823 4784 38875
rect 4784 38823 4798 38875
rect 4798 38823 4850 38875
rect 4850 38823 4864 38875
rect 4864 38823 4916 38875
rect 4916 38823 4930 38875
rect 4930 38823 4982 38875
rect 4982 38823 4996 38875
rect 4996 38823 5048 38875
rect 5048 38823 5062 38875
rect 5062 38823 5114 38875
rect 5114 38823 5128 38875
rect 5128 38823 5180 38875
rect 5180 38823 5194 38875
rect 5194 38823 5246 38875
rect 5246 38823 5260 38875
rect 5260 38823 5312 38875
rect 5312 38823 5326 38875
rect 5326 38823 5378 38875
rect 5378 38823 5392 38875
rect 5392 38823 5444 38875
rect 5444 38823 5551 38875
rect 4775 38811 5551 38823
rect 4775 38759 4784 38811
rect 4784 38759 4798 38811
rect 4798 38759 4850 38811
rect 4850 38759 4864 38811
rect 4864 38759 4916 38811
rect 4916 38759 4930 38811
rect 4930 38759 4982 38811
rect 4982 38759 4996 38811
rect 4996 38759 5048 38811
rect 5048 38759 5062 38811
rect 5062 38759 5114 38811
rect 5114 38759 5128 38811
rect 5128 38759 5180 38811
rect 5180 38759 5194 38811
rect 5194 38759 5246 38811
rect 5246 38759 5260 38811
rect 5260 38759 5312 38811
rect 5312 38759 5326 38811
rect 5326 38759 5378 38811
rect 5378 38759 5392 38811
rect 5392 38759 5444 38811
rect 5444 38759 5551 38811
rect 4775 38747 5551 38759
rect 4775 38695 4784 38747
rect 4784 38695 4798 38747
rect 4798 38695 4850 38747
rect 4850 38695 4864 38747
rect 4864 38695 4916 38747
rect 4916 38695 4930 38747
rect 4930 38695 4982 38747
rect 4982 38695 4996 38747
rect 4996 38695 5048 38747
rect 5048 38695 5062 38747
rect 5062 38695 5114 38747
rect 5114 38695 5128 38747
rect 5128 38695 5180 38747
rect 5180 38695 5194 38747
rect 5194 38695 5246 38747
rect 5246 38695 5260 38747
rect 5260 38695 5312 38747
rect 5312 38695 5326 38747
rect 5326 38695 5378 38747
rect 5378 38695 5392 38747
rect 5392 38695 5444 38747
rect 5444 38695 5551 38747
rect 4775 38683 5551 38695
rect 4775 38631 4784 38683
rect 4784 38631 4798 38683
rect 4798 38631 4850 38683
rect 4850 38631 4864 38683
rect 4864 38631 4916 38683
rect 4916 38631 4930 38683
rect 4930 38631 4982 38683
rect 4982 38631 4996 38683
rect 4996 38631 5048 38683
rect 5048 38631 5062 38683
rect 5062 38631 5114 38683
rect 5114 38631 5128 38683
rect 5128 38631 5180 38683
rect 5180 38631 5194 38683
rect 5194 38631 5246 38683
rect 5246 38631 5260 38683
rect 5260 38631 5312 38683
rect 5312 38631 5326 38683
rect 5326 38631 5378 38683
rect 5378 38631 5392 38683
rect 5392 38631 5444 38683
rect 5444 38631 5551 38683
rect 4775 38619 5551 38631
rect 4775 38567 4784 38619
rect 4784 38567 4798 38619
rect 4798 38567 4850 38619
rect 4850 38567 4864 38619
rect 4864 38567 4916 38619
rect 4916 38567 4930 38619
rect 4930 38567 4982 38619
rect 4982 38567 4996 38619
rect 4996 38567 5048 38619
rect 5048 38567 5062 38619
rect 5062 38567 5114 38619
rect 5114 38567 5128 38619
rect 5128 38567 5180 38619
rect 5180 38567 5194 38619
rect 5194 38567 5246 38619
rect 5246 38567 5260 38619
rect 5260 38567 5312 38619
rect 5312 38567 5326 38619
rect 5326 38567 5378 38619
rect 5378 38567 5392 38619
rect 5392 38567 5444 38619
rect 5444 38567 5551 38619
rect 4775 38555 5551 38567
rect 4775 38503 4784 38555
rect 4784 38503 4798 38555
rect 4798 38503 4850 38555
rect 4850 38503 4864 38555
rect 4864 38503 4916 38555
rect 4916 38503 4930 38555
rect 4930 38503 4982 38555
rect 4982 38503 4996 38555
rect 4996 38503 5048 38555
rect 5048 38503 5062 38555
rect 5062 38503 5114 38555
rect 5114 38503 5128 38555
rect 5128 38503 5180 38555
rect 5180 38503 5194 38555
rect 5194 38503 5246 38555
rect 5246 38503 5260 38555
rect 5260 38503 5312 38555
rect 5312 38503 5326 38555
rect 5326 38503 5378 38555
rect 5378 38503 5392 38555
rect 5392 38503 5444 38555
rect 5444 38503 5551 38555
rect 4775 38491 5551 38503
rect 4775 38439 4784 38491
rect 4784 38439 4798 38491
rect 4798 38439 4850 38491
rect 4850 38439 4864 38491
rect 4864 38439 4916 38491
rect 4916 38439 4930 38491
rect 4930 38439 4982 38491
rect 4982 38439 4996 38491
rect 4996 38439 5048 38491
rect 5048 38439 5062 38491
rect 5062 38439 5114 38491
rect 5114 38439 5128 38491
rect 5128 38439 5180 38491
rect 5180 38439 5194 38491
rect 5194 38439 5246 38491
rect 5246 38439 5260 38491
rect 5260 38439 5312 38491
rect 5312 38439 5326 38491
rect 5326 38439 5378 38491
rect 5378 38439 5392 38491
rect 5392 38439 5444 38491
rect 5444 38439 5551 38491
rect 4775 38427 5551 38439
rect 4775 38375 4784 38427
rect 4784 38375 4798 38427
rect 4798 38375 4850 38427
rect 4850 38375 4864 38427
rect 4864 38375 4916 38427
rect 4916 38375 4930 38427
rect 4930 38375 4982 38427
rect 4982 38375 4996 38427
rect 4996 38375 5048 38427
rect 5048 38375 5062 38427
rect 5062 38375 5114 38427
rect 5114 38375 5128 38427
rect 5128 38375 5180 38427
rect 5180 38375 5194 38427
rect 5194 38375 5246 38427
rect 5246 38375 5260 38427
rect 5260 38375 5312 38427
rect 5312 38375 5326 38427
rect 5326 38375 5378 38427
rect 5378 38375 5392 38427
rect 5392 38375 5444 38427
rect 5444 38375 5551 38427
rect 4775 38363 5551 38375
rect 4775 38311 4784 38363
rect 4784 38311 4798 38363
rect 4798 38311 4850 38363
rect 4850 38311 4864 38363
rect 4864 38311 4916 38363
rect 4916 38311 4930 38363
rect 4930 38311 4982 38363
rect 4982 38311 4996 38363
rect 4996 38311 5048 38363
rect 5048 38311 5062 38363
rect 5062 38311 5114 38363
rect 5114 38311 5128 38363
rect 5128 38311 5180 38363
rect 5180 38311 5194 38363
rect 5194 38311 5246 38363
rect 5246 38311 5260 38363
rect 5260 38311 5312 38363
rect 5312 38311 5326 38363
rect 5326 38311 5378 38363
rect 5378 38311 5392 38363
rect 5392 38311 5444 38363
rect 5444 38311 5551 38363
rect 4775 38299 5551 38311
rect 4775 38247 4784 38299
rect 4784 38247 4798 38299
rect 4798 38247 4850 38299
rect 4850 38247 4864 38299
rect 4864 38247 4916 38299
rect 4916 38247 4930 38299
rect 4930 38247 4982 38299
rect 4982 38247 4996 38299
rect 4996 38247 5048 38299
rect 5048 38247 5062 38299
rect 5062 38247 5114 38299
rect 5114 38247 5128 38299
rect 5128 38247 5180 38299
rect 5180 38247 5194 38299
rect 5194 38247 5246 38299
rect 5246 38247 5260 38299
rect 5260 38247 5312 38299
rect 5312 38247 5326 38299
rect 5326 38247 5378 38299
rect 5378 38247 5392 38299
rect 5392 38247 5444 38299
rect 5444 38247 5551 38299
rect 4775 38235 5551 38247
rect 4775 38183 4784 38235
rect 4784 38183 4798 38235
rect 4798 38183 4850 38235
rect 4850 38183 4864 38235
rect 4864 38183 4916 38235
rect 4916 38183 4930 38235
rect 4930 38183 4982 38235
rect 4982 38183 4996 38235
rect 4996 38183 5048 38235
rect 5048 38183 5062 38235
rect 5062 38183 5114 38235
rect 5114 38183 5128 38235
rect 5128 38183 5180 38235
rect 5180 38183 5194 38235
rect 5194 38183 5246 38235
rect 5246 38183 5260 38235
rect 5260 38183 5312 38235
rect 5312 38183 5326 38235
rect 5326 38183 5378 38235
rect 5378 38183 5392 38235
rect 5392 38183 5444 38235
rect 5444 38183 5551 38235
rect 4775 38171 5551 38183
rect 4775 38119 4784 38171
rect 4784 38119 4798 38171
rect 4798 38119 4850 38171
rect 4850 38119 4864 38171
rect 4864 38119 4916 38171
rect 4916 38119 4930 38171
rect 4930 38119 4982 38171
rect 4982 38119 4996 38171
rect 4996 38119 5048 38171
rect 5048 38119 5062 38171
rect 5062 38119 5114 38171
rect 5114 38119 5128 38171
rect 5128 38119 5180 38171
rect 5180 38119 5194 38171
rect 5194 38119 5246 38171
rect 5246 38119 5260 38171
rect 5260 38119 5312 38171
rect 5312 38119 5326 38171
rect 5326 38119 5378 38171
rect 5378 38119 5392 38171
rect 5392 38119 5444 38171
rect 5444 38119 5551 38171
rect 4775 38107 5551 38119
rect 4775 38055 4784 38107
rect 4784 38055 4798 38107
rect 4798 38055 4850 38107
rect 4850 38055 4864 38107
rect 4864 38055 4916 38107
rect 4916 38055 4930 38107
rect 4930 38055 4982 38107
rect 4982 38055 4996 38107
rect 4996 38055 5048 38107
rect 5048 38055 5062 38107
rect 5062 38055 5114 38107
rect 5114 38055 5128 38107
rect 5128 38055 5180 38107
rect 5180 38055 5194 38107
rect 5194 38055 5246 38107
rect 5246 38055 5260 38107
rect 5260 38055 5312 38107
rect 5312 38055 5326 38107
rect 5326 38055 5378 38107
rect 5378 38055 5392 38107
rect 5392 38055 5444 38107
rect 5444 38055 5551 38107
rect 4775 38043 5551 38055
rect 4775 37991 4784 38043
rect 4784 37991 4798 38043
rect 4798 37991 4850 38043
rect 4850 37991 4864 38043
rect 4864 37991 4916 38043
rect 4916 37991 4930 38043
rect 4930 37991 4982 38043
rect 4982 37991 4996 38043
rect 4996 37991 5048 38043
rect 5048 37991 5062 38043
rect 5062 37991 5114 38043
rect 5114 37991 5128 38043
rect 5128 37991 5180 38043
rect 5180 37991 5194 38043
rect 5194 37991 5246 38043
rect 5246 37991 5260 38043
rect 5260 37991 5312 38043
rect 5312 37991 5326 38043
rect 5326 37991 5378 38043
rect 5378 37991 5392 38043
rect 5392 37991 5444 38043
rect 5444 37991 5551 38043
rect 4775 37979 5551 37991
rect 4775 37927 4784 37979
rect 4784 37927 4798 37979
rect 4798 37927 4850 37979
rect 4850 37927 4864 37979
rect 4864 37927 4916 37979
rect 4916 37927 4930 37979
rect 4930 37927 4982 37979
rect 4982 37927 4996 37979
rect 4996 37927 5048 37979
rect 5048 37927 5062 37979
rect 5062 37927 5114 37979
rect 5114 37927 5128 37979
rect 5128 37927 5180 37979
rect 5180 37927 5194 37979
rect 5194 37927 5246 37979
rect 5246 37927 5260 37979
rect 5260 37927 5312 37979
rect 5312 37927 5326 37979
rect 5326 37927 5378 37979
rect 5378 37927 5392 37979
rect 5392 37927 5444 37979
rect 5444 37927 5551 37979
rect 4775 37915 5551 37927
rect 4775 37863 4784 37915
rect 4784 37863 4798 37915
rect 4798 37863 4850 37915
rect 4850 37863 4864 37915
rect 4864 37863 4916 37915
rect 4916 37863 4930 37915
rect 4930 37863 4982 37915
rect 4982 37863 4996 37915
rect 4996 37863 5048 37915
rect 5048 37863 5062 37915
rect 5062 37863 5114 37915
rect 5114 37863 5128 37915
rect 5128 37863 5180 37915
rect 5180 37863 5194 37915
rect 5194 37863 5246 37915
rect 5246 37863 5260 37915
rect 5260 37863 5312 37915
rect 5312 37863 5326 37915
rect 5326 37863 5378 37915
rect 5378 37863 5392 37915
rect 5392 37863 5444 37915
rect 5444 37863 5551 37915
rect 4775 37851 5551 37863
rect 4775 37799 4784 37851
rect 4784 37799 4798 37851
rect 4798 37799 4850 37851
rect 4850 37799 4864 37851
rect 4864 37799 4916 37851
rect 4916 37799 4930 37851
rect 4930 37799 4982 37851
rect 4982 37799 4996 37851
rect 4996 37799 5048 37851
rect 5048 37799 5062 37851
rect 5062 37799 5114 37851
rect 5114 37799 5128 37851
rect 5128 37799 5180 37851
rect 5180 37799 5194 37851
rect 5194 37799 5246 37851
rect 5246 37799 5260 37851
rect 5260 37799 5312 37851
rect 5312 37799 5326 37851
rect 5326 37799 5378 37851
rect 5378 37799 5392 37851
rect 5392 37799 5444 37851
rect 5444 37799 5551 37851
rect 4775 37787 5551 37799
rect 4775 37735 4784 37787
rect 4784 37735 4798 37787
rect 4798 37735 4850 37787
rect 4850 37735 4864 37787
rect 4864 37735 4916 37787
rect 4916 37735 4930 37787
rect 4930 37735 4982 37787
rect 4982 37735 4996 37787
rect 4996 37735 5048 37787
rect 5048 37735 5062 37787
rect 5062 37735 5114 37787
rect 5114 37735 5128 37787
rect 5128 37735 5180 37787
rect 5180 37735 5194 37787
rect 5194 37735 5246 37787
rect 5246 37735 5260 37787
rect 5260 37735 5312 37787
rect 5312 37735 5326 37787
rect 5326 37735 5378 37787
rect 5378 37735 5392 37787
rect 5392 37735 5444 37787
rect 5444 37735 5551 37787
rect 4775 37723 5551 37735
rect 4775 37671 4784 37723
rect 4784 37671 4798 37723
rect 4798 37671 4850 37723
rect 4850 37671 4864 37723
rect 4864 37671 4916 37723
rect 4916 37671 4930 37723
rect 4930 37671 4982 37723
rect 4982 37671 4996 37723
rect 4996 37671 5048 37723
rect 5048 37671 5062 37723
rect 5062 37671 5114 37723
rect 5114 37671 5128 37723
rect 5128 37671 5180 37723
rect 5180 37671 5194 37723
rect 5194 37671 5246 37723
rect 5246 37671 5260 37723
rect 5260 37671 5312 37723
rect 5312 37671 5326 37723
rect 5326 37671 5378 37723
rect 5378 37671 5392 37723
rect 5392 37671 5444 37723
rect 5444 37671 5551 37723
rect 4775 37659 5551 37671
rect 4775 37607 4784 37659
rect 4784 37607 4798 37659
rect 4798 37607 4850 37659
rect 4850 37607 4864 37659
rect 4864 37607 4916 37659
rect 4916 37607 4930 37659
rect 4930 37607 4982 37659
rect 4982 37607 4996 37659
rect 4996 37607 5048 37659
rect 5048 37607 5062 37659
rect 5062 37607 5114 37659
rect 5114 37607 5128 37659
rect 5128 37607 5180 37659
rect 5180 37607 5194 37659
rect 5194 37607 5246 37659
rect 5246 37607 5260 37659
rect 5260 37607 5312 37659
rect 5312 37607 5326 37659
rect 5326 37607 5378 37659
rect 5378 37607 5392 37659
rect 5392 37607 5444 37659
rect 5444 37607 5551 37659
rect 4775 37595 5551 37607
rect 4775 37543 4784 37595
rect 4784 37543 4798 37595
rect 4798 37543 4850 37595
rect 4850 37543 4864 37595
rect 4864 37543 4916 37595
rect 4916 37543 4930 37595
rect 4930 37543 4982 37595
rect 4982 37543 4996 37595
rect 4996 37543 5048 37595
rect 5048 37543 5062 37595
rect 5062 37543 5114 37595
rect 5114 37543 5128 37595
rect 5128 37543 5180 37595
rect 5180 37543 5194 37595
rect 5194 37543 5246 37595
rect 5246 37543 5260 37595
rect 5260 37543 5312 37595
rect 5312 37543 5326 37595
rect 5326 37543 5378 37595
rect 5378 37543 5392 37595
rect 5392 37543 5444 37595
rect 5444 37543 5551 37595
rect 4775 37531 5551 37543
rect 4775 37479 4784 37531
rect 4784 37479 4798 37531
rect 4798 37479 4850 37531
rect 4850 37479 4864 37531
rect 4864 37479 4916 37531
rect 4916 37479 4930 37531
rect 4930 37479 4982 37531
rect 4982 37479 4996 37531
rect 4996 37479 5048 37531
rect 5048 37479 5062 37531
rect 5062 37479 5114 37531
rect 5114 37479 5128 37531
rect 5128 37479 5180 37531
rect 5180 37479 5194 37531
rect 5194 37479 5246 37531
rect 5246 37479 5260 37531
rect 5260 37479 5312 37531
rect 5312 37479 5326 37531
rect 5326 37479 5378 37531
rect 5378 37479 5392 37531
rect 5392 37479 5444 37531
rect 5444 37479 5551 37531
rect 4775 37467 5551 37479
rect 4775 37415 4784 37467
rect 4784 37415 4798 37467
rect 4798 37415 4850 37467
rect 4850 37415 4864 37467
rect 4864 37415 4916 37467
rect 4916 37415 4930 37467
rect 4930 37415 4982 37467
rect 4982 37415 4996 37467
rect 4996 37415 5048 37467
rect 5048 37415 5062 37467
rect 5062 37415 5114 37467
rect 5114 37415 5128 37467
rect 5128 37415 5180 37467
rect 5180 37415 5194 37467
rect 5194 37415 5246 37467
rect 5246 37415 5260 37467
rect 5260 37415 5312 37467
rect 5312 37415 5326 37467
rect 5326 37415 5378 37467
rect 5378 37415 5392 37467
rect 5392 37415 5444 37467
rect 5444 37415 5551 37467
rect 4775 37403 5551 37415
rect 4775 37351 4784 37403
rect 4784 37351 4798 37403
rect 4798 37351 4850 37403
rect 4850 37351 4864 37403
rect 4864 37351 4916 37403
rect 4916 37351 4930 37403
rect 4930 37351 4982 37403
rect 4982 37351 4996 37403
rect 4996 37351 5048 37403
rect 5048 37351 5062 37403
rect 5062 37351 5114 37403
rect 5114 37351 5128 37403
rect 5128 37351 5180 37403
rect 5180 37351 5194 37403
rect 5194 37351 5246 37403
rect 5246 37351 5260 37403
rect 5260 37351 5312 37403
rect 5312 37351 5326 37403
rect 5326 37351 5378 37403
rect 5378 37351 5392 37403
rect 5392 37351 5444 37403
rect 5444 37351 5551 37403
rect 4775 37339 5551 37351
rect 4775 37287 4784 37339
rect 4784 37287 4798 37339
rect 4798 37287 4850 37339
rect 4850 37287 4864 37339
rect 4864 37287 4916 37339
rect 4916 37287 4930 37339
rect 4930 37287 4982 37339
rect 4982 37287 4996 37339
rect 4996 37287 5048 37339
rect 5048 37287 5062 37339
rect 5062 37287 5114 37339
rect 5114 37287 5128 37339
rect 5128 37287 5180 37339
rect 5180 37287 5194 37339
rect 5194 37287 5246 37339
rect 5246 37287 5260 37339
rect 5260 37287 5312 37339
rect 5312 37287 5326 37339
rect 5326 37287 5378 37339
rect 5378 37287 5392 37339
rect 5392 37287 5444 37339
rect 5444 37287 5551 37339
rect 4775 37275 5551 37287
rect 4775 37223 4784 37275
rect 4784 37223 4798 37275
rect 4798 37223 4850 37275
rect 4850 37223 4864 37275
rect 4864 37223 4916 37275
rect 4916 37223 4930 37275
rect 4930 37223 4982 37275
rect 4982 37223 4996 37275
rect 4996 37223 5048 37275
rect 5048 37223 5062 37275
rect 5062 37223 5114 37275
rect 5114 37223 5128 37275
rect 5128 37223 5180 37275
rect 5180 37223 5194 37275
rect 5194 37223 5246 37275
rect 5246 37223 5260 37275
rect 5260 37223 5312 37275
rect 5312 37223 5326 37275
rect 5326 37223 5378 37275
rect 5378 37223 5392 37275
rect 5392 37223 5444 37275
rect 5444 37223 5551 37275
rect 4775 37211 5551 37223
rect 4775 37159 4784 37211
rect 4784 37159 4798 37211
rect 4798 37159 4850 37211
rect 4850 37159 4864 37211
rect 4864 37159 4916 37211
rect 4916 37159 4930 37211
rect 4930 37159 4982 37211
rect 4982 37159 4996 37211
rect 4996 37159 5048 37211
rect 5048 37159 5062 37211
rect 5062 37159 5114 37211
rect 5114 37159 5128 37211
rect 5128 37159 5180 37211
rect 5180 37159 5194 37211
rect 5194 37159 5246 37211
rect 5246 37159 5260 37211
rect 5260 37159 5312 37211
rect 5312 37159 5326 37211
rect 5326 37159 5378 37211
rect 5378 37159 5392 37211
rect 5392 37159 5444 37211
rect 5444 37159 5551 37211
rect 4775 37147 5551 37159
rect 4775 37095 4784 37147
rect 4784 37095 4798 37147
rect 4798 37095 4850 37147
rect 4850 37095 4864 37147
rect 4864 37095 4916 37147
rect 4916 37095 4930 37147
rect 4930 37095 4982 37147
rect 4982 37095 4996 37147
rect 4996 37095 5048 37147
rect 5048 37095 5062 37147
rect 5062 37095 5114 37147
rect 5114 37095 5128 37147
rect 5128 37095 5180 37147
rect 5180 37095 5194 37147
rect 5194 37095 5246 37147
rect 5246 37095 5260 37147
rect 5260 37095 5312 37147
rect 5312 37095 5326 37147
rect 5326 37095 5378 37147
rect 5378 37095 5392 37147
rect 5392 37095 5444 37147
rect 5444 37095 5551 37147
rect 4775 37083 5551 37095
rect 4775 37031 4784 37083
rect 4784 37031 4798 37083
rect 4798 37031 4850 37083
rect 4850 37031 4864 37083
rect 4864 37031 4916 37083
rect 4916 37031 4930 37083
rect 4930 37031 4982 37083
rect 4982 37031 4996 37083
rect 4996 37031 5048 37083
rect 5048 37031 5062 37083
rect 5062 37031 5114 37083
rect 5114 37031 5128 37083
rect 5128 37031 5180 37083
rect 5180 37031 5194 37083
rect 5194 37031 5246 37083
rect 5246 37031 5260 37083
rect 5260 37031 5312 37083
rect 5312 37031 5326 37083
rect 5326 37031 5378 37083
rect 5378 37031 5392 37083
rect 5392 37031 5444 37083
rect 5444 37031 5551 37083
rect 4775 37019 5551 37031
rect 4775 36967 4784 37019
rect 4784 36967 4798 37019
rect 4798 36967 4850 37019
rect 4850 36967 4864 37019
rect 4864 36967 4916 37019
rect 4916 36967 4930 37019
rect 4930 36967 4982 37019
rect 4982 36967 4996 37019
rect 4996 36967 5048 37019
rect 5048 36967 5062 37019
rect 5062 36967 5114 37019
rect 5114 36967 5128 37019
rect 5128 36967 5180 37019
rect 5180 36967 5194 37019
rect 5194 36967 5246 37019
rect 5246 36967 5260 37019
rect 5260 36967 5312 37019
rect 5312 36967 5326 37019
rect 5326 36967 5378 37019
rect 5378 36967 5392 37019
rect 5392 36967 5444 37019
rect 5444 36967 5551 37019
rect 4775 36955 5551 36967
rect 4775 36903 4784 36955
rect 4784 36903 4798 36955
rect 4798 36903 4850 36955
rect 4850 36903 4864 36955
rect 4864 36903 4916 36955
rect 4916 36903 4930 36955
rect 4930 36903 4982 36955
rect 4982 36903 4996 36955
rect 4996 36903 5048 36955
rect 5048 36903 5062 36955
rect 5062 36903 5114 36955
rect 5114 36903 5128 36955
rect 5128 36903 5180 36955
rect 5180 36903 5194 36955
rect 5194 36903 5246 36955
rect 5246 36903 5260 36955
rect 5260 36903 5312 36955
rect 5312 36903 5326 36955
rect 5326 36903 5378 36955
rect 5378 36903 5392 36955
rect 5392 36903 5444 36955
rect 5444 36903 5551 36955
rect 4775 36891 5551 36903
rect 4775 36839 4784 36891
rect 4784 36839 4798 36891
rect 4798 36839 4850 36891
rect 4850 36839 4864 36891
rect 4864 36839 4916 36891
rect 4916 36839 4930 36891
rect 4930 36839 4982 36891
rect 4982 36839 4996 36891
rect 4996 36839 5048 36891
rect 5048 36839 5062 36891
rect 5062 36839 5114 36891
rect 5114 36839 5128 36891
rect 5128 36839 5180 36891
rect 5180 36839 5194 36891
rect 5194 36839 5246 36891
rect 5246 36839 5260 36891
rect 5260 36839 5312 36891
rect 5312 36839 5326 36891
rect 5326 36839 5378 36891
rect 5378 36839 5392 36891
rect 5392 36839 5444 36891
rect 5444 36839 5551 36891
rect 4775 36827 5551 36839
rect 4775 36775 4784 36827
rect 4784 36775 4798 36827
rect 4798 36775 4850 36827
rect 4850 36775 4864 36827
rect 4864 36775 4916 36827
rect 4916 36775 4930 36827
rect 4930 36775 4982 36827
rect 4982 36775 4996 36827
rect 4996 36775 5048 36827
rect 5048 36775 5062 36827
rect 5062 36775 5114 36827
rect 5114 36775 5128 36827
rect 5128 36775 5180 36827
rect 5180 36775 5194 36827
rect 5194 36775 5246 36827
rect 5246 36775 5260 36827
rect 5260 36775 5312 36827
rect 5312 36775 5326 36827
rect 5326 36775 5378 36827
rect 5378 36775 5392 36827
rect 5392 36775 5444 36827
rect 5444 36775 5551 36827
rect 4775 36763 5551 36775
rect 4775 36711 4784 36763
rect 4784 36711 4798 36763
rect 4798 36711 4850 36763
rect 4850 36711 4864 36763
rect 4864 36711 4916 36763
rect 4916 36711 4930 36763
rect 4930 36711 4982 36763
rect 4982 36711 4996 36763
rect 4996 36711 5048 36763
rect 5048 36711 5062 36763
rect 5062 36711 5114 36763
rect 5114 36711 5128 36763
rect 5128 36711 5180 36763
rect 5180 36711 5194 36763
rect 5194 36711 5246 36763
rect 5246 36711 5260 36763
rect 5260 36711 5312 36763
rect 5312 36711 5326 36763
rect 5326 36711 5378 36763
rect 5378 36711 5392 36763
rect 5392 36711 5444 36763
rect 5444 36711 5551 36763
rect 4775 36699 5551 36711
rect 4775 36647 4784 36699
rect 4784 36647 4798 36699
rect 4798 36647 4850 36699
rect 4850 36647 4864 36699
rect 4864 36647 4916 36699
rect 4916 36647 4930 36699
rect 4930 36647 4982 36699
rect 4982 36647 4996 36699
rect 4996 36647 5048 36699
rect 5048 36647 5062 36699
rect 5062 36647 5114 36699
rect 5114 36647 5128 36699
rect 5128 36647 5180 36699
rect 5180 36647 5194 36699
rect 5194 36647 5246 36699
rect 5246 36647 5260 36699
rect 5260 36647 5312 36699
rect 5312 36647 5326 36699
rect 5326 36647 5378 36699
rect 5378 36647 5392 36699
rect 5392 36647 5444 36699
rect 5444 36647 5551 36699
rect 4775 36635 5551 36647
rect 4775 36583 4784 36635
rect 4784 36583 4798 36635
rect 4798 36583 4850 36635
rect 4850 36583 4864 36635
rect 4864 36583 4916 36635
rect 4916 36583 4930 36635
rect 4930 36583 4982 36635
rect 4982 36583 4996 36635
rect 4996 36583 5048 36635
rect 5048 36583 5062 36635
rect 5062 36583 5114 36635
rect 5114 36583 5128 36635
rect 5128 36583 5180 36635
rect 5180 36583 5194 36635
rect 5194 36583 5246 36635
rect 5246 36583 5260 36635
rect 5260 36583 5312 36635
rect 5312 36583 5326 36635
rect 5326 36583 5378 36635
rect 5378 36583 5392 36635
rect 5392 36583 5444 36635
rect 5444 36583 5551 36635
rect 4775 36571 5551 36583
rect 4775 36519 4784 36571
rect 4784 36519 4798 36571
rect 4798 36519 4850 36571
rect 4850 36519 4864 36571
rect 4864 36519 4916 36571
rect 4916 36519 4930 36571
rect 4930 36519 4982 36571
rect 4982 36519 4996 36571
rect 4996 36519 5048 36571
rect 5048 36519 5062 36571
rect 5062 36519 5114 36571
rect 5114 36519 5128 36571
rect 5128 36519 5180 36571
rect 5180 36519 5194 36571
rect 5194 36519 5246 36571
rect 5246 36519 5260 36571
rect 5260 36519 5312 36571
rect 5312 36519 5326 36571
rect 5326 36519 5378 36571
rect 5378 36519 5392 36571
rect 5392 36519 5444 36571
rect 5444 36519 5551 36571
rect 4775 36507 5551 36519
rect 4775 36455 4784 36507
rect 4784 36455 4798 36507
rect 4798 36455 4850 36507
rect 4850 36455 4864 36507
rect 4864 36455 4916 36507
rect 4916 36455 4930 36507
rect 4930 36455 4982 36507
rect 4982 36455 4996 36507
rect 4996 36455 5048 36507
rect 5048 36455 5062 36507
rect 5062 36455 5114 36507
rect 5114 36455 5128 36507
rect 5128 36455 5180 36507
rect 5180 36455 5194 36507
rect 5194 36455 5246 36507
rect 5246 36455 5260 36507
rect 5260 36455 5312 36507
rect 5312 36455 5326 36507
rect 5326 36455 5378 36507
rect 5378 36455 5392 36507
rect 5392 36455 5444 36507
rect 5444 36455 5551 36507
rect 4775 36443 5551 36455
rect 4775 36416 4784 36443
rect 4784 36416 4798 36443
rect 4798 36416 4850 36443
rect 4850 36416 4864 36443
rect 4864 36416 4916 36443
rect 4916 36416 4930 36443
rect 4930 36416 4982 36443
rect 4982 36416 4996 36443
rect 4996 36416 5048 36443
rect 5048 36416 5062 36443
rect 5062 36416 5114 36443
rect 5114 36416 5128 36443
rect 5128 36416 5180 36443
rect 5180 36416 5194 36443
rect 5194 36416 5246 36443
rect 5246 36416 5260 36443
rect 5260 36416 5312 36443
rect 5312 36416 5326 36443
rect 5326 36416 5378 36443
rect 5378 36416 5392 36443
rect 5392 36416 5444 36443
rect 5444 36416 5551 36443
rect 4775 36379 4831 36391
rect 4855 36379 4911 36391
rect 4935 36379 4991 36391
rect 5015 36379 5071 36391
rect 5095 36379 5151 36391
rect 5175 36379 5231 36391
rect 5255 36379 5311 36391
rect 5335 36379 5391 36391
rect 5415 36379 5471 36391
rect 4775 36335 4784 36379
rect 4784 36335 4798 36379
rect 4798 36335 4831 36379
rect 4855 36335 4864 36379
rect 4864 36335 4911 36379
rect 4935 36335 4982 36379
rect 4982 36335 4991 36379
rect 5015 36335 5048 36379
rect 5048 36335 5062 36379
rect 5062 36335 5071 36379
rect 5095 36335 5114 36379
rect 5114 36335 5128 36379
rect 5128 36335 5151 36379
rect 5175 36335 5180 36379
rect 5180 36335 5194 36379
rect 5194 36335 5231 36379
rect 5255 36335 5260 36379
rect 5260 36335 5311 36379
rect 5335 36335 5378 36379
rect 5378 36335 5391 36379
rect 5415 36335 5444 36379
rect 5444 36335 5471 36379
rect 5495 36335 5551 36391
rect 4775 36263 4784 36310
rect 4784 36263 4798 36310
rect 4798 36263 4831 36310
rect 4855 36263 4864 36310
rect 4864 36263 4911 36310
rect 4935 36263 4982 36310
rect 4982 36263 4991 36310
rect 5015 36263 5048 36310
rect 5048 36263 5062 36310
rect 5062 36263 5071 36310
rect 5095 36263 5114 36310
rect 5114 36263 5128 36310
rect 5128 36263 5151 36310
rect 5175 36263 5180 36310
rect 5180 36263 5194 36310
rect 5194 36263 5231 36310
rect 5255 36263 5260 36310
rect 5260 36263 5311 36310
rect 5335 36263 5378 36310
rect 5378 36263 5391 36310
rect 5415 36263 5444 36310
rect 5444 36263 5471 36310
rect 4775 36254 4831 36263
rect 4855 36254 4911 36263
rect 4935 36254 4991 36263
rect 5015 36254 5071 36263
rect 5095 36254 5151 36263
rect 5175 36254 5231 36263
rect 5255 36254 5311 36263
rect 5335 36254 5391 36263
rect 5415 36254 5471 36263
rect 5495 36254 5551 36310
rect 4775 36199 4784 36229
rect 4784 36199 4798 36229
rect 4798 36199 4831 36229
rect 4855 36199 4864 36229
rect 4864 36199 4911 36229
rect 4935 36199 4982 36229
rect 4982 36199 4991 36229
rect 5015 36199 5048 36229
rect 5048 36199 5062 36229
rect 5062 36199 5071 36229
rect 5095 36199 5114 36229
rect 5114 36199 5128 36229
rect 5128 36199 5151 36229
rect 5175 36199 5180 36229
rect 5180 36199 5194 36229
rect 5194 36199 5231 36229
rect 5255 36199 5260 36229
rect 5260 36199 5311 36229
rect 5335 36199 5378 36229
rect 5378 36199 5391 36229
rect 5415 36199 5444 36229
rect 5444 36199 5471 36229
rect 4775 36187 4831 36199
rect 4855 36187 4911 36199
rect 4935 36187 4991 36199
rect 5015 36187 5071 36199
rect 5095 36187 5151 36199
rect 5175 36187 5231 36199
rect 5255 36187 5311 36199
rect 5335 36187 5391 36199
rect 5415 36187 5471 36199
rect 4775 36173 4784 36187
rect 4784 36173 4798 36187
rect 4798 36173 4831 36187
rect 4855 36173 4864 36187
rect 4864 36173 4911 36187
rect 4775 36135 4784 36148
rect 4784 36135 4798 36148
rect 4798 36135 4831 36148
rect 4855 36135 4864 36148
rect 4864 36135 4911 36148
rect 4935 36173 4982 36187
rect 4982 36173 4991 36187
rect 5015 36173 5048 36187
rect 5048 36173 5062 36187
rect 5062 36173 5071 36187
rect 5095 36173 5114 36187
rect 5114 36173 5128 36187
rect 5128 36173 5151 36187
rect 5175 36173 5180 36187
rect 5180 36173 5194 36187
rect 5194 36173 5231 36187
rect 5255 36173 5260 36187
rect 5260 36173 5311 36187
rect 4935 36135 4982 36148
rect 4982 36135 4991 36148
rect 5015 36135 5048 36148
rect 5048 36135 5062 36148
rect 5062 36135 5071 36148
rect 5095 36135 5114 36148
rect 5114 36135 5128 36148
rect 5128 36135 5151 36148
rect 5175 36135 5180 36148
rect 5180 36135 5194 36148
rect 5194 36135 5231 36148
rect 5255 36135 5260 36148
rect 5260 36135 5311 36148
rect 5335 36173 5378 36187
rect 5378 36173 5391 36187
rect 5415 36173 5444 36187
rect 5444 36173 5471 36187
rect 5495 36173 5551 36229
rect 5335 36135 5378 36148
rect 5378 36135 5391 36148
rect 5415 36135 5444 36148
rect 5444 36135 5471 36148
rect 4775 36123 4831 36135
rect 4855 36123 4911 36135
rect 4935 36123 4991 36135
rect 5015 36123 5071 36135
rect 5095 36123 5151 36135
rect 5175 36123 5231 36135
rect 5255 36123 5311 36135
rect 5335 36123 5391 36135
rect 5415 36123 5471 36135
rect 4775 36092 4784 36123
rect 4784 36092 4798 36123
rect 4798 36092 4831 36123
rect 4855 36092 4864 36123
rect 4864 36092 4911 36123
rect 4935 36092 4982 36123
rect 4982 36092 4991 36123
rect 5015 36092 5048 36123
rect 5048 36092 5062 36123
rect 5062 36092 5071 36123
rect 5095 36092 5114 36123
rect 5114 36092 5128 36123
rect 5128 36092 5151 36123
rect 5175 36092 5180 36123
rect 5180 36092 5194 36123
rect 5194 36092 5231 36123
rect 5255 36092 5260 36123
rect 5260 36092 5311 36123
rect 5335 36092 5378 36123
rect 5378 36092 5391 36123
rect 5415 36092 5444 36123
rect 5444 36092 5471 36123
rect 5495 36092 5551 36148
rect 4775 36059 4831 36067
rect 4855 36059 4911 36067
rect 4935 36059 4991 36067
rect 5015 36059 5071 36067
rect 5095 36059 5151 36067
rect 5175 36059 5231 36067
rect 5255 36059 5311 36067
rect 5335 36059 5391 36067
rect 5415 36059 5471 36067
rect 4775 36011 4784 36059
rect 4784 36011 4798 36059
rect 4798 36011 4831 36059
rect 4855 36011 4864 36059
rect 4864 36011 4911 36059
rect 4935 36011 4982 36059
rect 4982 36011 4991 36059
rect 5015 36011 5048 36059
rect 5048 36011 5062 36059
rect 5062 36011 5071 36059
rect 5095 36011 5114 36059
rect 5114 36011 5128 36059
rect 5128 36011 5151 36059
rect 5175 36011 5180 36059
rect 5180 36011 5194 36059
rect 5194 36011 5231 36059
rect 5255 36011 5260 36059
rect 5260 36011 5311 36059
rect 5335 36011 5378 36059
rect 5378 36011 5391 36059
rect 5415 36011 5444 36059
rect 5444 36011 5471 36059
rect 5495 36011 5551 36067
rect 4775 35943 4784 35986
rect 4784 35943 4798 35986
rect 4798 35943 4831 35986
rect 4855 35943 4864 35986
rect 4864 35943 4911 35986
rect 4935 35943 4982 35986
rect 4982 35943 4991 35986
rect 5015 35943 5048 35986
rect 5048 35943 5062 35986
rect 5062 35943 5071 35986
rect 5095 35943 5114 35986
rect 5114 35943 5128 35986
rect 5128 35943 5151 35986
rect 5175 35943 5180 35986
rect 5180 35943 5194 35986
rect 5194 35943 5231 35986
rect 5255 35943 5260 35986
rect 5260 35943 5311 35986
rect 5335 35943 5378 35986
rect 5378 35943 5391 35986
rect 5415 35943 5444 35986
rect 5444 35943 5471 35986
rect 4775 35931 4831 35943
rect 4855 35931 4911 35943
rect 4935 35931 4991 35943
rect 5015 35931 5071 35943
rect 5095 35931 5151 35943
rect 5175 35931 5231 35943
rect 5255 35931 5311 35943
rect 5335 35931 5391 35943
rect 5415 35931 5471 35943
rect 4775 35930 4784 35931
rect 4784 35930 4798 35931
rect 4798 35930 4831 35931
rect 4855 35930 4864 35931
rect 4864 35930 4911 35931
rect 4775 35879 4784 35905
rect 4784 35879 4798 35905
rect 4798 35879 4831 35905
rect 4855 35879 4864 35905
rect 4864 35879 4911 35905
rect 4935 35930 4982 35931
rect 4982 35930 4991 35931
rect 5015 35930 5048 35931
rect 5048 35930 5062 35931
rect 5062 35930 5071 35931
rect 5095 35930 5114 35931
rect 5114 35930 5128 35931
rect 5128 35930 5151 35931
rect 5175 35930 5180 35931
rect 5180 35930 5194 35931
rect 5194 35930 5231 35931
rect 5255 35930 5260 35931
rect 5260 35930 5311 35931
rect 4935 35879 4982 35905
rect 4982 35879 4991 35905
rect 5015 35879 5048 35905
rect 5048 35879 5062 35905
rect 5062 35879 5071 35905
rect 5095 35879 5114 35905
rect 5114 35879 5128 35905
rect 5128 35879 5151 35905
rect 5175 35879 5180 35905
rect 5180 35879 5194 35905
rect 5194 35879 5231 35905
rect 5255 35879 5260 35905
rect 5260 35879 5311 35905
rect 5335 35930 5378 35931
rect 5378 35930 5391 35931
rect 5415 35930 5444 35931
rect 5444 35930 5471 35931
rect 5495 35930 5551 35986
rect 5335 35879 5378 35905
rect 5378 35879 5391 35905
rect 5415 35879 5444 35905
rect 5444 35879 5471 35905
rect 4775 35867 4831 35879
rect 4855 35867 4911 35879
rect 4935 35867 4991 35879
rect 5015 35867 5071 35879
rect 5095 35867 5151 35879
rect 5175 35867 5231 35879
rect 5255 35867 5311 35879
rect 5335 35867 5391 35879
rect 5415 35867 5471 35879
rect 4775 35849 4784 35867
rect 4784 35849 4798 35867
rect 4798 35849 4831 35867
rect 4855 35849 4864 35867
rect 4864 35849 4911 35867
rect 4775 35815 4784 35824
rect 4784 35815 4798 35824
rect 4798 35815 4831 35824
rect 4855 35815 4864 35824
rect 4864 35815 4911 35824
rect 4935 35849 4982 35867
rect 4982 35849 4991 35867
rect 5015 35849 5048 35867
rect 5048 35849 5062 35867
rect 5062 35849 5071 35867
rect 5095 35849 5114 35867
rect 5114 35849 5128 35867
rect 5128 35849 5151 35867
rect 5175 35849 5180 35867
rect 5180 35849 5194 35867
rect 5194 35849 5231 35867
rect 5255 35849 5260 35867
rect 5260 35849 5311 35867
rect 4935 35815 4982 35824
rect 4982 35815 4991 35824
rect 5015 35815 5048 35824
rect 5048 35815 5062 35824
rect 5062 35815 5071 35824
rect 5095 35815 5114 35824
rect 5114 35815 5128 35824
rect 5128 35815 5151 35824
rect 5175 35815 5180 35824
rect 5180 35815 5194 35824
rect 5194 35815 5231 35824
rect 5255 35815 5260 35824
rect 5260 35815 5311 35824
rect 5335 35849 5378 35867
rect 5378 35849 5391 35867
rect 5415 35849 5444 35867
rect 5444 35849 5471 35867
rect 5495 35849 5551 35905
rect 5335 35815 5378 35824
rect 5378 35815 5391 35824
rect 5415 35815 5444 35824
rect 5444 35815 5471 35824
rect 4775 35803 4831 35815
rect 4855 35803 4911 35815
rect 4935 35803 4991 35815
rect 5015 35803 5071 35815
rect 5095 35803 5151 35815
rect 5175 35803 5231 35815
rect 5255 35803 5311 35815
rect 5335 35803 5391 35815
rect 5415 35803 5471 35815
rect 4775 35768 4784 35803
rect 4784 35768 4798 35803
rect 4798 35768 4831 35803
rect 4855 35768 4864 35803
rect 4864 35768 4911 35803
rect 4935 35768 4982 35803
rect 4982 35768 4991 35803
rect 5015 35768 5048 35803
rect 5048 35768 5062 35803
rect 5062 35768 5071 35803
rect 5095 35768 5114 35803
rect 5114 35768 5128 35803
rect 5128 35768 5151 35803
rect 5175 35768 5180 35803
rect 5180 35768 5194 35803
rect 5194 35768 5231 35803
rect 5255 35768 5260 35803
rect 5260 35768 5311 35803
rect 5335 35768 5378 35803
rect 5378 35768 5391 35803
rect 5415 35768 5444 35803
rect 5444 35768 5471 35803
rect 5495 35768 5551 35824
rect 4775 35739 4831 35743
rect 4855 35739 4911 35743
rect 4935 35739 4991 35743
rect 5015 35739 5071 35743
rect 5095 35739 5151 35743
rect 5175 35739 5231 35743
rect 5255 35739 5311 35743
rect 5335 35739 5391 35743
rect 5415 35739 5471 35743
rect 4775 35687 4784 35739
rect 4784 35687 4798 35739
rect 4798 35687 4831 35739
rect 4855 35687 4864 35739
rect 4864 35687 4911 35739
rect 4935 35687 4982 35739
rect 4982 35687 4991 35739
rect 5015 35687 5048 35739
rect 5048 35687 5062 35739
rect 5062 35687 5071 35739
rect 5095 35687 5114 35739
rect 5114 35687 5128 35739
rect 5128 35687 5151 35739
rect 5175 35687 5180 35739
rect 5180 35687 5194 35739
rect 5194 35687 5231 35739
rect 5255 35687 5260 35739
rect 5260 35687 5311 35739
rect 5335 35687 5378 35739
rect 5378 35687 5391 35739
rect 5415 35687 5444 35739
rect 5444 35687 5471 35739
rect 5495 35687 5551 35743
rect 4775 35623 4784 35662
rect 4784 35623 4798 35662
rect 4798 35623 4831 35662
rect 4855 35623 4864 35662
rect 4864 35623 4911 35662
rect 4935 35623 4982 35662
rect 4982 35623 4991 35662
rect 5015 35623 5048 35662
rect 5048 35623 5062 35662
rect 5062 35623 5071 35662
rect 5095 35623 5114 35662
rect 5114 35623 5128 35662
rect 5128 35623 5151 35662
rect 5175 35623 5180 35662
rect 5180 35623 5194 35662
rect 5194 35623 5231 35662
rect 5255 35623 5260 35662
rect 5260 35623 5311 35662
rect 5335 35623 5378 35662
rect 5378 35623 5391 35662
rect 5415 35623 5444 35662
rect 5444 35623 5471 35662
rect 4775 35611 4831 35623
rect 4855 35611 4911 35623
rect 4935 35611 4991 35623
rect 5015 35611 5071 35623
rect 5095 35611 5151 35623
rect 5175 35611 5231 35623
rect 5255 35611 5311 35623
rect 5335 35611 5391 35623
rect 5415 35611 5471 35623
rect 4775 35606 4784 35611
rect 4784 35606 4798 35611
rect 4798 35606 4831 35611
rect 4855 35606 4864 35611
rect 4864 35606 4911 35611
rect 4775 35559 4784 35581
rect 4784 35559 4798 35581
rect 4798 35559 4831 35581
rect 4855 35559 4864 35581
rect 4864 35559 4911 35581
rect 4935 35606 4982 35611
rect 4982 35606 4991 35611
rect 5015 35606 5048 35611
rect 5048 35606 5062 35611
rect 5062 35606 5071 35611
rect 5095 35606 5114 35611
rect 5114 35606 5128 35611
rect 5128 35606 5151 35611
rect 5175 35606 5180 35611
rect 5180 35606 5194 35611
rect 5194 35606 5231 35611
rect 5255 35606 5260 35611
rect 5260 35606 5311 35611
rect 4935 35559 4982 35581
rect 4982 35559 4991 35581
rect 5015 35559 5048 35581
rect 5048 35559 5062 35581
rect 5062 35559 5071 35581
rect 5095 35559 5114 35581
rect 5114 35559 5128 35581
rect 5128 35559 5151 35581
rect 5175 35559 5180 35581
rect 5180 35559 5194 35581
rect 5194 35559 5231 35581
rect 5255 35559 5260 35581
rect 5260 35559 5311 35581
rect 5335 35606 5378 35611
rect 5378 35606 5391 35611
rect 5415 35606 5444 35611
rect 5444 35606 5471 35611
rect 5495 35606 5551 35662
rect 5335 35559 5378 35581
rect 5378 35559 5391 35581
rect 5415 35559 5444 35581
rect 5444 35559 5471 35581
rect 4775 35547 4831 35559
rect 4855 35547 4911 35559
rect 4935 35547 4991 35559
rect 5015 35547 5071 35559
rect 5095 35547 5151 35559
rect 5175 35547 5231 35559
rect 5255 35547 5311 35559
rect 5335 35547 5391 35559
rect 5415 35547 5471 35559
rect 4775 35525 4784 35547
rect 4784 35525 4798 35547
rect 4798 35525 4831 35547
rect 4855 35525 4864 35547
rect 4864 35525 4911 35547
rect 4775 35495 4784 35500
rect 4784 35495 4798 35500
rect 4798 35495 4831 35500
rect 4855 35495 4864 35500
rect 4864 35495 4911 35500
rect 4935 35525 4982 35547
rect 4982 35525 4991 35547
rect 5015 35525 5048 35547
rect 5048 35525 5062 35547
rect 5062 35525 5071 35547
rect 5095 35525 5114 35547
rect 5114 35525 5128 35547
rect 5128 35525 5151 35547
rect 5175 35525 5180 35547
rect 5180 35525 5194 35547
rect 5194 35525 5231 35547
rect 5255 35525 5260 35547
rect 5260 35525 5311 35547
rect 4935 35495 4982 35500
rect 4982 35495 4991 35500
rect 5015 35495 5048 35500
rect 5048 35495 5062 35500
rect 5062 35495 5071 35500
rect 5095 35495 5114 35500
rect 5114 35495 5128 35500
rect 5128 35495 5151 35500
rect 5175 35495 5180 35500
rect 5180 35495 5194 35500
rect 5194 35495 5231 35500
rect 5255 35495 5260 35500
rect 5260 35495 5311 35500
rect 5335 35525 5378 35547
rect 5378 35525 5391 35547
rect 5415 35525 5444 35547
rect 5444 35525 5471 35547
rect 5495 35525 5551 35581
rect 5335 35495 5378 35500
rect 5378 35495 5391 35500
rect 5415 35495 5444 35500
rect 5444 35495 5471 35500
rect 4775 35483 4831 35495
rect 4855 35483 4911 35495
rect 4935 35483 4991 35495
rect 5015 35483 5071 35495
rect 5095 35483 5151 35495
rect 5175 35483 5231 35495
rect 5255 35483 5311 35495
rect 5335 35483 5391 35495
rect 5415 35483 5471 35495
rect 4775 35444 4784 35483
rect 4784 35444 4798 35483
rect 4798 35444 4831 35483
rect 4855 35444 4864 35483
rect 4864 35444 4911 35483
rect 4935 35444 4982 35483
rect 4982 35444 4991 35483
rect 5015 35444 5048 35483
rect 5048 35444 5062 35483
rect 5062 35444 5071 35483
rect 5095 35444 5114 35483
rect 5114 35444 5128 35483
rect 5128 35444 5151 35483
rect 5175 35444 5180 35483
rect 5180 35444 5194 35483
rect 5194 35444 5231 35483
rect 5255 35444 5260 35483
rect 5260 35444 5311 35483
rect 5335 35444 5378 35483
rect 5378 35444 5391 35483
rect 5415 35444 5444 35483
rect 5444 35444 5471 35483
rect 5495 35444 5551 35500
rect 4775 35367 4784 35419
rect 4784 35367 4798 35419
rect 4798 35367 4831 35419
rect 4855 35367 4864 35419
rect 4864 35367 4911 35419
rect 4935 35367 4982 35419
rect 4982 35367 4991 35419
rect 5015 35367 5048 35419
rect 5048 35367 5062 35419
rect 5062 35367 5071 35419
rect 5095 35367 5114 35419
rect 5114 35367 5128 35419
rect 5128 35367 5151 35419
rect 5175 35367 5180 35419
rect 5180 35367 5194 35419
rect 5194 35367 5231 35419
rect 5255 35367 5260 35419
rect 5260 35367 5311 35419
rect 5335 35367 5378 35419
rect 5378 35367 5391 35419
rect 5415 35367 5444 35419
rect 5444 35367 5471 35419
rect 4775 35363 4831 35367
rect 4855 35363 4911 35367
rect 4935 35363 4991 35367
rect 5015 35363 5071 35367
rect 5095 35363 5151 35367
rect 5175 35363 5231 35367
rect 5255 35363 5311 35367
rect 5335 35363 5391 35367
rect 5415 35363 5471 35367
rect 5495 35363 5551 35419
rect 4775 35303 4784 35338
rect 4784 35303 4798 35338
rect 4798 35303 4831 35338
rect 4855 35303 4864 35338
rect 4864 35303 4911 35338
rect 4935 35303 4982 35338
rect 4982 35303 4991 35338
rect 5015 35303 5048 35338
rect 5048 35303 5062 35338
rect 5062 35303 5071 35338
rect 5095 35303 5114 35338
rect 5114 35303 5128 35338
rect 5128 35303 5151 35338
rect 5175 35303 5180 35338
rect 5180 35303 5194 35338
rect 5194 35303 5231 35338
rect 5255 35303 5260 35338
rect 5260 35303 5311 35338
rect 5335 35303 5378 35338
rect 5378 35303 5391 35338
rect 5415 35303 5444 35338
rect 5444 35303 5471 35338
rect 4775 35291 4831 35303
rect 4855 35291 4911 35303
rect 4935 35291 4991 35303
rect 5015 35291 5071 35303
rect 5095 35291 5151 35303
rect 5175 35291 5231 35303
rect 5255 35291 5311 35303
rect 5335 35291 5391 35303
rect 5415 35291 5471 35303
rect 4775 35282 4784 35291
rect 4784 35282 4798 35291
rect 4798 35282 4831 35291
rect 4855 35282 4864 35291
rect 4864 35282 4911 35291
rect 4775 35239 4784 35257
rect 4784 35239 4798 35257
rect 4798 35239 4831 35257
rect 4855 35239 4864 35257
rect 4864 35239 4911 35257
rect 4935 35282 4982 35291
rect 4982 35282 4991 35291
rect 5015 35282 5048 35291
rect 5048 35282 5062 35291
rect 5062 35282 5071 35291
rect 5095 35282 5114 35291
rect 5114 35282 5128 35291
rect 5128 35282 5151 35291
rect 5175 35282 5180 35291
rect 5180 35282 5194 35291
rect 5194 35282 5231 35291
rect 5255 35282 5260 35291
rect 5260 35282 5311 35291
rect 4935 35239 4982 35257
rect 4982 35239 4991 35257
rect 5015 35239 5048 35257
rect 5048 35239 5062 35257
rect 5062 35239 5071 35257
rect 5095 35239 5114 35257
rect 5114 35239 5128 35257
rect 5128 35239 5151 35257
rect 5175 35239 5180 35257
rect 5180 35239 5194 35257
rect 5194 35239 5231 35257
rect 5255 35239 5260 35257
rect 5260 35239 5311 35257
rect 5335 35282 5378 35291
rect 5378 35282 5391 35291
rect 5415 35282 5444 35291
rect 5444 35282 5471 35291
rect 5495 35282 5551 35338
rect 5335 35239 5378 35257
rect 5378 35239 5391 35257
rect 5415 35239 5444 35257
rect 5444 35239 5471 35257
rect 4775 35227 4831 35239
rect 4855 35227 4911 35239
rect 4935 35227 4991 35239
rect 5015 35227 5071 35239
rect 5095 35227 5151 35239
rect 5175 35227 5231 35239
rect 5255 35227 5311 35239
rect 5335 35227 5391 35239
rect 5415 35227 5471 35239
rect 4775 35201 4784 35227
rect 4784 35201 4798 35227
rect 4798 35201 4831 35227
rect 4855 35201 4864 35227
rect 4864 35201 4911 35227
rect 4775 35175 4784 35176
rect 4784 35175 4798 35176
rect 4798 35175 4831 35176
rect 4855 35175 4864 35176
rect 4864 35175 4911 35176
rect 4935 35201 4982 35227
rect 4982 35201 4991 35227
rect 5015 35201 5048 35227
rect 5048 35201 5062 35227
rect 5062 35201 5071 35227
rect 5095 35201 5114 35227
rect 5114 35201 5128 35227
rect 5128 35201 5151 35227
rect 5175 35201 5180 35227
rect 5180 35201 5194 35227
rect 5194 35201 5231 35227
rect 5255 35201 5260 35227
rect 5260 35201 5311 35227
rect 4935 35175 4982 35176
rect 4982 35175 4991 35176
rect 5015 35175 5048 35176
rect 5048 35175 5062 35176
rect 5062 35175 5071 35176
rect 5095 35175 5114 35176
rect 5114 35175 5128 35176
rect 5128 35175 5151 35176
rect 5175 35175 5180 35176
rect 5180 35175 5194 35176
rect 5194 35175 5231 35176
rect 5255 35175 5260 35176
rect 5260 35175 5311 35176
rect 5335 35201 5378 35227
rect 5378 35201 5391 35227
rect 5415 35201 5444 35227
rect 5444 35201 5471 35227
rect 5495 35201 5551 35257
rect 5335 35175 5378 35176
rect 5378 35175 5391 35176
rect 5415 35175 5444 35176
rect 5444 35175 5471 35176
rect 4775 35163 4831 35175
rect 4855 35163 4911 35175
rect 4935 35163 4991 35175
rect 5015 35163 5071 35175
rect 5095 35163 5151 35175
rect 5175 35163 5231 35175
rect 5255 35163 5311 35175
rect 5335 35163 5391 35175
rect 5415 35163 5471 35175
rect 4775 35120 4784 35163
rect 4784 35120 4798 35163
rect 4798 35120 4831 35163
rect 4855 35120 4864 35163
rect 4864 35120 4911 35163
rect 4935 35120 4982 35163
rect 4982 35120 4991 35163
rect 5015 35120 5048 35163
rect 5048 35120 5062 35163
rect 5062 35120 5071 35163
rect 5095 35120 5114 35163
rect 5114 35120 5128 35163
rect 5128 35120 5151 35163
rect 5175 35120 5180 35163
rect 5180 35120 5194 35163
rect 5194 35120 5231 35163
rect 5255 35120 5260 35163
rect 5260 35120 5311 35163
rect 5335 35120 5378 35163
rect 5378 35120 5391 35163
rect 5415 35120 5444 35163
rect 5444 35120 5471 35163
rect 5495 35120 5551 35176
rect 4775 35047 4784 35095
rect 4784 35047 4798 35095
rect 4798 35047 4831 35095
rect 4855 35047 4864 35095
rect 4864 35047 4911 35095
rect 4935 35047 4982 35095
rect 4982 35047 4991 35095
rect 5015 35047 5048 35095
rect 5048 35047 5062 35095
rect 5062 35047 5071 35095
rect 5095 35047 5114 35095
rect 5114 35047 5128 35095
rect 5128 35047 5151 35095
rect 5175 35047 5180 35095
rect 5180 35047 5194 35095
rect 5194 35047 5231 35095
rect 5255 35047 5260 35095
rect 5260 35047 5311 35095
rect 5335 35047 5378 35095
rect 5378 35047 5391 35095
rect 5415 35047 5444 35095
rect 5444 35047 5471 35095
rect 4775 35039 4831 35047
rect 4855 35039 4911 35047
rect 4935 35039 4991 35047
rect 5015 35039 5071 35047
rect 5095 35039 5151 35047
rect 5175 35039 5231 35047
rect 5255 35039 5311 35047
rect 5335 35039 5391 35047
rect 5415 35039 5471 35047
rect 5495 35039 5551 35095
rect 4775 34983 4784 35014
rect 4784 34983 4798 35014
rect 4798 34983 4831 35014
rect 4855 34983 4864 35014
rect 4864 34983 4911 35014
rect 4935 34983 4982 35014
rect 4982 34983 4991 35014
rect 5015 34983 5048 35014
rect 5048 34983 5062 35014
rect 5062 34983 5071 35014
rect 5095 34983 5114 35014
rect 5114 34983 5128 35014
rect 5128 34983 5151 35014
rect 5175 34983 5180 35014
rect 5180 34983 5194 35014
rect 5194 34983 5231 35014
rect 5255 34983 5260 35014
rect 5260 34983 5311 35014
rect 5335 34983 5378 35014
rect 5378 34983 5391 35014
rect 5415 34983 5444 35014
rect 5444 34983 5471 35014
rect 4775 34971 4831 34983
rect 4855 34971 4911 34983
rect 4935 34971 4991 34983
rect 5015 34971 5071 34983
rect 5095 34971 5151 34983
rect 5175 34971 5231 34983
rect 5255 34971 5311 34983
rect 5335 34971 5391 34983
rect 5415 34971 5471 34983
rect 4775 34958 4784 34971
rect 4784 34958 4798 34971
rect 4798 34958 4831 34971
rect 4855 34958 4864 34971
rect 4864 34958 4911 34971
rect 4775 34919 4784 34933
rect 4784 34919 4798 34933
rect 4798 34919 4831 34933
rect 4855 34919 4864 34933
rect 4864 34919 4911 34933
rect 4935 34958 4982 34971
rect 4982 34958 4991 34971
rect 5015 34958 5048 34971
rect 5048 34958 5062 34971
rect 5062 34958 5071 34971
rect 5095 34958 5114 34971
rect 5114 34958 5128 34971
rect 5128 34958 5151 34971
rect 5175 34958 5180 34971
rect 5180 34958 5194 34971
rect 5194 34958 5231 34971
rect 5255 34958 5260 34971
rect 5260 34958 5311 34971
rect 4935 34919 4982 34933
rect 4982 34919 4991 34933
rect 5015 34919 5048 34933
rect 5048 34919 5062 34933
rect 5062 34919 5071 34933
rect 5095 34919 5114 34933
rect 5114 34919 5128 34933
rect 5128 34919 5151 34933
rect 5175 34919 5180 34933
rect 5180 34919 5194 34933
rect 5194 34919 5231 34933
rect 5255 34919 5260 34933
rect 5260 34919 5311 34933
rect 5335 34958 5378 34971
rect 5378 34958 5391 34971
rect 5415 34958 5444 34971
rect 5444 34958 5471 34971
rect 5495 34958 5551 35014
rect 5335 34919 5378 34933
rect 5378 34919 5391 34933
rect 5415 34919 5444 34933
rect 5444 34919 5471 34933
rect 4775 34907 4831 34919
rect 4855 34907 4911 34919
rect 4935 34907 4991 34919
rect 5015 34907 5071 34919
rect 5095 34907 5151 34919
rect 5175 34907 5231 34919
rect 5255 34907 5311 34919
rect 5335 34907 5391 34919
rect 5415 34907 5471 34919
rect 4775 34877 4784 34907
rect 4784 34877 4798 34907
rect 4798 34877 4831 34907
rect 4855 34877 4864 34907
rect 4864 34877 4911 34907
rect 4935 34877 4982 34907
rect 4982 34877 4991 34907
rect 5015 34877 5048 34907
rect 5048 34877 5062 34907
rect 5062 34877 5071 34907
rect 5095 34877 5114 34907
rect 5114 34877 5128 34907
rect 5128 34877 5151 34907
rect 5175 34877 5180 34907
rect 5180 34877 5194 34907
rect 5194 34877 5231 34907
rect 5255 34877 5260 34907
rect 5260 34877 5311 34907
rect 5335 34877 5378 34907
rect 5378 34877 5391 34907
rect 5415 34877 5444 34907
rect 5444 34877 5471 34907
rect 5495 34877 5551 34933
rect 4775 34843 4831 34852
rect 4855 34843 4911 34852
rect 4935 34843 4991 34852
rect 5015 34843 5071 34852
rect 5095 34843 5151 34852
rect 5175 34843 5231 34852
rect 5255 34843 5311 34852
rect 5335 34843 5391 34852
rect 5415 34843 5471 34852
rect 4775 34796 4784 34843
rect 4784 34796 4798 34843
rect 4798 34796 4831 34843
rect 4855 34796 4864 34843
rect 4864 34796 4911 34843
rect 4935 34796 4982 34843
rect 4982 34796 4991 34843
rect 5015 34796 5048 34843
rect 5048 34796 5062 34843
rect 5062 34796 5071 34843
rect 5095 34796 5114 34843
rect 5114 34796 5128 34843
rect 5128 34796 5151 34843
rect 5175 34796 5180 34843
rect 5180 34796 5194 34843
rect 5194 34796 5231 34843
rect 5255 34796 5260 34843
rect 5260 34796 5311 34843
rect 5335 34796 5378 34843
rect 5378 34796 5391 34843
rect 5415 34796 5444 34843
rect 5444 34796 5471 34843
rect 5495 34796 5551 34852
rect 4775 34727 4784 34771
rect 4784 34727 4798 34771
rect 4798 34727 4831 34771
rect 4855 34727 4864 34771
rect 4864 34727 4911 34771
rect 4935 34727 4982 34771
rect 4982 34727 4991 34771
rect 5015 34727 5048 34771
rect 5048 34727 5062 34771
rect 5062 34727 5071 34771
rect 5095 34727 5114 34771
rect 5114 34727 5128 34771
rect 5128 34727 5151 34771
rect 5175 34727 5180 34771
rect 5180 34727 5194 34771
rect 5194 34727 5231 34771
rect 5255 34727 5260 34771
rect 5260 34727 5311 34771
rect 5335 34727 5378 34771
rect 5378 34727 5391 34771
rect 5415 34727 5444 34771
rect 5444 34727 5471 34771
rect 4775 34715 4831 34727
rect 4855 34715 4911 34727
rect 4935 34715 4991 34727
rect 5015 34715 5071 34727
rect 5095 34715 5151 34727
rect 5175 34715 5231 34727
rect 5255 34715 5311 34727
rect 5335 34715 5391 34727
rect 5415 34715 5471 34727
rect 5495 34715 5551 34771
rect 4775 34663 4784 34690
rect 4784 34663 4798 34690
rect 4798 34663 4831 34690
rect 4855 34663 4864 34690
rect 4864 34663 4911 34690
rect 4935 34663 4982 34690
rect 4982 34663 4991 34690
rect 5015 34663 5048 34690
rect 5048 34663 5062 34690
rect 5062 34663 5071 34690
rect 5095 34663 5114 34690
rect 5114 34663 5128 34690
rect 5128 34663 5151 34690
rect 5175 34663 5180 34690
rect 5180 34663 5194 34690
rect 5194 34663 5231 34690
rect 5255 34663 5260 34690
rect 5260 34663 5311 34690
rect 5335 34663 5378 34690
rect 5378 34663 5391 34690
rect 5415 34663 5444 34690
rect 5444 34663 5471 34690
rect 4775 34651 4831 34663
rect 4855 34651 4911 34663
rect 4935 34651 4991 34663
rect 5015 34651 5071 34663
rect 5095 34651 5151 34663
rect 5175 34651 5231 34663
rect 5255 34651 5311 34663
rect 5335 34651 5391 34663
rect 5415 34651 5471 34663
rect 4775 34634 4784 34651
rect 4784 34634 4798 34651
rect 4798 34634 4831 34651
rect 4855 34634 4864 34651
rect 4864 34634 4911 34651
rect 4775 34599 4784 34609
rect 4784 34599 4798 34609
rect 4798 34599 4831 34609
rect 4855 34599 4864 34609
rect 4864 34599 4911 34609
rect 4935 34634 4982 34651
rect 4982 34634 4991 34651
rect 5015 34634 5048 34651
rect 5048 34634 5062 34651
rect 5062 34634 5071 34651
rect 5095 34634 5114 34651
rect 5114 34634 5128 34651
rect 5128 34634 5151 34651
rect 5175 34634 5180 34651
rect 5180 34634 5194 34651
rect 5194 34634 5231 34651
rect 5255 34634 5260 34651
rect 5260 34634 5311 34651
rect 4935 34599 4982 34609
rect 4982 34599 4991 34609
rect 5015 34599 5048 34609
rect 5048 34599 5062 34609
rect 5062 34599 5071 34609
rect 5095 34599 5114 34609
rect 5114 34599 5128 34609
rect 5128 34599 5151 34609
rect 5175 34599 5180 34609
rect 5180 34599 5194 34609
rect 5194 34599 5231 34609
rect 5255 34599 5260 34609
rect 5260 34599 5311 34609
rect 5335 34634 5378 34651
rect 5378 34634 5391 34651
rect 5415 34634 5444 34651
rect 5444 34634 5471 34651
rect 5495 34634 5551 34690
rect 5335 34599 5378 34609
rect 5378 34599 5391 34609
rect 5415 34599 5444 34609
rect 5444 34599 5471 34609
rect 4775 34587 4831 34599
rect 4855 34587 4911 34599
rect 4935 34587 4991 34599
rect 5015 34587 5071 34599
rect 5095 34587 5151 34599
rect 5175 34587 5231 34599
rect 5255 34587 5311 34599
rect 5335 34587 5391 34599
rect 5415 34587 5471 34599
rect 4775 34553 4784 34587
rect 4784 34553 4798 34587
rect 4798 34553 4831 34587
rect 4855 34553 4864 34587
rect 4864 34553 4911 34587
rect 4935 34553 4982 34587
rect 4982 34553 4991 34587
rect 5015 34553 5048 34587
rect 5048 34553 5062 34587
rect 5062 34553 5071 34587
rect 5095 34553 5114 34587
rect 5114 34553 5128 34587
rect 5128 34553 5151 34587
rect 5175 34553 5180 34587
rect 5180 34553 5194 34587
rect 5194 34553 5231 34587
rect 5255 34553 5260 34587
rect 5260 34553 5311 34587
rect 5335 34553 5378 34587
rect 5378 34553 5391 34587
rect 5415 34553 5444 34587
rect 5444 34553 5471 34587
rect 5495 34553 5551 34609
rect 4775 34523 4831 34528
rect 4855 34523 4911 34528
rect 4935 34523 4991 34528
rect 5015 34523 5071 34528
rect 5095 34523 5151 34528
rect 5175 34523 5231 34528
rect 5255 34523 5311 34528
rect 5335 34523 5391 34528
rect 5415 34523 5471 34528
rect 4775 34472 4784 34523
rect 4784 34472 4798 34523
rect 4798 34472 4831 34523
rect 4855 34472 4864 34523
rect 4864 34472 4911 34523
rect 4935 34472 4982 34523
rect 4982 34472 4991 34523
rect 5015 34472 5048 34523
rect 5048 34472 5062 34523
rect 5062 34472 5071 34523
rect 5095 34472 5114 34523
rect 5114 34472 5128 34523
rect 5128 34472 5151 34523
rect 5175 34472 5180 34523
rect 5180 34472 5194 34523
rect 5194 34472 5231 34523
rect 5255 34472 5260 34523
rect 5260 34472 5311 34523
rect 5335 34472 5378 34523
rect 5378 34472 5391 34523
rect 5415 34472 5444 34523
rect 5444 34472 5471 34523
rect 5495 34472 5551 34528
rect 4775 34407 4784 34447
rect 4784 34407 4798 34447
rect 4798 34407 4831 34447
rect 4855 34407 4864 34447
rect 4864 34407 4911 34447
rect 4935 34407 4982 34447
rect 4982 34407 4991 34447
rect 5015 34407 5048 34447
rect 5048 34407 5062 34447
rect 5062 34407 5071 34447
rect 5095 34407 5114 34447
rect 5114 34407 5128 34447
rect 5128 34407 5151 34447
rect 5175 34407 5180 34447
rect 5180 34407 5194 34447
rect 5194 34407 5231 34447
rect 5255 34407 5260 34447
rect 5260 34407 5311 34447
rect 5335 34407 5378 34447
rect 5378 34407 5391 34447
rect 5415 34407 5444 34447
rect 5444 34407 5471 34447
rect 4775 34395 4831 34407
rect 4855 34395 4911 34407
rect 4935 34395 4991 34407
rect 5015 34395 5071 34407
rect 5095 34395 5151 34407
rect 5175 34395 5231 34407
rect 5255 34395 5311 34407
rect 5335 34395 5391 34407
rect 5415 34395 5471 34407
rect 4775 34391 4784 34395
rect 4784 34391 4798 34395
rect 4798 34391 4831 34395
rect 4855 34391 4864 34395
rect 4864 34391 4911 34395
rect 4775 34343 4784 34366
rect 4784 34343 4798 34366
rect 4798 34343 4831 34366
rect 4855 34343 4864 34366
rect 4864 34343 4911 34366
rect 4935 34391 4982 34395
rect 4982 34391 4991 34395
rect 5015 34391 5048 34395
rect 5048 34391 5062 34395
rect 5062 34391 5071 34395
rect 5095 34391 5114 34395
rect 5114 34391 5128 34395
rect 5128 34391 5151 34395
rect 5175 34391 5180 34395
rect 5180 34391 5194 34395
rect 5194 34391 5231 34395
rect 5255 34391 5260 34395
rect 5260 34391 5311 34395
rect 4935 34343 4982 34366
rect 4982 34343 4991 34366
rect 5015 34343 5048 34366
rect 5048 34343 5062 34366
rect 5062 34343 5071 34366
rect 5095 34343 5114 34366
rect 5114 34343 5128 34366
rect 5128 34343 5151 34366
rect 5175 34343 5180 34366
rect 5180 34343 5194 34366
rect 5194 34343 5231 34366
rect 5255 34343 5260 34366
rect 5260 34343 5311 34366
rect 5335 34391 5378 34395
rect 5378 34391 5391 34395
rect 5415 34391 5444 34395
rect 5444 34391 5471 34395
rect 5495 34391 5551 34447
rect 5335 34343 5378 34366
rect 5378 34343 5391 34366
rect 5415 34343 5444 34366
rect 5444 34343 5471 34366
rect 4775 34331 4831 34343
rect 4855 34331 4911 34343
rect 4935 34331 4991 34343
rect 5015 34331 5071 34343
rect 5095 34331 5151 34343
rect 5175 34331 5231 34343
rect 5255 34331 5311 34343
rect 5335 34331 5391 34343
rect 5415 34331 5471 34343
rect 4775 34310 4784 34331
rect 4784 34310 4798 34331
rect 4798 34310 4831 34331
rect 4855 34310 4864 34331
rect 4864 34310 4911 34331
rect 4775 34279 4784 34285
rect 4784 34279 4798 34285
rect 4798 34279 4831 34285
rect 4855 34279 4864 34285
rect 4864 34279 4911 34285
rect 4935 34310 4982 34331
rect 4982 34310 4991 34331
rect 5015 34310 5048 34331
rect 5048 34310 5062 34331
rect 5062 34310 5071 34331
rect 5095 34310 5114 34331
rect 5114 34310 5128 34331
rect 5128 34310 5151 34331
rect 5175 34310 5180 34331
rect 5180 34310 5194 34331
rect 5194 34310 5231 34331
rect 5255 34310 5260 34331
rect 5260 34310 5311 34331
rect 4935 34279 4982 34285
rect 4982 34279 4991 34285
rect 5015 34279 5048 34285
rect 5048 34279 5062 34285
rect 5062 34279 5071 34285
rect 5095 34279 5114 34285
rect 5114 34279 5128 34285
rect 5128 34279 5151 34285
rect 5175 34279 5180 34285
rect 5180 34279 5194 34285
rect 5194 34279 5231 34285
rect 5255 34279 5260 34285
rect 5260 34279 5311 34285
rect 5335 34310 5378 34331
rect 5378 34310 5391 34331
rect 5415 34310 5444 34331
rect 5444 34310 5471 34331
rect 5495 34310 5551 34366
rect 5335 34279 5378 34285
rect 5378 34279 5391 34285
rect 5415 34279 5444 34285
rect 5444 34279 5471 34285
rect 4775 34267 4831 34279
rect 4855 34267 4911 34279
rect 4935 34267 4991 34279
rect 5015 34267 5071 34279
rect 5095 34267 5151 34279
rect 5175 34267 5231 34279
rect 5255 34267 5311 34279
rect 5335 34267 5391 34279
rect 5415 34267 5471 34279
rect 4775 34229 4784 34267
rect 4784 34229 4798 34267
rect 4798 34229 4831 34267
rect 4855 34229 4864 34267
rect 4864 34229 4911 34267
rect 4935 34229 4982 34267
rect 4982 34229 4991 34267
rect 5015 34229 5048 34267
rect 5048 34229 5062 34267
rect 5062 34229 5071 34267
rect 5095 34229 5114 34267
rect 5114 34229 5128 34267
rect 5128 34229 5151 34267
rect 5175 34229 5180 34267
rect 5180 34229 5194 34267
rect 5194 34229 5231 34267
rect 5255 34229 5260 34267
rect 5260 34229 5311 34267
rect 5335 34229 5378 34267
rect 5378 34229 5391 34267
rect 5415 34229 5444 34267
rect 5444 34229 5471 34267
rect 5495 34229 5551 34285
rect 4775 34203 4831 34204
rect 4855 34203 4911 34204
rect 4935 34203 4991 34204
rect 5015 34203 5071 34204
rect 5095 34203 5151 34204
rect 5175 34203 5231 34204
rect 5255 34203 5311 34204
rect 5335 34203 5391 34204
rect 5415 34203 5471 34204
rect 4775 34151 4784 34203
rect 4784 34151 4798 34203
rect 4798 34151 4831 34203
rect 4855 34151 4864 34203
rect 4864 34151 4911 34203
rect 4935 34151 4982 34203
rect 4982 34151 4991 34203
rect 5015 34151 5048 34203
rect 5048 34151 5062 34203
rect 5062 34151 5071 34203
rect 5095 34151 5114 34203
rect 5114 34151 5128 34203
rect 5128 34151 5151 34203
rect 5175 34151 5180 34203
rect 5180 34151 5194 34203
rect 5194 34151 5231 34203
rect 5255 34151 5260 34203
rect 5260 34151 5311 34203
rect 5335 34151 5378 34203
rect 5378 34151 5391 34203
rect 5415 34151 5444 34203
rect 5444 34151 5471 34203
rect 4775 34148 4831 34151
rect 4855 34148 4911 34151
rect 4935 34148 4991 34151
rect 5015 34148 5071 34151
rect 5095 34148 5151 34151
rect 5175 34148 5231 34151
rect 5255 34148 5311 34151
rect 5335 34148 5391 34151
rect 5415 34148 5471 34151
rect 5495 34148 5551 34204
rect 4775 34087 4784 34123
rect 4784 34087 4798 34123
rect 4798 34087 4831 34123
rect 4855 34087 4864 34123
rect 4864 34087 4911 34123
rect 4935 34087 4982 34123
rect 4982 34087 4991 34123
rect 5015 34087 5048 34123
rect 5048 34087 5062 34123
rect 5062 34087 5071 34123
rect 5095 34087 5114 34123
rect 5114 34087 5128 34123
rect 5128 34087 5151 34123
rect 5175 34087 5180 34123
rect 5180 34087 5194 34123
rect 5194 34087 5231 34123
rect 5255 34087 5260 34123
rect 5260 34087 5311 34123
rect 5335 34087 5378 34123
rect 5378 34087 5391 34123
rect 5415 34087 5444 34123
rect 5444 34087 5471 34123
rect 4775 34075 4831 34087
rect 4855 34075 4911 34087
rect 4935 34075 4991 34087
rect 5015 34075 5071 34087
rect 5095 34075 5151 34087
rect 5175 34075 5231 34087
rect 5255 34075 5311 34087
rect 5335 34075 5391 34087
rect 5415 34075 5471 34087
rect 4775 34067 4784 34075
rect 4784 34067 4798 34075
rect 4798 34067 4831 34075
rect 4855 34067 4864 34075
rect 4864 34067 4911 34075
rect 4775 34023 4784 34042
rect 4784 34023 4798 34042
rect 4798 34023 4831 34042
rect 4855 34023 4864 34042
rect 4864 34023 4911 34042
rect 4935 34067 4982 34075
rect 4982 34067 4991 34075
rect 5015 34067 5048 34075
rect 5048 34067 5062 34075
rect 5062 34067 5071 34075
rect 5095 34067 5114 34075
rect 5114 34067 5128 34075
rect 5128 34067 5151 34075
rect 5175 34067 5180 34075
rect 5180 34067 5194 34075
rect 5194 34067 5231 34075
rect 5255 34067 5260 34075
rect 5260 34067 5311 34075
rect 4935 34023 4982 34042
rect 4982 34023 4991 34042
rect 5015 34023 5048 34042
rect 5048 34023 5062 34042
rect 5062 34023 5071 34042
rect 5095 34023 5114 34042
rect 5114 34023 5128 34042
rect 5128 34023 5151 34042
rect 5175 34023 5180 34042
rect 5180 34023 5194 34042
rect 5194 34023 5231 34042
rect 5255 34023 5260 34042
rect 5260 34023 5311 34042
rect 5335 34067 5378 34075
rect 5378 34067 5391 34075
rect 5415 34067 5444 34075
rect 5444 34067 5471 34075
rect 5495 34067 5551 34123
rect 5335 34023 5378 34042
rect 5378 34023 5391 34042
rect 5415 34023 5444 34042
rect 5444 34023 5471 34042
rect 4775 34011 4831 34023
rect 4855 34011 4911 34023
rect 4935 34011 4991 34023
rect 5015 34011 5071 34023
rect 5095 34011 5151 34023
rect 5175 34011 5231 34023
rect 5255 34011 5311 34023
rect 5335 34011 5391 34023
rect 5415 34011 5471 34023
rect 4775 33986 4784 34011
rect 4784 33986 4798 34011
rect 4798 33986 4831 34011
rect 4855 33986 4864 34011
rect 4864 33986 4911 34011
rect 4775 33959 4784 33961
rect 4784 33959 4798 33961
rect 4798 33959 4831 33961
rect 4855 33959 4864 33961
rect 4864 33959 4911 33961
rect 4935 33986 4982 34011
rect 4982 33986 4991 34011
rect 5015 33986 5048 34011
rect 5048 33986 5062 34011
rect 5062 33986 5071 34011
rect 5095 33986 5114 34011
rect 5114 33986 5128 34011
rect 5128 33986 5151 34011
rect 5175 33986 5180 34011
rect 5180 33986 5194 34011
rect 5194 33986 5231 34011
rect 5255 33986 5260 34011
rect 5260 33986 5311 34011
rect 4935 33959 4982 33961
rect 4982 33959 4991 33961
rect 5015 33959 5048 33961
rect 5048 33959 5062 33961
rect 5062 33959 5071 33961
rect 5095 33959 5114 33961
rect 5114 33959 5128 33961
rect 5128 33959 5151 33961
rect 5175 33959 5180 33961
rect 5180 33959 5194 33961
rect 5194 33959 5231 33961
rect 5255 33959 5260 33961
rect 5260 33959 5311 33961
rect 5335 33986 5378 34011
rect 5378 33986 5391 34011
rect 5415 33986 5444 34011
rect 5444 33986 5471 34011
rect 5495 33986 5551 34042
rect 5335 33959 5378 33961
rect 5378 33959 5391 33961
rect 5415 33959 5444 33961
rect 5444 33959 5471 33961
rect 4775 33947 4831 33959
rect 4855 33947 4911 33959
rect 4935 33947 4991 33959
rect 5015 33947 5071 33959
rect 5095 33947 5151 33959
rect 5175 33947 5231 33959
rect 5255 33947 5311 33959
rect 5335 33947 5391 33959
rect 5415 33947 5471 33959
rect 4775 33905 4784 33947
rect 4784 33905 4798 33947
rect 4798 33905 4831 33947
rect 4855 33905 4864 33947
rect 4864 33905 4911 33947
rect 4935 33905 4982 33947
rect 4982 33905 4991 33947
rect 5015 33905 5048 33947
rect 5048 33905 5062 33947
rect 5062 33905 5071 33947
rect 5095 33905 5114 33947
rect 5114 33905 5128 33947
rect 5128 33905 5151 33947
rect 5175 33905 5180 33947
rect 5180 33905 5194 33947
rect 5194 33905 5231 33947
rect 5255 33905 5260 33947
rect 5260 33905 5311 33947
rect 5335 33905 5378 33947
rect 5378 33905 5391 33947
rect 5415 33905 5444 33947
rect 5444 33905 5471 33947
rect 5495 33905 5551 33961
rect 4775 33831 4784 33880
rect 4784 33831 4798 33880
rect 4798 33831 4831 33880
rect 4855 33831 4864 33880
rect 4864 33831 4911 33880
rect 4935 33831 4982 33880
rect 4982 33831 4991 33880
rect 5015 33831 5048 33880
rect 5048 33831 5062 33880
rect 5062 33831 5071 33880
rect 5095 33831 5114 33880
rect 5114 33831 5128 33880
rect 5128 33831 5151 33880
rect 5175 33831 5180 33880
rect 5180 33831 5194 33880
rect 5194 33831 5231 33880
rect 5255 33831 5260 33880
rect 5260 33831 5311 33880
rect 5335 33831 5378 33880
rect 5378 33831 5391 33880
rect 5415 33831 5444 33880
rect 5444 33831 5471 33880
rect 4775 33824 4831 33831
rect 4855 33824 4911 33831
rect 4935 33824 4991 33831
rect 5015 33824 5071 33831
rect 5095 33824 5151 33831
rect 5175 33824 5231 33831
rect 5255 33824 5311 33831
rect 5335 33824 5391 33831
rect 5415 33824 5471 33831
rect 5495 33824 5551 33880
rect 4775 33767 4784 33799
rect 4784 33767 4798 33799
rect 4798 33767 4831 33799
rect 4855 33767 4864 33799
rect 4864 33767 4911 33799
rect 4935 33767 4982 33799
rect 4982 33767 4991 33799
rect 5015 33767 5048 33799
rect 5048 33767 5062 33799
rect 5062 33767 5071 33799
rect 5095 33767 5114 33799
rect 5114 33767 5128 33799
rect 5128 33767 5151 33799
rect 5175 33767 5180 33799
rect 5180 33767 5194 33799
rect 5194 33767 5231 33799
rect 5255 33767 5260 33799
rect 5260 33767 5311 33799
rect 5335 33767 5378 33799
rect 5378 33767 5391 33799
rect 5415 33767 5444 33799
rect 5444 33767 5471 33799
rect 4775 33755 4831 33767
rect 4855 33755 4911 33767
rect 4935 33755 4991 33767
rect 5015 33755 5071 33767
rect 5095 33755 5151 33767
rect 5175 33755 5231 33767
rect 5255 33755 5311 33767
rect 5335 33755 5391 33767
rect 5415 33755 5471 33767
rect 4775 33743 4784 33755
rect 4784 33743 4798 33755
rect 4798 33743 4831 33755
rect 4855 33743 4864 33755
rect 4864 33743 4911 33755
rect 4775 33703 4784 33718
rect 4784 33703 4798 33718
rect 4798 33703 4831 33718
rect 4855 33703 4864 33718
rect 4864 33703 4911 33718
rect 4935 33743 4982 33755
rect 4982 33743 4991 33755
rect 5015 33743 5048 33755
rect 5048 33743 5062 33755
rect 5062 33743 5071 33755
rect 5095 33743 5114 33755
rect 5114 33743 5128 33755
rect 5128 33743 5151 33755
rect 5175 33743 5180 33755
rect 5180 33743 5194 33755
rect 5194 33743 5231 33755
rect 5255 33743 5260 33755
rect 5260 33743 5311 33755
rect 4935 33703 4982 33718
rect 4982 33703 4991 33718
rect 5015 33703 5048 33718
rect 5048 33703 5062 33718
rect 5062 33703 5071 33718
rect 5095 33703 5114 33718
rect 5114 33703 5128 33718
rect 5128 33703 5151 33718
rect 5175 33703 5180 33718
rect 5180 33703 5194 33718
rect 5194 33703 5231 33718
rect 5255 33703 5260 33718
rect 5260 33703 5311 33718
rect 5335 33743 5378 33755
rect 5378 33743 5391 33755
rect 5415 33743 5444 33755
rect 5444 33743 5471 33755
rect 5495 33743 5551 33799
rect 5335 33703 5378 33718
rect 5378 33703 5391 33718
rect 5415 33703 5444 33718
rect 5444 33703 5471 33718
rect 4775 33691 4831 33703
rect 4855 33691 4911 33703
rect 4935 33691 4991 33703
rect 5015 33691 5071 33703
rect 5095 33691 5151 33703
rect 5175 33691 5231 33703
rect 5255 33691 5311 33703
rect 5335 33691 5391 33703
rect 5415 33691 5471 33703
rect 4775 33662 4784 33691
rect 4784 33662 4798 33691
rect 4798 33662 4831 33691
rect 4855 33662 4864 33691
rect 4864 33662 4911 33691
rect 4935 33662 4982 33691
rect 4982 33662 4991 33691
rect 5015 33662 5048 33691
rect 5048 33662 5062 33691
rect 5062 33662 5071 33691
rect 5095 33662 5114 33691
rect 5114 33662 5128 33691
rect 5128 33662 5151 33691
rect 5175 33662 5180 33691
rect 5180 33662 5194 33691
rect 5194 33662 5231 33691
rect 5255 33662 5260 33691
rect 5260 33662 5311 33691
rect 5335 33662 5378 33691
rect 5378 33662 5391 33691
rect 5415 33662 5444 33691
rect 5444 33662 5471 33691
rect 5495 33662 5551 33718
rect 4775 33627 4831 33637
rect 4855 33627 4911 33637
rect 4935 33627 4991 33637
rect 5015 33627 5071 33637
rect 5095 33627 5151 33637
rect 5175 33627 5231 33637
rect 5255 33627 5311 33637
rect 5335 33627 5391 33637
rect 5415 33627 5471 33637
rect 4775 33581 4784 33627
rect 4784 33581 4798 33627
rect 4798 33581 4831 33627
rect 4855 33581 4864 33627
rect 4864 33581 4911 33627
rect 4935 33581 4982 33627
rect 4982 33581 4991 33627
rect 5015 33581 5048 33627
rect 5048 33581 5062 33627
rect 5062 33581 5071 33627
rect 5095 33581 5114 33627
rect 5114 33581 5128 33627
rect 5128 33581 5151 33627
rect 5175 33581 5180 33627
rect 5180 33581 5194 33627
rect 5194 33581 5231 33627
rect 5255 33581 5260 33627
rect 5260 33581 5311 33627
rect 5335 33581 5378 33627
rect 5378 33581 5391 33627
rect 5415 33581 5444 33627
rect 5444 33581 5471 33627
rect 5495 33581 5551 33637
rect 4775 33511 4784 33556
rect 4784 33511 4798 33556
rect 4798 33511 4831 33556
rect 4855 33511 4864 33556
rect 4864 33511 4911 33556
rect 4935 33511 4982 33556
rect 4982 33511 4991 33556
rect 5015 33511 5048 33556
rect 5048 33511 5062 33556
rect 5062 33511 5071 33556
rect 5095 33511 5114 33556
rect 5114 33511 5128 33556
rect 5128 33511 5151 33556
rect 5175 33511 5180 33556
rect 5180 33511 5194 33556
rect 5194 33511 5231 33556
rect 5255 33511 5260 33556
rect 5260 33511 5311 33556
rect 5335 33511 5378 33556
rect 5378 33511 5391 33556
rect 5415 33511 5444 33556
rect 5444 33511 5471 33556
rect 4775 33500 4831 33511
rect 4855 33500 4911 33511
rect 4935 33500 4991 33511
rect 5015 33500 5071 33511
rect 5095 33500 5151 33511
rect 5175 33500 5231 33511
rect 5255 33500 5311 33511
rect 5335 33500 5391 33511
rect 5415 33500 5471 33511
rect 5495 33500 5551 33556
rect 4775 33447 4784 33475
rect 4784 33447 4798 33475
rect 4798 33447 4831 33475
rect 4855 33447 4864 33475
rect 4864 33447 4911 33475
rect 4935 33447 4982 33475
rect 4982 33447 4991 33475
rect 5015 33447 5048 33475
rect 5048 33447 5062 33475
rect 5062 33447 5071 33475
rect 5095 33447 5114 33475
rect 5114 33447 5128 33475
rect 5128 33447 5151 33475
rect 5175 33447 5180 33475
rect 5180 33447 5194 33475
rect 5194 33447 5231 33475
rect 5255 33447 5260 33475
rect 5260 33447 5311 33475
rect 5335 33447 5378 33475
rect 5378 33447 5391 33475
rect 5415 33447 5444 33475
rect 5444 33447 5471 33475
rect 4775 33435 4831 33447
rect 4855 33435 4911 33447
rect 4935 33435 4991 33447
rect 5015 33435 5071 33447
rect 5095 33435 5151 33447
rect 5175 33435 5231 33447
rect 5255 33435 5311 33447
rect 5335 33435 5391 33447
rect 5415 33435 5471 33447
rect 4775 33419 4784 33435
rect 4784 33419 4798 33435
rect 4798 33419 4831 33435
rect 4855 33419 4864 33435
rect 4864 33419 4911 33435
rect 4775 33383 4784 33394
rect 4784 33383 4798 33394
rect 4798 33383 4831 33394
rect 4855 33383 4864 33394
rect 4864 33383 4911 33394
rect 4935 33419 4982 33435
rect 4982 33419 4991 33435
rect 5015 33419 5048 33435
rect 5048 33419 5062 33435
rect 5062 33419 5071 33435
rect 5095 33419 5114 33435
rect 5114 33419 5128 33435
rect 5128 33419 5151 33435
rect 5175 33419 5180 33435
rect 5180 33419 5194 33435
rect 5194 33419 5231 33435
rect 5255 33419 5260 33435
rect 5260 33419 5311 33435
rect 4935 33383 4982 33394
rect 4982 33383 4991 33394
rect 5015 33383 5048 33394
rect 5048 33383 5062 33394
rect 5062 33383 5071 33394
rect 5095 33383 5114 33394
rect 5114 33383 5128 33394
rect 5128 33383 5151 33394
rect 5175 33383 5180 33394
rect 5180 33383 5194 33394
rect 5194 33383 5231 33394
rect 5255 33383 5260 33394
rect 5260 33383 5311 33394
rect 5335 33419 5378 33435
rect 5378 33419 5391 33435
rect 5415 33419 5444 33435
rect 5444 33419 5471 33435
rect 5495 33419 5551 33475
rect 5335 33383 5378 33394
rect 5378 33383 5391 33394
rect 5415 33383 5444 33394
rect 5444 33383 5471 33394
rect 4775 33371 4831 33383
rect 4855 33371 4911 33383
rect 4935 33371 4991 33383
rect 5015 33371 5071 33383
rect 5095 33371 5151 33383
rect 5175 33371 5231 33383
rect 5255 33371 5311 33383
rect 5335 33371 5391 33383
rect 5415 33371 5471 33383
rect 4775 33338 4784 33371
rect 4784 33338 4798 33371
rect 4798 33338 4831 33371
rect 4855 33338 4864 33371
rect 4864 33338 4911 33371
rect 4935 33338 4982 33371
rect 4982 33338 4991 33371
rect 5015 33338 5048 33371
rect 5048 33338 5062 33371
rect 5062 33338 5071 33371
rect 5095 33338 5114 33371
rect 5114 33338 5128 33371
rect 5128 33338 5151 33371
rect 5175 33338 5180 33371
rect 5180 33338 5194 33371
rect 5194 33338 5231 33371
rect 5255 33338 5260 33371
rect 5260 33338 5311 33371
rect 5335 33338 5378 33371
rect 5378 33338 5391 33371
rect 5415 33338 5444 33371
rect 5444 33338 5471 33371
rect 5495 33338 5551 33394
rect 4775 33307 4831 33313
rect 4855 33307 4911 33313
rect 4935 33307 4991 33313
rect 5015 33307 5071 33313
rect 5095 33307 5151 33313
rect 5175 33307 5231 33313
rect 5255 33307 5311 33313
rect 5335 33307 5391 33313
rect 5415 33307 5471 33313
rect 4775 33257 4784 33307
rect 4784 33257 4798 33307
rect 4798 33257 4831 33307
rect 4855 33257 4864 33307
rect 4864 33257 4911 33307
rect 4935 33257 4982 33307
rect 4982 33257 4991 33307
rect 5015 33257 5048 33307
rect 5048 33257 5062 33307
rect 5062 33257 5071 33307
rect 5095 33257 5114 33307
rect 5114 33257 5128 33307
rect 5128 33257 5151 33307
rect 5175 33257 5180 33307
rect 5180 33257 5194 33307
rect 5194 33257 5231 33307
rect 5255 33257 5260 33307
rect 5260 33257 5311 33307
rect 5335 33257 5378 33307
rect 5378 33257 5391 33307
rect 5415 33257 5444 33307
rect 5444 33257 5471 33307
rect 5495 33257 5551 33313
rect 4775 33191 4784 33232
rect 4784 33191 4798 33232
rect 4798 33191 4831 33232
rect 4855 33191 4864 33232
rect 4864 33191 4911 33232
rect 4935 33191 4982 33232
rect 4982 33191 4991 33232
rect 5015 33191 5048 33232
rect 5048 33191 5062 33232
rect 5062 33191 5071 33232
rect 5095 33191 5114 33232
rect 5114 33191 5128 33232
rect 5128 33191 5151 33232
rect 5175 33191 5180 33232
rect 5180 33191 5194 33232
rect 5194 33191 5231 33232
rect 5255 33191 5260 33232
rect 5260 33191 5311 33232
rect 5335 33191 5378 33232
rect 5378 33191 5391 33232
rect 5415 33191 5444 33232
rect 5444 33191 5471 33232
rect 4775 33179 4831 33191
rect 4855 33179 4911 33191
rect 4935 33179 4991 33191
rect 5015 33179 5071 33191
rect 5095 33179 5151 33191
rect 5175 33179 5231 33191
rect 5255 33179 5311 33191
rect 5335 33179 5391 33191
rect 5415 33179 5471 33191
rect 4775 33176 4784 33179
rect 4784 33176 4798 33179
rect 4798 33176 4831 33179
rect 4855 33176 4864 33179
rect 4864 33176 4911 33179
rect 4775 33127 4784 33151
rect 4784 33127 4798 33151
rect 4798 33127 4831 33151
rect 4855 33127 4864 33151
rect 4864 33127 4911 33151
rect 4935 33176 4982 33179
rect 4982 33176 4991 33179
rect 5015 33176 5048 33179
rect 5048 33176 5062 33179
rect 5062 33176 5071 33179
rect 5095 33176 5114 33179
rect 5114 33176 5128 33179
rect 5128 33176 5151 33179
rect 5175 33176 5180 33179
rect 5180 33176 5194 33179
rect 5194 33176 5231 33179
rect 5255 33176 5260 33179
rect 5260 33176 5311 33179
rect 4935 33127 4982 33151
rect 4982 33127 4991 33151
rect 5015 33127 5048 33151
rect 5048 33127 5062 33151
rect 5062 33127 5071 33151
rect 5095 33127 5114 33151
rect 5114 33127 5128 33151
rect 5128 33127 5151 33151
rect 5175 33127 5180 33151
rect 5180 33127 5194 33151
rect 5194 33127 5231 33151
rect 5255 33127 5260 33151
rect 5260 33127 5311 33151
rect 5335 33176 5378 33179
rect 5378 33176 5391 33179
rect 5415 33176 5444 33179
rect 5444 33176 5471 33179
rect 5495 33176 5551 33232
rect 5335 33127 5378 33151
rect 5378 33127 5391 33151
rect 5415 33127 5444 33151
rect 5444 33127 5471 33151
rect 4775 33115 4831 33127
rect 4855 33115 4911 33127
rect 4935 33115 4991 33127
rect 5015 33115 5071 33127
rect 5095 33115 5151 33127
rect 5175 33115 5231 33127
rect 5255 33115 5311 33127
rect 5335 33115 5391 33127
rect 5415 33115 5471 33127
rect 4775 33095 4784 33115
rect 4784 33095 4798 33115
rect 4798 33095 4831 33115
rect 4855 33095 4864 33115
rect 4864 33095 4911 33115
rect 4775 33063 4784 33070
rect 4784 33063 4798 33070
rect 4798 33063 4831 33070
rect 4855 33063 4864 33070
rect 4864 33063 4911 33070
rect 4935 33095 4982 33115
rect 4982 33095 4991 33115
rect 5015 33095 5048 33115
rect 5048 33095 5062 33115
rect 5062 33095 5071 33115
rect 5095 33095 5114 33115
rect 5114 33095 5128 33115
rect 5128 33095 5151 33115
rect 5175 33095 5180 33115
rect 5180 33095 5194 33115
rect 5194 33095 5231 33115
rect 5255 33095 5260 33115
rect 5260 33095 5311 33115
rect 4935 33063 4982 33070
rect 4982 33063 4991 33070
rect 5015 33063 5048 33070
rect 5048 33063 5062 33070
rect 5062 33063 5071 33070
rect 5095 33063 5114 33070
rect 5114 33063 5128 33070
rect 5128 33063 5151 33070
rect 5175 33063 5180 33070
rect 5180 33063 5194 33070
rect 5194 33063 5231 33070
rect 5255 33063 5260 33070
rect 5260 33063 5311 33070
rect 5335 33095 5378 33115
rect 5378 33095 5391 33115
rect 5415 33095 5444 33115
rect 5444 33095 5471 33115
rect 5495 33095 5551 33151
rect 5335 33063 5378 33070
rect 5378 33063 5391 33070
rect 5415 33063 5444 33070
rect 5444 33063 5471 33070
rect 4775 33051 4831 33063
rect 4855 33051 4911 33063
rect 4935 33051 4991 33063
rect 5015 33051 5071 33063
rect 5095 33051 5151 33063
rect 5175 33051 5231 33063
rect 5255 33051 5311 33063
rect 5335 33051 5391 33063
rect 5415 33051 5471 33063
rect 4775 33014 4784 33051
rect 4784 33014 4798 33051
rect 4798 33014 4831 33051
rect 4855 33014 4864 33051
rect 4864 33014 4911 33051
rect 4935 33014 4982 33051
rect 4982 33014 4991 33051
rect 5015 33014 5048 33051
rect 5048 33014 5062 33051
rect 5062 33014 5071 33051
rect 5095 33014 5114 33051
rect 5114 33014 5128 33051
rect 5128 33014 5151 33051
rect 5175 33014 5180 33051
rect 5180 33014 5194 33051
rect 5194 33014 5231 33051
rect 5255 33014 5260 33051
rect 5260 33014 5311 33051
rect 5335 33014 5378 33051
rect 5378 33014 5391 33051
rect 5415 33014 5444 33051
rect 5444 33014 5471 33051
rect 5495 33014 5551 33070
rect 4775 32987 4831 32989
rect 4855 32987 4911 32989
rect 4935 32987 4991 32989
rect 5015 32987 5071 32989
rect 5095 32987 5151 32989
rect 5175 32987 5231 32989
rect 5255 32987 5311 32989
rect 5335 32987 5391 32989
rect 5415 32987 5471 32989
rect 4775 32935 4784 32987
rect 4784 32935 4798 32987
rect 4798 32935 4831 32987
rect 4855 32935 4864 32987
rect 4864 32935 4911 32987
rect 4935 32935 4982 32987
rect 4982 32935 4991 32987
rect 5015 32935 5048 32987
rect 5048 32935 5062 32987
rect 5062 32935 5071 32987
rect 5095 32935 5114 32987
rect 5114 32935 5128 32987
rect 5128 32935 5151 32987
rect 5175 32935 5180 32987
rect 5180 32935 5194 32987
rect 5194 32935 5231 32987
rect 5255 32935 5260 32987
rect 5260 32935 5311 32987
rect 5335 32935 5378 32987
rect 5378 32935 5391 32987
rect 5415 32935 5444 32987
rect 5444 32935 5471 32987
rect 4775 32933 4831 32935
rect 4855 32933 4911 32935
rect 4935 32933 4991 32935
rect 5015 32933 5071 32935
rect 5095 32933 5151 32935
rect 5175 32933 5231 32935
rect 5255 32933 5311 32935
rect 5335 32933 5391 32935
rect 5415 32933 5471 32935
rect 5495 32933 5551 32989
rect 4775 32871 4784 32908
rect 4784 32871 4798 32908
rect 4798 32871 4831 32908
rect 4855 32871 4864 32908
rect 4864 32871 4911 32908
rect 4935 32871 4982 32908
rect 4982 32871 4991 32908
rect 5015 32871 5048 32908
rect 5048 32871 5062 32908
rect 5062 32871 5071 32908
rect 5095 32871 5114 32908
rect 5114 32871 5128 32908
rect 5128 32871 5151 32908
rect 5175 32871 5180 32908
rect 5180 32871 5194 32908
rect 5194 32871 5231 32908
rect 5255 32871 5260 32908
rect 5260 32871 5311 32908
rect 5335 32871 5378 32908
rect 5378 32871 5391 32908
rect 5415 32871 5444 32908
rect 5444 32871 5471 32908
rect 4775 32859 4831 32871
rect 4855 32859 4911 32871
rect 4935 32859 4991 32871
rect 5015 32859 5071 32871
rect 5095 32859 5151 32871
rect 5175 32859 5231 32871
rect 5255 32859 5311 32871
rect 5335 32859 5391 32871
rect 5415 32859 5471 32871
rect 4775 32852 4784 32859
rect 4784 32852 4798 32859
rect 4798 32852 4831 32859
rect 4855 32852 4864 32859
rect 4864 32852 4911 32859
rect 4775 32807 4784 32827
rect 4784 32807 4798 32827
rect 4798 32807 4831 32827
rect 4855 32807 4864 32827
rect 4864 32807 4911 32827
rect 4935 32852 4982 32859
rect 4982 32852 4991 32859
rect 5015 32852 5048 32859
rect 5048 32852 5062 32859
rect 5062 32852 5071 32859
rect 5095 32852 5114 32859
rect 5114 32852 5128 32859
rect 5128 32852 5151 32859
rect 5175 32852 5180 32859
rect 5180 32852 5194 32859
rect 5194 32852 5231 32859
rect 5255 32852 5260 32859
rect 5260 32852 5311 32859
rect 4935 32807 4982 32827
rect 4982 32807 4991 32827
rect 5015 32807 5048 32827
rect 5048 32807 5062 32827
rect 5062 32807 5071 32827
rect 5095 32807 5114 32827
rect 5114 32807 5128 32827
rect 5128 32807 5151 32827
rect 5175 32807 5180 32827
rect 5180 32807 5194 32827
rect 5194 32807 5231 32827
rect 5255 32807 5260 32827
rect 5260 32807 5311 32827
rect 5335 32852 5378 32859
rect 5378 32852 5391 32859
rect 5415 32852 5444 32859
rect 5444 32852 5471 32859
rect 5495 32852 5551 32908
rect 5335 32807 5378 32827
rect 5378 32807 5391 32827
rect 5415 32807 5444 32827
rect 5444 32807 5471 32827
rect 4775 32795 4831 32807
rect 4855 32795 4911 32807
rect 4935 32795 4991 32807
rect 5015 32795 5071 32807
rect 5095 32795 5151 32807
rect 5175 32795 5231 32807
rect 5255 32795 5311 32807
rect 5335 32795 5391 32807
rect 5415 32795 5471 32807
rect 4775 32771 4784 32795
rect 4784 32771 4798 32795
rect 4798 32771 4831 32795
rect 4855 32771 4864 32795
rect 4864 32771 4911 32795
rect 4775 32743 4784 32746
rect 4784 32743 4798 32746
rect 4798 32743 4831 32746
rect 4855 32743 4864 32746
rect 4864 32743 4911 32746
rect 4935 32771 4982 32795
rect 4982 32771 4991 32795
rect 5015 32771 5048 32795
rect 5048 32771 5062 32795
rect 5062 32771 5071 32795
rect 5095 32771 5114 32795
rect 5114 32771 5128 32795
rect 5128 32771 5151 32795
rect 5175 32771 5180 32795
rect 5180 32771 5194 32795
rect 5194 32771 5231 32795
rect 5255 32771 5260 32795
rect 5260 32771 5311 32795
rect 4935 32743 4982 32746
rect 4982 32743 4991 32746
rect 5015 32743 5048 32746
rect 5048 32743 5062 32746
rect 5062 32743 5071 32746
rect 5095 32743 5114 32746
rect 5114 32743 5128 32746
rect 5128 32743 5151 32746
rect 5175 32743 5180 32746
rect 5180 32743 5194 32746
rect 5194 32743 5231 32746
rect 5255 32743 5260 32746
rect 5260 32743 5311 32746
rect 5335 32771 5378 32795
rect 5378 32771 5391 32795
rect 5415 32771 5444 32795
rect 5444 32771 5471 32795
rect 5495 32771 5551 32827
rect 5335 32743 5378 32746
rect 5378 32743 5391 32746
rect 5415 32743 5444 32746
rect 5444 32743 5471 32746
rect 4775 32730 4831 32743
rect 4855 32730 4911 32743
rect 4935 32730 4991 32743
rect 5015 32730 5071 32743
rect 5095 32730 5151 32743
rect 5175 32730 5231 32743
rect 5255 32730 5311 32743
rect 5335 32730 5391 32743
rect 5415 32730 5471 32743
rect 4775 32690 4784 32730
rect 4784 32690 4798 32730
rect 4798 32690 4831 32730
rect 4855 32690 4864 32730
rect 4864 32690 4911 32730
rect 4935 32690 4982 32730
rect 4982 32690 4991 32730
rect 5015 32690 5048 32730
rect 5048 32690 5062 32730
rect 5062 32690 5071 32730
rect 5095 32690 5114 32730
rect 5114 32690 5128 32730
rect 5128 32690 5151 32730
rect 5175 32690 5180 32730
rect 5180 32690 5194 32730
rect 5194 32690 5231 32730
rect 5255 32690 5260 32730
rect 5260 32690 5311 32730
rect 5335 32690 5378 32730
rect 5378 32690 5391 32730
rect 5415 32690 5444 32730
rect 5444 32690 5471 32730
rect 5495 32690 5551 32746
rect 4775 32613 4784 32665
rect 4784 32613 4798 32665
rect 4798 32613 4831 32665
rect 4855 32613 4864 32665
rect 4864 32613 4911 32665
rect 4935 32613 4982 32665
rect 4982 32613 4991 32665
rect 5015 32613 5048 32665
rect 5048 32613 5062 32665
rect 5062 32613 5071 32665
rect 5095 32613 5114 32665
rect 5114 32613 5128 32665
rect 5128 32613 5151 32665
rect 5175 32613 5180 32665
rect 5180 32613 5194 32665
rect 5194 32613 5231 32665
rect 5255 32613 5260 32665
rect 5260 32613 5311 32665
rect 5335 32613 5378 32665
rect 5378 32613 5391 32665
rect 5415 32613 5444 32665
rect 5444 32613 5471 32665
rect 4775 32609 4831 32613
rect 4855 32609 4911 32613
rect 4935 32609 4991 32613
rect 5015 32609 5071 32613
rect 5095 32609 5151 32613
rect 5175 32609 5231 32613
rect 5255 32609 5311 32613
rect 5335 32609 5391 32613
rect 5415 32609 5471 32613
rect 5495 32609 5551 32665
rect 4775 32548 4784 32584
rect 4784 32548 4798 32584
rect 4798 32548 4831 32584
rect 4855 32548 4864 32584
rect 4864 32548 4911 32584
rect 4935 32548 4982 32584
rect 4982 32548 4991 32584
rect 5015 32548 5048 32584
rect 5048 32548 5062 32584
rect 5062 32548 5071 32584
rect 5095 32548 5114 32584
rect 5114 32548 5128 32584
rect 5128 32548 5151 32584
rect 5175 32548 5180 32584
rect 5180 32548 5194 32584
rect 5194 32548 5231 32584
rect 5255 32548 5260 32584
rect 5260 32548 5311 32584
rect 5335 32548 5378 32584
rect 5378 32548 5391 32584
rect 5415 32548 5444 32584
rect 5444 32548 5471 32584
rect 4775 32535 4831 32548
rect 4855 32535 4911 32548
rect 4935 32535 4991 32548
rect 5015 32535 5071 32548
rect 5095 32535 5151 32548
rect 5175 32535 5231 32548
rect 5255 32535 5311 32548
rect 5335 32535 5391 32548
rect 5415 32535 5471 32548
rect 4775 32528 4784 32535
rect 4784 32528 4798 32535
rect 4798 32528 4831 32535
rect 4855 32528 4864 32535
rect 4864 32528 4911 32535
rect 4775 32483 4784 32503
rect 4784 32483 4798 32503
rect 4798 32483 4831 32503
rect 4855 32483 4864 32503
rect 4864 32483 4911 32503
rect 4935 32528 4982 32535
rect 4982 32528 4991 32535
rect 5015 32528 5048 32535
rect 5048 32528 5062 32535
rect 5062 32528 5071 32535
rect 5095 32528 5114 32535
rect 5114 32528 5128 32535
rect 5128 32528 5151 32535
rect 5175 32528 5180 32535
rect 5180 32528 5194 32535
rect 5194 32528 5231 32535
rect 5255 32528 5260 32535
rect 5260 32528 5311 32535
rect 4935 32483 4982 32503
rect 4982 32483 4991 32503
rect 5015 32483 5048 32503
rect 5048 32483 5062 32503
rect 5062 32483 5071 32503
rect 5095 32483 5114 32503
rect 5114 32483 5128 32503
rect 5128 32483 5151 32503
rect 5175 32483 5180 32503
rect 5180 32483 5194 32503
rect 5194 32483 5231 32503
rect 5255 32483 5260 32503
rect 5260 32483 5311 32503
rect 5335 32528 5378 32535
rect 5378 32528 5391 32535
rect 5415 32528 5444 32535
rect 5444 32528 5471 32535
rect 5495 32528 5551 32584
rect 5335 32483 5378 32503
rect 5378 32483 5391 32503
rect 5415 32483 5444 32503
rect 5444 32483 5471 32503
rect 4775 32470 4831 32483
rect 4855 32470 4911 32483
rect 4935 32470 4991 32483
rect 5015 32470 5071 32483
rect 5095 32470 5151 32483
rect 5175 32470 5231 32483
rect 5255 32470 5311 32483
rect 5335 32470 5391 32483
rect 5415 32470 5471 32483
rect 4775 32447 4784 32470
rect 4784 32447 4798 32470
rect 4798 32447 4831 32470
rect 4855 32447 4864 32470
rect 4864 32447 4911 32470
rect 4775 32418 4784 32422
rect 4784 32418 4798 32422
rect 4798 32418 4831 32422
rect 4855 32418 4864 32422
rect 4864 32418 4911 32422
rect 4935 32447 4982 32470
rect 4982 32447 4991 32470
rect 5015 32447 5048 32470
rect 5048 32447 5062 32470
rect 5062 32447 5071 32470
rect 5095 32447 5114 32470
rect 5114 32447 5128 32470
rect 5128 32447 5151 32470
rect 5175 32447 5180 32470
rect 5180 32447 5194 32470
rect 5194 32447 5231 32470
rect 5255 32447 5260 32470
rect 5260 32447 5311 32470
rect 4935 32418 4982 32422
rect 4982 32418 4991 32422
rect 5015 32418 5048 32422
rect 5048 32418 5062 32422
rect 5062 32418 5071 32422
rect 5095 32418 5114 32422
rect 5114 32418 5128 32422
rect 5128 32418 5151 32422
rect 5175 32418 5180 32422
rect 5180 32418 5194 32422
rect 5194 32418 5231 32422
rect 5255 32418 5260 32422
rect 5260 32418 5311 32422
rect 5335 32447 5378 32470
rect 5378 32447 5391 32470
rect 5415 32447 5444 32470
rect 5444 32447 5471 32470
rect 5495 32447 5551 32503
rect 5335 32418 5378 32422
rect 5378 32418 5391 32422
rect 5415 32418 5444 32422
rect 5444 32418 5471 32422
rect 4775 32405 4831 32418
rect 4855 32405 4911 32418
rect 4935 32405 4991 32418
rect 5015 32405 5071 32418
rect 5095 32405 5151 32418
rect 5175 32405 5231 32418
rect 5255 32405 5311 32418
rect 5335 32405 5391 32418
rect 5415 32405 5471 32418
rect 4775 32366 4784 32405
rect 4784 32366 4798 32405
rect 4798 32366 4831 32405
rect 4855 32366 4864 32405
rect 4864 32366 4911 32405
rect 4935 32366 4982 32405
rect 4982 32366 4991 32405
rect 5015 32366 5048 32405
rect 5048 32366 5062 32405
rect 5062 32366 5071 32405
rect 5095 32366 5114 32405
rect 5114 32366 5128 32405
rect 5128 32366 5151 32405
rect 5175 32366 5180 32405
rect 5180 32366 5194 32405
rect 5194 32366 5231 32405
rect 5255 32366 5260 32405
rect 5260 32366 5311 32405
rect 5335 32366 5378 32405
rect 5378 32366 5391 32405
rect 5415 32366 5444 32405
rect 5444 32366 5471 32405
rect 5495 32366 5551 32422
rect 4775 32340 4831 32341
rect 4855 32340 4911 32341
rect 4935 32340 4991 32341
rect 5015 32340 5071 32341
rect 5095 32340 5151 32341
rect 5175 32340 5231 32341
rect 5255 32340 5311 32341
rect 5335 32340 5391 32341
rect 5415 32340 5471 32341
rect 4775 32288 4784 32340
rect 4784 32288 4798 32340
rect 4798 32288 4831 32340
rect 4855 32288 4864 32340
rect 4864 32288 4911 32340
rect 4935 32288 4982 32340
rect 4982 32288 4991 32340
rect 5015 32288 5048 32340
rect 5048 32288 5062 32340
rect 5062 32288 5071 32340
rect 5095 32288 5114 32340
rect 5114 32288 5128 32340
rect 5128 32288 5151 32340
rect 5175 32288 5180 32340
rect 5180 32288 5194 32340
rect 5194 32288 5231 32340
rect 5255 32288 5260 32340
rect 5260 32288 5311 32340
rect 5335 32288 5378 32340
rect 5378 32288 5391 32340
rect 5415 32288 5444 32340
rect 5444 32288 5471 32340
rect 4775 32285 4831 32288
rect 4855 32285 4911 32288
rect 4935 32285 4991 32288
rect 5015 32285 5071 32288
rect 5095 32285 5151 32288
rect 5175 32285 5231 32288
rect 5255 32285 5311 32288
rect 5335 32285 5391 32288
rect 5415 32285 5471 32288
rect 5495 32285 5551 32341
rect 4775 32223 4784 32260
rect 4784 32223 4798 32260
rect 4798 32223 4831 32260
rect 4855 32223 4864 32260
rect 4864 32223 4911 32260
rect 4935 32223 4982 32260
rect 4982 32223 4991 32260
rect 5015 32223 5048 32260
rect 5048 32223 5062 32260
rect 5062 32223 5071 32260
rect 5095 32223 5114 32260
rect 5114 32223 5128 32260
rect 5128 32223 5151 32260
rect 5175 32223 5180 32260
rect 5180 32223 5194 32260
rect 5194 32223 5231 32260
rect 5255 32223 5260 32260
rect 5260 32223 5311 32260
rect 5335 32223 5378 32260
rect 5378 32223 5391 32260
rect 5415 32223 5444 32260
rect 5444 32223 5471 32260
rect 4775 32210 4831 32223
rect 4855 32210 4911 32223
rect 4935 32210 4991 32223
rect 5015 32210 5071 32223
rect 5095 32210 5151 32223
rect 5175 32210 5231 32223
rect 5255 32210 5311 32223
rect 5335 32210 5391 32223
rect 5415 32210 5471 32223
rect 4775 32204 4784 32210
rect 4784 32204 4798 32210
rect 4798 32204 4831 32210
rect 4855 32204 4864 32210
rect 4864 32204 4911 32210
rect 4775 32158 4784 32179
rect 4784 32158 4798 32179
rect 4798 32158 4831 32179
rect 4855 32158 4864 32179
rect 4864 32158 4911 32179
rect 4935 32204 4982 32210
rect 4982 32204 4991 32210
rect 5015 32204 5048 32210
rect 5048 32204 5062 32210
rect 5062 32204 5071 32210
rect 5095 32204 5114 32210
rect 5114 32204 5128 32210
rect 5128 32204 5151 32210
rect 5175 32204 5180 32210
rect 5180 32204 5194 32210
rect 5194 32204 5231 32210
rect 5255 32204 5260 32210
rect 5260 32204 5311 32210
rect 4935 32158 4982 32179
rect 4982 32158 4991 32179
rect 5015 32158 5048 32179
rect 5048 32158 5062 32179
rect 5062 32158 5071 32179
rect 5095 32158 5114 32179
rect 5114 32158 5128 32179
rect 5128 32158 5151 32179
rect 5175 32158 5180 32179
rect 5180 32158 5194 32179
rect 5194 32158 5231 32179
rect 5255 32158 5260 32179
rect 5260 32158 5311 32179
rect 5335 32204 5378 32210
rect 5378 32204 5391 32210
rect 5415 32204 5444 32210
rect 5444 32204 5471 32210
rect 5495 32204 5551 32260
rect 5335 32158 5378 32179
rect 5378 32158 5391 32179
rect 5415 32158 5444 32179
rect 5444 32158 5471 32179
rect 4775 32145 4831 32158
rect 4855 32145 4911 32158
rect 4935 32145 4991 32158
rect 5015 32145 5071 32158
rect 5095 32145 5151 32158
rect 5175 32145 5231 32158
rect 5255 32145 5311 32158
rect 5335 32145 5391 32158
rect 5415 32145 5471 32158
rect 4775 32123 4784 32145
rect 4784 32123 4798 32145
rect 4798 32123 4831 32145
rect 4855 32123 4864 32145
rect 4864 32123 4911 32145
rect 4775 32093 4784 32098
rect 4784 32093 4798 32098
rect 4798 32093 4831 32098
rect 4855 32093 4864 32098
rect 4864 32093 4911 32098
rect 4935 32123 4982 32145
rect 4982 32123 4991 32145
rect 5015 32123 5048 32145
rect 5048 32123 5062 32145
rect 5062 32123 5071 32145
rect 5095 32123 5114 32145
rect 5114 32123 5128 32145
rect 5128 32123 5151 32145
rect 5175 32123 5180 32145
rect 5180 32123 5194 32145
rect 5194 32123 5231 32145
rect 5255 32123 5260 32145
rect 5260 32123 5311 32145
rect 4935 32093 4982 32098
rect 4982 32093 4991 32098
rect 5015 32093 5048 32098
rect 5048 32093 5062 32098
rect 5062 32093 5071 32098
rect 5095 32093 5114 32098
rect 5114 32093 5128 32098
rect 5128 32093 5151 32098
rect 5175 32093 5180 32098
rect 5180 32093 5194 32098
rect 5194 32093 5231 32098
rect 5255 32093 5260 32098
rect 5260 32093 5311 32098
rect 5335 32123 5378 32145
rect 5378 32123 5391 32145
rect 5415 32123 5444 32145
rect 5444 32123 5471 32145
rect 5495 32123 5551 32179
rect 5335 32093 5378 32098
rect 5378 32093 5391 32098
rect 5415 32093 5444 32098
rect 5444 32093 5471 32098
rect 4775 32080 4831 32093
rect 4855 32080 4911 32093
rect 4935 32080 4991 32093
rect 5015 32080 5071 32093
rect 5095 32080 5151 32093
rect 5175 32080 5231 32093
rect 5255 32080 5311 32093
rect 5335 32080 5391 32093
rect 5415 32080 5471 32093
rect 4775 32042 4784 32080
rect 4784 32042 4798 32080
rect 4798 32042 4831 32080
rect 4855 32042 4864 32080
rect 4864 32042 4911 32080
rect 4935 32042 4982 32080
rect 4982 32042 4991 32080
rect 5015 32042 5048 32080
rect 5048 32042 5062 32080
rect 5062 32042 5071 32080
rect 5095 32042 5114 32080
rect 5114 32042 5128 32080
rect 5128 32042 5151 32080
rect 5175 32042 5180 32080
rect 5180 32042 5194 32080
rect 5194 32042 5231 32080
rect 5255 32042 5260 32080
rect 5260 32042 5311 32080
rect 5335 32042 5378 32080
rect 5378 32042 5391 32080
rect 5415 32042 5444 32080
rect 5444 32042 5471 32080
rect 5495 32042 5551 32098
rect 4775 32015 4831 32017
rect 4855 32015 4911 32017
rect 4935 32015 4991 32017
rect 5015 32015 5071 32017
rect 5095 32015 5151 32017
rect 5175 32015 5231 32017
rect 5255 32015 5311 32017
rect 5335 32015 5391 32017
rect 5415 32015 5471 32017
rect 4775 31963 4784 32015
rect 4784 31963 4798 32015
rect 4798 31963 4831 32015
rect 4855 31963 4864 32015
rect 4864 31963 4911 32015
rect 4935 31963 4982 32015
rect 4982 31963 4991 32015
rect 5015 31963 5048 32015
rect 5048 31963 5062 32015
rect 5062 31963 5071 32015
rect 5095 31963 5114 32015
rect 5114 31963 5128 32015
rect 5128 31963 5151 32015
rect 5175 31963 5180 32015
rect 5180 31963 5194 32015
rect 5194 31963 5231 32015
rect 5255 31963 5260 32015
rect 5260 31963 5311 32015
rect 5335 31963 5378 32015
rect 5378 31963 5391 32015
rect 5415 31963 5444 32015
rect 5444 31963 5471 32015
rect 4775 31961 4831 31963
rect 4855 31961 4911 31963
rect 4935 31961 4991 31963
rect 5015 31961 5071 31963
rect 5095 31961 5151 31963
rect 5175 31961 5231 31963
rect 5255 31961 5311 31963
rect 5335 31961 5391 31963
rect 5415 31961 5471 31963
rect 5495 31961 5551 32017
rect 4775 31898 4784 31936
rect 4784 31898 4798 31936
rect 4798 31898 4831 31936
rect 4855 31898 4864 31936
rect 4864 31898 4911 31936
rect 4935 31898 4982 31936
rect 4982 31898 4991 31936
rect 5015 31898 5048 31936
rect 5048 31898 5062 31936
rect 5062 31898 5071 31936
rect 5095 31898 5114 31936
rect 5114 31898 5128 31936
rect 5128 31898 5151 31936
rect 5175 31898 5180 31936
rect 5180 31898 5194 31936
rect 5194 31898 5231 31936
rect 5255 31898 5260 31936
rect 5260 31898 5311 31936
rect 5335 31898 5378 31936
rect 5378 31898 5391 31936
rect 5415 31898 5444 31936
rect 5444 31898 5471 31936
rect 4775 31885 4831 31898
rect 4855 31885 4911 31898
rect 4935 31885 4991 31898
rect 5015 31885 5071 31898
rect 5095 31885 5151 31898
rect 5175 31885 5231 31898
rect 5255 31885 5311 31898
rect 5335 31885 5391 31898
rect 5415 31885 5471 31898
rect 4775 31880 4784 31885
rect 4784 31880 4798 31885
rect 4798 31880 4831 31885
rect 4855 31880 4864 31885
rect 4864 31880 4911 31885
rect 4775 31833 4784 31855
rect 4784 31833 4798 31855
rect 4798 31833 4831 31855
rect 4855 31833 4864 31855
rect 4864 31833 4911 31855
rect 4935 31880 4982 31885
rect 4982 31880 4991 31885
rect 5015 31880 5048 31885
rect 5048 31880 5062 31885
rect 5062 31880 5071 31885
rect 5095 31880 5114 31885
rect 5114 31880 5128 31885
rect 5128 31880 5151 31885
rect 5175 31880 5180 31885
rect 5180 31880 5194 31885
rect 5194 31880 5231 31885
rect 5255 31880 5260 31885
rect 5260 31880 5311 31885
rect 4935 31833 4982 31855
rect 4982 31833 4991 31855
rect 5015 31833 5048 31855
rect 5048 31833 5062 31855
rect 5062 31833 5071 31855
rect 5095 31833 5114 31855
rect 5114 31833 5128 31855
rect 5128 31833 5151 31855
rect 5175 31833 5180 31855
rect 5180 31833 5194 31855
rect 5194 31833 5231 31855
rect 5255 31833 5260 31855
rect 5260 31833 5311 31855
rect 5335 31880 5378 31885
rect 5378 31880 5391 31885
rect 5415 31880 5444 31885
rect 5444 31880 5471 31885
rect 5495 31880 5551 31936
rect 5335 31833 5378 31855
rect 5378 31833 5391 31855
rect 5415 31833 5444 31855
rect 5444 31833 5471 31855
rect 4775 31820 4831 31833
rect 4855 31820 4911 31833
rect 4935 31820 4991 31833
rect 5015 31820 5071 31833
rect 5095 31820 5151 31833
rect 5175 31820 5231 31833
rect 5255 31820 5311 31833
rect 5335 31820 5391 31833
rect 5415 31820 5471 31833
rect 4775 31799 4784 31820
rect 4784 31799 4798 31820
rect 4798 31799 4831 31820
rect 4855 31799 4864 31820
rect 4864 31799 4911 31820
rect 4775 31768 4784 31774
rect 4784 31768 4798 31774
rect 4798 31768 4831 31774
rect 4855 31768 4864 31774
rect 4864 31768 4911 31774
rect 4935 31799 4982 31820
rect 4982 31799 4991 31820
rect 5015 31799 5048 31820
rect 5048 31799 5062 31820
rect 5062 31799 5071 31820
rect 5095 31799 5114 31820
rect 5114 31799 5128 31820
rect 5128 31799 5151 31820
rect 5175 31799 5180 31820
rect 5180 31799 5194 31820
rect 5194 31799 5231 31820
rect 5255 31799 5260 31820
rect 5260 31799 5311 31820
rect 4935 31768 4982 31774
rect 4982 31768 4991 31774
rect 5015 31768 5048 31774
rect 5048 31768 5062 31774
rect 5062 31768 5071 31774
rect 5095 31768 5114 31774
rect 5114 31768 5128 31774
rect 5128 31768 5151 31774
rect 5175 31768 5180 31774
rect 5180 31768 5194 31774
rect 5194 31768 5231 31774
rect 5255 31768 5260 31774
rect 5260 31768 5311 31774
rect 5335 31799 5378 31820
rect 5378 31799 5391 31820
rect 5415 31799 5444 31820
rect 5444 31799 5471 31820
rect 5495 31799 5551 31855
rect 5335 31768 5378 31774
rect 5378 31768 5391 31774
rect 5415 31768 5444 31774
rect 5444 31768 5471 31774
rect 4775 31755 4831 31768
rect 4855 31755 4911 31768
rect 4935 31755 4991 31768
rect 5015 31755 5071 31768
rect 5095 31755 5151 31768
rect 5175 31755 5231 31768
rect 5255 31755 5311 31768
rect 5335 31755 5391 31768
rect 5415 31755 5471 31768
rect 4775 31718 4784 31755
rect 4784 31718 4798 31755
rect 4798 31718 4831 31755
rect 4855 31718 4864 31755
rect 4864 31718 4911 31755
rect 4935 31718 4982 31755
rect 4982 31718 4991 31755
rect 5015 31718 5048 31755
rect 5048 31718 5062 31755
rect 5062 31718 5071 31755
rect 5095 31718 5114 31755
rect 5114 31718 5128 31755
rect 5128 31718 5151 31755
rect 5175 31718 5180 31755
rect 5180 31718 5194 31755
rect 5194 31718 5231 31755
rect 5255 31718 5260 31755
rect 5260 31718 5311 31755
rect 5335 31718 5378 31755
rect 5378 31718 5391 31755
rect 5415 31718 5444 31755
rect 5444 31718 5471 31755
rect 5495 31718 5551 31774
rect 4775 31690 4831 31693
rect 4855 31690 4911 31693
rect 4935 31690 4991 31693
rect 5015 31690 5071 31693
rect 5095 31690 5151 31693
rect 5175 31690 5231 31693
rect 5255 31690 5311 31693
rect 5335 31690 5391 31693
rect 5415 31690 5471 31693
rect 4775 31638 4784 31690
rect 4784 31638 4798 31690
rect 4798 31638 4831 31690
rect 4855 31638 4864 31690
rect 4864 31638 4911 31690
rect 4935 31638 4982 31690
rect 4982 31638 4991 31690
rect 5015 31638 5048 31690
rect 5048 31638 5062 31690
rect 5062 31638 5071 31690
rect 5095 31638 5114 31690
rect 5114 31638 5128 31690
rect 5128 31638 5151 31690
rect 5175 31638 5180 31690
rect 5180 31638 5194 31690
rect 5194 31638 5231 31690
rect 5255 31638 5260 31690
rect 5260 31638 5311 31690
rect 5335 31638 5378 31690
rect 5378 31638 5391 31690
rect 5415 31638 5444 31690
rect 5444 31638 5471 31690
rect 4775 31637 4831 31638
rect 4855 31637 4911 31638
rect 4935 31637 4991 31638
rect 5015 31637 5071 31638
rect 5095 31637 5151 31638
rect 5175 31637 5231 31638
rect 5255 31637 5311 31638
rect 5335 31637 5391 31638
rect 5415 31637 5471 31638
rect 5495 31637 5551 31693
rect 4775 31573 4784 31612
rect 4784 31573 4798 31612
rect 4798 31573 4831 31612
rect 4855 31573 4864 31612
rect 4864 31573 4911 31612
rect 4935 31573 4982 31612
rect 4982 31573 4991 31612
rect 5015 31573 5048 31612
rect 5048 31573 5062 31612
rect 5062 31573 5071 31612
rect 5095 31573 5114 31612
rect 5114 31573 5128 31612
rect 5128 31573 5151 31612
rect 5175 31573 5180 31612
rect 5180 31573 5194 31612
rect 5194 31573 5231 31612
rect 5255 31573 5260 31612
rect 5260 31573 5311 31612
rect 5335 31573 5378 31612
rect 5378 31573 5391 31612
rect 5415 31573 5444 31612
rect 5444 31573 5471 31612
rect 4775 31560 4831 31573
rect 4855 31560 4911 31573
rect 4935 31560 4991 31573
rect 5015 31560 5071 31573
rect 5095 31560 5151 31573
rect 5175 31560 5231 31573
rect 5255 31560 5311 31573
rect 5335 31560 5391 31573
rect 5415 31560 5471 31573
rect 4775 31556 4784 31560
rect 4784 31556 4798 31560
rect 4798 31556 4831 31560
rect 4855 31556 4864 31560
rect 4864 31556 4911 31560
rect 4775 31508 4784 31531
rect 4784 31508 4798 31531
rect 4798 31508 4831 31531
rect 4855 31508 4864 31531
rect 4864 31508 4911 31531
rect 4935 31556 4982 31560
rect 4982 31556 4991 31560
rect 5015 31556 5048 31560
rect 5048 31556 5062 31560
rect 5062 31556 5071 31560
rect 5095 31556 5114 31560
rect 5114 31556 5128 31560
rect 5128 31556 5151 31560
rect 5175 31556 5180 31560
rect 5180 31556 5194 31560
rect 5194 31556 5231 31560
rect 5255 31556 5260 31560
rect 5260 31556 5311 31560
rect 4935 31508 4982 31531
rect 4982 31508 4991 31531
rect 5015 31508 5048 31531
rect 5048 31508 5062 31531
rect 5062 31508 5071 31531
rect 5095 31508 5114 31531
rect 5114 31508 5128 31531
rect 5128 31508 5151 31531
rect 5175 31508 5180 31531
rect 5180 31508 5194 31531
rect 5194 31508 5231 31531
rect 5255 31508 5260 31531
rect 5260 31508 5311 31531
rect 5335 31556 5378 31560
rect 5378 31556 5391 31560
rect 5415 31556 5444 31560
rect 5444 31556 5471 31560
rect 5495 31556 5551 31612
rect 5335 31508 5378 31531
rect 5378 31508 5391 31531
rect 5415 31508 5444 31531
rect 5444 31508 5471 31531
rect 4775 31495 4831 31508
rect 4855 31495 4911 31508
rect 4935 31495 4991 31508
rect 5015 31495 5071 31508
rect 5095 31495 5151 31508
rect 5175 31495 5231 31508
rect 5255 31495 5311 31508
rect 5335 31495 5391 31508
rect 5415 31495 5471 31508
rect 4775 31475 4784 31495
rect 4784 31475 4798 31495
rect 4798 31475 4831 31495
rect 4855 31475 4864 31495
rect 4864 31475 4911 31495
rect 4775 31443 4784 31450
rect 4784 31443 4798 31450
rect 4798 31443 4831 31450
rect 4855 31443 4864 31450
rect 4864 31443 4911 31450
rect 4935 31475 4982 31495
rect 4982 31475 4991 31495
rect 5015 31475 5048 31495
rect 5048 31475 5062 31495
rect 5062 31475 5071 31495
rect 5095 31475 5114 31495
rect 5114 31475 5128 31495
rect 5128 31475 5151 31495
rect 5175 31475 5180 31495
rect 5180 31475 5194 31495
rect 5194 31475 5231 31495
rect 5255 31475 5260 31495
rect 5260 31475 5311 31495
rect 4935 31443 4982 31450
rect 4982 31443 4991 31450
rect 5015 31443 5048 31450
rect 5048 31443 5062 31450
rect 5062 31443 5071 31450
rect 5095 31443 5114 31450
rect 5114 31443 5128 31450
rect 5128 31443 5151 31450
rect 5175 31443 5180 31450
rect 5180 31443 5194 31450
rect 5194 31443 5231 31450
rect 5255 31443 5260 31450
rect 5260 31443 5311 31450
rect 5335 31475 5378 31495
rect 5378 31475 5391 31495
rect 5415 31475 5444 31495
rect 5444 31475 5471 31495
rect 5495 31475 5551 31531
rect 5335 31443 5378 31450
rect 5378 31443 5391 31450
rect 5415 31443 5444 31450
rect 5444 31443 5471 31450
rect 4775 31430 4831 31443
rect 4855 31430 4911 31443
rect 4935 31430 4991 31443
rect 5015 31430 5071 31443
rect 5095 31430 5151 31443
rect 5175 31430 5231 31443
rect 5255 31430 5311 31443
rect 5335 31430 5391 31443
rect 5415 31430 5471 31443
rect 4775 31394 4784 31430
rect 4784 31394 4798 31430
rect 4798 31394 4831 31430
rect 4855 31394 4864 31430
rect 4864 31394 4911 31430
rect 4935 31394 4982 31430
rect 4982 31394 4991 31430
rect 5015 31394 5048 31430
rect 5048 31394 5062 31430
rect 5062 31394 5071 31430
rect 5095 31394 5114 31430
rect 5114 31394 5128 31430
rect 5128 31394 5151 31430
rect 5175 31394 5180 31430
rect 5180 31394 5194 31430
rect 5194 31394 5231 31430
rect 5255 31394 5260 31430
rect 5260 31394 5311 31430
rect 5335 31394 5378 31430
rect 5378 31394 5391 31430
rect 5415 31394 5444 31430
rect 5444 31394 5471 31430
rect 5495 31394 5551 31450
rect 4775 31365 4831 31369
rect 4855 31365 4911 31369
rect 4935 31365 4991 31369
rect 5015 31365 5071 31369
rect 5095 31365 5151 31369
rect 5175 31365 5231 31369
rect 5255 31365 5311 31369
rect 5335 31365 5391 31369
rect 5415 31365 5471 31369
rect 4775 31313 4784 31365
rect 4784 31313 4798 31365
rect 4798 31313 4831 31365
rect 4855 31313 4864 31365
rect 4864 31313 4911 31365
rect 4935 31313 4982 31365
rect 4982 31313 4991 31365
rect 5015 31313 5048 31365
rect 5048 31313 5062 31365
rect 5062 31313 5071 31365
rect 5095 31313 5114 31365
rect 5114 31313 5128 31365
rect 5128 31313 5151 31365
rect 5175 31313 5180 31365
rect 5180 31313 5194 31365
rect 5194 31313 5231 31365
rect 5255 31313 5260 31365
rect 5260 31313 5311 31365
rect 5335 31313 5378 31365
rect 5378 31313 5391 31365
rect 5415 31313 5444 31365
rect 5444 31313 5471 31365
rect 5495 31313 5551 31369
rect 4775 31248 4784 31288
rect 4784 31248 4798 31288
rect 4798 31248 4831 31288
rect 4855 31248 4864 31288
rect 4864 31248 4911 31288
rect 4935 31248 4982 31288
rect 4982 31248 4991 31288
rect 5015 31248 5048 31288
rect 5048 31248 5062 31288
rect 5062 31248 5071 31288
rect 5095 31248 5114 31288
rect 5114 31248 5128 31288
rect 5128 31248 5151 31288
rect 5175 31248 5180 31288
rect 5180 31248 5194 31288
rect 5194 31248 5231 31288
rect 5255 31248 5260 31288
rect 5260 31248 5311 31288
rect 5335 31248 5378 31288
rect 5378 31248 5391 31288
rect 5415 31248 5444 31288
rect 5444 31248 5471 31288
rect 4775 31235 4831 31248
rect 4855 31235 4911 31248
rect 4935 31235 4991 31248
rect 5015 31235 5071 31248
rect 5095 31235 5151 31248
rect 5175 31235 5231 31248
rect 5255 31235 5311 31248
rect 5335 31235 5391 31248
rect 5415 31235 5471 31248
rect 4775 31232 4784 31235
rect 4784 31232 4798 31235
rect 4798 31232 4831 31235
rect 4855 31232 4864 31235
rect 4864 31232 4911 31235
rect 4775 31183 4784 31207
rect 4784 31183 4798 31207
rect 4798 31183 4831 31207
rect 4855 31183 4864 31207
rect 4864 31183 4911 31207
rect 4935 31232 4982 31235
rect 4982 31232 4991 31235
rect 5015 31232 5048 31235
rect 5048 31232 5062 31235
rect 5062 31232 5071 31235
rect 5095 31232 5114 31235
rect 5114 31232 5128 31235
rect 5128 31232 5151 31235
rect 5175 31232 5180 31235
rect 5180 31232 5194 31235
rect 5194 31232 5231 31235
rect 5255 31232 5260 31235
rect 5260 31232 5311 31235
rect 4935 31183 4982 31207
rect 4982 31183 4991 31207
rect 5015 31183 5048 31207
rect 5048 31183 5062 31207
rect 5062 31183 5071 31207
rect 5095 31183 5114 31207
rect 5114 31183 5128 31207
rect 5128 31183 5151 31207
rect 5175 31183 5180 31207
rect 5180 31183 5194 31207
rect 5194 31183 5231 31207
rect 5255 31183 5260 31207
rect 5260 31183 5311 31207
rect 5335 31232 5378 31235
rect 5378 31232 5391 31235
rect 5415 31232 5444 31235
rect 5444 31232 5471 31235
rect 5495 31232 5551 31288
rect 5335 31183 5378 31207
rect 5378 31183 5391 31207
rect 5415 31183 5444 31207
rect 5444 31183 5471 31207
rect 4775 31170 4831 31183
rect 4855 31170 4911 31183
rect 4935 31170 4991 31183
rect 5015 31170 5071 31183
rect 5095 31170 5151 31183
rect 5175 31170 5231 31183
rect 5255 31170 5311 31183
rect 5335 31170 5391 31183
rect 5415 31170 5471 31183
rect 4775 31151 4784 31170
rect 4784 31151 4798 31170
rect 4798 31151 4831 31170
rect 4855 31151 4864 31170
rect 4864 31151 4911 31170
rect 4775 31118 4784 31126
rect 4784 31118 4798 31126
rect 4798 31118 4831 31126
rect 4855 31118 4864 31126
rect 4864 31118 4911 31126
rect 4935 31151 4982 31170
rect 4982 31151 4991 31170
rect 5015 31151 5048 31170
rect 5048 31151 5062 31170
rect 5062 31151 5071 31170
rect 5095 31151 5114 31170
rect 5114 31151 5128 31170
rect 5128 31151 5151 31170
rect 5175 31151 5180 31170
rect 5180 31151 5194 31170
rect 5194 31151 5231 31170
rect 5255 31151 5260 31170
rect 5260 31151 5311 31170
rect 4935 31118 4982 31126
rect 4982 31118 4991 31126
rect 5015 31118 5048 31126
rect 5048 31118 5062 31126
rect 5062 31118 5071 31126
rect 5095 31118 5114 31126
rect 5114 31118 5128 31126
rect 5128 31118 5151 31126
rect 5175 31118 5180 31126
rect 5180 31118 5194 31126
rect 5194 31118 5231 31126
rect 5255 31118 5260 31126
rect 5260 31118 5311 31126
rect 5335 31151 5378 31170
rect 5378 31151 5391 31170
rect 5415 31151 5444 31170
rect 5444 31151 5471 31170
rect 5495 31151 5551 31207
rect 5335 31118 5378 31126
rect 5378 31118 5391 31126
rect 5415 31118 5444 31126
rect 5444 31118 5471 31126
rect 4775 31105 4831 31118
rect 4855 31105 4911 31118
rect 4935 31105 4991 31118
rect 5015 31105 5071 31118
rect 5095 31105 5151 31118
rect 5175 31105 5231 31118
rect 5255 31105 5311 31118
rect 5335 31105 5391 31118
rect 5415 31105 5471 31118
rect 4775 31070 4784 31105
rect 4784 31070 4798 31105
rect 4798 31070 4831 31105
rect 4855 31070 4864 31105
rect 4864 31070 4911 31105
rect 4935 31070 4982 31105
rect 4982 31070 4991 31105
rect 5015 31070 5048 31105
rect 5048 31070 5062 31105
rect 5062 31070 5071 31105
rect 5095 31070 5114 31105
rect 5114 31070 5128 31105
rect 5128 31070 5151 31105
rect 5175 31070 5180 31105
rect 5180 31070 5194 31105
rect 5194 31070 5231 31105
rect 5255 31070 5260 31105
rect 5260 31070 5311 31105
rect 5335 31070 5378 31105
rect 5378 31070 5391 31105
rect 5415 31070 5444 31105
rect 5444 31070 5471 31105
rect 5495 31070 5551 31126
rect 4775 31040 4831 31045
rect 4855 31040 4911 31045
rect 4935 31040 4991 31045
rect 5015 31040 5071 31045
rect 5095 31040 5151 31045
rect 5175 31040 5231 31045
rect 5255 31040 5311 31045
rect 5335 31040 5391 31045
rect 5415 31040 5471 31045
rect 4775 30989 4784 31040
rect 4784 30989 4798 31040
rect 4798 30989 4831 31040
rect 4855 30989 4864 31040
rect 4864 30989 4911 31040
rect 4935 30989 4982 31040
rect 4982 30989 4991 31040
rect 5015 30989 5048 31040
rect 5048 30989 5062 31040
rect 5062 30989 5071 31040
rect 5095 30989 5114 31040
rect 5114 30989 5128 31040
rect 5128 30989 5151 31040
rect 5175 30989 5180 31040
rect 5180 30989 5194 31040
rect 5194 30989 5231 31040
rect 5255 30989 5260 31040
rect 5260 30989 5311 31040
rect 5335 30989 5378 31040
rect 5378 30989 5391 31040
rect 5415 30989 5444 31040
rect 5444 30989 5471 31040
rect 5495 30989 5551 31045
rect 4775 30923 4784 30964
rect 4784 30923 4798 30964
rect 4798 30923 4831 30964
rect 4855 30923 4864 30964
rect 4864 30923 4911 30964
rect 4935 30923 4982 30964
rect 4982 30923 4991 30964
rect 5015 30923 5048 30964
rect 5048 30923 5062 30964
rect 5062 30923 5071 30964
rect 5095 30923 5114 30964
rect 5114 30923 5128 30964
rect 5128 30923 5151 30964
rect 5175 30923 5180 30964
rect 5180 30923 5194 30964
rect 5194 30923 5231 30964
rect 5255 30923 5260 30964
rect 5260 30923 5311 30964
rect 5335 30923 5378 30964
rect 5378 30923 5391 30964
rect 5415 30923 5444 30964
rect 5444 30923 5471 30964
rect 4775 30910 4831 30923
rect 4855 30910 4911 30923
rect 4935 30910 4991 30923
rect 5015 30910 5071 30923
rect 5095 30910 5151 30923
rect 5175 30910 5231 30923
rect 5255 30910 5311 30923
rect 5335 30910 5391 30923
rect 5415 30910 5471 30923
rect 4775 30908 4784 30910
rect 4784 30908 4798 30910
rect 4798 30908 4831 30910
rect 4855 30908 4864 30910
rect 4864 30908 4911 30910
rect 4775 30858 4784 30883
rect 4784 30858 4798 30883
rect 4798 30858 4831 30883
rect 4855 30858 4864 30883
rect 4864 30858 4911 30883
rect 4935 30908 4982 30910
rect 4982 30908 4991 30910
rect 5015 30908 5048 30910
rect 5048 30908 5062 30910
rect 5062 30908 5071 30910
rect 5095 30908 5114 30910
rect 5114 30908 5128 30910
rect 5128 30908 5151 30910
rect 5175 30908 5180 30910
rect 5180 30908 5194 30910
rect 5194 30908 5231 30910
rect 5255 30908 5260 30910
rect 5260 30908 5311 30910
rect 4935 30858 4982 30883
rect 4982 30858 4991 30883
rect 5015 30858 5048 30883
rect 5048 30858 5062 30883
rect 5062 30858 5071 30883
rect 5095 30858 5114 30883
rect 5114 30858 5128 30883
rect 5128 30858 5151 30883
rect 5175 30858 5180 30883
rect 5180 30858 5194 30883
rect 5194 30858 5231 30883
rect 5255 30858 5260 30883
rect 5260 30858 5311 30883
rect 5335 30908 5378 30910
rect 5378 30908 5391 30910
rect 5415 30908 5444 30910
rect 5444 30908 5471 30910
rect 5495 30908 5551 30964
rect 5335 30858 5378 30883
rect 5378 30858 5391 30883
rect 5415 30858 5444 30883
rect 5444 30858 5471 30883
rect 4775 30845 4831 30858
rect 4855 30845 4911 30858
rect 4935 30845 4991 30858
rect 5015 30845 5071 30858
rect 5095 30845 5151 30858
rect 5175 30845 5231 30858
rect 5255 30845 5311 30858
rect 5335 30845 5391 30858
rect 5415 30845 5471 30858
rect 4775 30827 4784 30845
rect 4784 30827 4798 30845
rect 4798 30827 4831 30845
rect 4855 30827 4864 30845
rect 4864 30827 4911 30845
rect 4775 30793 4784 30802
rect 4784 30793 4798 30802
rect 4798 30793 4831 30802
rect 4855 30793 4864 30802
rect 4864 30793 4911 30802
rect 4935 30827 4982 30845
rect 4982 30827 4991 30845
rect 5015 30827 5048 30845
rect 5048 30827 5062 30845
rect 5062 30827 5071 30845
rect 5095 30827 5114 30845
rect 5114 30827 5128 30845
rect 5128 30827 5151 30845
rect 5175 30827 5180 30845
rect 5180 30827 5194 30845
rect 5194 30827 5231 30845
rect 5255 30827 5260 30845
rect 5260 30827 5311 30845
rect 4935 30793 4982 30802
rect 4982 30793 4991 30802
rect 5015 30793 5048 30802
rect 5048 30793 5062 30802
rect 5062 30793 5071 30802
rect 5095 30793 5114 30802
rect 5114 30793 5128 30802
rect 5128 30793 5151 30802
rect 5175 30793 5180 30802
rect 5180 30793 5194 30802
rect 5194 30793 5231 30802
rect 5255 30793 5260 30802
rect 5260 30793 5311 30802
rect 5335 30827 5378 30845
rect 5378 30827 5391 30845
rect 5415 30827 5444 30845
rect 5444 30827 5471 30845
rect 5495 30827 5551 30883
rect 5335 30793 5378 30802
rect 5378 30793 5391 30802
rect 5415 30793 5444 30802
rect 5444 30793 5471 30802
rect 4775 30780 4831 30793
rect 4855 30780 4911 30793
rect 4935 30780 4991 30793
rect 5015 30780 5071 30793
rect 5095 30780 5151 30793
rect 5175 30780 5231 30793
rect 5255 30780 5311 30793
rect 5335 30780 5391 30793
rect 5415 30780 5471 30793
rect 4775 30746 4784 30780
rect 4784 30746 4798 30780
rect 4798 30746 4831 30780
rect 4855 30746 4864 30780
rect 4864 30746 4911 30780
rect 4935 30746 4982 30780
rect 4982 30746 4991 30780
rect 5015 30746 5048 30780
rect 5048 30746 5062 30780
rect 5062 30746 5071 30780
rect 5095 30746 5114 30780
rect 5114 30746 5128 30780
rect 5128 30746 5151 30780
rect 5175 30746 5180 30780
rect 5180 30746 5194 30780
rect 5194 30746 5231 30780
rect 5255 30746 5260 30780
rect 5260 30746 5311 30780
rect 5335 30746 5378 30780
rect 5378 30746 5391 30780
rect 5415 30746 5444 30780
rect 5444 30746 5471 30780
rect 5495 30746 5551 30802
rect 4775 30715 4831 30721
rect 4855 30715 4911 30721
rect 4935 30715 4991 30721
rect 5015 30715 5071 30721
rect 5095 30715 5151 30721
rect 5175 30715 5231 30721
rect 5255 30715 5311 30721
rect 5335 30715 5391 30721
rect 5415 30715 5471 30721
rect 4775 30665 4784 30715
rect 4784 30665 4798 30715
rect 4798 30665 4831 30715
rect 4855 30665 4864 30715
rect 4864 30665 4911 30715
rect 4935 30665 4982 30715
rect 4982 30665 4991 30715
rect 5015 30665 5048 30715
rect 5048 30665 5062 30715
rect 5062 30665 5071 30715
rect 5095 30665 5114 30715
rect 5114 30665 5128 30715
rect 5128 30665 5151 30715
rect 5175 30665 5180 30715
rect 5180 30665 5194 30715
rect 5194 30665 5231 30715
rect 5255 30665 5260 30715
rect 5260 30665 5311 30715
rect 5335 30665 5378 30715
rect 5378 30665 5391 30715
rect 5415 30665 5444 30715
rect 5444 30665 5471 30715
rect 5495 30665 5551 30721
rect 4775 30598 4784 30640
rect 4784 30598 4798 30640
rect 4798 30598 4831 30640
rect 4855 30598 4864 30640
rect 4864 30598 4911 30640
rect 4935 30598 4982 30640
rect 4982 30598 4991 30640
rect 5015 30598 5048 30640
rect 5048 30598 5062 30640
rect 5062 30598 5071 30640
rect 5095 30598 5114 30640
rect 5114 30598 5128 30640
rect 5128 30598 5151 30640
rect 5175 30598 5180 30640
rect 5180 30598 5194 30640
rect 5194 30598 5231 30640
rect 5255 30598 5260 30640
rect 5260 30598 5311 30640
rect 5335 30598 5378 30640
rect 5378 30598 5391 30640
rect 5415 30598 5444 30640
rect 5444 30598 5471 30640
rect 4775 30585 4831 30598
rect 4855 30585 4911 30598
rect 4935 30585 4991 30598
rect 5015 30585 5071 30598
rect 5095 30585 5151 30598
rect 5175 30585 5231 30598
rect 5255 30585 5311 30598
rect 5335 30585 5391 30598
rect 5415 30585 5471 30598
rect 4775 30584 4784 30585
rect 4784 30584 4798 30585
rect 4798 30584 4831 30585
rect 4855 30584 4864 30585
rect 4864 30584 4911 30585
rect 4775 30533 4784 30559
rect 4784 30533 4798 30559
rect 4798 30533 4831 30559
rect 4855 30533 4864 30559
rect 4864 30533 4911 30559
rect 4935 30584 4982 30585
rect 4982 30584 4991 30585
rect 5015 30584 5048 30585
rect 5048 30584 5062 30585
rect 5062 30584 5071 30585
rect 5095 30584 5114 30585
rect 5114 30584 5128 30585
rect 5128 30584 5151 30585
rect 5175 30584 5180 30585
rect 5180 30584 5194 30585
rect 5194 30584 5231 30585
rect 5255 30584 5260 30585
rect 5260 30584 5311 30585
rect 4935 30533 4982 30559
rect 4982 30533 4991 30559
rect 5015 30533 5048 30559
rect 5048 30533 5062 30559
rect 5062 30533 5071 30559
rect 5095 30533 5114 30559
rect 5114 30533 5128 30559
rect 5128 30533 5151 30559
rect 5175 30533 5180 30559
rect 5180 30533 5194 30559
rect 5194 30533 5231 30559
rect 5255 30533 5260 30559
rect 5260 30533 5311 30559
rect 5335 30584 5378 30585
rect 5378 30584 5391 30585
rect 5415 30584 5444 30585
rect 5444 30584 5471 30585
rect 5495 30584 5551 30640
rect 5335 30533 5378 30559
rect 5378 30533 5391 30559
rect 5415 30533 5444 30559
rect 5444 30533 5471 30559
rect 4775 30520 4831 30533
rect 4855 30520 4911 30533
rect 4935 30520 4991 30533
rect 5015 30520 5071 30533
rect 5095 30520 5151 30533
rect 5175 30520 5231 30533
rect 5255 30520 5311 30533
rect 5335 30520 5391 30533
rect 5415 30520 5471 30533
rect 4775 30503 4784 30520
rect 4784 30503 4798 30520
rect 4798 30503 4831 30520
rect 4855 30503 4864 30520
rect 4864 30503 4911 30520
rect 4775 30468 4784 30478
rect 4784 30468 4798 30478
rect 4798 30468 4831 30478
rect 4855 30468 4864 30478
rect 4864 30468 4911 30478
rect 4935 30503 4982 30520
rect 4982 30503 4991 30520
rect 5015 30503 5048 30520
rect 5048 30503 5062 30520
rect 5062 30503 5071 30520
rect 5095 30503 5114 30520
rect 5114 30503 5128 30520
rect 5128 30503 5151 30520
rect 5175 30503 5180 30520
rect 5180 30503 5194 30520
rect 5194 30503 5231 30520
rect 5255 30503 5260 30520
rect 5260 30503 5311 30520
rect 4935 30468 4982 30478
rect 4982 30468 4991 30478
rect 5015 30468 5048 30478
rect 5048 30468 5062 30478
rect 5062 30468 5071 30478
rect 5095 30468 5114 30478
rect 5114 30468 5128 30478
rect 5128 30468 5151 30478
rect 5175 30468 5180 30478
rect 5180 30468 5194 30478
rect 5194 30468 5231 30478
rect 5255 30468 5260 30478
rect 5260 30468 5311 30478
rect 5335 30503 5378 30520
rect 5378 30503 5391 30520
rect 5415 30503 5444 30520
rect 5444 30503 5471 30520
rect 5495 30503 5551 30559
rect 5335 30468 5378 30478
rect 5378 30468 5391 30478
rect 5415 30468 5444 30478
rect 5444 30468 5471 30478
rect 4775 30455 4831 30468
rect 4855 30455 4911 30468
rect 4935 30455 4991 30468
rect 5015 30455 5071 30468
rect 5095 30455 5151 30468
rect 5175 30455 5231 30468
rect 5255 30455 5311 30468
rect 5335 30455 5391 30468
rect 5415 30455 5471 30468
rect 4775 30422 4784 30455
rect 4784 30422 4798 30455
rect 4798 30422 4831 30455
rect 4855 30422 4864 30455
rect 4864 30422 4911 30455
rect 4935 30422 4982 30455
rect 4982 30422 4991 30455
rect 5015 30422 5048 30455
rect 5048 30422 5062 30455
rect 5062 30422 5071 30455
rect 5095 30422 5114 30455
rect 5114 30422 5128 30455
rect 5128 30422 5151 30455
rect 5175 30422 5180 30455
rect 5180 30422 5194 30455
rect 5194 30422 5231 30455
rect 5255 30422 5260 30455
rect 5260 30422 5311 30455
rect 5335 30422 5378 30455
rect 5378 30422 5391 30455
rect 5415 30422 5444 30455
rect 5444 30422 5471 30455
rect 5495 30422 5551 30478
rect 4775 30390 4831 30397
rect 4855 30390 4911 30397
rect 4935 30390 4991 30397
rect 5015 30390 5071 30397
rect 5095 30390 5151 30397
rect 5175 30390 5231 30397
rect 5255 30390 5311 30397
rect 5335 30390 5391 30397
rect 5415 30390 5471 30397
rect 4775 30341 4784 30390
rect 4784 30341 4798 30390
rect 4798 30341 4831 30390
rect 4855 30341 4864 30390
rect 4864 30341 4911 30390
rect 4935 30341 4982 30390
rect 4982 30341 4991 30390
rect 5015 30341 5048 30390
rect 5048 30341 5062 30390
rect 5062 30341 5071 30390
rect 5095 30341 5114 30390
rect 5114 30341 5128 30390
rect 5128 30341 5151 30390
rect 5175 30341 5180 30390
rect 5180 30341 5194 30390
rect 5194 30341 5231 30390
rect 5255 30341 5260 30390
rect 5260 30341 5311 30390
rect 5335 30341 5378 30390
rect 5378 30341 5391 30390
rect 5415 30341 5444 30390
rect 5444 30341 5471 30390
rect 5495 30341 5551 30397
rect 4672 29819 4728 29875
rect 4757 29819 4813 29875
rect 4842 29819 4898 29875
rect 4926 29819 4982 29875
rect 5010 29819 5066 29875
rect 5094 29819 5150 29875
rect 5178 29819 5234 29875
rect 5262 29853 5313 29875
rect 5313 29853 5318 29875
rect 5262 29841 5318 29853
rect 5262 29819 5313 29841
rect 5313 29819 5318 29841
rect 5346 29819 5402 29875
rect 5430 29819 5486 29875
rect 5514 29819 5570 29875
rect 5598 29819 5654 29875
rect 4672 28835 4728 28891
rect 4757 28835 4813 28891
rect 4842 28835 4898 28891
rect 4926 28835 4982 28891
rect 5010 28835 5066 28891
rect 5094 28835 5150 28891
rect 5178 28835 5234 28891
rect 5262 28869 5313 28891
rect 5313 28869 5318 28891
rect 5262 28857 5318 28869
rect 5262 28835 5313 28857
rect 5313 28835 5318 28857
rect 5346 28835 5402 28891
rect 5430 28835 5486 28891
rect 5514 28835 5570 28891
rect 5598 28835 5654 28891
rect 4672 28443 4728 28445
rect 4757 28443 4813 28445
rect 4842 28443 4898 28445
rect 4926 28443 4982 28445
rect 5010 28443 5066 28445
rect 5094 28443 5150 28445
rect 5178 28443 5234 28445
rect 5262 28443 5318 28445
rect 5346 28443 5402 28445
rect 5430 28443 5486 28445
rect 5514 28443 5570 28445
rect 5598 28443 5654 28445
rect 4672 28391 4721 28443
rect 4721 28391 4728 28443
rect 4757 28391 4788 28443
rect 4788 28391 4803 28443
rect 4803 28391 4813 28443
rect 4842 28391 4855 28443
rect 4855 28391 4870 28443
rect 4870 28391 4898 28443
rect 4926 28391 4937 28443
rect 4937 28391 4982 28443
rect 5010 28391 5056 28443
rect 5056 28391 5066 28443
rect 5094 28391 5123 28443
rect 5123 28391 5138 28443
rect 5138 28391 5150 28443
rect 5178 28391 5190 28443
rect 5190 28391 5205 28443
rect 5205 28391 5234 28443
rect 5262 28391 5272 28443
rect 5272 28391 5318 28443
rect 5346 28391 5391 28443
rect 5391 28391 5402 28443
rect 5430 28391 5458 28443
rect 5458 28391 5473 28443
rect 5473 28391 5486 28443
rect 5514 28391 5525 28443
rect 5525 28391 5539 28443
rect 5539 28391 5570 28443
rect 5598 28391 5605 28443
rect 5605 28391 5654 28443
rect 4672 28389 4728 28391
rect 4757 28389 4813 28391
rect 4842 28389 4898 28391
rect 4926 28389 4982 28391
rect 5010 28389 5066 28391
rect 5094 28389 5150 28391
rect 5178 28389 5234 28391
rect 5262 28389 5318 28391
rect 5346 28389 5402 28391
rect 5430 28389 5486 28391
rect 5514 28389 5570 28391
rect 5598 28389 5654 28391
rect 3712 28183 3768 28185
rect 3793 28183 3849 28185
rect 3874 28183 3930 28185
rect 3955 28183 4011 28185
rect 4036 28183 4092 28185
rect 4117 28183 4173 28185
rect 4198 28183 4254 28185
rect 4278 28183 4334 28185
rect 4358 28183 4414 28185
rect 4438 28183 4494 28185
rect 3712 28131 3761 28183
rect 3761 28131 3768 28183
rect 3793 28131 3828 28183
rect 3828 28131 3843 28183
rect 3843 28131 3849 28183
rect 3874 28131 3895 28183
rect 3895 28131 3910 28183
rect 3910 28131 3930 28183
rect 3955 28131 3962 28183
rect 3962 28131 3977 28183
rect 3977 28131 4011 28183
rect 4036 28131 4044 28183
rect 4044 28131 4092 28183
rect 4117 28131 4163 28183
rect 4163 28131 4173 28183
rect 4198 28131 4230 28183
rect 4230 28131 4245 28183
rect 4245 28131 4254 28183
rect 4278 28131 4297 28183
rect 4297 28131 4312 28183
rect 4312 28131 4334 28183
rect 4358 28131 4364 28183
rect 4364 28131 4379 28183
rect 4379 28131 4414 28183
rect 4438 28131 4445 28183
rect 4445 28131 4494 28183
rect 3712 28129 3768 28131
rect 3793 28129 3849 28131
rect 3874 28129 3930 28131
rect 3955 28129 4011 28131
rect 4036 28129 4092 28131
rect 4117 28129 4173 28131
rect 4198 28129 4254 28131
rect 4278 28129 4334 28131
rect 4358 28129 4414 28131
rect 4438 28129 4494 28131
rect 1592 25393 1648 25449
rect 1673 25393 1729 25449
rect 1754 25393 1810 25449
rect 1835 25393 1891 25449
rect 1916 25393 1972 25449
rect 1997 25393 2053 25449
rect 1592 25313 1648 25369
rect 1673 25313 1729 25369
rect 1754 25313 1810 25369
rect 1835 25313 1891 25369
rect 1916 25313 1972 25369
rect 1997 25313 2053 25369
rect 1592 25233 1648 25289
rect 1673 25233 1729 25289
rect 1754 25233 1810 25289
rect 1835 25233 1891 25289
rect 1916 25233 1972 25289
rect 1997 25233 2053 25289
rect 1592 25153 1648 25209
rect 1673 25153 1729 25209
rect 1754 25153 1810 25209
rect 1835 25153 1891 25209
rect 1916 25153 1972 25209
rect 1997 25153 2053 25209
rect 2078 25153 2374 25449
rect 3712 23758 3768 23814
rect 3793 23758 3849 23814
rect 3874 23758 3930 23814
rect 3955 23758 4011 23814
rect 4036 23758 4092 23814
rect 4117 23758 4173 23814
rect 4198 23758 4254 23814
rect 4278 23758 4334 23814
rect 4358 23758 4414 23814
rect 4438 23792 4451 23814
rect 4451 23792 4494 23814
rect 4438 23780 4494 23792
rect 4438 23758 4451 23780
rect 4451 23758 4494 23780
rect 3712 20363 3768 20419
rect 3793 20363 3849 20419
rect 3874 20363 3930 20419
rect 3955 20363 4011 20419
rect 4036 20363 4092 20419
rect 4117 20363 4173 20419
rect 4198 20363 4254 20419
rect 4278 20363 4334 20419
rect 4358 20363 4414 20419
rect 4438 20363 4494 20419
rect 3712 19968 3768 20024
rect 3793 19968 3849 20024
rect 3874 19968 3930 20024
rect 3955 19968 4011 20024
rect 4036 19968 4092 20024
rect 4117 19968 4173 20024
rect 4198 19968 4254 20024
rect 4278 19968 4334 20024
rect 4358 19968 4414 20024
rect 4438 19968 4472 20024
rect 4472 19968 4494 20024
rect 3712 18298 3768 18300
rect 3793 18298 3849 18300
rect 3874 18298 3930 18300
rect 3955 18298 4011 18300
rect 4036 18298 4092 18300
rect 4117 18298 4173 18300
rect 4198 18298 4254 18300
rect 4278 18298 4334 18300
rect 4358 18298 4414 18300
rect 4438 18298 4494 18300
rect 3712 18246 3761 18298
rect 3761 18246 3768 18298
rect 3793 18246 3828 18298
rect 3828 18246 3843 18298
rect 3843 18246 3849 18298
rect 3874 18246 3895 18298
rect 3895 18246 3910 18298
rect 3910 18246 3930 18298
rect 3955 18246 3962 18298
rect 3962 18246 3977 18298
rect 3977 18246 4011 18298
rect 4036 18246 4044 18298
rect 4044 18246 4092 18298
rect 4117 18246 4163 18298
rect 4163 18246 4173 18298
rect 4198 18246 4230 18298
rect 4230 18246 4245 18298
rect 4245 18246 4254 18298
rect 4278 18246 4297 18298
rect 4297 18246 4312 18298
rect 4312 18246 4334 18298
rect 4358 18246 4364 18298
rect 4364 18246 4379 18298
rect 4379 18246 4414 18298
rect 4438 18246 4445 18298
rect 4445 18246 4494 18298
rect 3712 18244 3768 18246
rect 3793 18244 3849 18246
rect 3874 18244 3930 18246
rect 3955 18244 4011 18246
rect 4036 18244 4092 18246
rect 4117 18244 4173 18246
rect 4198 18244 4254 18246
rect 4278 18244 4334 18246
rect 4358 18244 4414 18246
rect 4438 18244 4494 18246
rect 4672 17839 4728 17895
rect 4757 17839 4813 17895
rect 4842 17873 4891 17895
rect 4891 17873 4898 17895
rect 4842 17861 4898 17873
rect 4842 17839 4891 17861
rect 4891 17839 4898 17861
rect 4926 17839 4982 17895
rect 5010 17839 5066 17895
rect 5094 17839 5150 17895
rect 5178 17873 5203 17895
rect 5203 17873 5234 17895
rect 5178 17861 5234 17873
rect 5178 17839 5203 17861
rect 5203 17839 5234 17861
rect 5262 17839 5318 17895
rect 5346 17839 5402 17895
rect 5430 17873 5462 17895
rect 5462 17873 5486 17895
rect 5430 17861 5486 17873
rect 5430 17839 5462 17861
rect 5462 17839 5486 17861
rect 5514 17839 5570 17895
rect 5598 17839 5654 17895
rect 4672 14811 4728 14867
rect 4757 14811 4813 14867
rect 4842 14811 4898 14867
rect 4926 14811 4982 14867
rect 5010 14811 5066 14867
rect 5094 14811 5150 14867
rect 5178 14811 5234 14867
rect 5262 14811 5318 14867
rect 5346 14811 5402 14867
rect 5430 14811 5486 14867
rect 5514 14811 5570 14867
rect 5598 14811 5654 14867
rect 4672 14667 4728 14723
rect 4757 14667 4813 14723
rect 4842 14667 4898 14723
rect 4926 14667 4982 14723
rect 5010 14667 5066 14723
rect 5094 14667 5150 14723
rect 5178 14667 5234 14723
rect 5262 14667 5318 14723
rect 5346 14667 5402 14723
rect 5430 14667 5486 14723
rect 5514 14667 5570 14723
rect 5598 14667 5654 14723
<< metal3 >>
rect 1583 25449 2383 40000
rect 1583 25393 1592 25449
rect 1648 25393 1673 25449
rect 1729 25393 1754 25449
rect 1810 25393 1835 25449
rect 1891 25393 1916 25449
rect 1972 25393 1997 25449
rect 2053 25393 2078 25449
rect 1583 25369 2078 25393
rect 1583 25313 1592 25369
rect 1648 25313 1673 25369
rect 1729 25313 1754 25369
rect 1810 25313 1835 25369
rect 1891 25313 1916 25369
rect 1972 25313 1997 25369
rect 2053 25313 2078 25369
rect 1583 25289 2078 25313
rect 1583 25233 1592 25289
rect 1648 25233 1673 25289
rect 1729 25233 1754 25289
rect 1810 25233 1835 25289
rect 1891 25233 1916 25289
rect 1972 25233 1997 25289
rect 2053 25233 2078 25289
rect 1583 25209 2078 25233
rect 1583 25153 1592 25209
rect 1648 25153 1673 25209
rect 1729 25153 1754 25209
rect 1810 25153 1835 25209
rect 1891 25153 1916 25209
rect 1972 25153 1997 25209
rect 2053 25153 2078 25209
rect 2374 25153 2383 25449
rect 1583 0 2383 25153
rect 3703 28185 4503 40000
rect 3703 28129 3712 28185
rect 3768 28129 3793 28185
rect 3849 28129 3874 28185
rect 3930 28129 3955 28185
rect 4011 28129 4036 28185
rect 4092 28129 4117 28185
rect 4173 28129 4198 28185
rect 4254 28129 4278 28185
rect 4334 28129 4358 28185
rect 4414 28129 4438 28185
rect 4494 28129 4503 28185
rect 3703 23814 4503 28129
rect 3703 23758 3712 23814
rect 3768 23758 3793 23814
rect 3849 23758 3874 23814
rect 3930 23758 3955 23814
rect 4011 23758 4036 23814
rect 4092 23758 4117 23814
rect 4173 23758 4198 23814
rect 4254 23758 4278 23814
rect 4334 23758 4358 23814
rect 4414 23758 4438 23814
rect 4494 23758 4503 23814
rect 3703 20419 4503 23758
rect 3703 20363 3712 20419
rect 3768 20363 3793 20419
rect 3849 20363 3874 20419
rect 3930 20363 3955 20419
rect 4011 20363 4036 20419
rect 4092 20363 4117 20419
rect 4173 20363 4198 20419
rect 4254 20363 4278 20419
rect 4334 20363 4358 20419
rect 4414 20363 4438 20419
rect 4494 20363 4503 20419
rect 3703 20024 4503 20363
rect 3703 19968 3712 20024
rect 3768 19968 3793 20024
rect 3849 19968 3874 20024
rect 3930 19968 3955 20024
rect 4011 19968 4036 20024
rect 4092 19968 4117 20024
rect 4173 19968 4198 20024
rect 4254 19968 4278 20024
rect 4334 19968 4358 20024
rect 4414 19968 4438 20024
rect 4494 19968 4503 20024
rect 3703 18300 4503 19968
rect 3703 18244 3712 18300
rect 3768 18244 3793 18300
rect 3849 18244 3874 18300
rect 3930 18244 3955 18300
rect 4011 18244 4036 18300
rect 4092 18244 4117 18300
rect 4173 18244 4198 18300
rect 4254 18244 4278 18300
rect 4334 18244 4358 18300
rect 4414 18244 4438 18300
rect 4494 18244 4503 18300
rect 3703 0 4503 18244
rect 4663 39192 5663 40000
rect 4663 36416 4775 39192
rect 5551 36416 5663 39192
rect 4663 36391 5663 36416
rect 4663 36335 4775 36391
rect 4831 36335 4855 36391
rect 4911 36335 4935 36391
rect 4991 36335 5015 36391
rect 5071 36335 5095 36391
rect 5151 36335 5175 36391
rect 5231 36335 5255 36391
rect 5311 36335 5335 36391
rect 5391 36335 5415 36391
rect 5471 36335 5495 36391
rect 5551 36335 5663 36391
rect 4663 36310 5663 36335
rect 4663 36254 4775 36310
rect 4831 36254 4855 36310
rect 4911 36254 4935 36310
rect 4991 36254 5015 36310
rect 5071 36254 5095 36310
rect 5151 36254 5175 36310
rect 5231 36254 5255 36310
rect 5311 36254 5335 36310
rect 5391 36254 5415 36310
rect 5471 36254 5495 36310
rect 5551 36254 5663 36310
rect 4663 36229 5663 36254
rect 4663 36173 4775 36229
rect 4831 36173 4855 36229
rect 4911 36173 4935 36229
rect 4991 36173 5015 36229
rect 5071 36173 5095 36229
rect 5151 36173 5175 36229
rect 5231 36173 5255 36229
rect 5311 36173 5335 36229
rect 5391 36173 5415 36229
rect 5471 36173 5495 36229
rect 5551 36173 5663 36229
rect 4663 36148 5663 36173
rect 4663 36092 4775 36148
rect 4831 36092 4855 36148
rect 4911 36092 4935 36148
rect 4991 36092 5015 36148
rect 5071 36092 5095 36148
rect 5151 36092 5175 36148
rect 5231 36092 5255 36148
rect 5311 36092 5335 36148
rect 5391 36092 5415 36148
rect 5471 36092 5495 36148
rect 5551 36092 5663 36148
rect 4663 36067 5663 36092
rect 4663 36011 4775 36067
rect 4831 36011 4855 36067
rect 4911 36011 4935 36067
rect 4991 36011 5015 36067
rect 5071 36011 5095 36067
rect 5151 36011 5175 36067
rect 5231 36011 5255 36067
rect 5311 36011 5335 36067
rect 5391 36011 5415 36067
rect 5471 36011 5495 36067
rect 5551 36011 5663 36067
rect 4663 35986 5663 36011
rect 4663 35930 4775 35986
rect 4831 35930 4855 35986
rect 4911 35930 4935 35986
rect 4991 35930 5015 35986
rect 5071 35930 5095 35986
rect 5151 35930 5175 35986
rect 5231 35930 5255 35986
rect 5311 35930 5335 35986
rect 5391 35930 5415 35986
rect 5471 35930 5495 35986
rect 5551 35930 5663 35986
rect 4663 35905 5663 35930
rect 4663 35849 4775 35905
rect 4831 35849 4855 35905
rect 4911 35849 4935 35905
rect 4991 35849 5015 35905
rect 5071 35849 5095 35905
rect 5151 35849 5175 35905
rect 5231 35849 5255 35905
rect 5311 35849 5335 35905
rect 5391 35849 5415 35905
rect 5471 35849 5495 35905
rect 5551 35849 5663 35905
rect 4663 35824 5663 35849
rect 4663 35768 4775 35824
rect 4831 35768 4855 35824
rect 4911 35768 4935 35824
rect 4991 35768 5015 35824
rect 5071 35768 5095 35824
rect 5151 35768 5175 35824
rect 5231 35768 5255 35824
rect 5311 35768 5335 35824
rect 5391 35768 5415 35824
rect 5471 35768 5495 35824
rect 5551 35768 5663 35824
rect 4663 35743 5663 35768
rect 4663 35687 4775 35743
rect 4831 35687 4855 35743
rect 4911 35687 4935 35743
rect 4991 35687 5015 35743
rect 5071 35687 5095 35743
rect 5151 35687 5175 35743
rect 5231 35687 5255 35743
rect 5311 35687 5335 35743
rect 5391 35687 5415 35743
rect 5471 35687 5495 35743
rect 5551 35687 5663 35743
rect 4663 35662 5663 35687
rect 4663 35606 4775 35662
rect 4831 35606 4855 35662
rect 4911 35606 4935 35662
rect 4991 35606 5015 35662
rect 5071 35606 5095 35662
rect 5151 35606 5175 35662
rect 5231 35606 5255 35662
rect 5311 35606 5335 35662
rect 5391 35606 5415 35662
rect 5471 35606 5495 35662
rect 5551 35606 5663 35662
rect 4663 35581 5663 35606
rect 4663 35525 4775 35581
rect 4831 35525 4855 35581
rect 4911 35525 4935 35581
rect 4991 35525 5015 35581
rect 5071 35525 5095 35581
rect 5151 35525 5175 35581
rect 5231 35525 5255 35581
rect 5311 35525 5335 35581
rect 5391 35525 5415 35581
rect 5471 35525 5495 35581
rect 5551 35525 5663 35581
rect 4663 35500 5663 35525
rect 4663 35444 4775 35500
rect 4831 35444 4855 35500
rect 4911 35444 4935 35500
rect 4991 35444 5015 35500
rect 5071 35444 5095 35500
rect 5151 35444 5175 35500
rect 5231 35444 5255 35500
rect 5311 35444 5335 35500
rect 5391 35444 5415 35500
rect 5471 35444 5495 35500
rect 5551 35444 5663 35500
rect 4663 35419 5663 35444
rect 4663 35363 4775 35419
rect 4831 35363 4855 35419
rect 4911 35363 4935 35419
rect 4991 35363 5015 35419
rect 5071 35363 5095 35419
rect 5151 35363 5175 35419
rect 5231 35363 5255 35419
rect 5311 35363 5335 35419
rect 5391 35363 5415 35419
rect 5471 35363 5495 35419
rect 5551 35363 5663 35419
rect 4663 35338 5663 35363
rect 4663 35282 4775 35338
rect 4831 35282 4855 35338
rect 4911 35282 4935 35338
rect 4991 35282 5015 35338
rect 5071 35282 5095 35338
rect 5151 35282 5175 35338
rect 5231 35282 5255 35338
rect 5311 35282 5335 35338
rect 5391 35282 5415 35338
rect 5471 35282 5495 35338
rect 5551 35282 5663 35338
rect 4663 35257 5663 35282
rect 4663 35201 4775 35257
rect 4831 35201 4855 35257
rect 4911 35201 4935 35257
rect 4991 35201 5015 35257
rect 5071 35201 5095 35257
rect 5151 35201 5175 35257
rect 5231 35201 5255 35257
rect 5311 35201 5335 35257
rect 5391 35201 5415 35257
rect 5471 35201 5495 35257
rect 5551 35201 5663 35257
rect 4663 35176 5663 35201
rect 4663 35120 4775 35176
rect 4831 35120 4855 35176
rect 4911 35120 4935 35176
rect 4991 35120 5015 35176
rect 5071 35120 5095 35176
rect 5151 35120 5175 35176
rect 5231 35120 5255 35176
rect 5311 35120 5335 35176
rect 5391 35120 5415 35176
rect 5471 35120 5495 35176
rect 5551 35120 5663 35176
rect 4663 35095 5663 35120
rect 4663 35039 4775 35095
rect 4831 35039 4855 35095
rect 4911 35039 4935 35095
rect 4991 35039 5015 35095
rect 5071 35039 5095 35095
rect 5151 35039 5175 35095
rect 5231 35039 5255 35095
rect 5311 35039 5335 35095
rect 5391 35039 5415 35095
rect 5471 35039 5495 35095
rect 5551 35039 5663 35095
rect 4663 35014 5663 35039
rect 4663 34958 4775 35014
rect 4831 34958 4855 35014
rect 4911 34958 4935 35014
rect 4991 34958 5015 35014
rect 5071 34958 5095 35014
rect 5151 34958 5175 35014
rect 5231 34958 5255 35014
rect 5311 34958 5335 35014
rect 5391 34958 5415 35014
rect 5471 34958 5495 35014
rect 5551 34958 5663 35014
rect 4663 34933 5663 34958
rect 4663 34877 4775 34933
rect 4831 34877 4855 34933
rect 4911 34877 4935 34933
rect 4991 34877 5015 34933
rect 5071 34877 5095 34933
rect 5151 34877 5175 34933
rect 5231 34877 5255 34933
rect 5311 34877 5335 34933
rect 5391 34877 5415 34933
rect 5471 34877 5495 34933
rect 5551 34877 5663 34933
rect 4663 34852 5663 34877
rect 4663 34796 4775 34852
rect 4831 34796 4855 34852
rect 4911 34796 4935 34852
rect 4991 34796 5015 34852
rect 5071 34796 5095 34852
rect 5151 34796 5175 34852
rect 5231 34796 5255 34852
rect 5311 34796 5335 34852
rect 5391 34796 5415 34852
rect 5471 34796 5495 34852
rect 5551 34796 5663 34852
rect 4663 34771 5663 34796
rect 4663 34715 4775 34771
rect 4831 34715 4855 34771
rect 4911 34715 4935 34771
rect 4991 34715 5015 34771
rect 5071 34715 5095 34771
rect 5151 34715 5175 34771
rect 5231 34715 5255 34771
rect 5311 34715 5335 34771
rect 5391 34715 5415 34771
rect 5471 34715 5495 34771
rect 5551 34715 5663 34771
rect 4663 34690 5663 34715
rect 4663 34634 4775 34690
rect 4831 34634 4855 34690
rect 4911 34634 4935 34690
rect 4991 34634 5015 34690
rect 5071 34634 5095 34690
rect 5151 34634 5175 34690
rect 5231 34634 5255 34690
rect 5311 34634 5335 34690
rect 5391 34634 5415 34690
rect 5471 34634 5495 34690
rect 5551 34634 5663 34690
rect 4663 34609 5663 34634
rect 4663 34553 4775 34609
rect 4831 34553 4855 34609
rect 4911 34553 4935 34609
rect 4991 34553 5015 34609
rect 5071 34553 5095 34609
rect 5151 34553 5175 34609
rect 5231 34553 5255 34609
rect 5311 34553 5335 34609
rect 5391 34553 5415 34609
rect 5471 34553 5495 34609
rect 5551 34553 5663 34609
rect 4663 34528 5663 34553
rect 4663 34472 4775 34528
rect 4831 34472 4855 34528
rect 4911 34472 4935 34528
rect 4991 34472 5015 34528
rect 5071 34472 5095 34528
rect 5151 34472 5175 34528
rect 5231 34472 5255 34528
rect 5311 34472 5335 34528
rect 5391 34472 5415 34528
rect 5471 34472 5495 34528
rect 5551 34472 5663 34528
rect 4663 34447 5663 34472
rect 4663 34391 4775 34447
rect 4831 34391 4855 34447
rect 4911 34391 4935 34447
rect 4991 34391 5015 34447
rect 5071 34391 5095 34447
rect 5151 34391 5175 34447
rect 5231 34391 5255 34447
rect 5311 34391 5335 34447
rect 5391 34391 5415 34447
rect 5471 34391 5495 34447
rect 5551 34391 5663 34447
rect 4663 34366 5663 34391
rect 4663 34310 4775 34366
rect 4831 34310 4855 34366
rect 4911 34310 4935 34366
rect 4991 34310 5015 34366
rect 5071 34310 5095 34366
rect 5151 34310 5175 34366
rect 5231 34310 5255 34366
rect 5311 34310 5335 34366
rect 5391 34310 5415 34366
rect 5471 34310 5495 34366
rect 5551 34310 5663 34366
rect 4663 34285 5663 34310
rect 4663 34229 4775 34285
rect 4831 34229 4855 34285
rect 4911 34229 4935 34285
rect 4991 34229 5015 34285
rect 5071 34229 5095 34285
rect 5151 34229 5175 34285
rect 5231 34229 5255 34285
rect 5311 34229 5335 34285
rect 5391 34229 5415 34285
rect 5471 34229 5495 34285
rect 5551 34229 5663 34285
rect 4663 34204 5663 34229
rect 4663 34148 4775 34204
rect 4831 34148 4855 34204
rect 4911 34148 4935 34204
rect 4991 34148 5015 34204
rect 5071 34148 5095 34204
rect 5151 34148 5175 34204
rect 5231 34148 5255 34204
rect 5311 34148 5335 34204
rect 5391 34148 5415 34204
rect 5471 34148 5495 34204
rect 5551 34148 5663 34204
rect 4663 34123 5663 34148
rect 4663 34067 4775 34123
rect 4831 34067 4855 34123
rect 4911 34067 4935 34123
rect 4991 34067 5015 34123
rect 5071 34067 5095 34123
rect 5151 34067 5175 34123
rect 5231 34067 5255 34123
rect 5311 34067 5335 34123
rect 5391 34067 5415 34123
rect 5471 34067 5495 34123
rect 5551 34067 5663 34123
rect 4663 34042 5663 34067
rect 4663 33986 4775 34042
rect 4831 33986 4855 34042
rect 4911 33986 4935 34042
rect 4991 33986 5015 34042
rect 5071 33986 5095 34042
rect 5151 33986 5175 34042
rect 5231 33986 5255 34042
rect 5311 33986 5335 34042
rect 5391 33986 5415 34042
rect 5471 33986 5495 34042
rect 5551 33986 5663 34042
rect 4663 33961 5663 33986
rect 4663 33905 4775 33961
rect 4831 33905 4855 33961
rect 4911 33905 4935 33961
rect 4991 33905 5015 33961
rect 5071 33905 5095 33961
rect 5151 33905 5175 33961
rect 5231 33905 5255 33961
rect 5311 33905 5335 33961
rect 5391 33905 5415 33961
rect 5471 33905 5495 33961
rect 5551 33905 5663 33961
rect 4663 33880 5663 33905
rect 4663 33824 4775 33880
rect 4831 33824 4855 33880
rect 4911 33824 4935 33880
rect 4991 33824 5015 33880
rect 5071 33824 5095 33880
rect 5151 33824 5175 33880
rect 5231 33824 5255 33880
rect 5311 33824 5335 33880
rect 5391 33824 5415 33880
rect 5471 33824 5495 33880
rect 5551 33824 5663 33880
rect 4663 33799 5663 33824
rect 4663 33743 4775 33799
rect 4831 33743 4855 33799
rect 4911 33743 4935 33799
rect 4991 33743 5015 33799
rect 5071 33743 5095 33799
rect 5151 33743 5175 33799
rect 5231 33743 5255 33799
rect 5311 33743 5335 33799
rect 5391 33743 5415 33799
rect 5471 33743 5495 33799
rect 5551 33743 5663 33799
rect 4663 33718 5663 33743
rect 4663 33662 4775 33718
rect 4831 33662 4855 33718
rect 4911 33662 4935 33718
rect 4991 33662 5015 33718
rect 5071 33662 5095 33718
rect 5151 33662 5175 33718
rect 5231 33662 5255 33718
rect 5311 33662 5335 33718
rect 5391 33662 5415 33718
rect 5471 33662 5495 33718
rect 5551 33662 5663 33718
rect 4663 33637 5663 33662
rect 4663 33581 4775 33637
rect 4831 33581 4855 33637
rect 4911 33581 4935 33637
rect 4991 33581 5015 33637
rect 5071 33581 5095 33637
rect 5151 33581 5175 33637
rect 5231 33581 5255 33637
rect 5311 33581 5335 33637
rect 5391 33581 5415 33637
rect 5471 33581 5495 33637
rect 5551 33581 5663 33637
rect 4663 33556 5663 33581
rect 4663 33500 4775 33556
rect 4831 33500 4855 33556
rect 4911 33500 4935 33556
rect 4991 33500 5015 33556
rect 5071 33500 5095 33556
rect 5151 33500 5175 33556
rect 5231 33500 5255 33556
rect 5311 33500 5335 33556
rect 5391 33500 5415 33556
rect 5471 33500 5495 33556
rect 5551 33500 5663 33556
rect 4663 33475 5663 33500
rect 4663 33419 4775 33475
rect 4831 33419 4855 33475
rect 4911 33419 4935 33475
rect 4991 33419 5015 33475
rect 5071 33419 5095 33475
rect 5151 33419 5175 33475
rect 5231 33419 5255 33475
rect 5311 33419 5335 33475
rect 5391 33419 5415 33475
rect 5471 33419 5495 33475
rect 5551 33419 5663 33475
rect 4663 33394 5663 33419
rect 4663 33338 4775 33394
rect 4831 33338 4855 33394
rect 4911 33338 4935 33394
rect 4991 33338 5015 33394
rect 5071 33338 5095 33394
rect 5151 33338 5175 33394
rect 5231 33338 5255 33394
rect 5311 33338 5335 33394
rect 5391 33338 5415 33394
rect 5471 33338 5495 33394
rect 5551 33338 5663 33394
rect 4663 33313 5663 33338
rect 4663 33257 4775 33313
rect 4831 33257 4855 33313
rect 4911 33257 4935 33313
rect 4991 33257 5015 33313
rect 5071 33257 5095 33313
rect 5151 33257 5175 33313
rect 5231 33257 5255 33313
rect 5311 33257 5335 33313
rect 5391 33257 5415 33313
rect 5471 33257 5495 33313
rect 5551 33257 5663 33313
rect 4663 33232 5663 33257
rect 4663 33176 4775 33232
rect 4831 33176 4855 33232
rect 4911 33176 4935 33232
rect 4991 33176 5015 33232
rect 5071 33176 5095 33232
rect 5151 33176 5175 33232
rect 5231 33176 5255 33232
rect 5311 33176 5335 33232
rect 5391 33176 5415 33232
rect 5471 33176 5495 33232
rect 5551 33176 5663 33232
rect 4663 33151 5663 33176
rect 4663 33095 4775 33151
rect 4831 33095 4855 33151
rect 4911 33095 4935 33151
rect 4991 33095 5015 33151
rect 5071 33095 5095 33151
rect 5151 33095 5175 33151
rect 5231 33095 5255 33151
rect 5311 33095 5335 33151
rect 5391 33095 5415 33151
rect 5471 33095 5495 33151
rect 5551 33095 5663 33151
rect 4663 33070 5663 33095
rect 4663 33014 4775 33070
rect 4831 33014 4855 33070
rect 4911 33014 4935 33070
rect 4991 33014 5015 33070
rect 5071 33014 5095 33070
rect 5151 33014 5175 33070
rect 5231 33014 5255 33070
rect 5311 33014 5335 33070
rect 5391 33014 5415 33070
rect 5471 33014 5495 33070
rect 5551 33014 5663 33070
rect 4663 32989 5663 33014
rect 4663 32933 4775 32989
rect 4831 32933 4855 32989
rect 4911 32933 4935 32989
rect 4991 32933 5015 32989
rect 5071 32933 5095 32989
rect 5151 32933 5175 32989
rect 5231 32933 5255 32989
rect 5311 32933 5335 32989
rect 5391 32933 5415 32989
rect 5471 32933 5495 32989
rect 5551 32933 5663 32989
rect 4663 32908 5663 32933
rect 4663 32852 4775 32908
rect 4831 32852 4855 32908
rect 4911 32852 4935 32908
rect 4991 32852 5015 32908
rect 5071 32852 5095 32908
rect 5151 32852 5175 32908
rect 5231 32852 5255 32908
rect 5311 32852 5335 32908
rect 5391 32852 5415 32908
rect 5471 32852 5495 32908
rect 5551 32852 5663 32908
rect 4663 32827 5663 32852
rect 4663 32771 4775 32827
rect 4831 32771 4855 32827
rect 4911 32771 4935 32827
rect 4991 32771 5015 32827
rect 5071 32771 5095 32827
rect 5151 32771 5175 32827
rect 5231 32771 5255 32827
rect 5311 32771 5335 32827
rect 5391 32771 5415 32827
rect 5471 32771 5495 32827
rect 5551 32771 5663 32827
rect 4663 32746 5663 32771
rect 4663 32690 4775 32746
rect 4831 32690 4855 32746
rect 4911 32690 4935 32746
rect 4991 32690 5015 32746
rect 5071 32690 5095 32746
rect 5151 32690 5175 32746
rect 5231 32690 5255 32746
rect 5311 32690 5335 32746
rect 5391 32690 5415 32746
rect 5471 32690 5495 32746
rect 5551 32690 5663 32746
rect 4663 32665 5663 32690
rect 4663 32609 4775 32665
rect 4831 32609 4855 32665
rect 4911 32609 4935 32665
rect 4991 32609 5015 32665
rect 5071 32609 5095 32665
rect 5151 32609 5175 32665
rect 5231 32609 5255 32665
rect 5311 32609 5335 32665
rect 5391 32609 5415 32665
rect 5471 32609 5495 32665
rect 5551 32609 5663 32665
rect 4663 32584 5663 32609
rect 4663 32528 4775 32584
rect 4831 32528 4855 32584
rect 4911 32528 4935 32584
rect 4991 32528 5015 32584
rect 5071 32528 5095 32584
rect 5151 32528 5175 32584
rect 5231 32528 5255 32584
rect 5311 32528 5335 32584
rect 5391 32528 5415 32584
rect 5471 32528 5495 32584
rect 5551 32528 5663 32584
rect 4663 32503 5663 32528
rect 4663 32447 4775 32503
rect 4831 32447 4855 32503
rect 4911 32447 4935 32503
rect 4991 32447 5015 32503
rect 5071 32447 5095 32503
rect 5151 32447 5175 32503
rect 5231 32447 5255 32503
rect 5311 32447 5335 32503
rect 5391 32447 5415 32503
rect 5471 32447 5495 32503
rect 5551 32447 5663 32503
rect 4663 32422 5663 32447
rect 4663 32366 4775 32422
rect 4831 32366 4855 32422
rect 4911 32366 4935 32422
rect 4991 32366 5015 32422
rect 5071 32366 5095 32422
rect 5151 32366 5175 32422
rect 5231 32366 5255 32422
rect 5311 32366 5335 32422
rect 5391 32366 5415 32422
rect 5471 32366 5495 32422
rect 5551 32366 5663 32422
rect 4663 32341 5663 32366
rect 4663 32285 4775 32341
rect 4831 32285 4855 32341
rect 4911 32285 4935 32341
rect 4991 32285 5015 32341
rect 5071 32285 5095 32341
rect 5151 32285 5175 32341
rect 5231 32285 5255 32341
rect 5311 32285 5335 32341
rect 5391 32285 5415 32341
rect 5471 32285 5495 32341
rect 5551 32285 5663 32341
rect 4663 32260 5663 32285
rect 4663 32204 4775 32260
rect 4831 32204 4855 32260
rect 4911 32204 4935 32260
rect 4991 32204 5015 32260
rect 5071 32204 5095 32260
rect 5151 32204 5175 32260
rect 5231 32204 5255 32260
rect 5311 32204 5335 32260
rect 5391 32204 5415 32260
rect 5471 32204 5495 32260
rect 5551 32204 5663 32260
rect 4663 32179 5663 32204
rect 4663 32123 4775 32179
rect 4831 32123 4855 32179
rect 4911 32123 4935 32179
rect 4991 32123 5015 32179
rect 5071 32123 5095 32179
rect 5151 32123 5175 32179
rect 5231 32123 5255 32179
rect 5311 32123 5335 32179
rect 5391 32123 5415 32179
rect 5471 32123 5495 32179
rect 5551 32123 5663 32179
rect 4663 32098 5663 32123
rect 4663 32042 4775 32098
rect 4831 32042 4855 32098
rect 4911 32042 4935 32098
rect 4991 32042 5015 32098
rect 5071 32042 5095 32098
rect 5151 32042 5175 32098
rect 5231 32042 5255 32098
rect 5311 32042 5335 32098
rect 5391 32042 5415 32098
rect 5471 32042 5495 32098
rect 5551 32042 5663 32098
rect 4663 32017 5663 32042
rect 4663 31961 4775 32017
rect 4831 31961 4855 32017
rect 4911 31961 4935 32017
rect 4991 31961 5015 32017
rect 5071 31961 5095 32017
rect 5151 31961 5175 32017
rect 5231 31961 5255 32017
rect 5311 31961 5335 32017
rect 5391 31961 5415 32017
rect 5471 31961 5495 32017
rect 5551 31961 5663 32017
rect 4663 31936 5663 31961
rect 4663 31880 4775 31936
rect 4831 31880 4855 31936
rect 4911 31880 4935 31936
rect 4991 31880 5015 31936
rect 5071 31880 5095 31936
rect 5151 31880 5175 31936
rect 5231 31880 5255 31936
rect 5311 31880 5335 31936
rect 5391 31880 5415 31936
rect 5471 31880 5495 31936
rect 5551 31880 5663 31936
rect 4663 31855 5663 31880
rect 4663 31799 4775 31855
rect 4831 31799 4855 31855
rect 4911 31799 4935 31855
rect 4991 31799 5015 31855
rect 5071 31799 5095 31855
rect 5151 31799 5175 31855
rect 5231 31799 5255 31855
rect 5311 31799 5335 31855
rect 5391 31799 5415 31855
rect 5471 31799 5495 31855
rect 5551 31799 5663 31855
rect 4663 31774 5663 31799
rect 4663 31718 4775 31774
rect 4831 31718 4855 31774
rect 4911 31718 4935 31774
rect 4991 31718 5015 31774
rect 5071 31718 5095 31774
rect 5151 31718 5175 31774
rect 5231 31718 5255 31774
rect 5311 31718 5335 31774
rect 5391 31718 5415 31774
rect 5471 31718 5495 31774
rect 5551 31718 5663 31774
rect 4663 31693 5663 31718
rect 4663 31637 4775 31693
rect 4831 31637 4855 31693
rect 4911 31637 4935 31693
rect 4991 31637 5015 31693
rect 5071 31637 5095 31693
rect 5151 31637 5175 31693
rect 5231 31637 5255 31693
rect 5311 31637 5335 31693
rect 5391 31637 5415 31693
rect 5471 31637 5495 31693
rect 5551 31637 5663 31693
rect 4663 31612 5663 31637
rect 4663 31556 4775 31612
rect 4831 31556 4855 31612
rect 4911 31556 4935 31612
rect 4991 31556 5015 31612
rect 5071 31556 5095 31612
rect 5151 31556 5175 31612
rect 5231 31556 5255 31612
rect 5311 31556 5335 31612
rect 5391 31556 5415 31612
rect 5471 31556 5495 31612
rect 5551 31556 5663 31612
rect 4663 31531 5663 31556
rect 4663 31475 4775 31531
rect 4831 31475 4855 31531
rect 4911 31475 4935 31531
rect 4991 31475 5015 31531
rect 5071 31475 5095 31531
rect 5151 31475 5175 31531
rect 5231 31475 5255 31531
rect 5311 31475 5335 31531
rect 5391 31475 5415 31531
rect 5471 31475 5495 31531
rect 5551 31475 5663 31531
rect 4663 31450 5663 31475
rect 4663 31394 4775 31450
rect 4831 31394 4855 31450
rect 4911 31394 4935 31450
rect 4991 31394 5015 31450
rect 5071 31394 5095 31450
rect 5151 31394 5175 31450
rect 5231 31394 5255 31450
rect 5311 31394 5335 31450
rect 5391 31394 5415 31450
rect 5471 31394 5495 31450
rect 5551 31394 5663 31450
rect 4663 31369 5663 31394
rect 4663 31313 4775 31369
rect 4831 31313 4855 31369
rect 4911 31313 4935 31369
rect 4991 31313 5015 31369
rect 5071 31313 5095 31369
rect 5151 31313 5175 31369
rect 5231 31313 5255 31369
rect 5311 31313 5335 31369
rect 5391 31313 5415 31369
rect 5471 31313 5495 31369
rect 5551 31313 5663 31369
rect 4663 31288 5663 31313
rect 4663 31232 4775 31288
rect 4831 31232 4855 31288
rect 4911 31232 4935 31288
rect 4991 31232 5015 31288
rect 5071 31232 5095 31288
rect 5151 31232 5175 31288
rect 5231 31232 5255 31288
rect 5311 31232 5335 31288
rect 5391 31232 5415 31288
rect 5471 31232 5495 31288
rect 5551 31232 5663 31288
rect 4663 31207 5663 31232
rect 4663 31151 4775 31207
rect 4831 31151 4855 31207
rect 4911 31151 4935 31207
rect 4991 31151 5015 31207
rect 5071 31151 5095 31207
rect 5151 31151 5175 31207
rect 5231 31151 5255 31207
rect 5311 31151 5335 31207
rect 5391 31151 5415 31207
rect 5471 31151 5495 31207
rect 5551 31151 5663 31207
rect 4663 31126 5663 31151
rect 4663 31070 4775 31126
rect 4831 31070 4855 31126
rect 4911 31070 4935 31126
rect 4991 31070 5015 31126
rect 5071 31070 5095 31126
rect 5151 31070 5175 31126
rect 5231 31070 5255 31126
rect 5311 31070 5335 31126
rect 5391 31070 5415 31126
rect 5471 31070 5495 31126
rect 5551 31070 5663 31126
rect 4663 31045 5663 31070
rect 4663 30989 4775 31045
rect 4831 30989 4855 31045
rect 4911 30989 4935 31045
rect 4991 30989 5015 31045
rect 5071 30989 5095 31045
rect 5151 30989 5175 31045
rect 5231 30989 5255 31045
rect 5311 30989 5335 31045
rect 5391 30989 5415 31045
rect 5471 30989 5495 31045
rect 5551 30989 5663 31045
rect 4663 30964 5663 30989
rect 4663 30908 4775 30964
rect 4831 30908 4855 30964
rect 4911 30908 4935 30964
rect 4991 30908 5015 30964
rect 5071 30908 5095 30964
rect 5151 30908 5175 30964
rect 5231 30908 5255 30964
rect 5311 30908 5335 30964
rect 5391 30908 5415 30964
rect 5471 30908 5495 30964
rect 5551 30908 5663 30964
rect 4663 30883 5663 30908
rect 4663 30827 4775 30883
rect 4831 30827 4855 30883
rect 4911 30827 4935 30883
rect 4991 30827 5015 30883
rect 5071 30827 5095 30883
rect 5151 30827 5175 30883
rect 5231 30827 5255 30883
rect 5311 30827 5335 30883
rect 5391 30827 5415 30883
rect 5471 30827 5495 30883
rect 5551 30827 5663 30883
rect 4663 30802 5663 30827
rect 4663 30746 4775 30802
rect 4831 30746 4855 30802
rect 4911 30746 4935 30802
rect 4991 30746 5015 30802
rect 5071 30746 5095 30802
rect 5151 30746 5175 30802
rect 5231 30746 5255 30802
rect 5311 30746 5335 30802
rect 5391 30746 5415 30802
rect 5471 30746 5495 30802
rect 5551 30746 5663 30802
rect 4663 30721 5663 30746
rect 4663 30665 4775 30721
rect 4831 30665 4855 30721
rect 4911 30665 4935 30721
rect 4991 30665 5015 30721
rect 5071 30665 5095 30721
rect 5151 30665 5175 30721
rect 5231 30665 5255 30721
rect 5311 30665 5335 30721
rect 5391 30665 5415 30721
rect 5471 30665 5495 30721
rect 5551 30665 5663 30721
rect 4663 30640 5663 30665
rect 4663 30584 4775 30640
rect 4831 30584 4855 30640
rect 4911 30584 4935 30640
rect 4991 30584 5015 30640
rect 5071 30584 5095 30640
rect 5151 30584 5175 30640
rect 5231 30584 5255 30640
rect 5311 30584 5335 30640
rect 5391 30584 5415 30640
rect 5471 30584 5495 30640
rect 5551 30584 5663 30640
rect 4663 30559 5663 30584
rect 4663 30503 4775 30559
rect 4831 30503 4855 30559
rect 4911 30503 4935 30559
rect 4991 30503 5015 30559
rect 5071 30503 5095 30559
rect 5151 30503 5175 30559
rect 5231 30503 5255 30559
rect 5311 30503 5335 30559
rect 5391 30503 5415 30559
rect 5471 30503 5495 30559
rect 5551 30503 5663 30559
rect 4663 30478 5663 30503
rect 4663 30422 4775 30478
rect 4831 30422 4855 30478
rect 4911 30422 4935 30478
rect 4991 30422 5015 30478
rect 5071 30422 5095 30478
rect 5151 30422 5175 30478
rect 5231 30422 5255 30478
rect 5311 30422 5335 30478
rect 5391 30422 5415 30478
rect 5471 30422 5495 30478
rect 5551 30422 5663 30478
rect 4663 30397 5663 30422
rect 4663 30341 4775 30397
rect 4831 30341 4855 30397
rect 4911 30341 4935 30397
rect 4991 30341 5015 30397
rect 5071 30341 5095 30397
rect 5151 30341 5175 30397
rect 5231 30341 5255 30397
rect 5311 30341 5335 30397
rect 5391 30341 5415 30397
rect 5471 30341 5495 30397
rect 5551 30341 5663 30397
rect 4663 29875 5663 30341
rect 4663 29819 4672 29875
rect 4728 29819 4757 29875
rect 4813 29819 4842 29875
rect 4898 29819 4926 29875
rect 4982 29819 5010 29875
rect 5066 29819 5094 29875
rect 5150 29819 5178 29875
rect 5234 29819 5262 29875
rect 5318 29819 5346 29875
rect 5402 29819 5430 29875
rect 5486 29819 5514 29875
rect 5570 29819 5598 29875
rect 5654 29819 5663 29875
rect 4663 28891 5663 29819
rect 4663 28835 4672 28891
rect 4728 28835 4757 28891
rect 4813 28835 4842 28891
rect 4898 28835 4926 28891
rect 4982 28835 5010 28891
rect 5066 28835 5094 28891
rect 5150 28835 5178 28891
rect 5234 28835 5262 28891
rect 5318 28835 5346 28891
rect 5402 28835 5430 28891
rect 5486 28835 5514 28891
rect 5570 28835 5598 28891
rect 5654 28835 5663 28891
rect 4663 28445 5663 28835
rect 4663 28389 4672 28445
rect 4728 28389 4757 28445
rect 4813 28389 4842 28445
rect 4898 28389 4926 28445
rect 4982 28389 5010 28445
rect 5066 28389 5094 28445
rect 5150 28389 5178 28445
rect 5234 28389 5262 28445
rect 5318 28389 5346 28445
rect 5402 28389 5430 28445
rect 5486 28389 5514 28445
rect 5570 28389 5598 28445
rect 5654 28389 5663 28445
rect 4663 17895 5663 28389
rect 4663 17839 4672 17895
rect 4728 17839 4757 17895
rect 4813 17839 4842 17895
rect 4898 17839 4926 17895
rect 4982 17839 5010 17895
rect 5066 17839 5094 17895
rect 5150 17839 5178 17895
rect 5234 17839 5262 17895
rect 5318 17839 5346 17895
rect 5402 17839 5430 17895
rect 5486 17839 5514 17895
rect 5570 17839 5598 17895
rect 5654 17839 5663 17895
rect 4663 14867 5663 17839
rect 4663 14811 4672 14867
rect 4728 14811 4757 14867
rect 4813 14811 4842 14867
rect 4898 14811 4926 14867
rect 4982 14811 5010 14867
rect 5066 14811 5094 14867
rect 5150 14811 5178 14867
rect 5234 14811 5262 14867
rect 5318 14811 5346 14867
rect 5402 14811 5430 14867
rect 5486 14811 5514 14867
rect 5570 14811 5598 14867
rect 5654 14811 5663 14867
rect 4663 14723 5663 14811
rect 4663 14667 4672 14723
rect 4728 14667 4757 14723
rect 4813 14667 4842 14723
rect 4898 14667 4926 14723
rect 4982 14667 5010 14723
rect 5066 14667 5094 14723
rect 5150 14667 5178 14723
rect 5234 14667 5262 14723
rect 5318 14667 5346 14723
rect 5402 14667 5430 14723
rect 5486 14667 5514 14723
rect 5570 14667 5598 14723
rect 5654 14667 5663 14723
rect 4663 0 5663 14667
use DFL1_CDNS_52468879185881  DFL1_CDNS_52468879185881_0
timestamp 1707688321
transform 0 -1 5404 1 0 19596
box 0 0 1 1
use DFL1_CDNS_52468879185881  DFL1_CDNS_52468879185881_1
timestamp 1707688321
transform 0 -1 5148 1 0 19596
box 0 0 1 1
use DFL1_CDNS_52468879185881  DFL1_CDNS_52468879185881_2
timestamp 1707688321
transform 0 -1 5148 1 0 23788
box 0 0 1 1
use DFL1_CDNS_52468879185881  DFL1_CDNS_52468879185881_3
timestamp 1707688321
transform 0 -1 5404 1 0 23788
box 0 0 1 1
use nfet_CDNS_52468879185886  nfet_CDNS_52468879185886_0
timestamp 1707688321
transform 1 0 6255 0 -1 29806
box -82 -32 338 182
use nfet_CDNS_52468879185887  nfet_CDNS_52468879185887_0
timestamp 1707688321
transform -1 0 5835 0 1 15413
box -82 -32 1682 632
use nfet_CDNS_52468879185887  nfet_CDNS_52468879185887_1
timestamp 1707688321
transform -1 0 5835 0 1 16143
box -82 -32 1682 632
use nfet_CDNS_52468879185887  nfet_CDNS_52468879185887_2
timestamp 1707688321
transform -1 0 5835 0 1 14683
box -82 -32 1682 632
use nfet_CDNS_52468879185888  nfet_CDNS_52468879185888_0
timestamp 1707688321
transform 0 -1 3784 1 0 17132
box -82 -32 650 182
use nfet_CDNS_52468879185889  nfet_CDNS_52468879185889_0
timestamp 1707688321
transform 0 1 3196 1 0 16015
box -82 -32 1682 232
use nfet_CDNS_52468879185890  nfet_CDNS_52468879185890_0
timestamp 1707688321
transform -1 0 5461 0 -1 17915
box -82 -32 650 1032
use nfet_CDNS_52468879185890  nfet_CDNS_52468879185890_1
timestamp 1707688321
transform -1 0 4837 0 -1 17915
box -82 -32 650 1032
use nfet_CDNS_52468879185891  nfet_CDNS_52468879185891_0
timestamp 1707688321
transform 1 0 3604 0 -1 29617
box -82 -32 1738 332
use nfet_CDNS_52468879185891  nfet_CDNS_52468879185891_1
timestamp 1707688321
transform 1 0 3604 0 -1 30041
box -82 -32 1738 332
use nfet_CDNS_52468879185891  nfet_CDNS_52468879185891_2
timestamp 1707688321
transform 1 0 3604 0 -1 29057
box -82 -32 1738 332
use nfet_CDNS_52468879185893  nfet_CDNS_52468879185893_0
timestamp 1707688321
transform 0 -1 5256 1 0 30383
box -82 -32 9146 2032
use pfet_CDNS_52468879185894  pfet_CDNS_52468879185894_0
timestamp 1707688321
transform 1 0 5042 0 1 18786
box -122 -66 322 266
use pfet_CDNS_52468879185895  pfet_CDNS_52468879185895_0
timestamp 1707688321
transform 1 0 7381 0 1 21652
box -122 -66 378 366
use pfet_CDNS_52468879185896  pfet_CDNS_52468879185896_0
timestamp 1707688321
transform 0 -1 4851 -1 0 20048
box -119 -66 687 366
use pfet_CDNS_52468879185897  pfet_CDNS_52468879185897_0
timestamp 1707688321
transform 0 -1 4840 -1 0 23717
box -119 -66 3375 266
use pfet_CDNS_52468879185898  pfet_CDNS_52468879185898_0
timestamp 1707688321
transform -1 0 5590 0 1 24717
box -122 -66 1314 1466
use pfet_CDNS_52468879185899  pfet_CDNS_52468879185899_0
timestamp 1707688321
transform 0 -1 5404 -1 0 23717
box -119 -66 4119 150
use pfet_CDNS_52468879185899  pfet_CDNS_52468879185899_1
timestamp 1707688321
transform 0 -1 5148 -1 0 23717
box -119 -66 4119 150
use s8_esd_res250only_small  s8_esd_res250only_small_0
timestamp 1707688321
transform 0 -1 4236 1 0 18468
box 0 0 2270 404
use sky130_fd_io__top_pwrdetv2_res3  sky130_fd_io__top_pwrdetv2_res3_0
timestamp 1707688321
transform 1 0 2696 0 1 18525
box 0 0 952 7015
<< labels >>
flabel comment s 4895 28361 4895 28361 0 FreeSans 1000 0 0 0 condiode
flabel comment s 4895 18105 4895 18105 0 FreeSans 1000 0 0 0 condiode
flabel metal1 s 3926 18476 4192 18528 3 FreeSans 520 0 0 0 vddio_q
port 1 nsew
flabel metal1 s 8803 18983 8909 19117 3 FreeSans 520 0 0 0 out
port 2 nsew
flabel metal1 s 8226 23009 8347 23101 3 FreeSans 520 0 0 0 rst_por_hv_n
port 3 nsew
flabel metal1 s 952 16988 952 16988 3 FreeSans 520 0 0 0 vddio_b
flabel metal3 s 4663 39534 5658 39838 3 FreeSans 520 0 0 0 vssa
port 5 nsew
flabel metal3 s 3703 39640 4503 39938 3 FreeSans 520 0 0 0 vddd
port 6 nsew
flabel metal3 s 1583 39724 2383 39999 3 FreeSans 520 0 0 0 vccd
port 7 nsew
flabel metal2 s 3652 29440 3652 29440 3 FreeSans 520 0 0 0 pre_out
flabel metal2 s 2652 16387 2652 16387 3 FreeSans 520 0 0 0 vddio_r
<< properties >>
string GDS_END 6669256
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 6117744
string path 70.975 453.225 70.975 456.800 169.175 456.800 169.175 358.150 70.975 358.150 70.975 453.225 
<< end >>
