magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect 604 1268 820 1540
<< poly >>
rect 859 1256 1059 1278
rect 859 1222 911 1256
rect 945 1222 979 1256
rect 1013 1222 1059 1256
rect 859 1206 1059 1222
rect 1115 1220 1151 1279
rect 1207 1220 1243 1278
rect 1109 1204 1266 1220
rect 1109 1170 1125 1204
rect 1159 1170 1193 1204
rect 1227 1170 1266 1204
rect 1109 1154 1266 1170
rect 1230 1112 1266 1154
rect 974 838 1174 860
rect 974 804 1056 838
rect 1090 804 1124 838
rect 1158 804 1174 838
rect 974 788 1174 804
<< polycont >>
rect 911 1222 945 1256
rect 979 1222 1013 1256
rect 1125 1170 1159 1204
rect 1193 1170 1227 1204
rect 1056 804 1090 838
rect 1124 804 1158 838
<< locali >>
rect 141 1387 175 1421
rect 1070 1418 1104 1456
rect 1254 1418 1288 1456
rect 814 1226 848 1306
rect 1162 1272 1197 1306
rect 607 1188 848 1226
rect 895 1222 911 1256
rect 945 1222 979 1256
rect 1013 1222 1029 1256
rect 1162 1238 1311 1272
rect 1109 1188 1125 1204
rect 607 1170 1125 1188
rect 1159 1170 1193 1204
rect 1227 1170 1243 1204
rect 607 1154 1243 1170
rect 875 860 981 1096
rect 1277 1089 1311 1238
rect 1185 1012 1219 1050
rect 1185 940 1219 978
rect 451 826 489 860
rect 909 826 947 860
rect 1040 804 1056 838
rect 1090 804 1124 838
rect 1158 804 1174 838
rect 921 552 955 586
rect 262 16 295 50
rect 534 16 567 50
<< viali >>
rect 1070 1456 1104 1490
rect 1070 1384 1104 1418
rect 1254 1456 1288 1490
rect 1254 1384 1288 1418
rect 1185 1050 1219 1084
rect 1185 978 1219 1012
rect 1185 906 1219 940
rect 417 826 451 860
rect 489 826 523 860
rect 875 826 909 860
rect 947 826 981 860
<< metal1 >>
rect 85 1490 1332 1574
rect 85 1456 1070 1490
rect 1104 1456 1254 1490
rect 1288 1456 1332 1490
rect 85 1418 1332 1456
rect 85 1384 1070 1418
rect 1104 1384 1254 1418
rect 1288 1384 1332 1418
rect 85 1372 1332 1384
rect 8 894 33 1096
rect 834 1084 1283 1096
rect 834 1050 1185 1084
rect 1219 1050 1283 1084
rect 834 1012 1283 1050
rect 834 978 1185 1012
rect 1219 978 1283 1012
rect 834 940 1283 978
rect 834 906 1185 940
rect 1219 906 1283 940
rect 834 894 1283 906
rect 405 860 993 866
rect 405 826 417 860
rect 451 826 489 860
rect 523 826 875 860
rect 909 826 947 860
rect 981 826 993 860
rect 405 820 993 826
rect 398 44 439 74
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1707688321
transform 0 1 1070 -1 0 1490
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1707688321
transform 0 1 1254 -1 0 1490
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1707688321
transform -1 0 981 0 1 826
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1707688321
transform 1 0 417 0 1 826
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1707688321
transform 0 1 1185 -1 0 1084
box 0 0 1 1
use nfet_CDNS_524688791851207  nfet_CDNS_524688791851207_0
timestamp 1707688321
transform -1 0 1174 0 -1 1086
box -79 -26 279 226
use nfet_CDNS_524688791851208  nfet_CDNS_524688791851208_0
timestamp 1707688321
transform 1 0 1230 0 -1 1086
box -79 -26 115 226
use pfet_CDNS_524688791851209  pfet_CDNS_524688791851209_0
timestamp 1707688321
transform -1 0 1059 0 -1 1504
box -89 -36 289 236
use pfet_CDNS_524688791851210  pfet_CDNS_524688791851210_0
timestamp 1707688321
transform 1 0 1115 0 -1 1504
box -89 -36 217 236
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1707688321
transform 0 1 1109 1 0 1154
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_1
timestamp 1707688321
transform 0 1 895 1 0 1206
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_2
timestamp 1707688321
transform 0 -1 1174 1 0 788
box 0 0 1 1
use sky130_fd_io__sio_com_inbuf_ls  sky130_fd_io__sio_com_inbuf_ls_0
timestamp 1707688321
transform 1 0 8 0 1 0
box -51 0 973 1574
<< labels >>
flabel comment s 277 10 277 10 0 FreeSans 200 0 0 0 in_t
flabel comment s 551 11 551 11 0 FreeSans 200 0 0 0 in_c
flabel metal1 s 85 1372 108 1574 3 FreeSans 400 0 0 0 vpwr
port 2 nsew
flabel metal1 s 398 44 439 74 0 FreeSans 200 0 0 0 en_h
port 1 nsew
flabel metal1 s 8 894 33 1096 3 FreeSans 400 0 0 0 vgnd
port 3 nsew
flabel locali s 141 1387 175 1421 0 FreeSans 200 0 0 0 vpb
port 5 nsew
flabel locali s 1277 1174 1311 1206 0 FreeSans 200 0 0 0 out_ls
port 6 nsew
flabel locali s 921 552 955 586 0 FreeSans 200 0 0 0 vgnd
port 3 nsew
flabel locali s 262 16 295 50 0 FreeSans 600 0 0 0 in_t
port 7 nsew
flabel locali s 534 16 567 50 0 FreeSans 600 0 0 0 in_c
port 8 nsew
flabel locali s 1090 804 1124 838 0 FreeSans 600 0 0 0 en_n
port 9 nsew
flabel locali s 945 1222 979 1256 0 FreeSans 600 0 0 0 en
port 10 nsew
<< properties >>
string GDS_END 85572256
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85569008
<< end >>
