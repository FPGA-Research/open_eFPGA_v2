magic
tech sky130A
timestamp 1707688321
<< viali >>
rect 0 0 233 53
<< metal1 >>
rect -6 53 239 56
rect -6 0 0 53
rect 233 0 239 53
rect -6 -3 239 0
<< properties >>
string GDS_END 86915622
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86914594
<< end >>
