##
## LEF for PtnCells ;
## created by Innovus v15.20-p005_1 on Mon Jun 14 18:20:56 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO N_term_RAM_IO
  CLASS BLOCK ;
  SIZE 100.2800 BY 30.2600 ;
  FOREIGN N_term_RAM_IO 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.89 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.3725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7555 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.921 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.712 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.2038 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.224 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 31.828 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 168.025 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 7.9650 0.0000 8.1350 0.3300 ;
    END
  END N1END[3]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.23005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.153 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.6124 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 43.015 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.4664 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.096 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 19.0374 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 89.9969 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 7.0450 0.0000 7.2150 0.3300 ;
    END
  END N1END[2]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.38045 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.977 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.5616 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 27.7305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5976 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.87 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 5.10786 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 21.5157 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 6.1250 0.0000 6.2950 0.3300 ;
    END
  END N1END[1]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.47305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7644 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.785 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met1  ;
    ANTENNAMAXAREACAR 11.923 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 56.1635 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.181761 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 5.2050 0.0000 5.3750 0.3300 ;
    END
  END N1END[0]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9276 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.5605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6719 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1885 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.768 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.6936 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 52.64 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 69.7733 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 372.799 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 16.7050 0.0000 16.8750 0.3300 ;
    END
  END N2MID[7]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.461 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.0224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8525 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.056 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.0546 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.232 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 48.3374 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 258.761 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 15.3250 0.0000 15.4950 0.3300 ;
    END
  END N2MID[6]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08545 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.277 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.346 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 11.4487 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 52.7956 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 14.4050 0.0000 14.5750 0.3300 ;
    END
  END N2MID[5]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.3884 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.8645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1072 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.418 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 9.83113 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 39.327 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 13.4850 0.0000 13.6550 0.3300 ;
    END
  END N2MID[4]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.4356 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 27.1005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4321 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.9895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.781 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.7748 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.936 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 65.8846 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 352.028 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 12.1050 0.0000 12.2750 0.3300 ;
    END
  END N2MID[3]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.5036 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.4405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1476 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.502 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 15.9896 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 71.7327 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 11.1850 0.0000 11.3550 0.3300 ;
    END
  END N2MID[2]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.53085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.7242 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.584 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met1  ;
    ANTENNAMAXAREACAR 5.38082 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 23.4528 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.181761 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 10.2650 0.0000 10.4350 0.3300 ;
    END
  END N2MID[1]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.6328 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.0865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1688 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.726 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 9.66132 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 43.8585 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 9.3450 0.0000 9.5150 0.3300 ;
    END
  END N2MID[0]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.02765 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.209 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.4635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.1465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.31 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.2726 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 39.728 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 84.1236 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 452.047 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 24.9850 0.0000 25.1550 0.3300 ;
    END
  END N2END[7]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.6832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.3385 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5712 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.502 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.0764 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 84.4497 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 24.0650 0.0000 24.2350 0.3300 ;
    END
  END N2END[6]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8843 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.2505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.287 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.664 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 28.3362 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 149.673 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 22.6850 0.0000 22.8550 0.3300 ;
    END
  END N2END[5]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.202 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3765 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.14635 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.24 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.1584 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.256 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 71.9324 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 389.041 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 21.7650 0.0000 21.9350 0.3300 ;
    END
  END N2END[4]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.99025 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.165 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.4792 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 42.3185 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.6234 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.999 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 20.2186 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 96.6447 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 20.8450 0.0000 21.0150 0.3300 ;
    END
  END N2END[3]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.91205 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.073 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0732 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.298 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 6.90409 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 30.4969 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 19.4650 0.0000 19.6350 0.3300 ;
    END
  END N2END[2]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.02765 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.209 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.156 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 4.20975 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 17.0252 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 18.5450 0.0000 18.7150 0.3300 ;
    END
  END N2END[1]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.5708 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.5 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 23.8072 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 113.528 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 17.6250 0.0000 17.7950 0.3300 ;
    END
  END N2END[0]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.81685 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.961 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5884 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1476 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.502 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 10.7431 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 48.5252 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 41.5450 0.0000 41.7150 0.3300 ;
    END
  END N4END[15]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.58565 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.689 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.168 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.7625 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2164 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.964 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 8.99969 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 40.9748 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 40.6250 0.0000 40.7950 0.3300 ;
    END
  END N4END[14]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.132 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.5455 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.5528 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.174 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 38.8538 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 186.852 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 39.7050 0.0000 39.8750 0.3300 ;
    END
  END N4END[13]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08545 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.277 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.346 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 9.82862 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 44.695 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 38.7850 0.0000 38.9550 0.3300 ;
    END
  END N4END[12]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.3272 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5585 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8994 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.261 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 20.2525 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 96.0723 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 37.4050 0.0000 37.5750 0.3300 ;
    END
  END N4END[11]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.3916 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.8805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.026 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.012 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 12.7343 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 59.2233 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 36.4850 0.0000 36.6550 0.3300 ;
    END
  END N4END[10]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08545 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.277 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.346 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 8.18208 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 36.4623 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 35.5650 0.0000 35.7350 0.3300 ;
    END
  END N4END[9]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.24185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.461 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4072 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.918 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 4.87138 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.9088 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 34.1850 0.0000 34.3550 0.3300 ;
    END
  END N4END[8]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.41225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.485 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.026 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.012 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 23.9695 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 115.399 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 33.2650 0.0000 33.4350 0.3300 ;
    END
  END N4END[7]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96985 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.141 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7816 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.788 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.822 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 7.18711 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 31.4874 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 32.3450 0.0000 32.5150 0.3300 ;
    END
  END N4END[6]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.2368 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.137 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.346 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.9292 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 85.1981 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 31.4250 0.0000 31.5950 0.3300 ;
    END
  END N4END[5]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.18405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.2728 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 31.2865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4072 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.918 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 6.87767 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 26.9151 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 30.0450 0.0000 30.2150 0.3300 ;
    END
  END N4END[4]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2904 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.216 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 11.1758 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 46.2736 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 29.1250 0.0000 29.2950 0.3300 ;
    END
  END N4END[3]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2664 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1688 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.726 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 10.8764 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 49.934 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 28.2050 0.0000 28.3750 0.3300 ;
    END
  END N4END[2]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7172 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5085 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4241 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.782 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.6488 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 41.264 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 79.7047 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 424.456 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 26.8250 0.0000 26.9950 0.3300 ;
    END
  END N4END[1]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.6528 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.774 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 47.6726 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 233.915 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 25.9050 0.0000 26.0750 0.3300 ;
    END
  END N4END[0]
  PIN S1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.64345 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.757 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.5544 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.6945 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7404 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.584 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 45.6850 0.0000 45.8550 0.3300 ;
    END
  END S1BEG[3]
  PIN S1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08545 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.277 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.916 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 44.7650 0.0000 44.9350 0.3300 ;
    END
  END S1BEG[2]
  PIN S1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.5848 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.8465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.502 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.392 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 43.8450 0.0000 44.0150 0.3300 ;
    END
  END S1BEG[1]
  PIN S1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.778 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.8125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4544 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.154 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 42.9250 0.0000 43.0950 0.3300 ;
    END
  END S1BEG[0]
  PIN S2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.95285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.4392 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.1185 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.656 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 62.7050 0.0000 62.8750 0.3300 ;
    END
  END S2BEG[7]
  PIN S2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.8692 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 34.2685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1688 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.726 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 61.7850 0.0000 61.9550 0.3300 ;
    END
  END S2BEG[6]
  PIN S2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.2324 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.0845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.536 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 60.4050 0.0000 60.5750 0.3300 ;
    END
  END S2BEG[5]
  PIN S2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.7136 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.4905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7092 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.428 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 59.4850 0.0000 59.6550 0.3300 ;
    END
  END S2BEG[4]
  PIN S2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08545 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.277 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.204 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 58.5650 0.0000 58.7350 0.3300 ;
    END
  END S2BEG[3]
  PIN S2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.6776 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.2735 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.298 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 57.6450 0.0000 57.8150 0.3300 ;
    END
  END S2BEG[2]
  PIN S2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7816 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8356 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.06 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 56.2650 0.0000 56.4350 0.3300 ;
    END
  END S2BEG[1]
  PIN S2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.778 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.8125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6452 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.108 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 55.3450 0.0000 55.5150 0.3300 ;
    END
  END S2BEG[0]
  PIN S2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.1644 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.7445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3116 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.44 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 54.4250 0.0000 54.5950 0.3300 ;
    END
  END S2BEGb[7]
  PIN S2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.70125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.825 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.0052 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.9485 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6452 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.108 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 53.0450 0.0000 53.2150 0.3300 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.03 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.0355 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7404 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.584 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 52.1250 0.0000 52.2950 0.3300 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.3372 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.45 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 51.2050 0.0000 51.3750 0.3300 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.16 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.8084 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.9645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1688 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.726 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 50.2850 0.0000 50.4550 0.3300 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.2932 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.3885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.656 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 48.9050 0.0000 49.0750 0.3300 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08545 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.277 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3308 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.961 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.569 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 47.9850 0.0000 48.1550 0.3300 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0355 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.0065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 47.0650 0.0000 47.2350 0.3300 ;
    END
  END S2BEGb[0]
  PIN S4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.24185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.461 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.204 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 79.2650 0.0000 79.4350 0.3300 ;
    END
  END S4BEG[15]
  PIN S4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08545 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.277 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.026 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.012 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 78.3450 0.0000 78.5150 0.3300 ;
    END
  END S4BEG[14]
  PIN S4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.8316 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.922 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 77.4250 0.0000 77.5950 0.3300 ;
    END
  END S4BEG[13]
  PIN S4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08545 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.277 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.312 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.442 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 76.5050 0.0000 76.6750 0.3300 ;
    END
  END S4BEG[12]
  PIN S4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08545 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.277 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.204 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 75.1250 0.0000 75.2950 0.3300 ;
    END
  END S4BEG[11]
  PIN S4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5884 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.298 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 74.2050 0.0000 74.3750 0.3300 ;
    END
  END S4BEG[10]
  PIN S4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.5204 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.5245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0736 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.25 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 73.2850 0.0000 73.4550 0.3300 ;
    END
  END S4BEG[9]
  PIN S4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.24185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.461 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.4008 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.768 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 72.3650 0.0000 72.5350 0.3300 ;
    END
  END S4BEG[8]
  PIN S4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3308 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0436 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.982 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 70.9850 0.0000 71.1550 0.3300 ;
    END
  END S4BEG[7]
  PIN S4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.7512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6391 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.568 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 70.0650 0.0000 70.2350 0.3300 ;
    END
  END S4BEG[6]
  PIN S4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08545 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.277 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6452 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.108 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 69.1450 0.0000 69.3150 0.3300 ;
    END
  END S4BEG[5]
  PIN S4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96985 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.141 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1212 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.488 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 67.7650 0.0000 67.9350 0.3300 ;
    END
  END S4BEG[4]
  PIN S4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96985 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.141 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.134 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.5925 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7404 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.584 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 66.8450 0.0000 67.0150 0.3300 ;
    END
  END S4BEG[3]
  PIN S4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.8764 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.3045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.774 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 65.9250 0.0000 66.0950 0.3300 ;
    END
  END S4BEG[2]
  PIN S4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.5544 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.6945 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3369 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.9148 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.016 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 65.0050 0.0000 65.1750 0.3300 ;
    END
  END S4BEG[1]
  PIN S4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.24185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.461 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2213 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.6995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.735 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.72 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 63.6250 0.0000 63.7950 0.3300 ;
    END
  END S4BEG[0]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.002 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.9325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8352 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.058 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 12.8915 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 60.434 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 28.6450 0.3300 28.8150 ;
    END
  END FrameData[31]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8704 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.024 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.3376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 26.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3116 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.44 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.5557 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 78.3302 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 26.6050 0.3300 26.7750 ;
    END
  END FrameData[30]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.5036 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.4405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6616 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.19 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 13.1657 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 61.3805 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 24.9050 0.3300 25.0750 ;
    END
  END FrameData[29]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.1612 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.7285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1068 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.416 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 16.2915 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 77.0094 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 22.8650 0.3300 23.0350 ;
    END
  END FrameData[28]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.6932 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 28.3885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6448 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.106 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 23.7053 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 114.079 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 21.1650 0.3300 21.3350 ;
    END
  END FrameData[27]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1777 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.6748 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.736 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 59.6657 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 314.374 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 19.1250 0.3300 19.2950 ;
    END
  END FrameData[26]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.89 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.3725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.394 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 7.71541 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 34.1289 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 17.4250 0.3300 17.5950 ;
    END
  END FrameData[25]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2312 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.272 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.4392 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.1185 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8884 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.088 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 8.30283 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 35.5818 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 15.7250 0.3300 15.8950 ;
    END
  END FrameData[24]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.289 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.34 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.4032 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 51.9015 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1404 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.584 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.7972 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 84.5377 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 13.6850 0.3300 13.8550 ;
    END
  END FrameData[23]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2312 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.272 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2496 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.1705 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0751 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.7538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.824 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 72.2783 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 372.925 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 11.9850 0.3300 12.1550 ;
    END
  END FrameData[22]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.3612 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.7285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0048 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.788 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 7.66887 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 33.5786 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 10.2850 0.3300 10.4550 ;
    END
  END FrameData[21]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.3276 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.5605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3759 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.8968 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.92 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 63.172 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 323.327 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 8.2450 0.3300 8.4150 ;
    END
  END FrameData[20]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8632 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2385 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6855 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.2565 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.253 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.816 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 27.7374 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 148.11 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 6.5450 0.3300 6.7150 ;
    END
  END FrameData[19]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2312 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.272 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5884 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.8472 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 30.6877 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 143.833 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 4.5050 0.3300 4.6750 ;
    END
  END FrameData[18]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0842 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.452 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.4556 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.241 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met1  ;
    ANTENNAMAXAREACAR 22.5594 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 109.346 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.181761 LAYER via  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 2.8050 0.3300 2.9750 ;
    END
  END FrameData[17]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3418 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.108 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.6932 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 28.3885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9778 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.653 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 13.7884 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 64.1761 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 0.0000 1.1050 0.3300 1.2750 ;
    END
  END FrameData[16]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3948 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.748 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 24.8349 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 116.022 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 27.6400 0.4850 27.7800 ;
    END
  END FrameData[15]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8344 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.946 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 14.2525 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 66.1352 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 25.9400 0.4850 26.0800 ;
    END
  END FrameData[14]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.839 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.969 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 7.58711 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 32.8082 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 24.2400 0.4850 24.3800 ;
    END
  END FrameData[13]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3131 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4575 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 25.6959 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 124.094 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 22.5400 0.4850 22.6800 ;
    END
  END FrameData[12]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8908 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.228 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 6.95189 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 30.0566 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 20.8400 0.4850 20.9800 ;
    END
  END FrameData[11]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.151 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.411 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 8.58836 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.4969 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 19.1400 0.4850 19.2800 ;
    END
  END FrameData[10]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8169 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9235 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.014 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 75.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.7846 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 31.792 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 60.0129 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 319.075 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 17.4400 0.4850 17.5800 ;
    END
  END FrameData[9]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1589 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6335 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.8798 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.496 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 94.0607 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 491.289 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 15.7400 0.4850 15.8800 ;
    END
  END FrameData[8]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1659 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.37 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.8106 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.264 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 16.5186 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 89.2013 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 14.0400 0.4850 14.1800 ;
    END
  END FrameData[7]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2548 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.93 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 34.3355 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 165.808 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 12.3400 0.4850 12.4800 ;
    END
  END FrameData[6]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9028 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.17 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 15.8978 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 73.6195 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 10.6400 0.4850 10.7800 ;
    END
  END FrameData[5]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1715 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.4658 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.288 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 70.8267 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 374.252 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 8.9400 0.4850 9.0800 ;
    END
  END FrameData[4]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5448 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.616 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 21.6676 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 103.953 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 7.2400 0.4850 7.3800 ;
    END
  END FrameData[3]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4942 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.31 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.438 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.4914 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 36.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 46.8362 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 255.006 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 5.5400 0.4850 5.6800 ;
    END
  END FrameData[2]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5606 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.341 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 20.0349 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 93.5629 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 3.8400 0.4850 3.9800 ;
    END
  END FrameData[1]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2933 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.0208 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.248 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 88.872 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 465.642 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 0.0000 2.1400 0.4850 2.2800 ;
    END
  END FrameData[0]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9338 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.443 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 28.6600 100.2800 28.8000 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6174 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.926 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.413 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.4918 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.76 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 26.6200 100.2800 26.7600 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2156 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.852 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 24.9200 100.2800 25.0600 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5218 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.383 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 22.8800 100.2800 23.0200 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5631 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.5895 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 21.1800 100.2800 21.3200 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0227 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.8875 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 19.1400 100.2800 19.2800 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1295 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.372 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.7284 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 37.296 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 17.4400 100.2800 17.5800 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4148 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.848 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 15.7400 100.2800 15.8800 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.0468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.126 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 13.7000 100.2800 13.8400 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1701 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.24 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.08 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.2564 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.112 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 12.0000 100.2800 12.1400 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7956 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.752 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 10.3000 100.2800 10.4400 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1535 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6595 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 8.2600 100.2800 8.4000 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1504 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.29 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 6.5600 100.2800 6.7000 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0509 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.1465 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 4.5200 100.2800 4.6600 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3836 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.692 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 2.8200 100.2800 2.9600 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0204 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.758 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 99.7950 1.1200 100.2800 1.2600 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.5204 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.5245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7664 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.596 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 27.6250 100.2800 27.7950 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.12 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 50.5225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.216 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.962 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 25.9250 100.2800 26.0950 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7718 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.908 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 11.5368 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 57.6065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.846 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 24.2250 100.2800 24.3950 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.16 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.812 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.9825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0975 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.542 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.024 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.0928 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 27.632 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 22.5250 100.2800 22.6950 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.4184 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 32.0145 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1898 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.831 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 20.8250 100.2800 20.9950 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.6192 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.0185 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1751 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.1318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.84 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 19.1250 100.2800 19.2950 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.139 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.34 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 0.4455 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.2824 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.375 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 17.4250 100.2800 17.5950 ;
    END
  END FrameData_O[9]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2312 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.272 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2972 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4085 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7965 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.8115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.1788 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.424 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 15.7250 100.2800 15.8950 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.07565 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.089 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.4596 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2205 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3821 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7395 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.653 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.616 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.6004 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.28 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 14.0250 100.2800 14.1950 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 0.4455 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.5992 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.922 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 12.3250 100.2800 12.4950 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1156 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.7444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7404 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.584 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 10.6250 100.2800 10.7950 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.204 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 8.8296 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 44.0335 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8828 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.296 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 8.9250 100.2800 9.0950 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0578 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.068 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7144 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.4945 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2471 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9465 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 8.1228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.792 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 7.2250 100.2800 7.3950 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.431 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.86 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 0.4455 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.5404 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.665 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 5.5250 100.2800 5.6950 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2312 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.272 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.5004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.688 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.204 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 3.8250 100.2800 3.9950 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2312 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.272 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.9693 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.6755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.2988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 82.064 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 99.9500 2.1250 100.2800 2.2950 ;
    END
  END FrameData_O[0]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8207 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.8775 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 22.3752 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 106.748 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 97.6800 0.0000 97.8200 0.4850 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9568 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.623 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.335 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.92 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.2868 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 44.5531 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 236.217 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 96.7600 0.0000 96.9000 0.4850 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4917 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.2325 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 19.1965 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 90.8553 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 95.8400 0.0000 95.9800 0.4850 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8417 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.9825 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 20.5877 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 97.8113 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 94.9200 0.0000 95.0600 0.4850 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2371 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9065 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 8.8128 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 47.472 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 106.495 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 557.384 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 94.4600 0.0000 94.6000 0.4850 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.204 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.859 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.16 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.8476 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.128 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 32.0733 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 172.063 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 93.5400 0.0000 93.6800 0.4850 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6163 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.8555 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 18.3601 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 86.673 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 92.6200 0.0000 92.7600 0.4850 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.483 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.254 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.609 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.048 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.1318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.84 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 56.472 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 298.154 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 91.7000 0.0000 91.8400 0.4850 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3452 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.447 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.419 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.2194 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.248 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 52.1336 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 281.569 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 91.2400 0.0000 91.3800 0.4850 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.162 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.649 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.8366 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 42.736 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 128.68 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 685.846 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 90.3200 0.0000 90.4600 0.4850 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8755 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.2695 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 25.9865 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 125.547 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 89.4000 0.0000 89.5400 0.4850 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9683 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7335 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 14.2846 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 67.0377 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 88.4800 0.0000 88.6200 0.4850 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0803 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.2935 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 19.7701 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 94.4654 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 88.0200 0.0000 88.1600 0.4850 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0899 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.2235 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 17.0745 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 80.2453 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 87.1000 0.0000 87.2400 0.4850 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.288 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.8378 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.272 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 23.8708 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 125.138 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 86.1800 0.0000 86.3200 0.4850 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2443 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.8775 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 30.545 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 146.855 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 85.2600 0.0000 85.4000 0.4850 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6827 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3055 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 33.6645 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 163.937 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 84.8000 0.0000 84.9400 0.4850 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9458 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.45 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.3836 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.32 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 67.5248 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 364.654 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 83.8800 0.0000 84.0200 0.4850 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2402 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.922 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.4556 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.704 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 79.0645 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 422.465 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 82.9600 0.0000 83.1000 0.4850 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3538 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.608 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.125 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.8334 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.856 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 77.9324 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 420.61 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 82.5000 0.0000 82.6400 0.4850 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.2335 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.8235 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 97.6800 29.7750 97.8200 30.2600 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0899 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.2235 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 96.7600 29.7750 96.9000 30.2600 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1705 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.5085 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 95.8400 29.7750 95.9800 30.2600 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0324 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.001 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 9.8124 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 53.744 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 94.9200 29.7750 95.0600 30.2600 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9831 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.6895 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 94.4600 29.7750 94.6000 30.2600 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2338 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.008 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.781 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.2324 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 55.984 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 93.5400 29.7750 93.6800 30.2600 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4133 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8405 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 92.6200 29.7750 92.7600 30.2600 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1571 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.5595 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 91.7000 29.7750 91.8400 30.2600 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5874 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.593 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 91.2400 29.7750 91.3800 30.2600 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4091 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8195 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 90.3200 29.7750 90.4600 30.2600 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5875 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8295 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 89.4000 29.7750 89.5400 30.2600 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7327 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.5555 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 88.4800 29.7750 88.6200 30.2600 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4163 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.9735 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 88.0200 29.7750 88.1600 30.2600 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6595 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.9535 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 87.1000 29.7750 87.2400 30.2600 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.224 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.776 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 86.6400 29.7750 86.7800 30.2600 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.344 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.559 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.025 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.8476 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.128 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 85.7200 29.7750 85.8600 30.2600 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9061 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.3045 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 84.8000 29.7750 84.9400 30.2600 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5995 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.7715 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 83.8800 29.7750 84.0200 30.2600 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3447 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4975 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 82.9600 29.7750 83.1000 30.2600 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9681 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.6145 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 82.5000 29.7750 82.6400 30.2600 ;
    END
  END FrameStrobe_O[0]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 5.5600 4.0700 94.7200 6.0700 ;
        RECT 5.5600 23.0000 94.7200 25.0000 ;
        RECT 92.7200 15.0600 94.7200 15.5400 ;
        RECT 5.5600 15.0600 7.5600 15.5400 ;
        RECT 5.5600 9.6200 7.5600 10.1000 ;
        RECT 92.7200 9.6200 94.7200 10.1000 ;
        RECT 5.5600 20.5000 7.5600 20.9800 ;
        RECT 92.7200 20.5000 94.7200 20.9800 ;
      LAYER met4 ;
        RECT 5.5600 4.0700 7.5600 25.0000 ;
        RECT 92.7200 4.0700 94.7200 25.0000 ;
    END
# end of P/G power stripe data as pin

  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 2.5600 1.0700 97.7200 3.0700 ;
        RECT 2.5600 26.0000 97.7200 28.0000 ;
        RECT 2.5600 12.3400 4.5600 12.8200 ;
        RECT 2.5600 6.9000 4.5600 7.3800 ;
        RECT 95.7200 12.3400 97.7200 12.8200 ;
        RECT 95.7200 6.9000 97.7200 7.3800 ;
        RECT 2.5600 17.7800 4.5600 18.2600 ;
        RECT 95.7200 17.7800 97.7200 18.2600 ;
      LAYER met4 ;
        RECT 2.5600 1.0700 4.5600 28.0000 ;
        RECT 95.7200 1.0700 97.7200 28.0000 ;
    END
# end of P/G power stripe data as pin

  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.0000 28.9850 100.2800 30.2600 ;
      RECT 0.5000 28.4750 100.2800 28.9850 ;
      RECT 0.0000 27.9650 100.2800 28.4750 ;
      RECT 0.0000 27.4550 99.7800 27.9650 ;
      RECT 0.0000 26.9450 100.2800 27.4550 ;
      RECT 0.5000 26.4350 100.2800 26.9450 ;
      RECT 0.0000 26.2650 100.2800 26.4350 ;
      RECT 0.0000 25.7550 99.7800 26.2650 ;
      RECT 0.0000 25.2450 100.2800 25.7550 ;
      RECT 0.5000 24.7350 100.2800 25.2450 ;
      RECT 0.0000 24.5650 100.2800 24.7350 ;
      RECT 0.0000 24.0550 99.7800 24.5650 ;
      RECT 0.0000 23.2050 100.2800 24.0550 ;
      RECT 0.5000 22.8650 100.2800 23.2050 ;
      RECT 0.5000 22.6950 99.7800 22.8650 ;
      RECT 0.0000 22.3550 99.7800 22.6950 ;
      RECT 0.0000 21.5050 100.2800 22.3550 ;
      RECT 0.5000 21.1650 100.2800 21.5050 ;
      RECT 0.5000 20.9950 99.7800 21.1650 ;
      RECT 0.0000 20.6550 99.7800 20.9950 ;
      RECT 0.0000 19.4650 100.2800 20.6550 ;
      RECT 0.5000 18.9550 99.7800 19.4650 ;
      RECT 0.0000 17.7650 100.2800 18.9550 ;
      RECT 0.5000 17.2550 99.7800 17.7650 ;
      RECT 0.0000 16.0650 100.2800 17.2550 ;
      RECT 0.5000 15.5550 99.7800 16.0650 ;
      RECT 0.0000 14.3650 100.2800 15.5550 ;
      RECT 0.0000 14.0250 99.7800 14.3650 ;
      RECT 0.5000 13.8550 99.7800 14.0250 ;
      RECT 0.5000 13.5150 100.2800 13.8550 ;
      RECT 0.0000 12.6650 100.2800 13.5150 ;
      RECT 0.0000 12.3250 99.7800 12.6650 ;
      RECT 0.5000 12.1550 99.7800 12.3250 ;
      RECT 0.5000 11.8150 100.2800 12.1550 ;
      RECT 0.0000 10.9650 100.2800 11.8150 ;
      RECT 0.0000 10.6250 99.7800 10.9650 ;
      RECT 0.5000 10.4550 99.7800 10.6250 ;
      RECT 0.5000 10.1150 100.2800 10.4550 ;
      RECT 0.0000 9.2650 100.2800 10.1150 ;
      RECT 0.0000 8.7550 99.7800 9.2650 ;
      RECT 0.0000 8.5850 100.2800 8.7550 ;
      RECT 0.5000 8.0750 100.2800 8.5850 ;
      RECT 0.0000 7.5650 100.2800 8.0750 ;
      RECT 0.0000 7.0550 99.7800 7.5650 ;
      RECT 0.0000 6.8850 100.2800 7.0550 ;
      RECT 0.5000 6.3750 100.2800 6.8850 ;
      RECT 0.0000 5.8650 100.2800 6.3750 ;
      RECT 0.0000 5.3550 99.7800 5.8650 ;
      RECT 0.0000 4.8450 100.2800 5.3550 ;
      RECT 0.5000 4.3350 100.2800 4.8450 ;
      RECT 0.0000 4.1650 100.2800 4.3350 ;
      RECT 0.0000 3.6550 99.7800 4.1650 ;
      RECT 0.0000 3.1450 100.2800 3.6550 ;
      RECT 0.5000 2.6350 100.2800 3.1450 ;
      RECT 0.0000 2.4650 100.2800 2.6350 ;
      RECT 0.0000 1.9550 99.7800 2.4650 ;
      RECT 0.0000 1.4450 100.2800 1.9550 ;
      RECT 0.5000 0.9350 100.2800 1.4450 ;
      RECT 0.0000 0.5000 100.2800 0.9350 ;
      RECT 79.6050 0.0000 100.2800 0.5000 ;
      RECT 78.6850 0.0000 79.0950 0.5000 ;
      RECT 77.7650 0.0000 78.1750 0.5000 ;
      RECT 76.8450 0.0000 77.2550 0.5000 ;
      RECT 75.4650 0.0000 76.3350 0.5000 ;
      RECT 74.5450 0.0000 74.9550 0.5000 ;
      RECT 73.6250 0.0000 74.0350 0.5000 ;
      RECT 72.7050 0.0000 73.1150 0.5000 ;
      RECT 71.3250 0.0000 72.1950 0.5000 ;
      RECT 70.4050 0.0000 70.8150 0.5000 ;
      RECT 69.4850 0.0000 69.8950 0.5000 ;
      RECT 68.1050 0.0000 68.9750 0.5000 ;
      RECT 67.1850 0.0000 67.5950 0.5000 ;
      RECT 66.2650 0.0000 66.6750 0.5000 ;
      RECT 65.3450 0.0000 65.7550 0.5000 ;
      RECT 63.9650 0.0000 64.8350 0.5000 ;
      RECT 63.0450 0.0000 63.4550 0.5000 ;
      RECT 62.1250 0.0000 62.5350 0.5000 ;
      RECT 60.7450 0.0000 61.6150 0.5000 ;
      RECT 59.8250 0.0000 60.2350 0.5000 ;
      RECT 58.9050 0.0000 59.3150 0.5000 ;
      RECT 57.9850 0.0000 58.3950 0.5000 ;
      RECT 56.6050 0.0000 57.4750 0.5000 ;
      RECT 55.6850 0.0000 56.0950 0.5000 ;
      RECT 54.7650 0.0000 55.1750 0.5000 ;
      RECT 53.3850 0.0000 54.2550 0.5000 ;
      RECT 52.4650 0.0000 52.8750 0.5000 ;
      RECT 51.5450 0.0000 51.9550 0.5000 ;
      RECT 50.6250 0.0000 51.0350 0.5000 ;
      RECT 49.2450 0.0000 50.1150 0.5000 ;
      RECT 48.3250 0.0000 48.7350 0.5000 ;
      RECT 47.4050 0.0000 47.8150 0.5000 ;
      RECT 46.0250 0.0000 46.8950 0.5000 ;
      RECT 45.1050 0.0000 45.5150 0.5000 ;
      RECT 44.1850 0.0000 44.5950 0.5000 ;
      RECT 43.2650 0.0000 43.6750 0.5000 ;
      RECT 41.8850 0.0000 42.7550 0.5000 ;
      RECT 40.9650 0.0000 41.3750 0.5000 ;
      RECT 40.0450 0.0000 40.4550 0.5000 ;
      RECT 39.1250 0.0000 39.5350 0.5000 ;
      RECT 37.7450 0.0000 38.6150 0.5000 ;
      RECT 36.8250 0.0000 37.2350 0.5000 ;
      RECT 35.9050 0.0000 36.3150 0.5000 ;
      RECT 34.5250 0.0000 35.3950 0.5000 ;
      RECT 33.6050 0.0000 34.0150 0.5000 ;
      RECT 32.6850 0.0000 33.0950 0.5000 ;
      RECT 31.7650 0.0000 32.1750 0.5000 ;
      RECT 30.3850 0.0000 31.2550 0.5000 ;
      RECT 29.4650 0.0000 29.8750 0.5000 ;
      RECT 28.5450 0.0000 28.9550 0.5000 ;
      RECT 27.1650 0.0000 28.0350 0.5000 ;
      RECT 26.2450 0.0000 26.6550 0.5000 ;
      RECT 25.3250 0.0000 25.7350 0.5000 ;
      RECT 24.4050 0.0000 24.8150 0.5000 ;
      RECT 23.0250 0.0000 23.8950 0.5000 ;
      RECT 22.1050 0.0000 22.5150 0.5000 ;
      RECT 21.1850 0.0000 21.5950 0.5000 ;
      RECT 19.8050 0.0000 20.6750 0.5000 ;
      RECT 18.8850 0.0000 19.2950 0.5000 ;
      RECT 17.9650 0.0000 18.3750 0.5000 ;
      RECT 17.0450 0.0000 17.4550 0.5000 ;
      RECT 15.6650 0.0000 16.5350 0.5000 ;
      RECT 14.7450 0.0000 15.1550 0.5000 ;
      RECT 13.8250 0.0000 14.2350 0.5000 ;
      RECT 12.4450 0.0000 13.3150 0.5000 ;
      RECT 11.5250 0.0000 11.9350 0.5000 ;
      RECT 10.6050 0.0000 11.0150 0.5000 ;
      RECT 9.6850 0.0000 10.0950 0.5000 ;
      RECT 8.3050 0.0000 9.1750 0.5000 ;
      RECT 7.3850 0.0000 7.7950 0.5000 ;
      RECT 6.4650 0.0000 6.8750 0.5000 ;
      RECT 5.5450 0.0000 5.9550 0.5000 ;
      RECT 0.0000 0.0000 5.0350 0.5000 ;
    LAYER met1 ;
      RECT 0.0000 0.0000 100.2800 30.2600 ;
    LAYER met2 ;
      RECT 97.9600 29.6350 100.2800 30.2600 ;
      RECT 97.0400 29.6350 97.5400 30.2600 ;
      RECT 96.1200 29.6350 96.6200 30.2600 ;
      RECT 95.2000 29.6350 95.7000 30.2600 ;
      RECT 94.7400 29.6350 94.7800 30.2600 ;
      RECT 93.8200 29.6350 94.3200 30.2600 ;
      RECT 92.9000 29.6350 93.4000 30.2600 ;
      RECT 91.9800 29.6350 92.4800 30.2600 ;
      RECT 91.5200 29.6350 91.5600 30.2600 ;
      RECT 90.6000 29.6350 91.1000 30.2600 ;
      RECT 89.6800 29.6350 90.1800 30.2600 ;
      RECT 88.7600 29.6350 89.2600 30.2600 ;
      RECT 88.3000 29.6350 88.3400 30.2600 ;
      RECT 87.3800 29.6350 87.8800 30.2600 ;
      RECT 86.9200 29.6350 86.9600 30.2600 ;
      RECT 86.0000 29.6350 86.5000 30.2600 ;
      RECT 85.0800 29.6350 85.5800 30.2600 ;
      RECT 84.1600 29.6350 84.6600 30.2600 ;
      RECT 83.2400 29.6350 83.7400 30.2600 ;
      RECT 82.7800 29.6350 82.8200 30.2600 ;
      RECT 0.0000 29.6350 82.3600 30.2600 ;
      RECT 0.0000 28.9400 100.2800 29.6350 ;
      RECT 0.0000 28.5200 99.6550 28.9400 ;
      RECT 0.0000 27.9200 100.2800 28.5200 ;
      RECT 0.6250 27.5000 100.2800 27.9200 ;
      RECT 0.0000 26.9000 100.2800 27.5000 ;
      RECT 0.0000 26.4800 99.6550 26.9000 ;
      RECT 0.0000 26.2200 100.2800 26.4800 ;
      RECT 0.6250 25.8000 100.2800 26.2200 ;
      RECT 0.0000 25.2000 100.2800 25.8000 ;
      RECT 0.0000 24.7800 99.6550 25.2000 ;
      RECT 0.0000 24.5200 100.2800 24.7800 ;
      RECT 0.6250 24.1000 100.2800 24.5200 ;
      RECT 0.0000 23.1600 100.2800 24.1000 ;
      RECT 0.0000 22.8200 99.6550 23.1600 ;
      RECT 0.6250 22.7400 99.6550 22.8200 ;
      RECT 0.6250 22.4000 100.2800 22.7400 ;
      RECT 0.0000 21.4600 100.2800 22.4000 ;
      RECT 0.0000 21.1200 99.6550 21.4600 ;
      RECT 0.6250 21.0400 99.6550 21.1200 ;
      RECT 0.6250 20.7000 100.2800 21.0400 ;
      RECT 0.0000 19.4200 100.2800 20.7000 ;
      RECT 0.6250 19.0000 99.6550 19.4200 ;
      RECT 0.0000 17.7200 100.2800 19.0000 ;
      RECT 0.6250 17.3000 99.6550 17.7200 ;
      RECT 0.0000 16.0200 100.2800 17.3000 ;
      RECT 0.6250 15.6000 99.6550 16.0200 ;
      RECT 0.0000 14.3200 100.2800 15.6000 ;
      RECT 0.6250 13.9800 100.2800 14.3200 ;
      RECT 0.6250 13.9000 99.6550 13.9800 ;
      RECT 0.0000 13.5600 99.6550 13.9000 ;
      RECT 0.0000 12.6200 100.2800 13.5600 ;
      RECT 0.6250 12.2800 100.2800 12.6200 ;
      RECT 0.6250 12.2000 99.6550 12.2800 ;
      RECT 0.0000 11.8600 99.6550 12.2000 ;
      RECT 0.0000 10.9200 100.2800 11.8600 ;
      RECT 0.6250 10.5800 100.2800 10.9200 ;
      RECT 0.6250 10.5000 99.6550 10.5800 ;
      RECT 0.0000 10.1600 99.6550 10.5000 ;
      RECT 0.0000 9.2200 100.2800 10.1600 ;
      RECT 0.6250 8.8000 100.2800 9.2200 ;
      RECT 0.0000 8.5400 100.2800 8.8000 ;
      RECT 0.0000 8.1200 99.6550 8.5400 ;
      RECT 0.0000 7.5200 100.2800 8.1200 ;
      RECT 0.6250 7.1000 100.2800 7.5200 ;
      RECT 0.0000 6.8400 100.2800 7.1000 ;
      RECT 0.0000 6.4200 99.6550 6.8400 ;
      RECT 0.0000 5.8200 100.2800 6.4200 ;
      RECT 0.6250 5.4000 100.2800 5.8200 ;
      RECT 0.0000 4.8000 100.2800 5.4000 ;
      RECT 0.0000 4.3800 99.6550 4.8000 ;
      RECT 0.0000 4.1200 100.2800 4.3800 ;
      RECT 0.6250 3.7000 100.2800 4.1200 ;
      RECT 0.0000 3.1000 100.2800 3.7000 ;
      RECT 0.0000 2.6800 99.6550 3.1000 ;
      RECT 0.0000 2.4200 100.2800 2.6800 ;
      RECT 0.6250 2.0000 100.2800 2.4200 ;
      RECT 0.0000 1.4000 100.2800 2.0000 ;
      RECT 0.0000 0.9800 99.6550 1.4000 ;
      RECT 0.0000 0.6250 100.2800 0.9800 ;
      RECT 97.9600 0.0000 100.2800 0.6250 ;
      RECT 97.0400 0.0000 97.5400 0.6250 ;
      RECT 96.1200 0.0000 96.6200 0.6250 ;
      RECT 95.2000 0.0000 95.7000 0.6250 ;
      RECT 94.7400 0.0000 94.7800 0.6250 ;
      RECT 93.8200 0.0000 94.3200 0.6250 ;
      RECT 92.9000 0.0000 93.4000 0.6250 ;
      RECT 91.9800 0.0000 92.4800 0.6250 ;
      RECT 91.5200 0.0000 91.5600 0.6250 ;
      RECT 90.6000 0.0000 91.1000 0.6250 ;
      RECT 89.6800 0.0000 90.1800 0.6250 ;
      RECT 88.7600 0.0000 89.2600 0.6250 ;
      RECT 88.3000 0.0000 88.3400 0.6250 ;
      RECT 87.3800 0.0000 87.8800 0.6250 ;
      RECT 86.4600 0.0000 86.9600 0.6250 ;
      RECT 85.5400 0.0000 86.0400 0.6250 ;
      RECT 85.0800 0.0000 85.1200 0.6250 ;
      RECT 84.1600 0.0000 84.6600 0.6250 ;
      RECT 83.2400 0.0000 83.7400 0.6250 ;
      RECT 82.7800 0.0000 82.8200 0.6250 ;
      RECT 0.0000 0.0000 82.3600 0.6250 ;
    LAYER met3 ;
      RECT 0.0000 28.3000 100.2800 30.2600 ;
      RECT 98.0200 25.7000 100.2800 28.3000 ;
      RECT 0.0000 25.7000 2.2600 28.3000 ;
      RECT 0.0000 25.3000 100.2800 25.7000 ;
      RECT 95.0200 22.7000 100.2800 25.3000 ;
      RECT 0.0000 22.7000 5.2600 25.3000 ;
      RECT 0.0000 21.2800 100.2800 22.7000 ;
      RECT 95.0200 20.2000 100.2800 21.2800 ;
      RECT 7.8600 20.2000 92.4200 21.2800 ;
      RECT 0.0000 20.2000 5.2600 21.2800 ;
      RECT 0.0000 18.5600 100.2800 20.2000 ;
      RECT 98.0200 17.4800 100.2800 18.5600 ;
      RECT 4.8600 17.4800 95.4200 18.5600 ;
      RECT 0.0000 17.4800 2.2600 18.5600 ;
      RECT 0.0000 15.8400 100.2800 17.4800 ;
      RECT 95.0200 14.7600 100.2800 15.8400 ;
      RECT 7.8600 14.7600 92.4200 15.8400 ;
      RECT 0.0000 14.7600 5.2600 15.8400 ;
      RECT 0.0000 13.1200 100.2800 14.7600 ;
      RECT 98.0200 12.0400 100.2800 13.1200 ;
      RECT 4.8600 12.0400 95.4200 13.1200 ;
      RECT 0.0000 12.0400 2.2600 13.1200 ;
      RECT 0.0000 10.4000 100.2800 12.0400 ;
      RECT 95.0200 9.3200 100.2800 10.4000 ;
      RECT 7.8600 9.3200 92.4200 10.4000 ;
      RECT 0.0000 9.3200 5.2600 10.4000 ;
      RECT 0.0000 7.6800 100.2800 9.3200 ;
      RECT 98.0200 6.6000 100.2800 7.6800 ;
      RECT 4.8600 6.6000 95.4200 7.6800 ;
      RECT 0.0000 6.6000 2.2600 7.6800 ;
      RECT 0.0000 6.3700 100.2800 6.6000 ;
      RECT 95.0200 3.7700 100.2800 6.3700 ;
      RECT 0.0000 3.7700 5.2600 6.3700 ;
      RECT 0.0000 3.3700 100.2800 3.7700 ;
      RECT 98.0200 0.7700 100.2800 3.3700 ;
      RECT 0.0000 0.7700 2.2600 3.3700 ;
      RECT 0.0000 0.0000 100.2800 0.7700 ;
    LAYER met4 ;
      RECT 0.0000 28.3000 100.2800 30.2600 ;
      RECT 4.8600 25.3000 95.4200 28.3000 ;
      RECT 95.0200 3.7700 95.4200 25.3000 ;
      RECT 7.8600 3.7700 92.4200 25.3000 ;
      RECT 4.8600 3.7700 5.2600 25.3000 ;
      RECT 98.0200 0.7700 100.2800 28.3000 ;
      RECT 4.8600 0.7700 95.4200 3.7700 ;
      RECT 0.0000 0.7700 2.2600 28.3000 ;
      RECT 0.0000 0.0000 100.2800 0.7700 ;
  END
END N_term_RAM_IO

END LIBRARY
