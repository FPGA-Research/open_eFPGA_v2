magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -66 377 3426 897
<< pwell >>
rect 2641 283 2907 317
rect 545 217 1976 283
rect 2641 217 3356 283
rect 11 43 3356 217
rect -26 -43 3386 43
<< locali >>
rect 119 235 185 344
rect 596 301 733 424
rect 699 126 733 301
rect 770 162 833 421
rect 1433 365 1703 399
rect 1669 259 1703 365
rect 1291 225 1703 259
rect 1291 126 1325 225
rect 699 92 1325 126
rect 1669 87 1703 225
rect 2826 356 2876 751
rect 2302 226 2368 270
rect 2181 192 2368 226
rect 2809 299 2876 356
rect 2181 87 2215 192
rect 1669 53 2215 87
rect 2809 133 2885 299
rect 3268 103 3338 751
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3360 831
rect 119 735 297 741
rect 153 701 191 735
rect 225 701 263 735
rect 33 489 83 691
rect 119 525 297 701
rect 333 727 641 761
rect 333 489 367 727
rect 33 455 367 489
rect 33 199 83 455
rect 301 380 367 455
rect 403 310 455 691
rect 505 494 571 684
rect 607 564 641 727
rect 677 735 711 741
rect 677 600 711 701
rect 747 720 1113 754
rect 747 564 781 720
rect 817 600 903 684
rect 973 600 1043 684
rect 607 530 781 564
rect 869 494 903 600
rect 505 460 903 494
rect 403 199 437 310
rect 33 99 99 199
rect 135 113 325 199
rect 135 79 141 113
rect 175 79 213 113
rect 247 79 285 113
rect 319 79 325 113
rect 361 99 437 199
rect 473 113 663 265
rect 135 73 325 79
rect 473 79 479 113
rect 513 79 551 113
rect 585 79 623 113
rect 657 79 663 113
rect 869 265 903 460
rect 939 356 973 564
rect 1009 474 1043 600
rect 1079 609 1113 720
rect 1149 735 1337 741
rect 1149 701 1154 735
rect 1188 701 1226 735
rect 1260 701 1298 735
rect 1332 701 1337 735
rect 1149 645 1337 701
rect 1373 727 1547 761
rect 1373 609 1407 727
rect 1079 575 1407 609
rect 1079 510 1130 575
rect 1443 539 1477 691
rect 1513 574 1547 727
rect 1583 735 1773 741
rect 1583 701 1589 735
rect 1623 701 1661 735
rect 1695 701 1733 735
rect 1767 701 1773 735
rect 1583 610 1773 701
rect 2118 735 2308 741
rect 2118 701 2124 735
rect 2158 701 2196 735
rect 2230 701 2268 735
rect 2302 701 2308 735
rect 1513 540 1875 574
rect 1221 505 1477 539
rect 1221 474 1255 505
rect 1009 440 1255 474
rect 1739 469 1805 504
rect 1119 356 1185 404
rect 939 301 1185 356
rect 1221 329 1255 440
rect 1291 435 1805 469
rect 1291 365 1357 435
rect 1221 295 1633 329
rect 1221 265 1255 295
rect 869 165 931 265
rect 1054 231 1255 265
rect 1054 165 1120 231
rect 1443 113 1633 189
rect 473 73 663 79
rect 1443 79 1449 113
rect 1483 79 1521 113
rect 1555 79 1593 113
rect 1627 79 1633 113
rect 1443 73 1633 79
rect 1739 123 1805 435
rect 1841 280 1875 540
rect 1911 488 1961 670
rect 1911 454 2082 488
rect 2118 470 2308 701
rect 2612 735 2790 751
rect 2646 701 2684 735
rect 2718 701 2756 735
rect 2393 504 2459 554
rect 2393 470 2576 504
rect 2048 434 2082 454
rect 1945 316 2012 418
rect 2048 400 2506 434
rect 1841 246 2075 280
rect 2018 214 2075 246
rect 1916 157 1982 199
rect 2111 157 2145 400
rect 2440 376 2506 400
rect 2186 340 2252 364
rect 2542 340 2576 470
rect 2612 435 2790 701
rect 3035 735 3225 751
rect 3035 701 3041 735
rect 3075 701 3113 735
rect 3147 701 3185 735
rect 3219 701 3225 735
rect 2186 306 2576 340
rect 2186 262 2252 306
rect 1916 123 2145 157
rect 2542 195 2576 306
rect 2933 367 2999 601
rect 3035 435 3225 701
rect 2933 301 3232 367
rect 2251 113 2441 156
rect 2251 79 2257 113
rect 2291 79 2329 113
rect 2363 79 2401 113
rect 2435 79 2441 113
rect 2542 103 2615 195
rect 2651 113 2769 299
rect 2933 165 3003 301
rect 2251 73 2441 79
rect 2651 79 2657 113
rect 2691 79 2729 113
rect 2763 79 2769 113
rect 2651 73 2769 79
rect 3039 113 3229 265
rect 3039 79 3045 113
rect 3079 79 3117 113
rect 3151 79 3189 113
rect 3223 79 3229 113
rect 3039 73 3229 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3360 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 1663 797 1697 831
rect 1759 797 1793 831
rect 1855 797 1889 831
rect 1951 797 1985 831
rect 2047 797 2081 831
rect 2143 797 2177 831
rect 2239 797 2273 831
rect 2335 797 2369 831
rect 2431 797 2465 831
rect 2527 797 2561 831
rect 2623 797 2657 831
rect 2719 797 2753 831
rect 2815 797 2849 831
rect 2911 797 2945 831
rect 3007 797 3041 831
rect 3103 797 3137 831
rect 3199 797 3233 831
rect 3295 797 3329 831
rect 119 701 153 735
rect 191 701 225 735
rect 263 701 297 735
rect 677 701 711 735
rect 141 79 175 113
rect 213 79 247 113
rect 285 79 319 113
rect 479 79 513 113
rect 551 79 585 113
rect 623 79 657 113
rect 1154 701 1188 735
rect 1226 701 1260 735
rect 1298 701 1332 735
rect 1589 701 1623 735
rect 1661 701 1695 735
rect 1733 701 1767 735
rect 2124 701 2158 735
rect 2196 701 2230 735
rect 2268 701 2302 735
rect 1449 79 1483 113
rect 1521 79 1555 113
rect 1593 79 1627 113
rect 2612 701 2646 735
rect 2684 701 2718 735
rect 2756 701 2790 735
rect 3041 701 3075 735
rect 3113 701 3147 735
rect 3185 701 3219 735
rect 2257 79 2291 113
rect 2329 79 2363 113
rect 2401 79 2435 113
rect 2657 79 2691 113
rect 2729 79 2763 113
rect 3045 79 3079 113
rect 3117 79 3151 113
rect 3189 79 3223 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
<< metal1 >>
rect 0 831 3360 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1663 831
rect 1697 797 1759 831
rect 1793 797 1855 831
rect 1889 797 1951 831
rect 1985 797 2047 831
rect 2081 797 2143 831
rect 2177 797 2239 831
rect 2273 797 2335 831
rect 2369 797 2431 831
rect 2465 797 2527 831
rect 2561 797 2623 831
rect 2657 797 2719 831
rect 2753 797 2815 831
rect 2849 797 2911 831
rect 2945 797 3007 831
rect 3041 797 3103 831
rect 3137 797 3199 831
rect 3233 797 3295 831
rect 3329 797 3360 831
rect 0 791 3360 797
rect 0 735 3360 763
rect 0 701 119 735
rect 153 701 191 735
rect 225 701 263 735
rect 297 701 677 735
rect 711 701 1154 735
rect 1188 701 1226 735
rect 1260 701 1298 735
rect 1332 701 1589 735
rect 1623 701 1661 735
rect 1695 701 1733 735
rect 1767 701 2124 735
rect 2158 701 2196 735
rect 2230 701 2268 735
rect 2302 701 2612 735
rect 2646 701 2684 735
rect 2718 701 2756 735
rect 2790 701 3041 735
rect 3075 701 3113 735
rect 3147 701 3185 735
rect 3219 701 3360 735
rect 0 689 3360 701
rect 0 113 3360 125
rect 0 79 141 113
rect 175 79 213 113
rect 247 79 285 113
rect 319 79 479 113
rect 513 79 551 113
rect 585 79 623 113
rect 657 79 1449 113
rect 1483 79 1521 113
rect 1555 79 1593 113
rect 1627 79 2257 113
rect 2291 79 2329 113
rect 2363 79 2401 113
rect 2435 79 2657 113
rect 2691 79 2729 113
rect 2763 79 3045 113
rect 3079 79 3117 113
rect 3151 79 3189 113
rect 3223 79 3360 113
rect 0 51 3360 79
rect 0 17 3360 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3360 17
rect 0 -23 3360 -17
<< obsm1 >>
rect 403 347 461 356
rect 979 347 1037 356
rect 1939 347 1997 356
rect 403 319 1997 347
rect 403 310 461 319
rect 979 310 1037 319
rect 1939 310 1997 319
<< labels >>
rlabel locali s 119 235 185 344 6 CLK
port 1 nsew clock input
rlabel locali s 770 162 833 421 6 D
port 2 nsew signal input
rlabel locali s 1669 53 2215 87 6 RESET_B
port 3 nsew signal input
rlabel locali s 2181 87 2215 192 6 RESET_B
port 3 nsew signal input
rlabel locali s 2181 192 2368 226 6 RESET_B
port 3 nsew signal input
rlabel locali s 1669 87 1703 225 6 RESET_B
port 3 nsew signal input
rlabel locali s 699 92 1325 126 6 RESET_B
port 3 nsew signal input
rlabel locali s 1291 126 1325 225 6 RESET_B
port 3 nsew signal input
rlabel locali s 2302 226 2368 270 6 RESET_B
port 3 nsew signal input
rlabel locali s 1291 225 1703 259 6 RESET_B
port 3 nsew signal input
rlabel locali s 1669 259 1703 365 6 RESET_B
port 3 nsew signal input
rlabel locali s 699 126 733 301 6 RESET_B
port 3 nsew signal input
rlabel locali s 1433 365 1703 399 6 RESET_B
port 3 nsew signal input
rlabel locali s 596 301 733 424 6 RESET_B
port 3 nsew signal input
rlabel metal1 s 0 51 3360 125 6 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 -23 3360 23 8 VNB
port 5 nsew ground bidirectional
rlabel pwell s -26 -43 3386 43 8 VNB
port 5 nsew ground bidirectional
rlabel pwell s 11 43 3356 217 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 2641 217 3356 283 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 545 217 1976 283 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 2641 283 2907 317 6 VNB
port 5 nsew ground bidirectional
rlabel metal1 s 0 791 3360 837 6 VPB
port 6 nsew power bidirectional
rlabel nwell s -66 377 3426 897 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 689 3360 763 6 VPWR
port 7 nsew power bidirectional
rlabel locali s 3268 103 3338 751 6 Q
port 8 nsew signal output
rlabel locali s 2809 133 2885 299 6 Q_N
port 9 nsew signal output
rlabel locali s 2809 299 2876 356 6 Q_N
port 9 nsew signal output
rlabel locali s 2826 356 2876 751 6 Q_N
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 3360 814
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1031444
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 1000180
<< end >>
