magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -36 679 4724 1471
<< pwell >>
rect 4552 25 4654 159
<< psubdiff >>
rect 4578 109 4628 133
rect 4578 75 4586 109
rect 4620 75 4628 109
rect 4578 51 4628 75
<< nsubdiff >>
rect 4578 1339 4628 1363
rect 4578 1305 4586 1339
rect 4620 1305 4628 1339
rect 4578 1281 4628 1305
<< psubdiffcont >>
rect 4586 75 4620 109
<< nsubdiffcont >>
rect 4586 1305 4620 1339
<< poly >>
rect 114 740 144 907
rect 48 724 144 740
rect 48 690 64 724
rect 98 690 144 724
rect 48 674 144 690
rect 114 507 144 674
<< polycont >>
rect 64 690 98 724
<< locali >>
rect 0 1397 4688 1431
rect 62 1130 96 1397
rect 274 1130 308 1397
rect 490 1130 524 1397
rect 706 1130 740 1397
rect 922 1130 956 1397
rect 1138 1130 1172 1397
rect 1354 1130 1388 1397
rect 1570 1130 1604 1397
rect 1786 1130 1820 1397
rect 2002 1130 2036 1397
rect 2218 1130 2252 1397
rect 2434 1130 2468 1397
rect 2650 1130 2684 1397
rect 2866 1130 2900 1397
rect 3082 1130 3116 1397
rect 3298 1130 3332 1397
rect 3514 1130 3548 1397
rect 3730 1130 3764 1397
rect 3946 1130 3980 1397
rect 4162 1130 4196 1397
rect 4378 1130 4412 1397
rect 4586 1339 4620 1397
rect 4586 1289 4620 1305
rect 64 724 98 740
rect 64 674 98 690
rect 2324 724 2358 1096
rect 2324 690 2375 724
rect 2324 318 2358 690
rect 62 17 96 218
rect 274 17 308 218
rect 490 17 524 218
rect 706 17 740 218
rect 922 17 956 218
rect 1138 17 1172 218
rect 1354 17 1388 218
rect 1570 17 1604 218
rect 1786 17 1820 218
rect 2002 17 2036 218
rect 2218 17 2252 218
rect 2434 17 2468 218
rect 2650 17 2684 218
rect 2866 17 2900 218
rect 3082 17 3116 218
rect 3298 17 3332 218
rect 3514 17 3548 218
rect 3730 17 3764 218
rect 3946 17 3980 218
rect 4162 17 4196 218
rect 4378 17 4412 218
rect 4586 109 4620 125
rect 4586 17 4620 75
rect 0 -17 4688 17
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_16  sky130_sram_2kbyte_1rw1r_32x512_8_contact_16_0
timestamp 1707688321
transform 1 0 48 0 1 674
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_28  sky130_sram_2kbyte_1rw1r_32x512_8_contact_28_0
timestamp 1707688321
transform 1 0 4578 0 1 1281
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_29  sky130_sram_2kbyte_1rw1r_32x512_8_contact_29_0
timestamp 1707688321
transform 1 0 4578 0 1 51
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_nmos_m41_w2_000_sli_dli_da_p  sky130_sram_2kbyte_1rw1r_32x512_8_nmos_m41_w2_000_sli_dli_da_p_0
timestamp 1707688321
transform 1 0 54 0 1 51
box -26 -26 4496 456
use sky130_sram_2kbyte_1rw1r_32x512_8_pmos_m41_w2_000_sli_dli_da_p  sky130_sram_2kbyte_1rw1r_32x512_8_pmos_m41_w2_000_sli_dli_da_p_0
timestamp 1707688321
transform 1 0 54 0 1 963
box -59 -56 4529 454
<< labels >>
rlabel locali s 81 707 81 707 4 A
rlabel locali s 2358 707 2358 707 4 Z
rlabel locali s 2344 0 2344 0 4 gnd
rlabel locali s 2344 1414 2344 1414 4 vdd
<< properties >>
string FIXED_BBOX 0 0 4688 1414
string GDS_END 357800
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_START 353370
<< end >>
