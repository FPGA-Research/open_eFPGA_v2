magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -38 261 1878 582
<< pwell >>
rect 1 21 1822 157
rect 29 -17 63 21
<< scnmos >>
rect 80 47 110 131
rect 166 47 196 131
rect 252 47 282 131
rect 338 47 368 131
rect 424 47 454 131
rect 510 47 540 131
rect 596 47 626 131
rect 682 47 712 131
rect 768 47 798 131
rect 854 47 884 131
rect 940 47 970 131
rect 1026 47 1056 131
rect 1111 47 1141 131
rect 1197 47 1227 131
rect 1283 47 1313 131
rect 1369 47 1399 131
rect 1455 47 1485 131
rect 1541 47 1571 131
rect 1627 47 1657 131
rect 1713 47 1743 131
<< scpmoshvt >>
rect 80 297 110 497
rect 166 297 196 497
rect 252 297 282 497
rect 338 297 368 497
rect 424 297 454 497
rect 510 297 540 497
rect 596 297 626 497
rect 682 297 712 497
rect 768 297 798 497
rect 854 297 884 497
rect 940 297 970 497
rect 1026 297 1056 497
rect 1111 297 1141 497
rect 1197 297 1227 497
rect 1283 297 1313 497
rect 1369 297 1399 497
rect 1455 297 1485 497
rect 1541 297 1571 497
rect 1627 297 1657 497
rect 1713 297 1743 497
<< ndiff >>
rect 27 93 80 131
rect 27 59 35 93
rect 69 59 80 93
rect 27 47 80 59
rect 110 106 166 131
rect 110 72 121 106
rect 155 72 166 106
rect 110 47 166 72
rect 196 106 252 131
rect 196 72 207 106
rect 241 72 252 106
rect 196 47 252 72
rect 282 106 338 131
rect 282 72 293 106
rect 327 72 338 106
rect 282 47 338 72
rect 368 106 424 131
rect 368 72 379 106
rect 413 72 424 106
rect 368 47 424 72
rect 454 106 510 131
rect 454 72 465 106
rect 499 72 510 106
rect 454 47 510 72
rect 540 97 596 131
rect 540 63 551 97
rect 585 63 596 97
rect 540 47 596 63
rect 626 106 682 131
rect 626 72 637 106
rect 671 72 682 106
rect 626 47 682 72
rect 712 97 768 131
rect 712 63 723 97
rect 757 63 768 97
rect 712 47 768 63
rect 798 106 854 131
rect 798 72 809 106
rect 843 72 854 106
rect 798 47 854 72
rect 884 97 940 131
rect 884 63 895 97
rect 929 63 940 97
rect 884 47 940 63
rect 970 106 1026 131
rect 970 72 981 106
rect 1015 72 1026 106
rect 970 47 1026 72
rect 1056 97 1111 131
rect 1056 63 1067 97
rect 1101 63 1111 97
rect 1056 47 1111 63
rect 1141 106 1197 131
rect 1141 72 1152 106
rect 1186 72 1197 106
rect 1141 47 1197 72
rect 1227 97 1283 131
rect 1227 63 1238 97
rect 1272 63 1283 97
rect 1227 47 1283 63
rect 1313 106 1369 131
rect 1313 72 1324 106
rect 1358 72 1369 106
rect 1313 47 1369 72
rect 1399 97 1455 131
rect 1399 63 1410 97
rect 1444 63 1455 97
rect 1399 47 1455 63
rect 1485 106 1541 131
rect 1485 72 1496 106
rect 1530 72 1541 106
rect 1485 47 1541 72
rect 1571 97 1627 131
rect 1571 63 1582 97
rect 1616 63 1627 97
rect 1571 47 1627 63
rect 1657 106 1713 131
rect 1657 72 1668 106
rect 1702 72 1713 106
rect 1657 47 1713 72
rect 1743 97 1796 131
rect 1743 63 1754 97
rect 1788 63 1796 97
rect 1743 47 1796 63
<< pdiff >>
rect 27 485 80 497
rect 27 451 35 485
rect 69 451 80 485
rect 27 417 80 451
rect 27 383 35 417
rect 69 383 80 417
rect 27 349 80 383
rect 27 315 35 349
rect 69 315 80 349
rect 27 297 80 315
rect 110 476 166 497
rect 110 442 121 476
rect 155 442 166 476
rect 110 408 166 442
rect 110 374 121 408
rect 155 374 166 408
rect 110 340 166 374
rect 110 306 121 340
rect 155 306 166 340
rect 110 297 166 306
rect 196 485 252 497
rect 196 451 207 485
rect 241 451 252 485
rect 196 417 252 451
rect 196 383 207 417
rect 241 383 252 417
rect 196 349 252 383
rect 196 315 207 349
rect 241 315 252 349
rect 196 297 252 315
rect 282 476 338 497
rect 282 442 293 476
rect 327 442 338 476
rect 282 408 338 442
rect 282 374 293 408
rect 327 374 338 408
rect 282 340 338 374
rect 282 306 293 340
rect 327 306 338 340
rect 282 297 338 306
rect 368 485 424 497
rect 368 451 379 485
rect 413 451 424 485
rect 368 417 424 451
rect 368 383 379 417
rect 413 383 424 417
rect 368 349 424 383
rect 368 315 379 349
rect 413 315 424 349
rect 368 297 424 315
rect 454 476 510 497
rect 454 442 465 476
rect 499 442 510 476
rect 454 349 510 442
rect 454 315 465 349
rect 499 315 510 349
rect 454 297 510 315
rect 540 461 596 497
rect 540 427 551 461
rect 585 427 596 461
rect 540 297 596 427
rect 626 476 682 497
rect 626 442 637 476
rect 671 442 682 476
rect 626 349 682 442
rect 626 315 637 349
rect 671 315 682 349
rect 626 297 682 315
rect 712 461 768 497
rect 712 427 723 461
rect 757 427 768 461
rect 712 297 768 427
rect 798 476 854 497
rect 798 442 809 476
rect 843 442 854 476
rect 798 349 854 442
rect 798 315 809 349
rect 843 315 854 349
rect 798 297 854 315
rect 884 461 940 497
rect 884 427 895 461
rect 929 427 940 461
rect 884 297 940 427
rect 970 476 1026 497
rect 970 442 981 476
rect 1015 442 1026 476
rect 970 349 1026 442
rect 970 315 981 349
rect 1015 315 1026 349
rect 970 297 1026 315
rect 1056 461 1111 497
rect 1056 427 1067 461
rect 1101 427 1111 461
rect 1056 297 1111 427
rect 1141 476 1197 497
rect 1141 442 1152 476
rect 1186 442 1197 476
rect 1141 349 1197 442
rect 1141 315 1152 349
rect 1186 315 1197 349
rect 1141 297 1197 315
rect 1227 461 1283 497
rect 1227 427 1238 461
rect 1272 427 1283 461
rect 1227 297 1283 427
rect 1313 476 1369 497
rect 1313 442 1324 476
rect 1358 442 1369 476
rect 1313 349 1369 442
rect 1313 315 1324 349
rect 1358 315 1369 349
rect 1313 297 1369 315
rect 1399 461 1455 497
rect 1399 427 1410 461
rect 1444 427 1455 461
rect 1399 297 1455 427
rect 1485 476 1541 497
rect 1485 442 1496 476
rect 1530 442 1541 476
rect 1485 349 1541 442
rect 1485 315 1496 349
rect 1530 315 1541 349
rect 1485 297 1541 315
rect 1571 461 1627 497
rect 1571 427 1582 461
rect 1616 427 1627 461
rect 1571 297 1627 427
rect 1657 476 1713 497
rect 1657 442 1668 476
rect 1702 442 1713 476
rect 1657 349 1713 442
rect 1657 315 1668 349
rect 1702 315 1713 349
rect 1657 297 1713 315
rect 1743 461 1796 497
rect 1743 427 1754 461
rect 1788 427 1796 461
rect 1743 297 1796 427
<< ndiffc >>
rect 35 59 69 93
rect 121 72 155 106
rect 207 72 241 106
rect 293 72 327 106
rect 379 72 413 106
rect 465 72 499 106
rect 551 63 585 97
rect 637 72 671 106
rect 723 63 757 97
rect 809 72 843 106
rect 895 63 929 97
rect 981 72 1015 106
rect 1067 63 1101 97
rect 1152 72 1186 106
rect 1238 63 1272 97
rect 1324 72 1358 106
rect 1410 63 1444 97
rect 1496 72 1530 106
rect 1582 63 1616 97
rect 1668 72 1702 106
rect 1754 63 1788 97
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 121 442 155 476
rect 121 374 155 408
rect 121 306 155 340
rect 207 451 241 485
rect 207 383 241 417
rect 207 315 241 349
rect 293 442 327 476
rect 293 374 327 408
rect 293 306 327 340
rect 379 451 413 485
rect 379 383 413 417
rect 379 315 413 349
rect 465 442 499 476
rect 465 315 499 349
rect 551 427 585 461
rect 637 442 671 476
rect 637 315 671 349
rect 723 427 757 461
rect 809 442 843 476
rect 809 315 843 349
rect 895 427 929 461
rect 981 442 1015 476
rect 981 315 1015 349
rect 1067 427 1101 461
rect 1152 442 1186 476
rect 1152 315 1186 349
rect 1238 427 1272 461
rect 1324 442 1358 476
rect 1324 315 1358 349
rect 1410 427 1444 461
rect 1496 442 1530 476
rect 1496 315 1530 349
rect 1582 427 1616 461
rect 1668 442 1702 476
rect 1668 315 1702 349
rect 1754 427 1788 461
<< poly >>
rect 80 497 110 523
rect 166 497 196 523
rect 252 497 282 523
rect 338 497 368 523
rect 424 497 454 523
rect 510 497 540 523
rect 596 497 626 523
rect 682 497 712 523
rect 768 497 798 523
rect 854 497 884 523
rect 940 497 970 523
rect 1026 497 1056 523
rect 1111 497 1141 523
rect 1197 497 1227 523
rect 1283 497 1313 523
rect 1369 497 1399 523
rect 1455 497 1485 523
rect 1541 497 1571 523
rect 1627 497 1657 523
rect 1713 497 1743 523
rect 80 282 110 297
rect 166 282 196 297
rect 252 282 282 297
rect 338 282 368 297
rect 21 249 368 282
rect 21 215 37 249
rect 71 215 368 249
rect 21 180 368 215
rect 80 131 110 180
rect 166 131 196 180
rect 252 131 282 180
rect 338 131 368 180
rect 424 265 454 297
rect 510 265 540 297
rect 596 265 626 297
rect 682 265 712 297
rect 768 265 798 297
rect 854 265 884 297
rect 940 265 970 297
rect 1026 265 1056 297
rect 1111 265 1141 297
rect 1197 265 1227 297
rect 1283 265 1313 297
rect 1369 265 1399 297
rect 1455 265 1485 297
rect 1541 265 1571 297
rect 1627 265 1657 297
rect 1713 265 1743 297
rect 424 249 1743 265
rect 424 215 464 249
rect 498 215 532 249
rect 566 215 600 249
rect 634 215 668 249
rect 702 215 736 249
rect 770 215 804 249
rect 838 215 872 249
rect 906 215 940 249
rect 974 215 1008 249
rect 1042 215 1076 249
rect 1110 215 1144 249
rect 1178 215 1212 249
rect 1246 215 1280 249
rect 1314 215 1348 249
rect 1382 215 1416 249
rect 1450 215 1484 249
rect 1518 215 1743 249
rect 424 190 1743 215
rect 424 131 454 190
rect 510 131 540 190
rect 596 131 626 190
rect 682 131 712 190
rect 768 131 798 190
rect 854 131 884 190
rect 940 131 970 190
rect 1026 131 1056 190
rect 1111 131 1141 190
rect 1197 131 1227 190
rect 1283 131 1313 190
rect 1369 131 1399 190
rect 1455 131 1485 190
rect 1541 131 1571 190
rect 1627 131 1657 190
rect 1713 131 1743 190
rect 80 21 110 47
rect 166 21 196 47
rect 252 21 282 47
rect 338 21 368 47
rect 424 21 454 47
rect 510 21 540 47
rect 596 21 626 47
rect 682 21 712 47
rect 768 21 798 47
rect 854 21 884 47
rect 940 21 970 47
rect 1026 21 1056 47
rect 1111 21 1141 47
rect 1197 21 1227 47
rect 1283 21 1313 47
rect 1369 21 1399 47
rect 1455 21 1485 47
rect 1541 21 1571 47
rect 1627 21 1657 47
rect 1713 21 1743 47
<< polycont >>
rect 37 215 71 249
rect 464 215 498 249
rect 532 215 566 249
rect 600 215 634 249
rect 668 215 702 249
rect 736 215 770 249
rect 804 215 838 249
rect 872 215 906 249
rect 940 215 974 249
rect 1008 215 1042 249
rect 1076 215 1110 249
rect 1144 215 1178 249
rect 1212 215 1246 249
rect 1280 215 1314 249
rect 1348 215 1382 249
rect 1416 215 1450 249
rect 1484 215 1518 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 19 485 85 493
rect 19 425 35 485
rect 69 425 85 485
rect 19 417 85 425
rect 19 383 35 417
rect 69 383 85 417
rect 19 349 85 383
rect 19 315 35 349
rect 69 315 85 349
rect 19 299 85 315
rect 119 476 157 493
rect 119 442 121 476
rect 155 442 157 476
rect 119 408 157 442
rect 119 374 121 408
rect 155 374 157 408
rect 119 340 157 374
rect 119 306 121 340
rect 155 306 157 340
rect 119 265 157 306
rect 191 485 257 493
rect 191 425 207 485
rect 241 425 257 485
rect 191 417 257 425
rect 191 383 207 417
rect 241 383 257 417
rect 191 349 257 383
rect 191 315 207 349
rect 241 315 257 349
rect 191 299 257 315
rect 291 476 329 492
rect 291 442 293 476
rect 327 442 329 476
rect 291 408 329 442
rect 291 374 293 408
rect 327 374 329 408
rect 291 340 329 374
rect 291 306 293 340
rect 327 306 329 340
rect 291 265 329 306
rect 363 485 429 493
rect 363 459 379 485
rect 363 425 378 459
rect 413 451 429 485
rect 412 425 429 451
rect 363 417 429 425
rect 363 383 379 417
rect 413 383 429 417
rect 363 349 429 383
rect 363 315 379 349
rect 413 315 429 349
rect 363 299 429 315
rect 463 476 508 492
rect 463 442 465 476
rect 499 442 508 476
rect 463 349 508 442
rect 542 461 594 493
rect 542 459 551 461
rect 542 425 548 459
rect 585 427 594 461
rect 582 425 594 427
rect 542 381 594 425
rect 628 476 680 492
rect 628 442 637 476
rect 671 442 680 476
rect 463 315 465 349
rect 499 347 508 349
rect 628 349 680 442
rect 714 461 766 493
rect 714 427 723 461
rect 757 459 766 461
rect 714 425 724 427
rect 758 425 766 459
rect 714 381 766 425
rect 800 476 852 492
rect 800 442 809 476
rect 843 442 852 476
rect 628 347 637 349
rect 499 315 637 347
rect 671 347 680 349
rect 800 349 852 442
rect 886 461 938 493
rect 886 427 895 461
rect 929 459 938 461
rect 886 425 896 427
rect 930 425 938 459
rect 886 381 938 425
rect 972 476 1024 492
rect 972 442 981 476
rect 1015 442 1024 476
rect 800 347 809 349
rect 671 315 809 347
rect 843 347 852 349
rect 972 349 1024 442
rect 1058 461 1107 493
rect 1058 425 1067 461
rect 1101 425 1107 461
rect 1058 381 1107 425
rect 1141 476 1193 492
rect 1141 442 1152 476
rect 1186 442 1193 476
rect 972 347 981 349
rect 843 315 981 347
rect 1015 347 1024 349
rect 1141 349 1193 442
rect 1230 461 1279 493
rect 1230 427 1238 461
rect 1272 459 1279 461
rect 1230 425 1239 427
rect 1273 425 1279 459
rect 1230 381 1279 425
rect 1313 476 1365 492
rect 1313 442 1324 476
rect 1358 442 1365 476
rect 1141 347 1152 349
rect 1015 315 1152 347
rect 1186 347 1193 349
rect 1313 349 1365 442
rect 1402 461 1451 493
rect 1402 425 1410 461
rect 1444 425 1451 461
rect 1402 381 1451 425
rect 1485 476 1537 492
rect 1485 442 1496 476
rect 1530 442 1537 476
rect 1313 347 1324 349
rect 1186 315 1324 347
rect 1358 347 1365 349
rect 1485 349 1537 442
rect 1574 461 1625 493
rect 1574 459 1582 461
rect 1574 425 1580 459
rect 1616 427 1625 461
rect 1614 425 1625 427
rect 1574 381 1625 425
rect 1659 476 1717 492
rect 1659 442 1668 476
rect 1702 442 1717 476
rect 1485 347 1496 349
rect 1358 315 1496 347
rect 1530 344 1537 349
rect 1659 349 1717 442
rect 1751 461 1805 493
rect 1751 427 1754 461
rect 1788 459 1805 461
rect 1751 425 1756 427
rect 1790 425 1805 459
rect 1751 378 1805 425
rect 1659 344 1668 349
rect 1530 315 1668 344
rect 1702 344 1717 349
rect 1702 315 1805 344
rect 463 299 1805 315
rect 17 249 80 265
rect 17 215 37 249
rect 71 215 80 249
rect 17 153 80 215
rect 119 249 1538 265
rect 119 215 464 249
rect 498 215 532 249
rect 566 215 600 249
rect 634 215 668 249
rect 702 215 736 249
rect 770 215 804 249
rect 838 215 872 249
rect 906 215 940 249
rect 974 215 1008 249
rect 1042 215 1076 249
rect 1110 215 1144 249
rect 1178 215 1212 249
rect 1246 215 1280 249
rect 1314 215 1348 249
rect 1382 215 1416 249
rect 1450 215 1484 249
rect 1518 215 1538 249
rect 17 93 78 119
rect 17 59 35 93
rect 69 59 78 93
rect 17 17 78 59
rect 119 106 164 215
rect 119 72 121 106
rect 155 72 164 106
rect 119 53 164 72
rect 198 106 250 122
rect 198 72 207 106
rect 241 72 250 106
rect 198 17 250 72
rect 286 106 336 215
rect 1572 181 1805 299
rect 456 147 1805 181
rect 286 72 293 106
rect 327 72 336 106
rect 286 53 336 72
rect 370 106 422 129
rect 370 72 379 106
rect 413 72 422 106
rect 370 17 422 72
rect 456 106 508 147
rect 456 72 465 106
rect 499 72 508 106
rect 456 56 508 72
rect 542 97 594 113
rect 542 63 551 97
rect 585 63 594 97
rect 542 17 594 63
rect 628 106 680 147
rect 628 72 637 106
rect 671 72 680 106
rect 628 56 680 72
rect 714 97 766 113
rect 714 63 723 97
rect 757 63 766 97
rect 714 17 766 63
rect 800 106 852 147
rect 800 72 809 106
rect 843 72 852 106
rect 800 56 852 72
rect 886 97 935 113
rect 886 63 895 97
rect 929 63 935 97
rect 886 17 935 63
rect 969 106 1024 147
rect 969 72 981 106
rect 1015 72 1024 106
rect 969 56 1024 72
rect 1058 97 1107 113
rect 1058 63 1067 97
rect 1101 63 1107 97
rect 1058 17 1107 63
rect 1141 106 1193 147
rect 1141 72 1152 106
rect 1186 72 1193 106
rect 1141 56 1193 72
rect 1229 97 1279 113
rect 1229 63 1238 97
rect 1272 63 1279 97
rect 1229 17 1279 63
rect 1313 106 1365 147
rect 1313 72 1324 106
rect 1358 72 1365 106
rect 1313 56 1365 72
rect 1401 97 1451 113
rect 1401 63 1410 97
rect 1444 63 1451 97
rect 1401 17 1451 63
rect 1485 106 1537 147
rect 1485 72 1496 106
rect 1530 72 1537 106
rect 1485 56 1537 72
rect 1573 97 1625 113
rect 1573 63 1582 97
rect 1616 63 1625 97
rect 1573 17 1625 63
rect 1659 106 1711 147
rect 1659 72 1668 106
rect 1702 72 1711 106
rect 1659 56 1711 72
rect 1745 97 1805 113
rect 1745 63 1754 97
rect 1788 63 1805 97
rect 1745 17 1805 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 35 451 69 459
rect 35 425 69 451
rect 207 451 241 459
rect 207 425 241 451
rect 378 451 379 459
rect 379 451 412 459
rect 378 425 412 451
rect 548 427 551 459
rect 551 427 582 459
rect 548 425 582 427
rect 724 427 757 459
rect 757 427 758 459
rect 724 425 758 427
rect 896 427 929 459
rect 929 427 930 459
rect 896 425 930 427
rect 1067 427 1101 459
rect 1067 425 1101 427
rect 1239 427 1272 459
rect 1272 427 1273 459
rect 1239 425 1273 427
rect 1410 427 1444 459
rect 1410 425 1444 427
rect 1580 427 1582 459
rect 1582 427 1614 459
rect 1580 425 1614 427
rect 1756 427 1788 459
rect 1788 427 1790 459
rect 1756 425 1790 427
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
<< metal1 >>
rect 0 561 1840 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 0 496 1840 527
rect 14 459 1826 468
rect 14 428 35 459
rect 23 425 35 428
rect 69 428 207 459
rect 69 425 81 428
rect 23 416 81 425
rect 195 425 207 428
rect 241 428 378 459
rect 241 425 253 428
rect 195 416 253 425
rect 366 425 378 428
rect 412 428 548 459
rect 412 425 424 428
rect 366 416 424 425
rect 536 425 548 428
rect 582 428 724 459
rect 582 425 594 428
rect 536 416 594 425
rect 712 425 724 428
rect 758 428 896 459
rect 758 425 770 428
rect 712 416 770 425
rect 884 425 896 428
rect 930 428 1067 459
rect 930 425 942 428
rect 884 416 942 425
rect 1055 425 1067 428
rect 1101 428 1239 459
rect 1101 425 1113 428
rect 1055 416 1113 425
rect 1227 425 1239 428
rect 1273 428 1410 459
rect 1273 425 1285 428
rect 1227 416 1285 425
rect 1398 425 1410 428
rect 1444 428 1580 459
rect 1444 425 1456 428
rect 1398 416 1456 425
rect 1568 425 1580 428
rect 1614 428 1756 459
rect 1614 425 1626 428
rect 1568 416 1626 425
rect 1744 425 1756 428
rect 1790 428 1826 459
rect 1790 425 1802 428
rect 1744 416 1802 425
rect 0 17 1840 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
rect 0 -48 1840 -17
<< labels >>
flabel locali s 1593 289 1627 323 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 1685 289 1719 323 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 1685 221 1719 255 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 1593 221 1627 255 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 1593 153 1627 187 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 1685 153 1719 187 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 29 153 63 187 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel metal1 s 28 428 77 468 0 FreeSans 200 0 0 0 KAPWR
port 2 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 lpflow_clkbufkapwr_16
rlabel locali s 191 299 257 493 1 KAPWR
port 2 nsew power bidirectional abutment
rlabel locali s 363 299 429 493 1 KAPWR
port 2 nsew power bidirectional abutment
rlabel locali s 542 381 594 493 1 KAPWR
port 2 nsew power bidirectional abutment
rlabel locali s 714 381 766 493 1 KAPWR
port 2 nsew power bidirectional abutment
rlabel locali s 886 381 938 493 1 KAPWR
port 2 nsew power bidirectional abutment
rlabel locali s 1058 381 1107 493 1 KAPWR
port 2 nsew power bidirectional abutment
rlabel locali s 1230 381 1279 493 1 KAPWR
port 2 nsew power bidirectional abutment
rlabel locali s 1402 381 1451 493 1 KAPWR
port 2 nsew power bidirectional abutment
rlabel locali s 1574 381 1625 493 1 KAPWR
port 2 nsew power bidirectional abutment
rlabel locali s 1751 378 1805 493 1 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 1744 416 1802 428 1 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 1568 416 1626 428 1 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 1398 416 1456 428 1 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 1227 416 1285 428 1 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 1055 416 1113 428 1 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 884 416 942 428 1 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 712 416 770 428 1 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 536 416 594 428 1 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 366 416 424 428 1 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 195 416 253 428 1 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 23 416 81 428 1 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 14 428 1826 468 1 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 0 -48 1840 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1840 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1840 544
string GDS_END 2276556
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2261950
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
