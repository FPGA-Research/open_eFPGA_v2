magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect 7977 5506 8787 6258
<< pwell >>
rect 12973 3313 13195 4714
rect 12743 2714 13195 3313
rect 12973 2652 13195 2714
rect 15803 3583 16071 4714
rect 15803 3180 16174 3583
rect 15803 2661 16071 3180
rect 15123 1841 16025 1991
<< pdiff >>
rect 8919 4392 8957 4630
rect 10176 4392 10209 4630
<< psubdiff >>
rect 12999 4664 13169 4688
rect 13033 4630 13067 4664
rect 13101 4630 13135 4664
rect 12999 4595 13169 4630
rect 13033 4561 13067 4595
rect 13101 4561 13135 4595
rect 12999 4526 13169 4561
rect 13033 4492 13067 4526
rect 13101 4492 13135 4526
rect 12999 4457 13169 4492
rect 13033 4423 13067 4457
rect 13101 4423 13135 4457
rect 12999 4388 13169 4423
rect 13033 4354 13067 4388
rect 13101 4354 13135 4388
rect 12999 4319 13169 4354
rect 13033 4285 13067 4319
rect 13101 4285 13135 4319
rect 12999 4250 13169 4285
rect 13033 4216 13067 4250
rect 13101 4216 13135 4250
rect 12999 4181 13169 4216
rect 13033 4147 13067 4181
rect 13101 4147 13135 4181
rect 12999 4112 13169 4147
rect 13033 4078 13067 4112
rect 13101 4078 13135 4112
rect 12999 4043 13169 4078
rect 13033 4009 13067 4043
rect 13101 4009 13135 4043
rect 12999 3974 13169 4009
rect 13033 3940 13067 3974
rect 13101 3940 13135 3974
rect 12999 3905 13169 3940
rect 13033 3871 13067 3905
rect 13101 3871 13135 3905
rect 12999 3836 13169 3871
rect 13033 3802 13067 3836
rect 13101 3802 13135 3836
rect 12999 3767 13169 3802
rect 13033 3733 13067 3767
rect 13101 3733 13135 3767
rect 12999 3698 13169 3733
rect 13033 3664 13067 3698
rect 13101 3664 13135 3698
rect 12999 3629 13169 3664
rect 13033 3595 13067 3629
rect 13101 3595 13135 3629
rect 12999 3560 13169 3595
rect 13033 3526 13067 3560
rect 13101 3526 13135 3560
rect 12999 3491 13169 3526
rect 13033 3457 13067 3491
rect 13101 3457 13135 3491
rect 12999 3422 13169 3457
rect 13033 3388 13067 3422
rect 13101 3388 13135 3422
rect 12999 3353 13169 3388
rect 13033 3319 13067 3353
rect 13101 3319 13135 3353
rect 12999 3287 13169 3319
rect 12769 3284 13169 3287
rect 12769 3263 12999 3284
rect 12769 3229 12842 3263
rect 12876 3229 12910 3263
rect 12944 3250 12999 3263
rect 13033 3250 13067 3284
rect 13101 3250 13135 3284
rect 12944 3229 13169 3250
rect 12769 3215 13169 3229
rect 12769 3185 12999 3215
rect 12769 3151 12842 3185
rect 12876 3151 12910 3185
rect 12944 3181 12999 3185
rect 13033 3181 13067 3215
rect 13101 3181 13135 3215
rect 12944 3151 13169 3181
rect 12769 3146 13169 3151
rect 12769 3112 12999 3146
rect 13033 3112 13067 3146
rect 13101 3112 13135 3146
rect 12769 3107 13169 3112
rect 12769 3073 12842 3107
rect 12876 3073 12910 3107
rect 12944 3077 13169 3107
rect 12944 3073 12999 3077
rect 12769 3043 12999 3073
rect 13033 3043 13067 3077
rect 13101 3043 13135 3077
rect 12769 3029 13169 3043
rect 12769 2995 12842 3029
rect 12876 2995 12910 3029
rect 12944 3008 13169 3029
rect 12944 2995 12999 3008
rect 12769 2952 12999 2995
rect 12769 2918 12842 2952
rect 12876 2918 12910 2952
rect 12944 2918 12999 2952
rect 12769 2875 12999 2918
rect 12769 2841 12842 2875
rect 12876 2841 12910 2875
rect 12944 2841 12999 2875
rect 12769 2798 12999 2841
rect 12769 2764 12842 2798
rect 12876 2764 12910 2798
rect 12944 2764 12999 2798
rect 12769 2740 12999 2764
rect 12999 2678 13169 2702
rect 15829 4664 16045 4688
rect 15829 4630 15852 4664
rect 15886 4630 15920 4664
rect 15954 4630 15988 4664
rect 16022 4630 16045 4664
rect 15829 4595 16045 4630
rect 15829 4561 15852 4595
rect 15886 4561 15920 4595
rect 15954 4561 15988 4595
rect 16022 4561 16045 4595
rect 15829 4526 16045 4561
rect 15829 4492 15852 4526
rect 15886 4492 15920 4526
rect 15954 4492 15988 4526
rect 16022 4492 16045 4526
rect 15829 4457 16045 4492
rect 15829 4423 15852 4457
rect 15886 4423 15920 4457
rect 15954 4423 15988 4457
rect 16022 4423 16045 4457
rect 15829 4388 16045 4423
rect 15829 4354 15852 4388
rect 15886 4354 15920 4388
rect 15954 4354 15988 4388
rect 16022 4354 16045 4388
rect 15829 4319 16045 4354
rect 15829 4285 15852 4319
rect 15886 4285 15920 4319
rect 15954 4285 15988 4319
rect 16022 4285 16045 4319
rect 15829 4250 16045 4285
rect 15829 4216 15852 4250
rect 15886 4216 15920 4250
rect 15954 4216 15988 4250
rect 16022 4216 16045 4250
rect 15829 4181 16045 4216
rect 15829 4147 15852 4181
rect 15886 4147 15920 4181
rect 15954 4147 15988 4181
rect 16022 4147 16045 4181
rect 15829 4112 16045 4147
rect 15829 4078 15852 4112
rect 15886 4078 15920 4112
rect 15954 4078 15988 4112
rect 16022 4078 16045 4112
rect 15829 4043 16045 4078
rect 15829 4009 15852 4043
rect 15886 4009 15920 4043
rect 15954 4009 15988 4043
rect 16022 4009 16045 4043
rect 15829 3974 16045 4009
rect 15829 3940 15852 3974
rect 15886 3940 15920 3974
rect 15954 3940 15988 3974
rect 16022 3940 16045 3974
rect 15829 3905 16045 3940
rect 15829 3871 15852 3905
rect 15886 3871 15920 3905
rect 15954 3871 15988 3905
rect 16022 3871 16045 3905
rect 15829 3836 16045 3871
rect 15829 3802 15852 3836
rect 15886 3802 15920 3836
rect 15954 3802 15988 3836
rect 16022 3802 16045 3836
rect 15829 3767 16045 3802
rect 15829 3733 15852 3767
rect 15886 3733 15920 3767
rect 15954 3733 15988 3767
rect 16022 3733 16045 3767
rect 15829 3698 16045 3733
rect 15829 3664 15852 3698
rect 15886 3664 15920 3698
rect 15954 3664 15988 3698
rect 16022 3664 16045 3698
rect 15829 3629 16045 3664
rect 15829 2711 15852 3629
rect 16022 3557 16045 3629
rect 16022 3206 16148 3557
rect 16022 2711 16045 3206
rect 15829 2687 16045 2711
rect 15149 1901 15999 1965
rect 15149 1867 15173 1901
rect 15207 1867 15243 1901
rect 15277 1867 15313 1901
rect 15347 1867 15383 1901
rect 15417 1867 15453 1901
rect 15487 1867 15523 1901
rect 15557 1867 15593 1901
rect 15627 1867 15663 1901
rect 15697 1867 15733 1901
rect 15767 1867 15803 1901
rect 15837 1867 15872 1901
rect 15906 1867 15941 1901
rect 15975 1867 15999 1901
<< psubdiffcont >>
rect 12999 4630 13033 4664
rect 13067 4630 13101 4664
rect 13135 4630 13169 4664
rect 12999 4561 13033 4595
rect 13067 4561 13101 4595
rect 13135 4561 13169 4595
rect 12999 4492 13033 4526
rect 13067 4492 13101 4526
rect 13135 4492 13169 4526
rect 12999 4423 13033 4457
rect 13067 4423 13101 4457
rect 13135 4423 13169 4457
rect 12999 4354 13033 4388
rect 13067 4354 13101 4388
rect 13135 4354 13169 4388
rect 12999 4285 13033 4319
rect 13067 4285 13101 4319
rect 13135 4285 13169 4319
rect 12999 4216 13033 4250
rect 13067 4216 13101 4250
rect 13135 4216 13169 4250
rect 12999 4147 13033 4181
rect 13067 4147 13101 4181
rect 13135 4147 13169 4181
rect 12999 4078 13033 4112
rect 13067 4078 13101 4112
rect 13135 4078 13169 4112
rect 12999 4009 13033 4043
rect 13067 4009 13101 4043
rect 13135 4009 13169 4043
rect 12999 3940 13033 3974
rect 13067 3940 13101 3974
rect 13135 3940 13169 3974
rect 12999 3871 13033 3905
rect 13067 3871 13101 3905
rect 13135 3871 13169 3905
rect 12999 3802 13033 3836
rect 13067 3802 13101 3836
rect 13135 3802 13169 3836
rect 12999 3733 13033 3767
rect 13067 3733 13101 3767
rect 13135 3733 13169 3767
rect 12999 3664 13033 3698
rect 13067 3664 13101 3698
rect 13135 3664 13169 3698
rect 12999 3595 13033 3629
rect 13067 3595 13101 3629
rect 13135 3595 13169 3629
rect 12999 3526 13033 3560
rect 13067 3526 13101 3560
rect 13135 3526 13169 3560
rect 12999 3457 13033 3491
rect 13067 3457 13101 3491
rect 13135 3457 13169 3491
rect 12999 3388 13033 3422
rect 13067 3388 13101 3422
rect 13135 3388 13169 3422
rect 12999 3319 13033 3353
rect 13067 3319 13101 3353
rect 13135 3319 13169 3353
rect 12842 3229 12876 3263
rect 12910 3229 12944 3263
rect 12999 3250 13033 3284
rect 13067 3250 13101 3284
rect 13135 3250 13169 3284
rect 12842 3151 12876 3185
rect 12910 3151 12944 3185
rect 12999 3181 13033 3215
rect 13067 3181 13101 3215
rect 13135 3181 13169 3215
rect 12999 3112 13033 3146
rect 13067 3112 13101 3146
rect 13135 3112 13169 3146
rect 12842 3073 12876 3107
rect 12910 3073 12944 3107
rect 12999 3043 13033 3077
rect 13067 3043 13101 3077
rect 13135 3043 13169 3077
rect 12842 2995 12876 3029
rect 12910 2995 12944 3029
rect 12842 2918 12876 2952
rect 12910 2918 12944 2952
rect 12842 2841 12876 2875
rect 12910 2841 12944 2875
rect 12842 2764 12876 2798
rect 12910 2764 12944 2798
rect 12999 2702 13169 3008
rect 15852 4630 15886 4664
rect 15920 4630 15954 4664
rect 15988 4630 16022 4664
rect 15852 4561 15886 4595
rect 15920 4561 15954 4595
rect 15988 4561 16022 4595
rect 15852 4492 15886 4526
rect 15920 4492 15954 4526
rect 15988 4492 16022 4526
rect 15852 4423 15886 4457
rect 15920 4423 15954 4457
rect 15988 4423 16022 4457
rect 15852 4354 15886 4388
rect 15920 4354 15954 4388
rect 15988 4354 16022 4388
rect 15852 4285 15886 4319
rect 15920 4285 15954 4319
rect 15988 4285 16022 4319
rect 15852 4216 15886 4250
rect 15920 4216 15954 4250
rect 15988 4216 16022 4250
rect 15852 4147 15886 4181
rect 15920 4147 15954 4181
rect 15988 4147 16022 4181
rect 15852 4078 15886 4112
rect 15920 4078 15954 4112
rect 15988 4078 16022 4112
rect 15852 4009 15886 4043
rect 15920 4009 15954 4043
rect 15988 4009 16022 4043
rect 15852 3940 15886 3974
rect 15920 3940 15954 3974
rect 15988 3940 16022 3974
rect 15852 3871 15886 3905
rect 15920 3871 15954 3905
rect 15988 3871 16022 3905
rect 15852 3802 15886 3836
rect 15920 3802 15954 3836
rect 15988 3802 16022 3836
rect 15852 3733 15886 3767
rect 15920 3733 15954 3767
rect 15988 3733 16022 3767
rect 15852 3664 15886 3698
rect 15920 3664 15954 3698
rect 15988 3664 16022 3698
rect 15852 2711 16022 3629
rect 15173 1867 15207 1901
rect 15243 1867 15277 1901
rect 15313 1867 15347 1901
rect 15383 1867 15417 1901
rect 15453 1867 15487 1901
rect 15523 1867 15557 1901
rect 15593 1867 15627 1901
rect 15663 1867 15697 1901
rect 15733 1867 15767 1901
rect 15803 1867 15837 1901
rect 15872 1867 15906 1901
rect 15941 1867 15975 1901
<< locali >>
rect 7572 8847 7610 8881
rect 8183 8807 8385 8842
rect 8183 8773 8199 8807
rect 8233 8773 8271 8807
rect 8305 8773 8343 8807
rect 8377 8773 8385 8807
rect 13147 6070 13185 6104
rect 11424 6001 11458 6050
rect 14553 5946 14587 5989
rect 8839 5724 8873 5762
rect 10061 5724 10095 5762
rect 10413 5724 10447 5762
rect 7277 5268 7311 5306
rect 12999 4664 13229 4688
rect 13033 4630 13067 4664
rect 13101 4630 13135 4664
rect 13169 4630 13229 4664
rect 12999 4595 13229 4630
rect 13033 4561 13067 4595
rect 13101 4561 13135 4595
rect 13169 4561 13229 4595
rect 12999 4526 13229 4561
rect 13033 4492 13067 4526
rect 13101 4492 13135 4526
rect 13169 4492 13229 4526
rect 12999 4457 13229 4492
rect 13033 4423 13067 4457
rect 13101 4423 13135 4457
rect 13169 4423 13229 4457
rect 12999 4418 13229 4423
rect 13177 4312 13229 4418
rect 13033 4285 13067 4312
rect 13101 4285 13135 4312
rect 13169 4285 13229 4312
rect 12999 4250 13229 4285
rect 13033 4216 13067 4250
rect 13101 4216 13135 4250
rect 13169 4216 13229 4250
rect 12999 4181 13229 4216
rect 13033 4147 13067 4181
rect 13101 4147 13135 4181
rect 13169 4147 13229 4181
rect 12999 4112 13229 4147
rect 13033 4078 13067 4112
rect 13101 4078 13135 4112
rect 13169 4078 13229 4112
rect 12999 4043 13229 4078
rect 13033 4009 13067 4043
rect 13101 4009 13135 4043
rect 13169 4009 13229 4043
rect 12999 3974 13229 4009
rect 13033 3940 13067 3974
rect 13101 3940 13135 3974
rect 13169 3940 13229 3974
rect 12999 3905 13229 3940
rect 13033 3871 13067 3905
rect 13101 3871 13135 3905
rect 13169 3871 13229 3905
rect 12999 3836 13229 3871
rect 13033 3802 13067 3836
rect 13101 3802 13135 3836
rect 13169 3802 13229 3836
rect 12999 3767 13229 3802
rect 13033 3733 13067 3767
rect 13101 3733 13135 3767
rect 13169 3733 13229 3767
rect 12999 3698 13229 3733
rect 13033 3664 13067 3698
rect 13101 3664 13135 3698
rect 13169 3664 13229 3698
rect 12999 3629 13229 3664
rect 13033 3595 13067 3629
rect 13101 3595 13135 3629
rect 13169 3595 13229 3629
rect 6843 3551 6881 3585
rect 12999 3560 13229 3595
rect 13033 3526 13067 3560
rect 13101 3526 13135 3560
rect 13169 3526 13229 3560
rect 10175 3427 10209 3465
rect 10175 3355 10209 3393
rect 12999 3491 13229 3526
rect 13033 3457 13067 3491
rect 13101 3457 13135 3491
rect 13169 3457 13229 3491
rect 12999 3422 13229 3457
rect 13033 3388 13067 3422
rect 13101 3388 13135 3422
rect 13169 3388 13229 3422
rect 12999 3353 13229 3388
rect 6669 3287 6703 3321
rect 13033 3319 13067 3353
rect 13101 3319 13135 3353
rect 13169 3319 13229 3353
rect 12999 3287 13229 3319
rect 12754 3284 13229 3287
rect 12754 3263 12999 3284
rect 12754 3229 12842 3263
rect 12876 3229 12910 3263
rect 12944 3250 12999 3263
rect 13033 3250 13067 3284
rect 13101 3250 13135 3284
rect 13169 3250 13229 3284
rect 12944 3229 13229 3250
rect 12754 3215 13229 3229
rect 12754 3185 12999 3215
rect 12754 3151 12842 3185
rect 12876 3151 12910 3185
rect 12944 3181 12999 3185
rect 13033 3181 13067 3215
rect 13101 3181 13135 3215
rect 13169 3181 13229 3215
rect 12944 3151 13229 3181
rect 12754 3146 13229 3151
rect 12754 3112 12999 3146
rect 13033 3112 13067 3146
rect 13101 3112 13135 3146
rect 13169 3112 13229 3146
rect 12754 3107 13229 3112
rect 12754 3073 12842 3107
rect 12876 3073 12910 3107
rect 12944 3077 13229 3107
rect 12944 3073 12999 3077
rect 12754 3043 12999 3073
rect 13033 3043 13067 3077
rect 13101 3043 13135 3077
rect 13169 3043 13229 3077
rect 12754 3029 13229 3043
rect 12754 2995 12842 3029
rect 12876 2995 12910 3029
rect 12944 3008 13229 3029
rect 12944 2995 12999 3008
rect 12754 2952 12999 2995
rect 12754 2918 12842 2952
rect 12876 2918 12910 2952
rect 12944 2918 12999 2952
rect 12754 2875 12999 2918
rect 12754 2841 12842 2875
rect 12876 2841 12910 2875
rect 12944 2841 12999 2875
rect 12754 2798 12999 2841
rect 12754 2764 12842 2798
rect 12876 2764 12910 2798
rect 12944 2764 12999 2798
rect 12754 2740 12999 2764
rect 13169 2702 13229 3008
rect 12999 2678 13229 2702
rect 15829 4664 16045 4688
rect 15829 4630 15852 4664
rect 15886 4630 15920 4664
rect 15954 4630 15988 4664
rect 16022 4630 16045 4664
rect 15829 4595 16045 4630
rect 15829 4561 15852 4595
rect 15886 4561 15920 4595
rect 15954 4561 15988 4595
rect 16022 4561 16045 4595
rect 15829 4526 16045 4561
rect 15829 4492 15852 4526
rect 15886 4492 15920 4526
rect 15954 4492 15988 4526
rect 16022 4492 16045 4526
rect 15829 4457 16045 4492
rect 15829 4423 15852 4457
rect 15886 4423 15920 4457
rect 15954 4423 15988 4457
rect 16022 4423 16045 4457
rect 15829 4388 16045 4423
rect 15829 4354 15852 4388
rect 15886 4354 15920 4388
rect 15954 4354 15988 4388
rect 16022 4354 16045 4388
rect 15829 4319 16045 4354
rect 15829 4285 15852 4319
rect 15886 4285 15920 4319
rect 15954 4285 15988 4319
rect 16022 4285 16045 4319
rect 15829 4250 16045 4285
rect 15829 4216 15852 4250
rect 15886 4216 15920 4250
rect 15954 4216 15988 4250
rect 16022 4216 16045 4250
rect 15829 4181 16045 4216
rect 15829 4147 15852 4181
rect 15886 4147 15920 4181
rect 15954 4147 15988 4181
rect 16022 4147 16045 4181
rect 15829 4112 16045 4147
rect 15829 4078 15852 4112
rect 15886 4078 15920 4112
rect 15954 4078 15988 4112
rect 16022 4078 16045 4112
rect 15829 4043 16045 4078
rect 15829 4009 15852 4043
rect 15886 4009 15920 4043
rect 15954 4009 15988 4043
rect 16022 4009 16045 4043
rect 15829 3974 16045 4009
rect 15829 3940 15852 3974
rect 15886 3940 15920 3974
rect 15954 3940 15988 3974
rect 16022 3940 16045 3974
rect 15829 3910 16045 3940
rect 15829 3905 15954 3910
rect 15829 3871 15852 3905
rect 15886 3871 15920 3905
rect 15829 3836 15954 3871
rect 15829 3802 15852 3836
rect 15886 3802 15920 3836
rect 15954 3802 15988 3804
rect 16022 3802 16045 3804
rect 15829 3767 16045 3802
rect 15829 3733 15852 3767
rect 15886 3733 15920 3767
rect 15954 3733 15988 3767
rect 16022 3733 16045 3767
rect 15829 3698 16045 3733
rect 15829 3664 15852 3698
rect 15886 3664 15920 3698
rect 15954 3664 15988 3698
rect 16022 3664 16045 3698
rect 15829 3629 16045 3664
rect 15829 2711 15852 3629
rect 16022 3557 16045 3629
rect 16022 3186 16144 3557
rect 16022 2711 16045 3186
rect 15829 2687 16045 2711
rect 7511 2385 7552 2431
rect 8232 2385 8273 2431
rect 11576 2414 11616 2431
rect 11576 2384 11710 2414
rect 15149 1901 15999 1965
rect 15149 1867 15173 1901
rect 15207 1867 15243 1901
rect 15277 1867 15313 1901
rect 15347 1867 15383 1901
rect 15417 1867 15453 1901
rect 15487 1867 15523 1901
rect 15557 1867 15593 1901
rect 15627 1867 15663 1901
rect 15697 1867 15733 1901
rect 15767 1867 15803 1901
rect 15837 1867 15872 1901
rect 15906 1867 15941 1901
rect 15975 1867 15999 1901
<< viali >>
rect 7538 8847 7572 8881
rect 7610 8847 7644 8881
rect 8199 8773 8233 8807
rect 8271 8773 8305 8807
rect 8343 8773 8377 8807
rect 13113 6070 13147 6104
rect 13185 6070 13219 6104
rect 8839 5762 8873 5796
rect 5473 5693 5507 5727
rect 8839 5690 8873 5724
rect 10061 5762 10095 5796
rect 10061 5690 10095 5724
rect 10413 5762 10447 5796
rect 10413 5690 10447 5724
rect 7277 5306 7311 5340
rect 7277 5234 7311 5268
rect 12999 4388 13177 4418
rect 12999 4354 13033 4388
rect 13033 4354 13067 4388
rect 13067 4354 13101 4388
rect 13101 4354 13135 4388
rect 13135 4354 13169 4388
rect 13169 4354 13177 4388
rect 12999 4319 13177 4354
rect 12999 4312 13033 4319
rect 13033 4312 13067 4319
rect 13067 4312 13101 4319
rect 13101 4312 13135 4319
rect 13135 4312 13169 4319
rect 13169 4312 13177 4319
rect 6809 3551 6843 3585
rect 6881 3551 6915 3585
rect 10175 3465 10209 3499
rect 10175 3393 10209 3427
rect 10175 3321 10209 3355
rect 15954 3905 16060 3910
rect 15954 3871 15988 3905
rect 15988 3871 16022 3905
rect 16022 3871 16060 3905
rect 15954 3836 16060 3871
rect 15954 3804 15988 3836
rect 15988 3804 16022 3836
rect 16022 3804 16060 3836
<< metal1 >>
rect 8153 10649 8159 10673
rect 8108 10621 8159 10649
rect 8211 10621 8223 10673
rect 8275 10649 8281 10673
rect 8275 10621 14707 10649
rect -11 9733 -5 9849
rect 111 9733 117 9849
rect 8153 9669 8449 9675
rect 8205 9623 8397 9669
rect 8153 9605 8205 9617
rect 8153 9547 8205 9553
rect 8397 9605 8449 9617
rect 8397 9547 8449 9553
tri 7150 9466 7175 9491 ne
rect 7175 9467 7181 9519
rect 7233 9467 7239 9519
rect 7175 9455 7239 9467
tri 7239 9466 7264 9491 nw
rect 7175 9403 7181 9455
rect 7233 9403 7239 9455
rect 7872 9423 7906 9457
rect 9102 9417 9148 9463
rect 13703 9455 13742 9491
rect 10098 9375 10138 9421
rect 7668 9299 7708 9345
rect 9983 9341 10035 9347
tri 9958 9265 9983 9290 se
rect 9983 9277 10035 9289
rect 4190 9219 4230 9265
rect 5902 9219 5943 9265
tri 10035 9265 10060 9290 sw
rect 9983 9219 10035 9225
rect -11 9011 -5 9191
rect 111 9011 117 9191
rect 66 8909 607 8961
rect 659 8909 671 8961
rect 723 8909 729 8961
rect 6779 8840 6831 8846
rect 7015 8835 7021 8887
rect 7073 8835 7085 8887
rect 7137 8881 7656 8887
rect 7137 8847 7538 8881
rect 7572 8847 7610 8881
rect 7644 8847 7656 8881
rect 7137 8841 7656 8847
rect 7137 8835 7143 8841
tri 7143 8835 7149 8841 nw
rect 6779 8776 6831 8788
tri 6831 8773 6841 8783 sw
rect 6831 8761 6841 8773
tri 6841 8761 6853 8773 sw
rect 7445 8761 7451 8813
rect 7503 8761 7515 8813
rect 7567 8807 8389 8813
rect 7567 8773 8199 8807
rect 8233 8773 8271 8807
rect 8305 8773 8343 8807
rect 8377 8773 8389 8807
rect 7567 8761 8389 8773
rect 6831 8758 6853 8761
tri 6853 8758 6856 8761 sw
rect 6831 8733 6916 8758
tri 6916 8733 6941 8758 sw
tri 9739 8733 9764 8758 se
rect 9764 8757 9770 8809
rect 9822 8757 9828 8809
rect 9764 8745 9828 8757
rect 9764 8733 9770 8745
rect 6831 8724 9770 8733
rect 6779 8718 9770 8724
tri 6898 8693 6923 8718 ne
rect 6923 8693 9770 8718
rect 9822 8693 9828 8745
rect 7445 8331 7497 8337
rect 10333 8331 10385 8337
rect 7445 8267 7497 8279
tri 7497 8258 7522 8283 sw
tri 10308 8258 10333 8283 se
rect 10333 8267 10385 8279
rect 7497 8215 10333 8258
rect 7445 8209 10385 8215
rect 0 8051 42 8181
rect 9697 7593 9706 7645
rect 9758 7593 9770 7645
rect 9822 7593 9828 7645
rect 6755 7270 6807 7276
tri 6730 7200 6755 7225 se
rect 9535 7230 9575 7271
rect 6755 7206 6807 7218
rect 1393 7148 1399 7200
rect 1451 7148 1463 7200
rect 1515 7154 6755 7200
rect 1515 7148 6807 7154
rect -11 6860 -5 7040
rect 111 6860 117 7040
rect 5504 6542 5510 6594
rect 5562 6542 5574 6594
rect 5626 6542 7021 6594
rect 7073 6542 7085 6594
rect 7137 6542 7143 6594
rect 12223 6232 14428 6284
tri 14406 6219 14419 6232 ne
rect 14419 6219 14428 6232
tri 14428 6219 14493 6284 sw
tri 14419 6210 14428 6219 ne
rect 14428 6210 14493 6219
tri 14428 6197 14441 6210 ne
rect 2389 6066 2419 6096
rect 9432 6058 9438 6110
rect 9490 6104 13231 6110
rect 9490 6070 13113 6104
rect 13147 6070 13185 6104
rect 13219 6070 13231 6104
rect 9490 6058 13231 6070
rect 9432 6046 9496 6058
rect 9432 5994 9438 6046
rect 9490 5994 9496 6046
rect 223 5946 257 5982
rect 14441 5882 14493 6210
rect 15516 5934 15568 5940
tri 14441 5876 14447 5882 ne
rect 14447 5876 14493 5882
rect 2868 5841 2903 5876
tri 14447 5866 14457 5876 ne
rect 14457 5866 14493 5876
tri 14493 5866 14531 5904 sw
tri 15491 5866 15516 5891 se
rect 15516 5870 15568 5882
tri 14457 5841 14482 5866 ne
rect 14482 5841 15516 5866
tri 14482 5830 14493 5841 ne
rect 14493 5830 15516 5841
tri 14493 5814 14509 5830 ne
rect 14509 5818 15516 5830
rect 14509 5814 15568 5818
tri 15514 5812 15516 5814 ne
rect 15516 5812 15568 5814
rect 8830 5800 8882 5808
rect 563 5756 597 5790
rect 5460 5727 5510 5739
rect 5460 5693 5473 5727
rect 5507 5693 5510 5727
rect 5460 5687 5510 5693
rect 5562 5687 5568 5739
rect 8830 5736 8882 5748
rect 8830 5678 8882 5684
rect 10040 5802 10101 5808
rect 10092 5796 10101 5802
rect 10095 5762 10101 5796
rect 10092 5750 10101 5762
rect 10040 5738 10101 5750
rect 10092 5724 10101 5738
rect 10095 5690 10101 5724
rect 10092 5686 10101 5690
rect 10040 5678 10101 5686
rect 10333 5802 10453 5808
rect 10385 5796 10453 5802
rect 10385 5762 10413 5796
rect 10447 5762 10453 5796
rect 10385 5750 10453 5762
rect 10333 5738 10453 5750
rect 10385 5724 10453 5738
rect 10385 5690 10413 5724
rect 10447 5690 10453 5724
rect 10385 5686 10453 5690
rect 10333 5678 10453 5686
rect 7265 5294 7271 5346
rect 7323 5294 7329 5346
rect 7265 5282 7329 5294
rect 7265 5230 7271 5282
rect 7323 5230 7329 5282
rect 8988 5275 8994 5327
rect 9046 5275 9058 5327
rect 9110 5275 9374 5327
rect 9426 5275 9438 5327
rect 9490 5275 9496 5327
rect 7265 5228 7329 5230
tri 12954 5198 12979 5223 se
rect 12979 5152 12985 5268
rect 13101 5152 13107 5268
tri 13107 5198 13132 5223 sw
rect -54 5124 14914 5152
rect -54 4922 -29 5124
rect 349 4850 380 4883
rect 3400 4824 3434 4858
rect 4153 4697 4193 4737
rect -11 4458 0 4660
rect 6237 4458 6277 4660
rect 16029 4458 16040 4660
rect -17 4300 0 4430
rect 530 4305 536 4421
rect 652 4305 658 4421
rect 4622 4369 4628 4421
rect 4680 4369 4686 4421
rect 4622 4357 4686 4369
rect 4622 4305 4628 4357
rect 4680 4305 4686 4357
rect 12979 4314 12985 4430
rect 13101 4418 13183 4430
rect 12993 4312 12999 4314
rect 13177 4312 13183 4418
rect 12993 4300 13183 4312
rect 16023 4300 16040 4430
tri 13692 4275 13717 4300 ne
rect 13717 4192 13763 4300
tri 13763 4275 13788 4300 nw
rect 242 4122 708 4174
rect 760 4122 772 4174
rect 824 4122 1831 4174
rect 6787 4140 6793 4192
rect 6845 4140 6857 4192
rect 6909 4140 13121 4192
tri 13121 4140 13173 4192 sw
tri 13099 4126 13113 4140 ne
rect 13113 4126 13173 4140
tri 13173 4126 13187 4140 sw
tri 1675 4096 1701 4122 ne
rect 1701 4093 1831 4122
tri 13113 4118 13121 4126 ne
rect 13121 4118 13187 4126
tri 13121 4100 13139 4118 ne
rect 13139 4100 13187 4118
rect 12390 4048 12434 4100
tri 13139 4093 13146 4100 ne
rect 13146 4093 13187 4100
tri 13187 4093 13220 4126 sw
tri 13146 4052 13187 4093 ne
rect 13187 4052 13220 4093
tri 13220 4052 13261 4093 sw
rect 16030 4070 16040 4272
tri 13187 4048 13191 4052 ne
rect 13191 4048 13261 4052
tri 13191 3978 13261 4048 ne
tri 13261 4038 13275 4052 sw
rect 13261 4015 13275 4038
tri 13275 4015 13298 4038 sw
rect 15436 4032 15488 4038
rect 13261 3978 13298 4015
tri 13298 3978 13335 4015 sw
tri 15399 3978 15436 4015 se
rect 15436 3978 15488 3980
tri 13261 3962 13277 3978 ne
rect 13277 3962 14298 3978
tri 14298 3962 14314 3978 sw
tri 15383 3962 15399 3978 se
rect 15399 3968 15488 3978
rect 15399 3962 15436 3968
tri 13277 3926 13313 3962 ne
rect 13313 3926 15436 3962
tri 14276 3910 14292 3926 ne
rect 14292 3916 15436 3926
rect 14292 3910 15488 3916
rect 15944 3769 15950 3949
rect 16066 3769 16072 3949
rect 99 3667 133 3701
rect 4071 3667 4105 3701
rect 6797 3585 8994 3591
rect 6797 3551 6809 3585
rect 6843 3551 6881 3585
rect 6915 3551 8994 3585
rect 6797 3539 8994 3551
rect 9046 3539 9058 3591
rect 9110 3539 9116 3591
rect -51 3511 6306 3539
tri 6306 3511 6334 3539 sw
rect -51 3309 14 3511
rect 6237 3309 6277 3511
rect 6306 3505 6334 3511
tri 6334 3505 6340 3511 sw
rect 6306 3499 6340 3505
tri 6340 3499 6346 3505 sw
rect 10163 3499 10221 3505
rect 6306 3489 6346 3499
tri 6346 3489 6356 3499 sw
rect 6306 3465 6356 3489
tri 6356 3465 6380 3489 sw
rect 6306 3459 6380 3465
tri 6380 3459 6386 3465 sw
rect 6546 3437 6552 3489
rect 6604 3437 6610 3489
rect 6546 3425 6610 3437
rect 6546 3373 6552 3425
rect 6604 3373 6610 3425
rect 6546 3361 6610 3373
rect 6546 3309 6552 3361
rect 6604 3309 6610 3361
rect 10163 3465 10175 3499
rect 10209 3465 10221 3499
rect 10163 3427 10221 3465
rect 10163 3393 10175 3427
rect 10209 3393 10221 3427
rect 10163 3355 10221 3393
rect 10163 3321 10175 3355
rect 10209 3321 10221 3355
rect 10163 3315 10221 3321
rect 16027 3309 16081 3511
rect 21817 3309 21857 3511
rect 5404 3236 5438 3278
tri 6709 2961 6734 2986 sw
tri 6866 2961 6891 2986 se
rect 6709 2903 6891 2961
tri 12237 2961 12262 2986 sw
tri 12394 2961 12419 2986 se
rect 12237 2903 12419 2961
rect 12774 2903 12879 3249
rect 185 2664 196 2866
rect -2 2518 16 2636
rect 8956 2450 8989 2483
rect 10128 2450 10162 2484
rect 4759 2278 4826 2330
rect 4878 2278 4890 2330
rect 4942 2278 8160 2330
tri 16867 2278 16873 2284 se
rect 16873 2278 17554 2284
tri 16839 2250 16867 2278 se
rect 16867 2250 17554 2278
rect 15436 2244 17554 2250
rect 15488 2232 17554 2244
rect 15488 2198 16861 2232
tri 16861 2198 16895 2232 nw
rect 15436 2180 15488 2192
tri 15488 2173 15513 2198 nw
rect 15436 2122 15488 2128
rect 15516 2155 15568 2161
tri 15568 2124 15593 2149 sw
rect 15568 2103 17239 2124
rect 15516 2091 17239 2103
rect 15568 2072 17239 2091
tri 15568 2047 15593 2072 nw
rect 15516 2033 15568 2039
rect 16003 1997 16072 1998
rect 15944 1881 15950 1997
rect 16066 1881 16072 1997
rect 16003 1880 16072 1881
rect 16145 1842 16185 2044
rect 22257 1842 22297 2044
<< via1 >>
rect 8159 10621 8211 10673
rect 8223 10621 8275 10673
rect -5 9733 111 9849
rect 8153 9617 8205 9669
rect 8153 9553 8205 9605
rect 8397 9617 8449 9669
rect 8397 9553 8449 9605
rect 7181 9467 7233 9519
rect 7181 9403 7233 9455
rect 9983 9289 10035 9341
rect 9983 9225 10035 9277
rect -5 9011 111 9191
rect 607 8909 659 8961
rect 671 8909 723 8961
rect 6779 8788 6831 8840
rect 7021 8835 7073 8887
rect 7085 8835 7137 8887
rect 6779 8724 6831 8776
rect 7451 8761 7503 8813
rect 7515 8761 7567 8813
rect 9770 8757 9822 8809
rect 9770 8693 9822 8745
rect 7445 8279 7497 8331
rect 7445 8215 7497 8267
rect 10333 8279 10385 8331
rect 10333 8215 10385 8267
rect 9706 7593 9758 7645
rect 9770 7593 9822 7645
rect 6755 7218 6807 7270
rect 1399 7148 1451 7200
rect 1463 7148 1515 7200
rect 6755 7154 6807 7206
rect -5 6860 111 7040
rect 5510 6542 5562 6594
rect 5574 6542 5626 6594
rect 7021 6542 7073 6594
rect 7085 6542 7137 6594
rect 9438 6058 9490 6110
rect 9438 5994 9490 6046
rect 15516 5882 15568 5934
rect 15516 5818 15568 5870
rect 8830 5796 8882 5800
rect 8830 5762 8839 5796
rect 8839 5762 8873 5796
rect 8873 5762 8882 5796
rect 8830 5748 8882 5762
rect 5510 5687 5562 5739
rect 8830 5724 8882 5736
rect 8830 5690 8839 5724
rect 8839 5690 8873 5724
rect 8873 5690 8882 5724
rect 8830 5684 8882 5690
rect 10040 5796 10092 5802
rect 10040 5762 10061 5796
rect 10061 5762 10092 5796
rect 10040 5750 10092 5762
rect 10040 5724 10092 5738
rect 10040 5690 10061 5724
rect 10061 5690 10092 5724
rect 10040 5686 10092 5690
rect 10333 5750 10385 5802
rect 10333 5686 10385 5738
rect 7271 5340 7323 5346
rect 7271 5306 7277 5340
rect 7277 5306 7311 5340
rect 7311 5306 7323 5340
rect 7271 5294 7323 5306
rect 7271 5268 7323 5282
rect 7271 5234 7277 5268
rect 7277 5234 7311 5268
rect 7311 5234 7323 5268
rect 7271 5230 7323 5234
rect 8994 5275 9046 5327
rect 9058 5275 9110 5327
rect 9374 5275 9426 5327
rect 9438 5275 9490 5327
rect 12985 5152 13101 5268
rect 536 4305 652 4421
rect 4628 4369 4680 4421
rect 4628 4305 4680 4357
rect 12985 4418 13101 4430
rect 12985 4314 12999 4418
rect 12999 4314 13101 4418
rect 708 4122 760 4174
rect 772 4122 824 4174
rect 6793 4140 6845 4192
rect 6857 4140 6909 4192
rect 15436 3980 15488 4032
rect 15436 3916 15488 3968
rect 15950 3910 16066 3949
rect 15950 3804 15954 3910
rect 15954 3804 16060 3910
rect 16060 3804 16066 3910
rect 15950 3769 16066 3804
rect 8994 3539 9046 3591
rect 9058 3539 9110 3591
rect 6552 3437 6604 3489
rect 6552 3373 6604 3425
rect 6552 3309 6604 3361
rect 4826 2278 4878 2330
rect 4890 2278 4942 2330
rect 15436 2192 15488 2244
rect 15436 2128 15488 2180
rect 15516 2103 15568 2155
rect 15516 2039 15568 2091
rect 15950 1881 16066 1997
<< metal2 >>
rect 8153 10621 8159 10673
rect 8211 10621 8223 10673
rect 8275 10621 8281 10673
rect -11 9733 -5 9849
rect 111 9733 117 9849
rect -11 9191 117 9733
rect 8153 9669 8205 10621
rect 8153 9605 8205 9617
rect 8153 9547 8205 9553
rect 8397 9669 8449 9675
rect 8397 9605 8449 9617
rect 8397 9547 8449 9553
rect -11 9011 -5 9191
rect 111 9011 117 9191
rect -11 7040 117 9011
rect 7175 9467 7181 9519
rect 7233 9467 7239 9519
rect 7175 9455 7239 9467
rect 7175 9403 7181 9455
rect 7233 9403 7239 9455
rect 601 8909 607 8961
rect 659 8909 671 8961
rect 723 8909 729 8961
tri 652 8887 674 8909 ne
rect 674 8887 729 8909
tri 674 8884 677 8887 ne
rect -11 6860 -5 7040
rect 111 6860 117 7040
rect -11 5650 117 6860
rect 677 6131 729 8887
rect 6779 8840 6831 8846
rect 6875 8821 6927 8873
rect 7015 8835 7021 8887
rect 7073 8835 7085 8887
rect 7137 8835 7143 8887
tri 7066 8821 7080 8835 ne
rect 7080 8821 7143 8835
tri 7080 8813 7088 8821 ne
rect 7088 8813 7143 8821
tri 7088 8810 7091 8813 ne
rect 6779 8776 6831 8788
tri 6757 8553 6779 8575 se
rect 6779 8553 6831 8724
tri 6719 8515 6757 8553 se
rect 6757 8515 6771 8553
rect 6719 7803 6771 8515
tri 6771 8493 6831 8553 nw
tri 6809 7825 6821 7837 ne
rect 6821 7825 6887 7837
tri 6719 7789 6733 7803 ne
rect 6733 7789 6771 7803
tri 6771 7789 6807 7825 sw
tri 6821 7811 6835 7825 ne
tri 6733 7767 6755 7789 ne
rect 6755 7270 6807 7789
rect 6755 7206 6807 7218
rect 1393 7148 1399 7200
rect 1451 7148 1463 7200
rect 1515 7148 1521 7200
rect 6755 7148 6807 7154
tri 1371 6170 1393 6192 se
rect 1393 6170 1445 7148
tri 1445 7123 1470 7148 nw
tri 1364 6163 1371 6170 se
rect 1371 6163 1416 6170
tri 729 6131 740 6142 sw
rect 677 6110 740 6131
tri 740 6110 761 6131 sw
rect 677 6104 761 6110
tri 677 6058 723 6104 ne
rect 723 6058 761 6104
tri 761 6058 813 6110 sw
tri 723 6046 735 6058 ne
rect 735 6046 813 6058
tri 813 6046 825 6058 sw
tri 735 6041 740 6046 ne
rect 740 6041 825 6046
tri 825 6041 830 6046 sw
tri 740 6015 766 6041 ne
rect 566 5093 622 5102
rect 566 5013 622 5037
rect 566 4933 622 4957
rect 566 4853 622 4877
rect 566 4773 622 4797
rect 566 4693 622 4717
rect 566 4628 622 4637
rect 530 4305 536 4421
rect 652 4305 658 4421
tri 759 4192 766 4199 se
rect 766 4192 830 6041
rect 1364 4292 1416 6163
tri 1416 6141 1445 6170 nw
rect 5504 6542 5510 6594
rect 5562 6542 5574 6594
rect 5626 6542 5632 6594
rect 5504 5739 5568 6542
tri 5568 6517 5593 6542 nw
rect 5504 5687 5510 5739
rect 5562 5687 5568 5739
rect 3728 5093 3784 5102
rect 3728 5013 3784 5037
rect 3728 4933 3784 4957
rect 3728 4853 3784 4877
rect 3728 4773 3784 4797
rect 3728 4693 3784 4717
rect 3728 4628 3784 4637
rect 4626 5093 4682 5102
rect 4626 5013 4682 5037
rect 4626 4933 4682 4957
rect 4626 4853 4682 4877
rect 4626 4773 4682 4797
rect 4626 4693 4682 4717
rect 4626 4628 4682 4637
rect 4622 4369 4628 4421
rect 4680 4369 4686 4421
rect 4622 4357 4686 4369
rect 4622 4305 4628 4357
rect 4680 4305 4686 4357
tri 1416 4292 1422 4298 sw
rect 1364 4276 1422 4292
tri 1364 4218 1422 4276 ne
tri 1422 4218 1496 4292 sw
tri 1422 4217 1423 4218 ne
rect 1423 4217 1496 4218
tri 1423 4199 1441 4217 ne
rect 1441 4199 1496 4217
tri 1441 4196 1444 4199 ne
tri 741 4174 759 4192 se
rect 759 4174 830 4192
rect 702 4122 708 4174
rect 760 4122 772 4174
rect 824 4122 830 4174
rect 1444 4035 1496 4199
rect 4740 4140 4786 4688
tri 6834 4217 6835 4218 se
rect 6835 4217 6887 7825
tri 6887 7811 6913 7837 nw
tri 7066 6594 7091 6619 se
rect 7091 6594 7143 8813
rect 7015 6542 7021 6594
rect 7073 6542 7085 6594
rect 7137 6542 7143 6594
rect 7175 6198 7239 9403
rect 7445 8761 7451 8813
rect 7503 8761 7515 8813
rect 7567 8761 7573 8813
rect 7445 8757 7518 8761
tri 7518 8757 7522 8761 nw
rect 7445 8745 7506 8757
tri 7506 8745 7518 8757 nw
rect 7445 8331 7497 8745
tri 7497 8736 7506 8745 nw
rect 7445 8267 7497 8279
rect 7445 8209 7497 8215
rect 8397 7353 8425 9547
rect 9983 9341 10035 9347
rect 9983 9277 10035 9289
rect 9983 8809 10035 9225
rect 10365 8972 10384 8977
rect 10324 8909 10382 8961
tri 10035 8809 10048 8822 sw
rect 9764 8757 9770 8809
rect 9822 8757 9828 8809
rect 9983 8800 10048 8809
tri 9983 8765 10018 8800 ne
rect 10018 8765 10048 8800
tri 10048 8765 10092 8809 sw
rect 9764 8745 9828 8757
tri 10018 8748 10035 8765 ne
rect 10035 8748 10092 8765
rect 9764 8693 9770 8745
rect 9822 8693 9828 8745
tri 10035 8743 10040 8748 ne
tri 9739 7645 9764 7670 se
rect 9764 7645 9828 8693
rect 9700 7593 9706 7645
rect 9758 7593 9770 7645
rect 9822 7593 9828 7645
tri 8397 7352 8398 7353 ne
rect 8398 7352 8425 7353
tri 8425 7352 8448 7375 sw
tri 8398 7325 8425 7352 ne
rect 8425 7325 8448 7352
tri 8425 7302 8448 7325 ne
tri 8448 7302 8498 7352 sw
tri 8448 7280 8470 7302 ne
rect 8470 6279 8498 7302
tri 8498 6279 8508 6289 sw
rect 8470 6269 8508 6279
tri 8508 6269 8518 6279 sw
tri 8470 6231 8508 6269 ne
rect 8508 6259 8518 6269
tri 8518 6259 8528 6269 sw
rect 8508 6231 8866 6259
tri 7175 6141 7232 6198 ne
rect 7232 6141 7239 6198
tri 7239 6141 7322 6224 sw
tri 7232 6134 7239 6141 ne
rect 7239 6134 7322 6141
tri 7322 6134 7329 6141 sw
tri 7239 6110 7263 6134 ne
rect 7263 6110 7329 6134
tri 7263 6108 7265 6110 ne
rect 7265 5346 7329 6110
rect 8838 5806 8866 6231
rect 9432 6058 9438 6110
rect 9490 6058 9496 6110
rect 9432 6046 9496 6058
rect 9432 5994 9438 6046
rect 9490 5994 9496 6046
rect 8830 5800 8882 5806
rect 8830 5736 8882 5748
rect 8830 5678 8882 5684
rect 7265 5294 7271 5346
rect 7323 5294 7329 5346
rect 9432 5327 9496 5994
rect 10040 5802 10092 8748
rect 10040 5738 10092 5750
rect 10040 5680 10092 5686
rect 10333 8331 10385 8337
rect 10333 8267 10385 8279
rect 10333 5802 10385 8215
rect 10333 5738 10385 5750
rect 10333 5678 10385 5686
rect 15516 5934 15568 5940
rect 15516 5870 15568 5882
rect 7265 5282 7329 5294
rect 7265 5230 7271 5282
rect 7323 5230 7329 5282
rect 8988 5275 8994 5327
rect 9046 5275 9058 5327
rect 9110 5275 9116 5327
rect 9368 5275 9374 5327
rect 9426 5275 9438 5327
rect 9490 5275 9496 5327
tri 6809 4192 6834 4217 se
rect 6834 4199 6887 4217
tri 6887 4199 6905 4217 sw
rect 6834 4192 6905 4199
tri 6905 4192 6912 4199 sw
rect 6787 4140 6793 4192
rect 6845 4140 6857 4192
rect 6909 4140 6915 4192
tri 4791 4115 4816 4140 ne
tri 1496 4079 1521 4104 sw
tri 4750 3194 4816 3260 se
rect 4816 3240 4862 4140
tri 4862 4134 4868 4140 nw
rect 8988 3591 9040 5275
rect 12979 5152 12985 5268
rect 13101 5152 13107 5268
rect 12979 4430 13107 5152
rect 12979 4314 12985 4430
rect 13101 4314 13107 4430
rect 10805 4298 11362 4301
tri 11362 4298 11365 4301 nw
rect 10805 4292 11356 4298
tri 11356 4292 11362 4298 nw
rect 10805 4217 11281 4292
tri 11281 4217 11356 4292 nw
rect 10805 4199 11263 4217
tri 11263 4199 11281 4217 nw
rect 10805 4192 11256 4199
tri 11256 4192 11263 4199 nw
rect 10805 4140 11204 4192
tri 11204 4140 11256 4192 nw
rect 10805 4104 11168 4140
tri 11168 4104 11204 4140 nw
tri 9040 3591 9065 3616 sw
rect 8988 3539 8994 3591
rect 9046 3539 9058 3591
rect 9110 3539 9116 3591
rect 6546 3437 6552 3489
rect 6604 3437 6610 3489
rect 6546 3425 6610 3437
rect 6546 3373 6552 3425
rect 6604 3373 6610 3425
rect 6546 3361 6610 3373
rect 6546 3309 6552 3361
rect 6604 3309 6610 3361
rect 10805 3309 11165 4104
tri 11165 4101 11168 4104 nw
rect 15436 4032 15488 4038
rect 15436 3968 15488 3980
tri 4816 3194 4862 3240 nw
tri 4740 3184 4750 3194 se
rect 4750 3184 4806 3194
tri 4806 3184 4816 3194 nw
rect 4740 3054 4786 3184
tri 4786 3164 4806 3184 nw
tri 4786 3054 4806 3074 sw
tri 4740 2988 4806 3054 ne
tri 4806 2994 4866 3054 sw
rect 4806 2988 4866 2994
tri 4806 2974 4820 2988 ne
rect 4820 2330 4866 2988
tri 4866 2330 4891 2355 sw
rect 4820 2278 4826 2330
rect 4878 2278 4890 2330
rect 4942 2278 5014 2330
rect 12545 2303 12863 2335
rect 15436 2244 15488 3916
rect 15436 2180 15488 2192
rect 15436 2122 15488 2128
rect 15516 2155 15568 5818
rect 15944 3769 15950 3949
rect 16066 3769 16072 3949
rect 15991 3191 16025 3225
rect 15516 2091 15568 2103
rect 15516 2033 15568 2039
rect 15944 1997 16072 2894
rect 15944 1881 15950 1997
rect 16066 1881 16072 1997
<< via2 >>
rect 566 5037 622 5093
rect 566 4957 622 5013
rect 566 4877 622 4933
rect 566 4797 622 4853
rect 566 4717 622 4773
rect 566 4637 622 4693
rect 3728 5037 3784 5093
rect 3728 4957 3784 5013
rect 3728 4877 3784 4933
rect 3728 4797 3784 4853
rect 3728 4717 3784 4773
rect 3728 4637 3784 4693
rect 4626 5037 4682 5093
rect 4626 4957 4682 5013
rect 4626 4877 4682 4933
rect 4626 4797 4682 4853
rect 4626 4717 4682 4773
rect 4626 4637 4682 4693
<< metal3 >>
rect 561 5093 627 5098
rect 561 5037 566 5093
rect 622 5037 627 5093
rect 561 5013 627 5037
rect 561 4957 566 5013
rect 622 4957 627 5013
rect 561 4933 627 4957
rect 561 4877 566 4933
rect 622 4877 627 4933
rect 561 4853 627 4877
rect 561 4797 566 4853
rect 622 4797 627 4853
rect 561 4773 627 4797
rect 561 4717 566 4773
rect 622 4717 627 4773
rect 561 4693 627 4717
rect 561 4637 566 4693
rect 622 4637 627 4693
rect 561 4632 627 4637
rect 3723 5093 3789 5098
rect 3723 5037 3728 5093
rect 3784 5037 3789 5093
rect 3723 5013 3789 5037
rect 3723 4957 3728 5013
rect 3784 4957 3789 5013
rect 3723 4933 3789 4957
rect 3723 4877 3728 4933
rect 3784 4877 3789 4933
rect 3723 4853 3789 4877
rect 3723 4797 3728 4853
rect 3784 4797 3789 4853
rect 3723 4773 3789 4797
rect 3723 4717 3728 4773
rect 3784 4717 3789 4773
rect 3723 4693 3789 4717
rect 3723 4637 3728 4693
rect 3784 4637 3789 4693
rect 3723 4632 3789 4637
rect 4621 5093 4687 5098
rect 4621 5037 4626 5093
rect 4682 5037 4687 5093
rect 4621 5013 4687 5037
rect 4621 4957 4626 5013
rect 4682 4957 4687 5013
rect 4621 4933 4687 4957
rect 4621 4877 4626 4933
rect 4682 4877 4687 4933
rect 4621 4853 4687 4877
rect 4621 4797 4626 4853
rect 4682 4797 4687 4853
rect 4621 4773 4687 4797
rect 4621 4717 4626 4773
rect 4682 4717 4687 4773
rect 4621 4693 4687 4717
rect 4621 4637 4626 4693
rect 4682 4637 4687 4693
rect 4621 4632 4687 4637
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1707688321
transform 1 0 7277 0 -1 5340
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1707688321
transform 0 -1 10447 -1 0 5796
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1707688321
transform -1 0 6915 0 1 3551
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1707688321
transform 0 -1 10095 1 0 5690
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1707688321
transform 1 0 13113 0 -1 6104
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1707688321
transform 1 0 7538 0 1 8847
box 0 0 1 1
use L1M1_CDNS_5246887918558  L1M1_CDNS_5246887918558_0
timestamp 1707688321
transform 0 1 12999 -1 0 4418
box 0 0 1 1
use L1M1_CDNS_5246887918559  L1M1_CDNS_5246887918559_0
timestamp 1707688321
transform 0 1 15954 1 0 3804
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1707688321
transform 1 0 8199 0 1 8773
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_0
timestamp 1707688321
transform 1 0 10175 0 1 3321
box 0 0 1 1
use L1M1_CDNS_52468879185302  L1M1_CDNS_52468879185302_0
timestamp 1707688321
transform 1 0 12999 0 1 3317
box -12 -6 262 184
use L1M1_CDNS_52468879185449  L1M1_CDNS_52468879185449_0
timestamp 1707688321
transform 0 1 15817 -1 0 4418
box -12 -6 118 256
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_0
timestamp 1707688321
transform -1 0 5507 0 -1 5727
box 0 0 1 1
use L1M1_CDNS_524688791851397  L1M1_CDNS_524688791851397_0
timestamp 1707688321
transform -1 0 15991 0 -1 1992
box -12 -6 838 112
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1707688321
transform 0 -1 10092 -1 0 5808
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1707688321
transform 0 -1 10385 -1 0 5808
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1707688321
transform 0 -1 6807 -1 0 7276
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1707688321
transform 0 -1 6831 -1 0 8846
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1707688321
transform 0 -1 15488 -1 0 2250
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_5
timestamp 1707688321
transform 0 -1 15488 -1 0 4038
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_6
timestamp 1707688321
transform 0 1 15516 -1 0 2161
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_7
timestamp 1707688321
transform -1 0 9116 0 1 3539
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_8
timestamp 1707688321
transform -1 0 9116 0 -1 5327
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_9
timestamp 1707688321
transform -1 0 9496 0 -1 5327
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_10
timestamp 1707688321
transform 0 1 10333 1 0 8209
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_11
timestamp 1707688321
transform 0 -1 10035 1 0 9219
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_12
timestamp 1707688321
transform 0 -1 7497 1 0 8209
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_13
timestamp 1707688321
transform 0 -1 15568 1 0 5812
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_14
timestamp 1707688321
transform 1 0 6787 0 -1 4192
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_15
timestamp 1707688321
transform 1 0 4820 0 -1 2330
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_16
timestamp 1707688321
transform 1 0 7015 0 -1 6594
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_17
timestamp 1707688321
transform 1 0 702 0 1 4122
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_18
timestamp 1707688321
transform 1 0 601 0 1 8909
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_19
timestamp 1707688321
transform 1 0 5504 0 1 6542
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_20
timestamp 1707688321
transform 1 0 7015 0 1 8835
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_21
timestamp 1707688321
transform 1 0 7445 0 1 8761
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_22
timestamp 1707688321
transform 1 0 9700 0 1 7593
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_23
timestamp 1707688321
transform 1 0 1393 0 1 7148
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_0
timestamp 1707688321
transform -1 0 13107 0 -1 4430
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_1
timestamp 1707688321
transform -1 0 16072 0 -1 1997
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_2
timestamp 1707688321
transform 1 0 -11 0 -1 9849
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_3
timestamp 1707688321
transform 1 0 12979 0 1 5152
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_4
timestamp 1707688321
transform 1 0 530 0 1 4305
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_0
timestamp 1707688321
transform -1 0 16072 0 -1 3949
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_1
timestamp 1707688321
transform 1 0 -11 0 -1 7040
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_2
timestamp 1707688321
transform 1 0 -11 0 -1 9191
box 0 0 1 1
use M1M2_CDNS_52468879185201  M1M2_CDNS_52468879185201_0
timestamp 1707688321
transform 1 0 8015 0 1 4305
box 0 0 320 116
use M1M2_CDNS_52468879185201  M1M2_CDNS_52468879185201_1
timestamp 1707688321
transform 1 0 6987 0 1 4305
box 0 0 320 116
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_0
timestamp 1707688321
transform -1 0 9496 0 -1 6110
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_1
timestamp 1707688321
transform -1 0 9828 0 -1 8809
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_2
timestamp 1707688321
transform 1 0 7265 0 -1 5346
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_3
timestamp 1707688321
transform 1 0 7175 0 -1 9519
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_4
timestamp 1707688321
transform 1 0 4622 0 1 4305
box 0 0 1 1
use M1M2_CDNS_52468879185371  M1M2_CDNS_52468879185371_0
timestamp 1707688321
transform 1 0 6546 0 1 3309
box 0 0 1 1
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_0
timestamp 1707688321
transform 1 0 5504 0 -1 5739
box 0 0 1 1
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_0
timestamp 1707688321
transform 1 0 10825 0 1 3314
box 0 0 320 180
use M1M2_CDNS_524688791851177  M1M2_CDNS_524688791851177_0
timestamp 1707688321
transform 1 0 13682 0 1 4307
box 0 0 384 116
use M1M2_CDNS_524688791851250  M1M2_CDNS_524688791851250_0
timestamp 1707688321
transform 1 0 12411 0 1 3314
box 0 0 448 180
use M2M3_CDNS_524688791851395  M2M3_CDNS_524688791851395_0
timestamp 1707688321
transform 1 0 4626 0 1 4628
box 0 0 1 1
use M2M3_CDNS_524688791851395  M2M3_CDNS_524688791851395_1
timestamp 1707688321
transform 1 0 3728 0 1 4628
box 0 0 1 1
use M2M3_CDNS_524688791851395  M2M3_CDNS_524688791851395_2
timestamp 1707688321
transform 1 0 566 0 1 4628
box 0 0 1 1
use M2M3_CDNS_524688791851396  M2M3_CDNS_524688791851396_0
timestamp 1707688321
transform 1 0 8046 0 1 4628
box -5 0 301 474
use M2M3_CDNS_524688791851396  M2M3_CDNS_524688791851396_1
timestamp 1707688321
transform 1 0 6995 0 1 4628
box -5 0 301 474
use sky130_fd_io__sio_obpredrvr  sky130_fd_io__sio_obpredrvr_0
timestamp 1707688321
transform 1 0 0 0 1 5286
box -185 10 15401 5184
use sky130_fd_io__sio_octl_tsg4  sky130_fd_io__sio_octl_tsg4_0
timestamp 1707688321
transform 1 0 0 0 1 2446
box -84 -146 16041 3752
use sky130_fd_io__sio_opath_datoe  sky130_fd_io__sio_opath_datoe_0
timestamp 1707688321
transform 1 0 6416 0 1 2425
box -307 -1064 15881 2325
<< labels >>
flabel comment s 5171 2297 5171 2297 0 FreeSans 200 0 0 0 hld_i_h_n
flabel metal1 s 5404 3236 5438 3278 3 FreeSans 300 0 0 0 hld_i_vpwr
port 4 nsew
flabel metal1 s 21817 3309 21857 3511 3 FreeSans 300 180 0 0 vgnd
port 2 nsew
flabel metal1 s 16041 3309 16081 3511 3 FreeSans 300 0 0 0 vgnd
port 2 nsew
flabel metal1 s 6237 3309 6277 3511 3 FreeSans 300 180 0 0 vgnd
port 2 nsew
flabel metal1 s 22257 1842 22297 2044 3 FreeSans 300 180 0 0 vcc_io
port 3 nsew
flabel metal1 s 16145 1842 16185 2044 3 FreeSans 300 0 0 0 vcc_io
port 3 nsew
flabel metal1 s 6237 4458 6277 4660 3 FreeSans 300 180 0 0 vcc_io
port 3 nsew
flabel metal1 s 16030 4070 16040 4272 7 FreeSans 200 0 0 0 vpwr_ka
port 7 nsew
flabel metal1 s 16023 4300 16040 4430 7 FreeSans 200 0 0 0 vgnd
port 2 nsew
flabel metal1 s 16029 4458 16040 4660 7 FreeSans 200 0 0 0 vcc_io
port 3 nsew
flabel metal1 s -17 4300 0 4430 3 FreeSans 200 0 0 0 vgnd
port 2 nsew
flabel metal1 s 16027 3309 16041 3511 7 FreeSans 200 0 0 0 vgnd
port 2 nsew
flabel metal1 s -2 2518 16 2636 3 FreeSans 200 0 0 0 vpwr
port 8 nsew
flabel metal1 s 12390 4048 12434 4100 7 FreeSans 400 0 0 0 vreg_en_h
port 5 nsew
flabel metal1 s 4071 3667 4105 3701 0 FreeSans 200 0 0 0 vreg_en
port 6 nsew
flabel metal1 s 185 2664 196 2866 3 FreeSans 200 0 0 0 vpwr
port 8 nsew
flabel metal1 s 0 8051 42 8181 3 FreeSans 200 0 0 0 vgnd_io
port 9 nsew
flabel metal1 s 0 3309 14 3511 3 FreeSans 200 0 0 0 vgnd
port 2 nsew
flabel metal1 s -11 4458 0 4660 7 FreeSans 200 0 0 0 vcc_io
port 3 nsew
flabel metal1 s 5902 9219 5943 9265 3 FreeSans 300 0 0 0 pu_h_n<3>
port 11 nsew
flabel metal1 s 4190 9219 4230 9265 3 FreeSans 300 0 0 0 pu_h_n<2>
port 12 nsew
flabel metal1 s 10098 9375 10138 9421 3 FreeSans 300 0 0 0 pu_h_n<1>
port 13 nsew
flabel metal1 s 7668 9299 7708 9345 3 FreeSans 300 0 0 0 pu_h_n<0>
port 14 nsew
flabel metal1 s 9535 7230 9575 7271 0 FreeSans 200 0 0 0 pd_h<2>
port 15 nsew
flabel metal1 s 9102 9417 9148 9463 3 FreeSans 300 0 0 0 pd_h<1>
port 16 nsew
flabel metal1 s 7872 9423 7906 9457 5 FreeSans 200 0 0 0 pd_h<0>
port 17 nsew
flabel metal1 s 8956 2450 8989 2483 0 FreeSans 200 0 0 0 oe_n
port 19 nsew
flabel metal1 s 13703 9455 13742 9491 0 FreeSans 200 0 0 0 pd_h<4>
port 18 nsew
flabel metal1 s 4153 4697 4193 4737 3 FreeSans 400 0 0 0 od_h
port 20 nsew
flabel metal1 s 4972 2286 5009 2320 0 FreeSans 200 0 0 0 hld_i_h_n
port 21 nsew
flabel metal1 s 349 4850 380 4883 0 FreeSans 400 0 0 0 dm_h_n<2>
port 22 nsew
flabel metal1 s 223 5946 257 5982 3 FreeSans 400 0 0 0 dm_h_n<1>
port 23 nsew
flabel metal1 s 563 5756 597 5790 0 FreeSans 400 0 0 0 dm_h_n<0>
port 24 nsew
flabel metal1 s 3400 4824 3434 4858 0 FreeSans 400 0 0 0 dm_h<2>
port 25 nsew
flabel metal1 s 2868 5841 2903 5876 3 FreeSans 400 0 0 0 dm_h<1>
port 26 nsew
flabel metal1 s 2389 6066 2419 6096 0 FreeSans 400 0 0 0 dm_h<0>
port 27 nsew
flabel metal1 s 10128 2450 10162 2484 0 FreeSans 400 0 0 0 din
port 28 nsew
flabel metal1 s 1547 4124 1580 4167 0 FreeSans 200 0 0 0 slow_h_n
port 29 nsew
flabel metal1 s 99 3667 133 3701 0 FreeSans 400 0 0 0 slow
port 10 nsew
flabel locali s 11576 2385 11616 2431 7 FreeSans 300 0 0 0 od_h
port 20 nsew
flabel locali s 11424 6001 11458 6050 0 FreeSans 200 0 0 0 puen_h<2>
port 30 nsew
flabel locali s 14553 5946 14587 5989 0 FreeSans 200 0 0 0 oe_hs_h
port 31 nsew
flabel locali s 8232 2385 8273 2431 3 FreeSans 300 0 0 0 hld_i_ovr_h
port 32 nsew
flabel locali s 7511 2385 7552 2431 3 FreeSans 300 0 0 0 od_h
port 20 nsew
flabel metal2 s 12545 2303 12863 2335 0 FreeSans 200 0 0 0 vgnd
port 2 nsew
flabel metal2 s 1391 4741 1391 4741 0 FreeSans 200 0 0 0 slow_h
flabel metal2 s 7278 5367 7278 5367 3 FreeSans 300 0 0 0 puen_h<1>
flabel metal2 s 5529 6205 5529 6205 0 FreeSans 200 0 0 0 puen_h<0>
flabel metal2 s 10060 6204 10060 6204 0 FreeSans 200 0 0 0 pden_h_n<1>
flabel metal2 s 10357 5823 10357 5823 0 FreeSans 200 0 0 0 pden_h_n<0>
flabel metal2 s 12163 6257 12163 6257 0 FreeSans 200 0 0 0 drvlo_h_n
flabel metal2 s 15991 3191 16025 3225 0 FreeSans 200 0 0 0 vgnd
port 2 nsew
flabel metal2 s 10324 8909 10382 8961 3 FreeSans 300 0 0 0 pd_h<3>
port 33 nsew
flabel metal2 s 6875 8821 6927 8873 3 FreeSans 200 0 0 0 drvhi_h
port 34 nsew
<< properties >>
string GDS_END 88116650
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 88082900
string path 204.475 238.675 204.475 241.875 
<< end >>
