magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< dnwell >>
rect 1900 28993 7692 29425
rect 4958 1683 7599 16518
<< nwell >>
rect 1820 29073 7772 29345
rect 4878 16312 7679 16598
rect 4878 2736 5164 16312
rect 4878 1889 5234 2736
rect 7393 2735 7679 16312
rect 7348 1889 7679 2735
rect 4878 1603 7679 1889
<< pwell >>
rect 299 1 1745 40001
rect 7854 1 9300 40001
<< psubdiff >>
rect 325 39951 1719 39975
rect 359 39917 461 39951
rect 495 39917 597 39951
rect 631 39917 733 39951
rect 767 39917 869 39951
rect 903 39917 1005 39951
rect 1039 39917 1141 39951
rect 1175 39917 1277 39951
rect 1311 39917 1413 39951
rect 1447 39917 1549 39951
rect 1583 39917 1685 39951
rect 325 39815 1719 39917
rect 359 39781 461 39815
rect 495 39781 597 39815
rect 631 39781 733 39815
rect 767 39781 869 39815
rect 903 39781 1005 39815
rect 1039 39781 1141 39815
rect 1175 39781 1277 39815
rect 1311 39781 1413 39815
rect 1447 39781 1549 39815
rect 1583 39781 1685 39815
rect 325 39679 1719 39781
rect 359 39645 461 39679
rect 495 39645 597 39679
rect 631 39645 733 39679
rect 767 39645 869 39679
rect 903 39645 1005 39679
rect 1039 39645 1141 39679
rect 1175 39645 1277 39679
rect 1311 39645 1413 39679
rect 1447 39645 1549 39679
rect 1583 39645 1685 39679
rect 325 39543 1719 39645
rect 359 39509 461 39543
rect 495 39509 597 39543
rect 631 39509 733 39543
rect 767 39509 869 39543
rect 903 39509 1005 39543
rect 1039 39509 1141 39543
rect 1175 39509 1277 39543
rect 1311 39509 1413 39543
rect 1447 39509 1549 39543
rect 1583 39509 1685 39543
rect 325 39407 1719 39509
rect 359 39373 461 39407
rect 495 39373 597 39407
rect 631 39373 733 39407
rect 767 39373 869 39407
rect 903 39373 1005 39407
rect 1039 39373 1141 39407
rect 1175 39373 1277 39407
rect 1311 39373 1413 39407
rect 1447 39373 1549 39407
rect 1583 39373 1685 39407
rect 325 39271 1719 39373
rect 359 39237 461 39271
rect 495 39237 597 39271
rect 631 39237 733 39271
rect 767 39237 869 39271
rect 903 39237 1005 39271
rect 1039 39237 1141 39271
rect 1175 39237 1277 39271
rect 1311 39237 1413 39271
rect 1447 39237 1549 39271
rect 1583 39237 1685 39271
rect 325 39135 1719 39237
rect 359 39101 461 39135
rect 495 39101 597 39135
rect 631 39101 733 39135
rect 767 39101 869 39135
rect 903 39101 1005 39135
rect 1039 39101 1141 39135
rect 1175 39101 1277 39135
rect 1311 39101 1413 39135
rect 1447 39101 1549 39135
rect 1583 39101 1685 39135
rect 325 38999 1719 39101
rect 359 38965 461 38999
rect 495 38965 597 38999
rect 631 38965 733 38999
rect 767 38965 869 38999
rect 903 38965 1005 38999
rect 1039 38965 1141 38999
rect 1175 38965 1277 38999
rect 1311 38965 1413 38999
rect 1447 38965 1549 38999
rect 1583 38965 1685 38999
rect 325 38863 1719 38965
rect 359 38829 461 38863
rect 495 38829 597 38863
rect 631 38829 733 38863
rect 767 38829 869 38863
rect 903 38829 1005 38863
rect 1039 38829 1141 38863
rect 1175 38829 1277 38863
rect 1311 38829 1413 38863
rect 1447 38829 1549 38863
rect 1583 38829 1685 38863
rect 325 38727 1719 38829
rect 359 38693 461 38727
rect 495 38693 597 38727
rect 631 38693 733 38727
rect 767 38693 869 38727
rect 903 38693 1005 38727
rect 1039 38693 1141 38727
rect 1175 38693 1277 38727
rect 1311 38693 1413 38727
rect 1447 38693 1549 38727
rect 1583 38693 1685 38727
rect 325 38591 1719 38693
rect 359 38557 461 38591
rect 495 38557 597 38591
rect 631 38557 733 38591
rect 767 38557 869 38591
rect 903 38557 1005 38591
rect 1039 38557 1141 38591
rect 1175 38557 1277 38591
rect 1311 38557 1413 38591
rect 1447 38557 1549 38591
rect 1583 38557 1685 38591
rect 325 38455 1719 38557
rect 359 38421 461 38455
rect 495 38421 597 38455
rect 631 38421 733 38455
rect 767 38421 869 38455
rect 903 38421 1005 38455
rect 1039 38421 1141 38455
rect 1175 38421 1277 38455
rect 1311 38421 1413 38455
rect 1447 38421 1549 38455
rect 1583 38421 1685 38455
rect 325 38319 1719 38421
rect 359 38285 461 38319
rect 495 38285 597 38319
rect 631 38285 733 38319
rect 767 38285 869 38319
rect 903 38285 1005 38319
rect 1039 38285 1141 38319
rect 1175 38285 1277 38319
rect 1311 38285 1413 38319
rect 1447 38285 1549 38319
rect 1583 38285 1685 38319
rect 325 38183 1719 38285
rect 359 38149 461 38183
rect 495 38149 597 38183
rect 631 38149 733 38183
rect 767 38149 869 38183
rect 903 38149 1005 38183
rect 1039 38149 1141 38183
rect 1175 38149 1277 38183
rect 1311 38149 1413 38183
rect 1447 38149 1549 38183
rect 1583 38149 1685 38183
rect 325 38047 1719 38149
rect 359 38013 461 38047
rect 495 38013 597 38047
rect 631 38013 733 38047
rect 767 38013 869 38047
rect 903 38013 1005 38047
rect 1039 38013 1141 38047
rect 1175 38013 1277 38047
rect 1311 38013 1413 38047
rect 1447 38013 1549 38047
rect 1583 38013 1685 38047
rect 325 37911 1719 38013
rect 359 37877 461 37911
rect 495 37877 597 37911
rect 631 37877 733 37911
rect 767 37877 869 37911
rect 903 37877 1005 37911
rect 1039 37877 1141 37911
rect 1175 37877 1277 37911
rect 1311 37877 1413 37911
rect 1447 37877 1549 37911
rect 1583 37877 1685 37911
rect 325 37775 1719 37877
rect 359 37741 461 37775
rect 495 37741 597 37775
rect 631 37741 733 37775
rect 767 37741 869 37775
rect 903 37741 1005 37775
rect 1039 37741 1141 37775
rect 1175 37741 1277 37775
rect 1311 37741 1413 37775
rect 1447 37741 1549 37775
rect 1583 37741 1685 37775
rect 325 37639 1719 37741
rect 359 37605 461 37639
rect 495 37605 597 37639
rect 631 37605 733 37639
rect 767 37605 869 37639
rect 903 37605 1005 37639
rect 1039 37605 1141 37639
rect 1175 37605 1277 37639
rect 1311 37605 1413 37639
rect 1447 37605 1549 37639
rect 1583 37605 1685 37639
rect 325 37503 1719 37605
rect 359 37469 461 37503
rect 495 37469 597 37503
rect 631 37469 733 37503
rect 767 37469 869 37503
rect 903 37469 1005 37503
rect 1039 37469 1141 37503
rect 1175 37469 1277 37503
rect 1311 37469 1413 37503
rect 1447 37469 1549 37503
rect 1583 37469 1685 37503
rect 325 37367 1719 37469
rect 359 37333 461 37367
rect 495 37333 597 37367
rect 631 37333 733 37367
rect 767 37333 869 37367
rect 903 37333 1005 37367
rect 1039 37333 1141 37367
rect 1175 37333 1277 37367
rect 1311 37333 1413 37367
rect 1447 37333 1549 37367
rect 1583 37333 1685 37367
rect 325 37231 1719 37333
rect 359 37197 461 37231
rect 495 37197 597 37231
rect 631 37197 733 37231
rect 767 37197 869 37231
rect 903 37197 1005 37231
rect 1039 37197 1141 37231
rect 1175 37197 1277 37231
rect 1311 37197 1413 37231
rect 1447 37197 1549 37231
rect 1583 37197 1685 37231
rect 325 37095 1719 37197
rect 359 37061 461 37095
rect 495 37061 597 37095
rect 631 37061 733 37095
rect 767 37061 869 37095
rect 903 37061 1005 37095
rect 1039 37061 1141 37095
rect 1175 37061 1277 37095
rect 1311 37061 1413 37095
rect 1447 37061 1549 37095
rect 1583 37061 1685 37095
rect 325 36959 1719 37061
rect 359 36925 461 36959
rect 495 36925 597 36959
rect 631 36925 733 36959
rect 767 36925 869 36959
rect 903 36925 1005 36959
rect 1039 36925 1141 36959
rect 1175 36925 1277 36959
rect 1311 36925 1413 36959
rect 1447 36925 1549 36959
rect 1583 36925 1685 36959
rect 325 36823 1719 36925
rect 359 36789 461 36823
rect 495 36789 597 36823
rect 631 36789 733 36823
rect 767 36789 869 36823
rect 903 36789 1005 36823
rect 1039 36789 1141 36823
rect 1175 36789 1277 36823
rect 1311 36789 1413 36823
rect 1447 36789 1549 36823
rect 1583 36789 1685 36823
rect 325 36687 1719 36789
rect 359 36653 461 36687
rect 495 36653 597 36687
rect 631 36653 733 36687
rect 767 36653 869 36687
rect 903 36653 1005 36687
rect 1039 36653 1141 36687
rect 1175 36653 1277 36687
rect 1311 36653 1413 36687
rect 1447 36653 1549 36687
rect 1583 36653 1685 36687
rect 325 36551 1719 36653
rect 359 36517 461 36551
rect 495 36517 597 36551
rect 631 36517 733 36551
rect 767 36517 869 36551
rect 903 36517 1005 36551
rect 1039 36517 1141 36551
rect 1175 36517 1277 36551
rect 1311 36517 1413 36551
rect 1447 36517 1549 36551
rect 1583 36517 1685 36551
rect 325 36415 1719 36517
rect 359 36381 461 36415
rect 495 36381 597 36415
rect 631 36381 733 36415
rect 767 36381 869 36415
rect 903 36381 1005 36415
rect 1039 36381 1141 36415
rect 1175 36381 1277 36415
rect 1311 36381 1413 36415
rect 1447 36381 1549 36415
rect 1583 36381 1685 36415
rect 325 36279 1719 36381
rect 359 36245 461 36279
rect 495 36245 597 36279
rect 631 36245 733 36279
rect 767 36245 869 36279
rect 903 36245 1005 36279
rect 1039 36245 1141 36279
rect 1175 36245 1277 36279
rect 1311 36245 1413 36279
rect 1447 36245 1549 36279
rect 1583 36245 1685 36279
rect 325 36143 1719 36245
rect 359 36109 461 36143
rect 495 36109 597 36143
rect 631 36109 733 36143
rect 767 36109 869 36143
rect 903 36109 1005 36143
rect 1039 36109 1141 36143
rect 1175 36109 1277 36143
rect 1311 36109 1413 36143
rect 1447 36109 1549 36143
rect 1583 36109 1685 36143
rect 325 36007 1719 36109
rect 359 35973 461 36007
rect 495 35973 597 36007
rect 631 35973 733 36007
rect 767 35973 869 36007
rect 903 35973 1005 36007
rect 1039 35973 1141 36007
rect 1175 35973 1277 36007
rect 1311 35973 1413 36007
rect 1447 35973 1549 36007
rect 1583 35973 1685 36007
rect 325 35871 1719 35973
rect 359 35837 461 35871
rect 495 35837 597 35871
rect 631 35837 733 35871
rect 767 35837 869 35871
rect 903 35837 1005 35871
rect 1039 35837 1141 35871
rect 1175 35837 1277 35871
rect 1311 35837 1413 35871
rect 1447 35837 1549 35871
rect 1583 35837 1685 35871
rect 325 35735 1719 35837
rect 359 35701 461 35735
rect 495 35701 597 35735
rect 631 35701 733 35735
rect 767 35701 869 35735
rect 903 35701 1005 35735
rect 1039 35701 1141 35735
rect 1175 35701 1277 35735
rect 1311 35701 1413 35735
rect 1447 35701 1549 35735
rect 1583 35701 1685 35735
rect 325 35599 1719 35701
rect 359 35565 461 35599
rect 495 35565 597 35599
rect 631 35565 733 35599
rect 767 35565 869 35599
rect 903 35565 1005 35599
rect 1039 35565 1141 35599
rect 1175 35565 1277 35599
rect 1311 35565 1413 35599
rect 1447 35565 1549 35599
rect 1583 35565 1685 35599
rect 325 35463 1719 35565
rect 359 35429 461 35463
rect 495 35429 597 35463
rect 631 35429 733 35463
rect 767 35429 869 35463
rect 903 35429 1005 35463
rect 1039 35429 1141 35463
rect 1175 35429 1277 35463
rect 1311 35429 1413 35463
rect 1447 35429 1549 35463
rect 1583 35429 1685 35463
rect 325 35327 1719 35429
rect 359 35293 461 35327
rect 495 35293 597 35327
rect 631 35293 733 35327
rect 767 35293 869 35327
rect 903 35293 1005 35327
rect 1039 35293 1141 35327
rect 1175 35293 1277 35327
rect 1311 35293 1413 35327
rect 1447 35293 1549 35327
rect 1583 35293 1685 35327
rect 325 35191 1719 35293
rect 359 35157 461 35191
rect 495 35157 597 35191
rect 631 35157 733 35191
rect 767 35157 869 35191
rect 903 35157 1005 35191
rect 1039 35157 1141 35191
rect 1175 35157 1277 35191
rect 1311 35157 1413 35191
rect 1447 35157 1549 35191
rect 1583 35157 1685 35191
rect 325 35055 1719 35157
rect 359 35021 461 35055
rect 495 35021 597 35055
rect 631 35021 733 35055
rect 767 35021 869 35055
rect 903 35021 1005 35055
rect 1039 35021 1141 35055
rect 1175 35021 1277 35055
rect 1311 35021 1413 35055
rect 1447 35021 1549 35055
rect 1583 35021 1685 35055
rect 325 34919 1719 35021
rect 359 34885 461 34919
rect 495 34885 597 34919
rect 631 34885 733 34919
rect 767 34885 869 34919
rect 903 34885 1005 34919
rect 1039 34885 1141 34919
rect 1175 34885 1277 34919
rect 1311 34885 1413 34919
rect 1447 34885 1549 34919
rect 1583 34885 1685 34919
rect 325 34783 1719 34885
rect 359 34749 461 34783
rect 495 34749 597 34783
rect 631 34749 733 34783
rect 767 34749 869 34783
rect 903 34749 1005 34783
rect 1039 34749 1141 34783
rect 1175 34749 1277 34783
rect 1311 34749 1413 34783
rect 1447 34749 1549 34783
rect 1583 34749 1685 34783
rect 325 34647 1719 34749
rect 359 34613 461 34647
rect 495 34613 597 34647
rect 631 34613 733 34647
rect 767 34613 869 34647
rect 903 34613 1005 34647
rect 1039 34613 1141 34647
rect 1175 34613 1277 34647
rect 1311 34613 1413 34647
rect 1447 34613 1549 34647
rect 1583 34613 1685 34647
rect 325 34511 1719 34613
rect 359 34477 461 34511
rect 495 34477 597 34511
rect 631 34477 733 34511
rect 767 34477 869 34511
rect 903 34477 1005 34511
rect 1039 34477 1141 34511
rect 1175 34477 1277 34511
rect 1311 34477 1413 34511
rect 1447 34477 1549 34511
rect 1583 34477 1685 34511
rect 325 34375 1719 34477
rect 359 34341 461 34375
rect 495 34341 597 34375
rect 631 34341 733 34375
rect 767 34341 869 34375
rect 903 34341 1005 34375
rect 1039 34341 1141 34375
rect 1175 34341 1277 34375
rect 1311 34341 1413 34375
rect 1447 34341 1549 34375
rect 1583 34341 1685 34375
rect 325 34239 1719 34341
rect 359 34205 461 34239
rect 495 34205 597 34239
rect 631 34205 733 34239
rect 767 34205 869 34239
rect 903 34205 1005 34239
rect 1039 34205 1141 34239
rect 1175 34205 1277 34239
rect 1311 34205 1413 34239
rect 1447 34205 1549 34239
rect 1583 34205 1685 34239
rect 325 34103 1719 34205
rect 359 34069 461 34103
rect 495 34069 597 34103
rect 631 34069 733 34103
rect 767 34069 869 34103
rect 903 34069 1005 34103
rect 1039 34069 1141 34103
rect 1175 34069 1277 34103
rect 1311 34069 1413 34103
rect 1447 34069 1549 34103
rect 1583 34069 1685 34103
rect 325 33967 1719 34069
rect 359 33933 461 33967
rect 495 33933 597 33967
rect 631 33933 733 33967
rect 767 33933 869 33967
rect 903 33933 1005 33967
rect 1039 33933 1141 33967
rect 1175 33933 1277 33967
rect 1311 33933 1413 33967
rect 1447 33933 1549 33967
rect 1583 33933 1685 33967
rect 325 33831 1719 33933
rect 359 33797 461 33831
rect 495 33797 597 33831
rect 631 33797 733 33831
rect 767 33797 869 33831
rect 903 33797 1005 33831
rect 1039 33797 1141 33831
rect 1175 33797 1277 33831
rect 1311 33797 1413 33831
rect 1447 33797 1549 33831
rect 1583 33797 1685 33831
rect 325 33695 1719 33797
rect 359 33661 461 33695
rect 495 33661 597 33695
rect 631 33661 733 33695
rect 767 33661 869 33695
rect 903 33661 1005 33695
rect 1039 33661 1141 33695
rect 1175 33661 1277 33695
rect 1311 33661 1413 33695
rect 1447 33661 1549 33695
rect 1583 33661 1685 33695
rect 325 33559 1719 33661
rect 359 33525 461 33559
rect 495 33525 597 33559
rect 631 33525 733 33559
rect 767 33525 869 33559
rect 903 33525 1005 33559
rect 1039 33525 1141 33559
rect 1175 33525 1277 33559
rect 1311 33525 1413 33559
rect 1447 33525 1549 33559
rect 1583 33525 1685 33559
rect 325 33423 1719 33525
rect 359 33389 461 33423
rect 495 33389 597 33423
rect 631 33389 733 33423
rect 767 33389 869 33423
rect 903 33389 1005 33423
rect 1039 33389 1141 33423
rect 1175 33389 1277 33423
rect 1311 33389 1413 33423
rect 1447 33389 1549 33423
rect 1583 33389 1685 33423
rect 325 33287 1719 33389
rect 359 33253 461 33287
rect 495 33253 597 33287
rect 631 33253 733 33287
rect 767 33253 869 33287
rect 903 33253 1005 33287
rect 1039 33253 1141 33287
rect 1175 33253 1277 33287
rect 1311 33253 1413 33287
rect 1447 33253 1549 33287
rect 1583 33253 1685 33287
rect 325 33151 1719 33253
rect 359 33117 461 33151
rect 495 33117 597 33151
rect 631 33117 733 33151
rect 767 33117 869 33151
rect 903 33117 1005 33151
rect 1039 33117 1141 33151
rect 1175 33117 1277 33151
rect 1311 33117 1413 33151
rect 1447 33117 1549 33151
rect 1583 33117 1685 33151
rect 325 33015 1719 33117
rect 359 32981 461 33015
rect 495 32981 597 33015
rect 631 32981 733 33015
rect 767 32981 869 33015
rect 903 32981 1005 33015
rect 1039 32981 1141 33015
rect 1175 32981 1277 33015
rect 1311 32981 1413 33015
rect 1447 32981 1549 33015
rect 1583 32981 1685 33015
rect 325 32879 1719 32981
rect 359 32845 461 32879
rect 495 32845 597 32879
rect 631 32845 733 32879
rect 767 32845 869 32879
rect 903 32845 1005 32879
rect 1039 32845 1141 32879
rect 1175 32845 1277 32879
rect 1311 32845 1413 32879
rect 1447 32845 1549 32879
rect 1583 32845 1685 32879
rect 325 32743 1719 32845
rect 359 32709 461 32743
rect 495 32709 597 32743
rect 631 32709 733 32743
rect 767 32709 869 32743
rect 903 32709 1005 32743
rect 1039 32709 1141 32743
rect 1175 32709 1277 32743
rect 1311 32709 1413 32743
rect 1447 32709 1549 32743
rect 1583 32709 1685 32743
rect 325 32607 1719 32709
rect 359 32573 461 32607
rect 495 32573 597 32607
rect 631 32573 733 32607
rect 767 32573 869 32607
rect 903 32573 1005 32607
rect 1039 32573 1141 32607
rect 1175 32573 1277 32607
rect 1311 32573 1413 32607
rect 1447 32573 1549 32607
rect 1583 32573 1685 32607
rect 325 32471 1719 32573
rect 359 32437 461 32471
rect 495 32437 597 32471
rect 631 32437 733 32471
rect 767 32437 869 32471
rect 903 32437 1005 32471
rect 1039 32437 1141 32471
rect 1175 32437 1277 32471
rect 1311 32437 1413 32471
rect 1447 32437 1549 32471
rect 1583 32437 1685 32471
rect 325 32335 1719 32437
rect 359 32301 461 32335
rect 495 32301 597 32335
rect 631 32301 733 32335
rect 767 32301 869 32335
rect 903 32301 1005 32335
rect 1039 32301 1141 32335
rect 1175 32301 1277 32335
rect 1311 32301 1413 32335
rect 1447 32301 1549 32335
rect 1583 32301 1685 32335
rect 325 32199 1719 32301
rect 359 32165 461 32199
rect 495 32165 597 32199
rect 631 32165 733 32199
rect 767 32165 869 32199
rect 903 32165 1005 32199
rect 1039 32165 1141 32199
rect 1175 32165 1277 32199
rect 1311 32165 1413 32199
rect 1447 32165 1549 32199
rect 1583 32165 1685 32199
rect 325 32063 1719 32165
rect 359 32029 461 32063
rect 495 32029 597 32063
rect 631 32029 733 32063
rect 767 32029 869 32063
rect 903 32029 1005 32063
rect 1039 32029 1141 32063
rect 1175 32029 1277 32063
rect 1311 32029 1413 32063
rect 1447 32029 1549 32063
rect 1583 32029 1685 32063
rect 325 31927 1719 32029
rect 359 31893 461 31927
rect 495 31893 597 31927
rect 631 31893 733 31927
rect 767 31893 869 31927
rect 903 31893 1005 31927
rect 1039 31893 1141 31927
rect 1175 31893 1277 31927
rect 1311 31893 1413 31927
rect 1447 31893 1549 31927
rect 1583 31893 1685 31927
rect 325 31791 1719 31893
rect 359 31757 461 31791
rect 495 31757 597 31791
rect 631 31757 733 31791
rect 767 31757 869 31791
rect 903 31757 1005 31791
rect 1039 31757 1141 31791
rect 1175 31757 1277 31791
rect 1311 31757 1413 31791
rect 1447 31757 1549 31791
rect 1583 31757 1685 31791
rect 325 31655 1719 31757
rect 359 31621 461 31655
rect 495 31621 597 31655
rect 631 31621 733 31655
rect 767 31621 869 31655
rect 903 31621 1005 31655
rect 1039 31621 1141 31655
rect 1175 31621 1277 31655
rect 1311 31621 1413 31655
rect 1447 31621 1549 31655
rect 1583 31621 1685 31655
rect 325 31519 1719 31621
rect 359 31485 461 31519
rect 495 31485 597 31519
rect 631 31485 733 31519
rect 767 31485 869 31519
rect 903 31485 1005 31519
rect 1039 31485 1141 31519
rect 1175 31485 1277 31519
rect 1311 31485 1413 31519
rect 1447 31485 1549 31519
rect 1583 31485 1685 31519
rect 325 31383 1719 31485
rect 359 31349 461 31383
rect 495 31349 597 31383
rect 631 31349 733 31383
rect 767 31349 869 31383
rect 903 31349 1005 31383
rect 1039 31349 1141 31383
rect 1175 31349 1277 31383
rect 1311 31349 1413 31383
rect 1447 31349 1549 31383
rect 1583 31349 1685 31383
rect 325 31247 1719 31349
rect 359 31213 461 31247
rect 495 31213 597 31247
rect 631 31213 733 31247
rect 767 31213 869 31247
rect 903 31213 1005 31247
rect 1039 31213 1141 31247
rect 1175 31213 1277 31247
rect 1311 31213 1413 31247
rect 1447 31213 1549 31247
rect 1583 31213 1685 31247
rect 325 31111 1719 31213
rect 359 31077 461 31111
rect 495 31077 597 31111
rect 631 31077 733 31111
rect 767 31077 869 31111
rect 903 31077 1005 31111
rect 1039 31077 1141 31111
rect 1175 31077 1277 31111
rect 1311 31077 1413 31111
rect 1447 31077 1549 31111
rect 1583 31077 1685 31111
rect 325 30975 1719 31077
rect 359 30941 461 30975
rect 495 30941 597 30975
rect 631 30941 733 30975
rect 767 30941 869 30975
rect 903 30941 1005 30975
rect 1039 30941 1141 30975
rect 1175 30941 1277 30975
rect 1311 30941 1413 30975
rect 1447 30941 1549 30975
rect 1583 30941 1685 30975
rect 325 30839 1719 30941
rect 359 30805 461 30839
rect 495 30805 597 30839
rect 631 30805 733 30839
rect 767 30805 869 30839
rect 903 30805 1005 30839
rect 1039 30805 1141 30839
rect 1175 30805 1277 30839
rect 1311 30805 1413 30839
rect 1447 30805 1549 30839
rect 1583 30805 1685 30839
rect 325 30703 1719 30805
rect 359 30669 461 30703
rect 495 30669 597 30703
rect 631 30669 733 30703
rect 767 30669 869 30703
rect 903 30669 1005 30703
rect 1039 30669 1141 30703
rect 1175 30669 1277 30703
rect 1311 30669 1413 30703
rect 1447 30669 1549 30703
rect 1583 30669 1685 30703
rect 325 30567 1719 30669
rect 359 30533 461 30567
rect 495 30533 597 30567
rect 631 30533 733 30567
rect 767 30533 869 30567
rect 903 30533 1005 30567
rect 1039 30533 1141 30567
rect 1175 30533 1277 30567
rect 1311 30533 1413 30567
rect 1447 30533 1549 30567
rect 1583 30533 1685 30567
rect 325 30431 1719 30533
rect 359 30397 461 30431
rect 495 30397 597 30431
rect 631 30397 733 30431
rect 767 30397 869 30431
rect 903 30397 1005 30431
rect 1039 30397 1141 30431
rect 1175 30397 1277 30431
rect 1311 30397 1413 30431
rect 1447 30397 1549 30431
rect 1583 30397 1685 30431
rect 325 30295 1719 30397
rect 359 30261 461 30295
rect 495 30261 597 30295
rect 631 30261 733 30295
rect 767 30261 869 30295
rect 903 30261 1005 30295
rect 1039 30261 1141 30295
rect 1175 30261 1277 30295
rect 1311 30261 1413 30295
rect 1447 30261 1549 30295
rect 1583 30261 1685 30295
rect 325 30159 1719 30261
rect 359 30125 461 30159
rect 495 30125 597 30159
rect 631 30125 733 30159
rect 767 30125 869 30159
rect 903 30125 1005 30159
rect 1039 30125 1141 30159
rect 1175 30125 1277 30159
rect 1311 30125 1413 30159
rect 1447 30125 1549 30159
rect 1583 30125 1685 30159
rect 325 30023 1719 30125
rect 359 29989 461 30023
rect 495 29989 597 30023
rect 631 29989 733 30023
rect 767 29989 869 30023
rect 903 29989 1005 30023
rect 1039 29989 1141 30023
rect 1175 29989 1277 30023
rect 1311 29989 1413 30023
rect 1447 29989 1549 30023
rect 1583 29989 1685 30023
rect 325 29887 1719 29989
rect 359 29853 461 29887
rect 495 29853 597 29887
rect 631 29853 733 29887
rect 767 29853 869 29887
rect 903 29853 1005 29887
rect 1039 29853 1141 29887
rect 1175 29853 1277 29887
rect 1311 29853 1413 29887
rect 1447 29853 1549 29887
rect 1583 29853 1685 29887
rect 325 29751 1719 29853
rect 359 29717 461 29751
rect 495 29717 597 29751
rect 631 29717 733 29751
rect 767 29717 869 29751
rect 903 29717 1005 29751
rect 1039 29717 1141 29751
rect 1175 29717 1277 29751
rect 1311 29717 1413 29751
rect 1447 29717 1549 29751
rect 1583 29717 1685 29751
rect 325 29615 1719 29717
rect 359 29581 461 29615
rect 495 29581 597 29615
rect 631 29581 733 29615
rect 767 29581 869 29615
rect 903 29581 1005 29615
rect 1039 29581 1141 29615
rect 1175 29581 1277 29615
rect 1311 29581 1413 29615
rect 1447 29581 1549 29615
rect 1583 29581 1685 29615
rect 325 29479 1719 29581
rect 359 29445 461 29479
rect 495 29445 597 29479
rect 631 29445 733 29479
rect 767 29445 869 29479
rect 903 29445 1005 29479
rect 1039 29445 1141 29479
rect 1175 29445 1277 29479
rect 1311 29445 1413 29479
rect 1447 29445 1549 29479
rect 1583 29445 1685 29479
rect 325 29343 1719 29445
rect 359 29309 461 29343
rect 495 29309 597 29343
rect 631 29309 733 29343
rect 767 29309 869 29343
rect 903 29309 1005 29343
rect 1039 29309 1141 29343
rect 1175 29309 1277 29343
rect 1311 29309 1413 29343
rect 1447 29309 1549 29343
rect 1583 29309 1685 29343
rect 325 29207 1719 29309
rect 359 29173 461 29207
rect 495 29173 597 29207
rect 631 29173 733 29207
rect 767 29173 869 29207
rect 903 29173 1005 29207
rect 1039 29173 1141 29207
rect 1175 29173 1277 29207
rect 1311 29173 1413 29207
rect 1447 29173 1549 29207
rect 1583 29173 1685 29207
rect 325 29071 1719 29173
rect 359 29037 461 29071
rect 495 29037 597 29071
rect 631 29037 733 29071
rect 767 29037 869 29071
rect 903 29037 1005 29071
rect 1039 29037 1141 29071
rect 1175 29037 1277 29071
rect 1311 29037 1413 29071
rect 1447 29037 1549 29071
rect 1583 29037 1685 29071
rect 325 28935 1719 29037
rect 359 28901 461 28935
rect 495 28901 597 28935
rect 631 28901 733 28935
rect 767 28901 869 28935
rect 903 28901 1005 28935
rect 1039 28901 1141 28935
rect 1175 28901 1277 28935
rect 1311 28901 1413 28935
rect 1447 28901 1549 28935
rect 1583 28901 1685 28935
rect 325 28799 1719 28901
rect 359 28765 461 28799
rect 495 28765 597 28799
rect 631 28765 733 28799
rect 767 28765 869 28799
rect 903 28765 1005 28799
rect 1039 28765 1141 28799
rect 1175 28765 1277 28799
rect 1311 28765 1413 28799
rect 1447 28765 1549 28799
rect 1583 28765 1685 28799
rect 325 28663 1719 28765
rect 359 28629 461 28663
rect 495 28629 597 28663
rect 631 28629 733 28663
rect 767 28629 869 28663
rect 903 28629 1005 28663
rect 1039 28629 1141 28663
rect 1175 28629 1277 28663
rect 1311 28629 1413 28663
rect 1447 28629 1549 28663
rect 1583 28629 1685 28663
rect 325 28527 1719 28629
rect 359 28493 461 28527
rect 495 28493 597 28527
rect 631 28493 733 28527
rect 767 28493 869 28527
rect 903 28493 1005 28527
rect 1039 28493 1141 28527
rect 1175 28493 1277 28527
rect 1311 28493 1413 28527
rect 1447 28493 1549 28527
rect 1583 28493 1685 28527
rect 325 28391 1719 28493
rect 359 28357 461 28391
rect 495 28357 597 28391
rect 631 28357 733 28391
rect 767 28357 869 28391
rect 903 28357 1005 28391
rect 1039 28357 1141 28391
rect 1175 28357 1277 28391
rect 1311 28357 1413 28391
rect 1447 28357 1549 28391
rect 1583 28357 1685 28391
rect 325 28255 1719 28357
rect 359 28221 461 28255
rect 495 28221 597 28255
rect 631 28221 733 28255
rect 767 28221 869 28255
rect 903 28221 1005 28255
rect 1039 28221 1141 28255
rect 1175 28221 1277 28255
rect 1311 28221 1413 28255
rect 1447 28221 1549 28255
rect 1583 28221 1685 28255
rect 325 28119 1719 28221
rect 359 28085 461 28119
rect 495 28085 597 28119
rect 631 28085 733 28119
rect 767 28085 869 28119
rect 903 28085 1005 28119
rect 1039 28085 1141 28119
rect 1175 28085 1277 28119
rect 1311 28085 1413 28119
rect 1447 28085 1549 28119
rect 1583 28085 1685 28119
rect 325 27983 1719 28085
rect 359 27949 461 27983
rect 495 27949 597 27983
rect 631 27949 733 27983
rect 767 27949 869 27983
rect 903 27949 1005 27983
rect 1039 27949 1141 27983
rect 1175 27949 1277 27983
rect 1311 27949 1413 27983
rect 1447 27949 1549 27983
rect 1583 27949 1685 27983
rect 325 27847 1719 27949
rect 359 27813 461 27847
rect 495 27813 597 27847
rect 631 27813 733 27847
rect 767 27813 869 27847
rect 903 27813 1005 27847
rect 1039 27813 1141 27847
rect 1175 27813 1277 27847
rect 1311 27813 1413 27847
rect 1447 27813 1549 27847
rect 1583 27813 1685 27847
rect 325 27711 1719 27813
rect 359 27677 461 27711
rect 495 27677 597 27711
rect 631 27677 733 27711
rect 767 27677 869 27711
rect 903 27677 1005 27711
rect 1039 27677 1141 27711
rect 1175 27677 1277 27711
rect 1311 27677 1413 27711
rect 1447 27677 1549 27711
rect 1583 27677 1685 27711
rect 325 27575 1719 27677
rect 359 27541 461 27575
rect 495 27541 597 27575
rect 631 27541 733 27575
rect 767 27541 869 27575
rect 903 27541 1005 27575
rect 1039 27541 1141 27575
rect 1175 27541 1277 27575
rect 1311 27541 1413 27575
rect 1447 27541 1549 27575
rect 1583 27541 1685 27575
rect 325 27439 1719 27541
rect 359 27405 461 27439
rect 495 27405 597 27439
rect 631 27405 733 27439
rect 767 27405 869 27439
rect 903 27405 1005 27439
rect 1039 27405 1141 27439
rect 1175 27405 1277 27439
rect 1311 27405 1413 27439
rect 1447 27405 1549 27439
rect 1583 27405 1685 27439
rect 325 27303 1719 27405
rect 359 27269 461 27303
rect 495 27269 597 27303
rect 631 27269 733 27303
rect 767 27269 869 27303
rect 903 27269 1005 27303
rect 1039 27269 1141 27303
rect 1175 27269 1277 27303
rect 1311 27269 1413 27303
rect 1447 27269 1549 27303
rect 1583 27269 1685 27303
rect 325 27167 1719 27269
rect 359 27133 461 27167
rect 495 27133 597 27167
rect 631 27133 733 27167
rect 767 27133 869 27167
rect 903 27133 1005 27167
rect 1039 27133 1141 27167
rect 1175 27133 1277 27167
rect 1311 27133 1413 27167
rect 1447 27133 1549 27167
rect 1583 27133 1685 27167
rect 325 27031 1719 27133
rect 359 26997 461 27031
rect 495 26997 597 27031
rect 631 26997 733 27031
rect 767 26997 869 27031
rect 903 26997 1005 27031
rect 1039 26997 1141 27031
rect 1175 26997 1277 27031
rect 1311 26997 1413 27031
rect 1447 26997 1549 27031
rect 1583 26997 1685 27031
rect 325 26895 1719 26997
rect 359 26861 461 26895
rect 495 26861 597 26895
rect 631 26861 733 26895
rect 767 26861 869 26895
rect 903 26861 1005 26895
rect 1039 26861 1141 26895
rect 1175 26861 1277 26895
rect 1311 26861 1413 26895
rect 1447 26861 1549 26895
rect 1583 26861 1685 26895
rect 325 26759 1719 26861
rect 359 26725 461 26759
rect 495 26725 597 26759
rect 631 26725 733 26759
rect 767 26725 869 26759
rect 903 26725 1005 26759
rect 1039 26725 1141 26759
rect 1175 26725 1277 26759
rect 1311 26725 1413 26759
rect 1447 26725 1549 26759
rect 1583 26725 1685 26759
rect 325 26623 1719 26725
rect 359 26589 461 26623
rect 495 26589 597 26623
rect 631 26589 733 26623
rect 767 26589 869 26623
rect 903 26589 1005 26623
rect 1039 26589 1141 26623
rect 1175 26589 1277 26623
rect 1311 26589 1413 26623
rect 1447 26589 1549 26623
rect 1583 26589 1685 26623
rect 325 26487 1719 26589
rect 359 26453 461 26487
rect 495 26453 597 26487
rect 631 26453 733 26487
rect 767 26453 869 26487
rect 903 26453 1005 26487
rect 1039 26453 1141 26487
rect 1175 26453 1277 26487
rect 1311 26453 1413 26487
rect 1447 26453 1549 26487
rect 1583 26453 1685 26487
rect 325 26351 1719 26453
rect 359 26317 461 26351
rect 495 26317 597 26351
rect 631 26317 733 26351
rect 767 26317 869 26351
rect 903 26317 1005 26351
rect 1039 26317 1141 26351
rect 1175 26317 1277 26351
rect 1311 26317 1413 26351
rect 1447 26317 1549 26351
rect 1583 26317 1685 26351
rect 325 26215 1719 26317
rect 359 26181 461 26215
rect 495 26181 597 26215
rect 631 26181 733 26215
rect 767 26181 869 26215
rect 903 26181 1005 26215
rect 1039 26181 1141 26215
rect 1175 26181 1277 26215
rect 1311 26181 1413 26215
rect 1447 26181 1549 26215
rect 1583 26181 1685 26215
rect 325 26079 1719 26181
rect 359 26045 461 26079
rect 495 26045 597 26079
rect 631 26045 733 26079
rect 767 26045 869 26079
rect 903 26045 1005 26079
rect 1039 26045 1141 26079
rect 1175 26045 1277 26079
rect 1311 26045 1413 26079
rect 1447 26045 1549 26079
rect 1583 26045 1685 26079
rect 325 25943 1719 26045
rect 359 25909 461 25943
rect 495 25909 597 25943
rect 631 25909 733 25943
rect 767 25909 869 25943
rect 903 25909 1005 25943
rect 1039 25909 1141 25943
rect 1175 25909 1277 25943
rect 1311 25909 1413 25943
rect 1447 25909 1549 25943
rect 1583 25909 1685 25943
rect 325 25807 1719 25909
rect 359 25773 461 25807
rect 495 25773 597 25807
rect 631 25773 733 25807
rect 767 25773 869 25807
rect 903 25773 1005 25807
rect 1039 25773 1141 25807
rect 1175 25773 1277 25807
rect 1311 25773 1413 25807
rect 1447 25773 1549 25807
rect 1583 25773 1685 25807
rect 325 25671 1719 25773
rect 359 25637 461 25671
rect 495 25637 597 25671
rect 631 25637 733 25671
rect 767 25637 869 25671
rect 903 25637 1005 25671
rect 1039 25637 1141 25671
rect 1175 25637 1277 25671
rect 1311 25637 1413 25671
rect 1447 25637 1549 25671
rect 1583 25637 1685 25671
rect 325 25535 1719 25637
rect 359 25501 461 25535
rect 495 25501 597 25535
rect 631 25501 733 25535
rect 767 25501 869 25535
rect 903 25501 1005 25535
rect 1039 25501 1141 25535
rect 1175 25501 1277 25535
rect 1311 25501 1413 25535
rect 1447 25501 1549 25535
rect 1583 25501 1685 25535
rect 325 25399 1719 25501
rect 359 25365 461 25399
rect 495 25365 597 25399
rect 631 25365 733 25399
rect 767 25365 869 25399
rect 903 25365 1005 25399
rect 1039 25365 1141 25399
rect 1175 25365 1277 25399
rect 1311 25365 1413 25399
rect 1447 25365 1549 25399
rect 1583 25365 1685 25399
rect 325 25263 1719 25365
rect 359 25229 461 25263
rect 495 25229 597 25263
rect 631 25229 733 25263
rect 767 25229 869 25263
rect 903 25229 1005 25263
rect 1039 25229 1141 25263
rect 1175 25229 1277 25263
rect 1311 25229 1413 25263
rect 1447 25229 1549 25263
rect 1583 25229 1685 25263
rect 325 25127 1719 25229
rect 359 25093 461 25127
rect 495 25093 597 25127
rect 631 25093 733 25127
rect 767 25093 869 25127
rect 903 25093 1005 25127
rect 1039 25093 1141 25127
rect 1175 25093 1277 25127
rect 1311 25093 1413 25127
rect 1447 25093 1549 25127
rect 1583 25093 1685 25127
rect 325 24991 1719 25093
rect 359 24957 461 24991
rect 495 24957 597 24991
rect 631 24957 733 24991
rect 767 24957 869 24991
rect 903 24957 1005 24991
rect 1039 24957 1141 24991
rect 1175 24957 1277 24991
rect 1311 24957 1413 24991
rect 1447 24957 1549 24991
rect 1583 24957 1685 24991
rect 325 24855 1719 24957
rect 359 24821 461 24855
rect 495 24821 597 24855
rect 631 24821 733 24855
rect 767 24821 869 24855
rect 903 24821 1005 24855
rect 1039 24821 1141 24855
rect 1175 24821 1277 24855
rect 1311 24821 1413 24855
rect 1447 24821 1549 24855
rect 1583 24821 1685 24855
rect 325 24719 1719 24821
rect 359 24685 461 24719
rect 495 24685 597 24719
rect 631 24685 733 24719
rect 767 24685 869 24719
rect 903 24685 1005 24719
rect 1039 24685 1141 24719
rect 1175 24685 1277 24719
rect 1311 24685 1413 24719
rect 1447 24685 1549 24719
rect 1583 24685 1685 24719
rect 325 24583 1719 24685
rect 359 24549 461 24583
rect 495 24549 597 24583
rect 631 24549 733 24583
rect 767 24549 869 24583
rect 903 24549 1005 24583
rect 1039 24549 1141 24583
rect 1175 24549 1277 24583
rect 1311 24549 1413 24583
rect 1447 24549 1549 24583
rect 1583 24549 1685 24583
rect 325 24447 1719 24549
rect 359 24413 461 24447
rect 495 24413 597 24447
rect 631 24413 733 24447
rect 767 24413 869 24447
rect 903 24413 1005 24447
rect 1039 24413 1141 24447
rect 1175 24413 1277 24447
rect 1311 24413 1413 24447
rect 1447 24413 1549 24447
rect 1583 24413 1685 24447
rect 325 24311 1719 24413
rect 359 24277 461 24311
rect 495 24277 597 24311
rect 631 24277 733 24311
rect 767 24277 869 24311
rect 903 24277 1005 24311
rect 1039 24277 1141 24311
rect 1175 24277 1277 24311
rect 1311 24277 1413 24311
rect 1447 24277 1549 24311
rect 1583 24277 1685 24311
rect 325 24175 1719 24277
rect 359 24141 461 24175
rect 495 24141 597 24175
rect 631 24141 733 24175
rect 767 24141 869 24175
rect 903 24141 1005 24175
rect 1039 24141 1141 24175
rect 1175 24141 1277 24175
rect 1311 24141 1413 24175
rect 1447 24141 1549 24175
rect 1583 24141 1685 24175
rect 325 24039 1719 24141
rect 359 24005 461 24039
rect 495 24005 597 24039
rect 631 24005 733 24039
rect 767 24005 869 24039
rect 903 24005 1005 24039
rect 1039 24005 1141 24039
rect 1175 24005 1277 24039
rect 1311 24005 1413 24039
rect 1447 24005 1549 24039
rect 1583 24005 1685 24039
rect 325 23903 1719 24005
rect 359 23869 461 23903
rect 495 23869 597 23903
rect 631 23869 733 23903
rect 767 23869 869 23903
rect 903 23869 1005 23903
rect 1039 23869 1141 23903
rect 1175 23869 1277 23903
rect 1311 23869 1413 23903
rect 1447 23869 1549 23903
rect 1583 23869 1685 23903
rect 325 23767 1719 23869
rect 359 23733 461 23767
rect 495 23733 597 23767
rect 631 23733 733 23767
rect 767 23733 869 23767
rect 903 23733 1005 23767
rect 1039 23733 1141 23767
rect 1175 23733 1277 23767
rect 1311 23733 1413 23767
rect 1447 23733 1549 23767
rect 1583 23733 1685 23767
rect 325 23631 1719 23733
rect 359 23597 461 23631
rect 495 23597 597 23631
rect 631 23597 733 23631
rect 767 23597 869 23631
rect 903 23597 1005 23631
rect 1039 23597 1141 23631
rect 1175 23597 1277 23631
rect 1311 23597 1413 23631
rect 1447 23597 1549 23631
rect 1583 23597 1685 23631
rect 325 23495 1719 23597
rect 359 23461 461 23495
rect 495 23461 597 23495
rect 631 23461 733 23495
rect 767 23461 869 23495
rect 903 23461 1005 23495
rect 1039 23461 1141 23495
rect 1175 23461 1277 23495
rect 1311 23461 1413 23495
rect 1447 23461 1549 23495
rect 1583 23461 1685 23495
rect 325 23359 1719 23461
rect 359 23325 461 23359
rect 495 23325 597 23359
rect 631 23325 733 23359
rect 767 23325 869 23359
rect 903 23325 1005 23359
rect 1039 23325 1141 23359
rect 1175 23325 1277 23359
rect 1311 23325 1413 23359
rect 1447 23325 1549 23359
rect 1583 23325 1685 23359
rect 325 23223 1719 23325
rect 359 23189 461 23223
rect 495 23189 597 23223
rect 631 23189 733 23223
rect 767 23189 869 23223
rect 903 23189 1005 23223
rect 1039 23189 1141 23223
rect 1175 23189 1277 23223
rect 1311 23189 1413 23223
rect 1447 23189 1549 23223
rect 1583 23189 1685 23223
rect 325 23087 1719 23189
rect 359 23053 461 23087
rect 495 23053 597 23087
rect 631 23053 733 23087
rect 767 23053 869 23087
rect 903 23053 1005 23087
rect 1039 23053 1141 23087
rect 1175 23053 1277 23087
rect 1311 23053 1413 23087
rect 1447 23053 1549 23087
rect 1583 23053 1685 23087
rect 325 22951 1719 23053
rect 359 22917 461 22951
rect 495 22917 597 22951
rect 631 22917 733 22951
rect 767 22917 869 22951
rect 903 22917 1005 22951
rect 1039 22917 1141 22951
rect 1175 22917 1277 22951
rect 1311 22917 1413 22951
rect 1447 22917 1549 22951
rect 1583 22917 1685 22951
rect 325 22815 1719 22917
rect 359 22781 461 22815
rect 495 22781 597 22815
rect 631 22781 733 22815
rect 767 22781 869 22815
rect 903 22781 1005 22815
rect 1039 22781 1141 22815
rect 1175 22781 1277 22815
rect 1311 22781 1413 22815
rect 1447 22781 1549 22815
rect 1583 22781 1685 22815
rect 325 22679 1719 22781
rect 359 22645 461 22679
rect 495 22645 597 22679
rect 631 22645 733 22679
rect 767 22645 869 22679
rect 903 22645 1005 22679
rect 1039 22645 1141 22679
rect 1175 22645 1277 22679
rect 1311 22645 1413 22679
rect 1447 22645 1549 22679
rect 1583 22645 1685 22679
rect 325 22543 1719 22645
rect 359 22509 461 22543
rect 495 22509 597 22543
rect 631 22509 733 22543
rect 767 22509 869 22543
rect 903 22509 1005 22543
rect 1039 22509 1141 22543
rect 1175 22509 1277 22543
rect 1311 22509 1413 22543
rect 1447 22509 1549 22543
rect 1583 22509 1685 22543
rect 325 22407 1719 22509
rect 359 22373 461 22407
rect 495 22373 597 22407
rect 631 22373 733 22407
rect 767 22373 869 22407
rect 903 22373 1005 22407
rect 1039 22373 1141 22407
rect 1175 22373 1277 22407
rect 1311 22373 1413 22407
rect 1447 22373 1549 22407
rect 1583 22373 1685 22407
rect 325 22271 1719 22373
rect 359 22237 461 22271
rect 495 22237 597 22271
rect 631 22237 733 22271
rect 767 22237 869 22271
rect 903 22237 1005 22271
rect 1039 22237 1141 22271
rect 1175 22237 1277 22271
rect 1311 22237 1413 22271
rect 1447 22237 1549 22271
rect 1583 22237 1685 22271
rect 325 22135 1719 22237
rect 359 22101 461 22135
rect 495 22101 597 22135
rect 631 22101 733 22135
rect 767 22101 869 22135
rect 903 22101 1005 22135
rect 1039 22101 1141 22135
rect 1175 22101 1277 22135
rect 1311 22101 1413 22135
rect 1447 22101 1549 22135
rect 1583 22101 1685 22135
rect 325 21999 1719 22101
rect 359 21965 461 21999
rect 495 21965 597 21999
rect 631 21965 733 21999
rect 767 21965 869 21999
rect 903 21965 1005 21999
rect 1039 21965 1141 21999
rect 1175 21965 1277 21999
rect 1311 21965 1413 21999
rect 1447 21965 1549 21999
rect 1583 21965 1685 21999
rect 325 21863 1719 21965
rect 359 21829 461 21863
rect 495 21829 597 21863
rect 631 21829 733 21863
rect 767 21829 869 21863
rect 903 21829 1005 21863
rect 1039 21829 1141 21863
rect 1175 21829 1277 21863
rect 1311 21829 1413 21863
rect 1447 21829 1549 21863
rect 1583 21829 1685 21863
rect 325 21727 1719 21829
rect 359 21693 461 21727
rect 495 21693 597 21727
rect 631 21693 733 21727
rect 767 21693 869 21727
rect 903 21693 1005 21727
rect 1039 21693 1141 21727
rect 1175 21693 1277 21727
rect 1311 21693 1413 21727
rect 1447 21693 1549 21727
rect 1583 21693 1685 21727
rect 325 21591 1719 21693
rect 359 21557 461 21591
rect 495 21557 597 21591
rect 631 21557 733 21591
rect 767 21557 869 21591
rect 903 21557 1005 21591
rect 1039 21557 1141 21591
rect 1175 21557 1277 21591
rect 1311 21557 1413 21591
rect 1447 21557 1549 21591
rect 1583 21557 1685 21591
rect 325 21455 1719 21557
rect 359 21421 461 21455
rect 495 21421 597 21455
rect 631 21421 733 21455
rect 767 21421 869 21455
rect 903 21421 1005 21455
rect 1039 21421 1141 21455
rect 1175 21421 1277 21455
rect 1311 21421 1413 21455
rect 1447 21421 1549 21455
rect 1583 21421 1685 21455
rect 325 21319 1719 21421
rect 359 21285 461 21319
rect 495 21285 597 21319
rect 631 21285 733 21319
rect 767 21285 869 21319
rect 903 21285 1005 21319
rect 1039 21285 1141 21319
rect 1175 21285 1277 21319
rect 1311 21285 1413 21319
rect 1447 21285 1549 21319
rect 1583 21285 1685 21319
rect 325 21183 1719 21285
rect 359 21149 461 21183
rect 495 21149 597 21183
rect 631 21149 733 21183
rect 767 21149 869 21183
rect 903 21149 1005 21183
rect 1039 21149 1141 21183
rect 1175 21149 1277 21183
rect 1311 21149 1413 21183
rect 1447 21149 1549 21183
rect 1583 21149 1685 21183
rect 325 21047 1719 21149
rect 359 21013 461 21047
rect 495 21013 597 21047
rect 631 21013 733 21047
rect 767 21013 869 21047
rect 903 21013 1005 21047
rect 1039 21013 1141 21047
rect 1175 21013 1277 21047
rect 1311 21013 1413 21047
rect 1447 21013 1549 21047
rect 1583 21013 1685 21047
rect 325 20911 1719 21013
rect 359 20877 461 20911
rect 495 20877 597 20911
rect 631 20877 733 20911
rect 767 20877 869 20911
rect 903 20877 1005 20911
rect 1039 20877 1141 20911
rect 1175 20877 1277 20911
rect 1311 20877 1413 20911
rect 1447 20877 1549 20911
rect 1583 20877 1685 20911
rect 325 20775 1719 20877
rect 359 20741 461 20775
rect 495 20741 597 20775
rect 631 20741 733 20775
rect 767 20741 869 20775
rect 903 20741 1005 20775
rect 1039 20741 1141 20775
rect 1175 20741 1277 20775
rect 1311 20741 1413 20775
rect 1447 20741 1549 20775
rect 1583 20741 1685 20775
rect 325 20639 1719 20741
rect 359 20605 461 20639
rect 495 20605 597 20639
rect 631 20605 733 20639
rect 767 20605 869 20639
rect 903 20605 1005 20639
rect 1039 20605 1141 20639
rect 1175 20605 1277 20639
rect 1311 20605 1413 20639
rect 1447 20605 1549 20639
rect 1583 20605 1685 20639
rect 325 20503 1719 20605
rect 359 20469 461 20503
rect 495 20469 597 20503
rect 631 20469 733 20503
rect 767 20469 869 20503
rect 903 20469 1005 20503
rect 1039 20469 1141 20503
rect 1175 20469 1277 20503
rect 1311 20469 1413 20503
rect 1447 20469 1549 20503
rect 1583 20469 1685 20503
rect 325 20367 1719 20469
rect 359 20333 461 20367
rect 495 20333 597 20367
rect 631 20333 733 20367
rect 767 20333 869 20367
rect 903 20333 1005 20367
rect 1039 20333 1141 20367
rect 1175 20333 1277 20367
rect 1311 20333 1413 20367
rect 1447 20333 1549 20367
rect 1583 20333 1685 20367
rect 325 20231 1719 20333
rect 359 20197 461 20231
rect 495 20197 597 20231
rect 631 20197 733 20231
rect 767 20197 869 20231
rect 903 20197 1005 20231
rect 1039 20197 1141 20231
rect 1175 20197 1277 20231
rect 1311 20197 1413 20231
rect 1447 20197 1549 20231
rect 1583 20197 1685 20231
rect 325 20095 1719 20197
rect 359 20061 461 20095
rect 495 20061 597 20095
rect 631 20061 733 20095
rect 767 20061 869 20095
rect 903 20061 1005 20095
rect 1039 20061 1141 20095
rect 1175 20061 1277 20095
rect 1311 20061 1413 20095
rect 1447 20061 1549 20095
rect 1583 20061 1685 20095
rect 325 19959 1719 20061
rect 359 19925 461 19959
rect 495 19925 597 19959
rect 631 19925 733 19959
rect 767 19925 869 19959
rect 903 19925 1005 19959
rect 1039 19925 1141 19959
rect 1175 19925 1277 19959
rect 1311 19925 1413 19959
rect 1447 19925 1549 19959
rect 1583 19925 1685 19959
rect 325 19823 1719 19925
rect 359 19789 461 19823
rect 495 19789 597 19823
rect 631 19789 733 19823
rect 767 19789 869 19823
rect 903 19789 1005 19823
rect 1039 19789 1141 19823
rect 1175 19789 1277 19823
rect 1311 19789 1413 19823
rect 1447 19789 1549 19823
rect 1583 19789 1685 19823
rect 325 19687 1719 19789
rect 359 19653 461 19687
rect 495 19653 597 19687
rect 631 19653 733 19687
rect 767 19653 869 19687
rect 903 19653 1005 19687
rect 1039 19653 1141 19687
rect 1175 19653 1277 19687
rect 1311 19653 1413 19687
rect 1447 19653 1549 19687
rect 1583 19653 1685 19687
rect 325 19551 1719 19653
rect 359 19517 461 19551
rect 495 19517 597 19551
rect 631 19517 733 19551
rect 767 19517 869 19551
rect 903 19517 1005 19551
rect 1039 19517 1141 19551
rect 1175 19517 1277 19551
rect 1311 19517 1413 19551
rect 1447 19517 1549 19551
rect 1583 19517 1685 19551
rect 325 19415 1719 19517
rect 359 19381 461 19415
rect 495 19381 597 19415
rect 631 19381 733 19415
rect 767 19381 869 19415
rect 903 19381 1005 19415
rect 1039 19381 1141 19415
rect 1175 19381 1277 19415
rect 1311 19381 1413 19415
rect 1447 19381 1549 19415
rect 1583 19381 1685 19415
rect 325 19279 1719 19381
rect 359 19245 461 19279
rect 495 19245 597 19279
rect 631 19245 733 19279
rect 767 19245 869 19279
rect 903 19245 1005 19279
rect 1039 19245 1141 19279
rect 1175 19245 1277 19279
rect 1311 19245 1413 19279
rect 1447 19245 1549 19279
rect 1583 19245 1685 19279
rect 325 19143 1719 19245
rect 359 19109 461 19143
rect 495 19109 597 19143
rect 631 19109 733 19143
rect 767 19109 869 19143
rect 903 19109 1005 19143
rect 1039 19109 1141 19143
rect 1175 19109 1277 19143
rect 1311 19109 1413 19143
rect 1447 19109 1549 19143
rect 1583 19109 1685 19143
rect 325 19007 1719 19109
rect 359 18973 461 19007
rect 495 18973 597 19007
rect 631 18973 733 19007
rect 767 18973 869 19007
rect 903 18973 1005 19007
rect 1039 18973 1141 19007
rect 1175 18973 1277 19007
rect 1311 18973 1413 19007
rect 1447 18973 1549 19007
rect 1583 18973 1685 19007
rect 325 18871 1719 18973
rect 359 18837 461 18871
rect 495 18837 597 18871
rect 631 18837 733 18871
rect 767 18837 869 18871
rect 903 18837 1005 18871
rect 1039 18837 1141 18871
rect 1175 18837 1277 18871
rect 1311 18837 1413 18871
rect 1447 18837 1549 18871
rect 1583 18837 1685 18871
rect 325 18735 1719 18837
rect 359 18701 461 18735
rect 495 18701 597 18735
rect 631 18701 733 18735
rect 767 18701 869 18735
rect 903 18701 1005 18735
rect 1039 18701 1141 18735
rect 1175 18701 1277 18735
rect 1311 18701 1413 18735
rect 1447 18701 1549 18735
rect 1583 18701 1685 18735
rect 325 18599 1719 18701
rect 359 18565 461 18599
rect 495 18565 597 18599
rect 631 18565 733 18599
rect 767 18565 869 18599
rect 903 18565 1005 18599
rect 1039 18565 1141 18599
rect 1175 18565 1277 18599
rect 1311 18565 1413 18599
rect 1447 18565 1549 18599
rect 1583 18565 1685 18599
rect 325 18463 1719 18565
rect 359 18429 461 18463
rect 495 18429 597 18463
rect 631 18429 733 18463
rect 767 18429 869 18463
rect 903 18429 1005 18463
rect 1039 18429 1141 18463
rect 1175 18429 1277 18463
rect 1311 18429 1413 18463
rect 1447 18429 1549 18463
rect 1583 18429 1685 18463
rect 325 18327 1719 18429
rect 359 18293 461 18327
rect 495 18293 597 18327
rect 631 18293 733 18327
rect 767 18293 869 18327
rect 903 18293 1005 18327
rect 1039 18293 1141 18327
rect 1175 18293 1277 18327
rect 1311 18293 1413 18327
rect 1447 18293 1549 18327
rect 1583 18293 1685 18327
rect 325 18191 1719 18293
rect 359 18157 461 18191
rect 495 18157 597 18191
rect 631 18157 733 18191
rect 767 18157 869 18191
rect 903 18157 1005 18191
rect 1039 18157 1141 18191
rect 1175 18157 1277 18191
rect 1311 18157 1413 18191
rect 1447 18157 1549 18191
rect 1583 18157 1685 18191
rect 325 18055 1719 18157
rect 359 18021 461 18055
rect 495 18021 597 18055
rect 631 18021 733 18055
rect 767 18021 869 18055
rect 903 18021 1005 18055
rect 1039 18021 1141 18055
rect 1175 18021 1277 18055
rect 1311 18021 1413 18055
rect 1447 18021 1549 18055
rect 1583 18021 1685 18055
rect 325 17919 1719 18021
rect 359 17885 461 17919
rect 495 17885 597 17919
rect 631 17885 733 17919
rect 767 17885 869 17919
rect 903 17885 1005 17919
rect 1039 17885 1141 17919
rect 1175 17885 1277 17919
rect 1311 17885 1413 17919
rect 1447 17885 1549 17919
rect 1583 17885 1685 17919
rect 325 17783 1719 17885
rect 359 17749 461 17783
rect 495 17749 597 17783
rect 631 17749 733 17783
rect 767 17749 869 17783
rect 903 17749 1005 17783
rect 1039 17749 1141 17783
rect 1175 17749 1277 17783
rect 1311 17749 1413 17783
rect 1447 17749 1549 17783
rect 1583 17749 1685 17783
rect 325 17647 1719 17749
rect 359 17613 461 17647
rect 495 17613 597 17647
rect 631 17613 733 17647
rect 767 17613 869 17647
rect 903 17613 1005 17647
rect 1039 17613 1141 17647
rect 1175 17613 1277 17647
rect 1311 17613 1413 17647
rect 1447 17613 1549 17647
rect 1583 17613 1685 17647
rect 325 17511 1719 17613
rect 359 17477 461 17511
rect 495 17477 597 17511
rect 631 17477 733 17511
rect 767 17477 869 17511
rect 903 17477 1005 17511
rect 1039 17477 1141 17511
rect 1175 17477 1277 17511
rect 1311 17477 1413 17511
rect 1447 17477 1549 17511
rect 1583 17477 1685 17511
rect 325 17375 1719 17477
rect 359 17341 461 17375
rect 495 17341 597 17375
rect 631 17341 733 17375
rect 767 17341 869 17375
rect 903 17341 1005 17375
rect 1039 17341 1141 17375
rect 1175 17341 1277 17375
rect 1311 17341 1413 17375
rect 1447 17341 1549 17375
rect 1583 17341 1685 17375
rect 325 17239 1719 17341
rect 359 17205 461 17239
rect 495 17205 597 17239
rect 631 17205 733 17239
rect 767 17205 869 17239
rect 903 17205 1005 17239
rect 1039 17205 1141 17239
rect 1175 17205 1277 17239
rect 1311 17205 1413 17239
rect 1447 17205 1549 17239
rect 1583 17205 1685 17239
rect 325 17103 1719 17205
rect 359 17069 461 17103
rect 495 17069 597 17103
rect 631 17069 733 17103
rect 767 17069 869 17103
rect 903 17069 1005 17103
rect 1039 17069 1141 17103
rect 1175 17069 1277 17103
rect 1311 17069 1413 17103
rect 1447 17069 1549 17103
rect 1583 17069 1685 17103
rect 325 16967 1719 17069
rect 359 16933 461 16967
rect 495 16933 597 16967
rect 631 16933 733 16967
rect 767 16933 869 16967
rect 903 16933 1005 16967
rect 1039 16933 1141 16967
rect 1175 16933 1277 16967
rect 1311 16933 1413 16967
rect 1447 16933 1549 16967
rect 1583 16933 1685 16967
rect 325 16831 1719 16933
rect 359 16797 461 16831
rect 495 16797 597 16831
rect 631 16797 733 16831
rect 767 16797 869 16831
rect 903 16797 1005 16831
rect 1039 16797 1141 16831
rect 1175 16797 1277 16831
rect 1311 16797 1413 16831
rect 1447 16797 1549 16831
rect 1583 16797 1685 16831
rect 325 16695 1719 16797
rect 359 16661 461 16695
rect 495 16661 597 16695
rect 631 16661 733 16695
rect 767 16661 869 16695
rect 903 16661 1005 16695
rect 1039 16661 1141 16695
rect 1175 16661 1277 16695
rect 1311 16661 1413 16695
rect 1447 16661 1549 16695
rect 1583 16661 1685 16695
rect 325 16559 1719 16661
rect 359 16525 461 16559
rect 495 16525 597 16559
rect 631 16525 733 16559
rect 767 16525 869 16559
rect 903 16525 1005 16559
rect 1039 16525 1141 16559
rect 1175 16525 1277 16559
rect 1311 16525 1413 16559
rect 1447 16525 1549 16559
rect 1583 16525 1685 16559
rect 325 16423 1719 16525
rect 7880 39951 9274 39975
rect 7914 39917 8016 39951
rect 8050 39917 8152 39951
rect 8186 39917 8288 39951
rect 8322 39917 8424 39951
rect 8458 39917 8560 39951
rect 8594 39917 8696 39951
rect 8730 39917 8832 39951
rect 8866 39917 8968 39951
rect 9002 39917 9104 39951
rect 9138 39917 9240 39951
rect 7880 39815 9274 39917
rect 7914 39781 8016 39815
rect 8050 39781 8152 39815
rect 8186 39781 8288 39815
rect 8322 39781 8424 39815
rect 8458 39781 8560 39815
rect 8594 39781 8696 39815
rect 8730 39781 8832 39815
rect 8866 39781 8968 39815
rect 9002 39781 9104 39815
rect 9138 39781 9240 39815
rect 7880 39679 9274 39781
rect 7914 39645 8016 39679
rect 8050 39645 8152 39679
rect 8186 39645 8288 39679
rect 8322 39645 8424 39679
rect 8458 39645 8560 39679
rect 8594 39645 8696 39679
rect 8730 39645 8832 39679
rect 8866 39645 8968 39679
rect 9002 39645 9104 39679
rect 9138 39645 9240 39679
rect 7880 39543 9274 39645
rect 7914 39509 8016 39543
rect 8050 39509 8152 39543
rect 8186 39509 8288 39543
rect 8322 39509 8424 39543
rect 8458 39509 8560 39543
rect 8594 39509 8696 39543
rect 8730 39509 8832 39543
rect 8866 39509 8968 39543
rect 9002 39509 9104 39543
rect 9138 39509 9240 39543
rect 7880 39407 9274 39509
rect 7914 39373 8016 39407
rect 8050 39373 8152 39407
rect 8186 39373 8288 39407
rect 8322 39373 8424 39407
rect 8458 39373 8560 39407
rect 8594 39373 8696 39407
rect 8730 39373 8832 39407
rect 8866 39373 8968 39407
rect 9002 39373 9104 39407
rect 9138 39373 9240 39407
rect 7880 39271 9274 39373
rect 7914 39237 8016 39271
rect 8050 39237 8152 39271
rect 8186 39237 8288 39271
rect 8322 39237 8424 39271
rect 8458 39237 8560 39271
rect 8594 39237 8696 39271
rect 8730 39237 8832 39271
rect 8866 39237 8968 39271
rect 9002 39237 9104 39271
rect 9138 39237 9240 39271
rect 7880 39135 9274 39237
rect 7914 39101 8016 39135
rect 8050 39101 8152 39135
rect 8186 39101 8288 39135
rect 8322 39101 8424 39135
rect 8458 39101 8560 39135
rect 8594 39101 8696 39135
rect 8730 39101 8832 39135
rect 8866 39101 8968 39135
rect 9002 39101 9104 39135
rect 9138 39101 9240 39135
rect 7880 38999 9274 39101
rect 7914 38965 8016 38999
rect 8050 38965 8152 38999
rect 8186 38965 8288 38999
rect 8322 38965 8424 38999
rect 8458 38965 8560 38999
rect 8594 38965 8696 38999
rect 8730 38965 8832 38999
rect 8866 38965 8968 38999
rect 9002 38965 9104 38999
rect 9138 38965 9240 38999
rect 7880 38863 9274 38965
rect 7914 38829 8016 38863
rect 8050 38829 8152 38863
rect 8186 38829 8288 38863
rect 8322 38829 8424 38863
rect 8458 38829 8560 38863
rect 8594 38829 8696 38863
rect 8730 38829 8832 38863
rect 8866 38829 8968 38863
rect 9002 38829 9104 38863
rect 9138 38829 9240 38863
rect 7880 38727 9274 38829
rect 7914 38693 8016 38727
rect 8050 38693 8152 38727
rect 8186 38693 8288 38727
rect 8322 38693 8424 38727
rect 8458 38693 8560 38727
rect 8594 38693 8696 38727
rect 8730 38693 8832 38727
rect 8866 38693 8968 38727
rect 9002 38693 9104 38727
rect 9138 38693 9240 38727
rect 7880 38591 9274 38693
rect 7914 38557 8016 38591
rect 8050 38557 8152 38591
rect 8186 38557 8288 38591
rect 8322 38557 8424 38591
rect 8458 38557 8560 38591
rect 8594 38557 8696 38591
rect 8730 38557 8832 38591
rect 8866 38557 8968 38591
rect 9002 38557 9104 38591
rect 9138 38557 9240 38591
rect 7880 38455 9274 38557
rect 7914 38421 8016 38455
rect 8050 38421 8152 38455
rect 8186 38421 8288 38455
rect 8322 38421 8424 38455
rect 8458 38421 8560 38455
rect 8594 38421 8696 38455
rect 8730 38421 8832 38455
rect 8866 38421 8968 38455
rect 9002 38421 9104 38455
rect 9138 38421 9240 38455
rect 7880 38319 9274 38421
rect 7914 38285 8016 38319
rect 8050 38285 8152 38319
rect 8186 38285 8288 38319
rect 8322 38285 8424 38319
rect 8458 38285 8560 38319
rect 8594 38285 8696 38319
rect 8730 38285 8832 38319
rect 8866 38285 8968 38319
rect 9002 38285 9104 38319
rect 9138 38285 9240 38319
rect 7880 38183 9274 38285
rect 7914 38149 8016 38183
rect 8050 38149 8152 38183
rect 8186 38149 8288 38183
rect 8322 38149 8424 38183
rect 8458 38149 8560 38183
rect 8594 38149 8696 38183
rect 8730 38149 8832 38183
rect 8866 38149 8968 38183
rect 9002 38149 9104 38183
rect 9138 38149 9240 38183
rect 7880 38047 9274 38149
rect 7914 38013 8016 38047
rect 8050 38013 8152 38047
rect 8186 38013 8288 38047
rect 8322 38013 8424 38047
rect 8458 38013 8560 38047
rect 8594 38013 8696 38047
rect 8730 38013 8832 38047
rect 8866 38013 8968 38047
rect 9002 38013 9104 38047
rect 9138 38013 9240 38047
rect 7880 37911 9274 38013
rect 7914 37877 8016 37911
rect 8050 37877 8152 37911
rect 8186 37877 8288 37911
rect 8322 37877 8424 37911
rect 8458 37877 8560 37911
rect 8594 37877 8696 37911
rect 8730 37877 8832 37911
rect 8866 37877 8968 37911
rect 9002 37877 9104 37911
rect 9138 37877 9240 37911
rect 7880 37775 9274 37877
rect 7914 37741 8016 37775
rect 8050 37741 8152 37775
rect 8186 37741 8288 37775
rect 8322 37741 8424 37775
rect 8458 37741 8560 37775
rect 8594 37741 8696 37775
rect 8730 37741 8832 37775
rect 8866 37741 8968 37775
rect 9002 37741 9104 37775
rect 9138 37741 9240 37775
rect 7880 37639 9274 37741
rect 7914 37605 8016 37639
rect 8050 37605 8152 37639
rect 8186 37605 8288 37639
rect 8322 37605 8424 37639
rect 8458 37605 8560 37639
rect 8594 37605 8696 37639
rect 8730 37605 8832 37639
rect 8866 37605 8968 37639
rect 9002 37605 9104 37639
rect 9138 37605 9240 37639
rect 7880 37503 9274 37605
rect 7914 37469 8016 37503
rect 8050 37469 8152 37503
rect 8186 37469 8288 37503
rect 8322 37469 8424 37503
rect 8458 37469 8560 37503
rect 8594 37469 8696 37503
rect 8730 37469 8832 37503
rect 8866 37469 8968 37503
rect 9002 37469 9104 37503
rect 9138 37469 9240 37503
rect 7880 37367 9274 37469
rect 7914 37333 8016 37367
rect 8050 37333 8152 37367
rect 8186 37333 8288 37367
rect 8322 37333 8424 37367
rect 8458 37333 8560 37367
rect 8594 37333 8696 37367
rect 8730 37333 8832 37367
rect 8866 37333 8968 37367
rect 9002 37333 9104 37367
rect 9138 37333 9240 37367
rect 7880 37231 9274 37333
rect 7914 37197 8016 37231
rect 8050 37197 8152 37231
rect 8186 37197 8288 37231
rect 8322 37197 8424 37231
rect 8458 37197 8560 37231
rect 8594 37197 8696 37231
rect 8730 37197 8832 37231
rect 8866 37197 8968 37231
rect 9002 37197 9104 37231
rect 9138 37197 9240 37231
rect 7880 37095 9274 37197
rect 7914 37061 8016 37095
rect 8050 37061 8152 37095
rect 8186 37061 8288 37095
rect 8322 37061 8424 37095
rect 8458 37061 8560 37095
rect 8594 37061 8696 37095
rect 8730 37061 8832 37095
rect 8866 37061 8968 37095
rect 9002 37061 9104 37095
rect 9138 37061 9240 37095
rect 7880 36959 9274 37061
rect 7914 36925 8016 36959
rect 8050 36925 8152 36959
rect 8186 36925 8288 36959
rect 8322 36925 8424 36959
rect 8458 36925 8560 36959
rect 8594 36925 8696 36959
rect 8730 36925 8832 36959
rect 8866 36925 8968 36959
rect 9002 36925 9104 36959
rect 9138 36925 9240 36959
rect 7880 36823 9274 36925
rect 7914 36789 8016 36823
rect 8050 36789 8152 36823
rect 8186 36789 8288 36823
rect 8322 36789 8424 36823
rect 8458 36789 8560 36823
rect 8594 36789 8696 36823
rect 8730 36789 8832 36823
rect 8866 36789 8968 36823
rect 9002 36789 9104 36823
rect 9138 36789 9240 36823
rect 7880 36687 9274 36789
rect 7914 36653 8016 36687
rect 8050 36653 8152 36687
rect 8186 36653 8288 36687
rect 8322 36653 8424 36687
rect 8458 36653 8560 36687
rect 8594 36653 8696 36687
rect 8730 36653 8832 36687
rect 8866 36653 8968 36687
rect 9002 36653 9104 36687
rect 9138 36653 9240 36687
rect 7880 36551 9274 36653
rect 7914 36517 8016 36551
rect 8050 36517 8152 36551
rect 8186 36517 8288 36551
rect 8322 36517 8424 36551
rect 8458 36517 8560 36551
rect 8594 36517 8696 36551
rect 8730 36517 8832 36551
rect 8866 36517 8968 36551
rect 9002 36517 9104 36551
rect 9138 36517 9240 36551
rect 7880 36415 9274 36517
rect 7914 36381 8016 36415
rect 8050 36381 8152 36415
rect 8186 36381 8288 36415
rect 8322 36381 8424 36415
rect 8458 36381 8560 36415
rect 8594 36381 8696 36415
rect 8730 36381 8832 36415
rect 8866 36381 8968 36415
rect 9002 36381 9104 36415
rect 9138 36381 9240 36415
rect 7880 36279 9274 36381
rect 7914 36245 8016 36279
rect 8050 36245 8152 36279
rect 8186 36245 8288 36279
rect 8322 36245 8424 36279
rect 8458 36245 8560 36279
rect 8594 36245 8696 36279
rect 8730 36245 8832 36279
rect 8866 36245 8968 36279
rect 9002 36245 9104 36279
rect 9138 36245 9240 36279
rect 7880 36143 9274 36245
rect 7914 36109 8016 36143
rect 8050 36109 8152 36143
rect 8186 36109 8288 36143
rect 8322 36109 8424 36143
rect 8458 36109 8560 36143
rect 8594 36109 8696 36143
rect 8730 36109 8832 36143
rect 8866 36109 8968 36143
rect 9002 36109 9104 36143
rect 9138 36109 9240 36143
rect 7880 36007 9274 36109
rect 7914 35973 8016 36007
rect 8050 35973 8152 36007
rect 8186 35973 8288 36007
rect 8322 35973 8424 36007
rect 8458 35973 8560 36007
rect 8594 35973 8696 36007
rect 8730 35973 8832 36007
rect 8866 35973 8968 36007
rect 9002 35973 9104 36007
rect 9138 35973 9240 36007
rect 7880 35871 9274 35973
rect 7914 35837 8016 35871
rect 8050 35837 8152 35871
rect 8186 35837 8288 35871
rect 8322 35837 8424 35871
rect 8458 35837 8560 35871
rect 8594 35837 8696 35871
rect 8730 35837 8832 35871
rect 8866 35837 8968 35871
rect 9002 35837 9104 35871
rect 9138 35837 9240 35871
rect 7880 35735 9274 35837
rect 7914 35701 8016 35735
rect 8050 35701 8152 35735
rect 8186 35701 8288 35735
rect 8322 35701 8424 35735
rect 8458 35701 8560 35735
rect 8594 35701 8696 35735
rect 8730 35701 8832 35735
rect 8866 35701 8968 35735
rect 9002 35701 9104 35735
rect 9138 35701 9240 35735
rect 7880 35599 9274 35701
rect 7914 35565 8016 35599
rect 8050 35565 8152 35599
rect 8186 35565 8288 35599
rect 8322 35565 8424 35599
rect 8458 35565 8560 35599
rect 8594 35565 8696 35599
rect 8730 35565 8832 35599
rect 8866 35565 8968 35599
rect 9002 35565 9104 35599
rect 9138 35565 9240 35599
rect 7880 35463 9274 35565
rect 7914 35429 8016 35463
rect 8050 35429 8152 35463
rect 8186 35429 8288 35463
rect 8322 35429 8424 35463
rect 8458 35429 8560 35463
rect 8594 35429 8696 35463
rect 8730 35429 8832 35463
rect 8866 35429 8968 35463
rect 9002 35429 9104 35463
rect 9138 35429 9240 35463
rect 7880 35327 9274 35429
rect 7914 35293 8016 35327
rect 8050 35293 8152 35327
rect 8186 35293 8288 35327
rect 8322 35293 8424 35327
rect 8458 35293 8560 35327
rect 8594 35293 8696 35327
rect 8730 35293 8832 35327
rect 8866 35293 8968 35327
rect 9002 35293 9104 35327
rect 9138 35293 9240 35327
rect 7880 35191 9274 35293
rect 7914 35157 8016 35191
rect 8050 35157 8152 35191
rect 8186 35157 8288 35191
rect 8322 35157 8424 35191
rect 8458 35157 8560 35191
rect 8594 35157 8696 35191
rect 8730 35157 8832 35191
rect 8866 35157 8968 35191
rect 9002 35157 9104 35191
rect 9138 35157 9240 35191
rect 7880 35055 9274 35157
rect 7914 35021 8016 35055
rect 8050 35021 8152 35055
rect 8186 35021 8288 35055
rect 8322 35021 8424 35055
rect 8458 35021 8560 35055
rect 8594 35021 8696 35055
rect 8730 35021 8832 35055
rect 8866 35021 8968 35055
rect 9002 35021 9104 35055
rect 9138 35021 9240 35055
rect 7880 34919 9274 35021
rect 7914 34885 8016 34919
rect 8050 34885 8152 34919
rect 8186 34885 8288 34919
rect 8322 34885 8424 34919
rect 8458 34885 8560 34919
rect 8594 34885 8696 34919
rect 8730 34885 8832 34919
rect 8866 34885 8968 34919
rect 9002 34885 9104 34919
rect 9138 34885 9240 34919
rect 7880 34783 9274 34885
rect 7914 34749 8016 34783
rect 8050 34749 8152 34783
rect 8186 34749 8288 34783
rect 8322 34749 8424 34783
rect 8458 34749 8560 34783
rect 8594 34749 8696 34783
rect 8730 34749 8832 34783
rect 8866 34749 8968 34783
rect 9002 34749 9104 34783
rect 9138 34749 9240 34783
rect 7880 34647 9274 34749
rect 7914 34613 8016 34647
rect 8050 34613 8152 34647
rect 8186 34613 8288 34647
rect 8322 34613 8424 34647
rect 8458 34613 8560 34647
rect 8594 34613 8696 34647
rect 8730 34613 8832 34647
rect 8866 34613 8968 34647
rect 9002 34613 9104 34647
rect 9138 34613 9240 34647
rect 7880 34511 9274 34613
rect 7914 34477 8016 34511
rect 8050 34477 8152 34511
rect 8186 34477 8288 34511
rect 8322 34477 8424 34511
rect 8458 34477 8560 34511
rect 8594 34477 8696 34511
rect 8730 34477 8832 34511
rect 8866 34477 8968 34511
rect 9002 34477 9104 34511
rect 9138 34477 9240 34511
rect 7880 34375 9274 34477
rect 7914 34341 8016 34375
rect 8050 34341 8152 34375
rect 8186 34341 8288 34375
rect 8322 34341 8424 34375
rect 8458 34341 8560 34375
rect 8594 34341 8696 34375
rect 8730 34341 8832 34375
rect 8866 34341 8968 34375
rect 9002 34341 9104 34375
rect 9138 34341 9240 34375
rect 7880 34239 9274 34341
rect 7914 34205 8016 34239
rect 8050 34205 8152 34239
rect 8186 34205 8288 34239
rect 8322 34205 8424 34239
rect 8458 34205 8560 34239
rect 8594 34205 8696 34239
rect 8730 34205 8832 34239
rect 8866 34205 8968 34239
rect 9002 34205 9104 34239
rect 9138 34205 9240 34239
rect 7880 34103 9274 34205
rect 7914 34069 8016 34103
rect 8050 34069 8152 34103
rect 8186 34069 8288 34103
rect 8322 34069 8424 34103
rect 8458 34069 8560 34103
rect 8594 34069 8696 34103
rect 8730 34069 8832 34103
rect 8866 34069 8968 34103
rect 9002 34069 9104 34103
rect 9138 34069 9240 34103
rect 7880 33967 9274 34069
rect 7914 33933 8016 33967
rect 8050 33933 8152 33967
rect 8186 33933 8288 33967
rect 8322 33933 8424 33967
rect 8458 33933 8560 33967
rect 8594 33933 8696 33967
rect 8730 33933 8832 33967
rect 8866 33933 8968 33967
rect 9002 33933 9104 33967
rect 9138 33933 9240 33967
rect 7880 33831 9274 33933
rect 7914 33797 8016 33831
rect 8050 33797 8152 33831
rect 8186 33797 8288 33831
rect 8322 33797 8424 33831
rect 8458 33797 8560 33831
rect 8594 33797 8696 33831
rect 8730 33797 8832 33831
rect 8866 33797 8968 33831
rect 9002 33797 9104 33831
rect 9138 33797 9240 33831
rect 7880 33695 9274 33797
rect 7914 33661 8016 33695
rect 8050 33661 8152 33695
rect 8186 33661 8288 33695
rect 8322 33661 8424 33695
rect 8458 33661 8560 33695
rect 8594 33661 8696 33695
rect 8730 33661 8832 33695
rect 8866 33661 8968 33695
rect 9002 33661 9104 33695
rect 9138 33661 9240 33695
rect 7880 33559 9274 33661
rect 7914 33525 8016 33559
rect 8050 33525 8152 33559
rect 8186 33525 8288 33559
rect 8322 33525 8424 33559
rect 8458 33525 8560 33559
rect 8594 33525 8696 33559
rect 8730 33525 8832 33559
rect 8866 33525 8968 33559
rect 9002 33525 9104 33559
rect 9138 33525 9240 33559
rect 7880 33423 9274 33525
rect 7914 33389 8016 33423
rect 8050 33389 8152 33423
rect 8186 33389 8288 33423
rect 8322 33389 8424 33423
rect 8458 33389 8560 33423
rect 8594 33389 8696 33423
rect 8730 33389 8832 33423
rect 8866 33389 8968 33423
rect 9002 33389 9104 33423
rect 9138 33389 9240 33423
rect 7880 33287 9274 33389
rect 7914 33253 8016 33287
rect 8050 33253 8152 33287
rect 8186 33253 8288 33287
rect 8322 33253 8424 33287
rect 8458 33253 8560 33287
rect 8594 33253 8696 33287
rect 8730 33253 8832 33287
rect 8866 33253 8968 33287
rect 9002 33253 9104 33287
rect 9138 33253 9240 33287
rect 7880 33151 9274 33253
rect 7914 33117 8016 33151
rect 8050 33117 8152 33151
rect 8186 33117 8288 33151
rect 8322 33117 8424 33151
rect 8458 33117 8560 33151
rect 8594 33117 8696 33151
rect 8730 33117 8832 33151
rect 8866 33117 8968 33151
rect 9002 33117 9104 33151
rect 9138 33117 9240 33151
rect 7880 33015 9274 33117
rect 7914 32981 8016 33015
rect 8050 32981 8152 33015
rect 8186 32981 8288 33015
rect 8322 32981 8424 33015
rect 8458 32981 8560 33015
rect 8594 32981 8696 33015
rect 8730 32981 8832 33015
rect 8866 32981 8968 33015
rect 9002 32981 9104 33015
rect 9138 32981 9240 33015
rect 7880 32879 9274 32981
rect 7914 32845 8016 32879
rect 8050 32845 8152 32879
rect 8186 32845 8288 32879
rect 8322 32845 8424 32879
rect 8458 32845 8560 32879
rect 8594 32845 8696 32879
rect 8730 32845 8832 32879
rect 8866 32845 8968 32879
rect 9002 32845 9104 32879
rect 9138 32845 9240 32879
rect 7880 32743 9274 32845
rect 7914 32709 8016 32743
rect 8050 32709 8152 32743
rect 8186 32709 8288 32743
rect 8322 32709 8424 32743
rect 8458 32709 8560 32743
rect 8594 32709 8696 32743
rect 8730 32709 8832 32743
rect 8866 32709 8968 32743
rect 9002 32709 9104 32743
rect 9138 32709 9240 32743
rect 7880 32607 9274 32709
rect 7914 32573 8016 32607
rect 8050 32573 8152 32607
rect 8186 32573 8288 32607
rect 8322 32573 8424 32607
rect 8458 32573 8560 32607
rect 8594 32573 8696 32607
rect 8730 32573 8832 32607
rect 8866 32573 8968 32607
rect 9002 32573 9104 32607
rect 9138 32573 9240 32607
rect 7880 32471 9274 32573
rect 7914 32437 8016 32471
rect 8050 32437 8152 32471
rect 8186 32437 8288 32471
rect 8322 32437 8424 32471
rect 8458 32437 8560 32471
rect 8594 32437 8696 32471
rect 8730 32437 8832 32471
rect 8866 32437 8968 32471
rect 9002 32437 9104 32471
rect 9138 32437 9240 32471
rect 7880 32335 9274 32437
rect 7914 32301 8016 32335
rect 8050 32301 8152 32335
rect 8186 32301 8288 32335
rect 8322 32301 8424 32335
rect 8458 32301 8560 32335
rect 8594 32301 8696 32335
rect 8730 32301 8832 32335
rect 8866 32301 8968 32335
rect 9002 32301 9104 32335
rect 9138 32301 9240 32335
rect 7880 32199 9274 32301
rect 7914 32165 8016 32199
rect 8050 32165 8152 32199
rect 8186 32165 8288 32199
rect 8322 32165 8424 32199
rect 8458 32165 8560 32199
rect 8594 32165 8696 32199
rect 8730 32165 8832 32199
rect 8866 32165 8968 32199
rect 9002 32165 9104 32199
rect 9138 32165 9240 32199
rect 7880 32063 9274 32165
rect 7914 32029 8016 32063
rect 8050 32029 8152 32063
rect 8186 32029 8288 32063
rect 8322 32029 8424 32063
rect 8458 32029 8560 32063
rect 8594 32029 8696 32063
rect 8730 32029 8832 32063
rect 8866 32029 8968 32063
rect 9002 32029 9104 32063
rect 9138 32029 9240 32063
rect 7880 31927 9274 32029
rect 7914 31893 8016 31927
rect 8050 31893 8152 31927
rect 8186 31893 8288 31927
rect 8322 31893 8424 31927
rect 8458 31893 8560 31927
rect 8594 31893 8696 31927
rect 8730 31893 8832 31927
rect 8866 31893 8968 31927
rect 9002 31893 9104 31927
rect 9138 31893 9240 31927
rect 7880 31791 9274 31893
rect 7914 31757 8016 31791
rect 8050 31757 8152 31791
rect 8186 31757 8288 31791
rect 8322 31757 8424 31791
rect 8458 31757 8560 31791
rect 8594 31757 8696 31791
rect 8730 31757 8832 31791
rect 8866 31757 8968 31791
rect 9002 31757 9104 31791
rect 9138 31757 9240 31791
rect 7880 31655 9274 31757
rect 7914 31621 8016 31655
rect 8050 31621 8152 31655
rect 8186 31621 8288 31655
rect 8322 31621 8424 31655
rect 8458 31621 8560 31655
rect 8594 31621 8696 31655
rect 8730 31621 8832 31655
rect 8866 31621 8968 31655
rect 9002 31621 9104 31655
rect 9138 31621 9240 31655
rect 7880 31519 9274 31621
rect 7914 31485 8016 31519
rect 8050 31485 8152 31519
rect 8186 31485 8288 31519
rect 8322 31485 8424 31519
rect 8458 31485 8560 31519
rect 8594 31485 8696 31519
rect 8730 31485 8832 31519
rect 8866 31485 8968 31519
rect 9002 31485 9104 31519
rect 9138 31485 9240 31519
rect 7880 31383 9274 31485
rect 7914 31349 8016 31383
rect 8050 31349 8152 31383
rect 8186 31349 8288 31383
rect 8322 31349 8424 31383
rect 8458 31349 8560 31383
rect 8594 31349 8696 31383
rect 8730 31349 8832 31383
rect 8866 31349 8968 31383
rect 9002 31349 9104 31383
rect 9138 31349 9240 31383
rect 7880 31247 9274 31349
rect 7914 31213 8016 31247
rect 8050 31213 8152 31247
rect 8186 31213 8288 31247
rect 8322 31213 8424 31247
rect 8458 31213 8560 31247
rect 8594 31213 8696 31247
rect 8730 31213 8832 31247
rect 8866 31213 8968 31247
rect 9002 31213 9104 31247
rect 9138 31213 9240 31247
rect 7880 31111 9274 31213
rect 7914 31077 8016 31111
rect 8050 31077 8152 31111
rect 8186 31077 8288 31111
rect 8322 31077 8424 31111
rect 8458 31077 8560 31111
rect 8594 31077 8696 31111
rect 8730 31077 8832 31111
rect 8866 31077 8968 31111
rect 9002 31077 9104 31111
rect 9138 31077 9240 31111
rect 7880 30975 9274 31077
rect 7914 30941 8016 30975
rect 8050 30941 8152 30975
rect 8186 30941 8288 30975
rect 8322 30941 8424 30975
rect 8458 30941 8560 30975
rect 8594 30941 8696 30975
rect 8730 30941 8832 30975
rect 8866 30941 8968 30975
rect 9002 30941 9104 30975
rect 9138 30941 9240 30975
rect 7880 30839 9274 30941
rect 7914 30805 8016 30839
rect 8050 30805 8152 30839
rect 8186 30805 8288 30839
rect 8322 30805 8424 30839
rect 8458 30805 8560 30839
rect 8594 30805 8696 30839
rect 8730 30805 8832 30839
rect 8866 30805 8968 30839
rect 9002 30805 9104 30839
rect 9138 30805 9240 30839
rect 7880 30703 9274 30805
rect 7914 30669 8016 30703
rect 8050 30669 8152 30703
rect 8186 30669 8288 30703
rect 8322 30669 8424 30703
rect 8458 30669 8560 30703
rect 8594 30669 8696 30703
rect 8730 30669 8832 30703
rect 8866 30669 8968 30703
rect 9002 30669 9104 30703
rect 9138 30669 9240 30703
rect 7880 30567 9274 30669
rect 7914 30533 8016 30567
rect 8050 30533 8152 30567
rect 8186 30533 8288 30567
rect 8322 30533 8424 30567
rect 8458 30533 8560 30567
rect 8594 30533 8696 30567
rect 8730 30533 8832 30567
rect 8866 30533 8968 30567
rect 9002 30533 9104 30567
rect 9138 30533 9240 30567
rect 7880 30431 9274 30533
rect 7914 30397 8016 30431
rect 8050 30397 8152 30431
rect 8186 30397 8288 30431
rect 8322 30397 8424 30431
rect 8458 30397 8560 30431
rect 8594 30397 8696 30431
rect 8730 30397 8832 30431
rect 8866 30397 8968 30431
rect 9002 30397 9104 30431
rect 9138 30397 9240 30431
rect 7880 30295 9274 30397
rect 7914 30261 8016 30295
rect 8050 30261 8152 30295
rect 8186 30261 8288 30295
rect 8322 30261 8424 30295
rect 8458 30261 8560 30295
rect 8594 30261 8696 30295
rect 8730 30261 8832 30295
rect 8866 30261 8968 30295
rect 9002 30261 9104 30295
rect 9138 30261 9240 30295
rect 7880 30159 9274 30261
rect 7914 30125 8016 30159
rect 8050 30125 8152 30159
rect 8186 30125 8288 30159
rect 8322 30125 8424 30159
rect 8458 30125 8560 30159
rect 8594 30125 8696 30159
rect 8730 30125 8832 30159
rect 8866 30125 8968 30159
rect 9002 30125 9104 30159
rect 9138 30125 9240 30159
rect 7880 30023 9274 30125
rect 7914 29989 8016 30023
rect 8050 29989 8152 30023
rect 8186 29989 8288 30023
rect 8322 29989 8424 30023
rect 8458 29989 8560 30023
rect 8594 29989 8696 30023
rect 8730 29989 8832 30023
rect 8866 29989 8968 30023
rect 9002 29989 9104 30023
rect 9138 29989 9240 30023
rect 7880 29887 9274 29989
rect 7914 29853 8016 29887
rect 8050 29853 8152 29887
rect 8186 29853 8288 29887
rect 8322 29853 8424 29887
rect 8458 29853 8560 29887
rect 8594 29853 8696 29887
rect 8730 29853 8832 29887
rect 8866 29853 8968 29887
rect 9002 29853 9104 29887
rect 9138 29853 9240 29887
rect 7880 29751 9274 29853
rect 7914 29717 8016 29751
rect 8050 29717 8152 29751
rect 8186 29717 8288 29751
rect 8322 29717 8424 29751
rect 8458 29717 8560 29751
rect 8594 29717 8696 29751
rect 8730 29717 8832 29751
rect 8866 29717 8968 29751
rect 9002 29717 9104 29751
rect 9138 29717 9240 29751
rect 7880 29615 9274 29717
rect 7914 29581 8016 29615
rect 8050 29581 8152 29615
rect 8186 29581 8288 29615
rect 8322 29581 8424 29615
rect 8458 29581 8560 29615
rect 8594 29581 8696 29615
rect 8730 29581 8832 29615
rect 8866 29581 8968 29615
rect 9002 29581 9104 29615
rect 9138 29581 9240 29615
rect 7880 29479 9274 29581
rect 7914 29445 8016 29479
rect 8050 29445 8152 29479
rect 8186 29445 8288 29479
rect 8322 29445 8424 29479
rect 8458 29445 8560 29479
rect 8594 29445 8696 29479
rect 8730 29445 8832 29479
rect 8866 29445 8968 29479
rect 9002 29445 9104 29479
rect 9138 29445 9240 29479
rect 7880 29343 9274 29445
rect 7914 29309 8016 29343
rect 8050 29309 8152 29343
rect 8186 29309 8288 29343
rect 8322 29309 8424 29343
rect 8458 29309 8560 29343
rect 8594 29309 8696 29343
rect 8730 29309 8832 29343
rect 8866 29309 8968 29343
rect 9002 29309 9104 29343
rect 9138 29309 9240 29343
rect 7880 29207 9274 29309
rect 7914 29173 8016 29207
rect 8050 29173 8152 29207
rect 8186 29173 8288 29207
rect 8322 29173 8424 29207
rect 8458 29173 8560 29207
rect 8594 29173 8696 29207
rect 8730 29173 8832 29207
rect 8866 29173 8968 29207
rect 9002 29173 9104 29207
rect 9138 29173 9240 29207
rect 7880 29071 9274 29173
rect 7914 29037 8016 29071
rect 8050 29037 8152 29071
rect 8186 29037 8288 29071
rect 8322 29037 8424 29071
rect 8458 29037 8560 29071
rect 8594 29037 8696 29071
rect 8730 29037 8832 29071
rect 8866 29037 8968 29071
rect 9002 29037 9104 29071
rect 9138 29037 9240 29071
rect 7880 28935 9274 29037
rect 7914 28901 8016 28935
rect 8050 28901 8152 28935
rect 8186 28901 8288 28935
rect 8322 28901 8424 28935
rect 8458 28901 8560 28935
rect 8594 28901 8696 28935
rect 8730 28901 8832 28935
rect 8866 28901 8968 28935
rect 9002 28901 9104 28935
rect 9138 28901 9240 28935
rect 7880 28799 9274 28901
rect 7914 28765 8016 28799
rect 8050 28765 8152 28799
rect 8186 28765 8288 28799
rect 8322 28765 8424 28799
rect 8458 28765 8560 28799
rect 8594 28765 8696 28799
rect 8730 28765 8832 28799
rect 8866 28765 8968 28799
rect 9002 28765 9104 28799
rect 9138 28765 9240 28799
rect 7880 28663 9274 28765
rect 7914 28629 8016 28663
rect 8050 28629 8152 28663
rect 8186 28629 8288 28663
rect 8322 28629 8424 28663
rect 8458 28629 8560 28663
rect 8594 28629 8696 28663
rect 8730 28629 8832 28663
rect 8866 28629 8968 28663
rect 9002 28629 9104 28663
rect 9138 28629 9240 28663
rect 7880 28527 9274 28629
rect 7914 28493 8016 28527
rect 8050 28493 8152 28527
rect 8186 28493 8288 28527
rect 8322 28493 8424 28527
rect 8458 28493 8560 28527
rect 8594 28493 8696 28527
rect 8730 28493 8832 28527
rect 8866 28493 8968 28527
rect 9002 28493 9104 28527
rect 9138 28493 9240 28527
rect 7880 28391 9274 28493
rect 7914 28357 8016 28391
rect 8050 28357 8152 28391
rect 8186 28357 8288 28391
rect 8322 28357 8424 28391
rect 8458 28357 8560 28391
rect 8594 28357 8696 28391
rect 8730 28357 8832 28391
rect 8866 28357 8968 28391
rect 9002 28357 9104 28391
rect 9138 28357 9240 28391
rect 7880 28255 9274 28357
rect 7914 28221 8016 28255
rect 8050 28221 8152 28255
rect 8186 28221 8288 28255
rect 8322 28221 8424 28255
rect 8458 28221 8560 28255
rect 8594 28221 8696 28255
rect 8730 28221 8832 28255
rect 8866 28221 8968 28255
rect 9002 28221 9104 28255
rect 9138 28221 9240 28255
rect 7880 28119 9274 28221
rect 7914 28085 8016 28119
rect 8050 28085 8152 28119
rect 8186 28085 8288 28119
rect 8322 28085 8424 28119
rect 8458 28085 8560 28119
rect 8594 28085 8696 28119
rect 8730 28085 8832 28119
rect 8866 28085 8968 28119
rect 9002 28085 9104 28119
rect 9138 28085 9240 28119
rect 7880 27983 9274 28085
rect 7914 27949 8016 27983
rect 8050 27949 8152 27983
rect 8186 27949 8288 27983
rect 8322 27949 8424 27983
rect 8458 27949 8560 27983
rect 8594 27949 8696 27983
rect 8730 27949 8832 27983
rect 8866 27949 8968 27983
rect 9002 27949 9104 27983
rect 9138 27949 9240 27983
rect 7880 27847 9274 27949
rect 7914 27813 8016 27847
rect 8050 27813 8152 27847
rect 8186 27813 8288 27847
rect 8322 27813 8424 27847
rect 8458 27813 8560 27847
rect 8594 27813 8696 27847
rect 8730 27813 8832 27847
rect 8866 27813 8968 27847
rect 9002 27813 9104 27847
rect 9138 27813 9240 27847
rect 7880 27711 9274 27813
rect 7914 27677 8016 27711
rect 8050 27677 8152 27711
rect 8186 27677 8288 27711
rect 8322 27677 8424 27711
rect 8458 27677 8560 27711
rect 8594 27677 8696 27711
rect 8730 27677 8832 27711
rect 8866 27677 8968 27711
rect 9002 27677 9104 27711
rect 9138 27677 9240 27711
rect 7880 27575 9274 27677
rect 7914 27541 8016 27575
rect 8050 27541 8152 27575
rect 8186 27541 8288 27575
rect 8322 27541 8424 27575
rect 8458 27541 8560 27575
rect 8594 27541 8696 27575
rect 8730 27541 8832 27575
rect 8866 27541 8968 27575
rect 9002 27541 9104 27575
rect 9138 27541 9240 27575
rect 7880 27439 9274 27541
rect 7914 27405 8016 27439
rect 8050 27405 8152 27439
rect 8186 27405 8288 27439
rect 8322 27405 8424 27439
rect 8458 27405 8560 27439
rect 8594 27405 8696 27439
rect 8730 27405 8832 27439
rect 8866 27405 8968 27439
rect 9002 27405 9104 27439
rect 9138 27405 9240 27439
rect 7880 27303 9274 27405
rect 7914 27269 8016 27303
rect 8050 27269 8152 27303
rect 8186 27269 8288 27303
rect 8322 27269 8424 27303
rect 8458 27269 8560 27303
rect 8594 27269 8696 27303
rect 8730 27269 8832 27303
rect 8866 27269 8968 27303
rect 9002 27269 9104 27303
rect 9138 27269 9240 27303
rect 7880 27167 9274 27269
rect 7914 27133 8016 27167
rect 8050 27133 8152 27167
rect 8186 27133 8288 27167
rect 8322 27133 8424 27167
rect 8458 27133 8560 27167
rect 8594 27133 8696 27167
rect 8730 27133 8832 27167
rect 8866 27133 8968 27167
rect 9002 27133 9104 27167
rect 9138 27133 9240 27167
rect 7880 27031 9274 27133
rect 7914 26997 8016 27031
rect 8050 26997 8152 27031
rect 8186 26997 8288 27031
rect 8322 26997 8424 27031
rect 8458 26997 8560 27031
rect 8594 26997 8696 27031
rect 8730 26997 8832 27031
rect 8866 26997 8968 27031
rect 9002 26997 9104 27031
rect 9138 26997 9240 27031
rect 7880 26895 9274 26997
rect 7914 26861 8016 26895
rect 8050 26861 8152 26895
rect 8186 26861 8288 26895
rect 8322 26861 8424 26895
rect 8458 26861 8560 26895
rect 8594 26861 8696 26895
rect 8730 26861 8832 26895
rect 8866 26861 8968 26895
rect 9002 26861 9104 26895
rect 9138 26861 9240 26895
rect 7880 26759 9274 26861
rect 7914 26725 8016 26759
rect 8050 26725 8152 26759
rect 8186 26725 8288 26759
rect 8322 26725 8424 26759
rect 8458 26725 8560 26759
rect 8594 26725 8696 26759
rect 8730 26725 8832 26759
rect 8866 26725 8968 26759
rect 9002 26725 9104 26759
rect 9138 26725 9240 26759
rect 7880 26623 9274 26725
rect 7914 26589 8016 26623
rect 8050 26589 8152 26623
rect 8186 26589 8288 26623
rect 8322 26589 8424 26623
rect 8458 26589 8560 26623
rect 8594 26589 8696 26623
rect 8730 26589 8832 26623
rect 8866 26589 8968 26623
rect 9002 26589 9104 26623
rect 9138 26589 9240 26623
rect 7880 26487 9274 26589
rect 7914 26453 8016 26487
rect 8050 26453 8152 26487
rect 8186 26453 8288 26487
rect 8322 26453 8424 26487
rect 8458 26453 8560 26487
rect 8594 26453 8696 26487
rect 8730 26453 8832 26487
rect 8866 26453 8968 26487
rect 9002 26453 9104 26487
rect 9138 26453 9240 26487
rect 7880 26351 9274 26453
rect 7914 26317 8016 26351
rect 8050 26317 8152 26351
rect 8186 26317 8288 26351
rect 8322 26317 8424 26351
rect 8458 26317 8560 26351
rect 8594 26317 8696 26351
rect 8730 26317 8832 26351
rect 8866 26317 8968 26351
rect 9002 26317 9104 26351
rect 9138 26317 9240 26351
rect 7880 26215 9274 26317
rect 7914 26181 8016 26215
rect 8050 26181 8152 26215
rect 8186 26181 8288 26215
rect 8322 26181 8424 26215
rect 8458 26181 8560 26215
rect 8594 26181 8696 26215
rect 8730 26181 8832 26215
rect 8866 26181 8968 26215
rect 9002 26181 9104 26215
rect 9138 26181 9240 26215
rect 7880 26079 9274 26181
rect 7914 26045 8016 26079
rect 8050 26045 8152 26079
rect 8186 26045 8288 26079
rect 8322 26045 8424 26079
rect 8458 26045 8560 26079
rect 8594 26045 8696 26079
rect 8730 26045 8832 26079
rect 8866 26045 8968 26079
rect 9002 26045 9104 26079
rect 9138 26045 9240 26079
rect 7880 25943 9274 26045
rect 7914 25909 8016 25943
rect 8050 25909 8152 25943
rect 8186 25909 8288 25943
rect 8322 25909 8424 25943
rect 8458 25909 8560 25943
rect 8594 25909 8696 25943
rect 8730 25909 8832 25943
rect 8866 25909 8968 25943
rect 9002 25909 9104 25943
rect 9138 25909 9240 25943
rect 7880 25807 9274 25909
rect 7914 25773 8016 25807
rect 8050 25773 8152 25807
rect 8186 25773 8288 25807
rect 8322 25773 8424 25807
rect 8458 25773 8560 25807
rect 8594 25773 8696 25807
rect 8730 25773 8832 25807
rect 8866 25773 8968 25807
rect 9002 25773 9104 25807
rect 9138 25773 9240 25807
rect 7880 25671 9274 25773
rect 7914 25637 8016 25671
rect 8050 25637 8152 25671
rect 8186 25637 8288 25671
rect 8322 25637 8424 25671
rect 8458 25637 8560 25671
rect 8594 25637 8696 25671
rect 8730 25637 8832 25671
rect 8866 25637 8968 25671
rect 9002 25637 9104 25671
rect 9138 25637 9240 25671
rect 7880 25535 9274 25637
rect 7914 25501 8016 25535
rect 8050 25501 8152 25535
rect 8186 25501 8288 25535
rect 8322 25501 8424 25535
rect 8458 25501 8560 25535
rect 8594 25501 8696 25535
rect 8730 25501 8832 25535
rect 8866 25501 8968 25535
rect 9002 25501 9104 25535
rect 9138 25501 9240 25535
rect 7880 25399 9274 25501
rect 7914 25365 8016 25399
rect 8050 25365 8152 25399
rect 8186 25365 8288 25399
rect 8322 25365 8424 25399
rect 8458 25365 8560 25399
rect 8594 25365 8696 25399
rect 8730 25365 8832 25399
rect 8866 25365 8968 25399
rect 9002 25365 9104 25399
rect 9138 25365 9240 25399
rect 7880 25263 9274 25365
rect 7914 25229 8016 25263
rect 8050 25229 8152 25263
rect 8186 25229 8288 25263
rect 8322 25229 8424 25263
rect 8458 25229 8560 25263
rect 8594 25229 8696 25263
rect 8730 25229 8832 25263
rect 8866 25229 8968 25263
rect 9002 25229 9104 25263
rect 9138 25229 9240 25263
rect 7880 25127 9274 25229
rect 7914 25093 8016 25127
rect 8050 25093 8152 25127
rect 8186 25093 8288 25127
rect 8322 25093 8424 25127
rect 8458 25093 8560 25127
rect 8594 25093 8696 25127
rect 8730 25093 8832 25127
rect 8866 25093 8968 25127
rect 9002 25093 9104 25127
rect 9138 25093 9240 25127
rect 7880 24991 9274 25093
rect 7914 24957 8016 24991
rect 8050 24957 8152 24991
rect 8186 24957 8288 24991
rect 8322 24957 8424 24991
rect 8458 24957 8560 24991
rect 8594 24957 8696 24991
rect 8730 24957 8832 24991
rect 8866 24957 8968 24991
rect 9002 24957 9104 24991
rect 9138 24957 9240 24991
rect 7880 24855 9274 24957
rect 7914 24821 8016 24855
rect 8050 24821 8152 24855
rect 8186 24821 8288 24855
rect 8322 24821 8424 24855
rect 8458 24821 8560 24855
rect 8594 24821 8696 24855
rect 8730 24821 8832 24855
rect 8866 24821 8968 24855
rect 9002 24821 9104 24855
rect 9138 24821 9240 24855
rect 7880 24719 9274 24821
rect 7914 24685 8016 24719
rect 8050 24685 8152 24719
rect 8186 24685 8288 24719
rect 8322 24685 8424 24719
rect 8458 24685 8560 24719
rect 8594 24685 8696 24719
rect 8730 24685 8832 24719
rect 8866 24685 8968 24719
rect 9002 24685 9104 24719
rect 9138 24685 9240 24719
rect 7880 24583 9274 24685
rect 7914 24549 8016 24583
rect 8050 24549 8152 24583
rect 8186 24549 8288 24583
rect 8322 24549 8424 24583
rect 8458 24549 8560 24583
rect 8594 24549 8696 24583
rect 8730 24549 8832 24583
rect 8866 24549 8968 24583
rect 9002 24549 9104 24583
rect 9138 24549 9240 24583
rect 7880 24447 9274 24549
rect 7914 24413 8016 24447
rect 8050 24413 8152 24447
rect 8186 24413 8288 24447
rect 8322 24413 8424 24447
rect 8458 24413 8560 24447
rect 8594 24413 8696 24447
rect 8730 24413 8832 24447
rect 8866 24413 8968 24447
rect 9002 24413 9104 24447
rect 9138 24413 9240 24447
rect 7880 24311 9274 24413
rect 7914 24277 8016 24311
rect 8050 24277 8152 24311
rect 8186 24277 8288 24311
rect 8322 24277 8424 24311
rect 8458 24277 8560 24311
rect 8594 24277 8696 24311
rect 8730 24277 8832 24311
rect 8866 24277 8968 24311
rect 9002 24277 9104 24311
rect 9138 24277 9240 24311
rect 7880 24175 9274 24277
rect 7914 24141 8016 24175
rect 8050 24141 8152 24175
rect 8186 24141 8288 24175
rect 8322 24141 8424 24175
rect 8458 24141 8560 24175
rect 8594 24141 8696 24175
rect 8730 24141 8832 24175
rect 8866 24141 8968 24175
rect 9002 24141 9104 24175
rect 9138 24141 9240 24175
rect 7880 24039 9274 24141
rect 7914 24005 8016 24039
rect 8050 24005 8152 24039
rect 8186 24005 8288 24039
rect 8322 24005 8424 24039
rect 8458 24005 8560 24039
rect 8594 24005 8696 24039
rect 8730 24005 8832 24039
rect 8866 24005 8968 24039
rect 9002 24005 9104 24039
rect 9138 24005 9240 24039
rect 7880 23903 9274 24005
rect 7914 23869 8016 23903
rect 8050 23869 8152 23903
rect 8186 23869 8288 23903
rect 8322 23869 8424 23903
rect 8458 23869 8560 23903
rect 8594 23869 8696 23903
rect 8730 23869 8832 23903
rect 8866 23869 8968 23903
rect 9002 23869 9104 23903
rect 9138 23869 9240 23903
rect 7880 23767 9274 23869
rect 7914 23733 8016 23767
rect 8050 23733 8152 23767
rect 8186 23733 8288 23767
rect 8322 23733 8424 23767
rect 8458 23733 8560 23767
rect 8594 23733 8696 23767
rect 8730 23733 8832 23767
rect 8866 23733 8968 23767
rect 9002 23733 9104 23767
rect 9138 23733 9240 23767
rect 7880 23631 9274 23733
rect 7914 23597 8016 23631
rect 8050 23597 8152 23631
rect 8186 23597 8288 23631
rect 8322 23597 8424 23631
rect 8458 23597 8560 23631
rect 8594 23597 8696 23631
rect 8730 23597 8832 23631
rect 8866 23597 8968 23631
rect 9002 23597 9104 23631
rect 9138 23597 9240 23631
rect 7880 23495 9274 23597
rect 7914 23461 8016 23495
rect 8050 23461 8152 23495
rect 8186 23461 8288 23495
rect 8322 23461 8424 23495
rect 8458 23461 8560 23495
rect 8594 23461 8696 23495
rect 8730 23461 8832 23495
rect 8866 23461 8968 23495
rect 9002 23461 9104 23495
rect 9138 23461 9240 23495
rect 7880 23359 9274 23461
rect 7914 23325 8016 23359
rect 8050 23325 8152 23359
rect 8186 23325 8288 23359
rect 8322 23325 8424 23359
rect 8458 23325 8560 23359
rect 8594 23325 8696 23359
rect 8730 23325 8832 23359
rect 8866 23325 8968 23359
rect 9002 23325 9104 23359
rect 9138 23325 9240 23359
rect 7880 23223 9274 23325
rect 7914 23189 8016 23223
rect 8050 23189 8152 23223
rect 8186 23189 8288 23223
rect 8322 23189 8424 23223
rect 8458 23189 8560 23223
rect 8594 23189 8696 23223
rect 8730 23189 8832 23223
rect 8866 23189 8968 23223
rect 9002 23189 9104 23223
rect 9138 23189 9240 23223
rect 7880 23087 9274 23189
rect 7914 23053 8016 23087
rect 8050 23053 8152 23087
rect 8186 23053 8288 23087
rect 8322 23053 8424 23087
rect 8458 23053 8560 23087
rect 8594 23053 8696 23087
rect 8730 23053 8832 23087
rect 8866 23053 8968 23087
rect 9002 23053 9104 23087
rect 9138 23053 9240 23087
rect 7880 22951 9274 23053
rect 7914 22917 8016 22951
rect 8050 22917 8152 22951
rect 8186 22917 8288 22951
rect 8322 22917 8424 22951
rect 8458 22917 8560 22951
rect 8594 22917 8696 22951
rect 8730 22917 8832 22951
rect 8866 22917 8968 22951
rect 9002 22917 9104 22951
rect 9138 22917 9240 22951
rect 7880 22815 9274 22917
rect 7914 22781 8016 22815
rect 8050 22781 8152 22815
rect 8186 22781 8288 22815
rect 8322 22781 8424 22815
rect 8458 22781 8560 22815
rect 8594 22781 8696 22815
rect 8730 22781 8832 22815
rect 8866 22781 8968 22815
rect 9002 22781 9104 22815
rect 9138 22781 9240 22815
rect 7880 22679 9274 22781
rect 7914 22645 8016 22679
rect 8050 22645 8152 22679
rect 8186 22645 8288 22679
rect 8322 22645 8424 22679
rect 8458 22645 8560 22679
rect 8594 22645 8696 22679
rect 8730 22645 8832 22679
rect 8866 22645 8968 22679
rect 9002 22645 9104 22679
rect 9138 22645 9240 22679
rect 7880 22543 9274 22645
rect 7914 22509 8016 22543
rect 8050 22509 8152 22543
rect 8186 22509 8288 22543
rect 8322 22509 8424 22543
rect 8458 22509 8560 22543
rect 8594 22509 8696 22543
rect 8730 22509 8832 22543
rect 8866 22509 8968 22543
rect 9002 22509 9104 22543
rect 9138 22509 9240 22543
rect 7880 22407 9274 22509
rect 7914 22373 8016 22407
rect 8050 22373 8152 22407
rect 8186 22373 8288 22407
rect 8322 22373 8424 22407
rect 8458 22373 8560 22407
rect 8594 22373 8696 22407
rect 8730 22373 8832 22407
rect 8866 22373 8968 22407
rect 9002 22373 9104 22407
rect 9138 22373 9240 22407
rect 7880 22271 9274 22373
rect 7914 22237 8016 22271
rect 8050 22237 8152 22271
rect 8186 22237 8288 22271
rect 8322 22237 8424 22271
rect 8458 22237 8560 22271
rect 8594 22237 8696 22271
rect 8730 22237 8832 22271
rect 8866 22237 8968 22271
rect 9002 22237 9104 22271
rect 9138 22237 9240 22271
rect 7880 22135 9274 22237
rect 7914 22101 8016 22135
rect 8050 22101 8152 22135
rect 8186 22101 8288 22135
rect 8322 22101 8424 22135
rect 8458 22101 8560 22135
rect 8594 22101 8696 22135
rect 8730 22101 8832 22135
rect 8866 22101 8968 22135
rect 9002 22101 9104 22135
rect 9138 22101 9240 22135
rect 7880 21999 9274 22101
rect 7914 21965 8016 21999
rect 8050 21965 8152 21999
rect 8186 21965 8288 21999
rect 8322 21965 8424 21999
rect 8458 21965 8560 21999
rect 8594 21965 8696 21999
rect 8730 21965 8832 21999
rect 8866 21965 8968 21999
rect 9002 21965 9104 21999
rect 9138 21965 9240 21999
rect 7880 21863 9274 21965
rect 7914 21829 8016 21863
rect 8050 21829 8152 21863
rect 8186 21829 8288 21863
rect 8322 21829 8424 21863
rect 8458 21829 8560 21863
rect 8594 21829 8696 21863
rect 8730 21829 8832 21863
rect 8866 21829 8968 21863
rect 9002 21829 9104 21863
rect 9138 21829 9240 21863
rect 7880 21727 9274 21829
rect 7914 21693 8016 21727
rect 8050 21693 8152 21727
rect 8186 21693 8288 21727
rect 8322 21693 8424 21727
rect 8458 21693 8560 21727
rect 8594 21693 8696 21727
rect 8730 21693 8832 21727
rect 8866 21693 8968 21727
rect 9002 21693 9104 21727
rect 9138 21693 9240 21727
rect 7880 21591 9274 21693
rect 7914 21557 8016 21591
rect 8050 21557 8152 21591
rect 8186 21557 8288 21591
rect 8322 21557 8424 21591
rect 8458 21557 8560 21591
rect 8594 21557 8696 21591
rect 8730 21557 8832 21591
rect 8866 21557 8968 21591
rect 9002 21557 9104 21591
rect 9138 21557 9240 21591
rect 7880 21455 9274 21557
rect 7914 21421 8016 21455
rect 8050 21421 8152 21455
rect 8186 21421 8288 21455
rect 8322 21421 8424 21455
rect 8458 21421 8560 21455
rect 8594 21421 8696 21455
rect 8730 21421 8832 21455
rect 8866 21421 8968 21455
rect 9002 21421 9104 21455
rect 9138 21421 9240 21455
rect 7880 21319 9274 21421
rect 7914 21285 8016 21319
rect 8050 21285 8152 21319
rect 8186 21285 8288 21319
rect 8322 21285 8424 21319
rect 8458 21285 8560 21319
rect 8594 21285 8696 21319
rect 8730 21285 8832 21319
rect 8866 21285 8968 21319
rect 9002 21285 9104 21319
rect 9138 21285 9240 21319
rect 7880 21183 9274 21285
rect 7914 21149 8016 21183
rect 8050 21149 8152 21183
rect 8186 21149 8288 21183
rect 8322 21149 8424 21183
rect 8458 21149 8560 21183
rect 8594 21149 8696 21183
rect 8730 21149 8832 21183
rect 8866 21149 8968 21183
rect 9002 21149 9104 21183
rect 9138 21149 9240 21183
rect 7880 21047 9274 21149
rect 7914 21013 8016 21047
rect 8050 21013 8152 21047
rect 8186 21013 8288 21047
rect 8322 21013 8424 21047
rect 8458 21013 8560 21047
rect 8594 21013 8696 21047
rect 8730 21013 8832 21047
rect 8866 21013 8968 21047
rect 9002 21013 9104 21047
rect 9138 21013 9240 21047
rect 7880 20911 9274 21013
rect 7914 20877 8016 20911
rect 8050 20877 8152 20911
rect 8186 20877 8288 20911
rect 8322 20877 8424 20911
rect 8458 20877 8560 20911
rect 8594 20877 8696 20911
rect 8730 20877 8832 20911
rect 8866 20877 8968 20911
rect 9002 20877 9104 20911
rect 9138 20877 9240 20911
rect 7880 20775 9274 20877
rect 7914 20741 8016 20775
rect 8050 20741 8152 20775
rect 8186 20741 8288 20775
rect 8322 20741 8424 20775
rect 8458 20741 8560 20775
rect 8594 20741 8696 20775
rect 8730 20741 8832 20775
rect 8866 20741 8968 20775
rect 9002 20741 9104 20775
rect 9138 20741 9240 20775
rect 7880 20639 9274 20741
rect 7914 20605 8016 20639
rect 8050 20605 8152 20639
rect 8186 20605 8288 20639
rect 8322 20605 8424 20639
rect 8458 20605 8560 20639
rect 8594 20605 8696 20639
rect 8730 20605 8832 20639
rect 8866 20605 8968 20639
rect 9002 20605 9104 20639
rect 9138 20605 9240 20639
rect 7880 20503 9274 20605
rect 7914 20469 8016 20503
rect 8050 20469 8152 20503
rect 8186 20469 8288 20503
rect 8322 20469 8424 20503
rect 8458 20469 8560 20503
rect 8594 20469 8696 20503
rect 8730 20469 8832 20503
rect 8866 20469 8968 20503
rect 9002 20469 9104 20503
rect 9138 20469 9240 20503
rect 7880 20367 9274 20469
rect 7914 20333 8016 20367
rect 8050 20333 8152 20367
rect 8186 20333 8288 20367
rect 8322 20333 8424 20367
rect 8458 20333 8560 20367
rect 8594 20333 8696 20367
rect 8730 20333 8832 20367
rect 8866 20333 8968 20367
rect 9002 20333 9104 20367
rect 9138 20333 9240 20367
rect 7880 20231 9274 20333
rect 7914 20197 8016 20231
rect 8050 20197 8152 20231
rect 8186 20197 8288 20231
rect 8322 20197 8424 20231
rect 8458 20197 8560 20231
rect 8594 20197 8696 20231
rect 8730 20197 8832 20231
rect 8866 20197 8968 20231
rect 9002 20197 9104 20231
rect 9138 20197 9240 20231
rect 7880 20095 9274 20197
rect 7914 20061 8016 20095
rect 8050 20061 8152 20095
rect 8186 20061 8288 20095
rect 8322 20061 8424 20095
rect 8458 20061 8560 20095
rect 8594 20061 8696 20095
rect 8730 20061 8832 20095
rect 8866 20061 8968 20095
rect 9002 20061 9104 20095
rect 9138 20061 9240 20095
rect 7880 19959 9274 20061
rect 7914 19925 8016 19959
rect 8050 19925 8152 19959
rect 8186 19925 8288 19959
rect 8322 19925 8424 19959
rect 8458 19925 8560 19959
rect 8594 19925 8696 19959
rect 8730 19925 8832 19959
rect 8866 19925 8968 19959
rect 9002 19925 9104 19959
rect 9138 19925 9240 19959
rect 7880 19823 9274 19925
rect 7914 19789 8016 19823
rect 8050 19789 8152 19823
rect 8186 19789 8288 19823
rect 8322 19789 8424 19823
rect 8458 19789 8560 19823
rect 8594 19789 8696 19823
rect 8730 19789 8832 19823
rect 8866 19789 8968 19823
rect 9002 19789 9104 19823
rect 9138 19789 9240 19823
rect 7880 19687 9274 19789
rect 7914 19653 8016 19687
rect 8050 19653 8152 19687
rect 8186 19653 8288 19687
rect 8322 19653 8424 19687
rect 8458 19653 8560 19687
rect 8594 19653 8696 19687
rect 8730 19653 8832 19687
rect 8866 19653 8968 19687
rect 9002 19653 9104 19687
rect 9138 19653 9240 19687
rect 7880 19551 9274 19653
rect 7914 19517 8016 19551
rect 8050 19517 8152 19551
rect 8186 19517 8288 19551
rect 8322 19517 8424 19551
rect 8458 19517 8560 19551
rect 8594 19517 8696 19551
rect 8730 19517 8832 19551
rect 8866 19517 8968 19551
rect 9002 19517 9104 19551
rect 9138 19517 9240 19551
rect 7880 19415 9274 19517
rect 7914 19381 8016 19415
rect 8050 19381 8152 19415
rect 8186 19381 8288 19415
rect 8322 19381 8424 19415
rect 8458 19381 8560 19415
rect 8594 19381 8696 19415
rect 8730 19381 8832 19415
rect 8866 19381 8968 19415
rect 9002 19381 9104 19415
rect 9138 19381 9240 19415
rect 7880 19279 9274 19381
rect 7914 19245 8016 19279
rect 8050 19245 8152 19279
rect 8186 19245 8288 19279
rect 8322 19245 8424 19279
rect 8458 19245 8560 19279
rect 8594 19245 8696 19279
rect 8730 19245 8832 19279
rect 8866 19245 8968 19279
rect 9002 19245 9104 19279
rect 9138 19245 9240 19279
rect 7880 19143 9274 19245
rect 7914 19109 8016 19143
rect 8050 19109 8152 19143
rect 8186 19109 8288 19143
rect 8322 19109 8424 19143
rect 8458 19109 8560 19143
rect 8594 19109 8696 19143
rect 8730 19109 8832 19143
rect 8866 19109 8968 19143
rect 9002 19109 9104 19143
rect 9138 19109 9240 19143
rect 7880 19007 9274 19109
rect 7914 18973 8016 19007
rect 8050 18973 8152 19007
rect 8186 18973 8288 19007
rect 8322 18973 8424 19007
rect 8458 18973 8560 19007
rect 8594 18973 8696 19007
rect 8730 18973 8832 19007
rect 8866 18973 8968 19007
rect 9002 18973 9104 19007
rect 9138 18973 9240 19007
rect 7880 18871 9274 18973
rect 7914 18837 8016 18871
rect 8050 18837 8152 18871
rect 8186 18837 8288 18871
rect 8322 18837 8424 18871
rect 8458 18837 8560 18871
rect 8594 18837 8696 18871
rect 8730 18837 8832 18871
rect 8866 18837 8968 18871
rect 9002 18837 9104 18871
rect 9138 18837 9240 18871
rect 7880 18735 9274 18837
rect 7914 18701 8016 18735
rect 8050 18701 8152 18735
rect 8186 18701 8288 18735
rect 8322 18701 8424 18735
rect 8458 18701 8560 18735
rect 8594 18701 8696 18735
rect 8730 18701 8832 18735
rect 8866 18701 8968 18735
rect 9002 18701 9104 18735
rect 9138 18701 9240 18735
rect 7880 18599 9274 18701
rect 7914 18565 8016 18599
rect 8050 18565 8152 18599
rect 8186 18565 8288 18599
rect 8322 18565 8424 18599
rect 8458 18565 8560 18599
rect 8594 18565 8696 18599
rect 8730 18565 8832 18599
rect 8866 18565 8968 18599
rect 9002 18565 9104 18599
rect 9138 18565 9240 18599
rect 7880 18463 9274 18565
rect 7914 18429 8016 18463
rect 8050 18429 8152 18463
rect 8186 18429 8288 18463
rect 8322 18429 8424 18463
rect 8458 18429 8560 18463
rect 8594 18429 8696 18463
rect 8730 18429 8832 18463
rect 8866 18429 8968 18463
rect 9002 18429 9104 18463
rect 9138 18429 9240 18463
rect 7880 18327 9274 18429
rect 7914 18293 8016 18327
rect 8050 18293 8152 18327
rect 8186 18293 8288 18327
rect 8322 18293 8424 18327
rect 8458 18293 8560 18327
rect 8594 18293 8696 18327
rect 8730 18293 8832 18327
rect 8866 18293 8968 18327
rect 9002 18293 9104 18327
rect 9138 18293 9240 18327
rect 7880 18191 9274 18293
rect 7914 18157 8016 18191
rect 8050 18157 8152 18191
rect 8186 18157 8288 18191
rect 8322 18157 8424 18191
rect 8458 18157 8560 18191
rect 8594 18157 8696 18191
rect 8730 18157 8832 18191
rect 8866 18157 8968 18191
rect 9002 18157 9104 18191
rect 9138 18157 9240 18191
rect 7880 18055 9274 18157
rect 7914 18021 8016 18055
rect 8050 18021 8152 18055
rect 8186 18021 8288 18055
rect 8322 18021 8424 18055
rect 8458 18021 8560 18055
rect 8594 18021 8696 18055
rect 8730 18021 8832 18055
rect 8866 18021 8968 18055
rect 9002 18021 9104 18055
rect 9138 18021 9240 18055
rect 7880 17919 9274 18021
rect 7914 17885 8016 17919
rect 8050 17885 8152 17919
rect 8186 17885 8288 17919
rect 8322 17885 8424 17919
rect 8458 17885 8560 17919
rect 8594 17885 8696 17919
rect 8730 17885 8832 17919
rect 8866 17885 8968 17919
rect 9002 17885 9104 17919
rect 9138 17885 9240 17919
rect 7880 17783 9274 17885
rect 7914 17749 8016 17783
rect 8050 17749 8152 17783
rect 8186 17749 8288 17783
rect 8322 17749 8424 17783
rect 8458 17749 8560 17783
rect 8594 17749 8696 17783
rect 8730 17749 8832 17783
rect 8866 17749 8968 17783
rect 9002 17749 9104 17783
rect 9138 17749 9240 17783
rect 7880 17647 9274 17749
rect 7914 17613 8016 17647
rect 8050 17613 8152 17647
rect 8186 17613 8288 17647
rect 8322 17613 8424 17647
rect 8458 17613 8560 17647
rect 8594 17613 8696 17647
rect 8730 17613 8832 17647
rect 8866 17613 8968 17647
rect 9002 17613 9104 17647
rect 9138 17613 9240 17647
rect 7880 17511 9274 17613
rect 7914 17477 8016 17511
rect 8050 17477 8152 17511
rect 8186 17477 8288 17511
rect 8322 17477 8424 17511
rect 8458 17477 8560 17511
rect 8594 17477 8696 17511
rect 8730 17477 8832 17511
rect 8866 17477 8968 17511
rect 9002 17477 9104 17511
rect 9138 17477 9240 17511
rect 7880 17375 9274 17477
rect 7914 17341 8016 17375
rect 8050 17341 8152 17375
rect 8186 17341 8288 17375
rect 8322 17341 8424 17375
rect 8458 17341 8560 17375
rect 8594 17341 8696 17375
rect 8730 17341 8832 17375
rect 8866 17341 8968 17375
rect 9002 17341 9104 17375
rect 9138 17341 9240 17375
rect 7880 17239 9274 17341
rect 7914 17205 8016 17239
rect 8050 17205 8152 17239
rect 8186 17205 8288 17239
rect 8322 17205 8424 17239
rect 8458 17205 8560 17239
rect 8594 17205 8696 17239
rect 8730 17205 8832 17239
rect 8866 17205 8968 17239
rect 9002 17205 9104 17239
rect 9138 17205 9240 17239
rect 7880 17103 9274 17205
rect 7914 17069 8016 17103
rect 8050 17069 8152 17103
rect 8186 17069 8288 17103
rect 8322 17069 8424 17103
rect 8458 17069 8560 17103
rect 8594 17069 8696 17103
rect 8730 17069 8832 17103
rect 8866 17069 8968 17103
rect 9002 17069 9104 17103
rect 9138 17069 9240 17103
rect 7880 16967 9274 17069
rect 7914 16933 8016 16967
rect 8050 16933 8152 16967
rect 8186 16933 8288 16967
rect 8322 16933 8424 16967
rect 8458 16933 8560 16967
rect 8594 16933 8696 16967
rect 8730 16933 8832 16967
rect 8866 16933 8968 16967
rect 9002 16933 9104 16967
rect 9138 16933 9240 16967
rect 7880 16831 9274 16933
rect 7914 16797 8016 16831
rect 8050 16797 8152 16831
rect 8186 16797 8288 16831
rect 8322 16797 8424 16831
rect 8458 16797 8560 16831
rect 8594 16797 8696 16831
rect 8730 16797 8832 16831
rect 8866 16797 8968 16831
rect 9002 16797 9104 16831
rect 9138 16797 9240 16831
rect 7880 16695 9274 16797
rect 7914 16661 8016 16695
rect 8050 16661 8152 16695
rect 8186 16661 8288 16695
rect 8322 16661 8424 16695
rect 8458 16661 8560 16695
rect 8594 16661 8696 16695
rect 8730 16661 8832 16695
rect 8866 16661 8968 16695
rect 9002 16661 9104 16695
rect 9138 16661 9240 16695
rect 7880 16559 9274 16661
rect 7914 16525 8016 16559
rect 8050 16525 8152 16559
rect 8186 16525 8288 16559
rect 8322 16525 8424 16559
rect 8458 16525 8560 16559
rect 8594 16525 8696 16559
rect 8730 16525 8832 16559
rect 8866 16525 8968 16559
rect 9002 16525 9104 16559
rect 9138 16525 9240 16559
rect 359 16389 461 16423
rect 495 16389 597 16423
rect 631 16389 733 16423
rect 767 16389 869 16423
rect 903 16389 1005 16423
rect 1039 16389 1141 16423
rect 1175 16389 1277 16423
rect 1311 16389 1413 16423
rect 1447 16389 1549 16423
rect 1583 16389 1685 16423
rect 325 16287 1719 16389
rect 359 16253 461 16287
rect 495 16253 597 16287
rect 631 16253 733 16287
rect 767 16253 869 16287
rect 903 16253 1005 16287
rect 1039 16253 1141 16287
rect 1175 16253 1277 16287
rect 1311 16253 1413 16287
rect 1447 16253 1549 16287
rect 1583 16253 1685 16287
rect 325 16151 1719 16253
rect 359 16117 461 16151
rect 495 16117 597 16151
rect 631 16117 733 16151
rect 767 16117 869 16151
rect 903 16117 1005 16151
rect 1039 16117 1141 16151
rect 1175 16117 1277 16151
rect 1311 16117 1413 16151
rect 1447 16117 1549 16151
rect 1583 16117 1685 16151
rect 325 16015 1719 16117
rect 359 15981 461 16015
rect 495 15981 597 16015
rect 631 15981 733 16015
rect 767 15981 869 16015
rect 903 15981 1005 16015
rect 1039 15981 1141 16015
rect 1175 15981 1277 16015
rect 1311 15981 1413 16015
rect 1447 15981 1549 16015
rect 1583 15981 1685 16015
rect 325 15879 1719 15981
rect 359 15845 461 15879
rect 495 15845 597 15879
rect 631 15845 733 15879
rect 767 15845 869 15879
rect 903 15845 1005 15879
rect 1039 15845 1141 15879
rect 1175 15845 1277 15879
rect 1311 15845 1413 15879
rect 1447 15845 1549 15879
rect 1583 15845 1685 15879
rect 325 15743 1719 15845
rect 359 15709 461 15743
rect 495 15709 597 15743
rect 631 15709 733 15743
rect 767 15709 869 15743
rect 903 15709 1005 15743
rect 1039 15709 1141 15743
rect 1175 15709 1277 15743
rect 1311 15709 1413 15743
rect 1447 15709 1549 15743
rect 1583 15709 1685 15743
rect 325 15607 1719 15709
rect 359 15573 461 15607
rect 495 15573 597 15607
rect 631 15573 733 15607
rect 767 15573 869 15607
rect 903 15573 1005 15607
rect 1039 15573 1141 15607
rect 1175 15573 1277 15607
rect 1311 15573 1413 15607
rect 1447 15573 1549 15607
rect 1583 15573 1685 15607
rect 325 15471 1719 15573
rect 359 15437 461 15471
rect 495 15437 597 15471
rect 631 15437 733 15471
rect 767 15437 869 15471
rect 903 15437 1005 15471
rect 1039 15437 1141 15471
rect 1175 15437 1277 15471
rect 1311 15437 1413 15471
rect 1447 15437 1549 15471
rect 1583 15437 1685 15471
rect 325 15335 1719 15437
rect 359 15301 461 15335
rect 495 15301 597 15335
rect 631 15301 733 15335
rect 767 15301 869 15335
rect 903 15301 1005 15335
rect 1039 15301 1141 15335
rect 1175 15301 1277 15335
rect 1311 15301 1413 15335
rect 1447 15301 1549 15335
rect 1583 15301 1685 15335
rect 325 15199 1719 15301
rect 359 15165 461 15199
rect 495 15165 597 15199
rect 631 15165 733 15199
rect 767 15165 869 15199
rect 903 15165 1005 15199
rect 1039 15165 1141 15199
rect 1175 15165 1277 15199
rect 1311 15165 1413 15199
rect 1447 15165 1549 15199
rect 1583 15165 1685 15199
rect 325 15063 1719 15165
rect 359 15029 461 15063
rect 495 15029 597 15063
rect 631 15029 733 15063
rect 767 15029 869 15063
rect 903 15029 1005 15063
rect 1039 15029 1141 15063
rect 1175 15029 1277 15063
rect 1311 15029 1413 15063
rect 1447 15029 1549 15063
rect 1583 15029 1685 15063
rect 325 14927 1719 15029
rect 359 14893 461 14927
rect 495 14893 597 14927
rect 631 14893 733 14927
rect 767 14893 869 14927
rect 903 14893 1005 14927
rect 1039 14893 1141 14927
rect 1175 14893 1277 14927
rect 1311 14893 1413 14927
rect 1447 14893 1549 14927
rect 1583 14893 1685 14927
rect 325 14791 1719 14893
rect 359 14757 461 14791
rect 495 14757 597 14791
rect 631 14757 733 14791
rect 767 14757 869 14791
rect 903 14757 1005 14791
rect 1039 14757 1141 14791
rect 1175 14757 1277 14791
rect 1311 14757 1413 14791
rect 1447 14757 1549 14791
rect 1583 14757 1685 14791
rect 325 14655 1719 14757
rect 359 14621 461 14655
rect 495 14621 597 14655
rect 631 14621 733 14655
rect 767 14621 869 14655
rect 903 14621 1005 14655
rect 1039 14621 1141 14655
rect 1175 14621 1277 14655
rect 1311 14621 1413 14655
rect 1447 14621 1549 14655
rect 1583 14621 1685 14655
rect 325 14519 1719 14621
rect 359 14485 461 14519
rect 495 14485 597 14519
rect 631 14485 733 14519
rect 767 14485 869 14519
rect 903 14485 1005 14519
rect 1039 14485 1141 14519
rect 1175 14485 1277 14519
rect 1311 14485 1413 14519
rect 1447 14485 1549 14519
rect 1583 14485 1685 14519
rect 325 14383 1719 14485
rect 359 14349 461 14383
rect 495 14349 597 14383
rect 631 14349 733 14383
rect 767 14349 869 14383
rect 903 14349 1005 14383
rect 1039 14349 1141 14383
rect 1175 14349 1277 14383
rect 1311 14349 1413 14383
rect 1447 14349 1549 14383
rect 1583 14349 1685 14383
rect 325 14247 1719 14349
rect 359 14213 461 14247
rect 495 14213 597 14247
rect 631 14213 733 14247
rect 767 14213 869 14247
rect 903 14213 1005 14247
rect 1039 14213 1141 14247
rect 1175 14213 1277 14247
rect 1311 14213 1413 14247
rect 1447 14213 1549 14247
rect 1583 14213 1685 14247
rect 325 14111 1719 14213
rect 359 14077 461 14111
rect 495 14077 597 14111
rect 631 14077 733 14111
rect 767 14077 869 14111
rect 903 14077 1005 14111
rect 1039 14077 1141 14111
rect 1175 14077 1277 14111
rect 1311 14077 1413 14111
rect 1447 14077 1549 14111
rect 1583 14077 1685 14111
rect 325 13975 1719 14077
rect 359 13941 461 13975
rect 495 13941 597 13975
rect 631 13941 733 13975
rect 767 13941 869 13975
rect 903 13941 1005 13975
rect 1039 13941 1141 13975
rect 1175 13941 1277 13975
rect 1311 13941 1413 13975
rect 1447 13941 1549 13975
rect 1583 13941 1685 13975
rect 325 13839 1719 13941
rect 359 13805 461 13839
rect 495 13805 597 13839
rect 631 13805 733 13839
rect 767 13805 869 13839
rect 903 13805 1005 13839
rect 1039 13805 1141 13839
rect 1175 13805 1277 13839
rect 1311 13805 1413 13839
rect 1447 13805 1549 13839
rect 1583 13805 1685 13839
rect 325 13703 1719 13805
rect 359 13669 461 13703
rect 495 13669 597 13703
rect 631 13669 733 13703
rect 767 13669 869 13703
rect 903 13669 1005 13703
rect 1039 13669 1141 13703
rect 1175 13669 1277 13703
rect 1311 13669 1413 13703
rect 1447 13669 1549 13703
rect 1583 13669 1685 13703
rect 325 13567 1719 13669
rect 359 13533 461 13567
rect 495 13533 597 13567
rect 631 13533 733 13567
rect 767 13533 869 13567
rect 903 13533 1005 13567
rect 1039 13533 1141 13567
rect 1175 13533 1277 13567
rect 1311 13533 1413 13567
rect 1447 13533 1549 13567
rect 1583 13533 1685 13567
rect 325 13431 1719 13533
rect 359 13397 461 13431
rect 495 13397 597 13431
rect 631 13397 733 13431
rect 767 13397 869 13431
rect 903 13397 1005 13431
rect 1039 13397 1141 13431
rect 1175 13397 1277 13431
rect 1311 13397 1413 13431
rect 1447 13397 1549 13431
rect 1583 13397 1685 13431
rect 325 13295 1719 13397
rect 359 13261 461 13295
rect 495 13261 597 13295
rect 631 13261 733 13295
rect 767 13261 869 13295
rect 903 13261 1005 13295
rect 1039 13261 1141 13295
rect 1175 13261 1277 13295
rect 1311 13261 1413 13295
rect 1447 13261 1549 13295
rect 1583 13261 1685 13295
rect 325 13159 1719 13261
rect 359 13125 461 13159
rect 495 13125 597 13159
rect 631 13125 733 13159
rect 767 13125 869 13159
rect 903 13125 1005 13159
rect 1039 13125 1141 13159
rect 1175 13125 1277 13159
rect 1311 13125 1413 13159
rect 1447 13125 1549 13159
rect 1583 13125 1685 13159
rect 325 13023 1719 13125
rect 359 12989 461 13023
rect 495 12989 597 13023
rect 631 12989 733 13023
rect 767 12989 869 13023
rect 903 12989 1005 13023
rect 1039 12989 1141 13023
rect 1175 12989 1277 13023
rect 1311 12989 1413 13023
rect 1447 12989 1549 13023
rect 1583 12989 1685 13023
rect 325 12887 1719 12989
rect 359 12853 461 12887
rect 495 12853 597 12887
rect 631 12853 733 12887
rect 767 12853 869 12887
rect 903 12853 1005 12887
rect 1039 12853 1141 12887
rect 1175 12853 1277 12887
rect 1311 12853 1413 12887
rect 1447 12853 1549 12887
rect 1583 12853 1685 12887
rect 325 12751 1719 12853
rect 359 12717 461 12751
rect 495 12717 597 12751
rect 631 12717 733 12751
rect 767 12717 869 12751
rect 903 12717 1005 12751
rect 1039 12717 1141 12751
rect 1175 12717 1277 12751
rect 1311 12717 1413 12751
rect 1447 12717 1549 12751
rect 1583 12717 1685 12751
rect 325 12615 1719 12717
rect 359 12581 461 12615
rect 495 12581 597 12615
rect 631 12581 733 12615
rect 767 12581 869 12615
rect 903 12581 1005 12615
rect 1039 12581 1141 12615
rect 1175 12581 1277 12615
rect 1311 12581 1413 12615
rect 1447 12581 1549 12615
rect 1583 12581 1685 12615
rect 325 12479 1719 12581
rect 359 12445 461 12479
rect 495 12445 597 12479
rect 631 12445 733 12479
rect 767 12445 869 12479
rect 903 12445 1005 12479
rect 1039 12445 1141 12479
rect 1175 12445 1277 12479
rect 1311 12445 1413 12479
rect 1447 12445 1549 12479
rect 1583 12445 1685 12479
rect 325 12343 1719 12445
rect 359 12309 461 12343
rect 495 12309 597 12343
rect 631 12309 733 12343
rect 767 12309 869 12343
rect 903 12309 1005 12343
rect 1039 12309 1141 12343
rect 1175 12309 1277 12343
rect 1311 12309 1413 12343
rect 1447 12309 1549 12343
rect 1583 12309 1685 12343
rect 325 12207 1719 12309
rect 359 12173 461 12207
rect 495 12173 597 12207
rect 631 12173 733 12207
rect 767 12173 869 12207
rect 903 12173 1005 12207
rect 1039 12173 1141 12207
rect 1175 12173 1277 12207
rect 1311 12173 1413 12207
rect 1447 12173 1549 12207
rect 1583 12173 1685 12207
rect 325 12071 1719 12173
rect 359 12037 461 12071
rect 495 12037 597 12071
rect 631 12037 733 12071
rect 767 12037 869 12071
rect 903 12037 1005 12071
rect 1039 12037 1141 12071
rect 1175 12037 1277 12071
rect 1311 12037 1413 12071
rect 1447 12037 1549 12071
rect 1583 12037 1685 12071
rect 325 11935 1719 12037
rect 359 11901 461 11935
rect 495 11901 597 11935
rect 631 11901 733 11935
rect 767 11901 869 11935
rect 903 11901 1005 11935
rect 1039 11901 1141 11935
rect 1175 11901 1277 11935
rect 1311 11901 1413 11935
rect 1447 11901 1549 11935
rect 1583 11901 1685 11935
rect 325 11799 1719 11901
rect 359 11765 461 11799
rect 495 11765 597 11799
rect 631 11765 733 11799
rect 767 11765 869 11799
rect 903 11765 1005 11799
rect 1039 11765 1141 11799
rect 1175 11765 1277 11799
rect 1311 11765 1413 11799
rect 1447 11765 1549 11799
rect 1583 11765 1685 11799
rect 325 11663 1719 11765
rect 359 11629 461 11663
rect 495 11629 597 11663
rect 631 11629 733 11663
rect 767 11629 869 11663
rect 903 11629 1005 11663
rect 1039 11629 1141 11663
rect 1175 11629 1277 11663
rect 1311 11629 1413 11663
rect 1447 11629 1549 11663
rect 1583 11629 1685 11663
rect 325 11527 1719 11629
rect 359 11493 461 11527
rect 495 11493 597 11527
rect 631 11493 733 11527
rect 767 11493 869 11527
rect 903 11493 1005 11527
rect 1039 11493 1141 11527
rect 1175 11493 1277 11527
rect 1311 11493 1413 11527
rect 1447 11493 1549 11527
rect 1583 11493 1685 11527
rect 325 11391 1719 11493
rect 359 11357 461 11391
rect 495 11357 597 11391
rect 631 11357 733 11391
rect 767 11357 869 11391
rect 903 11357 1005 11391
rect 1039 11357 1141 11391
rect 1175 11357 1277 11391
rect 1311 11357 1413 11391
rect 1447 11357 1549 11391
rect 1583 11357 1685 11391
rect 325 11255 1719 11357
rect 359 11221 461 11255
rect 495 11221 597 11255
rect 631 11221 733 11255
rect 767 11221 869 11255
rect 903 11221 1005 11255
rect 1039 11221 1141 11255
rect 1175 11221 1277 11255
rect 1311 11221 1413 11255
rect 1447 11221 1549 11255
rect 1583 11221 1685 11255
rect 325 11119 1719 11221
rect 359 11085 461 11119
rect 495 11085 597 11119
rect 631 11085 733 11119
rect 767 11085 869 11119
rect 903 11085 1005 11119
rect 1039 11085 1141 11119
rect 1175 11085 1277 11119
rect 1311 11085 1413 11119
rect 1447 11085 1549 11119
rect 1583 11085 1685 11119
rect 325 10983 1719 11085
rect 359 10949 461 10983
rect 495 10949 597 10983
rect 631 10949 733 10983
rect 767 10949 869 10983
rect 903 10949 1005 10983
rect 1039 10949 1141 10983
rect 1175 10949 1277 10983
rect 1311 10949 1413 10983
rect 1447 10949 1549 10983
rect 1583 10949 1685 10983
rect 325 10847 1719 10949
rect 359 10813 461 10847
rect 495 10813 597 10847
rect 631 10813 733 10847
rect 767 10813 869 10847
rect 903 10813 1005 10847
rect 1039 10813 1141 10847
rect 1175 10813 1277 10847
rect 1311 10813 1413 10847
rect 1447 10813 1549 10847
rect 1583 10813 1685 10847
rect 325 10711 1719 10813
rect 359 10677 461 10711
rect 495 10677 597 10711
rect 631 10677 733 10711
rect 767 10677 869 10711
rect 903 10677 1005 10711
rect 1039 10677 1141 10711
rect 1175 10677 1277 10711
rect 1311 10677 1413 10711
rect 1447 10677 1549 10711
rect 1583 10677 1685 10711
rect 325 10575 1719 10677
rect 359 10541 461 10575
rect 495 10541 597 10575
rect 631 10541 733 10575
rect 767 10541 869 10575
rect 903 10541 1005 10575
rect 1039 10541 1141 10575
rect 1175 10541 1277 10575
rect 1311 10541 1413 10575
rect 1447 10541 1549 10575
rect 1583 10541 1685 10575
rect 325 10439 1719 10541
rect 359 10405 461 10439
rect 495 10405 597 10439
rect 631 10405 733 10439
rect 767 10405 869 10439
rect 903 10405 1005 10439
rect 1039 10405 1141 10439
rect 1175 10405 1277 10439
rect 1311 10405 1413 10439
rect 1447 10405 1549 10439
rect 1583 10405 1685 10439
rect 325 10303 1719 10405
rect 359 10269 461 10303
rect 495 10269 597 10303
rect 631 10269 733 10303
rect 767 10269 869 10303
rect 903 10269 1005 10303
rect 1039 10269 1141 10303
rect 1175 10269 1277 10303
rect 1311 10269 1413 10303
rect 1447 10269 1549 10303
rect 1583 10269 1685 10303
rect 325 10167 1719 10269
rect 359 10133 461 10167
rect 495 10133 597 10167
rect 631 10133 733 10167
rect 767 10133 869 10167
rect 903 10133 1005 10167
rect 1039 10133 1141 10167
rect 1175 10133 1277 10167
rect 1311 10133 1413 10167
rect 1447 10133 1549 10167
rect 1583 10133 1685 10167
rect 325 10031 1719 10133
rect 359 9997 461 10031
rect 495 9997 597 10031
rect 631 9997 733 10031
rect 767 9997 869 10031
rect 903 9997 1005 10031
rect 1039 9997 1141 10031
rect 1175 9997 1277 10031
rect 1311 9997 1413 10031
rect 1447 9997 1549 10031
rect 1583 9997 1685 10031
rect 325 9895 1719 9997
rect 359 9861 461 9895
rect 495 9861 597 9895
rect 631 9861 733 9895
rect 767 9861 869 9895
rect 903 9861 1005 9895
rect 1039 9861 1141 9895
rect 1175 9861 1277 9895
rect 1311 9861 1413 9895
rect 1447 9861 1549 9895
rect 1583 9861 1685 9895
rect 325 9759 1719 9861
rect 359 9725 461 9759
rect 495 9725 597 9759
rect 631 9725 733 9759
rect 767 9725 869 9759
rect 903 9725 1005 9759
rect 1039 9725 1141 9759
rect 1175 9725 1277 9759
rect 1311 9725 1413 9759
rect 1447 9725 1549 9759
rect 1583 9725 1685 9759
rect 325 9623 1719 9725
rect 359 9589 461 9623
rect 495 9589 597 9623
rect 631 9589 733 9623
rect 767 9589 869 9623
rect 903 9589 1005 9623
rect 1039 9589 1141 9623
rect 1175 9589 1277 9623
rect 1311 9589 1413 9623
rect 1447 9589 1549 9623
rect 1583 9589 1685 9623
rect 325 9487 1719 9589
rect 359 9453 461 9487
rect 495 9453 597 9487
rect 631 9453 733 9487
rect 767 9453 869 9487
rect 903 9453 1005 9487
rect 1039 9453 1141 9487
rect 1175 9453 1277 9487
rect 1311 9453 1413 9487
rect 1447 9453 1549 9487
rect 1583 9453 1685 9487
rect 325 9351 1719 9453
rect 359 9317 461 9351
rect 495 9317 597 9351
rect 631 9317 733 9351
rect 767 9317 869 9351
rect 903 9317 1005 9351
rect 1039 9317 1141 9351
rect 1175 9317 1277 9351
rect 1311 9317 1413 9351
rect 1447 9317 1549 9351
rect 1583 9317 1685 9351
rect 325 9215 1719 9317
rect 359 9181 461 9215
rect 495 9181 597 9215
rect 631 9181 733 9215
rect 767 9181 869 9215
rect 903 9181 1005 9215
rect 1039 9181 1141 9215
rect 1175 9181 1277 9215
rect 1311 9181 1413 9215
rect 1447 9181 1549 9215
rect 1583 9181 1685 9215
rect 325 9079 1719 9181
rect 359 9045 461 9079
rect 495 9045 597 9079
rect 631 9045 733 9079
rect 767 9045 869 9079
rect 903 9045 1005 9079
rect 1039 9045 1141 9079
rect 1175 9045 1277 9079
rect 1311 9045 1413 9079
rect 1447 9045 1549 9079
rect 1583 9045 1685 9079
rect 325 8943 1719 9045
rect 359 8909 461 8943
rect 495 8909 597 8943
rect 631 8909 733 8943
rect 767 8909 869 8943
rect 903 8909 1005 8943
rect 1039 8909 1141 8943
rect 1175 8909 1277 8943
rect 1311 8909 1413 8943
rect 1447 8909 1549 8943
rect 1583 8909 1685 8943
rect 325 8807 1719 8909
rect 359 8773 461 8807
rect 495 8773 597 8807
rect 631 8773 733 8807
rect 767 8773 869 8807
rect 903 8773 1005 8807
rect 1039 8773 1141 8807
rect 1175 8773 1277 8807
rect 1311 8773 1413 8807
rect 1447 8773 1549 8807
rect 1583 8773 1685 8807
rect 325 8671 1719 8773
rect 359 8637 461 8671
rect 495 8637 597 8671
rect 631 8637 733 8671
rect 767 8637 869 8671
rect 903 8637 1005 8671
rect 1039 8637 1141 8671
rect 1175 8637 1277 8671
rect 1311 8637 1413 8671
rect 1447 8637 1549 8671
rect 1583 8637 1685 8671
rect 325 8535 1719 8637
rect 359 8501 461 8535
rect 495 8501 597 8535
rect 631 8501 733 8535
rect 767 8501 869 8535
rect 903 8501 1005 8535
rect 1039 8501 1141 8535
rect 1175 8501 1277 8535
rect 1311 8501 1413 8535
rect 1447 8501 1549 8535
rect 1583 8501 1685 8535
rect 325 8399 1719 8501
rect 359 8365 461 8399
rect 495 8365 597 8399
rect 631 8365 733 8399
rect 767 8365 869 8399
rect 903 8365 1005 8399
rect 1039 8365 1141 8399
rect 1175 8365 1277 8399
rect 1311 8365 1413 8399
rect 1447 8365 1549 8399
rect 1583 8365 1685 8399
rect 325 8263 1719 8365
rect 359 8229 461 8263
rect 495 8229 597 8263
rect 631 8229 733 8263
rect 767 8229 869 8263
rect 903 8229 1005 8263
rect 1039 8229 1141 8263
rect 1175 8229 1277 8263
rect 1311 8229 1413 8263
rect 1447 8229 1549 8263
rect 1583 8229 1685 8263
rect 325 8127 1719 8229
rect 359 8093 461 8127
rect 495 8093 597 8127
rect 631 8093 733 8127
rect 767 8093 869 8127
rect 903 8093 1005 8127
rect 1039 8093 1141 8127
rect 1175 8093 1277 8127
rect 1311 8093 1413 8127
rect 1447 8093 1549 8127
rect 1583 8093 1685 8127
rect 325 7991 1719 8093
rect 359 7957 461 7991
rect 495 7957 597 7991
rect 631 7957 733 7991
rect 767 7957 869 7991
rect 903 7957 1005 7991
rect 1039 7957 1141 7991
rect 1175 7957 1277 7991
rect 1311 7957 1413 7991
rect 1447 7957 1549 7991
rect 1583 7957 1685 7991
rect 325 7855 1719 7957
rect 359 7821 461 7855
rect 495 7821 597 7855
rect 631 7821 733 7855
rect 767 7821 869 7855
rect 903 7821 1005 7855
rect 1039 7821 1141 7855
rect 1175 7821 1277 7855
rect 1311 7821 1413 7855
rect 1447 7821 1549 7855
rect 1583 7821 1685 7855
rect 325 7719 1719 7821
rect 359 7685 461 7719
rect 495 7685 597 7719
rect 631 7685 733 7719
rect 767 7685 869 7719
rect 903 7685 1005 7719
rect 1039 7685 1141 7719
rect 1175 7685 1277 7719
rect 1311 7685 1413 7719
rect 1447 7685 1549 7719
rect 1583 7685 1685 7719
rect 325 7583 1719 7685
rect 359 7549 461 7583
rect 495 7549 597 7583
rect 631 7549 733 7583
rect 767 7549 869 7583
rect 903 7549 1005 7583
rect 1039 7549 1141 7583
rect 1175 7549 1277 7583
rect 1311 7549 1413 7583
rect 1447 7549 1549 7583
rect 1583 7549 1685 7583
rect 325 7447 1719 7549
rect 359 7413 461 7447
rect 495 7413 597 7447
rect 631 7413 733 7447
rect 767 7413 869 7447
rect 903 7413 1005 7447
rect 1039 7413 1141 7447
rect 1175 7413 1277 7447
rect 1311 7413 1413 7447
rect 1447 7413 1549 7447
rect 1583 7413 1685 7447
rect 325 7311 1719 7413
rect 359 7277 461 7311
rect 495 7277 597 7311
rect 631 7277 733 7311
rect 767 7277 869 7311
rect 903 7277 1005 7311
rect 1039 7277 1141 7311
rect 1175 7277 1277 7311
rect 1311 7277 1413 7311
rect 1447 7277 1549 7311
rect 1583 7277 1685 7311
rect 325 7175 1719 7277
rect 359 7141 461 7175
rect 495 7141 597 7175
rect 631 7141 733 7175
rect 767 7141 869 7175
rect 903 7141 1005 7175
rect 1039 7141 1141 7175
rect 1175 7141 1277 7175
rect 1311 7141 1413 7175
rect 1447 7141 1549 7175
rect 1583 7141 1685 7175
rect 325 7039 1719 7141
rect 359 7005 461 7039
rect 495 7005 597 7039
rect 631 7005 733 7039
rect 767 7005 869 7039
rect 903 7005 1005 7039
rect 1039 7005 1141 7039
rect 1175 7005 1277 7039
rect 1311 7005 1413 7039
rect 1447 7005 1549 7039
rect 1583 7005 1685 7039
rect 325 6903 1719 7005
rect 359 6869 461 6903
rect 495 6869 597 6903
rect 631 6869 733 6903
rect 767 6869 869 6903
rect 903 6869 1005 6903
rect 1039 6869 1141 6903
rect 1175 6869 1277 6903
rect 1311 6869 1413 6903
rect 1447 6869 1549 6903
rect 1583 6869 1685 6903
rect 325 6767 1719 6869
rect 359 6733 461 6767
rect 495 6733 597 6767
rect 631 6733 733 6767
rect 767 6733 869 6767
rect 903 6733 1005 6767
rect 1039 6733 1141 6767
rect 1175 6733 1277 6767
rect 1311 6733 1413 6767
rect 1447 6733 1549 6767
rect 1583 6733 1685 6767
rect 325 6631 1719 6733
rect 359 6597 461 6631
rect 495 6597 597 6631
rect 631 6597 733 6631
rect 767 6597 869 6631
rect 903 6597 1005 6631
rect 1039 6597 1141 6631
rect 1175 6597 1277 6631
rect 1311 6597 1413 6631
rect 1447 6597 1549 6631
rect 1583 6597 1685 6631
rect 325 6495 1719 6597
rect 359 6461 461 6495
rect 495 6461 597 6495
rect 631 6461 733 6495
rect 767 6461 869 6495
rect 903 6461 1005 6495
rect 1039 6461 1141 6495
rect 1175 6461 1277 6495
rect 1311 6461 1413 6495
rect 1447 6461 1549 6495
rect 1583 6461 1685 6495
rect 325 6359 1719 6461
rect 359 6325 461 6359
rect 495 6325 597 6359
rect 631 6325 733 6359
rect 767 6325 869 6359
rect 903 6325 1005 6359
rect 1039 6325 1141 6359
rect 1175 6325 1277 6359
rect 1311 6325 1413 6359
rect 1447 6325 1549 6359
rect 1583 6325 1685 6359
rect 325 6223 1719 6325
rect 359 6189 461 6223
rect 495 6189 597 6223
rect 631 6189 733 6223
rect 767 6189 869 6223
rect 903 6189 1005 6223
rect 1039 6189 1141 6223
rect 1175 6189 1277 6223
rect 1311 6189 1413 6223
rect 1447 6189 1549 6223
rect 1583 6189 1685 6223
rect 325 6087 1719 6189
rect 359 6053 461 6087
rect 495 6053 597 6087
rect 631 6053 733 6087
rect 767 6053 869 6087
rect 903 6053 1005 6087
rect 1039 6053 1141 6087
rect 1175 6053 1277 6087
rect 1311 6053 1413 6087
rect 1447 6053 1549 6087
rect 1583 6053 1685 6087
rect 325 5951 1719 6053
rect 359 5917 461 5951
rect 495 5917 597 5951
rect 631 5917 733 5951
rect 767 5917 869 5951
rect 903 5917 1005 5951
rect 1039 5917 1141 5951
rect 1175 5917 1277 5951
rect 1311 5917 1413 5951
rect 1447 5917 1549 5951
rect 1583 5917 1685 5951
rect 325 5815 1719 5917
rect 359 5781 461 5815
rect 495 5781 597 5815
rect 631 5781 733 5815
rect 767 5781 869 5815
rect 903 5781 1005 5815
rect 1039 5781 1141 5815
rect 1175 5781 1277 5815
rect 1311 5781 1413 5815
rect 1447 5781 1549 5815
rect 1583 5781 1685 5815
rect 325 5679 1719 5781
rect 359 5645 461 5679
rect 495 5645 597 5679
rect 631 5645 733 5679
rect 767 5645 869 5679
rect 903 5645 1005 5679
rect 1039 5645 1141 5679
rect 1175 5645 1277 5679
rect 1311 5645 1413 5679
rect 1447 5645 1549 5679
rect 1583 5645 1685 5679
rect 325 5543 1719 5645
rect 359 5509 461 5543
rect 495 5509 597 5543
rect 631 5509 733 5543
rect 767 5509 869 5543
rect 903 5509 1005 5543
rect 1039 5509 1141 5543
rect 1175 5509 1277 5543
rect 1311 5509 1413 5543
rect 1447 5509 1549 5543
rect 1583 5509 1685 5543
rect 325 5407 1719 5509
rect 359 5373 461 5407
rect 495 5373 597 5407
rect 631 5373 733 5407
rect 767 5373 869 5407
rect 903 5373 1005 5407
rect 1039 5373 1141 5407
rect 1175 5373 1277 5407
rect 1311 5373 1413 5407
rect 1447 5373 1549 5407
rect 1583 5373 1685 5407
rect 325 5271 1719 5373
rect 359 5237 461 5271
rect 495 5237 597 5271
rect 631 5237 733 5271
rect 767 5237 869 5271
rect 903 5237 1005 5271
rect 1039 5237 1141 5271
rect 1175 5237 1277 5271
rect 1311 5237 1413 5271
rect 1447 5237 1549 5271
rect 1583 5237 1685 5271
rect 325 5135 1719 5237
rect 359 5101 461 5135
rect 495 5101 597 5135
rect 631 5101 733 5135
rect 767 5101 869 5135
rect 903 5101 1005 5135
rect 1039 5101 1141 5135
rect 1175 5101 1277 5135
rect 1311 5101 1413 5135
rect 1447 5101 1549 5135
rect 1583 5101 1685 5135
rect 325 4999 1719 5101
rect 359 4965 461 4999
rect 495 4965 597 4999
rect 631 4965 733 4999
rect 767 4965 869 4999
rect 903 4965 1005 4999
rect 1039 4965 1141 4999
rect 1175 4965 1277 4999
rect 1311 4965 1413 4999
rect 1447 4965 1549 4999
rect 1583 4965 1685 4999
rect 325 4863 1719 4965
rect 359 4829 461 4863
rect 495 4829 597 4863
rect 631 4829 733 4863
rect 767 4829 869 4863
rect 903 4829 1005 4863
rect 1039 4829 1141 4863
rect 1175 4829 1277 4863
rect 1311 4829 1413 4863
rect 1447 4829 1549 4863
rect 1583 4829 1685 4863
rect 325 4727 1719 4829
rect 359 4693 461 4727
rect 495 4693 597 4727
rect 631 4693 733 4727
rect 767 4693 869 4727
rect 903 4693 1005 4727
rect 1039 4693 1141 4727
rect 1175 4693 1277 4727
rect 1311 4693 1413 4727
rect 1447 4693 1549 4727
rect 1583 4693 1685 4727
rect 325 4591 1719 4693
rect 359 4557 461 4591
rect 495 4557 597 4591
rect 631 4557 733 4591
rect 767 4557 869 4591
rect 903 4557 1005 4591
rect 1039 4557 1141 4591
rect 1175 4557 1277 4591
rect 1311 4557 1413 4591
rect 1447 4557 1549 4591
rect 1583 4557 1685 4591
rect 325 4455 1719 4557
rect 359 4421 461 4455
rect 495 4421 597 4455
rect 631 4421 733 4455
rect 767 4421 869 4455
rect 903 4421 1005 4455
rect 1039 4421 1141 4455
rect 1175 4421 1277 4455
rect 1311 4421 1413 4455
rect 1447 4421 1549 4455
rect 1583 4421 1685 4455
rect 325 4319 1719 4421
rect 359 4285 461 4319
rect 495 4285 597 4319
rect 631 4285 733 4319
rect 767 4285 869 4319
rect 903 4285 1005 4319
rect 1039 4285 1141 4319
rect 1175 4285 1277 4319
rect 1311 4285 1413 4319
rect 1447 4285 1549 4319
rect 1583 4285 1685 4319
rect 325 4183 1719 4285
rect 359 4149 461 4183
rect 495 4149 597 4183
rect 631 4149 733 4183
rect 767 4149 869 4183
rect 903 4149 1005 4183
rect 1039 4149 1141 4183
rect 1175 4149 1277 4183
rect 1311 4149 1413 4183
rect 1447 4149 1549 4183
rect 1583 4149 1685 4183
rect 325 4047 1719 4149
rect 359 4013 461 4047
rect 495 4013 597 4047
rect 631 4013 733 4047
rect 767 4013 869 4047
rect 903 4013 1005 4047
rect 1039 4013 1141 4047
rect 1175 4013 1277 4047
rect 1311 4013 1413 4047
rect 1447 4013 1549 4047
rect 1583 4013 1685 4047
rect 325 3911 1719 4013
rect 359 3877 461 3911
rect 495 3877 597 3911
rect 631 3877 733 3911
rect 767 3877 869 3911
rect 903 3877 1005 3911
rect 1039 3877 1141 3911
rect 1175 3877 1277 3911
rect 1311 3877 1413 3911
rect 1447 3877 1549 3911
rect 1583 3877 1685 3911
rect 325 3775 1719 3877
rect 359 3741 461 3775
rect 495 3741 597 3775
rect 631 3741 733 3775
rect 767 3741 869 3775
rect 903 3741 1005 3775
rect 1039 3741 1141 3775
rect 1175 3741 1277 3775
rect 1311 3741 1413 3775
rect 1447 3741 1549 3775
rect 1583 3741 1685 3775
rect 325 3639 1719 3741
rect 359 3605 461 3639
rect 495 3605 597 3639
rect 631 3605 733 3639
rect 767 3605 869 3639
rect 903 3605 1005 3639
rect 1039 3605 1141 3639
rect 1175 3605 1277 3639
rect 1311 3605 1413 3639
rect 1447 3605 1549 3639
rect 1583 3605 1685 3639
rect 325 3503 1719 3605
rect 359 3469 461 3503
rect 495 3469 597 3503
rect 631 3469 733 3503
rect 767 3469 869 3503
rect 903 3469 1005 3503
rect 1039 3469 1141 3503
rect 1175 3469 1277 3503
rect 1311 3469 1413 3503
rect 1447 3469 1549 3503
rect 1583 3469 1685 3503
rect 325 3367 1719 3469
rect 359 3333 461 3367
rect 495 3333 597 3367
rect 631 3333 733 3367
rect 767 3333 869 3367
rect 903 3333 1005 3367
rect 1039 3333 1141 3367
rect 1175 3333 1277 3367
rect 1311 3333 1413 3367
rect 1447 3333 1549 3367
rect 1583 3333 1685 3367
rect 325 3231 1719 3333
rect 359 3197 461 3231
rect 495 3197 597 3231
rect 631 3197 733 3231
rect 767 3197 869 3231
rect 903 3197 1005 3231
rect 1039 3197 1141 3231
rect 1175 3197 1277 3231
rect 1311 3197 1413 3231
rect 1447 3197 1549 3231
rect 1583 3197 1685 3231
rect 325 3095 1719 3197
rect 359 3061 461 3095
rect 495 3061 597 3095
rect 631 3061 733 3095
rect 767 3061 869 3095
rect 903 3061 1005 3095
rect 1039 3061 1141 3095
rect 1175 3061 1277 3095
rect 1311 3061 1413 3095
rect 1447 3061 1549 3095
rect 1583 3061 1685 3095
rect 325 2959 1719 3061
rect 359 2925 461 2959
rect 495 2925 597 2959
rect 631 2925 733 2959
rect 767 2925 869 2959
rect 903 2925 1005 2959
rect 1039 2925 1141 2959
rect 1175 2925 1277 2959
rect 1311 2925 1413 2959
rect 1447 2925 1549 2959
rect 1583 2925 1685 2959
rect 325 2823 1719 2925
rect 359 2789 461 2823
rect 495 2789 597 2823
rect 631 2789 733 2823
rect 767 2789 869 2823
rect 903 2789 1005 2823
rect 1039 2789 1141 2823
rect 1175 2789 1277 2823
rect 1311 2789 1413 2823
rect 1447 2789 1549 2823
rect 1583 2789 1685 2823
rect 325 2687 1719 2789
rect 359 2653 461 2687
rect 495 2653 597 2687
rect 631 2653 733 2687
rect 767 2653 869 2687
rect 903 2653 1005 2687
rect 1039 2653 1141 2687
rect 1175 2653 1277 2687
rect 1311 2653 1413 2687
rect 1447 2653 1549 2687
rect 1583 2653 1685 2687
rect 325 2551 1719 2653
rect 359 2517 461 2551
rect 495 2517 597 2551
rect 631 2517 733 2551
rect 767 2517 869 2551
rect 903 2517 1005 2551
rect 1039 2517 1141 2551
rect 1175 2517 1277 2551
rect 1311 2517 1413 2551
rect 1447 2517 1549 2551
rect 1583 2517 1685 2551
rect 325 2414 1719 2517
rect 359 2380 461 2414
rect 495 2380 597 2414
rect 631 2380 733 2414
rect 767 2380 869 2414
rect 903 2380 1005 2414
rect 1039 2380 1141 2414
rect 1175 2380 1277 2414
rect 1311 2380 1413 2414
rect 1447 2380 1549 2414
rect 1583 2380 1685 2414
rect 325 2277 1719 2380
rect 359 2243 461 2277
rect 495 2243 597 2277
rect 631 2243 733 2277
rect 767 2243 869 2277
rect 903 2243 1005 2277
rect 1039 2243 1141 2277
rect 1175 2243 1277 2277
rect 1311 2243 1413 2277
rect 1447 2243 1549 2277
rect 1583 2243 1685 2277
rect 325 2140 1719 2243
rect 359 2106 461 2140
rect 495 2106 597 2140
rect 631 2106 733 2140
rect 767 2106 869 2140
rect 903 2106 1005 2140
rect 1039 2106 1141 2140
rect 1175 2106 1277 2140
rect 1311 2106 1413 2140
rect 1447 2106 1549 2140
rect 1583 2106 1685 2140
rect 325 2003 1719 2106
rect 359 1969 461 2003
rect 495 1969 597 2003
rect 631 1969 733 2003
rect 767 1969 869 2003
rect 903 1969 1005 2003
rect 1039 1969 1141 2003
rect 1175 1969 1277 2003
rect 1311 1969 1413 2003
rect 1447 1969 1549 2003
rect 1583 1969 1685 2003
rect 325 1866 1719 1969
rect 359 1832 461 1866
rect 495 1832 597 1866
rect 631 1832 733 1866
rect 767 1832 869 1866
rect 903 1832 1005 1866
rect 1039 1832 1141 1866
rect 1175 1832 1277 1866
rect 1311 1832 1413 1866
rect 1447 1832 1549 1866
rect 1583 1832 1685 1866
rect 325 1729 1719 1832
rect 7880 16423 9274 16525
rect 7914 16389 8016 16423
rect 8050 16389 8152 16423
rect 8186 16389 8288 16423
rect 8322 16389 8424 16423
rect 8458 16389 8560 16423
rect 8594 16389 8696 16423
rect 8730 16389 8832 16423
rect 8866 16389 8968 16423
rect 9002 16389 9104 16423
rect 9138 16389 9240 16423
rect 7880 16287 9274 16389
rect 7914 16253 8016 16287
rect 8050 16253 8152 16287
rect 8186 16253 8288 16287
rect 8322 16253 8424 16287
rect 8458 16253 8560 16287
rect 8594 16253 8696 16287
rect 8730 16253 8832 16287
rect 8866 16253 8968 16287
rect 9002 16253 9104 16287
rect 9138 16253 9240 16287
rect 7880 16151 9274 16253
rect 7914 16117 8016 16151
rect 8050 16117 8152 16151
rect 8186 16117 8288 16151
rect 8322 16117 8424 16151
rect 8458 16117 8560 16151
rect 8594 16117 8696 16151
rect 8730 16117 8832 16151
rect 8866 16117 8968 16151
rect 9002 16117 9104 16151
rect 9138 16117 9240 16151
rect 7880 16015 9274 16117
rect 7914 15981 8016 16015
rect 8050 15981 8152 16015
rect 8186 15981 8288 16015
rect 8322 15981 8424 16015
rect 8458 15981 8560 16015
rect 8594 15981 8696 16015
rect 8730 15981 8832 16015
rect 8866 15981 8968 16015
rect 9002 15981 9104 16015
rect 9138 15981 9240 16015
rect 7880 15879 9274 15981
rect 7914 15845 8016 15879
rect 8050 15845 8152 15879
rect 8186 15845 8288 15879
rect 8322 15845 8424 15879
rect 8458 15845 8560 15879
rect 8594 15845 8696 15879
rect 8730 15845 8832 15879
rect 8866 15845 8968 15879
rect 9002 15845 9104 15879
rect 9138 15845 9240 15879
rect 7880 15743 9274 15845
rect 7914 15709 8016 15743
rect 8050 15709 8152 15743
rect 8186 15709 8288 15743
rect 8322 15709 8424 15743
rect 8458 15709 8560 15743
rect 8594 15709 8696 15743
rect 8730 15709 8832 15743
rect 8866 15709 8968 15743
rect 9002 15709 9104 15743
rect 9138 15709 9240 15743
rect 7880 15607 9274 15709
rect 7914 15573 8016 15607
rect 8050 15573 8152 15607
rect 8186 15573 8288 15607
rect 8322 15573 8424 15607
rect 8458 15573 8560 15607
rect 8594 15573 8696 15607
rect 8730 15573 8832 15607
rect 8866 15573 8968 15607
rect 9002 15573 9104 15607
rect 9138 15573 9240 15607
rect 7880 15471 9274 15573
rect 7914 15437 8016 15471
rect 8050 15437 8152 15471
rect 8186 15437 8288 15471
rect 8322 15437 8424 15471
rect 8458 15437 8560 15471
rect 8594 15437 8696 15471
rect 8730 15437 8832 15471
rect 8866 15437 8968 15471
rect 9002 15437 9104 15471
rect 9138 15437 9240 15471
rect 7880 15335 9274 15437
rect 7914 15301 8016 15335
rect 8050 15301 8152 15335
rect 8186 15301 8288 15335
rect 8322 15301 8424 15335
rect 8458 15301 8560 15335
rect 8594 15301 8696 15335
rect 8730 15301 8832 15335
rect 8866 15301 8968 15335
rect 9002 15301 9104 15335
rect 9138 15301 9240 15335
rect 7880 15199 9274 15301
rect 7914 15165 8016 15199
rect 8050 15165 8152 15199
rect 8186 15165 8288 15199
rect 8322 15165 8424 15199
rect 8458 15165 8560 15199
rect 8594 15165 8696 15199
rect 8730 15165 8832 15199
rect 8866 15165 8968 15199
rect 9002 15165 9104 15199
rect 9138 15165 9240 15199
rect 7880 15063 9274 15165
rect 7914 15029 8016 15063
rect 8050 15029 8152 15063
rect 8186 15029 8288 15063
rect 8322 15029 8424 15063
rect 8458 15029 8560 15063
rect 8594 15029 8696 15063
rect 8730 15029 8832 15063
rect 8866 15029 8968 15063
rect 9002 15029 9104 15063
rect 9138 15029 9240 15063
rect 7880 14927 9274 15029
rect 7914 14893 8016 14927
rect 8050 14893 8152 14927
rect 8186 14893 8288 14927
rect 8322 14893 8424 14927
rect 8458 14893 8560 14927
rect 8594 14893 8696 14927
rect 8730 14893 8832 14927
rect 8866 14893 8968 14927
rect 9002 14893 9104 14927
rect 9138 14893 9240 14927
rect 7880 14791 9274 14893
rect 7914 14757 8016 14791
rect 8050 14757 8152 14791
rect 8186 14757 8288 14791
rect 8322 14757 8424 14791
rect 8458 14757 8560 14791
rect 8594 14757 8696 14791
rect 8730 14757 8832 14791
rect 8866 14757 8968 14791
rect 9002 14757 9104 14791
rect 9138 14757 9240 14791
rect 7880 14655 9274 14757
rect 7914 14621 8016 14655
rect 8050 14621 8152 14655
rect 8186 14621 8288 14655
rect 8322 14621 8424 14655
rect 8458 14621 8560 14655
rect 8594 14621 8696 14655
rect 8730 14621 8832 14655
rect 8866 14621 8968 14655
rect 9002 14621 9104 14655
rect 9138 14621 9240 14655
rect 7880 14519 9274 14621
rect 7914 14485 8016 14519
rect 8050 14485 8152 14519
rect 8186 14485 8288 14519
rect 8322 14485 8424 14519
rect 8458 14485 8560 14519
rect 8594 14485 8696 14519
rect 8730 14485 8832 14519
rect 8866 14485 8968 14519
rect 9002 14485 9104 14519
rect 9138 14485 9240 14519
rect 7880 14383 9274 14485
rect 7914 14349 8016 14383
rect 8050 14349 8152 14383
rect 8186 14349 8288 14383
rect 8322 14349 8424 14383
rect 8458 14349 8560 14383
rect 8594 14349 8696 14383
rect 8730 14349 8832 14383
rect 8866 14349 8968 14383
rect 9002 14349 9104 14383
rect 9138 14349 9240 14383
rect 7880 14247 9274 14349
rect 7914 14213 8016 14247
rect 8050 14213 8152 14247
rect 8186 14213 8288 14247
rect 8322 14213 8424 14247
rect 8458 14213 8560 14247
rect 8594 14213 8696 14247
rect 8730 14213 8832 14247
rect 8866 14213 8968 14247
rect 9002 14213 9104 14247
rect 9138 14213 9240 14247
rect 7880 14111 9274 14213
rect 7914 14077 8016 14111
rect 8050 14077 8152 14111
rect 8186 14077 8288 14111
rect 8322 14077 8424 14111
rect 8458 14077 8560 14111
rect 8594 14077 8696 14111
rect 8730 14077 8832 14111
rect 8866 14077 8968 14111
rect 9002 14077 9104 14111
rect 9138 14077 9240 14111
rect 7880 13975 9274 14077
rect 7914 13941 8016 13975
rect 8050 13941 8152 13975
rect 8186 13941 8288 13975
rect 8322 13941 8424 13975
rect 8458 13941 8560 13975
rect 8594 13941 8696 13975
rect 8730 13941 8832 13975
rect 8866 13941 8968 13975
rect 9002 13941 9104 13975
rect 9138 13941 9240 13975
rect 7880 13839 9274 13941
rect 7914 13805 8016 13839
rect 8050 13805 8152 13839
rect 8186 13805 8288 13839
rect 8322 13805 8424 13839
rect 8458 13805 8560 13839
rect 8594 13805 8696 13839
rect 8730 13805 8832 13839
rect 8866 13805 8968 13839
rect 9002 13805 9104 13839
rect 9138 13805 9240 13839
rect 7880 13703 9274 13805
rect 7914 13669 8016 13703
rect 8050 13669 8152 13703
rect 8186 13669 8288 13703
rect 8322 13669 8424 13703
rect 8458 13669 8560 13703
rect 8594 13669 8696 13703
rect 8730 13669 8832 13703
rect 8866 13669 8968 13703
rect 9002 13669 9104 13703
rect 9138 13669 9240 13703
rect 7880 13567 9274 13669
rect 7914 13533 8016 13567
rect 8050 13533 8152 13567
rect 8186 13533 8288 13567
rect 8322 13533 8424 13567
rect 8458 13533 8560 13567
rect 8594 13533 8696 13567
rect 8730 13533 8832 13567
rect 8866 13533 8968 13567
rect 9002 13533 9104 13567
rect 9138 13533 9240 13567
rect 7880 13431 9274 13533
rect 7914 13397 8016 13431
rect 8050 13397 8152 13431
rect 8186 13397 8288 13431
rect 8322 13397 8424 13431
rect 8458 13397 8560 13431
rect 8594 13397 8696 13431
rect 8730 13397 8832 13431
rect 8866 13397 8968 13431
rect 9002 13397 9104 13431
rect 9138 13397 9240 13431
rect 7880 13295 9274 13397
rect 7914 13261 8016 13295
rect 8050 13261 8152 13295
rect 8186 13261 8288 13295
rect 8322 13261 8424 13295
rect 8458 13261 8560 13295
rect 8594 13261 8696 13295
rect 8730 13261 8832 13295
rect 8866 13261 8968 13295
rect 9002 13261 9104 13295
rect 9138 13261 9240 13295
rect 7880 13159 9274 13261
rect 7914 13125 8016 13159
rect 8050 13125 8152 13159
rect 8186 13125 8288 13159
rect 8322 13125 8424 13159
rect 8458 13125 8560 13159
rect 8594 13125 8696 13159
rect 8730 13125 8832 13159
rect 8866 13125 8968 13159
rect 9002 13125 9104 13159
rect 9138 13125 9240 13159
rect 7880 13023 9274 13125
rect 7914 12989 8016 13023
rect 8050 12989 8152 13023
rect 8186 12989 8288 13023
rect 8322 12989 8424 13023
rect 8458 12989 8560 13023
rect 8594 12989 8696 13023
rect 8730 12989 8832 13023
rect 8866 12989 8968 13023
rect 9002 12989 9104 13023
rect 9138 12989 9240 13023
rect 7880 12887 9274 12989
rect 7914 12853 8016 12887
rect 8050 12853 8152 12887
rect 8186 12853 8288 12887
rect 8322 12853 8424 12887
rect 8458 12853 8560 12887
rect 8594 12853 8696 12887
rect 8730 12853 8832 12887
rect 8866 12853 8968 12887
rect 9002 12853 9104 12887
rect 9138 12853 9240 12887
rect 7880 12751 9274 12853
rect 7914 12717 8016 12751
rect 8050 12717 8152 12751
rect 8186 12717 8288 12751
rect 8322 12717 8424 12751
rect 8458 12717 8560 12751
rect 8594 12717 8696 12751
rect 8730 12717 8832 12751
rect 8866 12717 8968 12751
rect 9002 12717 9104 12751
rect 9138 12717 9240 12751
rect 7880 12615 9274 12717
rect 7914 12581 8016 12615
rect 8050 12581 8152 12615
rect 8186 12581 8288 12615
rect 8322 12581 8424 12615
rect 8458 12581 8560 12615
rect 8594 12581 8696 12615
rect 8730 12581 8832 12615
rect 8866 12581 8968 12615
rect 9002 12581 9104 12615
rect 9138 12581 9240 12615
rect 7880 12479 9274 12581
rect 7914 12445 8016 12479
rect 8050 12445 8152 12479
rect 8186 12445 8288 12479
rect 8322 12445 8424 12479
rect 8458 12445 8560 12479
rect 8594 12445 8696 12479
rect 8730 12445 8832 12479
rect 8866 12445 8968 12479
rect 9002 12445 9104 12479
rect 9138 12445 9240 12479
rect 7880 12343 9274 12445
rect 7914 12309 8016 12343
rect 8050 12309 8152 12343
rect 8186 12309 8288 12343
rect 8322 12309 8424 12343
rect 8458 12309 8560 12343
rect 8594 12309 8696 12343
rect 8730 12309 8832 12343
rect 8866 12309 8968 12343
rect 9002 12309 9104 12343
rect 9138 12309 9240 12343
rect 7880 12207 9274 12309
rect 7914 12173 8016 12207
rect 8050 12173 8152 12207
rect 8186 12173 8288 12207
rect 8322 12173 8424 12207
rect 8458 12173 8560 12207
rect 8594 12173 8696 12207
rect 8730 12173 8832 12207
rect 8866 12173 8968 12207
rect 9002 12173 9104 12207
rect 9138 12173 9240 12207
rect 7880 12071 9274 12173
rect 7914 12037 8016 12071
rect 8050 12037 8152 12071
rect 8186 12037 8288 12071
rect 8322 12037 8424 12071
rect 8458 12037 8560 12071
rect 8594 12037 8696 12071
rect 8730 12037 8832 12071
rect 8866 12037 8968 12071
rect 9002 12037 9104 12071
rect 9138 12037 9240 12071
rect 7880 11935 9274 12037
rect 7914 11901 8016 11935
rect 8050 11901 8152 11935
rect 8186 11901 8288 11935
rect 8322 11901 8424 11935
rect 8458 11901 8560 11935
rect 8594 11901 8696 11935
rect 8730 11901 8832 11935
rect 8866 11901 8968 11935
rect 9002 11901 9104 11935
rect 9138 11901 9240 11935
rect 7880 11799 9274 11901
rect 7914 11765 8016 11799
rect 8050 11765 8152 11799
rect 8186 11765 8288 11799
rect 8322 11765 8424 11799
rect 8458 11765 8560 11799
rect 8594 11765 8696 11799
rect 8730 11765 8832 11799
rect 8866 11765 8968 11799
rect 9002 11765 9104 11799
rect 9138 11765 9240 11799
rect 7880 11663 9274 11765
rect 7914 11629 8016 11663
rect 8050 11629 8152 11663
rect 8186 11629 8288 11663
rect 8322 11629 8424 11663
rect 8458 11629 8560 11663
rect 8594 11629 8696 11663
rect 8730 11629 8832 11663
rect 8866 11629 8968 11663
rect 9002 11629 9104 11663
rect 9138 11629 9240 11663
rect 7880 11527 9274 11629
rect 7914 11493 8016 11527
rect 8050 11493 8152 11527
rect 8186 11493 8288 11527
rect 8322 11493 8424 11527
rect 8458 11493 8560 11527
rect 8594 11493 8696 11527
rect 8730 11493 8832 11527
rect 8866 11493 8968 11527
rect 9002 11493 9104 11527
rect 9138 11493 9240 11527
rect 7880 11391 9274 11493
rect 7914 11357 8016 11391
rect 8050 11357 8152 11391
rect 8186 11357 8288 11391
rect 8322 11357 8424 11391
rect 8458 11357 8560 11391
rect 8594 11357 8696 11391
rect 8730 11357 8832 11391
rect 8866 11357 8968 11391
rect 9002 11357 9104 11391
rect 9138 11357 9240 11391
rect 7880 11255 9274 11357
rect 7914 11221 8016 11255
rect 8050 11221 8152 11255
rect 8186 11221 8288 11255
rect 8322 11221 8424 11255
rect 8458 11221 8560 11255
rect 8594 11221 8696 11255
rect 8730 11221 8832 11255
rect 8866 11221 8968 11255
rect 9002 11221 9104 11255
rect 9138 11221 9240 11255
rect 7880 11119 9274 11221
rect 7914 11085 8016 11119
rect 8050 11085 8152 11119
rect 8186 11085 8288 11119
rect 8322 11085 8424 11119
rect 8458 11085 8560 11119
rect 8594 11085 8696 11119
rect 8730 11085 8832 11119
rect 8866 11085 8968 11119
rect 9002 11085 9104 11119
rect 9138 11085 9240 11119
rect 7880 10983 9274 11085
rect 7914 10949 8016 10983
rect 8050 10949 8152 10983
rect 8186 10949 8288 10983
rect 8322 10949 8424 10983
rect 8458 10949 8560 10983
rect 8594 10949 8696 10983
rect 8730 10949 8832 10983
rect 8866 10949 8968 10983
rect 9002 10949 9104 10983
rect 9138 10949 9240 10983
rect 7880 10847 9274 10949
rect 7914 10813 8016 10847
rect 8050 10813 8152 10847
rect 8186 10813 8288 10847
rect 8322 10813 8424 10847
rect 8458 10813 8560 10847
rect 8594 10813 8696 10847
rect 8730 10813 8832 10847
rect 8866 10813 8968 10847
rect 9002 10813 9104 10847
rect 9138 10813 9240 10847
rect 7880 10711 9274 10813
rect 7914 10677 8016 10711
rect 8050 10677 8152 10711
rect 8186 10677 8288 10711
rect 8322 10677 8424 10711
rect 8458 10677 8560 10711
rect 8594 10677 8696 10711
rect 8730 10677 8832 10711
rect 8866 10677 8968 10711
rect 9002 10677 9104 10711
rect 9138 10677 9240 10711
rect 7880 10575 9274 10677
rect 7914 10541 8016 10575
rect 8050 10541 8152 10575
rect 8186 10541 8288 10575
rect 8322 10541 8424 10575
rect 8458 10541 8560 10575
rect 8594 10541 8696 10575
rect 8730 10541 8832 10575
rect 8866 10541 8968 10575
rect 9002 10541 9104 10575
rect 9138 10541 9240 10575
rect 7880 10439 9274 10541
rect 7914 10405 8016 10439
rect 8050 10405 8152 10439
rect 8186 10405 8288 10439
rect 8322 10405 8424 10439
rect 8458 10405 8560 10439
rect 8594 10405 8696 10439
rect 8730 10405 8832 10439
rect 8866 10405 8968 10439
rect 9002 10405 9104 10439
rect 9138 10405 9240 10439
rect 7880 10303 9274 10405
rect 7914 10269 8016 10303
rect 8050 10269 8152 10303
rect 8186 10269 8288 10303
rect 8322 10269 8424 10303
rect 8458 10269 8560 10303
rect 8594 10269 8696 10303
rect 8730 10269 8832 10303
rect 8866 10269 8968 10303
rect 9002 10269 9104 10303
rect 9138 10269 9240 10303
rect 7880 10167 9274 10269
rect 7914 10133 8016 10167
rect 8050 10133 8152 10167
rect 8186 10133 8288 10167
rect 8322 10133 8424 10167
rect 8458 10133 8560 10167
rect 8594 10133 8696 10167
rect 8730 10133 8832 10167
rect 8866 10133 8968 10167
rect 9002 10133 9104 10167
rect 9138 10133 9240 10167
rect 7880 10031 9274 10133
rect 7914 9997 8016 10031
rect 8050 9997 8152 10031
rect 8186 9997 8288 10031
rect 8322 9997 8424 10031
rect 8458 9997 8560 10031
rect 8594 9997 8696 10031
rect 8730 9997 8832 10031
rect 8866 9997 8968 10031
rect 9002 9997 9104 10031
rect 9138 9997 9240 10031
rect 7880 9895 9274 9997
rect 7914 9861 8016 9895
rect 8050 9861 8152 9895
rect 8186 9861 8288 9895
rect 8322 9861 8424 9895
rect 8458 9861 8560 9895
rect 8594 9861 8696 9895
rect 8730 9861 8832 9895
rect 8866 9861 8968 9895
rect 9002 9861 9104 9895
rect 9138 9861 9240 9895
rect 7880 9759 9274 9861
rect 7914 9725 8016 9759
rect 8050 9725 8152 9759
rect 8186 9725 8288 9759
rect 8322 9725 8424 9759
rect 8458 9725 8560 9759
rect 8594 9725 8696 9759
rect 8730 9725 8832 9759
rect 8866 9725 8968 9759
rect 9002 9725 9104 9759
rect 9138 9725 9240 9759
rect 7880 9623 9274 9725
rect 7914 9589 8016 9623
rect 8050 9589 8152 9623
rect 8186 9589 8288 9623
rect 8322 9589 8424 9623
rect 8458 9589 8560 9623
rect 8594 9589 8696 9623
rect 8730 9589 8832 9623
rect 8866 9589 8968 9623
rect 9002 9589 9104 9623
rect 9138 9589 9240 9623
rect 7880 9487 9274 9589
rect 7914 9453 8016 9487
rect 8050 9453 8152 9487
rect 8186 9453 8288 9487
rect 8322 9453 8424 9487
rect 8458 9453 8560 9487
rect 8594 9453 8696 9487
rect 8730 9453 8832 9487
rect 8866 9453 8968 9487
rect 9002 9453 9104 9487
rect 9138 9453 9240 9487
rect 7880 9351 9274 9453
rect 7914 9317 8016 9351
rect 8050 9317 8152 9351
rect 8186 9317 8288 9351
rect 8322 9317 8424 9351
rect 8458 9317 8560 9351
rect 8594 9317 8696 9351
rect 8730 9317 8832 9351
rect 8866 9317 8968 9351
rect 9002 9317 9104 9351
rect 9138 9317 9240 9351
rect 7880 9215 9274 9317
rect 7914 9181 8016 9215
rect 8050 9181 8152 9215
rect 8186 9181 8288 9215
rect 8322 9181 8424 9215
rect 8458 9181 8560 9215
rect 8594 9181 8696 9215
rect 8730 9181 8832 9215
rect 8866 9181 8968 9215
rect 9002 9181 9104 9215
rect 9138 9181 9240 9215
rect 7880 9079 9274 9181
rect 7914 9045 8016 9079
rect 8050 9045 8152 9079
rect 8186 9045 8288 9079
rect 8322 9045 8424 9079
rect 8458 9045 8560 9079
rect 8594 9045 8696 9079
rect 8730 9045 8832 9079
rect 8866 9045 8968 9079
rect 9002 9045 9104 9079
rect 9138 9045 9240 9079
rect 7880 8943 9274 9045
rect 7914 8909 8016 8943
rect 8050 8909 8152 8943
rect 8186 8909 8288 8943
rect 8322 8909 8424 8943
rect 8458 8909 8560 8943
rect 8594 8909 8696 8943
rect 8730 8909 8832 8943
rect 8866 8909 8968 8943
rect 9002 8909 9104 8943
rect 9138 8909 9240 8943
rect 7880 8807 9274 8909
rect 7914 8773 8016 8807
rect 8050 8773 8152 8807
rect 8186 8773 8288 8807
rect 8322 8773 8424 8807
rect 8458 8773 8560 8807
rect 8594 8773 8696 8807
rect 8730 8773 8832 8807
rect 8866 8773 8968 8807
rect 9002 8773 9104 8807
rect 9138 8773 9240 8807
rect 7880 8671 9274 8773
rect 7914 8637 8016 8671
rect 8050 8637 8152 8671
rect 8186 8637 8288 8671
rect 8322 8637 8424 8671
rect 8458 8637 8560 8671
rect 8594 8637 8696 8671
rect 8730 8637 8832 8671
rect 8866 8637 8968 8671
rect 9002 8637 9104 8671
rect 9138 8637 9240 8671
rect 7880 8535 9274 8637
rect 7914 8501 8016 8535
rect 8050 8501 8152 8535
rect 8186 8501 8288 8535
rect 8322 8501 8424 8535
rect 8458 8501 8560 8535
rect 8594 8501 8696 8535
rect 8730 8501 8832 8535
rect 8866 8501 8968 8535
rect 9002 8501 9104 8535
rect 9138 8501 9240 8535
rect 7880 8399 9274 8501
rect 7914 8365 8016 8399
rect 8050 8365 8152 8399
rect 8186 8365 8288 8399
rect 8322 8365 8424 8399
rect 8458 8365 8560 8399
rect 8594 8365 8696 8399
rect 8730 8365 8832 8399
rect 8866 8365 8968 8399
rect 9002 8365 9104 8399
rect 9138 8365 9240 8399
rect 7880 8263 9274 8365
rect 7914 8229 8016 8263
rect 8050 8229 8152 8263
rect 8186 8229 8288 8263
rect 8322 8229 8424 8263
rect 8458 8229 8560 8263
rect 8594 8229 8696 8263
rect 8730 8229 8832 8263
rect 8866 8229 8968 8263
rect 9002 8229 9104 8263
rect 9138 8229 9240 8263
rect 7880 8127 9274 8229
rect 7914 8093 8016 8127
rect 8050 8093 8152 8127
rect 8186 8093 8288 8127
rect 8322 8093 8424 8127
rect 8458 8093 8560 8127
rect 8594 8093 8696 8127
rect 8730 8093 8832 8127
rect 8866 8093 8968 8127
rect 9002 8093 9104 8127
rect 9138 8093 9240 8127
rect 7880 7991 9274 8093
rect 7914 7957 8016 7991
rect 8050 7957 8152 7991
rect 8186 7957 8288 7991
rect 8322 7957 8424 7991
rect 8458 7957 8560 7991
rect 8594 7957 8696 7991
rect 8730 7957 8832 7991
rect 8866 7957 8968 7991
rect 9002 7957 9104 7991
rect 9138 7957 9240 7991
rect 7880 7855 9274 7957
rect 7914 7821 8016 7855
rect 8050 7821 8152 7855
rect 8186 7821 8288 7855
rect 8322 7821 8424 7855
rect 8458 7821 8560 7855
rect 8594 7821 8696 7855
rect 8730 7821 8832 7855
rect 8866 7821 8968 7855
rect 9002 7821 9104 7855
rect 9138 7821 9240 7855
rect 7880 7719 9274 7821
rect 7914 7685 8016 7719
rect 8050 7685 8152 7719
rect 8186 7685 8288 7719
rect 8322 7685 8424 7719
rect 8458 7685 8560 7719
rect 8594 7685 8696 7719
rect 8730 7685 8832 7719
rect 8866 7685 8968 7719
rect 9002 7685 9104 7719
rect 9138 7685 9240 7719
rect 7880 7583 9274 7685
rect 7914 7549 8016 7583
rect 8050 7549 8152 7583
rect 8186 7549 8288 7583
rect 8322 7549 8424 7583
rect 8458 7549 8560 7583
rect 8594 7549 8696 7583
rect 8730 7549 8832 7583
rect 8866 7549 8968 7583
rect 9002 7549 9104 7583
rect 9138 7549 9240 7583
rect 7880 7447 9274 7549
rect 7914 7413 8016 7447
rect 8050 7413 8152 7447
rect 8186 7413 8288 7447
rect 8322 7413 8424 7447
rect 8458 7413 8560 7447
rect 8594 7413 8696 7447
rect 8730 7413 8832 7447
rect 8866 7413 8968 7447
rect 9002 7413 9104 7447
rect 9138 7413 9240 7447
rect 7880 7311 9274 7413
rect 7914 7277 8016 7311
rect 8050 7277 8152 7311
rect 8186 7277 8288 7311
rect 8322 7277 8424 7311
rect 8458 7277 8560 7311
rect 8594 7277 8696 7311
rect 8730 7277 8832 7311
rect 8866 7277 8968 7311
rect 9002 7277 9104 7311
rect 9138 7277 9240 7311
rect 7880 7175 9274 7277
rect 7914 7141 8016 7175
rect 8050 7141 8152 7175
rect 8186 7141 8288 7175
rect 8322 7141 8424 7175
rect 8458 7141 8560 7175
rect 8594 7141 8696 7175
rect 8730 7141 8832 7175
rect 8866 7141 8968 7175
rect 9002 7141 9104 7175
rect 9138 7141 9240 7175
rect 7880 7039 9274 7141
rect 7914 7005 8016 7039
rect 8050 7005 8152 7039
rect 8186 7005 8288 7039
rect 8322 7005 8424 7039
rect 8458 7005 8560 7039
rect 8594 7005 8696 7039
rect 8730 7005 8832 7039
rect 8866 7005 8968 7039
rect 9002 7005 9104 7039
rect 9138 7005 9240 7039
rect 7880 6903 9274 7005
rect 7914 6869 8016 6903
rect 8050 6869 8152 6903
rect 8186 6869 8288 6903
rect 8322 6869 8424 6903
rect 8458 6869 8560 6903
rect 8594 6869 8696 6903
rect 8730 6869 8832 6903
rect 8866 6869 8968 6903
rect 9002 6869 9104 6903
rect 9138 6869 9240 6903
rect 7880 6767 9274 6869
rect 7914 6733 8016 6767
rect 8050 6733 8152 6767
rect 8186 6733 8288 6767
rect 8322 6733 8424 6767
rect 8458 6733 8560 6767
rect 8594 6733 8696 6767
rect 8730 6733 8832 6767
rect 8866 6733 8968 6767
rect 9002 6733 9104 6767
rect 9138 6733 9240 6767
rect 7880 6631 9274 6733
rect 7914 6597 8016 6631
rect 8050 6597 8152 6631
rect 8186 6597 8288 6631
rect 8322 6597 8424 6631
rect 8458 6597 8560 6631
rect 8594 6597 8696 6631
rect 8730 6597 8832 6631
rect 8866 6597 8968 6631
rect 9002 6597 9104 6631
rect 9138 6597 9240 6631
rect 7880 6495 9274 6597
rect 7914 6461 8016 6495
rect 8050 6461 8152 6495
rect 8186 6461 8288 6495
rect 8322 6461 8424 6495
rect 8458 6461 8560 6495
rect 8594 6461 8696 6495
rect 8730 6461 8832 6495
rect 8866 6461 8968 6495
rect 9002 6461 9104 6495
rect 9138 6461 9240 6495
rect 7880 6359 9274 6461
rect 7914 6325 8016 6359
rect 8050 6325 8152 6359
rect 8186 6325 8288 6359
rect 8322 6325 8424 6359
rect 8458 6325 8560 6359
rect 8594 6325 8696 6359
rect 8730 6325 8832 6359
rect 8866 6325 8968 6359
rect 9002 6325 9104 6359
rect 9138 6325 9240 6359
rect 7880 6223 9274 6325
rect 7914 6189 8016 6223
rect 8050 6189 8152 6223
rect 8186 6189 8288 6223
rect 8322 6189 8424 6223
rect 8458 6189 8560 6223
rect 8594 6189 8696 6223
rect 8730 6189 8832 6223
rect 8866 6189 8968 6223
rect 9002 6189 9104 6223
rect 9138 6189 9240 6223
rect 7880 6087 9274 6189
rect 7914 6053 8016 6087
rect 8050 6053 8152 6087
rect 8186 6053 8288 6087
rect 8322 6053 8424 6087
rect 8458 6053 8560 6087
rect 8594 6053 8696 6087
rect 8730 6053 8832 6087
rect 8866 6053 8968 6087
rect 9002 6053 9104 6087
rect 9138 6053 9240 6087
rect 7880 5951 9274 6053
rect 7914 5917 8016 5951
rect 8050 5917 8152 5951
rect 8186 5917 8288 5951
rect 8322 5917 8424 5951
rect 8458 5917 8560 5951
rect 8594 5917 8696 5951
rect 8730 5917 8832 5951
rect 8866 5917 8968 5951
rect 9002 5917 9104 5951
rect 9138 5917 9240 5951
rect 7880 5815 9274 5917
rect 7914 5781 8016 5815
rect 8050 5781 8152 5815
rect 8186 5781 8288 5815
rect 8322 5781 8424 5815
rect 8458 5781 8560 5815
rect 8594 5781 8696 5815
rect 8730 5781 8832 5815
rect 8866 5781 8968 5815
rect 9002 5781 9104 5815
rect 9138 5781 9240 5815
rect 7880 5679 9274 5781
rect 7914 5645 8016 5679
rect 8050 5645 8152 5679
rect 8186 5645 8288 5679
rect 8322 5645 8424 5679
rect 8458 5645 8560 5679
rect 8594 5645 8696 5679
rect 8730 5645 8832 5679
rect 8866 5645 8968 5679
rect 9002 5645 9104 5679
rect 9138 5645 9240 5679
rect 7880 5543 9274 5645
rect 7914 5509 8016 5543
rect 8050 5509 8152 5543
rect 8186 5509 8288 5543
rect 8322 5509 8424 5543
rect 8458 5509 8560 5543
rect 8594 5509 8696 5543
rect 8730 5509 8832 5543
rect 8866 5509 8968 5543
rect 9002 5509 9104 5543
rect 9138 5509 9240 5543
rect 7880 5407 9274 5509
rect 7914 5373 8016 5407
rect 8050 5373 8152 5407
rect 8186 5373 8288 5407
rect 8322 5373 8424 5407
rect 8458 5373 8560 5407
rect 8594 5373 8696 5407
rect 8730 5373 8832 5407
rect 8866 5373 8968 5407
rect 9002 5373 9104 5407
rect 9138 5373 9240 5407
rect 7880 5271 9274 5373
rect 7914 5237 8016 5271
rect 8050 5237 8152 5271
rect 8186 5237 8288 5271
rect 8322 5237 8424 5271
rect 8458 5237 8560 5271
rect 8594 5237 8696 5271
rect 8730 5237 8832 5271
rect 8866 5237 8968 5271
rect 9002 5237 9104 5271
rect 9138 5237 9240 5271
rect 7880 5135 9274 5237
rect 7914 5101 8016 5135
rect 8050 5101 8152 5135
rect 8186 5101 8288 5135
rect 8322 5101 8424 5135
rect 8458 5101 8560 5135
rect 8594 5101 8696 5135
rect 8730 5101 8832 5135
rect 8866 5101 8968 5135
rect 9002 5101 9104 5135
rect 9138 5101 9240 5135
rect 7880 4999 9274 5101
rect 7914 4965 8016 4999
rect 8050 4965 8152 4999
rect 8186 4965 8288 4999
rect 8322 4965 8424 4999
rect 8458 4965 8560 4999
rect 8594 4965 8696 4999
rect 8730 4965 8832 4999
rect 8866 4965 8968 4999
rect 9002 4965 9104 4999
rect 9138 4965 9240 4999
rect 7880 4863 9274 4965
rect 7914 4829 8016 4863
rect 8050 4829 8152 4863
rect 8186 4829 8288 4863
rect 8322 4829 8424 4863
rect 8458 4829 8560 4863
rect 8594 4829 8696 4863
rect 8730 4829 8832 4863
rect 8866 4829 8968 4863
rect 9002 4829 9104 4863
rect 9138 4829 9240 4863
rect 7880 4727 9274 4829
rect 7914 4693 8016 4727
rect 8050 4693 8152 4727
rect 8186 4693 8288 4727
rect 8322 4693 8424 4727
rect 8458 4693 8560 4727
rect 8594 4693 8696 4727
rect 8730 4693 8832 4727
rect 8866 4693 8968 4727
rect 9002 4693 9104 4727
rect 9138 4693 9240 4727
rect 7880 4591 9274 4693
rect 7914 4557 8016 4591
rect 8050 4557 8152 4591
rect 8186 4557 8288 4591
rect 8322 4557 8424 4591
rect 8458 4557 8560 4591
rect 8594 4557 8696 4591
rect 8730 4557 8832 4591
rect 8866 4557 8968 4591
rect 9002 4557 9104 4591
rect 9138 4557 9240 4591
rect 7880 4455 9274 4557
rect 7914 4421 8016 4455
rect 8050 4421 8152 4455
rect 8186 4421 8288 4455
rect 8322 4421 8424 4455
rect 8458 4421 8560 4455
rect 8594 4421 8696 4455
rect 8730 4421 8832 4455
rect 8866 4421 8968 4455
rect 9002 4421 9104 4455
rect 9138 4421 9240 4455
rect 7880 4319 9274 4421
rect 7914 4285 8016 4319
rect 8050 4285 8152 4319
rect 8186 4285 8288 4319
rect 8322 4285 8424 4319
rect 8458 4285 8560 4319
rect 8594 4285 8696 4319
rect 8730 4285 8832 4319
rect 8866 4285 8968 4319
rect 9002 4285 9104 4319
rect 9138 4285 9240 4319
rect 7880 4183 9274 4285
rect 7914 4149 8016 4183
rect 8050 4149 8152 4183
rect 8186 4149 8288 4183
rect 8322 4149 8424 4183
rect 8458 4149 8560 4183
rect 8594 4149 8696 4183
rect 8730 4149 8832 4183
rect 8866 4149 8968 4183
rect 9002 4149 9104 4183
rect 9138 4149 9240 4183
rect 7880 4047 9274 4149
rect 7914 4013 8016 4047
rect 8050 4013 8152 4047
rect 8186 4013 8288 4047
rect 8322 4013 8424 4047
rect 8458 4013 8560 4047
rect 8594 4013 8696 4047
rect 8730 4013 8832 4047
rect 8866 4013 8968 4047
rect 9002 4013 9104 4047
rect 9138 4013 9240 4047
rect 7880 3911 9274 4013
rect 7914 3877 8016 3911
rect 8050 3877 8152 3911
rect 8186 3877 8288 3911
rect 8322 3877 8424 3911
rect 8458 3877 8560 3911
rect 8594 3877 8696 3911
rect 8730 3877 8832 3911
rect 8866 3877 8968 3911
rect 9002 3877 9104 3911
rect 9138 3877 9240 3911
rect 7880 3775 9274 3877
rect 7914 3741 8016 3775
rect 8050 3741 8152 3775
rect 8186 3741 8288 3775
rect 8322 3741 8424 3775
rect 8458 3741 8560 3775
rect 8594 3741 8696 3775
rect 8730 3741 8832 3775
rect 8866 3741 8968 3775
rect 9002 3741 9104 3775
rect 9138 3741 9240 3775
rect 7880 3639 9274 3741
rect 7914 3605 8016 3639
rect 8050 3605 8152 3639
rect 8186 3605 8288 3639
rect 8322 3605 8424 3639
rect 8458 3605 8560 3639
rect 8594 3605 8696 3639
rect 8730 3605 8832 3639
rect 8866 3605 8968 3639
rect 9002 3605 9104 3639
rect 9138 3605 9240 3639
rect 7880 3503 9274 3605
rect 7914 3469 8016 3503
rect 8050 3469 8152 3503
rect 8186 3469 8288 3503
rect 8322 3469 8424 3503
rect 8458 3469 8560 3503
rect 8594 3469 8696 3503
rect 8730 3469 8832 3503
rect 8866 3469 8968 3503
rect 9002 3469 9104 3503
rect 9138 3469 9240 3503
rect 7880 3367 9274 3469
rect 7914 3333 8016 3367
rect 8050 3333 8152 3367
rect 8186 3333 8288 3367
rect 8322 3333 8424 3367
rect 8458 3333 8560 3367
rect 8594 3333 8696 3367
rect 8730 3333 8832 3367
rect 8866 3333 8968 3367
rect 9002 3333 9104 3367
rect 9138 3333 9240 3367
rect 7880 3231 9274 3333
rect 7914 3197 8016 3231
rect 8050 3197 8152 3231
rect 8186 3197 8288 3231
rect 8322 3197 8424 3231
rect 8458 3197 8560 3231
rect 8594 3197 8696 3231
rect 8730 3197 8832 3231
rect 8866 3197 8968 3231
rect 9002 3197 9104 3231
rect 9138 3197 9240 3231
rect 7880 3095 9274 3197
rect 7914 3061 8016 3095
rect 8050 3061 8152 3095
rect 8186 3061 8288 3095
rect 8322 3061 8424 3095
rect 8458 3061 8560 3095
rect 8594 3061 8696 3095
rect 8730 3061 8832 3095
rect 8866 3061 8968 3095
rect 9002 3061 9104 3095
rect 9138 3061 9240 3095
rect 7880 2959 9274 3061
rect 7914 2925 8016 2959
rect 8050 2925 8152 2959
rect 8186 2925 8288 2959
rect 8322 2925 8424 2959
rect 8458 2925 8560 2959
rect 8594 2925 8696 2959
rect 8730 2925 8832 2959
rect 8866 2925 8968 2959
rect 9002 2925 9104 2959
rect 9138 2925 9240 2959
rect 7880 2823 9274 2925
rect 7914 2789 8016 2823
rect 8050 2789 8152 2823
rect 8186 2789 8288 2823
rect 8322 2789 8424 2823
rect 8458 2789 8560 2823
rect 8594 2789 8696 2823
rect 8730 2789 8832 2823
rect 8866 2789 8968 2823
rect 9002 2789 9104 2823
rect 9138 2789 9240 2823
rect 7880 2687 9274 2789
rect 7914 2653 8016 2687
rect 8050 2653 8152 2687
rect 8186 2653 8288 2687
rect 8322 2653 8424 2687
rect 8458 2653 8560 2687
rect 8594 2653 8696 2687
rect 8730 2653 8832 2687
rect 8866 2653 8968 2687
rect 9002 2653 9104 2687
rect 9138 2653 9240 2687
rect 7880 2551 9274 2653
rect 7914 2517 8016 2551
rect 8050 2517 8152 2551
rect 8186 2517 8288 2551
rect 8322 2517 8424 2551
rect 8458 2517 8560 2551
rect 8594 2517 8696 2551
rect 8730 2517 8832 2551
rect 8866 2517 8968 2551
rect 9002 2517 9104 2551
rect 9138 2517 9240 2551
rect 7880 2414 9274 2517
rect 7914 2380 8016 2414
rect 8050 2380 8152 2414
rect 8186 2380 8288 2414
rect 8322 2380 8424 2414
rect 8458 2380 8560 2414
rect 8594 2380 8696 2414
rect 8730 2380 8832 2414
rect 8866 2380 8968 2414
rect 9002 2380 9104 2414
rect 9138 2380 9240 2414
rect 7880 2277 9274 2380
rect 7914 2243 8016 2277
rect 8050 2243 8152 2277
rect 8186 2243 8288 2277
rect 8322 2243 8424 2277
rect 8458 2243 8560 2277
rect 8594 2243 8696 2277
rect 8730 2243 8832 2277
rect 8866 2243 8968 2277
rect 9002 2243 9104 2277
rect 9138 2243 9240 2277
rect 7880 2140 9274 2243
rect 7914 2106 8016 2140
rect 8050 2106 8152 2140
rect 8186 2106 8288 2140
rect 8322 2106 8424 2140
rect 8458 2106 8560 2140
rect 8594 2106 8696 2140
rect 8730 2106 8832 2140
rect 8866 2106 8968 2140
rect 9002 2106 9104 2140
rect 9138 2106 9240 2140
rect 7880 2003 9274 2106
rect 7914 1969 8016 2003
rect 8050 1969 8152 2003
rect 8186 1969 8288 2003
rect 8322 1969 8424 2003
rect 8458 1969 8560 2003
rect 8594 1969 8696 2003
rect 8730 1969 8832 2003
rect 8866 1969 8968 2003
rect 9002 1969 9104 2003
rect 9138 1969 9240 2003
rect 7880 1866 9274 1969
rect 7914 1832 8016 1866
rect 8050 1832 8152 1866
rect 8186 1832 8288 1866
rect 8322 1832 8424 1866
rect 8458 1832 8560 1866
rect 8594 1832 8696 1866
rect 8730 1832 8832 1866
rect 8866 1832 8968 1866
rect 9002 1832 9104 1866
rect 9138 1832 9240 1866
rect 7880 1729 9274 1832
rect 359 1695 461 1729
rect 495 1695 597 1729
rect 631 1695 733 1729
rect 767 1695 869 1729
rect 903 1695 1005 1729
rect 1039 1695 1141 1729
rect 1175 1695 1277 1729
rect 1311 1695 1413 1729
rect 1447 1695 1549 1729
rect 1583 1695 1685 1729
rect 325 1592 1719 1695
rect 359 1558 461 1592
rect 495 1558 597 1592
rect 631 1558 733 1592
rect 767 1558 869 1592
rect 903 1558 1005 1592
rect 1039 1558 1141 1592
rect 1175 1558 1277 1592
rect 1311 1558 1413 1592
rect 1447 1558 1549 1592
rect 1583 1558 1685 1592
rect 325 1455 1719 1558
rect 359 1421 461 1455
rect 495 1421 597 1455
rect 631 1421 733 1455
rect 767 1421 869 1455
rect 903 1421 1005 1455
rect 1039 1421 1141 1455
rect 1175 1421 1277 1455
rect 1311 1421 1413 1455
rect 1447 1421 1549 1455
rect 1583 1421 1685 1455
rect 325 1318 1719 1421
rect 359 1284 461 1318
rect 495 1284 597 1318
rect 631 1284 733 1318
rect 767 1284 869 1318
rect 903 1284 1005 1318
rect 1039 1284 1141 1318
rect 1175 1284 1277 1318
rect 1311 1284 1413 1318
rect 1447 1284 1549 1318
rect 1583 1284 1685 1318
rect 325 1181 1719 1284
rect 359 1147 461 1181
rect 495 1147 597 1181
rect 631 1147 733 1181
rect 767 1147 869 1181
rect 903 1147 1005 1181
rect 1039 1147 1141 1181
rect 1175 1147 1277 1181
rect 1311 1147 1413 1181
rect 1447 1147 1549 1181
rect 1583 1147 1685 1181
rect 325 1044 1719 1147
rect 359 1010 461 1044
rect 495 1010 597 1044
rect 631 1010 733 1044
rect 767 1010 869 1044
rect 903 1010 1005 1044
rect 1039 1010 1141 1044
rect 1175 1010 1277 1044
rect 1311 1010 1413 1044
rect 1447 1010 1549 1044
rect 1583 1010 1685 1044
rect 325 907 1719 1010
rect 359 873 461 907
rect 495 873 597 907
rect 631 873 733 907
rect 767 873 869 907
rect 903 873 1005 907
rect 1039 873 1141 907
rect 1175 873 1277 907
rect 1311 873 1413 907
rect 1447 873 1549 907
rect 1583 873 1685 907
rect 325 770 1719 873
rect 359 736 461 770
rect 495 736 597 770
rect 631 736 733 770
rect 767 736 869 770
rect 903 736 1005 770
rect 1039 736 1141 770
rect 1175 736 1277 770
rect 1311 736 1413 770
rect 1447 736 1549 770
rect 1583 736 1685 770
rect 325 633 1719 736
rect 359 599 461 633
rect 495 599 597 633
rect 631 599 733 633
rect 767 599 869 633
rect 903 599 1005 633
rect 1039 599 1141 633
rect 1175 599 1277 633
rect 1311 599 1413 633
rect 1447 599 1549 633
rect 1583 599 1685 633
rect 325 496 1719 599
rect 359 462 461 496
rect 495 462 597 496
rect 631 462 733 496
rect 767 462 869 496
rect 903 462 1005 496
rect 1039 462 1141 496
rect 1175 462 1277 496
rect 1311 462 1413 496
rect 1447 462 1549 496
rect 1583 462 1685 496
rect 325 359 1719 462
rect 359 325 461 359
rect 495 325 597 359
rect 631 325 733 359
rect 767 325 869 359
rect 903 325 1005 359
rect 1039 325 1141 359
rect 1175 325 1277 359
rect 1311 325 1413 359
rect 1447 325 1549 359
rect 1583 325 1685 359
rect 325 222 1719 325
rect 359 188 461 222
rect 495 188 597 222
rect 631 188 733 222
rect 767 188 869 222
rect 903 188 1005 222
rect 1039 188 1141 222
rect 1175 188 1277 222
rect 1311 188 1413 222
rect 1447 188 1549 222
rect 1583 188 1685 222
rect 325 85 1719 188
rect 359 51 461 85
rect 495 51 597 85
rect 631 51 733 85
rect 767 51 869 85
rect 903 51 1005 85
rect 1039 51 1141 85
rect 1175 51 1277 85
rect 1311 51 1413 85
rect 1447 51 1549 85
rect 1583 51 1685 85
rect 325 27 1719 51
rect 7914 1695 8016 1729
rect 8050 1695 8152 1729
rect 8186 1695 8288 1729
rect 8322 1695 8424 1729
rect 8458 1695 8560 1729
rect 8594 1695 8696 1729
rect 8730 1695 8832 1729
rect 8866 1695 8968 1729
rect 9002 1695 9104 1729
rect 9138 1695 9240 1729
rect 7880 1592 9274 1695
rect 7914 1558 8016 1592
rect 8050 1558 8152 1592
rect 8186 1558 8288 1592
rect 8322 1558 8424 1592
rect 8458 1558 8560 1592
rect 8594 1558 8696 1592
rect 8730 1558 8832 1592
rect 8866 1558 8968 1592
rect 9002 1558 9104 1592
rect 9138 1558 9240 1592
rect 7880 1455 9274 1558
rect 7914 1421 8016 1455
rect 8050 1421 8152 1455
rect 8186 1421 8288 1455
rect 8322 1421 8424 1455
rect 8458 1421 8560 1455
rect 8594 1421 8696 1455
rect 8730 1421 8832 1455
rect 8866 1421 8968 1455
rect 9002 1421 9104 1455
rect 9138 1421 9240 1455
rect 7880 1318 9274 1421
rect 7914 1284 8016 1318
rect 8050 1284 8152 1318
rect 8186 1284 8288 1318
rect 8322 1284 8424 1318
rect 8458 1284 8560 1318
rect 8594 1284 8696 1318
rect 8730 1284 8832 1318
rect 8866 1284 8968 1318
rect 9002 1284 9104 1318
rect 9138 1284 9240 1318
rect 7880 1181 9274 1284
rect 7914 1147 8016 1181
rect 8050 1147 8152 1181
rect 8186 1147 8288 1181
rect 8322 1147 8424 1181
rect 8458 1147 8560 1181
rect 8594 1147 8696 1181
rect 8730 1147 8832 1181
rect 8866 1147 8968 1181
rect 9002 1147 9104 1181
rect 9138 1147 9240 1181
rect 7880 1044 9274 1147
rect 7914 1010 8016 1044
rect 8050 1010 8152 1044
rect 8186 1010 8288 1044
rect 8322 1010 8424 1044
rect 8458 1010 8560 1044
rect 8594 1010 8696 1044
rect 8730 1010 8832 1044
rect 8866 1010 8968 1044
rect 9002 1010 9104 1044
rect 9138 1010 9240 1044
rect 7880 907 9274 1010
rect 7914 873 8016 907
rect 8050 873 8152 907
rect 8186 873 8288 907
rect 8322 873 8424 907
rect 8458 873 8560 907
rect 8594 873 8696 907
rect 8730 873 8832 907
rect 8866 873 8968 907
rect 9002 873 9104 907
rect 9138 873 9240 907
rect 7880 770 9274 873
rect 7914 736 8016 770
rect 8050 736 8152 770
rect 8186 736 8288 770
rect 8322 736 8424 770
rect 8458 736 8560 770
rect 8594 736 8696 770
rect 8730 736 8832 770
rect 8866 736 8968 770
rect 9002 736 9104 770
rect 9138 736 9240 770
rect 7880 633 9274 736
rect 7914 599 8016 633
rect 8050 599 8152 633
rect 8186 599 8288 633
rect 8322 599 8424 633
rect 8458 599 8560 633
rect 8594 599 8696 633
rect 8730 599 8832 633
rect 8866 599 8968 633
rect 9002 599 9104 633
rect 9138 599 9240 633
rect 7880 496 9274 599
rect 7914 462 8016 496
rect 8050 462 8152 496
rect 8186 462 8288 496
rect 8322 462 8424 496
rect 8458 462 8560 496
rect 8594 462 8696 496
rect 8730 462 8832 496
rect 8866 462 8968 496
rect 9002 462 9104 496
rect 9138 462 9240 496
rect 7880 359 9274 462
rect 7914 325 8016 359
rect 8050 325 8152 359
rect 8186 325 8288 359
rect 8322 325 8424 359
rect 8458 325 8560 359
rect 8594 325 8696 359
rect 8730 325 8832 359
rect 8866 325 8968 359
rect 9002 325 9104 359
rect 9138 325 9240 359
rect 7880 222 9274 325
rect 7914 188 8016 222
rect 8050 188 8152 222
rect 8186 188 8288 222
rect 8322 188 8424 222
rect 8458 188 8560 222
rect 8594 188 8696 222
rect 8730 188 8832 222
rect 8866 188 8968 222
rect 9002 188 9104 222
rect 9138 188 9240 222
rect 7880 85 9274 188
rect 7914 51 8016 85
rect 8050 51 8152 85
rect 8186 51 8288 85
rect 8322 51 8424 85
rect 8458 51 8560 85
rect 8594 51 8696 85
rect 8730 51 8832 85
rect 8866 51 8968 85
rect 9002 51 9104 85
rect 9138 51 9240 85
rect 7880 27 9274 51
<< mvnsubdiff >>
rect 5004 16438 5139 16472
rect 5173 16438 5207 16472
rect 5241 16438 5275 16472
rect 5309 16438 5343 16472
rect 5377 16438 5411 16472
rect 5445 16438 5479 16472
rect 5513 16438 5547 16472
rect 5581 16438 5615 16472
rect 5649 16438 5683 16472
rect 5717 16438 5751 16472
rect 5785 16438 5819 16472
rect 5853 16438 5887 16472
rect 5921 16438 5955 16472
rect 5989 16438 6023 16472
rect 6057 16438 6091 16472
rect 6125 16438 6159 16472
rect 6193 16438 6227 16472
rect 6261 16438 6295 16472
rect 6329 16438 6363 16472
rect 6397 16438 6431 16472
rect 6465 16438 6499 16472
rect 6533 16438 6567 16472
rect 6601 16438 6635 16472
rect 6669 16438 6703 16472
rect 6737 16438 6771 16472
rect 6805 16438 6839 16472
rect 6873 16438 6907 16472
rect 6941 16438 6975 16472
rect 7009 16438 7043 16472
rect 7077 16438 7111 16472
rect 7145 16438 7179 16472
rect 7213 16438 7247 16472
rect 7281 16438 7315 16472
rect 7349 16438 7383 16472
rect 7417 16438 7451 16472
rect 7485 16438 7553 16472
rect 5004 16404 5038 16438
rect 5004 16336 5038 16370
rect 5004 16268 5038 16302
rect 5004 16200 5038 16234
rect 5004 16132 5038 16166
rect 5004 16064 5038 16098
rect 5004 15996 5038 16030
rect 5004 15928 5038 15962
rect 5004 15860 5038 15894
rect 5004 15792 5038 15826
rect 5004 15724 5038 15758
rect 5004 15656 5038 15690
rect 5004 15588 5038 15622
rect 5004 15520 5038 15554
rect 5004 15452 5038 15486
rect 5004 15384 5038 15418
rect 5004 15316 5038 15350
rect 5004 15248 5038 15282
rect 5004 15180 5038 15214
rect 5004 15112 5038 15146
rect 5004 15044 5038 15078
rect 5004 14976 5038 15010
rect 5004 14908 5038 14942
rect 5004 14840 5038 14874
rect 5004 14772 5038 14806
rect 5004 14704 5038 14738
rect 5004 14636 5038 14670
rect 5004 14568 5038 14602
rect 5004 14500 5038 14534
rect 5004 14432 5038 14466
rect 5004 14364 5038 14398
rect 5004 14296 5038 14330
rect 5004 14228 5038 14262
rect 5004 14160 5038 14194
rect 5004 14092 5038 14126
rect 5004 14024 5038 14058
rect 5004 13956 5038 13990
rect 5004 13888 5038 13922
rect 5004 13820 5038 13854
rect 5004 13752 5038 13786
rect 5004 13684 5038 13718
rect 5004 13616 5038 13650
rect 5004 13548 5038 13582
rect 5004 13480 5038 13514
rect 5004 13412 5038 13446
rect 5004 13344 5038 13378
rect 5004 13276 5038 13310
rect 5004 13208 5038 13242
rect 5004 13140 5038 13174
rect 5004 13072 5038 13106
rect 5004 13004 5038 13038
rect 5004 12936 5038 12970
rect 5004 12868 5038 12902
rect 5004 12800 5038 12834
rect 5004 12732 5038 12766
rect 5004 12664 5038 12698
rect 5004 12596 5038 12630
rect 5004 12528 5038 12562
rect 5004 12460 5038 12494
rect 5004 12392 5038 12426
rect 5004 12324 5038 12358
rect 5004 12256 5038 12290
rect 5004 12188 5038 12222
rect 5004 12120 5038 12154
rect 5004 12052 5038 12086
rect 5004 11984 5038 12018
rect 5004 11916 5038 11950
rect 5004 11848 5038 11882
rect 5004 11780 5038 11814
rect 5004 11712 5038 11746
rect 5004 11644 5038 11678
rect 5004 11576 5038 11610
rect 5004 11508 5038 11542
rect 5004 11440 5038 11474
rect 5004 11372 5038 11406
rect 5004 11304 5038 11338
rect 5004 11236 5038 11270
rect 5004 11168 5038 11202
rect 5004 11100 5038 11134
rect 5004 11032 5038 11066
rect 5004 10964 5038 10998
rect 5004 10896 5038 10930
rect 5004 10828 5038 10862
rect 5004 10760 5038 10794
rect 5004 10692 5038 10726
rect 5004 10624 5038 10658
rect 5004 10556 5038 10590
rect 5004 10488 5038 10522
rect 5004 10420 5038 10454
rect 5004 10352 5038 10386
rect 5004 10284 5038 10318
rect 5004 10216 5038 10250
rect 5004 10148 5038 10182
rect 5004 10080 5038 10114
rect 5004 10012 5038 10046
rect 5004 9944 5038 9978
rect 5004 9876 5038 9910
rect 5004 9808 5038 9842
rect 5004 9740 5038 9774
rect 5004 9672 5038 9706
rect 5004 9604 5038 9638
rect 5004 9536 5038 9570
rect 5004 9468 5038 9502
rect 5004 9400 5038 9434
rect 5004 9332 5038 9366
rect 5004 9264 5038 9298
rect 5004 9196 5038 9230
rect 5004 9128 5038 9162
rect 5004 9060 5038 9094
rect 5004 8992 5038 9026
rect 5004 8924 5038 8958
rect 5004 8856 5038 8890
rect 5004 8788 5038 8822
rect 5004 8720 5038 8754
rect 5004 8652 5038 8686
rect 5004 8584 5038 8618
rect 5004 8516 5038 8550
rect 5004 8448 5038 8482
rect 5004 8380 5038 8414
rect 5004 8312 5038 8346
rect 5004 8244 5038 8278
rect 5004 8176 5038 8210
rect 5004 8108 5038 8142
rect 5004 8040 5038 8074
rect 5004 7972 5038 8006
rect 5004 7904 5038 7938
rect 5004 7836 5038 7870
rect 5004 7768 5038 7802
rect 5004 7700 5038 7734
rect 5004 7632 5038 7666
rect 5004 7564 5038 7598
rect 5004 7496 5038 7530
rect 5004 7428 5038 7462
rect 5004 7360 5038 7394
rect 5004 7292 5038 7326
rect 5004 7224 5038 7258
rect 5004 7156 5038 7190
rect 5004 7088 5038 7122
rect 5004 7020 5038 7054
rect 5004 6952 5038 6986
rect 5004 6884 5038 6918
rect 5004 6816 5038 6850
rect 5004 6748 5038 6782
rect 5004 6680 5038 6714
rect 5004 6612 5038 6646
rect 5004 6544 5038 6578
rect 5004 6476 5038 6510
rect 5004 6408 5038 6442
rect 5004 6340 5038 6374
rect 5004 6272 5038 6306
rect 5004 6204 5038 6238
rect 5004 6136 5038 6170
rect 5004 6068 5038 6102
rect 5004 6000 5038 6034
rect 5004 5932 5038 5966
rect 5004 5864 5038 5898
rect 5004 5796 5038 5830
rect 5004 5728 5038 5762
rect 5004 5660 5038 5694
rect 5004 5592 5038 5626
rect 5004 5524 5038 5558
rect 5004 5456 5038 5490
rect 5004 5388 5038 5422
rect 5004 5320 5038 5354
rect 5004 5252 5038 5286
rect 5004 5184 5038 5218
rect 5004 5116 5038 5150
rect 5004 5048 5038 5082
rect 5004 4980 5038 5014
rect 5004 4912 5038 4946
rect 5004 4844 5038 4878
rect 5004 4776 5038 4810
rect 5004 4708 5038 4742
rect 5004 4640 5038 4674
rect 5004 4572 5038 4606
rect 5004 4504 5038 4538
rect 5004 4436 5038 4470
rect 5004 4368 5038 4402
rect 5004 4300 5038 4334
rect 5004 4232 5038 4266
rect 5004 4164 5038 4198
rect 5004 4096 5038 4130
rect 5004 4028 5038 4062
rect 5004 3960 5038 3994
rect 5004 3892 5038 3926
rect 5004 3824 5038 3858
rect 5004 3756 5038 3790
rect 5004 3688 5038 3722
rect 5004 3620 5038 3654
rect 5004 3552 5038 3586
rect 5004 3484 5038 3518
rect 5004 3416 5038 3450
rect 5004 3348 5038 3382
rect 5004 3280 5038 3314
rect 5004 3212 5038 3246
rect 5004 3144 5038 3178
rect 5004 3076 5038 3110
rect 5004 3008 5038 3042
rect 5004 2940 5038 2974
rect 5004 2872 5038 2906
rect 5004 2804 5038 2838
rect 5004 2736 5038 2770
rect 5004 2668 5038 2702
rect 5004 2600 5038 2634
rect 5004 2532 5038 2566
rect 5004 2464 5038 2498
rect 5004 2396 5038 2430
rect 5004 2328 5038 2362
rect 5004 2260 5038 2294
rect 5004 2192 5038 2226
rect 5004 2124 5038 2158
rect 5004 2056 5038 2090
rect 5004 1988 5038 2022
rect 5004 1855 5038 1954
rect 5004 1763 5038 1821
rect 7519 16383 7553 16438
rect 7519 16315 7553 16349
rect 7519 16247 7553 16281
rect 7519 16179 7553 16213
rect 7519 16111 7553 16145
rect 7519 16043 7553 16077
rect 7519 15975 7553 16009
rect 7519 15907 7553 15941
rect 7519 15839 7553 15873
rect 7519 15771 7553 15805
rect 7519 15703 7553 15737
rect 7519 15635 7553 15669
rect 7519 15567 7553 15601
rect 7519 15499 7553 15533
rect 7519 15431 7553 15465
rect 7519 15363 7553 15397
rect 7519 15295 7553 15329
rect 7519 15227 7553 15261
rect 7519 15159 7553 15193
rect 7519 15091 7553 15125
rect 7519 15023 7553 15057
rect 7519 14955 7553 14989
rect 7519 14887 7553 14921
rect 7519 14819 7553 14853
rect 7519 14751 7553 14785
rect 7519 14683 7553 14717
rect 7519 14615 7553 14649
rect 7519 14547 7553 14581
rect 7519 14479 7553 14513
rect 7519 14411 7553 14445
rect 7519 14343 7553 14377
rect 7519 14275 7553 14309
rect 7519 14207 7553 14241
rect 7519 14139 7553 14173
rect 7519 14071 7553 14105
rect 7519 14003 7553 14037
rect 7519 13935 7553 13969
rect 7519 13867 7553 13901
rect 7519 13799 7553 13833
rect 7519 13731 7553 13765
rect 7519 13663 7553 13697
rect 7519 13595 7553 13629
rect 7519 13527 7553 13561
rect 7519 13459 7553 13493
rect 7519 13391 7553 13425
rect 7519 13323 7553 13357
rect 7519 13255 7553 13289
rect 7519 13187 7553 13221
rect 7519 13119 7553 13153
rect 7519 13051 7553 13085
rect 7519 12983 7553 13017
rect 7519 12915 7553 12949
rect 7519 12847 7553 12881
rect 7519 12779 7553 12813
rect 7519 12711 7553 12745
rect 7519 12643 7553 12677
rect 7519 12575 7553 12609
rect 7519 12507 7553 12541
rect 7519 12439 7553 12473
rect 7519 12371 7553 12405
rect 7519 12303 7553 12337
rect 7519 12235 7553 12269
rect 7519 12167 7553 12201
rect 7519 12099 7553 12133
rect 7519 12031 7553 12065
rect 7519 11963 7553 11997
rect 7519 11895 7553 11929
rect 7519 11827 7553 11861
rect 7519 11759 7553 11793
rect 7519 11691 7553 11725
rect 7519 11623 7553 11657
rect 7519 11555 7553 11589
rect 7519 11487 7553 11521
rect 7519 11419 7553 11453
rect 7519 11351 7553 11385
rect 7519 11283 7553 11317
rect 7519 11215 7553 11249
rect 7519 11147 7553 11181
rect 7519 11079 7553 11113
rect 7519 11011 7553 11045
rect 7519 10943 7553 10977
rect 7519 10875 7553 10909
rect 7519 10807 7553 10841
rect 7519 10739 7553 10773
rect 7519 10671 7553 10705
rect 7519 10603 7553 10637
rect 7519 10535 7553 10569
rect 7519 10467 7553 10501
rect 7519 10399 7553 10433
rect 7519 10331 7553 10365
rect 7519 10263 7553 10297
rect 7519 10195 7553 10229
rect 7519 10127 7553 10161
rect 7519 10059 7553 10093
rect 7519 9991 7553 10025
rect 7519 9923 7553 9957
rect 7519 9855 7553 9889
rect 7519 9787 7553 9821
rect 7519 9719 7553 9753
rect 7519 9651 7553 9685
rect 7519 9583 7553 9617
rect 7519 9515 7553 9549
rect 7519 9447 7553 9481
rect 7519 9379 7553 9413
rect 7519 9311 7553 9345
rect 7519 9243 7553 9277
rect 7519 9175 7553 9209
rect 7519 9107 7553 9141
rect 7519 9039 7553 9073
rect 7519 8971 7553 9005
rect 7519 8903 7553 8937
rect 7519 8835 7553 8869
rect 7519 8767 7553 8801
rect 7519 8699 7553 8733
rect 7519 8631 7553 8665
rect 7519 8563 7553 8597
rect 7519 8495 7553 8529
rect 7519 8427 7553 8461
rect 7519 8359 7553 8393
rect 7519 8291 7553 8325
rect 7519 8223 7553 8257
rect 7519 8155 7553 8189
rect 7519 8087 7553 8121
rect 7519 8019 7553 8053
rect 7519 7951 7553 7985
rect 7519 7883 7553 7917
rect 7519 7815 7553 7849
rect 7519 7747 7553 7781
rect 7519 7679 7553 7713
rect 7519 7611 7553 7645
rect 7519 7543 7553 7577
rect 7519 7475 7553 7509
rect 7519 7407 7553 7441
rect 7519 7339 7553 7373
rect 7519 7271 7553 7305
rect 7519 7203 7553 7237
rect 7519 7135 7553 7169
rect 7519 7067 7553 7101
rect 7519 6999 7553 7033
rect 7519 6931 7553 6965
rect 7519 6863 7553 6897
rect 7519 6795 7553 6829
rect 7519 6727 7553 6761
rect 7519 6659 7553 6693
rect 7519 6591 7553 6625
rect 7519 6523 7553 6557
rect 7519 6455 7553 6489
rect 7519 6387 7553 6421
rect 7519 6319 7553 6353
rect 7519 6251 7553 6285
rect 7519 6183 7553 6217
rect 7519 6115 7553 6149
rect 7519 6047 7553 6081
rect 7519 5979 7553 6013
rect 7519 5911 7553 5945
rect 7519 5843 7553 5877
rect 7519 5775 7553 5809
rect 7519 5707 7553 5741
rect 7519 5639 7553 5673
rect 7519 5571 7553 5605
rect 7519 5503 7553 5537
rect 7519 5435 7553 5469
rect 7519 5367 7553 5401
rect 7519 5299 7553 5333
rect 7519 5231 7553 5265
rect 7519 5163 7553 5197
rect 7519 5095 7553 5129
rect 7519 5027 7553 5061
rect 7519 4959 7553 4993
rect 7519 4891 7553 4925
rect 7519 4823 7553 4857
rect 7519 4755 7553 4789
rect 7519 4687 7553 4721
rect 7519 4619 7553 4653
rect 7519 4551 7553 4585
rect 7519 4483 7553 4517
rect 7519 4415 7553 4449
rect 7519 4347 7553 4381
rect 7519 4279 7553 4313
rect 7519 4211 7553 4245
rect 7519 4143 7553 4177
rect 7519 4075 7553 4109
rect 7519 4007 7553 4041
rect 7519 3939 7553 3973
rect 7519 3871 7553 3905
rect 7519 3803 7553 3837
rect 7519 3735 7553 3769
rect 7519 3667 7553 3701
rect 7519 3599 7553 3633
rect 7519 3531 7553 3565
rect 7519 3463 7553 3497
rect 7519 3395 7553 3429
rect 7519 3327 7553 3361
rect 7519 3259 7553 3293
rect 7519 3191 7553 3225
rect 7519 3123 7553 3157
rect 7519 3055 7553 3089
rect 7519 2987 7553 3021
rect 7519 2919 7553 2953
rect 7519 2851 7553 2885
rect 7519 2783 7553 2817
rect 7519 2715 7553 2749
rect 7519 2647 7553 2681
rect 7519 2579 7553 2613
rect 7519 2511 7553 2545
rect 7519 2443 7553 2477
rect 7519 2375 7553 2409
rect 7519 2307 7553 2341
rect 7519 2239 7553 2273
rect 7519 2171 7553 2205
rect 7519 2103 7553 2137
rect 7519 2035 7553 2069
rect 7519 1967 7553 2001
rect 7519 1899 7553 1933
rect 7519 1831 7553 1865
rect 7519 1763 7553 1797
rect 5004 1729 5072 1763
rect 5106 1729 5140 1763
rect 5174 1729 5208 1763
rect 5242 1729 5276 1763
rect 5310 1729 5344 1763
rect 5378 1729 5412 1763
rect 5446 1729 5480 1763
rect 5514 1729 5548 1763
rect 5582 1729 5616 1763
rect 5650 1729 5684 1763
rect 5718 1729 5752 1763
rect 5786 1729 5820 1763
rect 5854 1729 5888 1763
rect 5922 1729 5956 1763
rect 5990 1729 6024 1763
rect 6058 1729 6092 1763
rect 6126 1729 6160 1763
rect 6194 1729 6228 1763
rect 6262 1729 6296 1763
rect 6330 1729 6364 1763
rect 6398 1729 6432 1763
rect 6466 1729 6500 1763
rect 6534 1729 6568 1763
rect 6602 1729 6636 1763
rect 6670 1729 6704 1763
rect 6738 1729 6772 1763
rect 6806 1729 6840 1763
rect 6874 1729 6908 1763
rect 6942 1729 6976 1763
rect 7010 1729 7044 1763
rect 7078 1729 7112 1763
rect 7146 1729 7180 1763
rect 7214 1729 7248 1763
rect 7282 1729 7316 1763
rect 7350 1729 7384 1763
rect 7418 1729 7553 1763
<< psubdiffcont >>
rect 325 39917 359 39951
rect 461 39917 495 39951
rect 597 39917 631 39951
rect 733 39917 767 39951
rect 869 39917 903 39951
rect 1005 39917 1039 39951
rect 1141 39917 1175 39951
rect 1277 39917 1311 39951
rect 1413 39917 1447 39951
rect 1549 39917 1583 39951
rect 1685 39917 1719 39951
rect 325 39781 359 39815
rect 461 39781 495 39815
rect 597 39781 631 39815
rect 733 39781 767 39815
rect 869 39781 903 39815
rect 1005 39781 1039 39815
rect 1141 39781 1175 39815
rect 1277 39781 1311 39815
rect 1413 39781 1447 39815
rect 1549 39781 1583 39815
rect 1685 39781 1719 39815
rect 325 39645 359 39679
rect 461 39645 495 39679
rect 597 39645 631 39679
rect 733 39645 767 39679
rect 869 39645 903 39679
rect 1005 39645 1039 39679
rect 1141 39645 1175 39679
rect 1277 39645 1311 39679
rect 1413 39645 1447 39679
rect 1549 39645 1583 39679
rect 1685 39645 1719 39679
rect 325 39509 359 39543
rect 461 39509 495 39543
rect 597 39509 631 39543
rect 733 39509 767 39543
rect 869 39509 903 39543
rect 1005 39509 1039 39543
rect 1141 39509 1175 39543
rect 1277 39509 1311 39543
rect 1413 39509 1447 39543
rect 1549 39509 1583 39543
rect 1685 39509 1719 39543
rect 325 39373 359 39407
rect 461 39373 495 39407
rect 597 39373 631 39407
rect 733 39373 767 39407
rect 869 39373 903 39407
rect 1005 39373 1039 39407
rect 1141 39373 1175 39407
rect 1277 39373 1311 39407
rect 1413 39373 1447 39407
rect 1549 39373 1583 39407
rect 1685 39373 1719 39407
rect 325 39237 359 39271
rect 461 39237 495 39271
rect 597 39237 631 39271
rect 733 39237 767 39271
rect 869 39237 903 39271
rect 1005 39237 1039 39271
rect 1141 39237 1175 39271
rect 1277 39237 1311 39271
rect 1413 39237 1447 39271
rect 1549 39237 1583 39271
rect 1685 39237 1719 39271
rect 325 39101 359 39135
rect 461 39101 495 39135
rect 597 39101 631 39135
rect 733 39101 767 39135
rect 869 39101 903 39135
rect 1005 39101 1039 39135
rect 1141 39101 1175 39135
rect 1277 39101 1311 39135
rect 1413 39101 1447 39135
rect 1549 39101 1583 39135
rect 1685 39101 1719 39135
rect 325 38965 359 38999
rect 461 38965 495 38999
rect 597 38965 631 38999
rect 733 38965 767 38999
rect 869 38965 903 38999
rect 1005 38965 1039 38999
rect 1141 38965 1175 38999
rect 1277 38965 1311 38999
rect 1413 38965 1447 38999
rect 1549 38965 1583 38999
rect 1685 38965 1719 38999
rect 325 38829 359 38863
rect 461 38829 495 38863
rect 597 38829 631 38863
rect 733 38829 767 38863
rect 869 38829 903 38863
rect 1005 38829 1039 38863
rect 1141 38829 1175 38863
rect 1277 38829 1311 38863
rect 1413 38829 1447 38863
rect 1549 38829 1583 38863
rect 1685 38829 1719 38863
rect 325 38693 359 38727
rect 461 38693 495 38727
rect 597 38693 631 38727
rect 733 38693 767 38727
rect 869 38693 903 38727
rect 1005 38693 1039 38727
rect 1141 38693 1175 38727
rect 1277 38693 1311 38727
rect 1413 38693 1447 38727
rect 1549 38693 1583 38727
rect 1685 38693 1719 38727
rect 325 38557 359 38591
rect 461 38557 495 38591
rect 597 38557 631 38591
rect 733 38557 767 38591
rect 869 38557 903 38591
rect 1005 38557 1039 38591
rect 1141 38557 1175 38591
rect 1277 38557 1311 38591
rect 1413 38557 1447 38591
rect 1549 38557 1583 38591
rect 1685 38557 1719 38591
rect 325 38421 359 38455
rect 461 38421 495 38455
rect 597 38421 631 38455
rect 733 38421 767 38455
rect 869 38421 903 38455
rect 1005 38421 1039 38455
rect 1141 38421 1175 38455
rect 1277 38421 1311 38455
rect 1413 38421 1447 38455
rect 1549 38421 1583 38455
rect 1685 38421 1719 38455
rect 325 38285 359 38319
rect 461 38285 495 38319
rect 597 38285 631 38319
rect 733 38285 767 38319
rect 869 38285 903 38319
rect 1005 38285 1039 38319
rect 1141 38285 1175 38319
rect 1277 38285 1311 38319
rect 1413 38285 1447 38319
rect 1549 38285 1583 38319
rect 1685 38285 1719 38319
rect 325 38149 359 38183
rect 461 38149 495 38183
rect 597 38149 631 38183
rect 733 38149 767 38183
rect 869 38149 903 38183
rect 1005 38149 1039 38183
rect 1141 38149 1175 38183
rect 1277 38149 1311 38183
rect 1413 38149 1447 38183
rect 1549 38149 1583 38183
rect 1685 38149 1719 38183
rect 325 38013 359 38047
rect 461 38013 495 38047
rect 597 38013 631 38047
rect 733 38013 767 38047
rect 869 38013 903 38047
rect 1005 38013 1039 38047
rect 1141 38013 1175 38047
rect 1277 38013 1311 38047
rect 1413 38013 1447 38047
rect 1549 38013 1583 38047
rect 1685 38013 1719 38047
rect 325 37877 359 37911
rect 461 37877 495 37911
rect 597 37877 631 37911
rect 733 37877 767 37911
rect 869 37877 903 37911
rect 1005 37877 1039 37911
rect 1141 37877 1175 37911
rect 1277 37877 1311 37911
rect 1413 37877 1447 37911
rect 1549 37877 1583 37911
rect 1685 37877 1719 37911
rect 325 37741 359 37775
rect 461 37741 495 37775
rect 597 37741 631 37775
rect 733 37741 767 37775
rect 869 37741 903 37775
rect 1005 37741 1039 37775
rect 1141 37741 1175 37775
rect 1277 37741 1311 37775
rect 1413 37741 1447 37775
rect 1549 37741 1583 37775
rect 1685 37741 1719 37775
rect 325 37605 359 37639
rect 461 37605 495 37639
rect 597 37605 631 37639
rect 733 37605 767 37639
rect 869 37605 903 37639
rect 1005 37605 1039 37639
rect 1141 37605 1175 37639
rect 1277 37605 1311 37639
rect 1413 37605 1447 37639
rect 1549 37605 1583 37639
rect 1685 37605 1719 37639
rect 325 37469 359 37503
rect 461 37469 495 37503
rect 597 37469 631 37503
rect 733 37469 767 37503
rect 869 37469 903 37503
rect 1005 37469 1039 37503
rect 1141 37469 1175 37503
rect 1277 37469 1311 37503
rect 1413 37469 1447 37503
rect 1549 37469 1583 37503
rect 1685 37469 1719 37503
rect 325 37333 359 37367
rect 461 37333 495 37367
rect 597 37333 631 37367
rect 733 37333 767 37367
rect 869 37333 903 37367
rect 1005 37333 1039 37367
rect 1141 37333 1175 37367
rect 1277 37333 1311 37367
rect 1413 37333 1447 37367
rect 1549 37333 1583 37367
rect 1685 37333 1719 37367
rect 325 37197 359 37231
rect 461 37197 495 37231
rect 597 37197 631 37231
rect 733 37197 767 37231
rect 869 37197 903 37231
rect 1005 37197 1039 37231
rect 1141 37197 1175 37231
rect 1277 37197 1311 37231
rect 1413 37197 1447 37231
rect 1549 37197 1583 37231
rect 1685 37197 1719 37231
rect 325 37061 359 37095
rect 461 37061 495 37095
rect 597 37061 631 37095
rect 733 37061 767 37095
rect 869 37061 903 37095
rect 1005 37061 1039 37095
rect 1141 37061 1175 37095
rect 1277 37061 1311 37095
rect 1413 37061 1447 37095
rect 1549 37061 1583 37095
rect 1685 37061 1719 37095
rect 325 36925 359 36959
rect 461 36925 495 36959
rect 597 36925 631 36959
rect 733 36925 767 36959
rect 869 36925 903 36959
rect 1005 36925 1039 36959
rect 1141 36925 1175 36959
rect 1277 36925 1311 36959
rect 1413 36925 1447 36959
rect 1549 36925 1583 36959
rect 1685 36925 1719 36959
rect 325 36789 359 36823
rect 461 36789 495 36823
rect 597 36789 631 36823
rect 733 36789 767 36823
rect 869 36789 903 36823
rect 1005 36789 1039 36823
rect 1141 36789 1175 36823
rect 1277 36789 1311 36823
rect 1413 36789 1447 36823
rect 1549 36789 1583 36823
rect 1685 36789 1719 36823
rect 325 36653 359 36687
rect 461 36653 495 36687
rect 597 36653 631 36687
rect 733 36653 767 36687
rect 869 36653 903 36687
rect 1005 36653 1039 36687
rect 1141 36653 1175 36687
rect 1277 36653 1311 36687
rect 1413 36653 1447 36687
rect 1549 36653 1583 36687
rect 1685 36653 1719 36687
rect 325 36517 359 36551
rect 461 36517 495 36551
rect 597 36517 631 36551
rect 733 36517 767 36551
rect 869 36517 903 36551
rect 1005 36517 1039 36551
rect 1141 36517 1175 36551
rect 1277 36517 1311 36551
rect 1413 36517 1447 36551
rect 1549 36517 1583 36551
rect 1685 36517 1719 36551
rect 325 36381 359 36415
rect 461 36381 495 36415
rect 597 36381 631 36415
rect 733 36381 767 36415
rect 869 36381 903 36415
rect 1005 36381 1039 36415
rect 1141 36381 1175 36415
rect 1277 36381 1311 36415
rect 1413 36381 1447 36415
rect 1549 36381 1583 36415
rect 1685 36381 1719 36415
rect 325 36245 359 36279
rect 461 36245 495 36279
rect 597 36245 631 36279
rect 733 36245 767 36279
rect 869 36245 903 36279
rect 1005 36245 1039 36279
rect 1141 36245 1175 36279
rect 1277 36245 1311 36279
rect 1413 36245 1447 36279
rect 1549 36245 1583 36279
rect 1685 36245 1719 36279
rect 325 36109 359 36143
rect 461 36109 495 36143
rect 597 36109 631 36143
rect 733 36109 767 36143
rect 869 36109 903 36143
rect 1005 36109 1039 36143
rect 1141 36109 1175 36143
rect 1277 36109 1311 36143
rect 1413 36109 1447 36143
rect 1549 36109 1583 36143
rect 1685 36109 1719 36143
rect 325 35973 359 36007
rect 461 35973 495 36007
rect 597 35973 631 36007
rect 733 35973 767 36007
rect 869 35973 903 36007
rect 1005 35973 1039 36007
rect 1141 35973 1175 36007
rect 1277 35973 1311 36007
rect 1413 35973 1447 36007
rect 1549 35973 1583 36007
rect 1685 35973 1719 36007
rect 325 35837 359 35871
rect 461 35837 495 35871
rect 597 35837 631 35871
rect 733 35837 767 35871
rect 869 35837 903 35871
rect 1005 35837 1039 35871
rect 1141 35837 1175 35871
rect 1277 35837 1311 35871
rect 1413 35837 1447 35871
rect 1549 35837 1583 35871
rect 1685 35837 1719 35871
rect 325 35701 359 35735
rect 461 35701 495 35735
rect 597 35701 631 35735
rect 733 35701 767 35735
rect 869 35701 903 35735
rect 1005 35701 1039 35735
rect 1141 35701 1175 35735
rect 1277 35701 1311 35735
rect 1413 35701 1447 35735
rect 1549 35701 1583 35735
rect 1685 35701 1719 35735
rect 325 35565 359 35599
rect 461 35565 495 35599
rect 597 35565 631 35599
rect 733 35565 767 35599
rect 869 35565 903 35599
rect 1005 35565 1039 35599
rect 1141 35565 1175 35599
rect 1277 35565 1311 35599
rect 1413 35565 1447 35599
rect 1549 35565 1583 35599
rect 1685 35565 1719 35599
rect 325 35429 359 35463
rect 461 35429 495 35463
rect 597 35429 631 35463
rect 733 35429 767 35463
rect 869 35429 903 35463
rect 1005 35429 1039 35463
rect 1141 35429 1175 35463
rect 1277 35429 1311 35463
rect 1413 35429 1447 35463
rect 1549 35429 1583 35463
rect 1685 35429 1719 35463
rect 325 35293 359 35327
rect 461 35293 495 35327
rect 597 35293 631 35327
rect 733 35293 767 35327
rect 869 35293 903 35327
rect 1005 35293 1039 35327
rect 1141 35293 1175 35327
rect 1277 35293 1311 35327
rect 1413 35293 1447 35327
rect 1549 35293 1583 35327
rect 1685 35293 1719 35327
rect 325 35157 359 35191
rect 461 35157 495 35191
rect 597 35157 631 35191
rect 733 35157 767 35191
rect 869 35157 903 35191
rect 1005 35157 1039 35191
rect 1141 35157 1175 35191
rect 1277 35157 1311 35191
rect 1413 35157 1447 35191
rect 1549 35157 1583 35191
rect 1685 35157 1719 35191
rect 325 35021 359 35055
rect 461 35021 495 35055
rect 597 35021 631 35055
rect 733 35021 767 35055
rect 869 35021 903 35055
rect 1005 35021 1039 35055
rect 1141 35021 1175 35055
rect 1277 35021 1311 35055
rect 1413 35021 1447 35055
rect 1549 35021 1583 35055
rect 1685 35021 1719 35055
rect 325 34885 359 34919
rect 461 34885 495 34919
rect 597 34885 631 34919
rect 733 34885 767 34919
rect 869 34885 903 34919
rect 1005 34885 1039 34919
rect 1141 34885 1175 34919
rect 1277 34885 1311 34919
rect 1413 34885 1447 34919
rect 1549 34885 1583 34919
rect 1685 34885 1719 34919
rect 325 34749 359 34783
rect 461 34749 495 34783
rect 597 34749 631 34783
rect 733 34749 767 34783
rect 869 34749 903 34783
rect 1005 34749 1039 34783
rect 1141 34749 1175 34783
rect 1277 34749 1311 34783
rect 1413 34749 1447 34783
rect 1549 34749 1583 34783
rect 1685 34749 1719 34783
rect 325 34613 359 34647
rect 461 34613 495 34647
rect 597 34613 631 34647
rect 733 34613 767 34647
rect 869 34613 903 34647
rect 1005 34613 1039 34647
rect 1141 34613 1175 34647
rect 1277 34613 1311 34647
rect 1413 34613 1447 34647
rect 1549 34613 1583 34647
rect 1685 34613 1719 34647
rect 325 34477 359 34511
rect 461 34477 495 34511
rect 597 34477 631 34511
rect 733 34477 767 34511
rect 869 34477 903 34511
rect 1005 34477 1039 34511
rect 1141 34477 1175 34511
rect 1277 34477 1311 34511
rect 1413 34477 1447 34511
rect 1549 34477 1583 34511
rect 1685 34477 1719 34511
rect 325 34341 359 34375
rect 461 34341 495 34375
rect 597 34341 631 34375
rect 733 34341 767 34375
rect 869 34341 903 34375
rect 1005 34341 1039 34375
rect 1141 34341 1175 34375
rect 1277 34341 1311 34375
rect 1413 34341 1447 34375
rect 1549 34341 1583 34375
rect 1685 34341 1719 34375
rect 325 34205 359 34239
rect 461 34205 495 34239
rect 597 34205 631 34239
rect 733 34205 767 34239
rect 869 34205 903 34239
rect 1005 34205 1039 34239
rect 1141 34205 1175 34239
rect 1277 34205 1311 34239
rect 1413 34205 1447 34239
rect 1549 34205 1583 34239
rect 1685 34205 1719 34239
rect 325 34069 359 34103
rect 461 34069 495 34103
rect 597 34069 631 34103
rect 733 34069 767 34103
rect 869 34069 903 34103
rect 1005 34069 1039 34103
rect 1141 34069 1175 34103
rect 1277 34069 1311 34103
rect 1413 34069 1447 34103
rect 1549 34069 1583 34103
rect 1685 34069 1719 34103
rect 325 33933 359 33967
rect 461 33933 495 33967
rect 597 33933 631 33967
rect 733 33933 767 33967
rect 869 33933 903 33967
rect 1005 33933 1039 33967
rect 1141 33933 1175 33967
rect 1277 33933 1311 33967
rect 1413 33933 1447 33967
rect 1549 33933 1583 33967
rect 1685 33933 1719 33967
rect 325 33797 359 33831
rect 461 33797 495 33831
rect 597 33797 631 33831
rect 733 33797 767 33831
rect 869 33797 903 33831
rect 1005 33797 1039 33831
rect 1141 33797 1175 33831
rect 1277 33797 1311 33831
rect 1413 33797 1447 33831
rect 1549 33797 1583 33831
rect 1685 33797 1719 33831
rect 325 33661 359 33695
rect 461 33661 495 33695
rect 597 33661 631 33695
rect 733 33661 767 33695
rect 869 33661 903 33695
rect 1005 33661 1039 33695
rect 1141 33661 1175 33695
rect 1277 33661 1311 33695
rect 1413 33661 1447 33695
rect 1549 33661 1583 33695
rect 1685 33661 1719 33695
rect 325 33525 359 33559
rect 461 33525 495 33559
rect 597 33525 631 33559
rect 733 33525 767 33559
rect 869 33525 903 33559
rect 1005 33525 1039 33559
rect 1141 33525 1175 33559
rect 1277 33525 1311 33559
rect 1413 33525 1447 33559
rect 1549 33525 1583 33559
rect 1685 33525 1719 33559
rect 325 33389 359 33423
rect 461 33389 495 33423
rect 597 33389 631 33423
rect 733 33389 767 33423
rect 869 33389 903 33423
rect 1005 33389 1039 33423
rect 1141 33389 1175 33423
rect 1277 33389 1311 33423
rect 1413 33389 1447 33423
rect 1549 33389 1583 33423
rect 1685 33389 1719 33423
rect 325 33253 359 33287
rect 461 33253 495 33287
rect 597 33253 631 33287
rect 733 33253 767 33287
rect 869 33253 903 33287
rect 1005 33253 1039 33287
rect 1141 33253 1175 33287
rect 1277 33253 1311 33287
rect 1413 33253 1447 33287
rect 1549 33253 1583 33287
rect 1685 33253 1719 33287
rect 325 33117 359 33151
rect 461 33117 495 33151
rect 597 33117 631 33151
rect 733 33117 767 33151
rect 869 33117 903 33151
rect 1005 33117 1039 33151
rect 1141 33117 1175 33151
rect 1277 33117 1311 33151
rect 1413 33117 1447 33151
rect 1549 33117 1583 33151
rect 1685 33117 1719 33151
rect 325 32981 359 33015
rect 461 32981 495 33015
rect 597 32981 631 33015
rect 733 32981 767 33015
rect 869 32981 903 33015
rect 1005 32981 1039 33015
rect 1141 32981 1175 33015
rect 1277 32981 1311 33015
rect 1413 32981 1447 33015
rect 1549 32981 1583 33015
rect 1685 32981 1719 33015
rect 325 32845 359 32879
rect 461 32845 495 32879
rect 597 32845 631 32879
rect 733 32845 767 32879
rect 869 32845 903 32879
rect 1005 32845 1039 32879
rect 1141 32845 1175 32879
rect 1277 32845 1311 32879
rect 1413 32845 1447 32879
rect 1549 32845 1583 32879
rect 1685 32845 1719 32879
rect 325 32709 359 32743
rect 461 32709 495 32743
rect 597 32709 631 32743
rect 733 32709 767 32743
rect 869 32709 903 32743
rect 1005 32709 1039 32743
rect 1141 32709 1175 32743
rect 1277 32709 1311 32743
rect 1413 32709 1447 32743
rect 1549 32709 1583 32743
rect 1685 32709 1719 32743
rect 325 32573 359 32607
rect 461 32573 495 32607
rect 597 32573 631 32607
rect 733 32573 767 32607
rect 869 32573 903 32607
rect 1005 32573 1039 32607
rect 1141 32573 1175 32607
rect 1277 32573 1311 32607
rect 1413 32573 1447 32607
rect 1549 32573 1583 32607
rect 1685 32573 1719 32607
rect 325 32437 359 32471
rect 461 32437 495 32471
rect 597 32437 631 32471
rect 733 32437 767 32471
rect 869 32437 903 32471
rect 1005 32437 1039 32471
rect 1141 32437 1175 32471
rect 1277 32437 1311 32471
rect 1413 32437 1447 32471
rect 1549 32437 1583 32471
rect 1685 32437 1719 32471
rect 325 32301 359 32335
rect 461 32301 495 32335
rect 597 32301 631 32335
rect 733 32301 767 32335
rect 869 32301 903 32335
rect 1005 32301 1039 32335
rect 1141 32301 1175 32335
rect 1277 32301 1311 32335
rect 1413 32301 1447 32335
rect 1549 32301 1583 32335
rect 1685 32301 1719 32335
rect 325 32165 359 32199
rect 461 32165 495 32199
rect 597 32165 631 32199
rect 733 32165 767 32199
rect 869 32165 903 32199
rect 1005 32165 1039 32199
rect 1141 32165 1175 32199
rect 1277 32165 1311 32199
rect 1413 32165 1447 32199
rect 1549 32165 1583 32199
rect 1685 32165 1719 32199
rect 325 32029 359 32063
rect 461 32029 495 32063
rect 597 32029 631 32063
rect 733 32029 767 32063
rect 869 32029 903 32063
rect 1005 32029 1039 32063
rect 1141 32029 1175 32063
rect 1277 32029 1311 32063
rect 1413 32029 1447 32063
rect 1549 32029 1583 32063
rect 1685 32029 1719 32063
rect 325 31893 359 31927
rect 461 31893 495 31927
rect 597 31893 631 31927
rect 733 31893 767 31927
rect 869 31893 903 31927
rect 1005 31893 1039 31927
rect 1141 31893 1175 31927
rect 1277 31893 1311 31927
rect 1413 31893 1447 31927
rect 1549 31893 1583 31927
rect 1685 31893 1719 31927
rect 325 31757 359 31791
rect 461 31757 495 31791
rect 597 31757 631 31791
rect 733 31757 767 31791
rect 869 31757 903 31791
rect 1005 31757 1039 31791
rect 1141 31757 1175 31791
rect 1277 31757 1311 31791
rect 1413 31757 1447 31791
rect 1549 31757 1583 31791
rect 1685 31757 1719 31791
rect 325 31621 359 31655
rect 461 31621 495 31655
rect 597 31621 631 31655
rect 733 31621 767 31655
rect 869 31621 903 31655
rect 1005 31621 1039 31655
rect 1141 31621 1175 31655
rect 1277 31621 1311 31655
rect 1413 31621 1447 31655
rect 1549 31621 1583 31655
rect 1685 31621 1719 31655
rect 325 31485 359 31519
rect 461 31485 495 31519
rect 597 31485 631 31519
rect 733 31485 767 31519
rect 869 31485 903 31519
rect 1005 31485 1039 31519
rect 1141 31485 1175 31519
rect 1277 31485 1311 31519
rect 1413 31485 1447 31519
rect 1549 31485 1583 31519
rect 1685 31485 1719 31519
rect 325 31349 359 31383
rect 461 31349 495 31383
rect 597 31349 631 31383
rect 733 31349 767 31383
rect 869 31349 903 31383
rect 1005 31349 1039 31383
rect 1141 31349 1175 31383
rect 1277 31349 1311 31383
rect 1413 31349 1447 31383
rect 1549 31349 1583 31383
rect 1685 31349 1719 31383
rect 325 31213 359 31247
rect 461 31213 495 31247
rect 597 31213 631 31247
rect 733 31213 767 31247
rect 869 31213 903 31247
rect 1005 31213 1039 31247
rect 1141 31213 1175 31247
rect 1277 31213 1311 31247
rect 1413 31213 1447 31247
rect 1549 31213 1583 31247
rect 1685 31213 1719 31247
rect 325 31077 359 31111
rect 461 31077 495 31111
rect 597 31077 631 31111
rect 733 31077 767 31111
rect 869 31077 903 31111
rect 1005 31077 1039 31111
rect 1141 31077 1175 31111
rect 1277 31077 1311 31111
rect 1413 31077 1447 31111
rect 1549 31077 1583 31111
rect 1685 31077 1719 31111
rect 325 30941 359 30975
rect 461 30941 495 30975
rect 597 30941 631 30975
rect 733 30941 767 30975
rect 869 30941 903 30975
rect 1005 30941 1039 30975
rect 1141 30941 1175 30975
rect 1277 30941 1311 30975
rect 1413 30941 1447 30975
rect 1549 30941 1583 30975
rect 1685 30941 1719 30975
rect 325 30805 359 30839
rect 461 30805 495 30839
rect 597 30805 631 30839
rect 733 30805 767 30839
rect 869 30805 903 30839
rect 1005 30805 1039 30839
rect 1141 30805 1175 30839
rect 1277 30805 1311 30839
rect 1413 30805 1447 30839
rect 1549 30805 1583 30839
rect 1685 30805 1719 30839
rect 325 30669 359 30703
rect 461 30669 495 30703
rect 597 30669 631 30703
rect 733 30669 767 30703
rect 869 30669 903 30703
rect 1005 30669 1039 30703
rect 1141 30669 1175 30703
rect 1277 30669 1311 30703
rect 1413 30669 1447 30703
rect 1549 30669 1583 30703
rect 1685 30669 1719 30703
rect 325 30533 359 30567
rect 461 30533 495 30567
rect 597 30533 631 30567
rect 733 30533 767 30567
rect 869 30533 903 30567
rect 1005 30533 1039 30567
rect 1141 30533 1175 30567
rect 1277 30533 1311 30567
rect 1413 30533 1447 30567
rect 1549 30533 1583 30567
rect 1685 30533 1719 30567
rect 325 30397 359 30431
rect 461 30397 495 30431
rect 597 30397 631 30431
rect 733 30397 767 30431
rect 869 30397 903 30431
rect 1005 30397 1039 30431
rect 1141 30397 1175 30431
rect 1277 30397 1311 30431
rect 1413 30397 1447 30431
rect 1549 30397 1583 30431
rect 1685 30397 1719 30431
rect 325 30261 359 30295
rect 461 30261 495 30295
rect 597 30261 631 30295
rect 733 30261 767 30295
rect 869 30261 903 30295
rect 1005 30261 1039 30295
rect 1141 30261 1175 30295
rect 1277 30261 1311 30295
rect 1413 30261 1447 30295
rect 1549 30261 1583 30295
rect 1685 30261 1719 30295
rect 325 30125 359 30159
rect 461 30125 495 30159
rect 597 30125 631 30159
rect 733 30125 767 30159
rect 869 30125 903 30159
rect 1005 30125 1039 30159
rect 1141 30125 1175 30159
rect 1277 30125 1311 30159
rect 1413 30125 1447 30159
rect 1549 30125 1583 30159
rect 1685 30125 1719 30159
rect 325 29989 359 30023
rect 461 29989 495 30023
rect 597 29989 631 30023
rect 733 29989 767 30023
rect 869 29989 903 30023
rect 1005 29989 1039 30023
rect 1141 29989 1175 30023
rect 1277 29989 1311 30023
rect 1413 29989 1447 30023
rect 1549 29989 1583 30023
rect 1685 29989 1719 30023
rect 325 29853 359 29887
rect 461 29853 495 29887
rect 597 29853 631 29887
rect 733 29853 767 29887
rect 869 29853 903 29887
rect 1005 29853 1039 29887
rect 1141 29853 1175 29887
rect 1277 29853 1311 29887
rect 1413 29853 1447 29887
rect 1549 29853 1583 29887
rect 1685 29853 1719 29887
rect 325 29717 359 29751
rect 461 29717 495 29751
rect 597 29717 631 29751
rect 733 29717 767 29751
rect 869 29717 903 29751
rect 1005 29717 1039 29751
rect 1141 29717 1175 29751
rect 1277 29717 1311 29751
rect 1413 29717 1447 29751
rect 1549 29717 1583 29751
rect 1685 29717 1719 29751
rect 325 29581 359 29615
rect 461 29581 495 29615
rect 597 29581 631 29615
rect 733 29581 767 29615
rect 869 29581 903 29615
rect 1005 29581 1039 29615
rect 1141 29581 1175 29615
rect 1277 29581 1311 29615
rect 1413 29581 1447 29615
rect 1549 29581 1583 29615
rect 1685 29581 1719 29615
rect 325 29445 359 29479
rect 461 29445 495 29479
rect 597 29445 631 29479
rect 733 29445 767 29479
rect 869 29445 903 29479
rect 1005 29445 1039 29479
rect 1141 29445 1175 29479
rect 1277 29445 1311 29479
rect 1413 29445 1447 29479
rect 1549 29445 1583 29479
rect 1685 29445 1719 29479
rect 325 29309 359 29343
rect 461 29309 495 29343
rect 597 29309 631 29343
rect 733 29309 767 29343
rect 869 29309 903 29343
rect 1005 29309 1039 29343
rect 1141 29309 1175 29343
rect 1277 29309 1311 29343
rect 1413 29309 1447 29343
rect 1549 29309 1583 29343
rect 1685 29309 1719 29343
rect 325 29173 359 29207
rect 461 29173 495 29207
rect 597 29173 631 29207
rect 733 29173 767 29207
rect 869 29173 903 29207
rect 1005 29173 1039 29207
rect 1141 29173 1175 29207
rect 1277 29173 1311 29207
rect 1413 29173 1447 29207
rect 1549 29173 1583 29207
rect 1685 29173 1719 29207
rect 325 29037 359 29071
rect 461 29037 495 29071
rect 597 29037 631 29071
rect 733 29037 767 29071
rect 869 29037 903 29071
rect 1005 29037 1039 29071
rect 1141 29037 1175 29071
rect 1277 29037 1311 29071
rect 1413 29037 1447 29071
rect 1549 29037 1583 29071
rect 1685 29037 1719 29071
rect 325 28901 359 28935
rect 461 28901 495 28935
rect 597 28901 631 28935
rect 733 28901 767 28935
rect 869 28901 903 28935
rect 1005 28901 1039 28935
rect 1141 28901 1175 28935
rect 1277 28901 1311 28935
rect 1413 28901 1447 28935
rect 1549 28901 1583 28935
rect 1685 28901 1719 28935
rect 325 28765 359 28799
rect 461 28765 495 28799
rect 597 28765 631 28799
rect 733 28765 767 28799
rect 869 28765 903 28799
rect 1005 28765 1039 28799
rect 1141 28765 1175 28799
rect 1277 28765 1311 28799
rect 1413 28765 1447 28799
rect 1549 28765 1583 28799
rect 1685 28765 1719 28799
rect 325 28629 359 28663
rect 461 28629 495 28663
rect 597 28629 631 28663
rect 733 28629 767 28663
rect 869 28629 903 28663
rect 1005 28629 1039 28663
rect 1141 28629 1175 28663
rect 1277 28629 1311 28663
rect 1413 28629 1447 28663
rect 1549 28629 1583 28663
rect 1685 28629 1719 28663
rect 325 28493 359 28527
rect 461 28493 495 28527
rect 597 28493 631 28527
rect 733 28493 767 28527
rect 869 28493 903 28527
rect 1005 28493 1039 28527
rect 1141 28493 1175 28527
rect 1277 28493 1311 28527
rect 1413 28493 1447 28527
rect 1549 28493 1583 28527
rect 1685 28493 1719 28527
rect 325 28357 359 28391
rect 461 28357 495 28391
rect 597 28357 631 28391
rect 733 28357 767 28391
rect 869 28357 903 28391
rect 1005 28357 1039 28391
rect 1141 28357 1175 28391
rect 1277 28357 1311 28391
rect 1413 28357 1447 28391
rect 1549 28357 1583 28391
rect 1685 28357 1719 28391
rect 325 28221 359 28255
rect 461 28221 495 28255
rect 597 28221 631 28255
rect 733 28221 767 28255
rect 869 28221 903 28255
rect 1005 28221 1039 28255
rect 1141 28221 1175 28255
rect 1277 28221 1311 28255
rect 1413 28221 1447 28255
rect 1549 28221 1583 28255
rect 1685 28221 1719 28255
rect 325 28085 359 28119
rect 461 28085 495 28119
rect 597 28085 631 28119
rect 733 28085 767 28119
rect 869 28085 903 28119
rect 1005 28085 1039 28119
rect 1141 28085 1175 28119
rect 1277 28085 1311 28119
rect 1413 28085 1447 28119
rect 1549 28085 1583 28119
rect 1685 28085 1719 28119
rect 325 27949 359 27983
rect 461 27949 495 27983
rect 597 27949 631 27983
rect 733 27949 767 27983
rect 869 27949 903 27983
rect 1005 27949 1039 27983
rect 1141 27949 1175 27983
rect 1277 27949 1311 27983
rect 1413 27949 1447 27983
rect 1549 27949 1583 27983
rect 1685 27949 1719 27983
rect 325 27813 359 27847
rect 461 27813 495 27847
rect 597 27813 631 27847
rect 733 27813 767 27847
rect 869 27813 903 27847
rect 1005 27813 1039 27847
rect 1141 27813 1175 27847
rect 1277 27813 1311 27847
rect 1413 27813 1447 27847
rect 1549 27813 1583 27847
rect 1685 27813 1719 27847
rect 325 27677 359 27711
rect 461 27677 495 27711
rect 597 27677 631 27711
rect 733 27677 767 27711
rect 869 27677 903 27711
rect 1005 27677 1039 27711
rect 1141 27677 1175 27711
rect 1277 27677 1311 27711
rect 1413 27677 1447 27711
rect 1549 27677 1583 27711
rect 1685 27677 1719 27711
rect 325 27541 359 27575
rect 461 27541 495 27575
rect 597 27541 631 27575
rect 733 27541 767 27575
rect 869 27541 903 27575
rect 1005 27541 1039 27575
rect 1141 27541 1175 27575
rect 1277 27541 1311 27575
rect 1413 27541 1447 27575
rect 1549 27541 1583 27575
rect 1685 27541 1719 27575
rect 325 27405 359 27439
rect 461 27405 495 27439
rect 597 27405 631 27439
rect 733 27405 767 27439
rect 869 27405 903 27439
rect 1005 27405 1039 27439
rect 1141 27405 1175 27439
rect 1277 27405 1311 27439
rect 1413 27405 1447 27439
rect 1549 27405 1583 27439
rect 1685 27405 1719 27439
rect 325 27269 359 27303
rect 461 27269 495 27303
rect 597 27269 631 27303
rect 733 27269 767 27303
rect 869 27269 903 27303
rect 1005 27269 1039 27303
rect 1141 27269 1175 27303
rect 1277 27269 1311 27303
rect 1413 27269 1447 27303
rect 1549 27269 1583 27303
rect 1685 27269 1719 27303
rect 325 27133 359 27167
rect 461 27133 495 27167
rect 597 27133 631 27167
rect 733 27133 767 27167
rect 869 27133 903 27167
rect 1005 27133 1039 27167
rect 1141 27133 1175 27167
rect 1277 27133 1311 27167
rect 1413 27133 1447 27167
rect 1549 27133 1583 27167
rect 1685 27133 1719 27167
rect 325 26997 359 27031
rect 461 26997 495 27031
rect 597 26997 631 27031
rect 733 26997 767 27031
rect 869 26997 903 27031
rect 1005 26997 1039 27031
rect 1141 26997 1175 27031
rect 1277 26997 1311 27031
rect 1413 26997 1447 27031
rect 1549 26997 1583 27031
rect 1685 26997 1719 27031
rect 325 26861 359 26895
rect 461 26861 495 26895
rect 597 26861 631 26895
rect 733 26861 767 26895
rect 869 26861 903 26895
rect 1005 26861 1039 26895
rect 1141 26861 1175 26895
rect 1277 26861 1311 26895
rect 1413 26861 1447 26895
rect 1549 26861 1583 26895
rect 1685 26861 1719 26895
rect 325 26725 359 26759
rect 461 26725 495 26759
rect 597 26725 631 26759
rect 733 26725 767 26759
rect 869 26725 903 26759
rect 1005 26725 1039 26759
rect 1141 26725 1175 26759
rect 1277 26725 1311 26759
rect 1413 26725 1447 26759
rect 1549 26725 1583 26759
rect 1685 26725 1719 26759
rect 325 26589 359 26623
rect 461 26589 495 26623
rect 597 26589 631 26623
rect 733 26589 767 26623
rect 869 26589 903 26623
rect 1005 26589 1039 26623
rect 1141 26589 1175 26623
rect 1277 26589 1311 26623
rect 1413 26589 1447 26623
rect 1549 26589 1583 26623
rect 1685 26589 1719 26623
rect 325 26453 359 26487
rect 461 26453 495 26487
rect 597 26453 631 26487
rect 733 26453 767 26487
rect 869 26453 903 26487
rect 1005 26453 1039 26487
rect 1141 26453 1175 26487
rect 1277 26453 1311 26487
rect 1413 26453 1447 26487
rect 1549 26453 1583 26487
rect 1685 26453 1719 26487
rect 325 26317 359 26351
rect 461 26317 495 26351
rect 597 26317 631 26351
rect 733 26317 767 26351
rect 869 26317 903 26351
rect 1005 26317 1039 26351
rect 1141 26317 1175 26351
rect 1277 26317 1311 26351
rect 1413 26317 1447 26351
rect 1549 26317 1583 26351
rect 1685 26317 1719 26351
rect 325 26181 359 26215
rect 461 26181 495 26215
rect 597 26181 631 26215
rect 733 26181 767 26215
rect 869 26181 903 26215
rect 1005 26181 1039 26215
rect 1141 26181 1175 26215
rect 1277 26181 1311 26215
rect 1413 26181 1447 26215
rect 1549 26181 1583 26215
rect 1685 26181 1719 26215
rect 325 26045 359 26079
rect 461 26045 495 26079
rect 597 26045 631 26079
rect 733 26045 767 26079
rect 869 26045 903 26079
rect 1005 26045 1039 26079
rect 1141 26045 1175 26079
rect 1277 26045 1311 26079
rect 1413 26045 1447 26079
rect 1549 26045 1583 26079
rect 1685 26045 1719 26079
rect 325 25909 359 25943
rect 461 25909 495 25943
rect 597 25909 631 25943
rect 733 25909 767 25943
rect 869 25909 903 25943
rect 1005 25909 1039 25943
rect 1141 25909 1175 25943
rect 1277 25909 1311 25943
rect 1413 25909 1447 25943
rect 1549 25909 1583 25943
rect 1685 25909 1719 25943
rect 325 25773 359 25807
rect 461 25773 495 25807
rect 597 25773 631 25807
rect 733 25773 767 25807
rect 869 25773 903 25807
rect 1005 25773 1039 25807
rect 1141 25773 1175 25807
rect 1277 25773 1311 25807
rect 1413 25773 1447 25807
rect 1549 25773 1583 25807
rect 1685 25773 1719 25807
rect 325 25637 359 25671
rect 461 25637 495 25671
rect 597 25637 631 25671
rect 733 25637 767 25671
rect 869 25637 903 25671
rect 1005 25637 1039 25671
rect 1141 25637 1175 25671
rect 1277 25637 1311 25671
rect 1413 25637 1447 25671
rect 1549 25637 1583 25671
rect 1685 25637 1719 25671
rect 325 25501 359 25535
rect 461 25501 495 25535
rect 597 25501 631 25535
rect 733 25501 767 25535
rect 869 25501 903 25535
rect 1005 25501 1039 25535
rect 1141 25501 1175 25535
rect 1277 25501 1311 25535
rect 1413 25501 1447 25535
rect 1549 25501 1583 25535
rect 1685 25501 1719 25535
rect 325 25365 359 25399
rect 461 25365 495 25399
rect 597 25365 631 25399
rect 733 25365 767 25399
rect 869 25365 903 25399
rect 1005 25365 1039 25399
rect 1141 25365 1175 25399
rect 1277 25365 1311 25399
rect 1413 25365 1447 25399
rect 1549 25365 1583 25399
rect 1685 25365 1719 25399
rect 325 25229 359 25263
rect 461 25229 495 25263
rect 597 25229 631 25263
rect 733 25229 767 25263
rect 869 25229 903 25263
rect 1005 25229 1039 25263
rect 1141 25229 1175 25263
rect 1277 25229 1311 25263
rect 1413 25229 1447 25263
rect 1549 25229 1583 25263
rect 1685 25229 1719 25263
rect 325 25093 359 25127
rect 461 25093 495 25127
rect 597 25093 631 25127
rect 733 25093 767 25127
rect 869 25093 903 25127
rect 1005 25093 1039 25127
rect 1141 25093 1175 25127
rect 1277 25093 1311 25127
rect 1413 25093 1447 25127
rect 1549 25093 1583 25127
rect 1685 25093 1719 25127
rect 325 24957 359 24991
rect 461 24957 495 24991
rect 597 24957 631 24991
rect 733 24957 767 24991
rect 869 24957 903 24991
rect 1005 24957 1039 24991
rect 1141 24957 1175 24991
rect 1277 24957 1311 24991
rect 1413 24957 1447 24991
rect 1549 24957 1583 24991
rect 1685 24957 1719 24991
rect 325 24821 359 24855
rect 461 24821 495 24855
rect 597 24821 631 24855
rect 733 24821 767 24855
rect 869 24821 903 24855
rect 1005 24821 1039 24855
rect 1141 24821 1175 24855
rect 1277 24821 1311 24855
rect 1413 24821 1447 24855
rect 1549 24821 1583 24855
rect 1685 24821 1719 24855
rect 325 24685 359 24719
rect 461 24685 495 24719
rect 597 24685 631 24719
rect 733 24685 767 24719
rect 869 24685 903 24719
rect 1005 24685 1039 24719
rect 1141 24685 1175 24719
rect 1277 24685 1311 24719
rect 1413 24685 1447 24719
rect 1549 24685 1583 24719
rect 1685 24685 1719 24719
rect 325 24549 359 24583
rect 461 24549 495 24583
rect 597 24549 631 24583
rect 733 24549 767 24583
rect 869 24549 903 24583
rect 1005 24549 1039 24583
rect 1141 24549 1175 24583
rect 1277 24549 1311 24583
rect 1413 24549 1447 24583
rect 1549 24549 1583 24583
rect 1685 24549 1719 24583
rect 325 24413 359 24447
rect 461 24413 495 24447
rect 597 24413 631 24447
rect 733 24413 767 24447
rect 869 24413 903 24447
rect 1005 24413 1039 24447
rect 1141 24413 1175 24447
rect 1277 24413 1311 24447
rect 1413 24413 1447 24447
rect 1549 24413 1583 24447
rect 1685 24413 1719 24447
rect 325 24277 359 24311
rect 461 24277 495 24311
rect 597 24277 631 24311
rect 733 24277 767 24311
rect 869 24277 903 24311
rect 1005 24277 1039 24311
rect 1141 24277 1175 24311
rect 1277 24277 1311 24311
rect 1413 24277 1447 24311
rect 1549 24277 1583 24311
rect 1685 24277 1719 24311
rect 325 24141 359 24175
rect 461 24141 495 24175
rect 597 24141 631 24175
rect 733 24141 767 24175
rect 869 24141 903 24175
rect 1005 24141 1039 24175
rect 1141 24141 1175 24175
rect 1277 24141 1311 24175
rect 1413 24141 1447 24175
rect 1549 24141 1583 24175
rect 1685 24141 1719 24175
rect 325 24005 359 24039
rect 461 24005 495 24039
rect 597 24005 631 24039
rect 733 24005 767 24039
rect 869 24005 903 24039
rect 1005 24005 1039 24039
rect 1141 24005 1175 24039
rect 1277 24005 1311 24039
rect 1413 24005 1447 24039
rect 1549 24005 1583 24039
rect 1685 24005 1719 24039
rect 325 23869 359 23903
rect 461 23869 495 23903
rect 597 23869 631 23903
rect 733 23869 767 23903
rect 869 23869 903 23903
rect 1005 23869 1039 23903
rect 1141 23869 1175 23903
rect 1277 23869 1311 23903
rect 1413 23869 1447 23903
rect 1549 23869 1583 23903
rect 1685 23869 1719 23903
rect 325 23733 359 23767
rect 461 23733 495 23767
rect 597 23733 631 23767
rect 733 23733 767 23767
rect 869 23733 903 23767
rect 1005 23733 1039 23767
rect 1141 23733 1175 23767
rect 1277 23733 1311 23767
rect 1413 23733 1447 23767
rect 1549 23733 1583 23767
rect 1685 23733 1719 23767
rect 325 23597 359 23631
rect 461 23597 495 23631
rect 597 23597 631 23631
rect 733 23597 767 23631
rect 869 23597 903 23631
rect 1005 23597 1039 23631
rect 1141 23597 1175 23631
rect 1277 23597 1311 23631
rect 1413 23597 1447 23631
rect 1549 23597 1583 23631
rect 1685 23597 1719 23631
rect 325 23461 359 23495
rect 461 23461 495 23495
rect 597 23461 631 23495
rect 733 23461 767 23495
rect 869 23461 903 23495
rect 1005 23461 1039 23495
rect 1141 23461 1175 23495
rect 1277 23461 1311 23495
rect 1413 23461 1447 23495
rect 1549 23461 1583 23495
rect 1685 23461 1719 23495
rect 325 23325 359 23359
rect 461 23325 495 23359
rect 597 23325 631 23359
rect 733 23325 767 23359
rect 869 23325 903 23359
rect 1005 23325 1039 23359
rect 1141 23325 1175 23359
rect 1277 23325 1311 23359
rect 1413 23325 1447 23359
rect 1549 23325 1583 23359
rect 1685 23325 1719 23359
rect 325 23189 359 23223
rect 461 23189 495 23223
rect 597 23189 631 23223
rect 733 23189 767 23223
rect 869 23189 903 23223
rect 1005 23189 1039 23223
rect 1141 23189 1175 23223
rect 1277 23189 1311 23223
rect 1413 23189 1447 23223
rect 1549 23189 1583 23223
rect 1685 23189 1719 23223
rect 325 23053 359 23087
rect 461 23053 495 23087
rect 597 23053 631 23087
rect 733 23053 767 23087
rect 869 23053 903 23087
rect 1005 23053 1039 23087
rect 1141 23053 1175 23087
rect 1277 23053 1311 23087
rect 1413 23053 1447 23087
rect 1549 23053 1583 23087
rect 1685 23053 1719 23087
rect 325 22917 359 22951
rect 461 22917 495 22951
rect 597 22917 631 22951
rect 733 22917 767 22951
rect 869 22917 903 22951
rect 1005 22917 1039 22951
rect 1141 22917 1175 22951
rect 1277 22917 1311 22951
rect 1413 22917 1447 22951
rect 1549 22917 1583 22951
rect 1685 22917 1719 22951
rect 325 22781 359 22815
rect 461 22781 495 22815
rect 597 22781 631 22815
rect 733 22781 767 22815
rect 869 22781 903 22815
rect 1005 22781 1039 22815
rect 1141 22781 1175 22815
rect 1277 22781 1311 22815
rect 1413 22781 1447 22815
rect 1549 22781 1583 22815
rect 1685 22781 1719 22815
rect 325 22645 359 22679
rect 461 22645 495 22679
rect 597 22645 631 22679
rect 733 22645 767 22679
rect 869 22645 903 22679
rect 1005 22645 1039 22679
rect 1141 22645 1175 22679
rect 1277 22645 1311 22679
rect 1413 22645 1447 22679
rect 1549 22645 1583 22679
rect 1685 22645 1719 22679
rect 325 22509 359 22543
rect 461 22509 495 22543
rect 597 22509 631 22543
rect 733 22509 767 22543
rect 869 22509 903 22543
rect 1005 22509 1039 22543
rect 1141 22509 1175 22543
rect 1277 22509 1311 22543
rect 1413 22509 1447 22543
rect 1549 22509 1583 22543
rect 1685 22509 1719 22543
rect 325 22373 359 22407
rect 461 22373 495 22407
rect 597 22373 631 22407
rect 733 22373 767 22407
rect 869 22373 903 22407
rect 1005 22373 1039 22407
rect 1141 22373 1175 22407
rect 1277 22373 1311 22407
rect 1413 22373 1447 22407
rect 1549 22373 1583 22407
rect 1685 22373 1719 22407
rect 325 22237 359 22271
rect 461 22237 495 22271
rect 597 22237 631 22271
rect 733 22237 767 22271
rect 869 22237 903 22271
rect 1005 22237 1039 22271
rect 1141 22237 1175 22271
rect 1277 22237 1311 22271
rect 1413 22237 1447 22271
rect 1549 22237 1583 22271
rect 1685 22237 1719 22271
rect 325 22101 359 22135
rect 461 22101 495 22135
rect 597 22101 631 22135
rect 733 22101 767 22135
rect 869 22101 903 22135
rect 1005 22101 1039 22135
rect 1141 22101 1175 22135
rect 1277 22101 1311 22135
rect 1413 22101 1447 22135
rect 1549 22101 1583 22135
rect 1685 22101 1719 22135
rect 325 21965 359 21999
rect 461 21965 495 21999
rect 597 21965 631 21999
rect 733 21965 767 21999
rect 869 21965 903 21999
rect 1005 21965 1039 21999
rect 1141 21965 1175 21999
rect 1277 21965 1311 21999
rect 1413 21965 1447 21999
rect 1549 21965 1583 21999
rect 1685 21965 1719 21999
rect 325 21829 359 21863
rect 461 21829 495 21863
rect 597 21829 631 21863
rect 733 21829 767 21863
rect 869 21829 903 21863
rect 1005 21829 1039 21863
rect 1141 21829 1175 21863
rect 1277 21829 1311 21863
rect 1413 21829 1447 21863
rect 1549 21829 1583 21863
rect 1685 21829 1719 21863
rect 325 21693 359 21727
rect 461 21693 495 21727
rect 597 21693 631 21727
rect 733 21693 767 21727
rect 869 21693 903 21727
rect 1005 21693 1039 21727
rect 1141 21693 1175 21727
rect 1277 21693 1311 21727
rect 1413 21693 1447 21727
rect 1549 21693 1583 21727
rect 1685 21693 1719 21727
rect 325 21557 359 21591
rect 461 21557 495 21591
rect 597 21557 631 21591
rect 733 21557 767 21591
rect 869 21557 903 21591
rect 1005 21557 1039 21591
rect 1141 21557 1175 21591
rect 1277 21557 1311 21591
rect 1413 21557 1447 21591
rect 1549 21557 1583 21591
rect 1685 21557 1719 21591
rect 325 21421 359 21455
rect 461 21421 495 21455
rect 597 21421 631 21455
rect 733 21421 767 21455
rect 869 21421 903 21455
rect 1005 21421 1039 21455
rect 1141 21421 1175 21455
rect 1277 21421 1311 21455
rect 1413 21421 1447 21455
rect 1549 21421 1583 21455
rect 1685 21421 1719 21455
rect 325 21285 359 21319
rect 461 21285 495 21319
rect 597 21285 631 21319
rect 733 21285 767 21319
rect 869 21285 903 21319
rect 1005 21285 1039 21319
rect 1141 21285 1175 21319
rect 1277 21285 1311 21319
rect 1413 21285 1447 21319
rect 1549 21285 1583 21319
rect 1685 21285 1719 21319
rect 325 21149 359 21183
rect 461 21149 495 21183
rect 597 21149 631 21183
rect 733 21149 767 21183
rect 869 21149 903 21183
rect 1005 21149 1039 21183
rect 1141 21149 1175 21183
rect 1277 21149 1311 21183
rect 1413 21149 1447 21183
rect 1549 21149 1583 21183
rect 1685 21149 1719 21183
rect 325 21013 359 21047
rect 461 21013 495 21047
rect 597 21013 631 21047
rect 733 21013 767 21047
rect 869 21013 903 21047
rect 1005 21013 1039 21047
rect 1141 21013 1175 21047
rect 1277 21013 1311 21047
rect 1413 21013 1447 21047
rect 1549 21013 1583 21047
rect 1685 21013 1719 21047
rect 325 20877 359 20911
rect 461 20877 495 20911
rect 597 20877 631 20911
rect 733 20877 767 20911
rect 869 20877 903 20911
rect 1005 20877 1039 20911
rect 1141 20877 1175 20911
rect 1277 20877 1311 20911
rect 1413 20877 1447 20911
rect 1549 20877 1583 20911
rect 1685 20877 1719 20911
rect 325 20741 359 20775
rect 461 20741 495 20775
rect 597 20741 631 20775
rect 733 20741 767 20775
rect 869 20741 903 20775
rect 1005 20741 1039 20775
rect 1141 20741 1175 20775
rect 1277 20741 1311 20775
rect 1413 20741 1447 20775
rect 1549 20741 1583 20775
rect 1685 20741 1719 20775
rect 325 20605 359 20639
rect 461 20605 495 20639
rect 597 20605 631 20639
rect 733 20605 767 20639
rect 869 20605 903 20639
rect 1005 20605 1039 20639
rect 1141 20605 1175 20639
rect 1277 20605 1311 20639
rect 1413 20605 1447 20639
rect 1549 20605 1583 20639
rect 1685 20605 1719 20639
rect 325 20469 359 20503
rect 461 20469 495 20503
rect 597 20469 631 20503
rect 733 20469 767 20503
rect 869 20469 903 20503
rect 1005 20469 1039 20503
rect 1141 20469 1175 20503
rect 1277 20469 1311 20503
rect 1413 20469 1447 20503
rect 1549 20469 1583 20503
rect 1685 20469 1719 20503
rect 325 20333 359 20367
rect 461 20333 495 20367
rect 597 20333 631 20367
rect 733 20333 767 20367
rect 869 20333 903 20367
rect 1005 20333 1039 20367
rect 1141 20333 1175 20367
rect 1277 20333 1311 20367
rect 1413 20333 1447 20367
rect 1549 20333 1583 20367
rect 1685 20333 1719 20367
rect 325 20197 359 20231
rect 461 20197 495 20231
rect 597 20197 631 20231
rect 733 20197 767 20231
rect 869 20197 903 20231
rect 1005 20197 1039 20231
rect 1141 20197 1175 20231
rect 1277 20197 1311 20231
rect 1413 20197 1447 20231
rect 1549 20197 1583 20231
rect 1685 20197 1719 20231
rect 325 20061 359 20095
rect 461 20061 495 20095
rect 597 20061 631 20095
rect 733 20061 767 20095
rect 869 20061 903 20095
rect 1005 20061 1039 20095
rect 1141 20061 1175 20095
rect 1277 20061 1311 20095
rect 1413 20061 1447 20095
rect 1549 20061 1583 20095
rect 1685 20061 1719 20095
rect 325 19925 359 19959
rect 461 19925 495 19959
rect 597 19925 631 19959
rect 733 19925 767 19959
rect 869 19925 903 19959
rect 1005 19925 1039 19959
rect 1141 19925 1175 19959
rect 1277 19925 1311 19959
rect 1413 19925 1447 19959
rect 1549 19925 1583 19959
rect 1685 19925 1719 19959
rect 325 19789 359 19823
rect 461 19789 495 19823
rect 597 19789 631 19823
rect 733 19789 767 19823
rect 869 19789 903 19823
rect 1005 19789 1039 19823
rect 1141 19789 1175 19823
rect 1277 19789 1311 19823
rect 1413 19789 1447 19823
rect 1549 19789 1583 19823
rect 1685 19789 1719 19823
rect 325 19653 359 19687
rect 461 19653 495 19687
rect 597 19653 631 19687
rect 733 19653 767 19687
rect 869 19653 903 19687
rect 1005 19653 1039 19687
rect 1141 19653 1175 19687
rect 1277 19653 1311 19687
rect 1413 19653 1447 19687
rect 1549 19653 1583 19687
rect 1685 19653 1719 19687
rect 325 19517 359 19551
rect 461 19517 495 19551
rect 597 19517 631 19551
rect 733 19517 767 19551
rect 869 19517 903 19551
rect 1005 19517 1039 19551
rect 1141 19517 1175 19551
rect 1277 19517 1311 19551
rect 1413 19517 1447 19551
rect 1549 19517 1583 19551
rect 1685 19517 1719 19551
rect 325 19381 359 19415
rect 461 19381 495 19415
rect 597 19381 631 19415
rect 733 19381 767 19415
rect 869 19381 903 19415
rect 1005 19381 1039 19415
rect 1141 19381 1175 19415
rect 1277 19381 1311 19415
rect 1413 19381 1447 19415
rect 1549 19381 1583 19415
rect 1685 19381 1719 19415
rect 325 19245 359 19279
rect 461 19245 495 19279
rect 597 19245 631 19279
rect 733 19245 767 19279
rect 869 19245 903 19279
rect 1005 19245 1039 19279
rect 1141 19245 1175 19279
rect 1277 19245 1311 19279
rect 1413 19245 1447 19279
rect 1549 19245 1583 19279
rect 1685 19245 1719 19279
rect 325 19109 359 19143
rect 461 19109 495 19143
rect 597 19109 631 19143
rect 733 19109 767 19143
rect 869 19109 903 19143
rect 1005 19109 1039 19143
rect 1141 19109 1175 19143
rect 1277 19109 1311 19143
rect 1413 19109 1447 19143
rect 1549 19109 1583 19143
rect 1685 19109 1719 19143
rect 325 18973 359 19007
rect 461 18973 495 19007
rect 597 18973 631 19007
rect 733 18973 767 19007
rect 869 18973 903 19007
rect 1005 18973 1039 19007
rect 1141 18973 1175 19007
rect 1277 18973 1311 19007
rect 1413 18973 1447 19007
rect 1549 18973 1583 19007
rect 1685 18973 1719 19007
rect 325 18837 359 18871
rect 461 18837 495 18871
rect 597 18837 631 18871
rect 733 18837 767 18871
rect 869 18837 903 18871
rect 1005 18837 1039 18871
rect 1141 18837 1175 18871
rect 1277 18837 1311 18871
rect 1413 18837 1447 18871
rect 1549 18837 1583 18871
rect 1685 18837 1719 18871
rect 325 18701 359 18735
rect 461 18701 495 18735
rect 597 18701 631 18735
rect 733 18701 767 18735
rect 869 18701 903 18735
rect 1005 18701 1039 18735
rect 1141 18701 1175 18735
rect 1277 18701 1311 18735
rect 1413 18701 1447 18735
rect 1549 18701 1583 18735
rect 1685 18701 1719 18735
rect 325 18565 359 18599
rect 461 18565 495 18599
rect 597 18565 631 18599
rect 733 18565 767 18599
rect 869 18565 903 18599
rect 1005 18565 1039 18599
rect 1141 18565 1175 18599
rect 1277 18565 1311 18599
rect 1413 18565 1447 18599
rect 1549 18565 1583 18599
rect 1685 18565 1719 18599
rect 325 18429 359 18463
rect 461 18429 495 18463
rect 597 18429 631 18463
rect 733 18429 767 18463
rect 869 18429 903 18463
rect 1005 18429 1039 18463
rect 1141 18429 1175 18463
rect 1277 18429 1311 18463
rect 1413 18429 1447 18463
rect 1549 18429 1583 18463
rect 1685 18429 1719 18463
rect 325 18293 359 18327
rect 461 18293 495 18327
rect 597 18293 631 18327
rect 733 18293 767 18327
rect 869 18293 903 18327
rect 1005 18293 1039 18327
rect 1141 18293 1175 18327
rect 1277 18293 1311 18327
rect 1413 18293 1447 18327
rect 1549 18293 1583 18327
rect 1685 18293 1719 18327
rect 325 18157 359 18191
rect 461 18157 495 18191
rect 597 18157 631 18191
rect 733 18157 767 18191
rect 869 18157 903 18191
rect 1005 18157 1039 18191
rect 1141 18157 1175 18191
rect 1277 18157 1311 18191
rect 1413 18157 1447 18191
rect 1549 18157 1583 18191
rect 1685 18157 1719 18191
rect 325 18021 359 18055
rect 461 18021 495 18055
rect 597 18021 631 18055
rect 733 18021 767 18055
rect 869 18021 903 18055
rect 1005 18021 1039 18055
rect 1141 18021 1175 18055
rect 1277 18021 1311 18055
rect 1413 18021 1447 18055
rect 1549 18021 1583 18055
rect 1685 18021 1719 18055
rect 325 17885 359 17919
rect 461 17885 495 17919
rect 597 17885 631 17919
rect 733 17885 767 17919
rect 869 17885 903 17919
rect 1005 17885 1039 17919
rect 1141 17885 1175 17919
rect 1277 17885 1311 17919
rect 1413 17885 1447 17919
rect 1549 17885 1583 17919
rect 1685 17885 1719 17919
rect 325 17749 359 17783
rect 461 17749 495 17783
rect 597 17749 631 17783
rect 733 17749 767 17783
rect 869 17749 903 17783
rect 1005 17749 1039 17783
rect 1141 17749 1175 17783
rect 1277 17749 1311 17783
rect 1413 17749 1447 17783
rect 1549 17749 1583 17783
rect 1685 17749 1719 17783
rect 325 17613 359 17647
rect 461 17613 495 17647
rect 597 17613 631 17647
rect 733 17613 767 17647
rect 869 17613 903 17647
rect 1005 17613 1039 17647
rect 1141 17613 1175 17647
rect 1277 17613 1311 17647
rect 1413 17613 1447 17647
rect 1549 17613 1583 17647
rect 1685 17613 1719 17647
rect 325 17477 359 17511
rect 461 17477 495 17511
rect 597 17477 631 17511
rect 733 17477 767 17511
rect 869 17477 903 17511
rect 1005 17477 1039 17511
rect 1141 17477 1175 17511
rect 1277 17477 1311 17511
rect 1413 17477 1447 17511
rect 1549 17477 1583 17511
rect 1685 17477 1719 17511
rect 325 17341 359 17375
rect 461 17341 495 17375
rect 597 17341 631 17375
rect 733 17341 767 17375
rect 869 17341 903 17375
rect 1005 17341 1039 17375
rect 1141 17341 1175 17375
rect 1277 17341 1311 17375
rect 1413 17341 1447 17375
rect 1549 17341 1583 17375
rect 1685 17341 1719 17375
rect 325 17205 359 17239
rect 461 17205 495 17239
rect 597 17205 631 17239
rect 733 17205 767 17239
rect 869 17205 903 17239
rect 1005 17205 1039 17239
rect 1141 17205 1175 17239
rect 1277 17205 1311 17239
rect 1413 17205 1447 17239
rect 1549 17205 1583 17239
rect 1685 17205 1719 17239
rect 325 17069 359 17103
rect 461 17069 495 17103
rect 597 17069 631 17103
rect 733 17069 767 17103
rect 869 17069 903 17103
rect 1005 17069 1039 17103
rect 1141 17069 1175 17103
rect 1277 17069 1311 17103
rect 1413 17069 1447 17103
rect 1549 17069 1583 17103
rect 1685 17069 1719 17103
rect 325 16933 359 16967
rect 461 16933 495 16967
rect 597 16933 631 16967
rect 733 16933 767 16967
rect 869 16933 903 16967
rect 1005 16933 1039 16967
rect 1141 16933 1175 16967
rect 1277 16933 1311 16967
rect 1413 16933 1447 16967
rect 1549 16933 1583 16967
rect 1685 16933 1719 16967
rect 325 16797 359 16831
rect 461 16797 495 16831
rect 597 16797 631 16831
rect 733 16797 767 16831
rect 869 16797 903 16831
rect 1005 16797 1039 16831
rect 1141 16797 1175 16831
rect 1277 16797 1311 16831
rect 1413 16797 1447 16831
rect 1549 16797 1583 16831
rect 1685 16797 1719 16831
rect 325 16661 359 16695
rect 461 16661 495 16695
rect 597 16661 631 16695
rect 733 16661 767 16695
rect 869 16661 903 16695
rect 1005 16661 1039 16695
rect 1141 16661 1175 16695
rect 1277 16661 1311 16695
rect 1413 16661 1447 16695
rect 1549 16661 1583 16695
rect 1685 16661 1719 16695
rect 325 16525 359 16559
rect 461 16525 495 16559
rect 597 16525 631 16559
rect 733 16525 767 16559
rect 869 16525 903 16559
rect 1005 16525 1039 16559
rect 1141 16525 1175 16559
rect 1277 16525 1311 16559
rect 1413 16525 1447 16559
rect 1549 16525 1583 16559
rect 1685 16525 1719 16559
rect 7880 39917 7914 39951
rect 8016 39917 8050 39951
rect 8152 39917 8186 39951
rect 8288 39917 8322 39951
rect 8424 39917 8458 39951
rect 8560 39917 8594 39951
rect 8696 39917 8730 39951
rect 8832 39917 8866 39951
rect 8968 39917 9002 39951
rect 9104 39917 9138 39951
rect 9240 39917 9274 39951
rect 7880 39781 7914 39815
rect 8016 39781 8050 39815
rect 8152 39781 8186 39815
rect 8288 39781 8322 39815
rect 8424 39781 8458 39815
rect 8560 39781 8594 39815
rect 8696 39781 8730 39815
rect 8832 39781 8866 39815
rect 8968 39781 9002 39815
rect 9104 39781 9138 39815
rect 9240 39781 9274 39815
rect 7880 39645 7914 39679
rect 8016 39645 8050 39679
rect 8152 39645 8186 39679
rect 8288 39645 8322 39679
rect 8424 39645 8458 39679
rect 8560 39645 8594 39679
rect 8696 39645 8730 39679
rect 8832 39645 8866 39679
rect 8968 39645 9002 39679
rect 9104 39645 9138 39679
rect 9240 39645 9274 39679
rect 7880 39509 7914 39543
rect 8016 39509 8050 39543
rect 8152 39509 8186 39543
rect 8288 39509 8322 39543
rect 8424 39509 8458 39543
rect 8560 39509 8594 39543
rect 8696 39509 8730 39543
rect 8832 39509 8866 39543
rect 8968 39509 9002 39543
rect 9104 39509 9138 39543
rect 9240 39509 9274 39543
rect 7880 39373 7914 39407
rect 8016 39373 8050 39407
rect 8152 39373 8186 39407
rect 8288 39373 8322 39407
rect 8424 39373 8458 39407
rect 8560 39373 8594 39407
rect 8696 39373 8730 39407
rect 8832 39373 8866 39407
rect 8968 39373 9002 39407
rect 9104 39373 9138 39407
rect 9240 39373 9274 39407
rect 7880 39237 7914 39271
rect 8016 39237 8050 39271
rect 8152 39237 8186 39271
rect 8288 39237 8322 39271
rect 8424 39237 8458 39271
rect 8560 39237 8594 39271
rect 8696 39237 8730 39271
rect 8832 39237 8866 39271
rect 8968 39237 9002 39271
rect 9104 39237 9138 39271
rect 9240 39237 9274 39271
rect 7880 39101 7914 39135
rect 8016 39101 8050 39135
rect 8152 39101 8186 39135
rect 8288 39101 8322 39135
rect 8424 39101 8458 39135
rect 8560 39101 8594 39135
rect 8696 39101 8730 39135
rect 8832 39101 8866 39135
rect 8968 39101 9002 39135
rect 9104 39101 9138 39135
rect 9240 39101 9274 39135
rect 7880 38965 7914 38999
rect 8016 38965 8050 38999
rect 8152 38965 8186 38999
rect 8288 38965 8322 38999
rect 8424 38965 8458 38999
rect 8560 38965 8594 38999
rect 8696 38965 8730 38999
rect 8832 38965 8866 38999
rect 8968 38965 9002 38999
rect 9104 38965 9138 38999
rect 9240 38965 9274 38999
rect 7880 38829 7914 38863
rect 8016 38829 8050 38863
rect 8152 38829 8186 38863
rect 8288 38829 8322 38863
rect 8424 38829 8458 38863
rect 8560 38829 8594 38863
rect 8696 38829 8730 38863
rect 8832 38829 8866 38863
rect 8968 38829 9002 38863
rect 9104 38829 9138 38863
rect 9240 38829 9274 38863
rect 7880 38693 7914 38727
rect 8016 38693 8050 38727
rect 8152 38693 8186 38727
rect 8288 38693 8322 38727
rect 8424 38693 8458 38727
rect 8560 38693 8594 38727
rect 8696 38693 8730 38727
rect 8832 38693 8866 38727
rect 8968 38693 9002 38727
rect 9104 38693 9138 38727
rect 9240 38693 9274 38727
rect 7880 38557 7914 38591
rect 8016 38557 8050 38591
rect 8152 38557 8186 38591
rect 8288 38557 8322 38591
rect 8424 38557 8458 38591
rect 8560 38557 8594 38591
rect 8696 38557 8730 38591
rect 8832 38557 8866 38591
rect 8968 38557 9002 38591
rect 9104 38557 9138 38591
rect 9240 38557 9274 38591
rect 7880 38421 7914 38455
rect 8016 38421 8050 38455
rect 8152 38421 8186 38455
rect 8288 38421 8322 38455
rect 8424 38421 8458 38455
rect 8560 38421 8594 38455
rect 8696 38421 8730 38455
rect 8832 38421 8866 38455
rect 8968 38421 9002 38455
rect 9104 38421 9138 38455
rect 9240 38421 9274 38455
rect 7880 38285 7914 38319
rect 8016 38285 8050 38319
rect 8152 38285 8186 38319
rect 8288 38285 8322 38319
rect 8424 38285 8458 38319
rect 8560 38285 8594 38319
rect 8696 38285 8730 38319
rect 8832 38285 8866 38319
rect 8968 38285 9002 38319
rect 9104 38285 9138 38319
rect 9240 38285 9274 38319
rect 7880 38149 7914 38183
rect 8016 38149 8050 38183
rect 8152 38149 8186 38183
rect 8288 38149 8322 38183
rect 8424 38149 8458 38183
rect 8560 38149 8594 38183
rect 8696 38149 8730 38183
rect 8832 38149 8866 38183
rect 8968 38149 9002 38183
rect 9104 38149 9138 38183
rect 9240 38149 9274 38183
rect 7880 38013 7914 38047
rect 8016 38013 8050 38047
rect 8152 38013 8186 38047
rect 8288 38013 8322 38047
rect 8424 38013 8458 38047
rect 8560 38013 8594 38047
rect 8696 38013 8730 38047
rect 8832 38013 8866 38047
rect 8968 38013 9002 38047
rect 9104 38013 9138 38047
rect 9240 38013 9274 38047
rect 7880 37877 7914 37911
rect 8016 37877 8050 37911
rect 8152 37877 8186 37911
rect 8288 37877 8322 37911
rect 8424 37877 8458 37911
rect 8560 37877 8594 37911
rect 8696 37877 8730 37911
rect 8832 37877 8866 37911
rect 8968 37877 9002 37911
rect 9104 37877 9138 37911
rect 9240 37877 9274 37911
rect 7880 37741 7914 37775
rect 8016 37741 8050 37775
rect 8152 37741 8186 37775
rect 8288 37741 8322 37775
rect 8424 37741 8458 37775
rect 8560 37741 8594 37775
rect 8696 37741 8730 37775
rect 8832 37741 8866 37775
rect 8968 37741 9002 37775
rect 9104 37741 9138 37775
rect 9240 37741 9274 37775
rect 7880 37605 7914 37639
rect 8016 37605 8050 37639
rect 8152 37605 8186 37639
rect 8288 37605 8322 37639
rect 8424 37605 8458 37639
rect 8560 37605 8594 37639
rect 8696 37605 8730 37639
rect 8832 37605 8866 37639
rect 8968 37605 9002 37639
rect 9104 37605 9138 37639
rect 9240 37605 9274 37639
rect 7880 37469 7914 37503
rect 8016 37469 8050 37503
rect 8152 37469 8186 37503
rect 8288 37469 8322 37503
rect 8424 37469 8458 37503
rect 8560 37469 8594 37503
rect 8696 37469 8730 37503
rect 8832 37469 8866 37503
rect 8968 37469 9002 37503
rect 9104 37469 9138 37503
rect 9240 37469 9274 37503
rect 7880 37333 7914 37367
rect 8016 37333 8050 37367
rect 8152 37333 8186 37367
rect 8288 37333 8322 37367
rect 8424 37333 8458 37367
rect 8560 37333 8594 37367
rect 8696 37333 8730 37367
rect 8832 37333 8866 37367
rect 8968 37333 9002 37367
rect 9104 37333 9138 37367
rect 9240 37333 9274 37367
rect 7880 37197 7914 37231
rect 8016 37197 8050 37231
rect 8152 37197 8186 37231
rect 8288 37197 8322 37231
rect 8424 37197 8458 37231
rect 8560 37197 8594 37231
rect 8696 37197 8730 37231
rect 8832 37197 8866 37231
rect 8968 37197 9002 37231
rect 9104 37197 9138 37231
rect 9240 37197 9274 37231
rect 7880 37061 7914 37095
rect 8016 37061 8050 37095
rect 8152 37061 8186 37095
rect 8288 37061 8322 37095
rect 8424 37061 8458 37095
rect 8560 37061 8594 37095
rect 8696 37061 8730 37095
rect 8832 37061 8866 37095
rect 8968 37061 9002 37095
rect 9104 37061 9138 37095
rect 9240 37061 9274 37095
rect 7880 36925 7914 36959
rect 8016 36925 8050 36959
rect 8152 36925 8186 36959
rect 8288 36925 8322 36959
rect 8424 36925 8458 36959
rect 8560 36925 8594 36959
rect 8696 36925 8730 36959
rect 8832 36925 8866 36959
rect 8968 36925 9002 36959
rect 9104 36925 9138 36959
rect 9240 36925 9274 36959
rect 7880 36789 7914 36823
rect 8016 36789 8050 36823
rect 8152 36789 8186 36823
rect 8288 36789 8322 36823
rect 8424 36789 8458 36823
rect 8560 36789 8594 36823
rect 8696 36789 8730 36823
rect 8832 36789 8866 36823
rect 8968 36789 9002 36823
rect 9104 36789 9138 36823
rect 9240 36789 9274 36823
rect 7880 36653 7914 36687
rect 8016 36653 8050 36687
rect 8152 36653 8186 36687
rect 8288 36653 8322 36687
rect 8424 36653 8458 36687
rect 8560 36653 8594 36687
rect 8696 36653 8730 36687
rect 8832 36653 8866 36687
rect 8968 36653 9002 36687
rect 9104 36653 9138 36687
rect 9240 36653 9274 36687
rect 7880 36517 7914 36551
rect 8016 36517 8050 36551
rect 8152 36517 8186 36551
rect 8288 36517 8322 36551
rect 8424 36517 8458 36551
rect 8560 36517 8594 36551
rect 8696 36517 8730 36551
rect 8832 36517 8866 36551
rect 8968 36517 9002 36551
rect 9104 36517 9138 36551
rect 9240 36517 9274 36551
rect 7880 36381 7914 36415
rect 8016 36381 8050 36415
rect 8152 36381 8186 36415
rect 8288 36381 8322 36415
rect 8424 36381 8458 36415
rect 8560 36381 8594 36415
rect 8696 36381 8730 36415
rect 8832 36381 8866 36415
rect 8968 36381 9002 36415
rect 9104 36381 9138 36415
rect 9240 36381 9274 36415
rect 7880 36245 7914 36279
rect 8016 36245 8050 36279
rect 8152 36245 8186 36279
rect 8288 36245 8322 36279
rect 8424 36245 8458 36279
rect 8560 36245 8594 36279
rect 8696 36245 8730 36279
rect 8832 36245 8866 36279
rect 8968 36245 9002 36279
rect 9104 36245 9138 36279
rect 9240 36245 9274 36279
rect 7880 36109 7914 36143
rect 8016 36109 8050 36143
rect 8152 36109 8186 36143
rect 8288 36109 8322 36143
rect 8424 36109 8458 36143
rect 8560 36109 8594 36143
rect 8696 36109 8730 36143
rect 8832 36109 8866 36143
rect 8968 36109 9002 36143
rect 9104 36109 9138 36143
rect 9240 36109 9274 36143
rect 7880 35973 7914 36007
rect 8016 35973 8050 36007
rect 8152 35973 8186 36007
rect 8288 35973 8322 36007
rect 8424 35973 8458 36007
rect 8560 35973 8594 36007
rect 8696 35973 8730 36007
rect 8832 35973 8866 36007
rect 8968 35973 9002 36007
rect 9104 35973 9138 36007
rect 9240 35973 9274 36007
rect 7880 35837 7914 35871
rect 8016 35837 8050 35871
rect 8152 35837 8186 35871
rect 8288 35837 8322 35871
rect 8424 35837 8458 35871
rect 8560 35837 8594 35871
rect 8696 35837 8730 35871
rect 8832 35837 8866 35871
rect 8968 35837 9002 35871
rect 9104 35837 9138 35871
rect 9240 35837 9274 35871
rect 7880 35701 7914 35735
rect 8016 35701 8050 35735
rect 8152 35701 8186 35735
rect 8288 35701 8322 35735
rect 8424 35701 8458 35735
rect 8560 35701 8594 35735
rect 8696 35701 8730 35735
rect 8832 35701 8866 35735
rect 8968 35701 9002 35735
rect 9104 35701 9138 35735
rect 9240 35701 9274 35735
rect 7880 35565 7914 35599
rect 8016 35565 8050 35599
rect 8152 35565 8186 35599
rect 8288 35565 8322 35599
rect 8424 35565 8458 35599
rect 8560 35565 8594 35599
rect 8696 35565 8730 35599
rect 8832 35565 8866 35599
rect 8968 35565 9002 35599
rect 9104 35565 9138 35599
rect 9240 35565 9274 35599
rect 7880 35429 7914 35463
rect 8016 35429 8050 35463
rect 8152 35429 8186 35463
rect 8288 35429 8322 35463
rect 8424 35429 8458 35463
rect 8560 35429 8594 35463
rect 8696 35429 8730 35463
rect 8832 35429 8866 35463
rect 8968 35429 9002 35463
rect 9104 35429 9138 35463
rect 9240 35429 9274 35463
rect 7880 35293 7914 35327
rect 8016 35293 8050 35327
rect 8152 35293 8186 35327
rect 8288 35293 8322 35327
rect 8424 35293 8458 35327
rect 8560 35293 8594 35327
rect 8696 35293 8730 35327
rect 8832 35293 8866 35327
rect 8968 35293 9002 35327
rect 9104 35293 9138 35327
rect 9240 35293 9274 35327
rect 7880 35157 7914 35191
rect 8016 35157 8050 35191
rect 8152 35157 8186 35191
rect 8288 35157 8322 35191
rect 8424 35157 8458 35191
rect 8560 35157 8594 35191
rect 8696 35157 8730 35191
rect 8832 35157 8866 35191
rect 8968 35157 9002 35191
rect 9104 35157 9138 35191
rect 9240 35157 9274 35191
rect 7880 35021 7914 35055
rect 8016 35021 8050 35055
rect 8152 35021 8186 35055
rect 8288 35021 8322 35055
rect 8424 35021 8458 35055
rect 8560 35021 8594 35055
rect 8696 35021 8730 35055
rect 8832 35021 8866 35055
rect 8968 35021 9002 35055
rect 9104 35021 9138 35055
rect 9240 35021 9274 35055
rect 7880 34885 7914 34919
rect 8016 34885 8050 34919
rect 8152 34885 8186 34919
rect 8288 34885 8322 34919
rect 8424 34885 8458 34919
rect 8560 34885 8594 34919
rect 8696 34885 8730 34919
rect 8832 34885 8866 34919
rect 8968 34885 9002 34919
rect 9104 34885 9138 34919
rect 9240 34885 9274 34919
rect 7880 34749 7914 34783
rect 8016 34749 8050 34783
rect 8152 34749 8186 34783
rect 8288 34749 8322 34783
rect 8424 34749 8458 34783
rect 8560 34749 8594 34783
rect 8696 34749 8730 34783
rect 8832 34749 8866 34783
rect 8968 34749 9002 34783
rect 9104 34749 9138 34783
rect 9240 34749 9274 34783
rect 7880 34613 7914 34647
rect 8016 34613 8050 34647
rect 8152 34613 8186 34647
rect 8288 34613 8322 34647
rect 8424 34613 8458 34647
rect 8560 34613 8594 34647
rect 8696 34613 8730 34647
rect 8832 34613 8866 34647
rect 8968 34613 9002 34647
rect 9104 34613 9138 34647
rect 9240 34613 9274 34647
rect 7880 34477 7914 34511
rect 8016 34477 8050 34511
rect 8152 34477 8186 34511
rect 8288 34477 8322 34511
rect 8424 34477 8458 34511
rect 8560 34477 8594 34511
rect 8696 34477 8730 34511
rect 8832 34477 8866 34511
rect 8968 34477 9002 34511
rect 9104 34477 9138 34511
rect 9240 34477 9274 34511
rect 7880 34341 7914 34375
rect 8016 34341 8050 34375
rect 8152 34341 8186 34375
rect 8288 34341 8322 34375
rect 8424 34341 8458 34375
rect 8560 34341 8594 34375
rect 8696 34341 8730 34375
rect 8832 34341 8866 34375
rect 8968 34341 9002 34375
rect 9104 34341 9138 34375
rect 9240 34341 9274 34375
rect 7880 34205 7914 34239
rect 8016 34205 8050 34239
rect 8152 34205 8186 34239
rect 8288 34205 8322 34239
rect 8424 34205 8458 34239
rect 8560 34205 8594 34239
rect 8696 34205 8730 34239
rect 8832 34205 8866 34239
rect 8968 34205 9002 34239
rect 9104 34205 9138 34239
rect 9240 34205 9274 34239
rect 7880 34069 7914 34103
rect 8016 34069 8050 34103
rect 8152 34069 8186 34103
rect 8288 34069 8322 34103
rect 8424 34069 8458 34103
rect 8560 34069 8594 34103
rect 8696 34069 8730 34103
rect 8832 34069 8866 34103
rect 8968 34069 9002 34103
rect 9104 34069 9138 34103
rect 9240 34069 9274 34103
rect 7880 33933 7914 33967
rect 8016 33933 8050 33967
rect 8152 33933 8186 33967
rect 8288 33933 8322 33967
rect 8424 33933 8458 33967
rect 8560 33933 8594 33967
rect 8696 33933 8730 33967
rect 8832 33933 8866 33967
rect 8968 33933 9002 33967
rect 9104 33933 9138 33967
rect 9240 33933 9274 33967
rect 7880 33797 7914 33831
rect 8016 33797 8050 33831
rect 8152 33797 8186 33831
rect 8288 33797 8322 33831
rect 8424 33797 8458 33831
rect 8560 33797 8594 33831
rect 8696 33797 8730 33831
rect 8832 33797 8866 33831
rect 8968 33797 9002 33831
rect 9104 33797 9138 33831
rect 9240 33797 9274 33831
rect 7880 33661 7914 33695
rect 8016 33661 8050 33695
rect 8152 33661 8186 33695
rect 8288 33661 8322 33695
rect 8424 33661 8458 33695
rect 8560 33661 8594 33695
rect 8696 33661 8730 33695
rect 8832 33661 8866 33695
rect 8968 33661 9002 33695
rect 9104 33661 9138 33695
rect 9240 33661 9274 33695
rect 7880 33525 7914 33559
rect 8016 33525 8050 33559
rect 8152 33525 8186 33559
rect 8288 33525 8322 33559
rect 8424 33525 8458 33559
rect 8560 33525 8594 33559
rect 8696 33525 8730 33559
rect 8832 33525 8866 33559
rect 8968 33525 9002 33559
rect 9104 33525 9138 33559
rect 9240 33525 9274 33559
rect 7880 33389 7914 33423
rect 8016 33389 8050 33423
rect 8152 33389 8186 33423
rect 8288 33389 8322 33423
rect 8424 33389 8458 33423
rect 8560 33389 8594 33423
rect 8696 33389 8730 33423
rect 8832 33389 8866 33423
rect 8968 33389 9002 33423
rect 9104 33389 9138 33423
rect 9240 33389 9274 33423
rect 7880 33253 7914 33287
rect 8016 33253 8050 33287
rect 8152 33253 8186 33287
rect 8288 33253 8322 33287
rect 8424 33253 8458 33287
rect 8560 33253 8594 33287
rect 8696 33253 8730 33287
rect 8832 33253 8866 33287
rect 8968 33253 9002 33287
rect 9104 33253 9138 33287
rect 9240 33253 9274 33287
rect 7880 33117 7914 33151
rect 8016 33117 8050 33151
rect 8152 33117 8186 33151
rect 8288 33117 8322 33151
rect 8424 33117 8458 33151
rect 8560 33117 8594 33151
rect 8696 33117 8730 33151
rect 8832 33117 8866 33151
rect 8968 33117 9002 33151
rect 9104 33117 9138 33151
rect 9240 33117 9274 33151
rect 7880 32981 7914 33015
rect 8016 32981 8050 33015
rect 8152 32981 8186 33015
rect 8288 32981 8322 33015
rect 8424 32981 8458 33015
rect 8560 32981 8594 33015
rect 8696 32981 8730 33015
rect 8832 32981 8866 33015
rect 8968 32981 9002 33015
rect 9104 32981 9138 33015
rect 9240 32981 9274 33015
rect 7880 32845 7914 32879
rect 8016 32845 8050 32879
rect 8152 32845 8186 32879
rect 8288 32845 8322 32879
rect 8424 32845 8458 32879
rect 8560 32845 8594 32879
rect 8696 32845 8730 32879
rect 8832 32845 8866 32879
rect 8968 32845 9002 32879
rect 9104 32845 9138 32879
rect 9240 32845 9274 32879
rect 7880 32709 7914 32743
rect 8016 32709 8050 32743
rect 8152 32709 8186 32743
rect 8288 32709 8322 32743
rect 8424 32709 8458 32743
rect 8560 32709 8594 32743
rect 8696 32709 8730 32743
rect 8832 32709 8866 32743
rect 8968 32709 9002 32743
rect 9104 32709 9138 32743
rect 9240 32709 9274 32743
rect 7880 32573 7914 32607
rect 8016 32573 8050 32607
rect 8152 32573 8186 32607
rect 8288 32573 8322 32607
rect 8424 32573 8458 32607
rect 8560 32573 8594 32607
rect 8696 32573 8730 32607
rect 8832 32573 8866 32607
rect 8968 32573 9002 32607
rect 9104 32573 9138 32607
rect 9240 32573 9274 32607
rect 7880 32437 7914 32471
rect 8016 32437 8050 32471
rect 8152 32437 8186 32471
rect 8288 32437 8322 32471
rect 8424 32437 8458 32471
rect 8560 32437 8594 32471
rect 8696 32437 8730 32471
rect 8832 32437 8866 32471
rect 8968 32437 9002 32471
rect 9104 32437 9138 32471
rect 9240 32437 9274 32471
rect 7880 32301 7914 32335
rect 8016 32301 8050 32335
rect 8152 32301 8186 32335
rect 8288 32301 8322 32335
rect 8424 32301 8458 32335
rect 8560 32301 8594 32335
rect 8696 32301 8730 32335
rect 8832 32301 8866 32335
rect 8968 32301 9002 32335
rect 9104 32301 9138 32335
rect 9240 32301 9274 32335
rect 7880 32165 7914 32199
rect 8016 32165 8050 32199
rect 8152 32165 8186 32199
rect 8288 32165 8322 32199
rect 8424 32165 8458 32199
rect 8560 32165 8594 32199
rect 8696 32165 8730 32199
rect 8832 32165 8866 32199
rect 8968 32165 9002 32199
rect 9104 32165 9138 32199
rect 9240 32165 9274 32199
rect 7880 32029 7914 32063
rect 8016 32029 8050 32063
rect 8152 32029 8186 32063
rect 8288 32029 8322 32063
rect 8424 32029 8458 32063
rect 8560 32029 8594 32063
rect 8696 32029 8730 32063
rect 8832 32029 8866 32063
rect 8968 32029 9002 32063
rect 9104 32029 9138 32063
rect 9240 32029 9274 32063
rect 7880 31893 7914 31927
rect 8016 31893 8050 31927
rect 8152 31893 8186 31927
rect 8288 31893 8322 31927
rect 8424 31893 8458 31927
rect 8560 31893 8594 31927
rect 8696 31893 8730 31927
rect 8832 31893 8866 31927
rect 8968 31893 9002 31927
rect 9104 31893 9138 31927
rect 9240 31893 9274 31927
rect 7880 31757 7914 31791
rect 8016 31757 8050 31791
rect 8152 31757 8186 31791
rect 8288 31757 8322 31791
rect 8424 31757 8458 31791
rect 8560 31757 8594 31791
rect 8696 31757 8730 31791
rect 8832 31757 8866 31791
rect 8968 31757 9002 31791
rect 9104 31757 9138 31791
rect 9240 31757 9274 31791
rect 7880 31621 7914 31655
rect 8016 31621 8050 31655
rect 8152 31621 8186 31655
rect 8288 31621 8322 31655
rect 8424 31621 8458 31655
rect 8560 31621 8594 31655
rect 8696 31621 8730 31655
rect 8832 31621 8866 31655
rect 8968 31621 9002 31655
rect 9104 31621 9138 31655
rect 9240 31621 9274 31655
rect 7880 31485 7914 31519
rect 8016 31485 8050 31519
rect 8152 31485 8186 31519
rect 8288 31485 8322 31519
rect 8424 31485 8458 31519
rect 8560 31485 8594 31519
rect 8696 31485 8730 31519
rect 8832 31485 8866 31519
rect 8968 31485 9002 31519
rect 9104 31485 9138 31519
rect 9240 31485 9274 31519
rect 7880 31349 7914 31383
rect 8016 31349 8050 31383
rect 8152 31349 8186 31383
rect 8288 31349 8322 31383
rect 8424 31349 8458 31383
rect 8560 31349 8594 31383
rect 8696 31349 8730 31383
rect 8832 31349 8866 31383
rect 8968 31349 9002 31383
rect 9104 31349 9138 31383
rect 9240 31349 9274 31383
rect 7880 31213 7914 31247
rect 8016 31213 8050 31247
rect 8152 31213 8186 31247
rect 8288 31213 8322 31247
rect 8424 31213 8458 31247
rect 8560 31213 8594 31247
rect 8696 31213 8730 31247
rect 8832 31213 8866 31247
rect 8968 31213 9002 31247
rect 9104 31213 9138 31247
rect 9240 31213 9274 31247
rect 7880 31077 7914 31111
rect 8016 31077 8050 31111
rect 8152 31077 8186 31111
rect 8288 31077 8322 31111
rect 8424 31077 8458 31111
rect 8560 31077 8594 31111
rect 8696 31077 8730 31111
rect 8832 31077 8866 31111
rect 8968 31077 9002 31111
rect 9104 31077 9138 31111
rect 9240 31077 9274 31111
rect 7880 30941 7914 30975
rect 8016 30941 8050 30975
rect 8152 30941 8186 30975
rect 8288 30941 8322 30975
rect 8424 30941 8458 30975
rect 8560 30941 8594 30975
rect 8696 30941 8730 30975
rect 8832 30941 8866 30975
rect 8968 30941 9002 30975
rect 9104 30941 9138 30975
rect 9240 30941 9274 30975
rect 7880 30805 7914 30839
rect 8016 30805 8050 30839
rect 8152 30805 8186 30839
rect 8288 30805 8322 30839
rect 8424 30805 8458 30839
rect 8560 30805 8594 30839
rect 8696 30805 8730 30839
rect 8832 30805 8866 30839
rect 8968 30805 9002 30839
rect 9104 30805 9138 30839
rect 9240 30805 9274 30839
rect 7880 30669 7914 30703
rect 8016 30669 8050 30703
rect 8152 30669 8186 30703
rect 8288 30669 8322 30703
rect 8424 30669 8458 30703
rect 8560 30669 8594 30703
rect 8696 30669 8730 30703
rect 8832 30669 8866 30703
rect 8968 30669 9002 30703
rect 9104 30669 9138 30703
rect 9240 30669 9274 30703
rect 7880 30533 7914 30567
rect 8016 30533 8050 30567
rect 8152 30533 8186 30567
rect 8288 30533 8322 30567
rect 8424 30533 8458 30567
rect 8560 30533 8594 30567
rect 8696 30533 8730 30567
rect 8832 30533 8866 30567
rect 8968 30533 9002 30567
rect 9104 30533 9138 30567
rect 9240 30533 9274 30567
rect 7880 30397 7914 30431
rect 8016 30397 8050 30431
rect 8152 30397 8186 30431
rect 8288 30397 8322 30431
rect 8424 30397 8458 30431
rect 8560 30397 8594 30431
rect 8696 30397 8730 30431
rect 8832 30397 8866 30431
rect 8968 30397 9002 30431
rect 9104 30397 9138 30431
rect 9240 30397 9274 30431
rect 7880 30261 7914 30295
rect 8016 30261 8050 30295
rect 8152 30261 8186 30295
rect 8288 30261 8322 30295
rect 8424 30261 8458 30295
rect 8560 30261 8594 30295
rect 8696 30261 8730 30295
rect 8832 30261 8866 30295
rect 8968 30261 9002 30295
rect 9104 30261 9138 30295
rect 9240 30261 9274 30295
rect 7880 30125 7914 30159
rect 8016 30125 8050 30159
rect 8152 30125 8186 30159
rect 8288 30125 8322 30159
rect 8424 30125 8458 30159
rect 8560 30125 8594 30159
rect 8696 30125 8730 30159
rect 8832 30125 8866 30159
rect 8968 30125 9002 30159
rect 9104 30125 9138 30159
rect 9240 30125 9274 30159
rect 7880 29989 7914 30023
rect 8016 29989 8050 30023
rect 8152 29989 8186 30023
rect 8288 29989 8322 30023
rect 8424 29989 8458 30023
rect 8560 29989 8594 30023
rect 8696 29989 8730 30023
rect 8832 29989 8866 30023
rect 8968 29989 9002 30023
rect 9104 29989 9138 30023
rect 9240 29989 9274 30023
rect 7880 29853 7914 29887
rect 8016 29853 8050 29887
rect 8152 29853 8186 29887
rect 8288 29853 8322 29887
rect 8424 29853 8458 29887
rect 8560 29853 8594 29887
rect 8696 29853 8730 29887
rect 8832 29853 8866 29887
rect 8968 29853 9002 29887
rect 9104 29853 9138 29887
rect 9240 29853 9274 29887
rect 7880 29717 7914 29751
rect 8016 29717 8050 29751
rect 8152 29717 8186 29751
rect 8288 29717 8322 29751
rect 8424 29717 8458 29751
rect 8560 29717 8594 29751
rect 8696 29717 8730 29751
rect 8832 29717 8866 29751
rect 8968 29717 9002 29751
rect 9104 29717 9138 29751
rect 9240 29717 9274 29751
rect 7880 29581 7914 29615
rect 8016 29581 8050 29615
rect 8152 29581 8186 29615
rect 8288 29581 8322 29615
rect 8424 29581 8458 29615
rect 8560 29581 8594 29615
rect 8696 29581 8730 29615
rect 8832 29581 8866 29615
rect 8968 29581 9002 29615
rect 9104 29581 9138 29615
rect 9240 29581 9274 29615
rect 7880 29445 7914 29479
rect 8016 29445 8050 29479
rect 8152 29445 8186 29479
rect 8288 29445 8322 29479
rect 8424 29445 8458 29479
rect 8560 29445 8594 29479
rect 8696 29445 8730 29479
rect 8832 29445 8866 29479
rect 8968 29445 9002 29479
rect 9104 29445 9138 29479
rect 9240 29445 9274 29479
rect 7880 29309 7914 29343
rect 8016 29309 8050 29343
rect 8152 29309 8186 29343
rect 8288 29309 8322 29343
rect 8424 29309 8458 29343
rect 8560 29309 8594 29343
rect 8696 29309 8730 29343
rect 8832 29309 8866 29343
rect 8968 29309 9002 29343
rect 9104 29309 9138 29343
rect 9240 29309 9274 29343
rect 7880 29173 7914 29207
rect 8016 29173 8050 29207
rect 8152 29173 8186 29207
rect 8288 29173 8322 29207
rect 8424 29173 8458 29207
rect 8560 29173 8594 29207
rect 8696 29173 8730 29207
rect 8832 29173 8866 29207
rect 8968 29173 9002 29207
rect 9104 29173 9138 29207
rect 9240 29173 9274 29207
rect 7880 29037 7914 29071
rect 8016 29037 8050 29071
rect 8152 29037 8186 29071
rect 8288 29037 8322 29071
rect 8424 29037 8458 29071
rect 8560 29037 8594 29071
rect 8696 29037 8730 29071
rect 8832 29037 8866 29071
rect 8968 29037 9002 29071
rect 9104 29037 9138 29071
rect 9240 29037 9274 29071
rect 7880 28901 7914 28935
rect 8016 28901 8050 28935
rect 8152 28901 8186 28935
rect 8288 28901 8322 28935
rect 8424 28901 8458 28935
rect 8560 28901 8594 28935
rect 8696 28901 8730 28935
rect 8832 28901 8866 28935
rect 8968 28901 9002 28935
rect 9104 28901 9138 28935
rect 9240 28901 9274 28935
rect 7880 28765 7914 28799
rect 8016 28765 8050 28799
rect 8152 28765 8186 28799
rect 8288 28765 8322 28799
rect 8424 28765 8458 28799
rect 8560 28765 8594 28799
rect 8696 28765 8730 28799
rect 8832 28765 8866 28799
rect 8968 28765 9002 28799
rect 9104 28765 9138 28799
rect 9240 28765 9274 28799
rect 7880 28629 7914 28663
rect 8016 28629 8050 28663
rect 8152 28629 8186 28663
rect 8288 28629 8322 28663
rect 8424 28629 8458 28663
rect 8560 28629 8594 28663
rect 8696 28629 8730 28663
rect 8832 28629 8866 28663
rect 8968 28629 9002 28663
rect 9104 28629 9138 28663
rect 9240 28629 9274 28663
rect 7880 28493 7914 28527
rect 8016 28493 8050 28527
rect 8152 28493 8186 28527
rect 8288 28493 8322 28527
rect 8424 28493 8458 28527
rect 8560 28493 8594 28527
rect 8696 28493 8730 28527
rect 8832 28493 8866 28527
rect 8968 28493 9002 28527
rect 9104 28493 9138 28527
rect 9240 28493 9274 28527
rect 7880 28357 7914 28391
rect 8016 28357 8050 28391
rect 8152 28357 8186 28391
rect 8288 28357 8322 28391
rect 8424 28357 8458 28391
rect 8560 28357 8594 28391
rect 8696 28357 8730 28391
rect 8832 28357 8866 28391
rect 8968 28357 9002 28391
rect 9104 28357 9138 28391
rect 9240 28357 9274 28391
rect 7880 28221 7914 28255
rect 8016 28221 8050 28255
rect 8152 28221 8186 28255
rect 8288 28221 8322 28255
rect 8424 28221 8458 28255
rect 8560 28221 8594 28255
rect 8696 28221 8730 28255
rect 8832 28221 8866 28255
rect 8968 28221 9002 28255
rect 9104 28221 9138 28255
rect 9240 28221 9274 28255
rect 7880 28085 7914 28119
rect 8016 28085 8050 28119
rect 8152 28085 8186 28119
rect 8288 28085 8322 28119
rect 8424 28085 8458 28119
rect 8560 28085 8594 28119
rect 8696 28085 8730 28119
rect 8832 28085 8866 28119
rect 8968 28085 9002 28119
rect 9104 28085 9138 28119
rect 9240 28085 9274 28119
rect 7880 27949 7914 27983
rect 8016 27949 8050 27983
rect 8152 27949 8186 27983
rect 8288 27949 8322 27983
rect 8424 27949 8458 27983
rect 8560 27949 8594 27983
rect 8696 27949 8730 27983
rect 8832 27949 8866 27983
rect 8968 27949 9002 27983
rect 9104 27949 9138 27983
rect 9240 27949 9274 27983
rect 7880 27813 7914 27847
rect 8016 27813 8050 27847
rect 8152 27813 8186 27847
rect 8288 27813 8322 27847
rect 8424 27813 8458 27847
rect 8560 27813 8594 27847
rect 8696 27813 8730 27847
rect 8832 27813 8866 27847
rect 8968 27813 9002 27847
rect 9104 27813 9138 27847
rect 9240 27813 9274 27847
rect 7880 27677 7914 27711
rect 8016 27677 8050 27711
rect 8152 27677 8186 27711
rect 8288 27677 8322 27711
rect 8424 27677 8458 27711
rect 8560 27677 8594 27711
rect 8696 27677 8730 27711
rect 8832 27677 8866 27711
rect 8968 27677 9002 27711
rect 9104 27677 9138 27711
rect 9240 27677 9274 27711
rect 7880 27541 7914 27575
rect 8016 27541 8050 27575
rect 8152 27541 8186 27575
rect 8288 27541 8322 27575
rect 8424 27541 8458 27575
rect 8560 27541 8594 27575
rect 8696 27541 8730 27575
rect 8832 27541 8866 27575
rect 8968 27541 9002 27575
rect 9104 27541 9138 27575
rect 9240 27541 9274 27575
rect 7880 27405 7914 27439
rect 8016 27405 8050 27439
rect 8152 27405 8186 27439
rect 8288 27405 8322 27439
rect 8424 27405 8458 27439
rect 8560 27405 8594 27439
rect 8696 27405 8730 27439
rect 8832 27405 8866 27439
rect 8968 27405 9002 27439
rect 9104 27405 9138 27439
rect 9240 27405 9274 27439
rect 7880 27269 7914 27303
rect 8016 27269 8050 27303
rect 8152 27269 8186 27303
rect 8288 27269 8322 27303
rect 8424 27269 8458 27303
rect 8560 27269 8594 27303
rect 8696 27269 8730 27303
rect 8832 27269 8866 27303
rect 8968 27269 9002 27303
rect 9104 27269 9138 27303
rect 9240 27269 9274 27303
rect 7880 27133 7914 27167
rect 8016 27133 8050 27167
rect 8152 27133 8186 27167
rect 8288 27133 8322 27167
rect 8424 27133 8458 27167
rect 8560 27133 8594 27167
rect 8696 27133 8730 27167
rect 8832 27133 8866 27167
rect 8968 27133 9002 27167
rect 9104 27133 9138 27167
rect 9240 27133 9274 27167
rect 7880 26997 7914 27031
rect 8016 26997 8050 27031
rect 8152 26997 8186 27031
rect 8288 26997 8322 27031
rect 8424 26997 8458 27031
rect 8560 26997 8594 27031
rect 8696 26997 8730 27031
rect 8832 26997 8866 27031
rect 8968 26997 9002 27031
rect 9104 26997 9138 27031
rect 9240 26997 9274 27031
rect 7880 26861 7914 26895
rect 8016 26861 8050 26895
rect 8152 26861 8186 26895
rect 8288 26861 8322 26895
rect 8424 26861 8458 26895
rect 8560 26861 8594 26895
rect 8696 26861 8730 26895
rect 8832 26861 8866 26895
rect 8968 26861 9002 26895
rect 9104 26861 9138 26895
rect 9240 26861 9274 26895
rect 7880 26725 7914 26759
rect 8016 26725 8050 26759
rect 8152 26725 8186 26759
rect 8288 26725 8322 26759
rect 8424 26725 8458 26759
rect 8560 26725 8594 26759
rect 8696 26725 8730 26759
rect 8832 26725 8866 26759
rect 8968 26725 9002 26759
rect 9104 26725 9138 26759
rect 9240 26725 9274 26759
rect 7880 26589 7914 26623
rect 8016 26589 8050 26623
rect 8152 26589 8186 26623
rect 8288 26589 8322 26623
rect 8424 26589 8458 26623
rect 8560 26589 8594 26623
rect 8696 26589 8730 26623
rect 8832 26589 8866 26623
rect 8968 26589 9002 26623
rect 9104 26589 9138 26623
rect 9240 26589 9274 26623
rect 7880 26453 7914 26487
rect 8016 26453 8050 26487
rect 8152 26453 8186 26487
rect 8288 26453 8322 26487
rect 8424 26453 8458 26487
rect 8560 26453 8594 26487
rect 8696 26453 8730 26487
rect 8832 26453 8866 26487
rect 8968 26453 9002 26487
rect 9104 26453 9138 26487
rect 9240 26453 9274 26487
rect 7880 26317 7914 26351
rect 8016 26317 8050 26351
rect 8152 26317 8186 26351
rect 8288 26317 8322 26351
rect 8424 26317 8458 26351
rect 8560 26317 8594 26351
rect 8696 26317 8730 26351
rect 8832 26317 8866 26351
rect 8968 26317 9002 26351
rect 9104 26317 9138 26351
rect 9240 26317 9274 26351
rect 7880 26181 7914 26215
rect 8016 26181 8050 26215
rect 8152 26181 8186 26215
rect 8288 26181 8322 26215
rect 8424 26181 8458 26215
rect 8560 26181 8594 26215
rect 8696 26181 8730 26215
rect 8832 26181 8866 26215
rect 8968 26181 9002 26215
rect 9104 26181 9138 26215
rect 9240 26181 9274 26215
rect 7880 26045 7914 26079
rect 8016 26045 8050 26079
rect 8152 26045 8186 26079
rect 8288 26045 8322 26079
rect 8424 26045 8458 26079
rect 8560 26045 8594 26079
rect 8696 26045 8730 26079
rect 8832 26045 8866 26079
rect 8968 26045 9002 26079
rect 9104 26045 9138 26079
rect 9240 26045 9274 26079
rect 7880 25909 7914 25943
rect 8016 25909 8050 25943
rect 8152 25909 8186 25943
rect 8288 25909 8322 25943
rect 8424 25909 8458 25943
rect 8560 25909 8594 25943
rect 8696 25909 8730 25943
rect 8832 25909 8866 25943
rect 8968 25909 9002 25943
rect 9104 25909 9138 25943
rect 9240 25909 9274 25943
rect 7880 25773 7914 25807
rect 8016 25773 8050 25807
rect 8152 25773 8186 25807
rect 8288 25773 8322 25807
rect 8424 25773 8458 25807
rect 8560 25773 8594 25807
rect 8696 25773 8730 25807
rect 8832 25773 8866 25807
rect 8968 25773 9002 25807
rect 9104 25773 9138 25807
rect 9240 25773 9274 25807
rect 7880 25637 7914 25671
rect 8016 25637 8050 25671
rect 8152 25637 8186 25671
rect 8288 25637 8322 25671
rect 8424 25637 8458 25671
rect 8560 25637 8594 25671
rect 8696 25637 8730 25671
rect 8832 25637 8866 25671
rect 8968 25637 9002 25671
rect 9104 25637 9138 25671
rect 9240 25637 9274 25671
rect 7880 25501 7914 25535
rect 8016 25501 8050 25535
rect 8152 25501 8186 25535
rect 8288 25501 8322 25535
rect 8424 25501 8458 25535
rect 8560 25501 8594 25535
rect 8696 25501 8730 25535
rect 8832 25501 8866 25535
rect 8968 25501 9002 25535
rect 9104 25501 9138 25535
rect 9240 25501 9274 25535
rect 7880 25365 7914 25399
rect 8016 25365 8050 25399
rect 8152 25365 8186 25399
rect 8288 25365 8322 25399
rect 8424 25365 8458 25399
rect 8560 25365 8594 25399
rect 8696 25365 8730 25399
rect 8832 25365 8866 25399
rect 8968 25365 9002 25399
rect 9104 25365 9138 25399
rect 9240 25365 9274 25399
rect 7880 25229 7914 25263
rect 8016 25229 8050 25263
rect 8152 25229 8186 25263
rect 8288 25229 8322 25263
rect 8424 25229 8458 25263
rect 8560 25229 8594 25263
rect 8696 25229 8730 25263
rect 8832 25229 8866 25263
rect 8968 25229 9002 25263
rect 9104 25229 9138 25263
rect 9240 25229 9274 25263
rect 7880 25093 7914 25127
rect 8016 25093 8050 25127
rect 8152 25093 8186 25127
rect 8288 25093 8322 25127
rect 8424 25093 8458 25127
rect 8560 25093 8594 25127
rect 8696 25093 8730 25127
rect 8832 25093 8866 25127
rect 8968 25093 9002 25127
rect 9104 25093 9138 25127
rect 9240 25093 9274 25127
rect 7880 24957 7914 24991
rect 8016 24957 8050 24991
rect 8152 24957 8186 24991
rect 8288 24957 8322 24991
rect 8424 24957 8458 24991
rect 8560 24957 8594 24991
rect 8696 24957 8730 24991
rect 8832 24957 8866 24991
rect 8968 24957 9002 24991
rect 9104 24957 9138 24991
rect 9240 24957 9274 24991
rect 7880 24821 7914 24855
rect 8016 24821 8050 24855
rect 8152 24821 8186 24855
rect 8288 24821 8322 24855
rect 8424 24821 8458 24855
rect 8560 24821 8594 24855
rect 8696 24821 8730 24855
rect 8832 24821 8866 24855
rect 8968 24821 9002 24855
rect 9104 24821 9138 24855
rect 9240 24821 9274 24855
rect 7880 24685 7914 24719
rect 8016 24685 8050 24719
rect 8152 24685 8186 24719
rect 8288 24685 8322 24719
rect 8424 24685 8458 24719
rect 8560 24685 8594 24719
rect 8696 24685 8730 24719
rect 8832 24685 8866 24719
rect 8968 24685 9002 24719
rect 9104 24685 9138 24719
rect 9240 24685 9274 24719
rect 7880 24549 7914 24583
rect 8016 24549 8050 24583
rect 8152 24549 8186 24583
rect 8288 24549 8322 24583
rect 8424 24549 8458 24583
rect 8560 24549 8594 24583
rect 8696 24549 8730 24583
rect 8832 24549 8866 24583
rect 8968 24549 9002 24583
rect 9104 24549 9138 24583
rect 9240 24549 9274 24583
rect 7880 24413 7914 24447
rect 8016 24413 8050 24447
rect 8152 24413 8186 24447
rect 8288 24413 8322 24447
rect 8424 24413 8458 24447
rect 8560 24413 8594 24447
rect 8696 24413 8730 24447
rect 8832 24413 8866 24447
rect 8968 24413 9002 24447
rect 9104 24413 9138 24447
rect 9240 24413 9274 24447
rect 7880 24277 7914 24311
rect 8016 24277 8050 24311
rect 8152 24277 8186 24311
rect 8288 24277 8322 24311
rect 8424 24277 8458 24311
rect 8560 24277 8594 24311
rect 8696 24277 8730 24311
rect 8832 24277 8866 24311
rect 8968 24277 9002 24311
rect 9104 24277 9138 24311
rect 9240 24277 9274 24311
rect 7880 24141 7914 24175
rect 8016 24141 8050 24175
rect 8152 24141 8186 24175
rect 8288 24141 8322 24175
rect 8424 24141 8458 24175
rect 8560 24141 8594 24175
rect 8696 24141 8730 24175
rect 8832 24141 8866 24175
rect 8968 24141 9002 24175
rect 9104 24141 9138 24175
rect 9240 24141 9274 24175
rect 7880 24005 7914 24039
rect 8016 24005 8050 24039
rect 8152 24005 8186 24039
rect 8288 24005 8322 24039
rect 8424 24005 8458 24039
rect 8560 24005 8594 24039
rect 8696 24005 8730 24039
rect 8832 24005 8866 24039
rect 8968 24005 9002 24039
rect 9104 24005 9138 24039
rect 9240 24005 9274 24039
rect 7880 23869 7914 23903
rect 8016 23869 8050 23903
rect 8152 23869 8186 23903
rect 8288 23869 8322 23903
rect 8424 23869 8458 23903
rect 8560 23869 8594 23903
rect 8696 23869 8730 23903
rect 8832 23869 8866 23903
rect 8968 23869 9002 23903
rect 9104 23869 9138 23903
rect 9240 23869 9274 23903
rect 7880 23733 7914 23767
rect 8016 23733 8050 23767
rect 8152 23733 8186 23767
rect 8288 23733 8322 23767
rect 8424 23733 8458 23767
rect 8560 23733 8594 23767
rect 8696 23733 8730 23767
rect 8832 23733 8866 23767
rect 8968 23733 9002 23767
rect 9104 23733 9138 23767
rect 9240 23733 9274 23767
rect 7880 23597 7914 23631
rect 8016 23597 8050 23631
rect 8152 23597 8186 23631
rect 8288 23597 8322 23631
rect 8424 23597 8458 23631
rect 8560 23597 8594 23631
rect 8696 23597 8730 23631
rect 8832 23597 8866 23631
rect 8968 23597 9002 23631
rect 9104 23597 9138 23631
rect 9240 23597 9274 23631
rect 7880 23461 7914 23495
rect 8016 23461 8050 23495
rect 8152 23461 8186 23495
rect 8288 23461 8322 23495
rect 8424 23461 8458 23495
rect 8560 23461 8594 23495
rect 8696 23461 8730 23495
rect 8832 23461 8866 23495
rect 8968 23461 9002 23495
rect 9104 23461 9138 23495
rect 9240 23461 9274 23495
rect 7880 23325 7914 23359
rect 8016 23325 8050 23359
rect 8152 23325 8186 23359
rect 8288 23325 8322 23359
rect 8424 23325 8458 23359
rect 8560 23325 8594 23359
rect 8696 23325 8730 23359
rect 8832 23325 8866 23359
rect 8968 23325 9002 23359
rect 9104 23325 9138 23359
rect 9240 23325 9274 23359
rect 7880 23189 7914 23223
rect 8016 23189 8050 23223
rect 8152 23189 8186 23223
rect 8288 23189 8322 23223
rect 8424 23189 8458 23223
rect 8560 23189 8594 23223
rect 8696 23189 8730 23223
rect 8832 23189 8866 23223
rect 8968 23189 9002 23223
rect 9104 23189 9138 23223
rect 9240 23189 9274 23223
rect 7880 23053 7914 23087
rect 8016 23053 8050 23087
rect 8152 23053 8186 23087
rect 8288 23053 8322 23087
rect 8424 23053 8458 23087
rect 8560 23053 8594 23087
rect 8696 23053 8730 23087
rect 8832 23053 8866 23087
rect 8968 23053 9002 23087
rect 9104 23053 9138 23087
rect 9240 23053 9274 23087
rect 7880 22917 7914 22951
rect 8016 22917 8050 22951
rect 8152 22917 8186 22951
rect 8288 22917 8322 22951
rect 8424 22917 8458 22951
rect 8560 22917 8594 22951
rect 8696 22917 8730 22951
rect 8832 22917 8866 22951
rect 8968 22917 9002 22951
rect 9104 22917 9138 22951
rect 9240 22917 9274 22951
rect 7880 22781 7914 22815
rect 8016 22781 8050 22815
rect 8152 22781 8186 22815
rect 8288 22781 8322 22815
rect 8424 22781 8458 22815
rect 8560 22781 8594 22815
rect 8696 22781 8730 22815
rect 8832 22781 8866 22815
rect 8968 22781 9002 22815
rect 9104 22781 9138 22815
rect 9240 22781 9274 22815
rect 7880 22645 7914 22679
rect 8016 22645 8050 22679
rect 8152 22645 8186 22679
rect 8288 22645 8322 22679
rect 8424 22645 8458 22679
rect 8560 22645 8594 22679
rect 8696 22645 8730 22679
rect 8832 22645 8866 22679
rect 8968 22645 9002 22679
rect 9104 22645 9138 22679
rect 9240 22645 9274 22679
rect 7880 22509 7914 22543
rect 8016 22509 8050 22543
rect 8152 22509 8186 22543
rect 8288 22509 8322 22543
rect 8424 22509 8458 22543
rect 8560 22509 8594 22543
rect 8696 22509 8730 22543
rect 8832 22509 8866 22543
rect 8968 22509 9002 22543
rect 9104 22509 9138 22543
rect 9240 22509 9274 22543
rect 7880 22373 7914 22407
rect 8016 22373 8050 22407
rect 8152 22373 8186 22407
rect 8288 22373 8322 22407
rect 8424 22373 8458 22407
rect 8560 22373 8594 22407
rect 8696 22373 8730 22407
rect 8832 22373 8866 22407
rect 8968 22373 9002 22407
rect 9104 22373 9138 22407
rect 9240 22373 9274 22407
rect 7880 22237 7914 22271
rect 8016 22237 8050 22271
rect 8152 22237 8186 22271
rect 8288 22237 8322 22271
rect 8424 22237 8458 22271
rect 8560 22237 8594 22271
rect 8696 22237 8730 22271
rect 8832 22237 8866 22271
rect 8968 22237 9002 22271
rect 9104 22237 9138 22271
rect 9240 22237 9274 22271
rect 7880 22101 7914 22135
rect 8016 22101 8050 22135
rect 8152 22101 8186 22135
rect 8288 22101 8322 22135
rect 8424 22101 8458 22135
rect 8560 22101 8594 22135
rect 8696 22101 8730 22135
rect 8832 22101 8866 22135
rect 8968 22101 9002 22135
rect 9104 22101 9138 22135
rect 9240 22101 9274 22135
rect 7880 21965 7914 21999
rect 8016 21965 8050 21999
rect 8152 21965 8186 21999
rect 8288 21965 8322 21999
rect 8424 21965 8458 21999
rect 8560 21965 8594 21999
rect 8696 21965 8730 21999
rect 8832 21965 8866 21999
rect 8968 21965 9002 21999
rect 9104 21965 9138 21999
rect 9240 21965 9274 21999
rect 7880 21829 7914 21863
rect 8016 21829 8050 21863
rect 8152 21829 8186 21863
rect 8288 21829 8322 21863
rect 8424 21829 8458 21863
rect 8560 21829 8594 21863
rect 8696 21829 8730 21863
rect 8832 21829 8866 21863
rect 8968 21829 9002 21863
rect 9104 21829 9138 21863
rect 9240 21829 9274 21863
rect 7880 21693 7914 21727
rect 8016 21693 8050 21727
rect 8152 21693 8186 21727
rect 8288 21693 8322 21727
rect 8424 21693 8458 21727
rect 8560 21693 8594 21727
rect 8696 21693 8730 21727
rect 8832 21693 8866 21727
rect 8968 21693 9002 21727
rect 9104 21693 9138 21727
rect 9240 21693 9274 21727
rect 7880 21557 7914 21591
rect 8016 21557 8050 21591
rect 8152 21557 8186 21591
rect 8288 21557 8322 21591
rect 8424 21557 8458 21591
rect 8560 21557 8594 21591
rect 8696 21557 8730 21591
rect 8832 21557 8866 21591
rect 8968 21557 9002 21591
rect 9104 21557 9138 21591
rect 9240 21557 9274 21591
rect 7880 21421 7914 21455
rect 8016 21421 8050 21455
rect 8152 21421 8186 21455
rect 8288 21421 8322 21455
rect 8424 21421 8458 21455
rect 8560 21421 8594 21455
rect 8696 21421 8730 21455
rect 8832 21421 8866 21455
rect 8968 21421 9002 21455
rect 9104 21421 9138 21455
rect 9240 21421 9274 21455
rect 7880 21285 7914 21319
rect 8016 21285 8050 21319
rect 8152 21285 8186 21319
rect 8288 21285 8322 21319
rect 8424 21285 8458 21319
rect 8560 21285 8594 21319
rect 8696 21285 8730 21319
rect 8832 21285 8866 21319
rect 8968 21285 9002 21319
rect 9104 21285 9138 21319
rect 9240 21285 9274 21319
rect 7880 21149 7914 21183
rect 8016 21149 8050 21183
rect 8152 21149 8186 21183
rect 8288 21149 8322 21183
rect 8424 21149 8458 21183
rect 8560 21149 8594 21183
rect 8696 21149 8730 21183
rect 8832 21149 8866 21183
rect 8968 21149 9002 21183
rect 9104 21149 9138 21183
rect 9240 21149 9274 21183
rect 7880 21013 7914 21047
rect 8016 21013 8050 21047
rect 8152 21013 8186 21047
rect 8288 21013 8322 21047
rect 8424 21013 8458 21047
rect 8560 21013 8594 21047
rect 8696 21013 8730 21047
rect 8832 21013 8866 21047
rect 8968 21013 9002 21047
rect 9104 21013 9138 21047
rect 9240 21013 9274 21047
rect 7880 20877 7914 20911
rect 8016 20877 8050 20911
rect 8152 20877 8186 20911
rect 8288 20877 8322 20911
rect 8424 20877 8458 20911
rect 8560 20877 8594 20911
rect 8696 20877 8730 20911
rect 8832 20877 8866 20911
rect 8968 20877 9002 20911
rect 9104 20877 9138 20911
rect 9240 20877 9274 20911
rect 7880 20741 7914 20775
rect 8016 20741 8050 20775
rect 8152 20741 8186 20775
rect 8288 20741 8322 20775
rect 8424 20741 8458 20775
rect 8560 20741 8594 20775
rect 8696 20741 8730 20775
rect 8832 20741 8866 20775
rect 8968 20741 9002 20775
rect 9104 20741 9138 20775
rect 9240 20741 9274 20775
rect 7880 20605 7914 20639
rect 8016 20605 8050 20639
rect 8152 20605 8186 20639
rect 8288 20605 8322 20639
rect 8424 20605 8458 20639
rect 8560 20605 8594 20639
rect 8696 20605 8730 20639
rect 8832 20605 8866 20639
rect 8968 20605 9002 20639
rect 9104 20605 9138 20639
rect 9240 20605 9274 20639
rect 7880 20469 7914 20503
rect 8016 20469 8050 20503
rect 8152 20469 8186 20503
rect 8288 20469 8322 20503
rect 8424 20469 8458 20503
rect 8560 20469 8594 20503
rect 8696 20469 8730 20503
rect 8832 20469 8866 20503
rect 8968 20469 9002 20503
rect 9104 20469 9138 20503
rect 9240 20469 9274 20503
rect 7880 20333 7914 20367
rect 8016 20333 8050 20367
rect 8152 20333 8186 20367
rect 8288 20333 8322 20367
rect 8424 20333 8458 20367
rect 8560 20333 8594 20367
rect 8696 20333 8730 20367
rect 8832 20333 8866 20367
rect 8968 20333 9002 20367
rect 9104 20333 9138 20367
rect 9240 20333 9274 20367
rect 7880 20197 7914 20231
rect 8016 20197 8050 20231
rect 8152 20197 8186 20231
rect 8288 20197 8322 20231
rect 8424 20197 8458 20231
rect 8560 20197 8594 20231
rect 8696 20197 8730 20231
rect 8832 20197 8866 20231
rect 8968 20197 9002 20231
rect 9104 20197 9138 20231
rect 9240 20197 9274 20231
rect 7880 20061 7914 20095
rect 8016 20061 8050 20095
rect 8152 20061 8186 20095
rect 8288 20061 8322 20095
rect 8424 20061 8458 20095
rect 8560 20061 8594 20095
rect 8696 20061 8730 20095
rect 8832 20061 8866 20095
rect 8968 20061 9002 20095
rect 9104 20061 9138 20095
rect 9240 20061 9274 20095
rect 7880 19925 7914 19959
rect 8016 19925 8050 19959
rect 8152 19925 8186 19959
rect 8288 19925 8322 19959
rect 8424 19925 8458 19959
rect 8560 19925 8594 19959
rect 8696 19925 8730 19959
rect 8832 19925 8866 19959
rect 8968 19925 9002 19959
rect 9104 19925 9138 19959
rect 9240 19925 9274 19959
rect 7880 19789 7914 19823
rect 8016 19789 8050 19823
rect 8152 19789 8186 19823
rect 8288 19789 8322 19823
rect 8424 19789 8458 19823
rect 8560 19789 8594 19823
rect 8696 19789 8730 19823
rect 8832 19789 8866 19823
rect 8968 19789 9002 19823
rect 9104 19789 9138 19823
rect 9240 19789 9274 19823
rect 7880 19653 7914 19687
rect 8016 19653 8050 19687
rect 8152 19653 8186 19687
rect 8288 19653 8322 19687
rect 8424 19653 8458 19687
rect 8560 19653 8594 19687
rect 8696 19653 8730 19687
rect 8832 19653 8866 19687
rect 8968 19653 9002 19687
rect 9104 19653 9138 19687
rect 9240 19653 9274 19687
rect 7880 19517 7914 19551
rect 8016 19517 8050 19551
rect 8152 19517 8186 19551
rect 8288 19517 8322 19551
rect 8424 19517 8458 19551
rect 8560 19517 8594 19551
rect 8696 19517 8730 19551
rect 8832 19517 8866 19551
rect 8968 19517 9002 19551
rect 9104 19517 9138 19551
rect 9240 19517 9274 19551
rect 7880 19381 7914 19415
rect 8016 19381 8050 19415
rect 8152 19381 8186 19415
rect 8288 19381 8322 19415
rect 8424 19381 8458 19415
rect 8560 19381 8594 19415
rect 8696 19381 8730 19415
rect 8832 19381 8866 19415
rect 8968 19381 9002 19415
rect 9104 19381 9138 19415
rect 9240 19381 9274 19415
rect 7880 19245 7914 19279
rect 8016 19245 8050 19279
rect 8152 19245 8186 19279
rect 8288 19245 8322 19279
rect 8424 19245 8458 19279
rect 8560 19245 8594 19279
rect 8696 19245 8730 19279
rect 8832 19245 8866 19279
rect 8968 19245 9002 19279
rect 9104 19245 9138 19279
rect 9240 19245 9274 19279
rect 7880 19109 7914 19143
rect 8016 19109 8050 19143
rect 8152 19109 8186 19143
rect 8288 19109 8322 19143
rect 8424 19109 8458 19143
rect 8560 19109 8594 19143
rect 8696 19109 8730 19143
rect 8832 19109 8866 19143
rect 8968 19109 9002 19143
rect 9104 19109 9138 19143
rect 9240 19109 9274 19143
rect 7880 18973 7914 19007
rect 8016 18973 8050 19007
rect 8152 18973 8186 19007
rect 8288 18973 8322 19007
rect 8424 18973 8458 19007
rect 8560 18973 8594 19007
rect 8696 18973 8730 19007
rect 8832 18973 8866 19007
rect 8968 18973 9002 19007
rect 9104 18973 9138 19007
rect 9240 18973 9274 19007
rect 7880 18837 7914 18871
rect 8016 18837 8050 18871
rect 8152 18837 8186 18871
rect 8288 18837 8322 18871
rect 8424 18837 8458 18871
rect 8560 18837 8594 18871
rect 8696 18837 8730 18871
rect 8832 18837 8866 18871
rect 8968 18837 9002 18871
rect 9104 18837 9138 18871
rect 9240 18837 9274 18871
rect 7880 18701 7914 18735
rect 8016 18701 8050 18735
rect 8152 18701 8186 18735
rect 8288 18701 8322 18735
rect 8424 18701 8458 18735
rect 8560 18701 8594 18735
rect 8696 18701 8730 18735
rect 8832 18701 8866 18735
rect 8968 18701 9002 18735
rect 9104 18701 9138 18735
rect 9240 18701 9274 18735
rect 7880 18565 7914 18599
rect 8016 18565 8050 18599
rect 8152 18565 8186 18599
rect 8288 18565 8322 18599
rect 8424 18565 8458 18599
rect 8560 18565 8594 18599
rect 8696 18565 8730 18599
rect 8832 18565 8866 18599
rect 8968 18565 9002 18599
rect 9104 18565 9138 18599
rect 9240 18565 9274 18599
rect 7880 18429 7914 18463
rect 8016 18429 8050 18463
rect 8152 18429 8186 18463
rect 8288 18429 8322 18463
rect 8424 18429 8458 18463
rect 8560 18429 8594 18463
rect 8696 18429 8730 18463
rect 8832 18429 8866 18463
rect 8968 18429 9002 18463
rect 9104 18429 9138 18463
rect 9240 18429 9274 18463
rect 7880 18293 7914 18327
rect 8016 18293 8050 18327
rect 8152 18293 8186 18327
rect 8288 18293 8322 18327
rect 8424 18293 8458 18327
rect 8560 18293 8594 18327
rect 8696 18293 8730 18327
rect 8832 18293 8866 18327
rect 8968 18293 9002 18327
rect 9104 18293 9138 18327
rect 9240 18293 9274 18327
rect 7880 18157 7914 18191
rect 8016 18157 8050 18191
rect 8152 18157 8186 18191
rect 8288 18157 8322 18191
rect 8424 18157 8458 18191
rect 8560 18157 8594 18191
rect 8696 18157 8730 18191
rect 8832 18157 8866 18191
rect 8968 18157 9002 18191
rect 9104 18157 9138 18191
rect 9240 18157 9274 18191
rect 7880 18021 7914 18055
rect 8016 18021 8050 18055
rect 8152 18021 8186 18055
rect 8288 18021 8322 18055
rect 8424 18021 8458 18055
rect 8560 18021 8594 18055
rect 8696 18021 8730 18055
rect 8832 18021 8866 18055
rect 8968 18021 9002 18055
rect 9104 18021 9138 18055
rect 9240 18021 9274 18055
rect 7880 17885 7914 17919
rect 8016 17885 8050 17919
rect 8152 17885 8186 17919
rect 8288 17885 8322 17919
rect 8424 17885 8458 17919
rect 8560 17885 8594 17919
rect 8696 17885 8730 17919
rect 8832 17885 8866 17919
rect 8968 17885 9002 17919
rect 9104 17885 9138 17919
rect 9240 17885 9274 17919
rect 7880 17749 7914 17783
rect 8016 17749 8050 17783
rect 8152 17749 8186 17783
rect 8288 17749 8322 17783
rect 8424 17749 8458 17783
rect 8560 17749 8594 17783
rect 8696 17749 8730 17783
rect 8832 17749 8866 17783
rect 8968 17749 9002 17783
rect 9104 17749 9138 17783
rect 9240 17749 9274 17783
rect 7880 17613 7914 17647
rect 8016 17613 8050 17647
rect 8152 17613 8186 17647
rect 8288 17613 8322 17647
rect 8424 17613 8458 17647
rect 8560 17613 8594 17647
rect 8696 17613 8730 17647
rect 8832 17613 8866 17647
rect 8968 17613 9002 17647
rect 9104 17613 9138 17647
rect 9240 17613 9274 17647
rect 7880 17477 7914 17511
rect 8016 17477 8050 17511
rect 8152 17477 8186 17511
rect 8288 17477 8322 17511
rect 8424 17477 8458 17511
rect 8560 17477 8594 17511
rect 8696 17477 8730 17511
rect 8832 17477 8866 17511
rect 8968 17477 9002 17511
rect 9104 17477 9138 17511
rect 9240 17477 9274 17511
rect 7880 17341 7914 17375
rect 8016 17341 8050 17375
rect 8152 17341 8186 17375
rect 8288 17341 8322 17375
rect 8424 17341 8458 17375
rect 8560 17341 8594 17375
rect 8696 17341 8730 17375
rect 8832 17341 8866 17375
rect 8968 17341 9002 17375
rect 9104 17341 9138 17375
rect 9240 17341 9274 17375
rect 7880 17205 7914 17239
rect 8016 17205 8050 17239
rect 8152 17205 8186 17239
rect 8288 17205 8322 17239
rect 8424 17205 8458 17239
rect 8560 17205 8594 17239
rect 8696 17205 8730 17239
rect 8832 17205 8866 17239
rect 8968 17205 9002 17239
rect 9104 17205 9138 17239
rect 9240 17205 9274 17239
rect 7880 17069 7914 17103
rect 8016 17069 8050 17103
rect 8152 17069 8186 17103
rect 8288 17069 8322 17103
rect 8424 17069 8458 17103
rect 8560 17069 8594 17103
rect 8696 17069 8730 17103
rect 8832 17069 8866 17103
rect 8968 17069 9002 17103
rect 9104 17069 9138 17103
rect 9240 17069 9274 17103
rect 7880 16933 7914 16967
rect 8016 16933 8050 16967
rect 8152 16933 8186 16967
rect 8288 16933 8322 16967
rect 8424 16933 8458 16967
rect 8560 16933 8594 16967
rect 8696 16933 8730 16967
rect 8832 16933 8866 16967
rect 8968 16933 9002 16967
rect 9104 16933 9138 16967
rect 9240 16933 9274 16967
rect 7880 16797 7914 16831
rect 8016 16797 8050 16831
rect 8152 16797 8186 16831
rect 8288 16797 8322 16831
rect 8424 16797 8458 16831
rect 8560 16797 8594 16831
rect 8696 16797 8730 16831
rect 8832 16797 8866 16831
rect 8968 16797 9002 16831
rect 9104 16797 9138 16831
rect 9240 16797 9274 16831
rect 7880 16661 7914 16695
rect 8016 16661 8050 16695
rect 8152 16661 8186 16695
rect 8288 16661 8322 16695
rect 8424 16661 8458 16695
rect 8560 16661 8594 16695
rect 8696 16661 8730 16695
rect 8832 16661 8866 16695
rect 8968 16661 9002 16695
rect 9104 16661 9138 16695
rect 9240 16661 9274 16695
rect 7880 16525 7914 16559
rect 8016 16525 8050 16559
rect 8152 16525 8186 16559
rect 8288 16525 8322 16559
rect 8424 16525 8458 16559
rect 8560 16525 8594 16559
rect 8696 16525 8730 16559
rect 8832 16525 8866 16559
rect 8968 16525 9002 16559
rect 9104 16525 9138 16559
rect 9240 16525 9274 16559
rect 325 16389 359 16423
rect 461 16389 495 16423
rect 597 16389 631 16423
rect 733 16389 767 16423
rect 869 16389 903 16423
rect 1005 16389 1039 16423
rect 1141 16389 1175 16423
rect 1277 16389 1311 16423
rect 1413 16389 1447 16423
rect 1549 16389 1583 16423
rect 1685 16389 1719 16423
rect 325 16253 359 16287
rect 461 16253 495 16287
rect 597 16253 631 16287
rect 733 16253 767 16287
rect 869 16253 903 16287
rect 1005 16253 1039 16287
rect 1141 16253 1175 16287
rect 1277 16253 1311 16287
rect 1413 16253 1447 16287
rect 1549 16253 1583 16287
rect 1685 16253 1719 16287
rect 325 16117 359 16151
rect 461 16117 495 16151
rect 597 16117 631 16151
rect 733 16117 767 16151
rect 869 16117 903 16151
rect 1005 16117 1039 16151
rect 1141 16117 1175 16151
rect 1277 16117 1311 16151
rect 1413 16117 1447 16151
rect 1549 16117 1583 16151
rect 1685 16117 1719 16151
rect 325 15981 359 16015
rect 461 15981 495 16015
rect 597 15981 631 16015
rect 733 15981 767 16015
rect 869 15981 903 16015
rect 1005 15981 1039 16015
rect 1141 15981 1175 16015
rect 1277 15981 1311 16015
rect 1413 15981 1447 16015
rect 1549 15981 1583 16015
rect 1685 15981 1719 16015
rect 325 15845 359 15879
rect 461 15845 495 15879
rect 597 15845 631 15879
rect 733 15845 767 15879
rect 869 15845 903 15879
rect 1005 15845 1039 15879
rect 1141 15845 1175 15879
rect 1277 15845 1311 15879
rect 1413 15845 1447 15879
rect 1549 15845 1583 15879
rect 1685 15845 1719 15879
rect 325 15709 359 15743
rect 461 15709 495 15743
rect 597 15709 631 15743
rect 733 15709 767 15743
rect 869 15709 903 15743
rect 1005 15709 1039 15743
rect 1141 15709 1175 15743
rect 1277 15709 1311 15743
rect 1413 15709 1447 15743
rect 1549 15709 1583 15743
rect 1685 15709 1719 15743
rect 325 15573 359 15607
rect 461 15573 495 15607
rect 597 15573 631 15607
rect 733 15573 767 15607
rect 869 15573 903 15607
rect 1005 15573 1039 15607
rect 1141 15573 1175 15607
rect 1277 15573 1311 15607
rect 1413 15573 1447 15607
rect 1549 15573 1583 15607
rect 1685 15573 1719 15607
rect 325 15437 359 15471
rect 461 15437 495 15471
rect 597 15437 631 15471
rect 733 15437 767 15471
rect 869 15437 903 15471
rect 1005 15437 1039 15471
rect 1141 15437 1175 15471
rect 1277 15437 1311 15471
rect 1413 15437 1447 15471
rect 1549 15437 1583 15471
rect 1685 15437 1719 15471
rect 325 15301 359 15335
rect 461 15301 495 15335
rect 597 15301 631 15335
rect 733 15301 767 15335
rect 869 15301 903 15335
rect 1005 15301 1039 15335
rect 1141 15301 1175 15335
rect 1277 15301 1311 15335
rect 1413 15301 1447 15335
rect 1549 15301 1583 15335
rect 1685 15301 1719 15335
rect 325 15165 359 15199
rect 461 15165 495 15199
rect 597 15165 631 15199
rect 733 15165 767 15199
rect 869 15165 903 15199
rect 1005 15165 1039 15199
rect 1141 15165 1175 15199
rect 1277 15165 1311 15199
rect 1413 15165 1447 15199
rect 1549 15165 1583 15199
rect 1685 15165 1719 15199
rect 325 15029 359 15063
rect 461 15029 495 15063
rect 597 15029 631 15063
rect 733 15029 767 15063
rect 869 15029 903 15063
rect 1005 15029 1039 15063
rect 1141 15029 1175 15063
rect 1277 15029 1311 15063
rect 1413 15029 1447 15063
rect 1549 15029 1583 15063
rect 1685 15029 1719 15063
rect 325 14893 359 14927
rect 461 14893 495 14927
rect 597 14893 631 14927
rect 733 14893 767 14927
rect 869 14893 903 14927
rect 1005 14893 1039 14927
rect 1141 14893 1175 14927
rect 1277 14893 1311 14927
rect 1413 14893 1447 14927
rect 1549 14893 1583 14927
rect 1685 14893 1719 14927
rect 325 14757 359 14791
rect 461 14757 495 14791
rect 597 14757 631 14791
rect 733 14757 767 14791
rect 869 14757 903 14791
rect 1005 14757 1039 14791
rect 1141 14757 1175 14791
rect 1277 14757 1311 14791
rect 1413 14757 1447 14791
rect 1549 14757 1583 14791
rect 1685 14757 1719 14791
rect 325 14621 359 14655
rect 461 14621 495 14655
rect 597 14621 631 14655
rect 733 14621 767 14655
rect 869 14621 903 14655
rect 1005 14621 1039 14655
rect 1141 14621 1175 14655
rect 1277 14621 1311 14655
rect 1413 14621 1447 14655
rect 1549 14621 1583 14655
rect 1685 14621 1719 14655
rect 325 14485 359 14519
rect 461 14485 495 14519
rect 597 14485 631 14519
rect 733 14485 767 14519
rect 869 14485 903 14519
rect 1005 14485 1039 14519
rect 1141 14485 1175 14519
rect 1277 14485 1311 14519
rect 1413 14485 1447 14519
rect 1549 14485 1583 14519
rect 1685 14485 1719 14519
rect 325 14349 359 14383
rect 461 14349 495 14383
rect 597 14349 631 14383
rect 733 14349 767 14383
rect 869 14349 903 14383
rect 1005 14349 1039 14383
rect 1141 14349 1175 14383
rect 1277 14349 1311 14383
rect 1413 14349 1447 14383
rect 1549 14349 1583 14383
rect 1685 14349 1719 14383
rect 325 14213 359 14247
rect 461 14213 495 14247
rect 597 14213 631 14247
rect 733 14213 767 14247
rect 869 14213 903 14247
rect 1005 14213 1039 14247
rect 1141 14213 1175 14247
rect 1277 14213 1311 14247
rect 1413 14213 1447 14247
rect 1549 14213 1583 14247
rect 1685 14213 1719 14247
rect 325 14077 359 14111
rect 461 14077 495 14111
rect 597 14077 631 14111
rect 733 14077 767 14111
rect 869 14077 903 14111
rect 1005 14077 1039 14111
rect 1141 14077 1175 14111
rect 1277 14077 1311 14111
rect 1413 14077 1447 14111
rect 1549 14077 1583 14111
rect 1685 14077 1719 14111
rect 325 13941 359 13975
rect 461 13941 495 13975
rect 597 13941 631 13975
rect 733 13941 767 13975
rect 869 13941 903 13975
rect 1005 13941 1039 13975
rect 1141 13941 1175 13975
rect 1277 13941 1311 13975
rect 1413 13941 1447 13975
rect 1549 13941 1583 13975
rect 1685 13941 1719 13975
rect 325 13805 359 13839
rect 461 13805 495 13839
rect 597 13805 631 13839
rect 733 13805 767 13839
rect 869 13805 903 13839
rect 1005 13805 1039 13839
rect 1141 13805 1175 13839
rect 1277 13805 1311 13839
rect 1413 13805 1447 13839
rect 1549 13805 1583 13839
rect 1685 13805 1719 13839
rect 325 13669 359 13703
rect 461 13669 495 13703
rect 597 13669 631 13703
rect 733 13669 767 13703
rect 869 13669 903 13703
rect 1005 13669 1039 13703
rect 1141 13669 1175 13703
rect 1277 13669 1311 13703
rect 1413 13669 1447 13703
rect 1549 13669 1583 13703
rect 1685 13669 1719 13703
rect 325 13533 359 13567
rect 461 13533 495 13567
rect 597 13533 631 13567
rect 733 13533 767 13567
rect 869 13533 903 13567
rect 1005 13533 1039 13567
rect 1141 13533 1175 13567
rect 1277 13533 1311 13567
rect 1413 13533 1447 13567
rect 1549 13533 1583 13567
rect 1685 13533 1719 13567
rect 325 13397 359 13431
rect 461 13397 495 13431
rect 597 13397 631 13431
rect 733 13397 767 13431
rect 869 13397 903 13431
rect 1005 13397 1039 13431
rect 1141 13397 1175 13431
rect 1277 13397 1311 13431
rect 1413 13397 1447 13431
rect 1549 13397 1583 13431
rect 1685 13397 1719 13431
rect 325 13261 359 13295
rect 461 13261 495 13295
rect 597 13261 631 13295
rect 733 13261 767 13295
rect 869 13261 903 13295
rect 1005 13261 1039 13295
rect 1141 13261 1175 13295
rect 1277 13261 1311 13295
rect 1413 13261 1447 13295
rect 1549 13261 1583 13295
rect 1685 13261 1719 13295
rect 325 13125 359 13159
rect 461 13125 495 13159
rect 597 13125 631 13159
rect 733 13125 767 13159
rect 869 13125 903 13159
rect 1005 13125 1039 13159
rect 1141 13125 1175 13159
rect 1277 13125 1311 13159
rect 1413 13125 1447 13159
rect 1549 13125 1583 13159
rect 1685 13125 1719 13159
rect 325 12989 359 13023
rect 461 12989 495 13023
rect 597 12989 631 13023
rect 733 12989 767 13023
rect 869 12989 903 13023
rect 1005 12989 1039 13023
rect 1141 12989 1175 13023
rect 1277 12989 1311 13023
rect 1413 12989 1447 13023
rect 1549 12989 1583 13023
rect 1685 12989 1719 13023
rect 325 12853 359 12887
rect 461 12853 495 12887
rect 597 12853 631 12887
rect 733 12853 767 12887
rect 869 12853 903 12887
rect 1005 12853 1039 12887
rect 1141 12853 1175 12887
rect 1277 12853 1311 12887
rect 1413 12853 1447 12887
rect 1549 12853 1583 12887
rect 1685 12853 1719 12887
rect 325 12717 359 12751
rect 461 12717 495 12751
rect 597 12717 631 12751
rect 733 12717 767 12751
rect 869 12717 903 12751
rect 1005 12717 1039 12751
rect 1141 12717 1175 12751
rect 1277 12717 1311 12751
rect 1413 12717 1447 12751
rect 1549 12717 1583 12751
rect 1685 12717 1719 12751
rect 325 12581 359 12615
rect 461 12581 495 12615
rect 597 12581 631 12615
rect 733 12581 767 12615
rect 869 12581 903 12615
rect 1005 12581 1039 12615
rect 1141 12581 1175 12615
rect 1277 12581 1311 12615
rect 1413 12581 1447 12615
rect 1549 12581 1583 12615
rect 1685 12581 1719 12615
rect 325 12445 359 12479
rect 461 12445 495 12479
rect 597 12445 631 12479
rect 733 12445 767 12479
rect 869 12445 903 12479
rect 1005 12445 1039 12479
rect 1141 12445 1175 12479
rect 1277 12445 1311 12479
rect 1413 12445 1447 12479
rect 1549 12445 1583 12479
rect 1685 12445 1719 12479
rect 325 12309 359 12343
rect 461 12309 495 12343
rect 597 12309 631 12343
rect 733 12309 767 12343
rect 869 12309 903 12343
rect 1005 12309 1039 12343
rect 1141 12309 1175 12343
rect 1277 12309 1311 12343
rect 1413 12309 1447 12343
rect 1549 12309 1583 12343
rect 1685 12309 1719 12343
rect 325 12173 359 12207
rect 461 12173 495 12207
rect 597 12173 631 12207
rect 733 12173 767 12207
rect 869 12173 903 12207
rect 1005 12173 1039 12207
rect 1141 12173 1175 12207
rect 1277 12173 1311 12207
rect 1413 12173 1447 12207
rect 1549 12173 1583 12207
rect 1685 12173 1719 12207
rect 325 12037 359 12071
rect 461 12037 495 12071
rect 597 12037 631 12071
rect 733 12037 767 12071
rect 869 12037 903 12071
rect 1005 12037 1039 12071
rect 1141 12037 1175 12071
rect 1277 12037 1311 12071
rect 1413 12037 1447 12071
rect 1549 12037 1583 12071
rect 1685 12037 1719 12071
rect 325 11901 359 11935
rect 461 11901 495 11935
rect 597 11901 631 11935
rect 733 11901 767 11935
rect 869 11901 903 11935
rect 1005 11901 1039 11935
rect 1141 11901 1175 11935
rect 1277 11901 1311 11935
rect 1413 11901 1447 11935
rect 1549 11901 1583 11935
rect 1685 11901 1719 11935
rect 325 11765 359 11799
rect 461 11765 495 11799
rect 597 11765 631 11799
rect 733 11765 767 11799
rect 869 11765 903 11799
rect 1005 11765 1039 11799
rect 1141 11765 1175 11799
rect 1277 11765 1311 11799
rect 1413 11765 1447 11799
rect 1549 11765 1583 11799
rect 1685 11765 1719 11799
rect 325 11629 359 11663
rect 461 11629 495 11663
rect 597 11629 631 11663
rect 733 11629 767 11663
rect 869 11629 903 11663
rect 1005 11629 1039 11663
rect 1141 11629 1175 11663
rect 1277 11629 1311 11663
rect 1413 11629 1447 11663
rect 1549 11629 1583 11663
rect 1685 11629 1719 11663
rect 325 11493 359 11527
rect 461 11493 495 11527
rect 597 11493 631 11527
rect 733 11493 767 11527
rect 869 11493 903 11527
rect 1005 11493 1039 11527
rect 1141 11493 1175 11527
rect 1277 11493 1311 11527
rect 1413 11493 1447 11527
rect 1549 11493 1583 11527
rect 1685 11493 1719 11527
rect 325 11357 359 11391
rect 461 11357 495 11391
rect 597 11357 631 11391
rect 733 11357 767 11391
rect 869 11357 903 11391
rect 1005 11357 1039 11391
rect 1141 11357 1175 11391
rect 1277 11357 1311 11391
rect 1413 11357 1447 11391
rect 1549 11357 1583 11391
rect 1685 11357 1719 11391
rect 325 11221 359 11255
rect 461 11221 495 11255
rect 597 11221 631 11255
rect 733 11221 767 11255
rect 869 11221 903 11255
rect 1005 11221 1039 11255
rect 1141 11221 1175 11255
rect 1277 11221 1311 11255
rect 1413 11221 1447 11255
rect 1549 11221 1583 11255
rect 1685 11221 1719 11255
rect 325 11085 359 11119
rect 461 11085 495 11119
rect 597 11085 631 11119
rect 733 11085 767 11119
rect 869 11085 903 11119
rect 1005 11085 1039 11119
rect 1141 11085 1175 11119
rect 1277 11085 1311 11119
rect 1413 11085 1447 11119
rect 1549 11085 1583 11119
rect 1685 11085 1719 11119
rect 325 10949 359 10983
rect 461 10949 495 10983
rect 597 10949 631 10983
rect 733 10949 767 10983
rect 869 10949 903 10983
rect 1005 10949 1039 10983
rect 1141 10949 1175 10983
rect 1277 10949 1311 10983
rect 1413 10949 1447 10983
rect 1549 10949 1583 10983
rect 1685 10949 1719 10983
rect 325 10813 359 10847
rect 461 10813 495 10847
rect 597 10813 631 10847
rect 733 10813 767 10847
rect 869 10813 903 10847
rect 1005 10813 1039 10847
rect 1141 10813 1175 10847
rect 1277 10813 1311 10847
rect 1413 10813 1447 10847
rect 1549 10813 1583 10847
rect 1685 10813 1719 10847
rect 325 10677 359 10711
rect 461 10677 495 10711
rect 597 10677 631 10711
rect 733 10677 767 10711
rect 869 10677 903 10711
rect 1005 10677 1039 10711
rect 1141 10677 1175 10711
rect 1277 10677 1311 10711
rect 1413 10677 1447 10711
rect 1549 10677 1583 10711
rect 1685 10677 1719 10711
rect 325 10541 359 10575
rect 461 10541 495 10575
rect 597 10541 631 10575
rect 733 10541 767 10575
rect 869 10541 903 10575
rect 1005 10541 1039 10575
rect 1141 10541 1175 10575
rect 1277 10541 1311 10575
rect 1413 10541 1447 10575
rect 1549 10541 1583 10575
rect 1685 10541 1719 10575
rect 325 10405 359 10439
rect 461 10405 495 10439
rect 597 10405 631 10439
rect 733 10405 767 10439
rect 869 10405 903 10439
rect 1005 10405 1039 10439
rect 1141 10405 1175 10439
rect 1277 10405 1311 10439
rect 1413 10405 1447 10439
rect 1549 10405 1583 10439
rect 1685 10405 1719 10439
rect 325 10269 359 10303
rect 461 10269 495 10303
rect 597 10269 631 10303
rect 733 10269 767 10303
rect 869 10269 903 10303
rect 1005 10269 1039 10303
rect 1141 10269 1175 10303
rect 1277 10269 1311 10303
rect 1413 10269 1447 10303
rect 1549 10269 1583 10303
rect 1685 10269 1719 10303
rect 325 10133 359 10167
rect 461 10133 495 10167
rect 597 10133 631 10167
rect 733 10133 767 10167
rect 869 10133 903 10167
rect 1005 10133 1039 10167
rect 1141 10133 1175 10167
rect 1277 10133 1311 10167
rect 1413 10133 1447 10167
rect 1549 10133 1583 10167
rect 1685 10133 1719 10167
rect 325 9997 359 10031
rect 461 9997 495 10031
rect 597 9997 631 10031
rect 733 9997 767 10031
rect 869 9997 903 10031
rect 1005 9997 1039 10031
rect 1141 9997 1175 10031
rect 1277 9997 1311 10031
rect 1413 9997 1447 10031
rect 1549 9997 1583 10031
rect 1685 9997 1719 10031
rect 325 9861 359 9895
rect 461 9861 495 9895
rect 597 9861 631 9895
rect 733 9861 767 9895
rect 869 9861 903 9895
rect 1005 9861 1039 9895
rect 1141 9861 1175 9895
rect 1277 9861 1311 9895
rect 1413 9861 1447 9895
rect 1549 9861 1583 9895
rect 1685 9861 1719 9895
rect 325 9725 359 9759
rect 461 9725 495 9759
rect 597 9725 631 9759
rect 733 9725 767 9759
rect 869 9725 903 9759
rect 1005 9725 1039 9759
rect 1141 9725 1175 9759
rect 1277 9725 1311 9759
rect 1413 9725 1447 9759
rect 1549 9725 1583 9759
rect 1685 9725 1719 9759
rect 325 9589 359 9623
rect 461 9589 495 9623
rect 597 9589 631 9623
rect 733 9589 767 9623
rect 869 9589 903 9623
rect 1005 9589 1039 9623
rect 1141 9589 1175 9623
rect 1277 9589 1311 9623
rect 1413 9589 1447 9623
rect 1549 9589 1583 9623
rect 1685 9589 1719 9623
rect 325 9453 359 9487
rect 461 9453 495 9487
rect 597 9453 631 9487
rect 733 9453 767 9487
rect 869 9453 903 9487
rect 1005 9453 1039 9487
rect 1141 9453 1175 9487
rect 1277 9453 1311 9487
rect 1413 9453 1447 9487
rect 1549 9453 1583 9487
rect 1685 9453 1719 9487
rect 325 9317 359 9351
rect 461 9317 495 9351
rect 597 9317 631 9351
rect 733 9317 767 9351
rect 869 9317 903 9351
rect 1005 9317 1039 9351
rect 1141 9317 1175 9351
rect 1277 9317 1311 9351
rect 1413 9317 1447 9351
rect 1549 9317 1583 9351
rect 1685 9317 1719 9351
rect 325 9181 359 9215
rect 461 9181 495 9215
rect 597 9181 631 9215
rect 733 9181 767 9215
rect 869 9181 903 9215
rect 1005 9181 1039 9215
rect 1141 9181 1175 9215
rect 1277 9181 1311 9215
rect 1413 9181 1447 9215
rect 1549 9181 1583 9215
rect 1685 9181 1719 9215
rect 325 9045 359 9079
rect 461 9045 495 9079
rect 597 9045 631 9079
rect 733 9045 767 9079
rect 869 9045 903 9079
rect 1005 9045 1039 9079
rect 1141 9045 1175 9079
rect 1277 9045 1311 9079
rect 1413 9045 1447 9079
rect 1549 9045 1583 9079
rect 1685 9045 1719 9079
rect 325 8909 359 8943
rect 461 8909 495 8943
rect 597 8909 631 8943
rect 733 8909 767 8943
rect 869 8909 903 8943
rect 1005 8909 1039 8943
rect 1141 8909 1175 8943
rect 1277 8909 1311 8943
rect 1413 8909 1447 8943
rect 1549 8909 1583 8943
rect 1685 8909 1719 8943
rect 325 8773 359 8807
rect 461 8773 495 8807
rect 597 8773 631 8807
rect 733 8773 767 8807
rect 869 8773 903 8807
rect 1005 8773 1039 8807
rect 1141 8773 1175 8807
rect 1277 8773 1311 8807
rect 1413 8773 1447 8807
rect 1549 8773 1583 8807
rect 1685 8773 1719 8807
rect 325 8637 359 8671
rect 461 8637 495 8671
rect 597 8637 631 8671
rect 733 8637 767 8671
rect 869 8637 903 8671
rect 1005 8637 1039 8671
rect 1141 8637 1175 8671
rect 1277 8637 1311 8671
rect 1413 8637 1447 8671
rect 1549 8637 1583 8671
rect 1685 8637 1719 8671
rect 325 8501 359 8535
rect 461 8501 495 8535
rect 597 8501 631 8535
rect 733 8501 767 8535
rect 869 8501 903 8535
rect 1005 8501 1039 8535
rect 1141 8501 1175 8535
rect 1277 8501 1311 8535
rect 1413 8501 1447 8535
rect 1549 8501 1583 8535
rect 1685 8501 1719 8535
rect 325 8365 359 8399
rect 461 8365 495 8399
rect 597 8365 631 8399
rect 733 8365 767 8399
rect 869 8365 903 8399
rect 1005 8365 1039 8399
rect 1141 8365 1175 8399
rect 1277 8365 1311 8399
rect 1413 8365 1447 8399
rect 1549 8365 1583 8399
rect 1685 8365 1719 8399
rect 325 8229 359 8263
rect 461 8229 495 8263
rect 597 8229 631 8263
rect 733 8229 767 8263
rect 869 8229 903 8263
rect 1005 8229 1039 8263
rect 1141 8229 1175 8263
rect 1277 8229 1311 8263
rect 1413 8229 1447 8263
rect 1549 8229 1583 8263
rect 1685 8229 1719 8263
rect 325 8093 359 8127
rect 461 8093 495 8127
rect 597 8093 631 8127
rect 733 8093 767 8127
rect 869 8093 903 8127
rect 1005 8093 1039 8127
rect 1141 8093 1175 8127
rect 1277 8093 1311 8127
rect 1413 8093 1447 8127
rect 1549 8093 1583 8127
rect 1685 8093 1719 8127
rect 325 7957 359 7991
rect 461 7957 495 7991
rect 597 7957 631 7991
rect 733 7957 767 7991
rect 869 7957 903 7991
rect 1005 7957 1039 7991
rect 1141 7957 1175 7991
rect 1277 7957 1311 7991
rect 1413 7957 1447 7991
rect 1549 7957 1583 7991
rect 1685 7957 1719 7991
rect 325 7821 359 7855
rect 461 7821 495 7855
rect 597 7821 631 7855
rect 733 7821 767 7855
rect 869 7821 903 7855
rect 1005 7821 1039 7855
rect 1141 7821 1175 7855
rect 1277 7821 1311 7855
rect 1413 7821 1447 7855
rect 1549 7821 1583 7855
rect 1685 7821 1719 7855
rect 325 7685 359 7719
rect 461 7685 495 7719
rect 597 7685 631 7719
rect 733 7685 767 7719
rect 869 7685 903 7719
rect 1005 7685 1039 7719
rect 1141 7685 1175 7719
rect 1277 7685 1311 7719
rect 1413 7685 1447 7719
rect 1549 7685 1583 7719
rect 1685 7685 1719 7719
rect 325 7549 359 7583
rect 461 7549 495 7583
rect 597 7549 631 7583
rect 733 7549 767 7583
rect 869 7549 903 7583
rect 1005 7549 1039 7583
rect 1141 7549 1175 7583
rect 1277 7549 1311 7583
rect 1413 7549 1447 7583
rect 1549 7549 1583 7583
rect 1685 7549 1719 7583
rect 325 7413 359 7447
rect 461 7413 495 7447
rect 597 7413 631 7447
rect 733 7413 767 7447
rect 869 7413 903 7447
rect 1005 7413 1039 7447
rect 1141 7413 1175 7447
rect 1277 7413 1311 7447
rect 1413 7413 1447 7447
rect 1549 7413 1583 7447
rect 1685 7413 1719 7447
rect 325 7277 359 7311
rect 461 7277 495 7311
rect 597 7277 631 7311
rect 733 7277 767 7311
rect 869 7277 903 7311
rect 1005 7277 1039 7311
rect 1141 7277 1175 7311
rect 1277 7277 1311 7311
rect 1413 7277 1447 7311
rect 1549 7277 1583 7311
rect 1685 7277 1719 7311
rect 325 7141 359 7175
rect 461 7141 495 7175
rect 597 7141 631 7175
rect 733 7141 767 7175
rect 869 7141 903 7175
rect 1005 7141 1039 7175
rect 1141 7141 1175 7175
rect 1277 7141 1311 7175
rect 1413 7141 1447 7175
rect 1549 7141 1583 7175
rect 1685 7141 1719 7175
rect 325 7005 359 7039
rect 461 7005 495 7039
rect 597 7005 631 7039
rect 733 7005 767 7039
rect 869 7005 903 7039
rect 1005 7005 1039 7039
rect 1141 7005 1175 7039
rect 1277 7005 1311 7039
rect 1413 7005 1447 7039
rect 1549 7005 1583 7039
rect 1685 7005 1719 7039
rect 325 6869 359 6903
rect 461 6869 495 6903
rect 597 6869 631 6903
rect 733 6869 767 6903
rect 869 6869 903 6903
rect 1005 6869 1039 6903
rect 1141 6869 1175 6903
rect 1277 6869 1311 6903
rect 1413 6869 1447 6903
rect 1549 6869 1583 6903
rect 1685 6869 1719 6903
rect 325 6733 359 6767
rect 461 6733 495 6767
rect 597 6733 631 6767
rect 733 6733 767 6767
rect 869 6733 903 6767
rect 1005 6733 1039 6767
rect 1141 6733 1175 6767
rect 1277 6733 1311 6767
rect 1413 6733 1447 6767
rect 1549 6733 1583 6767
rect 1685 6733 1719 6767
rect 325 6597 359 6631
rect 461 6597 495 6631
rect 597 6597 631 6631
rect 733 6597 767 6631
rect 869 6597 903 6631
rect 1005 6597 1039 6631
rect 1141 6597 1175 6631
rect 1277 6597 1311 6631
rect 1413 6597 1447 6631
rect 1549 6597 1583 6631
rect 1685 6597 1719 6631
rect 325 6461 359 6495
rect 461 6461 495 6495
rect 597 6461 631 6495
rect 733 6461 767 6495
rect 869 6461 903 6495
rect 1005 6461 1039 6495
rect 1141 6461 1175 6495
rect 1277 6461 1311 6495
rect 1413 6461 1447 6495
rect 1549 6461 1583 6495
rect 1685 6461 1719 6495
rect 325 6325 359 6359
rect 461 6325 495 6359
rect 597 6325 631 6359
rect 733 6325 767 6359
rect 869 6325 903 6359
rect 1005 6325 1039 6359
rect 1141 6325 1175 6359
rect 1277 6325 1311 6359
rect 1413 6325 1447 6359
rect 1549 6325 1583 6359
rect 1685 6325 1719 6359
rect 325 6189 359 6223
rect 461 6189 495 6223
rect 597 6189 631 6223
rect 733 6189 767 6223
rect 869 6189 903 6223
rect 1005 6189 1039 6223
rect 1141 6189 1175 6223
rect 1277 6189 1311 6223
rect 1413 6189 1447 6223
rect 1549 6189 1583 6223
rect 1685 6189 1719 6223
rect 325 6053 359 6087
rect 461 6053 495 6087
rect 597 6053 631 6087
rect 733 6053 767 6087
rect 869 6053 903 6087
rect 1005 6053 1039 6087
rect 1141 6053 1175 6087
rect 1277 6053 1311 6087
rect 1413 6053 1447 6087
rect 1549 6053 1583 6087
rect 1685 6053 1719 6087
rect 325 5917 359 5951
rect 461 5917 495 5951
rect 597 5917 631 5951
rect 733 5917 767 5951
rect 869 5917 903 5951
rect 1005 5917 1039 5951
rect 1141 5917 1175 5951
rect 1277 5917 1311 5951
rect 1413 5917 1447 5951
rect 1549 5917 1583 5951
rect 1685 5917 1719 5951
rect 325 5781 359 5815
rect 461 5781 495 5815
rect 597 5781 631 5815
rect 733 5781 767 5815
rect 869 5781 903 5815
rect 1005 5781 1039 5815
rect 1141 5781 1175 5815
rect 1277 5781 1311 5815
rect 1413 5781 1447 5815
rect 1549 5781 1583 5815
rect 1685 5781 1719 5815
rect 325 5645 359 5679
rect 461 5645 495 5679
rect 597 5645 631 5679
rect 733 5645 767 5679
rect 869 5645 903 5679
rect 1005 5645 1039 5679
rect 1141 5645 1175 5679
rect 1277 5645 1311 5679
rect 1413 5645 1447 5679
rect 1549 5645 1583 5679
rect 1685 5645 1719 5679
rect 325 5509 359 5543
rect 461 5509 495 5543
rect 597 5509 631 5543
rect 733 5509 767 5543
rect 869 5509 903 5543
rect 1005 5509 1039 5543
rect 1141 5509 1175 5543
rect 1277 5509 1311 5543
rect 1413 5509 1447 5543
rect 1549 5509 1583 5543
rect 1685 5509 1719 5543
rect 325 5373 359 5407
rect 461 5373 495 5407
rect 597 5373 631 5407
rect 733 5373 767 5407
rect 869 5373 903 5407
rect 1005 5373 1039 5407
rect 1141 5373 1175 5407
rect 1277 5373 1311 5407
rect 1413 5373 1447 5407
rect 1549 5373 1583 5407
rect 1685 5373 1719 5407
rect 325 5237 359 5271
rect 461 5237 495 5271
rect 597 5237 631 5271
rect 733 5237 767 5271
rect 869 5237 903 5271
rect 1005 5237 1039 5271
rect 1141 5237 1175 5271
rect 1277 5237 1311 5271
rect 1413 5237 1447 5271
rect 1549 5237 1583 5271
rect 1685 5237 1719 5271
rect 325 5101 359 5135
rect 461 5101 495 5135
rect 597 5101 631 5135
rect 733 5101 767 5135
rect 869 5101 903 5135
rect 1005 5101 1039 5135
rect 1141 5101 1175 5135
rect 1277 5101 1311 5135
rect 1413 5101 1447 5135
rect 1549 5101 1583 5135
rect 1685 5101 1719 5135
rect 325 4965 359 4999
rect 461 4965 495 4999
rect 597 4965 631 4999
rect 733 4965 767 4999
rect 869 4965 903 4999
rect 1005 4965 1039 4999
rect 1141 4965 1175 4999
rect 1277 4965 1311 4999
rect 1413 4965 1447 4999
rect 1549 4965 1583 4999
rect 1685 4965 1719 4999
rect 325 4829 359 4863
rect 461 4829 495 4863
rect 597 4829 631 4863
rect 733 4829 767 4863
rect 869 4829 903 4863
rect 1005 4829 1039 4863
rect 1141 4829 1175 4863
rect 1277 4829 1311 4863
rect 1413 4829 1447 4863
rect 1549 4829 1583 4863
rect 1685 4829 1719 4863
rect 325 4693 359 4727
rect 461 4693 495 4727
rect 597 4693 631 4727
rect 733 4693 767 4727
rect 869 4693 903 4727
rect 1005 4693 1039 4727
rect 1141 4693 1175 4727
rect 1277 4693 1311 4727
rect 1413 4693 1447 4727
rect 1549 4693 1583 4727
rect 1685 4693 1719 4727
rect 325 4557 359 4591
rect 461 4557 495 4591
rect 597 4557 631 4591
rect 733 4557 767 4591
rect 869 4557 903 4591
rect 1005 4557 1039 4591
rect 1141 4557 1175 4591
rect 1277 4557 1311 4591
rect 1413 4557 1447 4591
rect 1549 4557 1583 4591
rect 1685 4557 1719 4591
rect 325 4421 359 4455
rect 461 4421 495 4455
rect 597 4421 631 4455
rect 733 4421 767 4455
rect 869 4421 903 4455
rect 1005 4421 1039 4455
rect 1141 4421 1175 4455
rect 1277 4421 1311 4455
rect 1413 4421 1447 4455
rect 1549 4421 1583 4455
rect 1685 4421 1719 4455
rect 325 4285 359 4319
rect 461 4285 495 4319
rect 597 4285 631 4319
rect 733 4285 767 4319
rect 869 4285 903 4319
rect 1005 4285 1039 4319
rect 1141 4285 1175 4319
rect 1277 4285 1311 4319
rect 1413 4285 1447 4319
rect 1549 4285 1583 4319
rect 1685 4285 1719 4319
rect 325 4149 359 4183
rect 461 4149 495 4183
rect 597 4149 631 4183
rect 733 4149 767 4183
rect 869 4149 903 4183
rect 1005 4149 1039 4183
rect 1141 4149 1175 4183
rect 1277 4149 1311 4183
rect 1413 4149 1447 4183
rect 1549 4149 1583 4183
rect 1685 4149 1719 4183
rect 325 4013 359 4047
rect 461 4013 495 4047
rect 597 4013 631 4047
rect 733 4013 767 4047
rect 869 4013 903 4047
rect 1005 4013 1039 4047
rect 1141 4013 1175 4047
rect 1277 4013 1311 4047
rect 1413 4013 1447 4047
rect 1549 4013 1583 4047
rect 1685 4013 1719 4047
rect 325 3877 359 3911
rect 461 3877 495 3911
rect 597 3877 631 3911
rect 733 3877 767 3911
rect 869 3877 903 3911
rect 1005 3877 1039 3911
rect 1141 3877 1175 3911
rect 1277 3877 1311 3911
rect 1413 3877 1447 3911
rect 1549 3877 1583 3911
rect 1685 3877 1719 3911
rect 325 3741 359 3775
rect 461 3741 495 3775
rect 597 3741 631 3775
rect 733 3741 767 3775
rect 869 3741 903 3775
rect 1005 3741 1039 3775
rect 1141 3741 1175 3775
rect 1277 3741 1311 3775
rect 1413 3741 1447 3775
rect 1549 3741 1583 3775
rect 1685 3741 1719 3775
rect 325 3605 359 3639
rect 461 3605 495 3639
rect 597 3605 631 3639
rect 733 3605 767 3639
rect 869 3605 903 3639
rect 1005 3605 1039 3639
rect 1141 3605 1175 3639
rect 1277 3605 1311 3639
rect 1413 3605 1447 3639
rect 1549 3605 1583 3639
rect 1685 3605 1719 3639
rect 325 3469 359 3503
rect 461 3469 495 3503
rect 597 3469 631 3503
rect 733 3469 767 3503
rect 869 3469 903 3503
rect 1005 3469 1039 3503
rect 1141 3469 1175 3503
rect 1277 3469 1311 3503
rect 1413 3469 1447 3503
rect 1549 3469 1583 3503
rect 1685 3469 1719 3503
rect 325 3333 359 3367
rect 461 3333 495 3367
rect 597 3333 631 3367
rect 733 3333 767 3367
rect 869 3333 903 3367
rect 1005 3333 1039 3367
rect 1141 3333 1175 3367
rect 1277 3333 1311 3367
rect 1413 3333 1447 3367
rect 1549 3333 1583 3367
rect 1685 3333 1719 3367
rect 325 3197 359 3231
rect 461 3197 495 3231
rect 597 3197 631 3231
rect 733 3197 767 3231
rect 869 3197 903 3231
rect 1005 3197 1039 3231
rect 1141 3197 1175 3231
rect 1277 3197 1311 3231
rect 1413 3197 1447 3231
rect 1549 3197 1583 3231
rect 1685 3197 1719 3231
rect 325 3061 359 3095
rect 461 3061 495 3095
rect 597 3061 631 3095
rect 733 3061 767 3095
rect 869 3061 903 3095
rect 1005 3061 1039 3095
rect 1141 3061 1175 3095
rect 1277 3061 1311 3095
rect 1413 3061 1447 3095
rect 1549 3061 1583 3095
rect 1685 3061 1719 3095
rect 325 2925 359 2959
rect 461 2925 495 2959
rect 597 2925 631 2959
rect 733 2925 767 2959
rect 869 2925 903 2959
rect 1005 2925 1039 2959
rect 1141 2925 1175 2959
rect 1277 2925 1311 2959
rect 1413 2925 1447 2959
rect 1549 2925 1583 2959
rect 1685 2925 1719 2959
rect 325 2789 359 2823
rect 461 2789 495 2823
rect 597 2789 631 2823
rect 733 2789 767 2823
rect 869 2789 903 2823
rect 1005 2789 1039 2823
rect 1141 2789 1175 2823
rect 1277 2789 1311 2823
rect 1413 2789 1447 2823
rect 1549 2789 1583 2823
rect 1685 2789 1719 2823
rect 325 2653 359 2687
rect 461 2653 495 2687
rect 597 2653 631 2687
rect 733 2653 767 2687
rect 869 2653 903 2687
rect 1005 2653 1039 2687
rect 1141 2653 1175 2687
rect 1277 2653 1311 2687
rect 1413 2653 1447 2687
rect 1549 2653 1583 2687
rect 1685 2653 1719 2687
rect 325 2517 359 2551
rect 461 2517 495 2551
rect 597 2517 631 2551
rect 733 2517 767 2551
rect 869 2517 903 2551
rect 1005 2517 1039 2551
rect 1141 2517 1175 2551
rect 1277 2517 1311 2551
rect 1413 2517 1447 2551
rect 1549 2517 1583 2551
rect 1685 2517 1719 2551
rect 325 2380 359 2414
rect 461 2380 495 2414
rect 597 2380 631 2414
rect 733 2380 767 2414
rect 869 2380 903 2414
rect 1005 2380 1039 2414
rect 1141 2380 1175 2414
rect 1277 2380 1311 2414
rect 1413 2380 1447 2414
rect 1549 2380 1583 2414
rect 1685 2380 1719 2414
rect 325 2243 359 2277
rect 461 2243 495 2277
rect 597 2243 631 2277
rect 733 2243 767 2277
rect 869 2243 903 2277
rect 1005 2243 1039 2277
rect 1141 2243 1175 2277
rect 1277 2243 1311 2277
rect 1413 2243 1447 2277
rect 1549 2243 1583 2277
rect 1685 2243 1719 2277
rect 325 2106 359 2140
rect 461 2106 495 2140
rect 597 2106 631 2140
rect 733 2106 767 2140
rect 869 2106 903 2140
rect 1005 2106 1039 2140
rect 1141 2106 1175 2140
rect 1277 2106 1311 2140
rect 1413 2106 1447 2140
rect 1549 2106 1583 2140
rect 1685 2106 1719 2140
rect 325 1969 359 2003
rect 461 1969 495 2003
rect 597 1969 631 2003
rect 733 1969 767 2003
rect 869 1969 903 2003
rect 1005 1969 1039 2003
rect 1141 1969 1175 2003
rect 1277 1969 1311 2003
rect 1413 1969 1447 2003
rect 1549 1969 1583 2003
rect 1685 1969 1719 2003
rect 325 1832 359 1866
rect 461 1832 495 1866
rect 597 1832 631 1866
rect 733 1832 767 1866
rect 869 1832 903 1866
rect 1005 1832 1039 1866
rect 1141 1832 1175 1866
rect 1277 1832 1311 1866
rect 1413 1832 1447 1866
rect 1549 1832 1583 1866
rect 1685 1832 1719 1866
rect 7880 16389 7914 16423
rect 8016 16389 8050 16423
rect 8152 16389 8186 16423
rect 8288 16389 8322 16423
rect 8424 16389 8458 16423
rect 8560 16389 8594 16423
rect 8696 16389 8730 16423
rect 8832 16389 8866 16423
rect 8968 16389 9002 16423
rect 9104 16389 9138 16423
rect 9240 16389 9274 16423
rect 7880 16253 7914 16287
rect 8016 16253 8050 16287
rect 8152 16253 8186 16287
rect 8288 16253 8322 16287
rect 8424 16253 8458 16287
rect 8560 16253 8594 16287
rect 8696 16253 8730 16287
rect 8832 16253 8866 16287
rect 8968 16253 9002 16287
rect 9104 16253 9138 16287
rect 9240 16253 9274 16287
rect 7880 16117 7914 16151
rect 8016 16117 8050 16151
rect 8152 16117 8186 16151
rect 8288 16117 8322 16151
rect 8424 16117 8458 16151
rect 8560 16117 8594 16151
rect 8696 16117 8730 16151
rect 8832 16117 8866 16151
rect 8968 16117 9002 16151
rect 9104 16117 9138 16151
rect 9240 16117 9274 16151
rect 7880 15981 7914 16015
rect 8016 15981 8050 16015
rect 8152 15981 8186 16015
rect 8288 15981 8322 16015
rect 8424 15981 8458 16015
rect 8560 15981 8594 16015
rect 8696 15981 8730 16015
rect 8832 15981 8866 16015
rect 8968 15981 9002 16015
rect 9104 15981 9138 16015
rect 9240 15981 9274 16015
rect 7880 15845 7914 15879
rect 8016 15845 8050 15879
rect 8152 15845 8186 15879
rect 8288 15845 8322 15879
rect 8424 15845 8458 15879
rect 8560 15845 8594 15879
rect 8696 15845 8730 15879
rect 8832 15845 8866 15879
rect 8968 15845 9002 15879
rect 9104 15845 9138 15879
rect 9240 15845 9274 15879
rect 7880 15709 7914 15743
rect 8016 15709 8050 15743
rect 8152 15709 8186 15743
rect 8288 15709 8322 15743
rect 8424 15709 8458 15743
rect 8560 15709 8594 15743
rect 8696 15709 8730 15743
rect 8832 15709 8866 15743
rect 8968 15709 9002 15743
rect 9104 15709 9138 15743
rect 9240 15709 9274 15743
rect 7880 15573 7914 15607
rect 8016 15573 8050 15607
rect 8152 15573 8186 15607
rect 8288 15573 8322 15607
rect 8424 15573 8458 15607
rect 8560 15573 8594 15607
rect 8696 15573 8730 15607
rect 8832 15573 8866 15607
rect 8968 15573 9002 15607
rect 9104 15573 9138 15607
rect 9240 15573 9274 15607
rect 7880 15437 7914 15471
rect 8016 15437 8050 15471
rect 8152 15437 8186 15471
rect 8288 15437 8322 15471
rect 8424 15437 8458 15471
rect 8560 15437 8594 15471
rect 8696 15437 8730 15471
rect 8832 15437 8866 15471
rect 8968 15437 9002 15471
rect 9104 15437 9138 15471
rect 9240 15437 9274 15471
rect 7880 15301 7914 15335
rect 8016 15301 8050 15335
rect 8152 15301 8186 15335
rect 8288 15301 8322 15335
rect 8424 15301 8458 15335
rect 8560 15301 8594 15335
rect 8696 15301 8730 15335
rect 8832 15301 8866 15335
rect 8968 15301 9002 15335
rect 9104 15301 9138 15335
rect 9240 15301 9274 15335
rect 7880 15165 7914 15199
rect 8016 15165 8050 15199
rect 8152 15165 8186 15199
rect 8288 15165 8322 15199
rect 8424 15165 8458 15199
rect 8560 15165 8594 15199
rect 8696 15165 8730 15199
rect 8832 15165 8866 15199
rect 8968 15165 9002 15199
rect 9104 15165 9138 15199
rect 9240 15165 9274 15199
rect 7880 15029 7914 15063
rect 8016 15029 8050 15063
rect 8152 15029 8186 15063
rect 8288 15029 8322 15063
rect 8424 15029 8458 15063
rect 8560 15029 8594 15063
rect 8696 15029 8730 15063
rect 8832 15029 8866 15063
rect 8968 15029 9002 15063
rect 9104 15029 9138 15063
rect 9240 15029 9274 15063
rect 7880 14893 7914 14927
rect 8016 14893 8050 14927
rect 8152 14893 8186 14927
rect 8288 14893 8322 14927
rect 8424 14893 8458 14927
rect 8560 14893 8594 14927
rect 8696 14893 8730 14927
rect 8832 14893 8866 14927
rect 8968 14893 9002 14927
rect 9104 14893 9138 14927
rect 9240 14893 9274 14927
rect 7880 14757 7914 14791
rect 8016 14757 8050 14791
rect 8152 14757 8186 14791
rect 8288 14757 8322 14791
rect 8424 14757 8458 14791
rect 8560 14757 8594 14791
rect 8696 14757 8730 14791
rect 8832 14757 8866 14791
rect 8968 14757 9002 14791
rect 9104 14757 9138 14791
rect 9240 14757 9274 14791
rect 7880 14621 7914 14655
rect 8016 14621 8050 14655
rect 8152 14621 8186 14655
rect 8288 14621 8322 14655
rect 8424 14621 8458 14655
rect 8560 14621 8594 14655
rect 8696 14621 8730 14655
rect 8832 14621 8866 14655
rect 8968 14621 9002 14655
rect 9104 14621 9138 14655
rect 9240 14621 9274 14655
rect 7880 14485 7914 14519
rect 8016 14485 8050 14519
rect 8152 14485 8186 14519
rect 8288 14485 8322 14519
rect 8424 14485 8458 14519
rect 8560 14485 8594 14519
rect 8696 14485 8730 14519
rect 8832 14485 8866 14519
rect 8968 14485 9002 14519
rect 9104 14485 9138 14519
rect 9240 14485 9274 14519
rect 7880 14349 7914 14383
rect 8016 14349 8050 14383
rect 8152 14349 8186 14383
rect 8288 14349 8322 14383
rect 8424 14349 8458 14383
rect 8560 14349 8594 14383
rect 8696 14349 8730 14383
rect 8832 14349 8866 14383
rect 8968 14349 9002 14383
rect 9104 14349 9138 14383
rect 9240 14349 9274 14383
rect 7880 14213 7914 14247
rect 8016 14213 8050 14247
rect 8152 14213 8186 14247
rect 8288 14213 8322 14247
rect 8424 14213 8458 14247
rect 8560 14213 8594 14247
rect 8696 14213 8730 14247
rect 8832 14213 8866 14247
rect 8968 14213 9002 14247
rect 9104 14213 9138 14247
rect 9240 14213 9274 14247
rect 7880 14077 7914 14111
rect 8016 14077 8050 14111
rect 8152 14077 8186 14111
rect 8288 14077 8322 14111
rect 8424 14077 8458 14111
rect 8560 14077 8594 14111
rect 8696 14077 8730 14111
rect 8832 14077 8866 14111
rect 8968 14077 9002 14111
rect 9104 14077 9138 14111
rect 9240 14077 9274 14111
rect 7880 13941 7914 13975
rect 8016 13941 8050 13975
rect 8152 13941 8186 13975
rect 8288 13941 8322 13975
rect 8424 13941 8458 13975
rect 8560 13941 8594 13975
rect 8696 13941 8730 13975
rect 8832 13941 8866 13975
rect 8968 13941 9002 13975
rect 9104 13941 9138 13975
rect 9240 13941 9274 13975
rect 7880 13805 7914 13839
rect 8016 13805 8050 13839
rect 8152 13805 8186 13839
rect 8288 13805 8322 13839
rect 8424 13805 8458 13839
rect 8560 13805 8594 13839
rect 8696 13805 8730 13839
rect 8832 13805 8866 13839
rect 8968 13805 9002 13839
rect 9104 13805 9138 13839
rect 9240 13805 9274 13839
rect 7880 13669 7914 13703
rect 8016 13669 8050 13703
rect 8152 13669 8186 13703
rect 8288 13669 8322 13703
rect 8424 13669 8458 13703
rect 8560 13669 8594 13703
rect 8696 13669 8730 13703
rect 8832 13669 8866 13703
rect 8968 13669 9002 13703
rect 9104 13669 9138 13703
rect 9240 13669 9274 13703
rect 7880 13533 7914 13567
rect 8016 13533 8050 13567
rect 8152 13533 8186 13567
rect 8288 13533 8322 13567
rect 8424 13533 8458 13567
rect 8560 13533 8594 13567
rect 8696 13533 8730 13567
rect 8832 13533 8866 13567
rect 8968 13533 9002 13567
rect 9104 13533 9138 13567
rect 9240 13533 9274 13567
rect 7880 13397 7914 13431
rect 8016 13397 8050 13431
rect 8152 13397 8186 13431
rect 8288 13397 8322 13431
rect 8424 13397 8458 13431
rect 8560 13397 8594 13431
rect 8696 13397 8730 13431
rect 8832 13397 8866 13431
rect 8968 13397 9002 13431
rect 9104 13397 9138 13431
rect 9240 13397 9274 13431
rect 7880 13261 7914 13295
rect 8016 13261 8050 13295
rect 8152 13261 8186 13295
rect 8288 13261 8322 13295
rect 8424 13261 8458 13295
rect 8560 13261 8594 13295
rect 8696 13261 8730 13295
rect 8832 13261 8866 13295
rect 8968 13261 9002 13295
rect 9104 13261 9138 13295
rect 9240 13261 9274 13295
rect 7880 13125 7914 13159
rect 8016 13125 8050 13159
rect 8152 13125 8186 13159
rect 8288 13125 8322 13159
rect 8424 13125 8458 13159
rect 8560 13125 8594 13159
rect 8696 13125 8730 13159
rect 8832 13125 8866 13159
rect 8968 13125 9002 13159
rect 9104 13125 9138 13159
rect 9240 13125 9274 13159
rect 7880 12989 7914 13023
rect 8016 12989 8050 13023
rect 8152 12989 8186 13023
rect 8288 12989 8322 13023
rect 8424 12989 8458 13023
rect 8560 12989 8594 13023
rect 8696 12989 8730 13023
rect 8832 12989 8866 13023
rect 8968 12989 9002 13023
rect 9104 12989 9138 13023
rect 9240 12989 9274 13023
rect 7880 12853 7914 12887
rect 8016 12853 8050 12887
rect 8152 12853 8186 12887
rect 8288 12853 8322 12887
rect 8424 12853 8458 12887
rect 8560 12853 8594 12887
rect 8696 12853 8730 12887
rect 8832 12853 8866 12887
rect 8968 12853 9002 12887
rect 9104 12853 9138 12887
rect 9240 12853 9274 12887
rect 7880 12717 7914 12751
rect 8016 12717 8050 12751
rect 8152 12717 8186 12751
rect 8288 12717 8322 12751
rect 8424 12717 8458 12751
rect 8560 12717 8594 12751
rect 8696 12717 8730 12751
rect 8832 12717 8866 12751
rect 8968 12717 9002 12751
rect 9104 12717 9138 12751
rect 9240 12717 9274 12751
rect 7880 12581 7914 12615
rect 8016 12581 8050 12615
rect 8152 12581 8186 12615
rect 8288 12581 8322 12615
rect 8424 12581 8458 12615
rect 8560 12581 8594 12615
rect 8696 12581 8730 12615
rect 8832 12581 8866 12615
rect 8968 12581 9002 12615
rect 9104 12581 9138 12615
rect 9240 12581 9274 12615
rect 7880 12445 7914 12479
rect 8016 12445 8050 12479
rect 8152 12445 8186 12479
rect 8288 12445 8322 12479
rect 8424 12445 8458 12479
rect 8560 12445 8594 12479
rect 8696 12445 8730 12479
rect 8832 12445 8866 12479
rect 8968 12445 9002 12479
rect 9104 12445 9138 12479
rect 9240 12445 9274 12479
rect 7880 12309 7914 12343
rect 8016 12309 8050 12343
rect 8152 12309 8186 12343
rect 8288 12309 8322 12343
rect 8424 12309 8458 12343
rect 8560 12309 8594 12343
rect 8696 12309 8730 12343
rect 8832 12309 8866 12343
rect 8968 12309 9002 12343
rect 9104 12309 9138 12343
rect 9240 12309 9274 12343
rect 7880 12173 7914 12207
rect 8016 12173 8050 12207
rect 8152 12173 8186 12207
rect 8288 12173 8322 12207
rect 8424 12173 8458 12207
rect 8560 12173 8594 12207
rect 8696 12173 8730 12207
rect 8832 12173 8866 12207
rect 8968 12173 9002 12207
rect 9104 12173 9138 12207
rect 9240 12173 9274 12207
rect 7880 12037 7914 12071
rect 8016 12037 8050 12071
rect 8152 12037 8186 12071
rect 8288 12037 8322 12071
rect 8424 12037 8458 12071
rect 8560 12037 8594 12071
rect 8696 12037 8730 12071
rect 8832 12037 8866 12071
rect 8968 12037 9002 12071
rect 9104 12037 9138 12071
rect 9240 12037 9274 12071
rect 7880 11901 7914 11935
rect 8016 11901 8050 11935
rect 8152 11901 8186 11935
rect 8288 11901 8322 11935
rect 8424 11901 8458 11935
rect 8560 11901 8594 11935
rect 8696 11901 8730 11935
rect 8832 11901 8866 11935
rect 8968 11901 9002 11935
rect 9104 11901 9138 11935
rect 9240 11901 9274 11935
rect 7880 11765 7914 11799
rect 8016 11765 8050 11799
rect 8152 11765 8186 11799
rect 8288 11765 8322 11799
rect 8424 11765 8458 11799
rect 8560 11765 8594 11799
rect 8696 11765 8730 11799
rect 8832 11765 8866 11799
rect 8968 11765 9002 11799
rect 9104 11765 9138 11799
rect 9240 11765 9274 11799
rect 7880 11629 7914 11663
rect 8016 11629 8050 11663
rect 8152 11629 8186 11663
rect 8288 11629 8322 11663
rect 8424 11629 8458 11663
rect 8560 11629 8594 11663
rect 8696 11629 8730 11663
rect 8832 11629 8866 11663
rect 8968 11629 9002 11663
rect 9104 11629 9138 11663
rect 9240 11629 9274 11663
rect 7880 11493 7914 11527
rect 8016 11493 8050 11527
rect 8152 11493 8186 11527
rect 8288 11493 8322 11527
rect 8424 11493 8458 11527
rect 8560 11493 8594 11527
rect 8696 11493 8730 11527
rect 8832 11493 8866 11527
rect 8968 11493 9002 11527
rect 9104 11493 9138 11527
rect 9240 11493 9274 11527
rect 7880 11357 7914 11391
rect 8016 11357 8050 11391
rect 8152 11357 8186 11391
rect 8288 11357 8322 11391
rect 8424 11357 8458 11391
rect 8560 11357 8594 11391
rect 8696 11357 8730 11391
rect 8832 11357 8866 11391
rect 8968 11357 9002 11391
rect 9104 11357 9138 11391
rect 9240 11357 9274 11391
rect 7880 11221 7914 11255
rect 8016 11221 8050 11255
rect 8152 11221 8186 11255
rect 8288 11221 8322 11255
rect 8424 11221 8458 11255
rect 8560 11221 8594 11255
rect 8696 11221 8730 11255
rect 8832 11221 8866 11255
rect 8968 11221 9002 11255
rect 9104 11221 9138 11255
rect 9240 11221 9274 11255
rect 7880 11085 7914 11119
rect 8016 11085 8050 11119
rect 8152 11085 8186 11119
rect 8288 11085 8322 11119
rect 8424 11085 8458 11119
rect 8560 11085 8594 11119
rect 8696 11085 8730 11119
rect 8832 11085 8866 11119
rect 8968 11085 9002 11119
rect 9104 11085 9138 11119
rect 9240 11085 9274 11119
rect 7880 10949 7914 10983
rect 8016 10949 8050 10983
rect 8152 10949 8186 10983
rect 8288 10949 8322 10983
rect 8424 10949 8458 10983
rect 8560 10949 8594 10983
rect 8696 10949 8730 10983
rect 8832 10949 8866 10983
rect 8968 10949 9002 10983
rect 9104 10949 9138 10983
rect 9240 10949 9274 10983
rect 7880 10813 7914 10847
rect 8016 10813 8050 10847
rect 8152 10813 8186 10847
rect 8288 10813 8322 10847
rect 8424 10813 8458 10847
rect 8560 10813 8594 10847
rect 8696 10813 8730 10847
rect 8832 10813 8866 10847
rect 8968 10813 9002 10847
rect 9104 10813 9138 10847
rect 9240 10813 9274 10847
rect 7880 10677 7914 10711
rect 8016 10677 8050 10711
rect 8152 10677 8186 10711
rect 8288 10677 8322 10711
rect 8424 10677 8458 10711
rect 8560 10677 8594 10711
rect 8696 10677 8730 10711
rect 8832 10677 8866 10711
rect 8968 10677 9002 10711
rect 9104 10677 9138 10711
rect 9240 10677 9274 10711
rect 7880 10541 7914 10575
rect 8016 10541 8050 10575
rect 8152 10541 8186 10575
rect 8288 10541 8322 10575
rect 8424 10541 8458 10575
rect 8560 10541 8594 10575
rect 8696 10541 8730 10575
rect 8832 10541 8866 10575
rect 8968 10541 9002 10575
rect 9104 10541 9138 10575
rect 9240 10541 9274 10575
rect 7880 10405 7914 10439
rect 8016 10405 8050 10439
rect 8152 10405 8186 10439
rect 8288 10405 8322 10439
rect 8424 10405 8458 10439
rect 8560 10405 8594 10439
rect 8696 10405 8730 10439
rect 8832 10405 8866 10439
rect 8968 10405 9002 10439
rect 9104 10405 9138 10439
rect 9240 10405 9274 10439
rect 7880 10269 7914 10303
rect 8016 10269 8050 10303
rect 8152 10269 8186 10303
rect 8288 10269 8322 10303
rect 8424 10269 8458 10303
rect 8560 10269 8594 10303
rect 8696 10269 8730 10303
rect 8832 10269 8866 10303
rect 8968 10269 9002 10303
rect 9104 10269 9138 10303
rect 9240 10269 9274 10303
rect 7880 10133 7914 10167
rect 8016 10133 8050 10167
rect 8152 10133 8186 10167
rect 8288 10133 8322 10167
rect 8424 10133 8458 10167
rect 8560 10133 8594 10167
rect 8696 10133 8730 10167
rect 8832 10133 8866 10167
rect 8968 10133 9002 10167
rect 9104 10133 9138 10167
rect 9240 10133 9274 10167
rect 7880 9997 7914 10031
rect 8016 9997 8050 10031
rect 8152 9997 8186 10031
rect 8288 9997 8322 10031
rect 8424 9997 8458 10031
rect 8560 9997 8594 10031
rect 8696 9997 8730 10031
rect 8832 9997 8866 10031
rect 8968 9997 9002 10031
rect 9104 9997 9138 10031
rect 9240 9997 9274 10031
rect 7880 9861 7914 9895
rect 8016 9861 8050 9895
rect 8152 9861 8186 9895
rect 8288 9861 8322 9895
rect 8424 9861 8458 9895
rect 8560 9861 8594 9895
rect 8696 9861 8730 9895
rect 8832 9861 8866 9895
rect 8968 9861 9002 9895
rect 9104 9861 9138 9895
rect 9240 9861 9274 9895
rect 7880 9725 7914 9759
rect 8016 9725 8050 9759
rect 8152 9725 8186 9759
rect 8288 9725 8322 9759
rect 8424 9725 8458 9759
rect 8560 9725 8594 9759
rect 8696 9725 8730 9759
rect 8832 9725 8866 9759
rect 8968 9725 9002 9759
rect 9104 9725 9138 9759
rect 9240 9725 9274 9759
rect 7880 9589 7914 9623
rect 8016 9589 8050 9623
rect 8152 9589 8186 9623
rect 8288 9589 8322 9623
rect 8424 9589 8458 9623
rect 8560 9589 8594 9623
rect 8696 9589 8730 9623
rect 8832 9589 8866 9623
rect 8968 9589 9002 9623
rect 9104 9589 9138 9623
rect 9240 9589 9274 9623
rect 7880 9453 7914 9487
rect 8016 9453 8050 9487
rect 8152 9453 8186 9487
rect 8288 9453 8322 9487
rect 8424 9453 8458 9487
rect 8560 9453 8594 9487
rect 8696 9453 8730 9487
rect 8832 9453 8866 9487
rect 8968 9453 9002 9487
rect 9104 9453 9138 9487
rect 9240 9453 9274 9487
rect 7880 9317 7914 9351
rect 8016 9317 8050 9351
rect 8152 9317 8186 9351
rect 8288 9317 8322 9351
rect 8424 9317 8458 9351
rect 8560 9317 8594 9351
rect 8696 9317 8730 9351
rect 8832 9317 8866 9351
rect 8968 9317 9002 9351
rect 9104 9317 9138 9351
rect 9240 9317 9274 9351
rect 7880 9181 7914 9215
rect 8016 9181 8050 9215
rect 8152 9181 8186 9215
rect 8288 9181 8322 9215
rect 8424 9181 8458 9215
rect 8560 9181 8594 9215
rect 8696 9181 8730 9215
rect 8832 9181 8866 9215
rect 8968 9181 9002 9215
rect 9104 9181 9138 9215
rect 9240 9181 9274 9215
rect 7880 9045 7914 9079
rect 8016 9045 8050 9079
rect 8152 9045 8186 9079
rect 8288 9045 8322 9079
rect 8424 9045 8458 9079
rect 8560 9045 8594 9079
rect 8696 9045 8730 9079
rect 8832 9045 8866 9079
rect 8968 9045 9002 9079
rect 9104 9045 9138 9079
rect 9240 9045 9274 9079
rect 7880 8909 7914 8943
rect 8016 8909 8050 8943
rect 8152 8909 8186 8943
rect 8288 8909 8322 8943
rect 8424 8909 8458 8943
rect 8560 8909 8594 8943
rect 8696 8909 8730 8943
rect 8832 8909 8866 8943
rect 8968 8909 9002 8943
rect 9104 8909 9138 8943
rect 9240 8909 9274 8943
rect 7880 8773 7914 8807
rect 8016 8773 8050 8807
rect 8152 8773 8186 8807
rect 8288 8773 8322 8807
rect 8424 8773 8458 8807
rect 8560 8773 8594 8807
rect 8696 8773 8730 8807
rect 8832 8773 8866 8807
rect 8968 8773 9002 8807
rect 9104 8773 9138 8807
rect 9240 8773 9274 8807
rect 7880 8637 7914 8671
rect 8016 8637 8050 8671
rect 8152 8637 8186 8671
rect 8288 8637 8322 8671
rect 8424 8637 8458 8671
rect 8560 8637 8594 8671
rect 8696 8637 8730 8671
rect 8832 8637 8866 8671
rect 8968 8637 9002 8671
rect 9104 8637 9138 8671
rect 9240 8637 9274 8671
rect 7880 8501 7914 8535
rect 8016 8501 8050 8535
rect 8152 8501 8186 8535
rect 8288 8501 8322 8535
rect 8424 8501 8458 8535
rect 8560 8501 8594 8535
rect 8696 8501 8730 8535
rect 8832 8501 8866 8535
rect 8968 8501 9002 8535
rect 9104 8501 9138 8535
rect 9240 8501 9274 8535
rect 7880 8365 7914 8399
rect 8016 8365 8050 8399
rect 8152 8365 8186 8399
rect 8288 8365 8322 8399
rect 8424 8365 8458 8399
rect 8560 8365 8594 8399
rect 8696 8365 8730 8399
rect 8832 8365 8866 8399
rect 8968 8365 9002 8399
rect 9104 8365 9138 8399
rect 9240 8365 9274 8399
rect 7880 8229 7914 8263
rect 8016 8229 8050 8263
rect 8152 8229 8186 8263
rect 8288 8229 8322 8263
rect 8424 8229 8458 8263
rect 8560 8229 8594 8263
rect 8696 8229 8730 8263
rect 8832 8229 8866 8263
rect 8968 8229 9002 8263
rect 9104 8229 9138 8263
rect 9240 8229 9274 8263
rect 7880 8093 7914 8127
rect 8016 8093 8050 8127
rect 8152 8093 8186 8127
rect 8288 8093 8322 8127
rect 8424 8093 8458 8127
rect 8560 8093 8594 8127
rect 8696 8093 8730 8127
rect 8832 8093 8866 8127
rect 8968 8093 9002 8127
rect 9104 8093 9138 8127
rect 9240 8093 9274 8127
rect 7880 7957 7914 7991
rect 8016 7957 8050 7991
rect 8152 7957 8186 7991
rect 8288 7957 8322 7991
rect 8424 7957 8458 7991
rect 8560 7957 8594 7991
rect 8696 7957 8730 7991
rect 8832 7957 8866 7991
rect 8968 7957 9002 7991
rect 9104 7957 9138 7991
rect 9240 7957 9274 7991
rect 7880 7821 7914 7855
rect 8016 7821 8050 7855
rect 8152 7821 8186 7855
rect 8288 7821 8322 7855
rect 8424 7821 8458 7855
rect 8560 7821 8594 7855
rect 8696 7821 8730 7855
rect 8832 7821 8866 7855
rect 8968 7821 9002 7855
rect 9104 7821 9138 7855
rect 9240 7821 9274 7855
rect 7880 7685 7914 7719
rect 8016 7685 8050 7719
rect 8152 7685 8186 7719
rect 8288 7685 8322 7719
rect 8424 7685 8458 7719
rect 8560 7685 8594 7719
rect 8696 7685 8730 7719
rect 8832 7685 8866 7719
rect 8968 7685 9002 7719
rect 9104 7685 9138 7719
rect 9240 7685 9274 7719
rect 7880 7549 7914 7583
rect 8016 7549 8050 7583
rect 8152 7549 8186 7583
rect 8288 7549 8322 7583
rect 8424 7549 8458 7583
rect 8560 7549 8594 7583
rect 8696 7549 8730 7583
rect 8832 7549 8866 7583
rect 8968 7549 9002 7583
rect 9104 7549 9138 7583
rect 9240 7549 9274 7583
rect 7880 7413 7914 7447
rect 8016 7413 8050 7447
rect 8152 7413 8186 7447
rect 8288 7413 8322 7447
rect 8424 7413 8458 7447
rect 8560 7413 8594 7447
rect 8696 7413 8730 7447
rect 8832 7413 8866 7447
rect 8968 7413 9002 7447
rect 9104 7413 9138 7447
rect 9240 7413 9274 7447
rect 7880 7277 7914 7311
rect 8016 7277 8050 7311
rect 8152 7277 8186 7311
rect 8288 7277 8322 7311
rect 8424 7277 8458 7311
rect 8560 7277 8594 7311
rect 8696 7277 8730 7311
rect 8832 7277 8866 7311
rect 8968 7277 9002 7311
rect 9104 7277 9138 7311
rect 9240 7277 9274 7311
rect 7880 7141 7914 7175
rect 8016 7141 8050 7175
rect 8152 7141 8186 7175
rect 8288 7141 8322 7175
rect 8424 7141 8458 7175
rect 8560 7141 8594 7175
rect 8696 7141 8730 7175
rect 8832 7141 8866 7175
rect 8968 7141 9002 7175
rect 9104 7141 9138 7175
rect 9240 7141 9274 7175
rect 7880 7005 7914 7039
rect 8016 7005 8050 7039
rect 8152 7005 8186 7039
rect 8288 7005 8322 7039
rect 8424 7005 8458 7039
rect 8560 7005 8594 7039
rect 8696 7005 8730 7039
rect 8832 7005 8866 7039
rect 8968 7005 9002 7039
rect 9104 7005 9138 7039
rect 9240 7005 9274 7039
rect 7880 6869 7914 6903
rect 8016 6869 8050 6903
rect 8152 6869 8186 6903
rect 8288 6869 8322 6903
rect 8424 6869 8458 6903
rect 8560 6869 8594 6903
rect 8696 6869 8730 6903
rect 8832 6869 8866 6903
rect 8968 6869 9002 6903
rect 9104 6869 9138 6903
rect 9240 6869 9274 6903
rect 7880 6733 7914 6767
rect 8016 6733 8050 6767
rect 8152 6733 8186 6767
rect 8288 6733 8322 6767
rect 8424 6733 8458 6767
rect 8560 6733 8594 6767
rect 8696 6733 8730 6767
rect 8832 6733 8866 6767
rect 8968 6733 9002 6767
rect 9104 6733 9138 6767
rect 9240 6733 9274 6767
rect 7880 6597 7914 6631
rect 8016 6597 8050 6631
rect 8152 6597 8186 6631
rect 8288 6597 8322 6631
rect 8424 6597 8458 6631
rect 8560 6597 8594 6631
rect 8696 6597 8730 6631
rect 8832 6597 8866 6631
rect 8968 6597 9002 6631
rect 9104 6597 9138 6631
rect 9240 6597 9274 6631
rect 7880 6461 7914 6495
rect 8016 6461 8050 6495
rect 8152 6461 8186 6495
rect 8288 6461 8322 6495
rect 8424 6461 8458 6495
rect 8560 6461 8594 6495
rect 8696 6461 8730 6495
rect 8832 6461 8866 6495
rect 8968 6461 9002 6495
rect 9104 6461 9138 6495
rect 9240 6461 9274 6495
rect 7880 6325 7914 6359
rect 8016 6325 8050 6359
rect 8152 6325 8186 6359
rect 8288 6325 8322 6359
rect 8424 6325 8458 6359
rect 8560 6325 8594 6359
rect 8696 6325 8730 6359
rect 8832 6325 8866 6359
rect 8968 6325 9002 6359
rect 9104 6325 9138 6359
rect 9240 6325 9274 6359
rect 7880 6189 7914 6223
rect 8016 6189 8050 6223
rect 8152 6189 8186 6223
rect 8288 6189 8322 6223
rect 8424 6189 8458 6223
rect 8560 6189 8594 6223
rect 8696 6189 8730 6223
rect 8832 6189 8866 6223
rect 8968 6189 9002 6223
rect 9104 6189 9138 6223
rect 9240 6189 9274 6223
rect 7880 6053 7914 6087
rect 8016 6053 8050 6087
rect 8152 6053 8186 6087
rect 8288 6053 8322 6087
rect 8424 6053 8458 6087
rect 8560 6053 8594 6087
rect 8696 6053 8730 6087
rect 8832 6053 8866 6087
rect 8968 6053 9002 6087
rect 9104 6053 9138 6087
rect 9240 6053 9274 6087
rect 7880 5917 7914 5951
rect 8016 5917 8050 5951
rect 8152 5917 8186 5951
rect 8288 5917 8322 5951
rect 8424 5917 8458 5951
rect 8560 5917 8594 5951
rect 8696 5917 8730 5951
rect 8832 5917 8866 5951
rect 8968 5917 9002 5951
rect 9104 5917 9138 5951
rect 9240 5917 9274 5951
rect 7880 5781 7914 5815
rect 8016 5781 8050 5815
rect 8152 5781 8186 5815
rect 8288 5781 8322 5815
rect 8424 5781 8458 5815
rect 8560 5781 8594 5815
rect 8696 5781 8730 5815
rect 8832 5781 8866 5815
rect 8968 5781 9002 5815
rect 9104 5781 9138 5815
rect 9240 5781 9274 5815
rect 7880 5645 7914 5679
rect 8016 5645 8050 5679
rect 8152 5645 8186 5679
rect 8288 5645 8322 5679
rect 8424 5645 8458 5679
rect 8560 5645 8594 5679
rect 8696 5645 8730 5679
rect 8832 5645 8866 5679
rect 8968 5645 9002 5679
rect 9104 5645 9138 5679
rect 9240 5645 9274 5679
rect 7880 5509 7914 5543
rect 8016 5509 8050 5543
rect 8152 5509 8186 5543
rect 8288 5509 8322 5543
rect 8424 5509 8458 5543
rect 8560 5509 8594 5543
rect 8696 5509 8730 5543
rect 8832 5509 8866 5543
rect 8968 5509 9002 5543
rect 9104 5509 9138 5543
rect 9240 5509 9274 5543
rect 7880 5373 7914 5407
rect 8016 5373 8050 5407
rect 8152 5373 8186 5407
rect 8288 5373 8322 5407
rect 8424 5373 8458 5407
rect 8560 5373 8594 5407
rect 8696 5373 8730 5407
rect 8832 5373 8866 5407
rect 8968 5373 9002 5407
rect 9104 5373 9138 5407
rect 9240 5373 9274 5407
rect 7880 5237 7914 5271
rect 8016 5237 8050 5271
rect 8152 5237 8186 5271
rect 8288 5237 8322 5271
rect 8424 5237 8458 5271
rect 8560 5237 8594 5271
rect 8696 5237 8730 5271
rect 8832 5237 8866 5271
rect 8968 5237 9002 5271
rect 9104 5237 9138 5271
rect 9240 5237 9274 5271
rect 7880 5101 7914 5135
rect 8016 5101 8050 5135
rect 8152 5101 8186 5135
rect 8288 5101 8322 5135
rect 8424 5101 8458 5135
rect 8560 5101 8594 5135
rect 8696 5101 8730 5135
rect 8832 5101 8866 5135
rect 8968 5101 9002 5135
rect 9104 5101 9138 5135
rect 9240 5101 9274 5135
rect 7880 4965 7914 4999
rect 8016 4965 8050 4999
rect 8152 4965 8186 4999
rect 8288 4965 8322 4999
rect 8424 4965 8458 4999
rect 8560 4965 8594 4999
rect 8696 4965 8730 4999
rect 8832 4965 8866 4999
rect 8968 4965 9002 4999
rect 9104 4965 9138 4999
rect 9240 4965 9274 4999
rect 7880 4829 7914 4863
rect 8016 4829 8050 4863
rect 8152 4829 8186 4863
rect 8288 4829 8322 4863
rect 8424 4829 8458 4863
rect 8560 4829 8594 4863
rect 8696 4829 8730 4863
rect 8832 4829 8866 4863
rect 8968 4829 9002 4863
rect 9104 4829 9138 4863
rect 9240 4829 9274 4863
rect 7880 4693 7914 4727
rect 8016 4693 8050 4727
rect 8152 4693 8186 4727
rect 8288 4693 8322 4727
rect 8424 4693 8458 4727
rect 8560 4693 8594 4727
rect 8696 4693 8730 4727
rect 8832 4693 8866 4727
rect 8968 4693 9002 4727
rect 9104 4693 9138 4727
rect 9240 4693 9274 4727
rect 7880 4557 7914 4591
rect 8016 4557 8050 4591
rect 8152 4557 8186 4591
rect 8288 4557 8322 4591
rect 8424 4557 8458 4591
rect 8560 4557 8594 4591
rect 8696 4557 8730 4591
rect 8832 4557 8866 4591
rect 8968 4557 9002 4591
rect 9104 4557 9138 4591
rect 9240 4557 9274 4591
rect 7880 4421 7914 4455
rect 8016 4421 8050 4455
rect 8152 4421 8186 4455
rect 8288 4421 8322 4455
rect 8424 4421 8458 4455
rect 8560 4421 8594 4455
rect 8696 4421 8730 4455
rect 8832 4421 8866 4455
rect 8968 4421 9002 4455
rect 9104 4421 9138 4455
rect 9240 4421 9274 4455
rect 7880 4285 7914 4319
rect 8016 4285 8050 4319
rect 8152 4285 8186 4319
rect 8288 4285 8322 4319
rect 8424 4285 8458 4319
rect 8560 4285 8594 4319
rect 8696 4285 8730 4319
rect 8832 4285 8866 4319
rect 8968 4285 9002 4319
rect 9104 4285 9138 4319
rect 9240 4285 9274 4319
rect 7880 4149 7914 4183
rect 8016 4149 8050 4183
rect 8152 4149 8186 4183
rect 8288 4149 8322 4183
rect 8424 4149 8458 4183
rect 8560 4149 8594 4183
rect 8696 4149 8730 4183
rect 8832 4149 8866 4183
rect 8968 4149 9002 4183
rect 9104 4149 9138 4183
rect 9240 4149 9274 4183
rect 7880 4013 7914 4047
rect 8016 4013 8050 4047
rect 8152 4013 8186 4047
rect 8288 4013 8322 4047
rect 8424 4013 8458 4047
rect 8560 4013 8594 4047
rect 8696 4013 8730 4047
rect 8832 4013 8866 4047
rect 8968 4013 9002 4047
rect 9104 4013 9138 4047
rect 9240 4013 9274 4047
rect 7880 3877 7914 3911
rect 8016 3877 8050 3911
rect 8152 3877 8186 3911
rect 8288 3877 8322 3911
rect 8424 3877 8458 3911
rect 8560 3877 8594 3911
rect 8696 3877 8730 3911
rect 8832 3877 8866 3911
rect 8968 3877 9002 3911
rect 9104 3877 9138 3911
rect 9240 3877 9274 3911
rect 7880 3741 7914 3775
rect 8016 3741 8050 3775
rect 8152 3741 8186 3775
rect 8288 3741 8322 3775
rect 8424 3741 8458 3775
rect 8560 3741 8594 3775
rect 8696 3741 8730 3775
rect 8832 3741 8866 3775
rect 8968 3741 9002 3775
rect 9104 3741 9138 3775
rect 9240 3741 9274 3775
rect 7880 3605 7914 3639
rect 8016 3605 8050 3639
rect 8152 3605 8186 3639
rect 8288 3605 8322 3639
rect 8424 3605 8458 3639
rect 8560 3605 8594 3639
rect 8696 3605 8730 3639
rect 8832 3605 8866 3639
rect 8968 3605 9002 3639
rect 9104 3605 9138 3639
rect 9240 3605 9274 3639
rect 7880 3469 7914 3503
rect 8016 3469 8050 3503
rect 8152 3469 8186 3503
rect 8288 3469 8322 3503
rect 8424 3469 8458 3503
rect 8560 3469 8594 3503
rect 8696 3469 8730 3503
rect 8832 3469 8866 3503
rect 8968 3469 9002 3503
rect 9104 3469 9138 3503
rect 9240 3469 9274 3503
rect 7880 3333 7914 3367
rect 8016 3333 8050 3367
rect 8152 3333 8186 3367
rect 8288 3333 8322 3367
rect 8424 3333 8458 3367
rect 8560 3333 8594 3367
rect 8696 3333 8730 3367
rect 8832 3333 8866 3367
rect 8968 3333 9002 3367
rect 9104 3333 9138 3367
rect 9240 3333 9274 3367
rect 7880 3197 7914 3231
rect 8016 3197 8050 3231
rect 8152 3197 8186 3231
rect 8288 3197 8322 3231
rect 8424 3197 8458 3231
rect 8560 3197 8594 3231
rect 8696 3197 8730 3231
rect 8832 3197 8866 3231
rect 8968 3197 9002 3231
rect 9104 3197 9138 3231
rect 9240 3197 9274 3231
rect 7880 3061 7914 3095
rect 8016 3061 8050 3095
rect 8152 3061 8186 3095
rect 8288 3061 8322 3095
rect 8424 3061 8458 3095
rect 8560 3061 8594 3095
rect 8696 3061 8730 3095
rect 8832 3061 8866 3095
rect 8968 3061 9002 3095
rect 9104 3061 9138 3095
rect 9240 3061 9274 3095
rect 7880 2925 7914 2959
rect 8016 2925 8050 2959
rect 8152 2925 8186 2959
rect 8288 2925 8322 2959
rect 8424 2925 8458 2959
rect 8560 2925 8594 2959
rect 8696 2925 8730 2959
rect 8832 2925 8866 2959
rect 8968 2925 9002 2959
rect 9104 2925 9138 2959
rect 9240 2925 9274 2959
rect 7880 2789 7914 2823
rect 8016 2789 8050 2823
rect 8152 2789 8186 2823
rect 8288 2789 8322 2823
rect 8424 2789 8458 2823
rect 8560 2789 8594 2823
rect 8696 2789 8730 2823
rect 8832 2789 8866 2823
rect 8968 2789 9002 2823
rect 9104 2789 9138 2823
rect 9240 2789 9274 2823
rect 7880 2653 7914 2687
rect 8016 2653 8050 2687
rect 8152 2653 8186 2687
rect 8288 2653 8322 2687
rect 8424 2653 8458 2687
rect 8560 2653 8594 2687
rect 8696 2653 8730 2687
rect 8832 2653 8866 2687
rect 8968 2653 9002 2687
rect 9104 2653 9138 2687
rect 9240 2653 9274 2687
rect 7880 2517 7914 2551
rect 8016 2517 8050 2551
rect 8152 2517 8186 2551
rect 8288 2517 8322 2551
rect 8424 2517 8458 2551
rect 8560 2517 8594 2551
rect 8696 2517 8730 2551
rect 8832 2517 8866 2551
rect 8968 2517 9002 2551
rect 9104 2517 9138 2551
rect 9240 2517 9274 2551
rect 7880 2380 7914 2414
rect 8016 2380 8050 2414
rect 8152 2380 8186 2414
rect 8288 2380 8322 2414
rect 8424 2380 8458 2414
rect 8560 2380 8594 2414
rect 8696 2380 8730 2414
rect 8832 2380 8866 2414
rect 8968 2380 9002 2414
rect 9104 2380 9138 2414
rect 9240 2380 9274 2414
rect 7880 2243 7914 2277
rect 8016 2243 8050 2277
rect 8152 2243 8186 2277
rect 8288 2243 8322 2277
rect 8424 2243 8458 2277
rect 8560 2243 8594 2277
rect 8696 2243 8730 2277
rect 8832 2243 8866 2277
rect 8968 2243 9002 2277
rect 9104 2243 9138 2277
rect 9240 2243 9274 2277
rect 7880 2106 7914 2140
rect 8016 2106 8050 2140
rect 8152 2106 8186 2140
rect 8288 2106 8322 2140
rect 8424 2106 8458 2140
rect 8560 2106 8594 2140
rect 8696 2106 8730 2140
rect 8832 2106 8866 2140
rect 8968 2106 9002 2140
rect 9104 2106 9138 2140
rect 9240 2106 9274 2140
rect 7880 1969 7914 2003
rect 8016 1969 8050 2003
rect 8152 1969 8186 2003
rect 8288 1969 8322 2003
rect 8424 1969 8458 2003
rect 8560 1969 8594 2003
rect 8696 1969 8730 2003
rect 8832 1969 8866 2003
rect 8968 1969 9002 2003
rect 9104 1969 9138 2003
rect 9240 1969 9274 2003
rect 7880 1832 7914 1866
rect 8016 1832 8050 1866
rect 8152 1832 8186 1866
rect 8288 1832 8322 1866
rect 8424 1832 8458 1866
rect 8560 1832 8594 1866
rect 8696 1832 8730 1866
rect 8832 1832 8866 1866
rect 8968 1832 9002 1866
rect 9104 1832 9138 1866
rect 9240 1832 9274 1866
rect 325 1695 359 1729
rect 461 1695 495 1729
rect 597 1695 631 1729
rect 733 1695 767 1729
rect 869 1695 903 1729
rect 1005 1695 1039 1729
rect 1141 1695 1175 1729
rect 1277 1695 1311 1729
rect 1413 1695 1447 1729
rect 1549 1695 1583 1729
rect 1685 1695 1719 1729
rect 325 1558 359 1592
rect 461 1558 495 1592
rect 597 1558 631 1592
rect 733 1558 767 1592
rect 869 1558 903 1592
rect 1005 1558 1039 1592
rect 1141 1558 1175 1592
rect 1277 1558 1311 1592
rect 1413 1558 1447 1592
rect 1549 1558 1583 1592
rect 1685 1558 1719 1592
rect 325 1421 359 1455
rect 461 1421 495 1455
rect 597 1421 631 1455
rect 733 1421 767 1455
rect 869 1421 903 1455
rect 1005 1421 1039 1455
rect 1141 1421 1175 1455
rect 1277 1421 1311 1455
rect 1413 1421 1447 1455
rect 1549 1421 1583 1455
rect 1685 1421 1719 1455
rect 325 1284 359 1318
rect 461 1284 495 1318
rect 597 1284 631 1318
rect 733 1284 767 1318
rect 869 1284 903 1318
rect 1005 1284 1039 1318
rect 1141 1284 1175 1318
rect 1277 1284 1311 1318
rect 1413 1284 1447 1318
rect 1549 1284 1583 1318
rect 1685 1284 1719 1318
rect 325 1147 359 1181
rect 461 1147 495 1181
rect 597 1147 631 1181
rect 733 1147 767 1181
rect 869 1147 903 1181
rect 1005 1147 1039 1181
rect 1141 1147 1175 1181
rect 1277 1147 1311 1181
rect 1413 1147 1447 1181
rect 1549 1147 1583 1181
rect 1685 1147 1719 1181
rect 325 1010 359 1044
rect 461 1010 495 1044
rect 597 1010 631 1044
rect 733 1010 767 1044
rect 869 1010 903 1044
rect 1005 1010 1039 1044
rect 1141 1010 1175 1044
rect 1277 1010 1311 1044
rect 1413 1010 1447 1044
rect 1549 1010 1583 1044
rect 1685 1010 1719 1044
rect 325 873 359 907
rect 461 873 495 907
rect 597 873 631 907
rect 733 873 767 907
rect 869 873 903 907
rect 1005 873 1039 907
rect 1141 873 1175 907
rect 1277 873 1311 907
rect 1413 873 1447 907
rect 1549 873 1583 907
rect 1685 873 1719 907
rect 325 736 359 770
rect 461 736 495 770
rect 597 736 631 770
rect 733 736 767 770
rect 869 736 903 770
rect 1005 736 1039 770
rect 1141 736 1175 770
rect 1277 736 1311 770
rect 1413 736 1447 770
rect 1549 736 1583 770
rect 1685 736 1719 770
rect 325 599 359 633
rect 461 599 495 633
rect 597 599 631 633
rect 733 599 767 633
rect 869 599 903 633
rect 1005 599 1039 633
rect 1141 599 1175 633
rect 1277 599 1311 633
rect 1413 599 1447 633
rect 1549 599 1583 633
rect 1685 599 1719 633
rect 325 462 359 496
rect 461 462 495 496
rect 597 462 631 496
rect 733 462 767 496
rect 869 462 903 496
rect 1005 462 1039 496
rect 1141 462 1175 496
rect 1277 462 1311 496
rect 1413 462 1447 496
rect 1549 462 1583 496
rect 1685 462 1719 496
rect 325 325 359 359
rect 461 325 495 359
rect 597 325 631 359
rect 733 325 767 359
rect 869 325 903 359
rect 1005 325 1039 359
rect 1141 325 1175 359
rect 1277 325 1311 359
rect 1413 325 1447 359
rect 1549 325 1583 359
rect 1685 325 1719 359
rect 325 188 359 222
rect 461 188 495 222
rect 597 188 631 222
rect 733 188 767 222
rect 869 188 903 222
rect 1005 188 1039 222
rect 1141 188 1175 222
rect 1277 188 1311 222
rect 1413 188 1447 222
rect 1549 188 1583 222
rect 1685 188 1719 222
rect 325 51 359 85
rect 461 51 495 85
rect 597 51 631 85
rect 733 51 767 85
rect 869 51 903 85
rect 1005 51 1039 85
rect 1141 51 1175 85
rect 1277 51 1311 85
rect 1413 51 1447 85
rect 1549 51 1583 85
rect 1685 51 1719 85
rect 7880 1695 7914 1729
rect 8016 1695 8050 1729
rect 8152 1695 8186 1729
rect 8288 1695 8322 1729
rect 8424 1695 8458 1729
rect 8560 1695 8594 1729
rect 8696 1695 8730 1729
rect 8832 1695 8866 1729
rect 8968 1695 9002 1729
rect 9104 1695 9138 1729
rect 9240 1695 9274 1729
rect 7880 1558 7914 1592
rect 8016 1558 8050 1592
rect 8152 1558 8186 1592
rect 8288 1558 8322 1592
rect 8424 1558 8458 1592
rect 8560 1558 8594 1592
rect 8696 1558 8730 1592
rect 8832 1558 8866 1592
rect 8968 1558 9002 1592
rect 9104 1558 9138 1592
rect 9240 1558 9274 1592
rect 7880 1421 7914 1455
rect 8016 1421 8050 1455
rect 8152 1421 8186 1455
rect 8288 1421 8322 1455
rect 8424 1421 8458 1455
rect 8560 1421 8594 1455
rect 8696 1421 8730 1455
rect 8832 1421 8866 1455
rect 8968 1421 9002 1455
rect 9104 1421 9138 1455
rect 9240 1421 9274 1455
rect 7880 1284 7914 1318
rect 8016 1284 8050 1318
rect 8152 1284 8186 1318
rect 8288 1284 8322 1318
rect 8424 1284 8458 1318
rect 8560 1284 8594 1318
rect 8696 1284 8730 1318
rect 8832 1284 8866 1318
rect 8968 1284 9002 1318
rect 9104 1284 9138 1318
rect 9240 1284 9274 1318
rect 7880 1147 7914 1181
rect 8016 1147 8050 1181
rect 8152 1147 8186 1181
rect 8288 1147 8322 1181
rect 8424 1147 8458 1181
rect 8560 1147 8594 1181
rect 8696 1147 8730 1181
rect 8832 1147 8866 1181
rect 8968 1147 9002 1181
rect 9104 1147 9138 1181
rect 9240 1147 9274 1181
rect 7880 1010 7914 1044
rect 8016 1010 8050 1044
rect 8152 1010 8186 1044
rect 8288 1010 8322 1044
rect 8424 1010 8458 1044
rect 8560 1010 8594 1044
rect 8696 1010 8730 1044
rect 8832 1010 8866 1044
rect 8968 1010 9002 1044
rect 9104 1010 9138 1044
rect 9240 1010 9274 1044
rect 7880 873 7914 907
rect 8016 873 8050 907
rect 8152 873 8186 907
rect 8288 873 8322 907
rect 8424 873 8458 907
rect 8560 873 8594 907
rect 8696 873 8730 907
rect 8832 873 8866 907
rect 8968 873 9002 907
rect 9104 873 9138 907
rect 9240 873 9274 907
rect 7880 736 7914 770
rect 8016 736 8050 770
rect 8152 736 8186 770
rect 8288 736 8322 770
rect 8424 736 8458 770
rect 8560 736 8594 770
rect 8696 736 8730 770
rect 8832 736 8866 770
rect 8968 736 9002 770
rect 9104 736 9138 770
rect 9240 736 9274 770
rect 7880 599 7914 633
rect 8016 599 8050 633
rect 8152 599 8186 633
rect 8288 599 8322 633
rect 8424 599 8458 633
rect 8560 599 8594 633
rect 8696 599 8730 633
rect 8832 599 8866 633
rect 8968 599 9002 633
rect 9104 599 9138 633
rect 9240 599 9274 633
rect 7880 462 7914 496
rect 8016 462 8050 496
rect 8152 462 8186 496
rect 8288 462 8322 496
rect 8424 462 8458 496
rect 8560 462 8594 496
rect 8696 462 8730 496
rect 8832 462 8866 496
rect 8968 462 9002 496
rect 9104 462 9138 496
rect 9240 462 9274 496
rect 7880 325 7914 359
rect 8016 325 8050 359
rect 8152 325 8186 359
rect 8288 325 8322 359
rect 8424 325 8458 359
rect 8560 325 8594 359
rect 8696 325 8730 359
rect 8832 325 8866 359
rect 8968 325 9002 359
rect 9104 325 9138 359
rect 9240 325 9274 359
rect 7880 188 7914 222
rect 8016 188 8050 222
rect 8152 188 8186 222
rect 8288 188 8322 222
rect 8424 188 8458 222
rect 8560 188 8594 222
rect 8696 188 8730 222
rect 8832 188 8866 222
rect 8968 188 9002 222
rect 9104 188 9138 222
rect 9240 188 9274 222
rect 7880 51 7914 85
rect 8016 51 8050 85
rect 8152 51 8186 85
rect 8288 51 8322 85
rect 8424 51 8458 85
rect 8560 51 8594 85
rect 8696 51 8730 85
rect 8832 51 8866 85
rect 8968 51 9002 85
rect 9104 51 9138 85
rect 9240 51 9274 85
<< mvnsubdiffcont >>
rect 5139 16438 5173 16472
rect 5207 16438 5241 16472
rect 5275 16438 5309 16472
rect 5343 16438 5377 16472
rect 5411 16438 5445 16472
rect 5479 16438 5513 16472
rect 5547 16438 5581 16472
rect 5615 16438 5649 16472
rect 5683 16438 5717 16472
rect 5751 16438 5785 16472
rect 5819 16438 5853 16472
rect 5887 16438 5921 16472
rect 5955 16438 5989 16472
rect 6023 16438 6057 16472
rect 6091 16438 6125 16472
rect 6159 16438 6193 16472
rect 6227 16438 6261 16472
rect 6295 16438 6329 16472
rect 6363 16438 6397 16472
rect 6431 16438 6465 16472
rect 6499 16438 6533 16472
rect 6567 16438 6601 16472
rect 6635 16438 6669 16472
rect 6703 16438 6737 16472
rect 6771 16438 6805 16472
rect 6839 16438 6873 16472
rect 6907 16438 6941 16472
rect 6975 16438 7009 16472
rect 7043 16438 7077 16472
rect 7111 16438 7145 16472
rect 7179 16438 7213 16472
rect 7247 16438 7281 16472
rect 7315 16438 7349 16472
rect 7383 16438 7417 16472
rect 7451 16438 7485 16472
rect 5004 16370 5038 16404
rect 5004 16302 5038 16336
rect 5004 16234 5038 16268
rect 5004 16166 5038 16200
rect 5004 16098 5038 16132
rect 5004 16030 5038 16064
rect 5004 15962 5038 15996
rect 5004 15894 5038 15928
rect 5004 15826 5038 15860
rect 5004 15758 5038 15792
rect 5004 15690 5038 15724
rect 5004 15622 5038 15656
rect 5004 15554 5038 15588
rect 5004 15486 5038 15520
rect 5004 15418 5038 15452
rect 5004 15350 5038 15384
rect 5004 15282 5038 15316
rect 5004 15214 5038 15248
rect 5004 15146 5038 15180
rect 5004 15078 5038 15112
rect 5004 15010 5038 15044
rect 5004 14942 5038 14976
rect 5004 14874 5038 14908
rect 5004 14806 5038 14840
rect 5004 14738 5038 14772
rect 5004 14670 5038 14704
rect 5004 14602 5038 14636
rect 5004 14534 5038 14568
rect 5004 14466 5038 14500
rect 5004 14398 5038 14432
rect 5004 14330 5038 14364
rect 5004 14262 5038 14296
rect 5004 14194 5038 14228
rect 5004 14126 5038 14160
rect 5004 14058 5038 14092
rect 5004 13990 5038 14024
rect 5004 13922 5038 13956
rect 5004 13854 5038 13888
rect 5004 13786 5038 13820
rect 5004 13718 5038 13752
rect 5004 13650 5038 13684
rect 5004 13582 5038 13616
rect 5004 13514 5038 13548
rect 5004 13446 5038 13480
rect 5004 13378 5038 13412
rect 5004 13310 5038 13344
rect 5004 13242 5038 13276
rect 5004 13174 5038 13208
rect 5004 13106 5038 13140
rect 5004 13038 5038 13072
rect 5004 12970 5038 13004
rect 5004 12902 5038 12936
rect 5004 12834 5038 12868
rect 5004 12766 5038 12800
rect 5004 12698 5038 12732
rect 5004 12630 5038 12664
rect 5004 12562 5038 12596
rect 5004 12494 5038 12528
rect 5004 12426 5038 12460
rect 5004 12358 5038 12392
rect 5004 12290 5038 12324
rect 5004 12222 5038 12256
rect 5004 12154 5038 12188
rect 5004 12086 5038 12120
rect 5004 12018 5038 12052
rect 5004 11950 5038 11984
rect 5004 11882 5038 11916
rect 5004 11814 5038 11848
rect 5004 11746 5038 11780
rect 5004 11678 5038 11712
rect 5004 11610 5038 11644
rect 5004 11542 5038 11576
rect 5004 11474 5038 11508
rect 5004 11406 5038 11440
rect 5004 11338 5038 11372
rect 5004 11270 5038 11304
rect 5004 11202 5038 11236
rect 5004 11134 5038 11168
rect 5004 11066 5038 11100
rect 5004 10998 5038 11032
rect 5004 10930 5038 10964
rect 5004 10862 5038 10896
rect 5004 10794 5038 10828
rect 5004 10726 5038 10760
rect 5004 10658 5038 10692
rect 5004 10590 5038 10624
rect 5004 10522 5038 10556
rect 5004 10454 5038 10488
rect 5004 10386 5038 10420
rect 5004 10318 5038 10352
rect 5004 10250 5038 10284
rect 5004 10182 5038 10216
rect 5004 10114 5038 10148
rect 5004 10046 5038 10080
rect 5004 9978 5038 10012
rect 5004 9910 5038 9944
rect 5004 9842 5038 9876
rect 5004 9774 5038 9808
rect 5004 9706 5038 9740
rect 5004 9638 5038 9672
rect 5004 9570 5038 9604
rect 5004 9502 5038 9536
rect 5004 9434 5038 9468
rect 5004 9366 5038 9400
rect 5004 9298 5038 9332
rect 5004 9230 5038 9264
rect 5004 9162 5038 9196
rect 5004 9094 5038 9128
rect 5004 9026 5038 9060
rect 5004 8958 5038 8992
rect 5004 8890 5038 8924
rect 5004 8822 5038 8856
rect 5004 8754 5038 8788
rect 5004 8686 5038 8720
rect 5004 8618 5038 8652
rect 5004 8550 5038 8584
rect 5004 8482 5038 8516
rect 5004 8414 5038 8448
rect 5004 8346 5038 8380
rect 5004 8278 5038 8312
rect 5004 8210 5038 8244
rect 5004 8142 5038 8176
rect 5004 8074 5038 8108
rect 5004 8006 5038 8040
rect 5004 7938 5038 7972
rect 5004 7870 5038 7904
rect 5004 7802 5038 7836
rect 5004 7734 5038 7768
rect 5004 7666 5038 7700
rect 5004 7598 5038 7632
rect 5004 7530 5038 7564
rect 5004 7462 5038 7496
rect 5004 7394 5038 7428
rect 5004 7326 5038 7360
rect 5004 7258 5038 7292
rect 5004 7190 5038 7224
rect 5004 7122 5038 7156
rect 5004 7054 5038 7088
rect 5004 6986 5038 7020
rect 5004 6918 5038 6952
rect 5004 6850 5038 6884
rect 5004 6782 5038 6816
rect 5004 6714 5038 6748
rect 5004 6646 5038 6680
rect 5004 6578 5038 6612
rect 5004 6510 5038 6544
rect 5004 6442 5038 6476
rect 5004 6374 5038 6408
rect 5004 6306 5038 6340
rect 5004 6238 5038 6272
rect 5004 6170 5038 6204
rect 5004 6102 5038 6136
rect 5004 6034 5038 6068
rect 5004 5966 5038 6000
rect 5004 5898 5038 5932
rect 5004 5830 5038 5864
rect 5004 5762 5038 5796
rect 5004 5694 5038 5728
rect 5004 5626 5038 5660
rect 5004 5558 5038 5592
rect 5004 5490 5038 5524
rect 5004 5422 5038 5456
rect 5004 5354 5038 5388
rect 5004 5286 5038 5320
rect 5004 5218 5038 5252
rect 5004 5150 5038 5184
rect 5004 5082 5038 5116
rect 5004 5014 5038 5048
rect 5004 4946 5038 4980
rect 5004 4878 5038 4912
rect 5004 4810 5038 4844
rect 5004 4742 5038 4776
rect 5004 4674 5038 4708
rect 5004 4606 5038 4640
rect 5004 4538 5038 4572
rect 5004 4470 5038 4504
rect 5004 4402 5038 4436
rect 5004 4334 5038 4368
rect 5004 4266 5038 4300
rect 5004 4198 5038 4232
rect 5004 4130 5038 4164
rect 5004 4062 5038 4096
rect 5004 3994 5038 4028
rect 5004 3926 5038 3960
rect 5004 3858 5038 3892
rect 5004 3790 5038 3824
rect 5004 3722 5038 3756
rect 5004 3654 5038 3688
rect 5004 3586 5038 3620
rect 5004 3518 5038 3552
rect 5004 3450 5038 3484
rect 5004 3382 5038 3416
rect 5004 3314 5038 3348
rect 5004 3246 5038 3280
rect 5004 3178 5038 3212
rect 5004 3110 5038 3144
rect 5004 3042 5038 3076
rect 5004 2974 5038 3008
rect 5004 2906 5038 2940
rect 5004 2838 5038 2872
rect 5004 2770 5038 2804
rect 5004 2702 5038 2736
rect 5004 2634 5038 2668
rect 5004 2566 5038 2600
rect 5004 2498 5038 2532
rect 5004 2430 5038 2464
rect 5004 2362 5038 2396
rect 5004 2294 5038 2328
rect 5004 2226 5038 2260
rect 5004 2158 5038 2192
rect 5004 2090 5038 2124
rect 5004 2022 5038 2056
rect 5004 1954 5038 1988
rect 5004 1821 5038 1855
rect 7519 16349 7553 16383
rect 7519 16281 7553 16315
rect 7519 16213 7553 16247
rect 7519 16145 7553 16179
rect 7519 16077 7553 16111
rect 7519 16009 7553 16043
rect 7519 15941 7553 15975
rect 7519 15873 7553 15907
rect 7519 15805 7553 15839
rect 7519 15737 7553 15771
rect 7519 15669 7553 15703
rect 7519 15601 7553 15635
rect 7519 15533 7553 15567
rect 7519 15465 7553 15499
rect 7519 15397 7553 15431
rect 7519 15329 7553 15363
rect 7519 15261 7553 15295
rect 7519 15193 7553 15227
rect 7519 15125 7553 15159
rect 7519 15057 7553 15091
rect 7519 14989 7553 15023
rect 7519 14921 7553 14955
rect 7519 14853 7553 14887
rect 7519 14785 7553 14819
rect 7519 14717 7553 14751
rect 7519 14649 7553 14683
rect 7519 14581 7553 14615
rect 7519 14513 7553 14547
rect 7519 14445 7553 14479
rect 7519 14377 7553 14411
rect 7519 14309 7553 14343
rect 7519 14241 7553 14275
rect 7519 14173 7553 14207
rect 7519 14105 7553 14139
rect 7519 14037 7553 14071
rect 7519 13969 7553 14003
rect 7519 13901 7553 13935
rect 7519 13833 7553 13867
rect 7519 13765 7553 13799
rect 7519 13697 7553 13731
rect 7519 13629 7553 13663
rect 7519 13561 7553 13595
rect 7519 13493 7553 13527
rect 7519 13425 7553 13459
rect 7519 13357 7553 13391
rect 7519 13289 7553 13323
rect 7519 13221 7553 13255
rect 7519 13153 7553 13187
rect 7519 13085 7553 13119
rect 7519 13017 7553 13051
rect 7519 12949 7553 12983
rect 7519 12881 7553 12915
rect 7519 12813 7553 12847
rect 7519 12745 7553 12779
rect 7519 12677 7553 12711
rect 7519 12609 7553 12643
rect 7519 12541 7553 12575
rect 7519 12473 7553 12507
rect 7519 12405 7553 12439
rect 7519 12337 7553 12371
rect 7519 12269 7553 12303
rect 7519 12201 7553 12235
rect 7519 12133 7553 12167
rect 7519 12065 7553 12099
rect 7519 11997 7553 12031
rect 7519 11929 7553 11963
rect 7519 11861 7553 11895
rect 7519 11793 7553 11827
rect 7519 11725 7553 11759
rect 7519 11657 7553 11691
rect 7519 11589 7553 11623
rect 7519 11521 7553 11555
rect 7519 11453 7553 11487
rect 7519 11385 7553 11419
rect 7519 11317 7553 11351
rect 7519 11249 7553 11283
rect 7519 11181 7553 11215
rect 7519 11113 7553 11147
rect 7519 11045 7553 11079
rect 7519 10977 7553 11011
rect 7519 10909 7553 10943
rect 7519 10841 7553 10875
rect 7519 10773 7553 10807
rect 7519 10705 7553 10739
rect 7519 10637 7553 10671
rect 7519 10569 7553 10603
rect 7519 10501 7553 10535
rect 7519 10433 7553 10467
rect 7519 10365 7553 10399
rect 7519 10297 7553 10331
rect 7519 10229 7553 10263
rect 7519 10161 7553 10195
rect 7519 10093 7553 10127
rect 7519 10025 7553 10059
rect 7519 9957 7553 9991
rect 7519 9889 7553 9923
rect 7519 9821 7553 9855
rect 7519 9753 7553 9787
rect 7519 9685 7553 9719
rect 7519 9617 7553 9651
rect 7519 9549 7553 9583
rect 7519 9481 7553 9515
rect 7519 9413 7553 9447
rect 7519 9345 7553 9379
rect 7519 9277 7553 9311
rect 7519 9209 7553 9243
rect 7519 9141 7553 9175
rect 7519 9073 7553 9107
rect 7519 9005 7553 9039
rect 7519 8937 7553 8971
rect 7519 8869 7553 8903
rect 7519 8801 7553 8835
rect 7519 8733 7553 8767
rect 7519 8665 7553 8699
rect 7519 8597 7553 8631
rect 7519 8529 7553 8563
rect 7519 8461 7553 8495
rect 7519 8393 7553 8427
rect 7519 8325 7553 8359
rect 7519 8257 7553 8291
rect 7519 8189 7553 8223
rect 7519 8121 7553 8155
rect 7519 8053 7553 8087
rect 7519 7985 7553 8019
rect 7519 7917 7553 7951
rect 7519 7849 7553 7883
rect 7519 7781 7553 7815
rect 7519 7713 7553 7747
rect 7519 7645 7553 7679
rect 7519 7577 7553 7611
rect 7519 7509 7553 7543
rect 7519 7441 7553 7475
rect 7519 7373 7553 7407
rect 7519 7305 7553 7339
rect 7519 7237 7553 7271
rect 7519 7169 7553 7203
rect 7519 7101 7553 7135
rect 7519 7033 7553 7067
rect 7519 6965 7553 6999
rect 7519 6897 7553 6931
rect 7519 6829 7553 6863
rect 7519 6761 7553 6795
rect 7519 6693 7553 6727
rect 7519 6625 7553 6659
rect 7519 6557 7553 6591
rect 7519 6489 7553 6523
rect 7519 6421 7553 6455
rect 7519 6353 7553 6387
rect 7519 6285 7553 6319
rect 7519 6217 7553 6251
rect 7519 6149 7553 6183
rect 7519 6081 7553 6115
rect 7519 6013 7553 6047
rect 7519 5945 7553 5979
rect 7519 5877 7553 5911
rect 7519 5809 7553 5843
rect 7519 5741 7553 5775
rect 7519 5673 7553 5707
rect 7519 5605 7553 5639
rect 7519 5537 7553 5571
rect 7519 5469 7553 5503
rect 7519 5401 7553 5435
rect 7519 5333 7553 5367
rect 7519 5265 7553 5299
rect 7519 5197 7553 5231
rect 7519 5129 7553 5163
rect 7519 5061 7553 5095
rect 7519 4993 7553 5027
rect 7519 4925 7553 4959
rect 7519 4857 7553 4891
rect 7519 4789 7553 4823
rect 7519 4721 7553 4755
rect 7519 4653 7553 4687
rect 7519 4585 7553 4619
rect 7519 4517 7553 4551
rect 7519 4449 7553 4483
rect 7519 4381 7553 4415
rect 7519 4313 7553 4347
rect 7519 4245 7553 4279
rect 7519 4177 7553 4211
rect 7519 4109 7553 4143
rect 7519 4041 7553 4075
rect 7519 3973 7553 4007
rect 7519 3905 7553 3939
rect 7519 3837 7553 3871
rect 7519 3769 7553 3803
rect 7519 3701 7553 3735
rect 7519 3633 7553 3667
rect 7519 3565 7553 3599
rect 7519 3497 7553 3531
rect 7519 3429 7553 3463
rect 7519 3361 7553 3395
rect 7519 3293 7553 3327
rect 7519 3225 7553 3259
rect 7519 3157 7553 3191
rect 7519 3089 7553 3123
rect 7519 3021 7553 3055
rect 7519 2953 7553 2987
rect 7519 2885 7553 2919
rect 7519 2817 7553 2851
rect 7519 2749 7553 2783
rect 7519 2681 7553 2715
rect 7519 2613 7553 2647
rect 7519 2545 7553 2579
rect 7519 2477 7553 2511
rect 7519 2409 7553 2443
rect 7519 2341 7553 2375
rect 7519 2273 7553 2307
rect 7519 2205 7553 2239
rect 7519 2137 7553 2171
rect 7519 2069 7553 2103
rect 7519 2001 7553 2035
rect 7519 1933 7553 1967
rect 7519 1865 7553 1899
rect 7519 1797 7553 1831
rect 5072 1729 5106 1763
rect 5140 1729 5174 1763
rect 5208 1729 5242 1763
rect 5276 1729 5310 1763
rect 5344 1729 5378 1763
rect 5412 1729 5446 1763
rect 5480 1729 5514 1763
rect 5548 1729 5582 1763
rect 5616 1729 5650 1763
rect 5684 1729 5718 1763
rect 5752 1729 5786 1763
rect 5820 1729 5854 1763
rect 5888 1729 5922 1763
rect 5956 1729 5990 1763
rect 6024 1729 6058 1763
rect 6092 1729 6126 1763
rect 6160 1729 6194 1763
rect 6228 1729 6262 1763
rect 6296 1729 6330 1763
rect 6364 1729 6398 1763
rect 6432 1729 6466 1763
rect 6500 1729 6534 1763
rect 6568 1729 6602 1763
rect 6636 1729 6670 1763
rect 6704 1729 6738 1763
rect 6772 1729 6806 1763
rect 6840 1729 6874 1763
rect 6908 1729 6942 1763
rect 6976 1729 7010 1763
rect 7044 1729 7078 1763
rect 7112 1729 7146 1763
rect 7180 1729 7214 1763
rect 7248 1729 7282 1763
rect 7316 1729 7350 1763
rect 7384 1729 7418 1763
<< locali >>
rect 315 39951 1729 39975
rect 315 39943 325 39951
rect 359 39943 461 39951
rect 495 39943 597 39951
rect 631 39943 733 39951
rect 767 39943 869 39951
rect 903 39943 1005 39951
rect 1039 39943 1141 39951
rect 1175 39943 1277 39951
rect 1311 39943 1413 39951
rect 1447 39943 1549 39951
rect 1583 39943 1685 39951
rect 1719 39943 1729 39951
rect 315 33357 321 39943
rect 1723 33357 1729 39943
rect 315 33318 1729 33357
rect 315 33284 321 33318
rect 355 33287 393 33318
rect 359 33284 393 33287
rect 427 33287 465 33318
rect 427 33284 461 33287
rect 499 33284 537 33318
rect 571 33287 609 33318
rect 571 33284 597 33287
rect 643 33284 681 33318
rect 715 33287 753 33318
rect 715 33284 733 33287
rect 787 33284 825 33318
rect 859 33287 897 33318
rect 859 33284 869 33287
rect 931 33284 969 33318
rect 1003 33287 1041 33318
rect 1003 33284 1005 33287
rect 315 33253 325 33284
rect 359 33253 461 33284
rect 495 33253 597 33284
rect 631 33253 733 33284
rect 767 33253 869 33284
rect 903 33253 1005 33284
rect 1039 33284 1041 33287
rect 1075 33284 1113 33318
rect 1147 33287 1185 33318
rect 1175 33284 1185 33287
rect 1219 33284 1257 33318
rect 1291 33287 1329 33318
rect 1311 33284 1329 33287
rect 1363 33284 1401 33318
rect 1435 33287 1473 33318
rect 1447 33284 1473 33287
rect 1507 33284 1545 33318
rect 1579 33287 1617 33318
rect 1583 33284 1617 33287
rect 1651 33287 1689 33318
rect 1651 33284 1685 33287
rect 1723 33284 1729 33318
rect 1039 33253 1141 33284
rect 1175 33253 1277 33284
rect 1311 33253 1413 33284
rect 1447 33253 1549 33284
rect 1583 33253 1685 33284
rect 1719 33253 1729 33284
rect 315 33245 1729 33253
rect 315 33211 321 33245
rect 355 33211 393 33245
rect 427 33211 465 33245
rect 499 33211 537 33245
rect 571 33211 609 33245
rect 643 33211 681 33245
rect 715 33211 753 33245
rect 787 33211 825 33245
rect 859 33211 897 33245
rect 931 33211 969 33245
rect 1003 33211 1041 33245
rect 1075 33211 1113 33245
rect 1147 33211 1185 33245
rect 1219 33211 1257 33245
rect 1291 33211 1329 33245
rect 1363 33211 1401 33245
rect 1435 33211 1473 33245
rect 1507 33211 1545 33245
rect 1579 33211 1617 33245
rect 1651 33211 1689 33245
rect 1723 33211 1729 33245
rect 315 33172 1729 33211
rect 315 33138 321 33172
rect 355 33151 393 33172
rect 359 33138 393 33151
rect 427 33151 465 33172
rect 427 33138 461 33151
rect 499 33138 537 33172
rect 571 33151 609 33172
rect 571 33138 597 33151
rect 643 33138 681 33172
rect 715 33151 753 33172
rect 715 33138 733 33151
rect 787 33138 825 33172
rect 859 33151 897 33172
rect 859 33138 869 33151
rect 931 33138 969 33172
rect 1003 33151 1041 33172
rect 1003 33138 1005 33151
rect 315 33117 325 33138
rect 359 33117 461 33138
rect 495 33117 597 33138
rect 631 33117 733 33138
rect 767 33117 869 33138
rect 903 33117 1005 33138
rect 1039 33138 1041 33151
rect 1075 33138 1113 33172
rect 1147 33151 1185 33172
rect 1175 33138 1185 33151
rect 1219 33138 1257 33172
rect 1291 33151 1329 33172
rect 1311 33138 1329 33151
rect 1363 33138 1401 33172
rect 1435 33151 1473 33172
rect 1447 33138 1473 33151
rect 1507 33138 1545 33172
rect 1579 33151 1617 33172
rect 1583 33138 1617 33151
rect 1651 33151 1689 33172
rect 1651 33138 1685 33151
rect 1723 33138 1729 33172
rect 1039 33117 1141 33138
rect 1175 33117 1277 33138
rect 1311 33117 1413 33138
rect 1447 33117 1549 33138
rect 1583 33117 1685 33138
rect 1719 33117 1729 33138
rect 315 33099 1729 33117
rect 315 33065 321 33099
rect 355 33065 393 33099
rect 427 33065 465 33099
rect 499 33065 537 33099
rect 571 33065 609 33099
rect 643 33065 681 33099
rect 715 33065 753 33099
rect 787 33065 825 33099
rect 859 33065 897 33099
rect 931 33065 969 33099
rect 1003 33065 1041 33099
rect 1075 33065 1113 33099
rect 1147 33065 1185 33099
rect 1219 33065 1257 33099
rect 1291 33065 1329 33099
rect 1363 33065 1401 33099
rect 1435 33065 1473 33099
rect 1507 33065 1545 33099
rect 1579 33065 1617 33099
rect 1651 33065 1689 33099
rect 1723 33065 1729 33099
rect 315 33026 1729 33065
rect 315 32992 321 33026
rect 355 33015 393 33026
rect 359 32992 393 33015
rect 427 33015 465 33026
rect 427 32992 461 33015
rect 499 32992 537 33026
rect 571 33015 609 33026
rect 571 32992 597 33015
rect 643 32992 681 33026
rect 715 33015 753 33026
rect 715 32992 733 33015
rect 787 32992 825 33026
rect 859 33015 897 33026
rect 859 32992 869 33015
rect 931 32992 969 33026
rect 1003 33015 1041 33026
rect 1003 32992 1005 33015
rect 315 32981 325 32992
rect 359 32981 461 32992
rect 495 32981 597 32992
rect 631 32981 733 32992
rect 767 32981 869 32992
rect 903 32981 1005 32992
rect 1039 32992 1041 33015
rect 1075 32992 1113 33026
rect 1147 33015 1185 33026
rect 1175 32992 1185 33015
rect 1219 32992 1257 33026
rect 1291 33015 1329 33026
rect 1311 32992 1329 33015
rect 1363 32992 1401 33026
rect 1435 33015 1473 33026
rect 1447 32992 1473 33015
rect 1507 32992 1545 33026
rect 1579 33015 1617 33026
rect 1583 32992 1617 33015
rect 1651 33015 1689 33026
rect 1651 32992 1685 33015
rect 1723 32992 1729 33026
rect 1039 32981 1141 32992
rect 1175 32981 1277 32992
rect 1311 32981 1413 32992
rect 1447 32981 1549 32992
rect 1583 32981 1685 32992
rect 1719 32981 1729 32992
rect 315 32953 1729 32981
rect 315 32919 321 32953
rect 355 32919 393 32953
rect 427 32919 465 32953
rect 499 32919 537 32953
rect 571 32919 609 32953
rect 643 32919 681 32953
rect 715 32919 753 32953
rect 787 32919 825 32953
rect 859 32919 897 32953
rect 931 32919 969 32953
rect 1003 32919 1041 32953
rect 1075 32919 1113 32953
rect 1147 32919 1185 32953
rect 1219 32919 1257 32953
rect 1291 32919 1329 32953
rect 1363 32919 1401 32953
rect 1435 32919 1473 32953
rect 1507 32919 1545 32953
rect 1579 32919 1617 32953
rect 1651 32919 1689 32953
rect 1723 32919 1729 32953
rect 315 32880 1729 32919
rect 315 32846 321 32880
rect 355 32879 393 32880
rect 359 32846 393 32879
rect 427 32879 465 32880
rect 427 32846 461 32879
rect 499 32846 537 32880
rect 571 32879 609 32880
rect 571 32846 597 32879
rect 643 32846 681 32880
rect 715 32879 753 32880
rect 715 32846 733 32879
rect 787 32846 825 32880
rect 859 32879 897 32880
rect 859 32846 869 32879
rect 931 32846 969 32880
rect 1003 32879 1041 32880
rect 1003 32846 1005 32879
rect 315 32845 325 32846
rect 359 32845 461 32846
rect 495 32845 597 32846
rect 631 32845 733 32846
rect 767 32845 869 32846
rect 903 32845 1005 32846
rect 1039 32846 1041 32879
rect 1075 32846 1113 32880
rect 1147 32879 1185 32880
rect 1175 32846 1185 32879
rect 1219 32846 1257 32880
rect 1291 32879 1329 32880
rect 1311 32846 1329 32879
rect 1363 32846 1401 32880
rect 1435 32879 1473 32880
rect 1447 32846 1473 32879
rect 1507 32846 1545 32880
rect 1579 32879 1617 32880
rect 1583 32846 1617 32879
rect 1651 32879 1689 32880
rect 1651 32846 1685 32879
rect 1723 32846 1729 32880
rect 1039 32845 1141 32846
rect 1175 32845 1277 32846
rect 1311 32845 1413 32846
rect 1447 32845 1549 32846
rect 1583 32845 1685 32846
rect 1719 32845 1729 32846
rect 315 32807 1729 32845
rect 315 32773 321 32807
rect 355 32773 393 32807
rect 427 32773 465 32807
rect 499 32773 537 32807
rect 571 32773 609 32807
rect 643 32773 681 32807
rect 715 32773 753 32807
rect 787 32773 825 32807
rect 859 32773 897 32807
rect 931 32773 969 32807
rect 1003 32773 1041 32807
rect 1075 32773 1113 32807
rect 1147 32773 1185 32807
rect 1219 32773 1257 32807
rect 1291 32773 1329 32807
rect 1363 32773 1401 32807
rect 1435 32773 1473 32807
rect 1507 32773 1545 32807
rect 1579 32773 1617 32807
rect 1651 32773 1689 32807
rect 1723 32773 1729 32807
rect 315 32743 1729 32773
rect 315 32734 325 32743
rect 359 32734 461 32743
rect 495 32734 597 32743
rect 631 32734 733 32743
rect 767 32734 869 32743
rect 903 32734 1005 32743
rect 315 32700 321 32734
rect 359 32709 393 32734
rect 355 32700 393 32709
rect 427 32709 461 32734
rect 427 32700 465 32709
rect 499 32700 537 32734
rect 571 32709 597 32734
rect 571 32700 609 32709
rect 643 32700 681 32734
rect 715 32709 733 32734
rect 715 32700 753 32709
rect 787 32700 825 32734
rect 859 32709 869 32734
rect 859 32700 897 32709
rect 931 32700 969 32734
rect 1003 32709 1005 32734
rect 1039 32734 1141 32743
rect 1175 32734 1277 32743
rect 1311 32734 1413 32743
rect 1447 32734 1549 32743
rect 1583 32734 1685 32743
rect 1719 32734 1729 32743
rect 1039 32709 1041 32734
rect 1003 32700 1041 32709
rect 1075 32700 1113 32734
rect 1175 32709 1185 32734
rect 1147 32700 1185 32709
rect 1219 32700 1257 32734
rect 1311 32709 1329 32734
rect 1291 32700 1329 32709
rect 1363 32700 1401 32734
rect 1447 32709 1473 32734
rect 1435 32700 1473 32709
rect 1507 32700 1545 32734
rect 1583 32709 1617 32734
rect 1579 32700 1617 32709
rect 1651 32709 1685 32734
rect 1651 32700 1689 32709
rect 1723 32700 1729 32734
rect 315 32661 1729 32700
rect 315 32627 321 32661
rect 355 32627 393 32661
rect 427 32627 465 32661
rect 499 32627 537 32661
rect 571 32627 609 32661
rect 643 32627 681 32661
rect 715 32627 753 32661
rect 787 32627 825 32661
rect 859 32627 897 32661
rect 931 32627 969 32661
rect 1003 32627 1041 32661
rect 1075 32627 1113 32661
rect 1147 32627 1185 32661
rect 1219 32627 1257 32661
rect 1291 32627 1329 32661
rect 1363 32627 1401 32661
rect 1435 32627 1473 32661
rect 1507 32627 1545 32661
rect 1579 32627 1617 32661
rect 1651 32627 1689 32661
rect 1723 32627 1729 32661
rect 315 32607 1729 32627
rect 315 32588 325 32607
rect 359 32588 461 32607
rect 495 32588 597 32607
rect 631 32588 733 32607
rect 767 32588 869 32607
rect 903 32588 1005 32607
rect 315 32554 321 32588
rect 359 32573 393 32588
rect 355 32554 393 32573
rect 427 32573 461 32588
rect 427 32554 465 32573
rect 499 32554 537 32588
rect 571 32573 597 32588
rect 571 32554 609 32573
rect 643 32554 681 32588
rect 715 32573 733 32588
rect 715 32554 753 32573
rect 787 32554 825 32588
rect 859 32573 869 32588
rect 859 32554 897 32573
rect 931 32554 969 32588
rect 1003 32573 1005 32588
rect 1039 32588 1141 32607
rect 1175 32588 1277 32607
rect 1311 32588 1413 32607
rect 1447 32588 1549 32607
rect 1583 32588 1685 32607
rect 1719 32588 1729 32607
rect 1039 32573 1041 32588
rect 1003 32554 1041 32573
rect 1075 32554 1113 32588
rect 1175 32573 1185 32588
rect 1147 32554 1185 32573
rect 1219 32554 1257 32588
rect 1311 32573 1329 32588
rect 1291 32554 1329 32573
rect 1363 32554 1401 32588
rect 1447 32573 1473 32588
rect 1435 32554 1473 32573
rect 1507 32554 1545 32588
rect 1583 32573 1617 32588
rect 1579 32554 1617 32573
rect 1651 32573 1685 32588
rect 1651 32554 1689 32573
rect 1723 32554 1729 32588
rect 315 32515 1729 32554
rect 315 32481 321 32515
rect 355 32481 393 32515
rect 427 32481 465 32515
rect 499 32481 537 32515
rect 571 32481 609 32515
rect 643 32481 681 32515
rect 715 32481 753 32515
rect 787 32481 825 32515
rect 859 32481 897 32515
rect 931 32481 969 32515
rect 1003 32481 1041 32515
rect 1075 32481 1113 32515
rect 1147 32481 1185 32515
rect 1219 32481 1257 32515
rect 1291 32481 1329 32515
rect 1363 32481 1401 32515
rect 1435 32481 1473 32515
rect 1507 32481 1545 32515
rect 1579 32481 1617 32515
rect 1651 32481 1689 32515
rect 1723 32481 1729 32515
rect 315 32471 1729 32481
rect 315 32442 325 32471
rect 359 32442 461 32471
rect 495 32442 597 32471
rect 631 32442 733 32471
rect 767 32442 869 32471
rect 903 32442 1005 32471
rect 315 32408 321 32442
rect 359 32437 393 32442
rect 355 32408 393 32437
rect 427 32437 461 32442
rect 427 32408 465 32437
rect 499 32408 537 32442
rect 571 32437 597 32442
rect 571 32408 609 32437
rect 643 32408 681 32442
rect 715 32437 733 32442
rect 715 32408 753 32437
rect 787 32408 825 32442
rect 859 32437 869 32442
rect 859 32408 897 32437
rect 931 32408 969 32442
rect 1003 32437 1005 32442
rect 1039 32442 1141 32471
rect 1175 32442 1277 32471
rect 1311 32442 1413 32471
rect 1447 32442 1549 32471
rect 1583 32442 1685 32471
rect 1719 32442 1729 32471
rect 1039 32437 1041 32442
rect 1003 32408 1041 32437
rect 1075 32408 1113 32442
rect 1175 32437 1185 32442
rect 1147 32408 1185 32437
rect 1219 32408 1257 32442
rect 1311 32437 1329 32442
rect 1291 32408 1329 32437
rect 1363 32408 1401 32442
rect 1447 32437 1473 32442
rect 1435 32408 1473 32437
rect 1507 32408 1545 32442
rect 1583 32437 1617 32442
rect 1579 32408 1617 32437
rect 1651 32437 1685 32442
rect 1651 32408 1689 32437
rect 1723 32408 1729 32442
rect 315 32369 1729 32408
rect 315 32335 321 32369
rect 355 32335 393 32369
rect 427 32335 465 32369
rect 499 32335 537 32369
rect 571 32335 609 32369
rect 643 32335 681 32369
rect 715 32335 753 32369
rect 787 32335 825 32369
rect 859 32335 897 32369
rect 931 32335 969 32369
rect 1003 32335 1041 32369
rect 1075 32335 1113 32369
rect 1147 32335 1185 32369
rect 1219 32335 1257 32369
rect 1291 32335 1329 32369
rect 1363 32335 1401 32369
rect 1435 32335 1473 32369
rect 1507 32335 1545 32369
rect 1579 32335 1617 32369
rect 1651 32335 1689 32369
rect 1723 32335 1729 32369
rect 315 32301 325 32335
rect 359 32301 461 32335
rect 495 32301 597 32335
rect 631 32301 733 32335
rect 767 32301 869 32335
rect 903 32301 1005 32335
rect 1039 32301 1141 32335
rect 1175 32301 1277 32335
rect 1311 32301 1413 32335
rect 1447 32301 1549 32335
rect 1583 32301 1685 32335
rect 1719 32301 1729 32335
rect 315 32296 1729 32301
rect 315 32262 321 32296
rect 355 32262 393 32296
rect 427 32262 465 32296
rect 499 32262 537 32296
rect 571 32262 609 32296
rect 643 32262 681 32296
rect 715 32262 753 32296
rect 787 32262 825 32296
rect 859 32262 897 32296
rect 931 32262 969 32296
rect 1003 32262 1041 32296
rect 1075 32262 1113 32296
rect 1147 32262 1185 32296
rect 1219 32262 1257 32296
rect 1291 32262 1329 32296
rect 1363 32262 1401 32296
rect 1435 32262 1473 32296
rect 1507 32262 1545 32296
rect 1579 32262 1617 32296
rect 1651 32262 1689 32296
rect 1723 32262 1729 32296
rect 315 32223 1729 32262
rect 315 32189 321 32223
rect 355 32199 393 32223
rect 359 32189 393 32199
rect 427 32199 465 32223
rect 427 32189 461 32199
rect 499 32189 537 32223
rect 571 32199 609 32223
rect 571 32189 597 32199
rect 643 32189 681 32223
rect 715 32199 753 32223
rect 715 32189 733 32199
rect 787 32189 825 32223
rect 859 32199 897 32223
rect 859 32189 869 32199
rect 931 32189 969 32223
rect 1003 32199 1041 32223
rect 1003 32189 1005 32199
rect 315 32165 325 32189
rect 359 32165 461 32189
rect 495 32165 597 32189
rect 631 32165 733 32189
rect 767 32165 869 32189
rect 903 32165 1005 32189
rect 1039 32189 1041 32199
rect 1075 32189 1113 32223
rect 1147 32199 1185 32223
rect 1175 32189 1185 32199
rect 1219 32189 1257 32223
rect 1291 32199 1329 32223
rect 1311 32189 1329 32199
rect 1363 32189 1401 32223
rect 1435 32199 1473 32223
rect 1447 32189 1473 32199
rect 1507 32189 1545 32223
rect 1579 32199 1617 32223
rect 1583 32189 1617 32199
rect 1651 32199 1689 32223
rect 1651 32189 1685 32199
rect 1723 32189 1729 32223
rect 1039 32165 1141 32189
rect 1175 32165 1277 32189
rect 1311 32165 1413 32189
rect 1447 32165 1549 32189
rect 1583 32165 1685 32189
rect 1719 32165 1729 32189
rect 315 32150 1729 32165
rect 315 32116 321 32150
rect 355 32116 393 32150
rect 427 32116 465 32150
rect 499 32116 537 32150
rect 571 32116 609 32150
rect 643 32116 681 32150
rect 715 32116 753 32150
rect 787 32116 825 32150
rect 859 32116 897 32150
rect 931 32116 969 32150
rect 1003 32116 1041 32150
rect 1075 32116 1113 32150
rect 1147 32116 1185 32150
rect 1219 32116 1257 32150
rect 1291 32116 1329 32150
rect 1363 32116 1401 32150
rect 1435 32116 1473 32150
rect 1507 32116 1545 32150
rect 1579 32116 1617 32150
rect 1651 32116 1689 32150
rect 1723 32116 1729 32150
rect 315 32077 1729 32116
rect 315 32043 321 32077
rect 355 32063 393 32077
rect 359 32043 393 32063
rect 427 32063 465 32077
rect 427 32043 461 32063
rect 499 32043 537 32077
rect 571 32063 609 32077
rect 571 32043 597 32063
rect 643 32043 681 32077
rect 715 32063 753 32077
rect 715 32043 733 32063
rect 787 32043 825 32077
rect 859 32063 897 32077
rect 859 32043 869 32063
rect 931 32043 969 32077
rect 1003 32063 1041 32077
rect 1003 32043 1005 32063
rect 315 32029 325 32043
rect 359 32029 461 32043
rect 495 32029 597 32043
rect 631 32029 733 32043
rect 767 32029 869 32043
rect 903 32029 1005 32043
rect 1039 32043 1041 32063
rect 1075 32043 1113 32077
rect 1147 32063 1185 32077
rect 1175 32043 1185 32063
rect 1219 32043 1257 32077
rect 1291 32063 1329 32077
rect 1311 32043 1329 32063
rect 1363 32043 1401 32077
rect 1435 32063 1473 32077
rect 1447 32043 1473 32063
rect 1507 32043 1545 32077
rect 1579 32063 1617 32077
rect 1583 32043 1617 32063
rect 1651 32063 1689 32077
rect 1651 32043 1685 32063
rect 1723 32043 1729 32077
rect 1039 32029 1141 32043
rect 1175 32029 1277 32043
rect 1311 32029 1413 32043
rect 1447 32029 1549 32043
rect 1583 32029 1685 32043
rect 1719 32029 1729 32043
rect 315 32004 1729 32029
rect 315 31970 321 32004
rect 355 31970 393 32004
rect 427 31970 465 32004
rect 499 31970 537 32004
rect 571 31970 609 32004
rect 643 31970 681 32004
rect 715 31970 753 32004
rect 787 31970 825 32004
rect 859 31970 897 32004
rect 931 31970 969 32004
rect 1003 31970 1041 32004
rect 1075 31970 1113 32004
rect 1147 31970 1185 32004
rect 1219 31970 1257 32004
rect 1291 31970 1329 32004
rect 1363 31970 1401 32004
rect 1435 31970 1473 32004
rect 1507 31970 1545 32004
rect 1579 31970 1617 32004
rect 1651 31970 1689 32004
rect 1723 31970 1729 32004
rect 315 31931 1729 31970
rect 315 31897 321 31931
rect 355 31927 393 31931
rect 359 31897 393 31927
rect 427 31927 465 31931
rect 427 31897 461 31927
rect 499 31897 537 31931
rect 571 31927 609 31931
rect 571 31897 597 31927
rect 643 31897 681 31931
rect 715 31927 753 31931
rect 715 31897 733 31927
rect 787 31897 825 31931
rect 859 31927 897 31931
rect 859 31897 869 31927
rect 931 31897 969 31931
rect 1003 31927 1041 31931
rect 1003 31897 1005 31927
rect 315 31893 325 31897
rect 359 31893 461 31897
rect 495 31893 597 31897
rect 631 31893 733 31897
rect 767 31893 869 31897
rect 903 31893 1005 31897
rect 1039 31897 1041 31927
rect 1075 31897 1113 31931
rect 1147 31927 1185 31931
rect 1175 31897 1185 31927
rect 1219 31897 1257 31931
rect 1291 31927 1329 31931
rect 1311 31897 1329 31927
rect 1363 31897 1401 31931
rect 1435 31927 1473 31931
rect 1447 31897 1473 31927
rect 1507 31897 1545 31931
rect 1579 31927 1617 31931
rect 1583 31897 1617 31927
rect 1651 31927 1689 31931
rect 1651 31897 1685 31927
rect 1723 31897 1729 31931
rect 1039 31893 1141 31897
rect 1175 31893 1277 31897
rect 1311 31893 1413 31897
rect 1447 31893 1549 31897
rect 1583 31893 1685 31897
rect 1719 31893 1729 31897
rect 315 31858 1729 31893
rect 315 31824 321 31858
rect 355 31824 393 31858
rect 427 31824 465 31858
rect 499 31824 537 31858
rect 571 31824 609 31858
rect 643 31824 681 31858
rect 715 31824 753 31858
rect 787 31824 825 31858
rect 859 31824 897 31858
rect 931 31824 969 31858
rect 1003 31824 1041 31858
rect 1075 31824 1113 31858
rect 1147 31824 1185 31858
rect 1219 31824 1257 31858
rect 1291 31824 1329 31858
rect 1363 31824 1401 31858
rect 1435 31824 1473 31858
rect 1507 31824 1545 31858
rect 1579 31824 1617 31858
rect 1651 31824 1689 31858
rect 1723 31824 1729 31858
rect 315 31791 1729 31824
rect 315 31785 325 31791
rect 359 31785 461 31791
rect 495 31785 597 31791
rect 631 31785 733 31791
rect 767 31785 869 31791
rect 903 31785 1005 31791
rect 315 31751 321 31785
rect 359 31757 393 31785
rect 355 31751 393 31757
rect 427 31757 461 31785
rect 427 31751 465 31757
rect 499 31751 537 31785
rect 571 31757 597 31785
rect 571 31751 609 31757
rect 643 31751 681 31785
rect 715 31757 733 31785
rect 715 31751 753 31757
rect 787 31751 825 31785
rect 859 31757 869 31785
rect 859 31751 897 31757
rect 931 31751 969 31785
rect 1003 31757 1005 31785
rect 1039 31785 1141 31791
rect 1175 31785 1277 31791
rect 1311 31785 1413 31791
rect 1447 31785 1549 31791
rect 1583 31785 1685 31791
rect 1719 31785 1729 31791
rect 1039 31757 1041 31785
rect 1003 31751 1041 31757
rect 1075 31751 1113 31785
rect 1175 31757 1185 31785
rect 1147 31751 1185 31757
rect 1219 31751 1257 31785
rect 1311 31757 1329 31785
rect 1291 31751 1329 31757
rect 1363 31751 1401 31785
rect 1447 31757 1473 31785
rect 1435 31751 1473 31757
rect 1507 31751 1545 31785
rect 1583 31757 1617 31785
rect 1579 31751 1617 31757
rect 1651 31757 1685 31785
rect 1651 31751 1689 31757
rect 1723 31751 1729 31785
rect 315 31712 1729 31751
rect 315 31678 321 31712
rect 355 31678 393 31712
rect 427 31678 465 31712
rect 499 31678 537 31712
rect 571 31678 609 31712
rect 643 31678 681 31712
rect 715 31678 753 31712
rect 787 31678 825 31712
rect 859 31678 897 31712
rect 931 31678 969 31712
rect 1003 31678 1041 31712
rect 1075 31678 1113 31712
rect 1147 31678 1185 31712
rect 1219 31678 1257 31712
rect 1291 31678 1329 31712
rect 1363 31678 1401 31712
rect 1435 31678 1473 31712
rect 1507 31678 1545 31712
rect 1579 31678 1617 31712
rect 1651 31678 1689 31712
rect 1723 31678 1729 31712
rect 315 31655 1729 31678
rect 315 31639 325 31655
rect 359 31639 461 31655
rect 495 31639 597 31655
rect 631 31639 733 31655
rect 767 31639 869 31655
rect 903 31639 1005 31655
rect 315 31605 321 31639
rect 359 31621 393 31639
rect 355 31605 393 31621
rect 427 31621 461 31639
rect 427 31605 465 31621
rect 499 31605 537 31639
rect 571 31621 597 31639
rect 571 31605 609 31621
rect 643 31605 681 31639
rect 715 31621 733 31639
rect 715 31605 753 31621
rect 787 31605 825 31639
rect 859 31621 869 31639
rect 859 31605 897 31621
rect 931 31605 969 31639
rect 1003 31621 1005 31639
rect 1039 31639 1141 31655
rect 1175 31639 1277 31655
rect 1311 31639 1413 31655
rect 1447 31639 1549 31655
rect 1583 31639 1685 31655
rect 1719 31639 1729 31655
rect 1039 31621 1041 31639
rect 1003 31605 1041 31621
rect 1075 31605 1113 31639
rect 1175 31621 1185 31639
rect 1147 31605 1185 31621
rect 1219 31605 1257 31639
rect 1311 31621 1329 31639
rect 1291 31605 1329 31621
rect 1363 31605 1401 31639
rect 1447 31621 1473 31639
rect 1435 31605 1473 31621
rect 1507 31605 1545 31639
rect 1583 31621 1617 31639
rect 1579 31605 1617 31621
rect 1651 31621 1685 31639
rect 1651 31605 1689 31621
rect 1723 31605 1729 31639
rect 315 31566 1729 31605
rect 315 31532 321 31566
rect 355 31532 393 31566
rect 427 31532 465 31566
rect 499 31532 537 31566
rect 571 31532 609 31566
rect 643 31532 681 31566
rect 715 31532 753 31566
rect 787 31532 825 31566
rect 859 31532 897 31566
rect 931 31532 969 31566
rect 1003 31532 1041 31566
rect 1075 31532 1113 31566
rect 1147 31532 1185 31566
rect 1219 31532 1257 31566
rect 1291 31532 1329 31566
rect 1363 31532 1401 31566
rect 1435 31532 1473 31566
rect 1507 31532 1545 31566
rect 1579 31532 1617 31566
rect 1651 31532 1689 31566
rect 1723 31532 1729 31566
rect 315 31519 1729 31532
rect 315 31493 325 31519
rect 359 31493 461 31519
rect 495 31493 597 31519
rect 631 31493 733 31519
rect 767 31493 869 31519
rect 903 31493 1005 31519
rect 315 31459 321 31493
rect 359 31485 393 31493
rect 355 31459 393 31485
rect 427 31485 461 31493
rect 427 31459 465 31485
rect 499 31459 537 31493
rect 571 31485 597 31493
rect 571 31459 609 31485
rect 643 31459 681 31493
rect 715 31485 733 31493
rect 715 31459 753 31485
rect 787 31459 825 31493
rect 859 31485 869 31493
rect 859 31459 897 31485
rect 931 31459 969 31493
rect 1003 31485 1005 31493
rect 1039 31493 1141 31519
rect 1175 31493 1277 31519
rect 1311 31493 1413 31519
rect 1447 31493 1549 31519
rect 1583 31493 1685 31519
rect 1719 31493 1729 31519
rect 1039 31485 1041 31493
rect 1003 31459 1041 31485
rect 1075 31459 1113 31493
rect 1175 31485 1185 31493
rect 1147 31459 1185 31485
rect 1219 31459 1257 31493
rect 1311 31485 1329 31493
rect 1291 31459 1329 31485
rect 1363 31459 1401 31493
rect 1447 31485 1473 31493
rect 1435 31459 1473 31485
rect 1507 31459 1545 31493
rect 1583 31485 1617 31493
rect 1579 31459 1617 31485
rect 1651 31485 1685 31493
rect 1651 31459 1689 31485
rect 1723 31459 1729 31493
rect 315 31420 1729 31459
rect 315 31386 321 31420
rect 355 31386 393 31420
rect 427 31386 465 31420
rect 499 31386 537 31420
rect 571 31386 609 31420
rect 643 31386 681 31420
rect 715 31386 753 31420
rect 787 31386 825 31420
rect 859 31386 897 31420
rect 931 31386 969 31420
rect 1003 31386 1041 31420
rect 1075 31386 1113 31420
rect 1147 31386 1185 31420
rect 1219 31386 1257 31420
rect 1291 31386 1329 31420
rect 1363 31386 1401 31420
rect 1435 31386 1473 31420
rect 1507 31386 1545 31420
rect 1579 31386 1617 31420
rect 1651 31386 1689 31420
rect 1723 31386 1729 31420
rect 315 31383 1729 31386
rect 315 31349 325 31383
rect 359 31349 461 31383
rect 495 31349 597 31383
rect 631 31349 733 31383
rect 767 31349 869 31383
rect 903 31349 1005 31383
rect 1039 31349 1141 31383
rect 1175 31349 1277 31383
rect 1311 31349 1413 31383
rect 1447 31349 1549 31383
rect 1583 31349 1685 31383
rect 1719 31349 1729 31383
rect 315 31347 1729 31349
rect 315 31313 321 31347
rect 355 31313 393 31347
rect 427 31313 465 31347
rect 499 31313 537 31347
rect 571 31313 609 31347
rect 643 31313 681 31347
rect 715 31313 753 31347
rect 787 31313 825 31347
rect 859 31313 897 31347
rect 931 31313 969 31347
rect 1003 31313 1041 31347
rect 1075 31313 1113 31347
rect 1147 31313 1185 31347
rect 1219 31313 1257 31347
rect 1291 31313 1329 31347
rect 1363 31313 1401 31347
rect 1435 31313 1473 31347
rect 1507 31313 1545 31347
rect 1579 31313 1617 31347
rect 1651 31313 1689 31347
rect 1723 31313 1729 31347
rect 315 31274 1729 31313
rect 315 31240 321 31274
rect 355 31247 393 31274
rect 359 31240 393 31247
rect 427 31247 465 31274
rect 427 31240 461 31247
rect 499 31240 537 31274
rect 571 31247 609 31274
rect 571 31240 597 31247
rect 643 31240 681 31274
rect 715 31247 753 31274
rect 715 31240 733 31247
rect 787 31240 825 31274
rect 859 31247 897 31274
rect 859 31240 869 31247
rect 931 31240 969 31274
rect 1003 31247 1041 31274
rect 1003 31240 1005 31247
rect 315 31213 325 31240
rect 359 31213 461 31240
rect 495 31213 597 31240
rect 631 31213 733 31240
rect 767 31213 869 31240
rect 903 31213 1005 31240
rect 1039 31240 1041 31247
rect 1075 31240 1113 31274
rect 1147 31247 1185 31274
rect 1175 31240 1185 31247
rect 1219 31240 1257 31274
rect 1291 31247 1329 31274
rect 1311 31240 1329 31247
rect 1363 31240 1401 31274
rect 1435 31247 1473 31274
rect 1447 31240 1473 31247
rect 1507 31240 1545 31274
rect 1579 31247 1617 31274
rect 1583 31240 1617 31247
rect 1651 31247 1689 31274
rect 1651 31240 1685 31247
rect 1723 31240 1729 31274
rect 1039 31213 1141 31240
rect 1175 31213 1277 31240
rect 1311 31213 1413 31240
rect 1447 31213 1549 31240
rect 1583 31213 1685 31240
rect 1719 31213 1729 31240
rect 315 31201 1729 31213
rect 315 31167 321 31201
rect 355 31167 393 31201
rect 427 31167 465 31201
rect 499 31167 537 31201
rect 571 31167 609 31201
rect 643 31167 681 31201
rect 715 31167 753 31201
rect 787 31167 825 31201
rect 859 31167 897 31201
rect 931 31167 969 31201
rect 1003 31167 1041 31201
rect 1075 31167 1113 31201
rect 1147 31167 1185 31201
rect 1219 31167 1257 31201
rect 1291 31167 1329 31201
rect 1363 31167 1401 31201
rect 1435 31167 1473 31201
rect 1507 31167 1545 31201
rect 1579 31167 1617 31201
rect 1651 31167 1689 31201
rect 1723 31167 1729 31201
rect 315 31128 1729 31167
rect 315 31094 321 31128
rect 355 31111 393 31128
rect 359 31094 393 31111
rect 427 31111 465 31128
rect 427 31094 461 31111
rect 499 31094 537 31128
rect 571 31111 609 31128
rect 571 31094 597 31111
rect 643 31094 681 31128
rect 715 31111 753 31128
rect 715 31094 733 31111
rect 787 31094 825 31128
rect 859 31111 897 31128
rect 859 31094 869 31111
rect 931 31094 969 31128
rect 1003 31111 1041 31128
rect 1003 31094 1005 31111
rect 315 31077 325 31094
rect 359 31077 461 31094
rect 495 31077 597 31094
rect 631 31077 733 31094
rect 767 31077 869 31094
rect 903 31077 1005 31094
rect 1039 31094 1041 31111
rect 1075 31094 1113 31128
rect 1147 31111 1185 31128
rect 1175 31094 1185 31111
rect 1219 31094 1257 31128
rect 1291 31111 1329 31128
rect 1311 31094 1329 31111
rect 1363 31094 1401 31128
rect 1435 31111 1473 31128
rect 1447 31094 1473 31111
rect 1507 31094 1545 31128
rect 1579 31111 1617 31128
rect 1583 31094 1617 31111
rect 1651 31111 1689 31128
rect 1651 31094 1685 31111
rect 1723 31094 1729 31128
rect 1039 31077 1141 31094
rect 1175 31077 1277 31094
rect 1311 31077 1413 31094
rect 1447 31077 1549 31094
rect 1583 31077 1685 31094
rect 1719 31077 1729 31094
rect 315 31055 1729 31077
rect 315 31021 321 31055
rect 355 31021 393 31055
rect 427 31021 465 31055
rect 499 31021 537 31055
rect 571 31021 609 31055
rect 643 31021 681 31055
rect 715 31021 753 31055
rect 787 31021 825 31055
rect 859 31021 897 31055
rect 931 31021 969 31055
rect 1003 31021 1041 31055
rect 1075 31021 1113 31055
rect 1147 31021 1185 31055
rect 1219 31021 1257 31055
rect 1291 31021 1329 31055
rect 1363 31021 1401 31055
rect 1435 31021 1473 31055
rect 1507 31021 1545 31055
rect 1579 31021 1617 31055
rect 1651 31021 1689 31055
rect 1723 31021 1729 31055
rect 315 30982 1729 31021
rect 315 30948 321 30982
rect 355 30975 393 30982
rect 359 30948 393 30975
rect 427 30975 465 30982
rect 427 30948 461 30975
rect 499 30948 537 30982
rect 571 30975 609 30982
rect 571 30948 597 30975
rect 643 30948 681 30982
rect 715 30975 753 30982
rect 715 30948 733 30975
rect 787 30948 825 30982
rect 859 30975 897 30982
rect 859 30948 869 30975
rect 931 30948 969 30982
rect 1003 30975 1041 30982
rect 1003 30948 1005 30975
rect 315 30941 325 30948
rect 359 30941 461 30948
rect 495 30941 597 30948
rect 631 30941 733 30948
rect 767 30941 869 30948
rect 903 30941 1005 30948
rect 1039 30948 1041 30975
rect 1075 30948 1113 30982
rect 1147 30975 1185 30982
rect 1175 30948 1185 30975
rect 1219 30948 1257 30982
rect 1291 30975 1329 30982
rect 1311 30948 1329 30975
rect 1363 30948 1401 30982
rect 1435 30975 1473 30982
rect 1447 30948 1473 30975
rect 1507 30948 1545 30982
rect 1579 30975 1617 30982
rect 1583 30948 1617 30975
rect 1651 30975 1689 30982
rect 1651 30948 1685 30975
rect 1723 30948 1729 30982
rect 1039 30941 1141 30948
rect 1175 30941 1277 30948
rect 1311 30941 1413 30948
rect 1447 30941 1549 30948
rect 1583 30941 1685 30948
rect 1719 30941 1729 30948
rect 315 30909 1729 30941
rect 315 30875 321 30909
rect 355 30875 393 30909
rect 427 30875 465 30909
rect 499 30875 537 30909
rect 571 30875 609 30909
rect 643 30875 681 30909
rect 715 30875 753 30909
rect 787 30875 825 30909
rect 859 30875 897 30909
rect 931 30875 969 30909
rect 1003 30875 1041 30909
rect 1075 30875 1113 30909
rect 1147 30875 1185 30909
rect 1219 30875 1257 30909
rect 1291 30875 1329 30909
rect 1363 30875 1401 30909
rect 1435 30875 1473 30909
rect 1507 30875 1545 30909
rect 1579 30875 1617 30909
rect 1651 30875 1689 30909
rect 1723 30875 1729 30909
rect 315 30839 1729 30875
rect 315 30836 325 30839
rect 359 30836 461 30839
rect 495 30836 597 30839
rect 631 30836 733 30839
rect 767 30836 869 30839
rect 903 30836 1005 30839
rect 315 30802 321 30836
rect 359 30805 393 30836
rect 355 30802 393 30805
rect 427 30805 461 30836
rect 427 30802 465 30805
rect 499 30802 537 30836
rect 571 30805 597 30836
rect 571 30802 609 30805
rect 643 30802 681 30836
rect 715 30805 733 30836
rect 715 30802 753 30805
rect 787 30802 825 30836
rect 859 30805 869 30836
rect 859 30802 897 30805
rect 931 30802 969 30836
rect 1003 30805 1005 30836
rect 1039 30836 1141 30839
rect 1175 30836 1277 30839
rect 1311 30836 1413 30839
rect 1447 30836 1549 30839
rect 1583 30836 1685 30839
rect 1719 30836 1729 30839
rect 1039 30805 1041 30836
rect 1003 30802 1041 30805
rect 1075 30802 1113 30836
rect 1175 30805 1185 30836
rect 1147 30802 1185 30805
rect 1219 30802 1257 30836
rect 1311 30805 1329 30836
rect 1291 30802 1329 30805
rect 1363 30802 1401 30836
rect 1447 30805 1473 30836
rect 1435 30802 1473 30805
rect 1507 30802 1545 30836
rect 1583 30805 1617 30836
rect 1579 30802 1617 30805
rect 1651 30805 1685 30836
rect 1651 30802 1689 30805
rect 1723 30802 1729 30836
rect 315 30763 1729 30802
rect 315 30729 321 30763
rect 355 30729 393 30763
rect 427 30729 465 30763
rect 499 30729 537 30763
rect 571 30729 609 30763
rect 643 30729 681 30763
rect 715 30729 753 30763
rect 787 30729 825 30763
rect 859 30729 897 30763
rect 931 30729 969 30763
rect 1003 30729 1041 30763
rect 1075 30729 1113 30763
rect 1147 30729 1185 30763
rect 1219 30729 1257 30763
rect 1291 30729 1329 30763
rect 1363 30729 1401 30763
rect 1435 30729 1473 30763
rect 1507 30729 1545 30763
rect 1579 30729 1617 30763
rect 1651 30729 1689 30763
rect 1723 30729 1729 30763
rect 315 30703 1729 30729
rect 315 30690 325 30703
rect 359 30690 461 30703
rect 495 30690 597 30703
rect 631 30690 733 30703
rect 767 30690 869 30703
rect 903 30690 1005 30703
rect 315 30656 321 30690
rect 359 30669 393 30690
rect 355 30656 393 30669
rect 427 30669 461 30690
rect 427 30656 465 30669
rect 499 30656 537 30690
rect 571 30669 597 30690
rect 571 30656 609 30669
rect 643 30656 681 30690
rect 715 30669 733 30690
rect 715 30656 753 30669
rect 787 30656 825 30690
rect 859 30669 869 30690
rect 859 30656 897 30669
rect 931 30656 969 30690
rect 1003 30669 1005 30690
rect 1039 30690 1141 30703
rect 1175 30690 1277 30703
rect 1311 30690 1413 30703
rect 1447 30690 1549 30703
rect 1583 30690 1685 30703
rect 1719 30690 1729 30703
rect 1039 30669 1041 30690
rect 1003 30656 1041 30669
rect 1075 30656 1113 30690
rect 1175 30669 1185 30690
rect 1147 30656 1185 30669
rect 1219 30656 1257 30690
rect 1311 30669 1329 30690
rect 1291 30656 1329 30669
rect 1363 30656 1401 30690
rect 1447 30669 1473 30690
rect 1435 30656 1473 30669
rect 1507 30656 1545 30690
rect 1583 30669 1617 30690
rect 1579 30656 1617 30669
rect 1651 30669 1685 30690
rect 1651 30656 1689 30669
rect 1723 30656 1729 30690
rect 315 30617 1729 30656
rect 315 30583 321 30617
rect 355 30583 393 30617
rect 427 30583 465 30617
rect 499 30583 537 30617
rect 571 30583 609 30617
rect 643 30583 681 30617
rect 715 30583 753 30617
rect 787 30583 825 30617
rect 859 30583 897 30617
rect 931 30583 969 30617
rect 1003 30583 1041 30617
rect 1075 30583 1113 30617
rect 1147 30583 1185 30617
rect 1219 30583 1257 30617
rect 1291 30583 1329 30617
rect 1363 30583 1401 30617
rect 1435 30583 1473 30617
rect 1507 30583 1545 30617
rect 1579 30583 1617 30617
rect 1651 30583 1689 30617
rect 1723 30583 1729 30617
rect 315 30567 1729 30583
rect 315 30544 325 30567
rect 359 30544 461 30567
rect 495 30544 597 30567
rect 631 30544 733 30567
rect 767 30544 869 30567
rect 903 30544 1005 30567
rect 315 30510 321 30544
rect 359 30533 393 30544
rect 355 30510 393 30533
rect 427 30533 461 30544
rect 427 30510 465 30533
rect 499 30510 537 30544
rect 571 30533 597 30544
rect 571 30510 609 30533
rect 643 30510 681 30544
rect 715 30533 733 30544
rect 715 30510 753 30533
rect 787 30510 825 30544
rect 859 30533 869 30544
rect 859 30510 897 30533
rect 931 30510 969 30544
rect 1003 30533 1005 30544
rect 1039 30544 1141 30567
rect 1175 30544 1277 30567
rect 1311 30544 1413 30567
rect 1447 30544 1549 30567
rect 1583 30544 1685 30567
rect 1719 30544 1729 30567
rect 1039 30533 1041 30544
rect 1003 30510 1041 30533
rect 1075 30510 1113 30544
rect 1175 30533 1185 30544
rect 1147 30510 1185 30533
rect 1219 30510 1257 30544
rect 1311 30533 1329 30544
rect 1291 30510 1329 30533
rect 1363 30510 1401 30544
rect 1447 30533 1473 30544
rect 1435 30510 1473 30533
rect 1507 30510 1545 30544
rect 1583 30533 1617 30544
rect 1579 30510 1617 30533
rect 1651 30533 1685 30544
rect 1651 30510 1689 30533
rect 1723 30510 1729 30544
rect 315 30471 1729 30510
rect 315 30437 321 30471
rect 355 30437 393 30471
rect 427 30437 465 30471
rect 499 30437 537 30471
rect 571 30437 609 30471
rect 643 30437 681 30471
rect 715 30437 753 30471
rect 787 30437 825 30471
rect 859 30437 897 30471
rect 931 30437 969 30471
rect 1003 30437 1041 30471
rect 1075 30437 1113 30471
rect 1147 30437 1185 30471
rect 1219 30437 1257 30471
rect 1291 30437 1329 30471
rect 1363 30437 1401 30471
rect 1435 30437 1473 30471
rect 1507 30437 1545 30471
rect 1579 30437 1617 30471
rect 1651 30437 1689 30471
rect 1723 30437 1729 30471
rect 315 30431 1729 30437
rect 315 30398 325 30431
rect 359 30398 461 30431
rect 495 30398 597 30431
rect 631 30398 733 30431
rect 767 30398 869 30431
rect 903 30398 1005 30431
rect 315 30364 321 30398
rect 359 30397 393 30398
rect 355 30364 393 30397
rect 427 30397 461 30398
rect 427 30364 465 30397
rect 499 30364 537 30398
rect 571 30397 597 30398
rect 571 30364 609 30397
rect 643 30364 681 30398
rect 715 30397 733 30398
rect 715 30364 753 30397
rect 787 30364 825 30398
rect 859 30397 869 30398
rect 859 30364 897 30397
rect 931 30364 969 30398
rect 1003 30397 1005 30398
rect 1039 30398 1141 30431
rect 1175 30398 1277 30431
rect 1311 30398 1413 30431
rect 1447 30398 1549 30431
rect 1583 30398 1685 30431
rect 1719 30398 1729 30431
rect 1039 30397 1041 30398
rect 1003 30364 1041 30397
rect 1075 30364 1113 30398
rect 1175 30397 1185 30398
rect 1147 30364 1185 30397
rect 1219 30364 1257 30398
rect 1311 30397 1329 30398
rect 1291 30364 1329 30397
rect 1363 30364 1401 30398
rect 1447 30397 1473 30398
rect 1435 30364 1473 30397
rect 1507 30364 1545 30398
rect 1583 30397 1617 30398
rect 1579 30364 1617 30397
rect 1651 30397 1685 30398
rect 1651 30364 1689 30397
rect 1723 30364 1729 30398
rect 315 30325 1729 30364
rect 315 30291 321 30325
rect 355 30295 393 30325
rect 359 30291 393 30295
rect 427 30295 465 30325
rect 427 30291 461 30295
rect 499 30291 537 30325
rect 571 30295 609 30325
rect 571 30291 597 30295
rect 643 30291 681 30325
rect 715 30295 753 30325
rect 715 30291 733 30295
rect 787 30291 825 30325
rect 859 30295 897 30325
rect 859 30291 869 30295
rect 931 30291 969 30325
rect 1003 30295 1041 30325
rect 1003 30291 1005 30295
rect 315 30261 325 30291
rect 359 30261 461 30291
rect 495 30261 597 30291
rect 631 30261 733 30291
rect 767 30261 869 30291
rect 903 30261 1005 30291
rect 1039 30291 1041 30295
rect 1075 30291 1113 30325
rect 1147 30295 1185 30325
rect 1175 30291 1185 30295
rect 1219 30291 1257 30325
rect 1291 30295 1329 30325
rect 1311 30291 1329 30295
rect 1363 30291 1401 30325
rect 1435 30295 1473 30325
rect 1447 30291 1473 30295
rect 1507 30291 1545 30325
rect 1579 30295 1617 30325
rect 1583 30291 1617 30295
rect 1651 30295 1689 30325
rect 1651 30291 1685 30295
rect 1723 30291 1729 30325
rect 1039 30261 1141 30291
rect 1175 30261 1277 30291
rect 1311 30261 1413 30291
rect 1447 30261 1549 30291
rect 1583 30261 1685 30291
rect 1719 30261 1729 30291
rect 315 30252 1729 30261
rect 315 30218 321 30252
rect 355 30218 393 30252
rect 427 30218 465 30252
rect 499 30218 537 30252
rect 571 30218 609 30252
rect 643 30218 681 30252
rect 715 30218 753 30252
rect 787 30218 825 30252
rect 859 30218 897 30252
rect 931 30218 969 30252
rect 1003 30218 1041 30252
rect 1075 30218 1113 30252
rect 1147 30218 1185 30252
rect 1219 30218 1257 30252
rect 1291 30218 1329 30252
rect 1363 30218 1401 30252
rect 1435 30218 1473 30252
rect 1507 30218 1545 30252
rect 1579 30218 1617 30252
rect 1651 30218 1689 30252
rect 1723 30218 1729 30252
rect 315 30179 1729 30218
rect 315 30145 321 30179
rect 355 30159 393 30179
rect 359 30145 393 30159
rect 427 30159 465 30179
rect 427 30145 461 30159
rect 499 30145 537 30179
rect 571 30159 609 30179
rect 571 30145 597 30159
rect 643 30145 681 30179
rect 715 30159 753 30179
rect 715 30145 733 30159
rect 787 30145 825 30179
rect 859 30159 897 30179
rect 859 30145 869 30159
rect 931 30145 969 30179
rect 1003 30159 1041 30179
rect 1003 30145 1005 30159
rect 315 30125 325 30145
rect 359 30125 461 30145
rect 495 30125 597 30145
rect 631 30125 733 30145
rect 767 30125 869 30145
rect 903 30125 1005 30145
rect 1039 30145 1041 30159
rect 1075 30145 1113 30179
rect 1147 30159 1185 30179
rect 1175 30145 1185 30159
rect 1219 30145 1257 30179
rect 1291 30159 1329 30179
rect 1311 30145 1329 30159
rect 1363 30145 1401 30179
rect 1435 30159 1473 30179
rect 1447 30145 1473 30159
rect 1507 30145 1545 30179
rect 1579 30159 1617 30179
rect 1583 30145 1617 30159
rect 1651 30159 1689 30179
rect 1651 30145 1685 30159
rect 1723 30145 1729 30179
rect 1039 30125 1141 30145
rect 1175 30125 1277 30145
rect 1311 30125 1413 30145
rect 1447 30125 1549 30145
rect 1583 30125 1685 30145
rect 1719 30125 1729 30145
rect 315 30106 1729 30125
rect 315 30072 321 30106
rect 355 30072 393 30106
rect 427 30072 465 30106
rect 499 30072 537 30106
rect 571 30072 609 30106
rect 643 30072 681 30106
rect 715 30072 753 30106
rect 787 30072 825 30106
rect 859 30072 897 30106
rect 931 30072 969 30106
rect 1003 30072 1041 30106
rect 1075 30072 1113 30106
rect 1147 30072 1185 30106
rect 1219 30072 1257 30106
rect 1291 30072 1329 30106
rect 1363 30072 1401 30106
rect 1435 30072 1473 30106
rect 1507 30072 1545 30106
rect 1579 30072 1617 30106
rect 1651 30072 1689 30106
rect 1723 30072 1729 30106
rect 315 30033 1729 30072
rect 315 29999 321 30033
rect 355 30023 393 30033
rect 359 29999 393 30023
rect 427 30023 465 30033
rect 427 29999 461 30023
rect 499 29999 537 30033
rect 571 30023 609 30033
rect 571 29999 597 30023
rect 643 29999 681 30033
rect 715 30023 753 30033
rect 715 29999 733 30023
rect 787 29999 825 30033
rect 859 30023 897 30033
rect 859 29999 869 30023
rect 931 29999 969 30033
rect 1003 30023 1041 30033
rect 1003 29999 1005 30023
rect 315 29989 325 29999
rect 359 29989 461 29999
rect 495 29989 597 29999
rect 631 29989 733 29999
rect 767 29989 869 29999
rect 903 29989 1005 29999
rect 1039 29999 1041 30023
rect 1075 29999 1113 30033
rect 1147 30023 1185 30033
rect 1175 29999 1185 30023
rect 1219 29999 1257 30033
rect 1291 30023 1329 30033
rect 1311 29999 1329 30023
rect 1363 29999 1401 30033
rect 1435 30023 1473 30033
rect 1447 29999 1473 30023
rect 1507 29999 1545 30033
rect 1579 30023 1617 30033
rect 1583 29999 1617 30023
rect 1651 30023 1689 30033
rect 1651 29999 1685 30023
rect 1723 29999 1729 30033
rect 1039 29989 1141 29999
rect 1175 29989 1277 29999
rect 1311 29989 1413 29999
rect 1447 29989 1549 29999
rect 1583 29989 1685 29999
rect 1719 29989 1729 29999
rect 315 29960 1729 29989
rect 315 29926 321 29960
rect 355 29926 393 29960
rect 427 29926 465 29960
rect 499 29926 537 29960
rect 571 29926 609 29960
rect 643 29926 681 29960
rect 715 29926 753 29960
rect 787 29926 825 29960
rect 859 29926 897 29960
rect 931 29926 969 29960
rect 1003 29926 1041 29960
rect 1075 29926 1113 29960
rect 1147 29926 1185 29960
rect 1219 29926 1257 29960
rect 1291 29926 1329 29960
rect 1363 29926 1401 29960
rect 1435 29926 1473 29960
rect 1507 29926 1545 29960
rect 1579 29926 1617 29960
rect 1651 29926 1689 29960
rect 1723 29926 1729 29960
rect 315 29887 1729 29926
rect 315 29853 321 29887
rect 359 29853 393 29887
rect 427 29853 461 29887
rect 499 29853 537 29887
rect 571 29853 597 29887
rect 643 29853 681 29887
rect 715 29853 733 29887
rect 787 29853 825 29887
rect 859 29853 869 29887
rect 931 29853 969 29887
rect 1003 29853 1005 29887
rect 1039 29853 1041 29887
rect 1075 29853 1113 29887
rect 1175 29853 1185 29887
rect 1219 29853 1257 29887
rect 1311 29853 1329 29887
rect 1363 29853 1401 29887
rect 1447 29853 1473 29887
rect 1507 29853 1545 29887
rect 1583 29853 1617 29887
rect 1651 29853 1685 29887
rect 1723 29853 1729 29887
rect 315 29814 1729 29853
rect 315 29780 321 29814
rect 355 29780 393 29814
rect 427 29780 465 29814
rect 499 29780 537 29814
rect 571 29780 609 29814
rect 643 29780 681 29814
rect 715 29780 753 29814
rect 787 29780 825 29814
rect 859 29780 897 29814
rect 931 29780 969 29814
rect 1003 29780 1041 29814
rect 1075 29780 1113 29814
rect 1147 29780 1185 29814
rect 1219 29780 1257 29814
rect 1291 29780 1329 29814
rect 1363 29780 1401 29814
rect 1435 29780 1473 29814
rect 1507 29780 1545 29814
rect 1579 29780 1617 29814
rect 1651 29780 1689 29814
rect 1723 29780 1729 29814
rect 315 29751 1729 29780
rect 315 29741 325 29751
rect 359 29741 461 29751
rect 495 29741 597 29751
rect 631 29741 733 29751
rect 767 29741 869 29751
rect 903 29741 1005 29751
rect 315 29707 321 29741
rect 359 29717 393 29741
rect 355 29707 393 29717
rect 427 29717 461 29741
rect 427 29707 465 29717
rect 499 29707 537 29741
rect 571 29717 597 29741
rect 571 29707 609 29717
rect 643 29707 681 29741
rect 715 29717 733 29741
rect 715 29707 753 29717
rect 787 29707 825 29741
rect 859 29717 869 29741
rect 859 29707 897 29717
rect 931 29707 969 29741
rect 1003 29717 1005 29741
rect 1039 29741 1141 29751
rect 1175 29741 1277 29751
rect 1311 29741 1413 29751
rect 1447 29741 1549 29751
rect 1583 29741 1685 29751
rect 1719 29741 1729 29751
rect 1039 29717 1041 29741
rect 1003 29707 1041 29717
rect 1075 29707 1113 29741
rect 1175 29717 1185 29741
rect 1147 29707 1185 29717
rect 1219 29707 1257 29741
rect 1311 29717 1329 29741
rect 1291 29707 1329 29717
rect 1363 29707 1401 29741
rect 1447 29717 1473 29741
rect 1435 29707 1473 29717
rect 1507 29707 1545 29741
rect 1583 29717 1617 29741
rect 1579 29707 1617 29717
rect 1651 29717 1685 29741
rect 1651 29707 1689 29717
rect 1723 29707 1729 29741
rect 315 29668 1729 29707
rect 315 29634 321 29668
rect 355 29634 393 29668
rect 427 29634 465 29668
rect 499 29634 537 29668
rect 571 29634 609 29668
rect 643 29634 681 29668
rect 715 29634 753 29668
rect 787 29634 825 29668
rect 859 29634 897 29668
rect 931 29634 969 29668
rect 1003 29634 1041 29668
rect 1075 29634 1113 29668
rect 1147 29634 1185 29668
rect 1219 29634 1257 29668
rect 1291 29634 1329 29668
rect 1363 29634 1401 29668
rect 1435 29634 1473 29668
rect 1507 29634 1545 29668
rect 1579 29634 1617 29668
rect 1651 29634 1689 29668
rect 1723 29634 1729 29668
rect 315 29615 1729 29634
rect 315 29602 325 29615
rect 359 29581 461 29615
rect 495 29581 597 29615
rect 631 29581 733 29615
rect 767 29581 869 29615
rect 903 29581 1005 29615
rect 1039 29581 1141 29615
rect 1175 29581 1277 29615
rect 1311 29581 1413 29615
rect 1447 29581 1549 29615
rect 1583 29581 1685 29615
rect 1719 29602 1729 29615
rect 7870 39951 9284 39975
rect 7870 39943 7880 39951
rect 7914 39943 8016 39951
rect 8050 39943 8152 39951
rect 8186 39943 8288 39951
rect 8322 39943 8424 39951
rect 8458 39943 8560 39951
rect 8594 39943 8696 39951
rect 8730 39943 8832 39951
rect 8866 39943 8968 39951
rect 9002 39943 9104 39951
rect 9138 39943 9240 39951
rect 9274 39943 9284 39951
rect 7870 33357 7876 39943
rect 9278 33357 9284 39943
rect 7870 33318 9284 33357
rect 7870 33284 7876 33318
rect 7910 33287 7948 33318
rect 7914 33284 7948 33287
rect 7982 33287 8020 33318
rect 7982 33284 8016 33287
rect 8054 33284 8092 33318
rect 8126 33287 8164 33318
rect 8126 33284 8152 33287
rect 8198 33284 8236 33318
rect 8270 33287 8308 33318
rect 8270 33284 8288 33287
rect 8342 33284 8380 33318
rect 8414 33287 8452 33318
rect 8414 33284 8424 33287
rect 8486 33284 8524 33318
rect 8558 33287 8596 33318
rect 8558 33284 8560 33287
rect 7870 33253 7880 33284
rect 7914 33253 8016 33284
rect 8050 33253 8152 33284
rect 8186 33253 8288 33284
rect 8322 33253 8424 33284
rect 8458 33253 8560 33284
rect 8594 33284 8596 33287
rect 8630 33284 8668 33318
rect 8702 33287 8740 33318
rect 8730 33284 8740 33287
rect 8774 33284 8812 33318
rect 8846 33287 8884 33318
rect 8866 33284 8884 33287
rect 8918 33284 8956 33318
rect 8990 33287 9028 33318
rect 9002 33284 9028 33287
rect 9062 33284 9100 33318
rect 9134 33287 9172 33318
rect 9138 33284 9172 33287
rect 9206 33287 9244 33318
rect 9206 33284 9240 33287
rect 9278 33284 9284 33318
rect 8594 33253 8696 33284
rect 8730 33253 8832 33284
rect 8866 33253 8968 33284
rect 9002 33253 9104 33284
rect 9138 33253 9240 33284
rect 9274 33253 9284 33284
rect 7870 33245 9284 33253
rect 7870 33211 7876 33245
rect 7910 33211 7948 33245
rect 7982 33211 8020 33245
rect 8054 33211 8092 33245
rect 8126 33211 8164 33245
rect 8198 33211 8236 33245
rect 8270 33211 8308 33245
rect 8342 33211 8380 33245
rect 8414 33211 8452 33245
rect 8486 33211 8524 33245
rect 8558 33211 8596 33245
rect 8630 33211 8668 33245
rect 8702 33211 8740 33245
rect 8774 33211 8812 33245
rect 8846 33211 8884 33245
rect 8918 33211 8956 33245
rect 8990 33211 9028 33245
rect 9062 33211 9100 33245
rect 9134 33211 9172 33245
rect 9206 33211 9244 33245
rect 9278 33211 9284 33245
rect 7870 33172 9284 33211
rect 7870 33138 7876 33172
rect 7910 33151 7948 33172
rect 7914 33138 7948 33151
rect 7982 33151 8020 33172
rect 7982 33138 8016 33151
rect 8054 33138 8092 33172
rect 8126 33151 8164 33172
rect 8126 33138 8152 33151
rect 8198 33138 8236 33172
rect 8270 33151 8308 33172
rect 8270 33138 8288 33151
rect 8342 33138 8380 33172
rect 8414 33151 8452 33172
rect 8414 33138 8424 33151
rect 8486 33138 8524 33172
rect 8558 33151 8596 33172
rect 8558 33138 8560 33151
rect 7870 33117 7880 33138
rect 7914 33117 8016 33138
rect 8050 33117 8152 33138
rect 8186 33117 8288 33138
rect 8322 33117 8424 33138
rect 8458 33117 8560 33138
rect 8594 33138 8596 33151
rect 8630 33138 8668 33172
rect 8702 33151 8740 33172
rect 8730 33138 8740 33151
rect 8774 33138 8812 33172
rect 8846 33151 8884 33172
rect 8866 33138 8884 33151
rect 8918 33138 8956 33172
rect 8990 33151 9028 33172
rect 9002 33138 9028 33151
rect 9062 33138 9100 33172
rect 9134 33151 9172 33172
rect 9138 33138 9172 33151
rect 9206 33151 9244 33172
rect 9206 33138 9240 33151
rect 9278 33138 9284 33172
rect 8594 33117 8696 33138
rect 8730 33117 8832 33138
rect 8866 33117 8968 33138
rect 9002 33117 9104 33138
rect 9138 33117 9240 33138
rect 9274 33117 9284 33138
rect 7870 33099 9284 33117
rect 7870 33065 7876 33099
rect 7910 33065 7948 33099
rect 7982 33065 8020 33099
rect 8054 33065 8092 33099
rect 8126 33065 8164 33099
rect 8198 33065 8236 33099
rect 8270 33065 8308 33099
rect 8342 33065 8380 33099
rect 8414 33065 8452 33099
rect 8486 33065 8524 33099
rect 8558 33065 8596 33099
rect 8630 33065 8668 33099
rect 8702 33065 8740 33099
rect 8774 33065 8812 33099
rect 8846 33065 8884 33099
rect 8918 33065 8956 33099
rect 8990 33065 9028 33099
rect 9062 33065 9100 33099
rect 9134 33065 9172 33099
rect 9206 33065 9244 33099
rect 9278 33065 9284 33099
rect 7870 33026 9284 33065
rect 7870 32992 7876 33026
rect 7910 33015 7948 33026
rect 7914 32992 7948 33015
rect 7982 33015 8020 33026
rect 7982 32992 8016 33015
rect 8054 32992 8092 33026
rect 8126 33015 8164 33026
rect 8126 32992 8152 33015
rect 8198 32992 8236 33026
rect 8270 33015 8308 33026
rect 8270 32992 8288 33015
rect 8342 32992 8380 33026
rect 8414 33015 8452 33026
rect 8414 32992 8424 33015
rect 8486 32992 8524 33026
rect 8558 33015 8596 33026
rect 8558 32992 8560 33015
rect 7870 32981 7880 32992
rect 7914 32981 8016 32992
rect 8050 32981 8152 32992
rect 8186 32981 8288 32992
rect 8322 32981 8424 32992
rect 8458 32981 8560 32992
rect 8594 32992 8596 33015
rect 8630 32992 8668 33026
rect 8702 33015 8740 33026
rect 8730 32992 8740 33015
rect 8774 32992 8812 33026
rect 8846 33015 8884 33026
rect 8866 32992 8884 33015
rect 8918 32992 8956 33026
rect 8990 33015 9028 33026
rect 9002 32992 9028 33015
rect 9062 32992 9100 33026
rect 9134 33015 9172 33026
rect 9138 32992 9172 33015
rect 9206 33015 9244 33026
rect 9206 32992 9240 33015
rect 9278 32992 9284 33026
rect 8594 32981 8696 32992
rect 8730 32981 8832 32992
rect 8866 32981 8968 32992
rect 9002 32981 9104 32992
rect 9138 32981 9240 32992
rect 9274 32981 9284 32992
rect 7870 32953 9284 32981
rect 7870 32919 7876 32953
rect 7910 32919 7948 32953
rect 7982 32919 8020 32953
rect 8054 32919 8092 32953
rect 8126 32919 8164 32953
rect 8198 32919 8236 32953
rect 8270 32919 8308 32953
rect 8342 32919 8380 32953
rect 8414 32919 8452 32953
rect 8486 32919 8524 32953
rect 8558 32919 8596 32953
rect 8630 32919 8668 32953
rect 8702 32919 8740 32953
rect 8774 32919 8812 32953
rect 8846 32919 8884 32953
rect 8918 32919 8956 32953
rect 8990 32919 9028 32953
rect 9062 32919 9100 32953
rect 9134 32919 9172 32953
rect 9206 32919 9244 32953
rect 9278 32919 9284 32953
rect 7870 32880 9284 32919
rect 7870 32846 7876 32880
rect 7910 32879 7948 32880
rect 7914 32846 7948 32879
rect 7982 32879 8020 32880
rect 7982 32846 8016 32879
rect 8054 32846 8092 32880
rect 8126 32879 8164 32880
rect 8126 32846 8152 32879
rect 8198 32846 8236 32880
rect 8270 32879 8308 32880
rect 8270 32846 8288 32879
rect 8342 32846 8380 32880
rect 8414 32879 8452 32880
rect 8414 32846 8424 32879
rect 8486 32846 8524 32880
rect 8558 32879 8596 32880
rect 8558 32846 8560 32879
rect 7870 32845 7880 32846
rect 7914 32845 8016 32846
rect 8050 32845 8152 32846
rect 8186 32845 8288 32846
rect 8322 32845 8424 32846
rect 8458 32845 8560 32846
rect 8594 32846 8596 32879
rect 8630 32846 8668 32880
rect 8702 32879 8740 32880
rect 8730 32846 8740 32879
rect 8774 32846 8812 32880
rect 8846 32879 8884 32880
rect 8866 32846 8884 32879
rect 8918 32846 8956 32880
rect 8990 32879 9028 32880
rect 9002 32846 9028 32879
rect 9062 32846 9100 32880
rect 9134 32879 9172 32880
rect 9138 32846 9172 32879
rect 9206 32879 9244 32880
rect 9206 32846 9240 32879
rect 9278 32846 9284 32880
rect 8594 32845 8696 32846
rect 8730 32845 8832 32846
rect 8866 32845 8968 32846
rect 9002 32845 9104 32846
rect 9138 32845 9240 32846
rect 9274 32845 9284 32846
rect 7870 32807 9284 32845
rect 7870 32773 7876 32807
rect 7910 32773 7948 32807
rect 7982 32773 8020 32807
rect 8054 32773 8092 32807
rect 8126 32773 8164 32807
rect 8198 32773 8236 32807
rect 8270 32773 8308 32807
rect 8342 32773 8380 32807
rect 8414 32773 8452 32807
rect 8486 32773 8524 32807
rect 8558 32773 8596 32807
rect 8630 32773 8668 32807
rect 8702 32773 8740 32807
rect 8774 32773 8812 32807
rect 8846 32773 8884 32807
rect 8918 32773 8956 32807
rect 8990 32773 9028 32807
rect 9062 32773 9100 32807
rect 9134 32773 9172 32807
rect 9206 32773 9244 32807
rect 9278 32773 9284 32807
rect 7870 32743 9284 32773
rect 7870 32734 7880 32743
rect 7914 32734 8016 32743
rect 8050 32734 8152 32743
rect 8186 32734 8288 32743
rect 8322 32734 8424 32743
rect 8458 32734 8560 32743
rect 7870 32700 7876 32734
rect 7914 32709 7948 32734
rect 7910 32700 7948 32709
rect 7982 32709 8016 32734
rect 7982 32700 8020 32709
rect 8054 32700 8092 32734
rect 8126 32709 8152 32734
rect 8126 32700 8164 32709
rect 8198 32700 8236 32734
rect 8270 32709 8288 32734
rect 8270 32700 8308 32709
rect 8342 32700 8380 32734
rect 8414 32709 8424 32734
rect 8414 32700 8452 32709
rect 8486 32700 8524 32734
rect 8558 32709 8560 32734
rect 8594 32734 8696 32743
rect 8730 32734 8832 32743
rect 8866 32734 8968 32743
rect 9002 32734 9104 32743
rect 9138 32734 9240 32743
rect 9274 32734 9284 32743
rect 8594 32709 8596 32734
rect 8558 32700 8596 32709
rect 8630 32700 8668 32734
rect 8730 32709 8740 32734
rect 8702 32700 8740 32709
rect 8774 32700 8812 32734
rect 8866 32709 8884 32734
rect 8846 32700 8884 32709
rect 8918 32700 8956 32734
rect 9002 32709 9028 32734
rect 8990 32700 9028 32709
rect 9062 32700 9100 32734
rect 9138 32709 9172 32734
rect 9134 32700 9172 32709
rect 9206 32709 9240 32734
rect 9206 32700 9244 32709
rect 9278 32700 9284 32734
rect 7870 32661 9284 32700
rect 7870 32627 7876 32661
rect 7910 32627 7948 32661
rect 7982 32627 8020 32661
rect 8054 32627 8092 32661
rect 8126 32627 8164 32661
rect 8198 32627 8236 32661
rect 8270 32627 8308 32661
rect 8342 32627 8380 32661
rect 8414 32627 8452 32661
rect 8486 32627 8524 32661
rect 8558 32627 8596 32661
rect 8630 32627 8668 32661
rect 8702 32627 8740 32661
rect 8774 32627 8812 32661
rect 8846 32627 8884 32661
rect 8918 32627 8956 32661
rect 8990 32627 9028 32661
rect 9062 32627 9100 32661
rect 9134 32627 9172 32661
rect 9206 32627 9244 32661
rect 9278 32627 9284 32661
rect 7870 32607 9284 32627
rect 7870 32588 7880 32607
rect 7914 32588 8016 32607
rect 8050 32588 8152 32607
rect 8186 32588 8288 32607
rect 8322 32588 8424 32607
rect 8458 32588 8560 32607
rect 7870 32554 7876 32588
rect 7914 32573 7948 32588
rect 7910 32554 7948 32573
rect 7982 32573 8016 32588
rect 7982 32554 8020 32573
rect 8054 32554 8092 32588
rect 8126 32573 8152 32588
rect 8126 32554 8164 32573
rect 8198 32554 8236 32588
rect 8270 32573 8288 32588
rect 8270 32554 8308 32573
rect 8342 32554 8380 32588
rect 8414 32573 8424 32588
rect 8414 32554 8452 32573
rect 8486 32554 8524 32588
rect 8558 32573 8560 32588
rect 8594 32588 8696 32607
rect 8730 32588 8832 32607
rect 8866 32588 8968 32607
rect 9002 32588 9104 32607
rect 9138 32588 9240 32607
rect 9274 32588 9284 32607
rect 8594 32573 8596 32588
rect 8558 32554 8596 32573
rect 8630 32554 8668 32588
rect 8730 32573 8740 32588
rect 8702 32554 8740 32573
rect 8774 32554 8812 32588
rect 8866 32573 8884 32588
rect 8846 32554 8884 32573
rect 8918 32554 8956 32588
rect 9002 32573 9028 32588
rect 8990 32554 9028 32573
rect 9062 32554 9100 32588
rect 9138 32573 9172 32588
rect 9134 32554 9172 32573
rect 9206 32573 9240 32588
rect 9206 32554 9244 32573
rect 9278 32554 9284 32588
rect 7870 32515 9284 32554
rect 7870 32481 7876 32515
rect 7910 32481 7948 32515
rect 7982 32481 8020 32515
rect 8054 32481 8092 32515
rect 8126 32481 8164 32515
rect 8198 32481 8236 32515
rect 8270 32481 8308 32515
rect 8342 32481 8380 32515
rect 8414 32481 8452 32515
rect 8486 32481 8524 32515
rect 8558 32481 8596 32515
rect 8630 32481 8668 32515
rect 8702 32481 8740 32515
rect 8774 32481 8812 32515
rect 8846 32481 8884 32515
rect 8918 32481 8956 32515
rect 8990 32481 9028 32515
rect 9062 32481 9100 32515
rect 9134 32481 9172 32515
rect 9206 32481 9244 32515
rect 9278 32481 9284 32515
rect 7870 32471 9284 32481
rect 7870 32442 7880 32471
rect 7914 32442 8016 32471
rect 8050 32442 8152 32471
rect 8186 32442 8288 32471
rect 8322 32442 8424 32471
rect 8458 32442 8560 32471
rect 7870 32408 7876 32442
rect 7914 32437 7948 32442
rect 7910 32408 7948 32437
rect 7982 32437 8016 32442
rect 7982 32408 8020 32437
rect 8054 32408 8092 32442
rect 8126 32437 8152 32442
rect 8126 32408 8164 32437
rect 8198 32408 8236 32442
rect 8270 32437 8288 32442
rect 8270 32408 8308 32437
rect 8342 32408 8380 32442
rect 8414 32437 8424 32442
rect 8414 32408 8452 32437
rect 8486 32408 8524 32442
rect 8558 32437 8560 32442
rect 8594 32442 8696 32471
rect 8730 32442 8832 32471
rect 8866 32442 8968 32471
rect 9002 32442 9104 32471
rect 9138 32442 9240 32471
rect 9274 32442 9284 32471
rect 8594 32437 8596 32442
rect 8558 32408 8596 32437
rect 8630 32408 8668 32442
rect 8730 32437 8740 32442
rect 8702 32408 8740 32437
rect 8774 32408 8812 32442
rect 8866 32437 8884 32442
rect 8846 32408 8884 32437
rect 8918 32408 8956 32442
rect 9002 32437 9028 32442
rect 8990 32408 9028 32437
rect 9062 32408 9100 32442
rect 9138 32437 9172 32442
rect 9134 32408 9172 32437
rect 9206 32437 9240 32442
rect 9206 32408 9244 32437
rect 9278 32408 9284 32442
rect 7870 32369 9284 32408
rect 7870 32335 7876 32369
rect 7910 32335 7948 32369
rect 7982 32335 8020 32369
rect 8054 32335 8092 32369
rect 8126 32335 8164 32369
rect 8198 32335 8236 32369
rect 8270 32335 8308 32369
rect 8342 32335 8380 32369
rect 8414 32335 8452 32369
rect 8486 32335 8524 32369
rect 8558 32335 8596 32369
rect 8630 32335 8668 32369
rect 8702 32335 8740 32369
rect 8774 32335 8812 32369
rect 8846 32335 8884 32369
rect 8918 32335 8956 32369
rect 8990 32335 9028 32369
rect 9062 32335 9100 32369
rect 9134 32335 9172 32369
rect 9206 32335 9244 32369
rect 9278 32335 9284 32369
rect 7870 32301 7880 32335
rect 7914 32301 8016 32335
rect 8050 32301 8152 32335
rect 8186 32301 8288 32335
rect 8322 32301 8424 32335
rect 8458 32301 8560 32335
rect 8594 32301 8696 32335
rect 8730 32301 8832 32335
rect 8866 32301 8968 32335
rect 9002 32301 9104 32335
rect 9138 32301 9240 32335
rect 9274 32301 9284 32335
rect 7870 32296 9284 32301
rect 7870 32262 7876 32296
rect 7910 32262 7948 32296
rect 7982 32262 8020 32296
rect 8054 32262 8092 32296
rect 8126 32262 8164 32296
rect 8198 32262 8236 32296
rect 8270 32262 8308 32296
rect 8342 32262 8380 32296
rect 8414 32262 8452 32296
rect 8486 32262 8524 32296
rect 8558 32262 8596 32296
rect 8630 32262 8668 32296
rect 8702 32262 8740 32296
rect 8774 32262 8812 32296
rect 8846 32262 8884 32296
rect 8918 32262 8956 32296
rect 8990 32262 9028 32296
rect 9062 32262 9100 32296
rect 9134 32262 9172 32296
rect 9206 32262 9244 32296
rect 9278 32262 9284 32296
rect 7870 32223 9284 32262
rect 7870 32189 7876 32223
rect 7910 32199 7948 32223
rect 7914 32189 7948 32199
rect 7982 32199 8020 32223
rect 7982 32189 8016 32199
rect 8054 32189 8092 32223
rect 8126 32199 8164 32223
rect 8126 32189 8152 32199
rect 8198 32189 8236 32223
rect 8270 32199 8308 32223
rect 8270 32189 8288 32199
rect 8342 32189 8380 32223
rect 8414 32199 8452 32223
rect 8414 32189 8424 32199
rect 8486 32189 8524 32223
rect 8558 32199 8596 32223
rect 8558 32189 8560 32199
rect 7870 32165 7880 32189
rect 7914 32165 8016 32189
rect 8050 32165 8152 32189
rect 8186 32165 8288 32189
rect 8322 32165 8424 32189
rect 8458 32165 8560 32189
rect 8594 32189 8596 32199
rect 8630 32189 8668 32223
rect 8702 32199 8740 32223
rect 8730 32189 8740 32199
rect 8774 32189 8812 32223
rect 8846 32199 8884 32223
rect 8866 32189 8884 32199
rect 8918 32189 8956 32223
rect 8990 32199 9028 32223
rect 9002 32189 9028 32199
rect 9062 32189 9100 32223
rect 9134 32199 9172 32223
rect 9138 32189 9172 32199
rect 9206 32199 9244 32223
rect 9206 32189 9240 32199
rect 9278 32189 9284 32223
rect 8594 32165 8696 32189
rect 8730 32165 8832 32189
rect 8866 32165 8968 32189
rect 9002 32165 9104 32189
rect 9138 32165 9240 32189
rect 9274 32165 9284 32189
rect 7870 32150 9284 32165
rect 7870 32116 7876 32150
rect 7910 32116 7948 32150
rect 7982 32116 8020 32150
rect 8054 32116 8092 32150
rect 8126 32116 8164 32150
rect 8198 32116 8236 32150
rect 8270 32116 8308 32150
rect 8342 32116 8380 32150
rect 8414 32116 8452 32150
rect 8486 32116 8524 32150
rect 8558 32116 8596 32150
rect 8630 32116 8668 32150
rect 8702 32116 8740 32150
rect 8774 32116 8812 32150
rect 8846 32116 8884 32150
rect 8918 32116 8956 32150
rect 8990 32116 9028 32150
rect 9062 32116 9100 32150
rect 9134 32116 9172 32150
rect 9206 32116 9244 32150
rect 9278 32116 9284 32150
rect 7870 32077 9284 32116
rect 7870 32043 7876 32077
rect 7910 32063 7948 32077
rect 7914 32043 7948 32063
rect 7982 32063 8020 32077
rect 7982 32043 8016 32063
rect 8054 32043 8092 32077
rect 8126 32063 8164 32077
rect 8126 32043 8152 32063
rect 8198 32043 8236 32077
rect 8270 32063 8308 32077
rect 8270 32043 8288 32063
rect 8342 32043 8380 32077
rect 8414 32063 8452 32077
rect 8414 32043 8424 32063
rect 8486 32043 8524 32077
rect 8558 32063 8596 32077
rect 8558 32043 8560 32063
rect 7870 32029 7880 32043
rect 7914 32029 8016 32043
rect 8050 32029 8152 32043
rect 8186 32029 8288 32043
rect 8322 32029 8424 32043
rect 8458 32029 8560 32043
rect 8594 32043 8596 32063
rect 8630 32043 8668 32077
rect 8702 32063 8740 32077
rect 8730 32043 8740 32063
rect 8774 32043 8812 32077
rect 8846 32063 8884 32077
rect 8866 32043 8884 32063
rect 8918 32043 8956 32077
rect 8990 32063 9028 32077
rect 9002 32043 9028 32063
rect 9062 32043 9100 32077
rect 9134 32063 9172 32077
rect 9138 32043 9172 32063
rect 9206 32063 9244 32077
rect 9206 32043 9240 32063
rect 9278 32043 9284 32077
rect 8594 32029 8696 32043
rect 8730 32029 8832 32043
rect 8866 32029 8968 32043
rect 9002 32029 9104 32043
rect 9138 32029 9240 32043
rect 9274 32029 9284 32043
rect 7870 32004 9284 32029
rect 7870 31970 7876 32004
rect 7910 31970 7948 32004
rect 7982 31970 8020 32004
rect 8054 31970 8092 32004
rect 8126 31970 8164 32004
rect 8198 31970 8236 32004
rect 8270 31970 8308 32004
rect 8342 31970 8380 32004
rect 8414 31970 8452 32004
rect 8486 31970 8524 32004
rect 8558 31970 8596 32004
rect 8630 31970 8668 32004
rect 8702 31970 8740 32004
rect 8774 31970 8812 32004
rect 8846 31970 8884 32004
rect 8918 31970 8956 32004
rect 8990 31970 9028 32004
rect 9062 31970 9100 32004
rect 9134 31970 9172 32004
rect 9206 31970 9244 32004
rect 9278 31970 9284 32004
rect 7870 31931 9284 31970
rect 7870 31897 7876 31931
rect 7910 31927 7948 31931
rect 7914 31897 7948 31927
rect 7982 31927 8020 31931
rect 7982 31897 8016 31927
rect 8054 31897 8092 31931
rect 8126 31927 8164 31931
rect 8126 31897 8152 31927
rect 8198 31897 8236 31931
rect 8270 31927 8308 31931
rect 8270 31897 8288 31927
rect 8342 31897 8380 31931
rect 8414 31927 8452 31931
rect 8414 31897 8424 31927
rect 8486 31897 8524 31931
rect 8558 31927 8596 31931
rect 8558 31897 8560 31927
rect 7870 31893 7880 31897
rect 7914 31893 8016 31897
rect 8050 31893 8152 31897
rect 8186 31893 8288 31897
rect 8322 31893 8424 31897
rect 8458 31893 8560 31897
rect 8594 31897 8596 31927
rect 8630 31897 8668 31931
rect 8702 31927 8740 31931
rect 8730 31897 8740 31927
rect 8774 31897 8812 31931
rect 8846 31927 8884 31931
rect 8866 31897 8884 31927
rect 8918 31897 8956 31931
rect 8990 31927 9028 31931
rect 9002 31897 9028 31927
rect 9062 31897 9100 31931
rect 9134 31927 9172 31931
rect 9138 31897 9172 31927
rect 9206 31927 9244 31931
rect 9206 31897 9240 31927
rect 9278 31897 9284 31931
rect 8594 31893 8696 31897
rect 8730 31893 8832 31897
rect 8866 31893 8968 31897
rect 9002 31893 9104 31897
rect 9138 31893 9240 31897
rect 9274 31893 9284 31897
rect 7870 31858 9284 31893
rect 7870 31824 7876 31858
rect 7910 31824 7948 31858
rect 7982 31824 8020 31858
rect 8054 31824 8092 31858
rect 8126 31824 8164 31858
rect 8198 31824 8236 31858
rect 8270 31824 8308 31858
rect 8342 31824 8380 31858
rect 8414 31824 8452 31858
rect 8486 31824 8524 31858
rect 8558 31824 8596 31858
rect 8630 31824 8668 31858
rect 8702 31824 8740 31858
rect 8774 31824 8812 31858
rect 8846 31824 8884 31858
rect 8918 31824 8956 31858
rect 8990 31824 9028 31858
rect 9062 31824 9100 31858
rect 9134 31824 9172 31858
rect 9206 31824 9244 31858
rect 9278 31824 9284 31858
rect 7870 31791 9284 31824
rect 7870 31785 7880 31791
rect 7914 31785 8016 31791
rect 8050 31785 8152 31791
rect 8186 31785 8288 31791
rect 8322 31785 8424 31791
rect 8458 31785 8560 31791
rect 7870 31751 7876 31785
rect 7914 31757 7948 31785
rect 7910 31751 7948 31757
rect 7982 31757 8016 31785
rect 7982 31751 8020 31757
rect 8054 31751 8092 31785
rect 8126 31757 8152 31785
rect 8126 31751 8164 31757
rect 8198 31751 8236 31785
rect 8270 31757 8288 31785
rect 8270 31751 8308 31757
rect 8342 31751 8380 31785
rect 8414 31757 8424 31785
rect 8414 31751 8452 31757
rect 8486 31751 8524 31785
rect 8558 31757 8560 31785
rect 8594 31785 8696 31791
rect 8730 31785 8832 31791
rect 8866 31785 8968 31791
rect 9002 31785 9104 31791
rect 9138 31785 9240 31791
rect 9274 31785 9284 31791
rect 8594 31757 8596 31785
rect 8558 31751 8596 31757
rect 8630 31751 8668 31785
rect 8730 31757 8740 31785
rect 8702 31751 8740 31757
rect 8774 31751 8812 31785
rect 8866 31757 8884 31785
rect 8846 31751 8884 31757
rect 8918 31751 8956 31785
rect 9002 31757 9028 31785
rect 8990 31751 9028 31757
rect 9062 31751 9100 31785
rect 9138 31757 9172 31785
rect 9134 31751 9172 31757
rect 9206 31757 9240 31785
rect 9206 31751 9244 31757
rect 9278 31751 9284 31785
rect 7870 31712 9284 31751
rect 7870 31678 7876 31712
rect 7910 31678 7948 31712
rect 7982 31678 8020 31712
rect 8054 31678 8092 31712
rect 8126 31678 8164 31712
rect 8198 31678 8236 31712
rect 8270 31678 8308 31712
rect 8342 31678 8380 31712
rect 8414 31678 8452 31712
rect 8486 31678 8524 31712
rect 8558 31678 8596 31712
rect 8630 31678 8668 31712
rect 8702 31678 8740 31712
rect 8774 31678 8812 31712
rect 8846 31678 8884 31712
rect 8918 31678 8956 31712
rect 8990 31678 9028 31712
rect 9062 31678 9100 31712
rect 9134 31678 9172 31712
rect 9206 31678 9244 31712
rect 9278 31678 9284 31712
rect 7870 31655 9284 31678
rect 7870 31639 7880 31655
rect 7914 31639 8016 31655
rect 8050 31639 8152 31655
rect 8186 31639 8288 31655
rect 8322 31639 8424 31655
rect 8458 31639 8560 31655
rect 7870 31605 7876 31639
rect 7914 31621 7948 31639
rect 7910 31605 7948 31621
rect 7982 31621 8016 31639
rect 7982 31605 8020 31621
rect 8054 31605 8092 31639
rect 8126 31621 8152 31639
rect 8126 31605 8164 31621
rect 8198 31605 8236 31639
rect 8270 31621 8288 31639
rect 8270 31605 8308 31621
rect 8342 31605 8380 31639
rect 8414 31621 8424 31639
rect 8414 31605 8452 31621
rect 8486 31605 8524 31639
rect 8558 31621 8560 31639
rect 8594 31639 8696 31655
rect 8730 31639 8832 31655
rect 8866 31639 8968 31655
rect 9002 31639 9104 31655
rect 9138 31639 9240 31655
rect 9274 31639 9284 31655
rect 8594 31621 8596 31639
rect 8558 31605 8596 31621
rect 8630 31605 8668 31639
rect 8730 31621 8740 31639
rect 8702 31605 8740 31621
rect 8774 31605 8812 31639
rect 8866 31621 8884 31639
rect 8846 31605 8884 31621
rect 8918 31605 8956 31639
rect 9002 31621 9028 31639
rect 8990 31605 9028 31621
rect 9062 31605 9100 31639
rect 9138 31621 9172 31639
rect 9134 31605 9172 31621
rect 9206 31621 9240 31639
rect 9206 31605 9244 31621
rect 9278 31605 9284 31639
rect 7870 31566 9284 31605
rect 7870 31532 7876 31566
rect 7910 31532 7948 31566
rect 7982 31532 8020 31566
rect 8054 31532 8092 31566
rect 8126 31532 8164 31566
rect 8198 31532 8236 31566
rect 8270 31532 8308 31566
rect 8342 31532 8380 31566
rect 8414 31532 8452 31566
rect 8486 31532 8524 31566
rect 8558 31532 8596 31566
rect 8630 31532 8668 31566
rect 8702 31532 8740 31566
rect 8774 31532 8812 31566
rect 8846 31532 8884 31566
rect 8918 31532 8956 31566
rect 8990 31532 9028 31566
rect 9062 31532 9100 31566
rect 9134 31532 9172 31566
rect 9206 31532 9244 31566
rect 9278 31532 9284 31566
rect 7870 31519 9284 31532
rect 7870 31493 7880 31519
rect 7914 31493 8016 31519
rect 8050 31493 8152 31519
rect 8186 31493 8288 31519
rect 8322 31493 8424 31519
rect 8458 31493 8560 31519
rect 7870 31459 7876 31493
rect 7914 31485 7948 31493
rect 7910 31459 7948 31485
rect 7982 31485 8016 31493
rect 7982 31459 8020 31485
rect 8054 31459 8092 31493
rect 8126 31485 8152 31493
rect 8126 31459 8164 31485
rect 8198 31459 8236 31493
rect 8270 31485 8288 31493
rect 8270 31459 8308 31485
rect 8342 31459 8380 31493
rect 8414 31485 8424 31493
rect 8414 31459 8452 31485
rect 8486 31459 8524 31493
rect 8558 31485 8560 31493
rect 8594 31493 8696 31519
rect 8730 31493 8832 31519
rect 8866 31493 8968 31519
rect 9002 31493 9104 31519
rect 9138 31493 9240 31519
rect 9274 31493 9284 31519
rect 8594 31485 8596 31493
rect 8558 31459 8596 31485
rect 8630 31459 8668 31493
rect 8730 31485 8740 31493
rect 8702 31459 8740 31485
rect 8774 31459 8812 31493
rect 8866 31485 8884 31493
rect 8846 31459 8884 31485
rect 8918 31459 8956 31493
rect 9002 31485 9028 31493
rect 8990 31459 9028 31485
rect 9062 31459 9100 31493
rect 9138 31485 9172 31493
rect 9134 31459 9172 31485
rect 9206 31485 9240 31493
rect 9206 31459 9244 31485
rect 9278 31459 9284 31493
rect 7870 31420 9284 31459
rect 7870 31386 7876 31420
rect 7910 31386 7948 31420
rect 7982 31386 8020 31420
rect 8054 31386 8092 31420
rect 8126 31386 8164 31420
rect 8198 31386 8236 31420
rect 8270 31386 8308 31420
rect 8342 31386 8380 31420
rect 8414 31386 8452 31420
rect 8486 31386 8524 31420
rect 8558 31386 8596 31420
rect 8630 31386 8668 31420
rect 8702 31386 8740 31420
rect 8774 31386 8812 31420
rect 8846 31386 8884 31420
rect 8918 31386 8956 31420
rect 8990 31386 9028 31420
rect 9062 31386 9100 31420
rect 9134 31386 9172 31420
rect 9206 31386 9244 31420
rect 9278 31386 9284 31420
rect 7870 31383 9284 31386
rect 7870 31349 7880 31383
rect 7914 31349 8016 31383
rect 8050 31349 8152 31383
rect 8186 31349 8288 31383
rect 8322 31349 8424 31383
rect 8458 31349 8560 31383
rect 8594 31349 8696 31383
rect 8730 31349 8832 31383
rect 8866 31349 8968 31383
rect 9002 31349 9104 31383
rect 9138 31349 9240 31383
rect 9274 31349 9284 31383
rect 7870 31347 9284 31349
rect 7870 31313 7876 31347
rect 7910 31313 7948 31347
rect 7982 31313 8020 31347
rect 8054 31313 8092 31347
rect 8126 31313 8164 31347
rect 8198 31313 8236 31347
rect 8270 31313 8308 31347
rect 8342 31313 8380 31347
rect 8414 31313 8452 31347
rect 8486 31313 8524 31347
rect 8558 31313 8596 31347
rect 8630 31313 8668 31347
rect 8702 31313 8740 31347
rect 8774 31313 8812 31347
rect 8846 31313 8884 31347
rect 8918 31313 8956 31347
rect 8990 31313 9028 31347
rect 9062 31313 9100 31347
rect 9134 31313 9172 31347
rect 9206 31313 9244 31347
rect 9278 31313 9284 31347
rect 7870 31274 9284 31313
rect 7870 31240 7876 31274
rect 7910 31247 7948 31274
rect 7914 31240 7948 31247
rect 7982 31247 8020 31274
rect 7982 31240 8016 31247
rect 8054 31240 8092 31274
rect 8126 31247 8164 31274
rect 8126 31240 8152 31247
rect 8198 31240 8236 31274
rect 8270 31247 8308 31274
rect 8270 31240 8288 31247
rect 8342 31240 8380 31274
rect 8414 31247 8452 31274
rect 8414 31240 8424 31247
rect 8486 31240 8524 31274
rect 8558 31247 8596 31274
rect 8558 31240 8560 31247
rect 7870 31213 7880 31240
rect 7914 31213 8016 31240
rect 8050 31213 8152 31240
rect 8186 31213 8288 31240
rect 8322 31213 8424 31240
rect 8458 31213 8560 31240
rect 8594 31240 8596 31247
rect 8630 31240 8668 31274
rect 8702 31247 8740 31274
rect 8730 31240 8740 31247
rect 8774 31240 8812 31274
rect 8846 31247 8884 31274
rect 8866 31240 8884 31247
rect 8918 31240 8956 31274
rect 8990 31247 9028 31274
rect 9002 31240 9028 31247
rect 9062 31240 9100 31274
rect 9134 31247 9172 31274
rect 9138 31240 9172 31247
rect 9206 31247 9244 31274
rect 9206 31240 9240 31247
rect 9278 31240 9284 31274
rect 8594 31213 8696 31240
rect 8730 31213 8832 31240
rect 8866 31213 8968 31240
rect 9002 31213 9104 31240
rect 9138 31213 9240 31240
rect 9274 31213 9284 31240
rect 7870 31201 9284 31213
rect 7870 31167 7876 31201
rect 7910 31167 7948 31201
rect 7982 31167 8020 31201
rect 8054 31167 8092 31201
rect 8126 31167 8164 31201
rect 8198 31167 8236 31201
rect 8270 31167 8308 31201
rect 8342 31167 8380 31201
rect 8414 31167 8452 31201
rect 8486 31167 8524 31201
rect 8558 31167 8596 31201
rect 8630 31167 8668 31201
rect 8702 31167 8740 31201
rect 8774 31167 8812 31201
rect 8846 31167 8884 31201
rect 8918 31167 8956 31201
rect 8990 31167 9028 31201
rect 9062 31167 9100 31201
rect 9134 31167 9172 31201
rect 9206 31167 9244 31201
rect 9278 31167 9284 31201
rect 7870 31128 9284 31167
rect 7870 31094 7876 31128
rect 7910 31111 7948 31128
rect 7914 31094 7948 31111
rect 7982 31111 8020 31128
rect 7982 31094 8016 31111
rect 8054 31094 8092 31128
rect 8126 31111 8164 31128
rect 8126 31094 8152 31111
rect 8198 31094 8236 31128
rect 8270 31111 8308 31128
rect 8270 31094 8288 31111
rect 8342 31094 8380 31128
rect 8414 31111 8452 31128
rect 8414 31094 8424 31111
rect 8486 31094 8524 31128
rect 8558 31111 8596 31128
rect 8558 31094 8560 31111
rect 7870 31077 7880 31094
rect 7914 31077 8016 31094
rect 8050 31077 8152 31094
rect 8186 31077 8288 31094
rect 8322 31077 8424 31094
rect 8458 31077 8560 31094
rect 8594 31094 8596 31111
rect 8630 31094 8668 31128
rect 8702 31111 8740 31128
rect 8730 31094 8740 31111
rect 8774 31094 8812 31128
rect 8846 31111 8884 31128
rect 8866 31094 8884 31111
rect 8918 31094 8956 31128
rect 8990 31111 9028 31128
rect 9002 31094 9028 31111
rect 9062 31094 9100 31128
rect 9134 31111 9172 31128
rect 9138 31094 9172 31111
rect 9206 31111 9244 31128
rect 9206 31094 9240 31111
rect 9278 31094 9284 31128
rect 8594 31077 8696 31094
rect 8730 31077 8832 31094
rect 8866 31077 8968 31094
rect 9002 31077 9104 31094
rect 9138 31077 9240 31094
rect 9274 31077 9284 31094
rect 7870 31055 9284 31077
rect 7870 31021 7876 31055
rect 7910 31021 7948 31055
rect 7982 31021 8020 31055
rect 8054 31021 8092 31055
rect 8126 31021 8164 31055
rect 8198 31021 8236 31055
rect 8270 31021 8308 31055
rect 8342 31021 8380 31055
rect 8414 31021 8452 31055
rect 8486 31021 8524 31055
rect 8558 31021 8596 31055
rect 8630 31021 8668 31055
rect 8702 31021 8740 31055
rect 8774 31021 8812 31055
rect 8846 31021 8884 31055
rect 8918 31021 8956 31055
rect 8990 31021 9028 31055
rect 9062 31021 9100 31055
rect 9134 31021 9172 31055
rect 9206 31021 9244 31055
rect 9278 31021 9284 31055
rect 7870 30982 9284 31021
rect 7870 30948 7876 30982
rect 7910 30975 7948 30982
rect 7914 30948 7948 30975
rect 7982 30975 8020 30982
rect 7982 30948 8016 30975
rect 8054 30948 8092 30982
rect 8126 30975 8164 30982
rect 8126 30948 8152 30975
rect 8198 30948 8236 30982
rect 8270 30975 8308 30982
rect 8270 30948 8288 30975
rect 8342 30948 8380 30982
rect 8414 30975 8452 30982
rect 8414 30948 8424 30975
rect 8486 30948 8524 30982
rect 8558 30975 8596 30982
rect 8558 30948 8560 30975
rect 7870 30941 7880 30948
rect 7914 30941 8016 30948
rect 8050 30941 8152 30948
rect 8186 30941 8288 30948
rect 8322 30941 8424 30948
rect 8458 30941 8560 30948
rect 8594 30948 8596 30975
rect 8630 30948 8668 30982
rect 8702 30975 8740 30982
rect 8730 30948 8740 30975
rect 8774 30948 8812 30982
rect 8846 30975 8884 30982
rect 8866 30948 8884 30975
rect 8918 30948 8956 30982
rect 8990 30975 9028 30982
rect 9002 30948 9028 30975
rect 9062 30948 9100 30982
rect 9134 30975 9172 30982
rect 9138 30948 9172 30975
rect 9206 30975 9244 30982
rect 9206 30948 9240 30975
rect 9278 30948 9284 30982
rect 8594 30941 8696 30948
rect 8730 30941 8832 30948
rect 8866 30941 8968 30948
rect 9002 30941 9104 30948
rect 9138 30941 9240 30948
rect 9274 30941 9284 30948
rect 7870 30909 9284 30941
rect 7870 30875 7876 30909
rect 7910 30875 7948 30909
rect 7982 30875 8020 30909
rect 8054 30875 8092 30909
rect 8126 30875 8164 30909
rect 8198 30875 8236 30909
rect 8270 30875 8308 30909
rect 8342 30875 8380 30909
rect 8414 30875 8452 30909
rect 8486 30875 8524 30909
rect 8558 30875 8596 30909
rect 8630 30875 8668 30909
rect 8702 30875 8740 30909
rect 8774 30875 8812 30909
rect 8846 30875 8884 30909
rect 8918 30875 8956 30909
rect 8990 30875 9028 30909
rect 9062 30875 9100 30909
rect 9134 30875 9172 30909
rect 9206 30875 9244 30909
rect 9278 30875 9284 30909
rect 7870 30839 9284 30875
rect 7870 30836 7880 30839
rect 7914 30836 8016 30839
rect 8050 30836 8152 30839
rect 8186 30836 8288 30839
rect 8322 30836 8424 30839
rect 8458 30836 8560 30839
rect 7870 30802 7876 30836
rect 7914 30805 7948 30836
rect 7910 30802 7948 30805
rect 7982 30805 8016 30836
rect 7982 30802 8020 30805
rect 8054 30802 8092 30836
rect 8126 30805 8152 30836
rect 8126 30802 8164 30805
rect 8198 30802 8236 30836
rect 8270 30805 8288 30836
rect 8270 30802 8308 30805
rect 8342 30802 8380 30836
rect 8414 30805 8424 30836
rect 8414 30802 8452 30805
rect 8486 30802 8524 30836
rect 8558 30805 8560 30836
rect 8594 30836 8696 30839
rect 8730 30836 8832 30839
rect 8866 30836 8968 30839
rect 9002 30836 9104 30839
rect 9138 30836 9240 30839
rect 9274 30836 9284 30839
rect 8594 30805 8596 30836
rect 8558 30802 8596 30805
rect 8630 30802 8668 30836
rect 8730 30805 8740 30836
rect 8702 30802 8740 30805
rect 8774 30802 8812 30836
rect 8866 30805 8884 30836
rect 8846 30802 8884 30805
rect 8918 30802 8956 30836
rect 9002 30805 9028 30836
rect 8990 30802 9028 30805
rect 9062 30802 9100 30836
rect 9138 30805 9172 30836
rect 9134 30802 9172 30805
rect 9206 30805 9240 30836
rect 9206 30802 9244 30805
rect 9278 30802 9284 30836
rect 7870 30763 9284 30802
rect 7870 30729 7876 30763
rect 7910 30729 7948 30763
rect 7982 30729 8020 30763
rect 8054 30729 8092 30763
rect 8126 30729 8164 30763
rect 8198 30729 8236 30763
rect 8270 30729 8308 30763
rect 8342 30729 8380 30763
rect 8414 30729 8452 30763
rect 8486 30729 8524 30763
rect 8558 30729 8596 30763
rect 8630 30729 8668 30763
rect 8702 30729 8740 30763
rect 8774 30729 8812 30763
rect 8846 30729 8884 30763
rect 8918 30729 8956 30763
rect 8990 30729 9028 30763
rect 9062 30729 9100 30763
rect 9134 30729 9172 30763
rect 9206 30729 9244 30763
rect 9278 30729 9284 30763
rect 7870 30703 9284 30729
rect 7870 30690 7880 30703
rect 7914 30690 8016 30703
rect 8050 30690 8152 30703
rect 8186 30690 8288 30703
rect 8322 30690 8424 30703
rect 8458 30690 8560 30703
rect 7870 30656 7876 30690
rect 7914 30669 7948 30690
rect 7910 30656 7948 30669
rect 7982 30669 8016 30690
rect 7982 30656 8020 30669
rect 8054 30656 8092 30690
rect 8126 30669 8152 30690
rect 8126 30656 8164 30669
rect 8198 30656 8236 30690
rect 8270 30669 8288 30690
rect 8270 30656 8308 30669
rect 8342 30656 8380 30690
rect 8414 30669 8424 30690
rect 8414 30656 8452 30669
rect 8486 30656 8524 30690
rect 8558 30669 8560 30690
rect 8594 30690 8696 30703
rect 8730 30690 8832 30703
rect 8866 30690 8968 30703
rect 9002 30690 9104 30703
rect 9138 30690 9240 30703
rect 9274 30690 9284 30703
rect 8594 30669 8596 30690
rect 8558 30656 8596 30669
rect 8630 30656 8668 30690
rect 8730 30669 8740 30690
rect 8702 30656 8740 30669
rect 8774 30656 8812 30690
rect 8866 30669 8884 30690
rect 8846 30656 8884 30669
rect 8918 30656 8956 30690
rect 9002 30669 9028 30690
rect 8990 30656 9028 30669
rect 9062 30656 9100 30690
rect 9138 30669 9172 30690
rect 9134 30656 9172 30669
rect 9206 30669 9240 30690
rect 9206 30656 9244 30669
rect 9278 30656 9284 30690
rect 7870 30617 9284 30656
rect 7870 30583 7876 30617
rect 7910 30583 7948 30617
rect 7982 30583 8020 30617
rect 8054 30583 8092 30617
rect 8126 30583 8164 30617
rect 8198 30583 8236 30617
rect 8270 30583 8308 30617
rect 8342 30583 8380 30617
rect 8414 30583 8452 30617
rect 8486 30583 8524 30617
rect 8558 30583 8596 30617
rect 8630 30583 8668 30617
rect 8702 30583 8740 30617
rect 8774 30583 8812 30617
rect 8846 30583 8884 30617
rect 8918 30583 8956 30617
rect 8990 30583 9028 30617
rect 9062 30583 9100 30617
rect 9134 30583 9172 30617
rect 9206 30583 9244 30617
rect 9278 30583 9284 30617
rect 7870 30567 9284 30583
rect 7870 30544 7880 30567
rect 7914 30544 8016 30567
rect 8050 30544 8152 30567
rect 8186 30544 8288 30567
rect 8322 30544 8424 30567
rect 8458 30544 8560 30567
rect 7870 30510 7876 30544
rect 7914 30533 7948 30544
rect 7910 30510 7948 30533
rect 7982 30533 8016 30544
rect 7982 30510 8020 30533
rect 8054 30510 8092 30544
rect 8126 30533 8152 30544
rect 8126 30510 8164 30533
rect 8198 30510 8236 30544
rect 8270 30533 8288 30544
rect 8270 30510 8308 30533
rect 8342 30510 8380 30544
rect 8414 30533 8424 30544
rect 8414 30510 8452 30533
rect 8486 30510 8524 30544
rect 8558 30533 8560 30544
rect 8594 30544 8696 30567
rect 8730 30544 8832 30567
rect 8866 30544 8968 30567
rect 9002 30544 9104 30567
rect 9138 30544 9240 30567
rect 9274 30544 9284 30567
rect 8594 30533 8596 30544
rect 8558 30510 8596 30533
rect 8630 30510 8668 30544
rect 8730 30533 8740 30544
rect 8702 30510 8740 30533
rect 8774 30510 8812 30544
rect 8866 30533 8884 30544
rect 8846 30510 8884 30533
rect 8918 30510 8956 30544
rect 9002 30533 9028 30544
rect 8990 30510 9028 30533
rect 9062 30510 9100 30544
rect 9138 30533 9172 30544
rect 9134 30510 9172 30533
rect 9206 30533 9240 30544
rect 9206 30510 9244 30533
rect 9278 30510 9284 30544
rect 7870 30471 9284 30510
rect 7870 30437 7876 30471
rect 7910 30437 7948 30471
rect 7982 30437 8020 30471
rect 8054 30437 8092 30471
rect 8126 30437 8164 30471
rect 8198 30437 8236 30471
rect 8270 30437 8308 30471
rect 8342 30437 8380 30471
rect 8414 30437 8452 30471
rect 8486 30437 8524 30471
rect 8558 30437 8596 30471
rect 8630 30437 8668 30471
rect 8702 30437 8740 30471
rect 8774 30437 8812 30471
rect 8846 30437 8884 30471
rect 8918 30437 8956 30471
rect 8990 30437 9028 30471
rect 9062 30437 9100 30471
rect 9134 30437 9172 30471
rect 9206 30437 9244 30471
rect 9278 30437 9284 30471
rect 7870 30431 9284 30437
rect 7870 30398 7880 30431
rect 7914 30398 8016 30431
rect 8050 30398 8152 30431
rect 8186 30398 8288 30431
rect 8322 30398 8424 30431
rect 8458 30398 8560 30431
rect 7870 30364 7876 30398
rect 7914 30397 7948 30398
rect 7910 30364 7948 30397
rect 7982 30397 8016 30398
rect 7982 30364 8020 30397
rect 8054 30364 8092 30398
rect 8126 30397 8152 30398
rect 8126 30364 8164 30397
rect 8198 30364 8236 30398
rect 8270 30397 8288 30398
rect 8270 30364 8308 30397
rect 8342 30364 8380 30398
rect 8414 30397 8424 30398
rect 8414 30364 8452 30397
rect 8486 30364 8524 30398
rect 8558 30397 8560 30398
rect 8594 30398 8696 30431
rect 8730 30398 8832 30431
rect 8866 30398 8968 30431
rect 9002 30398 9104 30431
rect 9138 30398 9240 30431
rect 9274 30398 9284 30431
rect 8594 30397 8596 30398
rect 8558 30364 8596 30397
rect 8630 30364 8668 30398
rect 8730 30397 8740 30398
rect 8702 30364 8740 30397
rect 8774 30364 8812 30398
rect 8866 30397 8884 30398
rect 8846 30364 8884 30397
rect 8918 30364 8956 30398
rect 9002 30397 9028 30398
rect 8990 30364 9028 30397
rect 9062 30364 9100 30398
rect 9138 30397 9172 30398
rect 9134 30364 9172 30397
rect 9206 30397 9240 30398
rect 9206 30364 9244 30397
rect 9278 30364 9284 30398
rect 7870 30325 9284 30364
rect 7870 30291 7876 30325
rect 7910 30295 7948 30325
rect 7914 30291 7948 30295
rect 7982 30295 8020 30325
rect 7982 30291 8016 30295
rect 8054 30291 8092 30325
rect 8126 30295 8164 30325
rect 8126 30291 8152 30295
rect 8198 30291 8236 30325
rect 8270 30295 8308 30325
rect 8270 30291 8288 30295
rect 8342 30291 8380 30325
rect 8414 30295 8452 30325
rect 8414 30291 8424 30295
rect 8486 30291 8524 30325
rect 8558 30295 8596 30325
rect 8558 30291 8560 30295
rect 7870 30261 7880 30291
rect 7914 30261 8016 30291
rect 8050 30261 8152 30291
rect 8186 30261 8288 30291
rect 8322 30261 8424 30291
rect 8458 30261 8560 30291
rect 8594 30291 8596 30295
rect 8630 30291 8668 30325
rect 8702 30295 8740 30325
rect 8730 30291 8740 30295
rect 8774 30291 8812 30325
rect 8846 30295 8884 30325
rect 8866 30291 8884 30295
rect 8918 30291 8956 30325
rect 8990 30295 9028 30325
rect 9002 30291 9028 30295
rect 9062 30291 9100 30325
rect 9134 30295 9172 30325
rect 9138 30291 9172 30295
rect 9206 30295 9244 30325
rect 9206 30291 9240 30295
rect 9278 30291 9284 30325
rect 8594 30261 8696 30291
rect 8730 30261 8832 30291
rect 8866 30261 8968 30291
rect 9002 30261 9104 30291
rect 9138 30261 9240 30291
rect 9274 30261 9284 30291
rect 7870 30252 9284 30261
rect 7870 30218 7876 30252
rect 7910 30218 7948 30252
rect 7982 30218 8020 30252
rect 8054 30218 8092 30252
rect 8126 30218 8164 30252
rect 8198 30218 8236 30252
rect 8270 30218 8308 30252
rect 8342 30218 8380 30252
rect 8414 30218 8452 30252
rect 8486 30218 8524 30252
rect 8558 30218 8596 30252
rect 8630 30218 8668 30252
rect 8702 30218 8740 30252
rect 8774 30218 8812 30252
rect 8846 30218 8884 30252
rect 8918 30218 8956 30252
rect 8990 30218 9028 30252
rect 9062 30218 9100 30252
rect 9134 30218 9172 30252
rect 9206 30218 9244 30252
rect 9278 30218 9284 30252
rect 7870 30179 9284 30218
rect 7870 30145 7876 30179
rect 7910 30159 7948 30179
rect 7914 30145 7948 30159
rect 7982 30159 8020 30179
rect 7982 30145 8016 30159
rect 8054 30145 8092 30179
rect 8126 30159 8164 30179
rect 8126 30145 8152 30159
rect 8198 30145 8236 30179
rect 8270 30159 8308 30179
rect 8270 30145 8288 30159
rect 8342 30145 8380 30179
rect 8414 30159 8452 30179
rect 8414 30145 8424 30159
rect 8486 30145 8524 30179
rect 8558 30159 8596 30179
rect 8558 30145 8560 30159
rect 7870 30125 7880 30145
rect 7914 30125 8016 30145
rect 8050 30125 8152 30145
rect 8186 30125 8288 30145
rect 8322 30125 8424 30145
rect 8458 30125 8560 30145
rect 8594 30145 8596 30159
rect 8630 30145 8668 30179
rect 8702 30159 8740 30179
rect 8730 30145 8740 30159
rect 8774 30145 8812 30179
rect 8846 30159 8884 30179
rect 8866 30145 8884 30159
rect 8918 30145 8956 30179
rect 8990 30159 9028 30179
rect 9002 30145 9028 30159
rect 9062 30145 9100 30179
rect 9134 30159 9172 30179
rect 9138 30145 9172 30159
rect 9206 30159 9244 30179
rect 9206 30145 9240 30159
rect 9278 30145 9284 30179
rect 8594 30125 8696 30145
rect 8730 30125 8832 30145
rect 8866 30125 8968 30145
rect 9002 30125 9104 30145
rect 9138 30125 9240 30145
rect 9274 30125 9284 30145
rect 7870 30106 9284 30125
rect 7870 30072 7876 30106
rect 7910 30072 7948 30106
rect 7982 30072 8020 30106
rect 8054 30072 8092 30106
rect 8126 30072 8164 30106
rect 8198 30072 8236 30106
rect 8270 30072 8308 30106
rect 8342 30072 8380 30106
rect 8414 30072 8452 30106
rect 8486 30072 8524 30106
rect 8558 30072 8596 30106
rect 8630 30072 8668 30106
rect 8702 30072 8740 30106
rect 8774 30072 8812 30106
rect 8846 30072 8884 30106
rect 8918 30072 8956 30106
rect 8990 30072 9028 30106
rect 9062 30072 9100 30106
rect 9134 30072 9172 30106
rect 9206 30072 9244 30106
rect 9278 30072 9284 30106
rect 7870 30033 9284 30072
rect 7870 29999 7876 30033
rect 7910 30023 7948 30033
rect 7914 29999 7948 30023
rect 7982 30023 8020 30033
rect 7982 29999 8016 30023
rect 8054 29999 8092 30033
rect 8126 30023 8164 30033
rect 8126 29999 8152 30023
rect 8198 29999 8236 30033
rect 8270 30023 8308 30033
rect 8270 29999 8288 30023
rect 8342 29999 8380 30033
rect 8414 30023 8452 30033
rect 8414 29999 8424 30023
rect 8486 29999 8524 30033
rect 8558 30023 8596 30033
rect 8558 29999 8560 30023
rect 7870 29989 7880 29999
rect 7914 29989 8016 29999
rect 8050 29989 8152 29999
rect 8186 29989 8288 29999
rect 8322 29989 8424 29999
rect 8458 29989 8560 29999
rect 8594 29999 8596 30023
rect 8630 29999 8668 30033
rect 8702 30023 8740 30033
rect 8730 29999 8740 30023
rect 8774 29999 8812 30033
rect 8846 30023 8884 30033
rect 8866 29999 8884 30023
rect 8918 29999 8956 30033
rect 8990 30023 9028 30033
rect 9002 29999 9028 30023
rect 9062 29999 9100 30033
rect 9134 30023 9172 30033
rect 9138 29999 9172 30023
rect 9206 30023 9244 30033
rect 9206 29999 9240 30023
rect 9278 29999 9284 30033
rect 8594 29989 8696 29999
rect 8730 29989 8832 29999
rect 8866 29989 8968 29999
rect 9002 29989 9104 29999
rect 9138 29989 9240 29999
rect 9274 29989 9284 29999
rect 7870 29960 9284 29989
rect 7870 29926 7876 29960
rect 7910 29926 7948 29960
rect 7982 29926 8020 29960
rect 8054 29926 8092 29960
rect 8126 29926 8164 29960
rect 8198 29926 8236 29960
rect 8270 29926 8308 29960
rect 8342 29926 8380 29960
rect 8414 29926 8452 29960
rect 8486 29926 8524 29960
rect 8558 29926 8596 29960
rect 8630 29926 8668 29960
rect 8702 29926 8740 29960
rect 8774 29926 8812 29960
rect 8846 29926 8884 29960
rect 8918 29926 8956 29960
rect 8990 29926 9028 29960
rect 9062 29926 9100 29960
rect 9134 29926 9172 29960
rect 9206 29926 9244 29960
rect 9278 29926 9284 29960
rect 7870 29887 9284 29926
rect 7870 29853 7876 29887
rect 7914 29853 7948 29887
rect 7982 29853 8016 29887
rect 8054 29853 8092 29887
rect 8126 29853 8152 29887
rect 8198 29853 8236 29887
rect 8270 29853 8288 29887
rect 8342 29853 8380 29887
rect 8414 29853 8424 29887
rect 8486 29853 8524 29887
rect 8558 29853 8560 29887
rect 8594 29853 8596 29887
rect 8630 29853 8668 29887
rect 8730 29853 8740 29887
rect 8774 29853 8812 29887
rect 8866 29853 8884 29887
rect 8918 29853 8956 29887
rect 9002 29853 9028 29887
rect 9062 29853 9100 29887
rect 9138 29853 9172 29887
rect 9206 29853 9240 29887
rect 9278 29853 9284 29887
rect 7870 29814 9284 29853
rect 7870 29780 7876 29814
rect 7910 29780 7948 29814
rect 7982 29780 8020 29814
rect 8054 29780 8092 29814
rect 8126 29780 8164 29814
rect 8198 29780 8236 29814
rect 8270 29780 8308 29814
rect 8342 29780 8380 29814
rect 8414 29780 8452 29814
rect 8486 29780 8524 29814
rect 8558 29780 8596 29814
rect 8630 29780 8668 29814
rect 8702 29780 8740 29814
rect 8774 29780 8812 29814
rect 8846 29780 8884 29814
rect 8918 29780 8956 29814
rect 8990 29780 9028 29814
rect 9062 29780 9100 29814
rect 9134 29780 9172 29814
rect 9206 29780 9244 29814
rect 9278 29780 9284 29814
rect 7870 29751 9284 29780
rect 7870 29741 7880 29751
rect 7914 29741 8016 29751
rect 8050 29741 8152 29751
rect 8186 29741 8288 29751
rect 8322 29741 8424 29751
rect 8458 29741 8560 29751
rect 7870 29707 7876 29741
rect 7914 29717 7948 29741
rect 7910 29707 7948 29717
rect 7982 29717 8016 29741
rect 7982 29707 8020 29717
rect 8054 29707 8092 29741
rect 8126 29717 8152 29741
rect 8126 29707 8164 29717
rect 8198 29707 8236 29741
rect 8270 29717 8288 29741
rect 8270 29707 8308 29717
rect 8342 29707 8380 29741
rect 8414 29717 8424 29741
rect 8414 29707 8452 29717
rect 8486 29707 8524 29741
rect 8558 29717 8560 29741
rect 8594 29741 8696 29751
rect 8730 29741 8832 29751
rect 8866 29741 8968 29751
rect 9002 29741 9104 29751
rect 9138 29741 9240 29751
rect 9274 29741 9284 29751
rect 8594 29717 8596 29741
rect 8558 29707 8596 29717
rect 8630 29707 8668 29741
rect 8730 29717 8740 29741
rect 8702 29707 8740 29717
rect 8774 29707 8812 29741
rect 8866 29717 8884 29741
rect 8846 29707 8884 29717
rect 8918 29707 8956 29741
rect 9002 29717 9028 29741
rect 8990 29707 9028 29717
rect 9062 29707 9100 29741
rect 9138 29717 9172 29741
rect 9134 29707 9172 29717
rect 9206 29717 9240 29741
rect 9206 29707 9244 29717
rect 9278 29707 9284 29741
rect 7870 29668 9284 29707
rect 7870 29634 7876 29668
rect 7910 29634 7948 29668
rect 7982 29634 8020 29668
rect 8054 29634 8092 29668
rect 8126 29634 8164 29668
rect 8198 29634 8236 29668
rect 8270 29634 8308 29668
rect 8342 29634 8380 29668
rect 8414 29634 8452 29668
rect 8486 29634 8524 29668
rect 8558 29634 8596 29668
rect 8630 29634 8668 29668
rect 8702 29634 8740 29668
rect 8774 29634 8812 29668
rect 8846 29634 8884 29668
rect 8918 29634 8956 29668
rect 8990 29634 9028 29668
rect 9062 29634 9100 29668
rect 9134 29634 9172 29668
rect 9206 29634 9244 29668
rect 9278 29634 9284 29668
rect 7870 29615 9284 29634
rect 7870 29602 7880 29615
rect 325 29543 1719 29581
rect 315 29511 1719 29543
rect 315 3125 321 29511
rect 1003 29479 1719 29511
rect 1003 29445 1005 29479
rect 1039 29445 1141 29479
rect 1175 29445 1277 29479
rect 1311 29445 1413 29479
rect 1447 29445 1549 29479
rect 1583 29445 1685 29479
rect 1003 29343 1719 29445
rect 1003 29309 1005 29343
rect 1039 29309 1141 29343
rect 1175 29309 1277 29343
rect 1311 29309 1413 29343
rect 1447 29309 1549 29343
rect 1583 29309 1685 29343
rect 1003 29207 1719 29309
rect 1003 29173 1005 29207
rect 1039 29173 1141 29207
rect 1175 29173 1277 29207
rect 1311 29173 1413 29207
rect 1447 29173 1549 29207
rect 1583 29173 1685 29207
rect 1003 29071 1719 29173
rect 1003 29037 1005 29071
rect 1039 29037 1141 29071
rect 1175 29037 1277 29071
rect 1311 29037 1413 29071
rect 1447 29037 1549 29071
rect 1583 29037 1685 29071
rect 1003 28935 1719 29037
rect 1003 28901 1005 28935
rect 1039 28901 1141 28935
rect 1175 28901 1277 28935
rect 1311 28901 1413 28935
rect 1447 28901 1549 28935
rect 1583 28901 1685 28935
rect 1003 28799 1719 28901
rect 1003 28765 1005 28799
rect 1039 28765 1141 28799
rect 1175 28765 1277 28799
rect 1311 28765 1413 28799
rect 1447 28765 1549 28799
rect 1583 28765 1685 28799
rect 1003 28663 1719 28765
rect 1003 28629 1005 28663
rect 1039 28629 1141 28663
rect 1175 28629 1277 28663
rect 1311 28629 1413 28663
rect 1447 28629 1549 28663
rect 1583 28629 1685 28663
rect 1003 28527 1719 28629
rect 1003 28493 1005 28527
rect 1039 28493 1141 28527
rect 1175 28493 1277 28527
rect 1311 28493 1413 28527
rect 1447 28493 1549 28527
rect 1583 28493 1685 28527
rect 1003 28391 1719 28493
rect 1003 28357 1005 28391
rect 1039 28357 1141 28391
rect 1175 28357 1277 28391
rect 1311 28357 1413 28391
rect 1447 28357 1549 28391
rect 1583 28357 1685 28391
rect 1003 28255 1719 28357
rect 1003 28221 1005 28255
rect 1039 28221 1141 28255
rect 1175 28221 1277 28255
rect 1311 28221 1413 28255
rect 1447 28221 1549 28255
rect 1583 28221 1685 28255
rect 1003 28119 1719 28221
rect 1003 28085 1005 28119
rect 1039 28085 1141 28119
rect 1175 28085 1277 28119
rect 1311 28085 1413 28119
rect 1447 28085 1549 28119
rect 1583 28085 1685 28119
rect 1003 27983 1719 28085
rect 1003 27949 1005 27983
rect 1039 27949 1141 27983
rect 1175 27949 1277 27983
rect 1311 27949 1413 27983
rect 1447 27949 1549 27983
rect 1583 27949 1685 27983
rect 1003 27847 1719 27949
rect 1003 27813 1005 27847
rect 1039 27813 1141 27847
rect 1175 27813 1277 27847
rect 1311 27813 1413 27847
rect 1447 27813 1549 27847
rect 1583 27813 1685 27847
rect 1003 27711 1719 27813
rect 1003 27677 1005 27711
rect 1039 27677 1141 27711
rect 1175 27677 1277 27711
rect 1311 27677 1413 27711
rect 1447 27677 1549 27711
rect 1583 27677 1685 27711
rect 1003 27575 1719 27677
rect 1003 27541 1005 27575
rect 1039 27541 1141 27575
rect 1175 27541 1277 27575
rect 1311 27541 1413 27575
rect 1447 27541 1549 27575
rect 1583 27541 1685 27575
rect 1003 27439 1719 27541
rect 1003 27405 1005 27439
rect 1039 27405 1141 27439
rect 1175 27405 1277 27439
rect 1311 27405 1413 27439
rect 1447 27405 1549 27439
rect 1583 27405 1685 27439
rect 1003 27303 1719 27405
rect 1003 27269 1005 27303
rect 1039 27269 1141 27303
rect 1175 27269 1277 27303
rect 1311 27269 1413 27303
rect 1447 27269 1549 27303
rect 1583 27269 1685 27303
rect 1003 27167 1719 27269
rect 1003 27133 1005 27167
rect 1039 27133 1141 27167
rect 1175 27133 1277 27167
rect 1311 27133 1413 27167
rect 1447 27133 1549 27167
rect 1583 27133 1685 27167
rect 1003 27031 1719 27133
rect 1003 26997 1005 27031
rect 1039 26997 1141 27031
rect 1175 26997 1277 27031
rect 1311 26997 1413 27031
rect 1447 26997 1549 27031
rect 1583 26997 1685 27031
rect 1003 26895 1719 26997
rect 1003 26861 1005 26895
rect 1039 26861 1141 26895
rect 1175 26861 1277 26895
rect 1311 26861 1413 26895
rect 1447 26861 1549 26895
rect 1583 26861 1685 26895
rect 1003 26759 1719 26861
rect 1003 26725 1005 26759
rect 1039 26725 1141 26759
rect 1175 26725 1277 26759
rect 1311 26725 1413 26759
rect 1447 26725 1549 26759
rect 1583 26725 1685 26759
rect 1003 26623 1719 26725
rect 1003 26589 1005 26623
rect 1039 26589 1141 26623
rect 1175 26589 1277 26623
rect 1311 26589 1413 26623
rect 1447 26589 1549 26623
rect 1583 26589 1685 26623
rect 1003 26487 1719 26589
rect 1003 26453 1005 26487
rect 1039 26453 1141 26487
rect 1175 26453 1277 26487
rect 1311 26453 1413 26487
rect 1447 26453 1549 26487
rect 1583 26453 1685 26487
rect 1003 26351 1719 26453
rect 1003 26317 1005 26351
rect 1039 26317 1141 26351
rect 1175 26317 1277 26351
rect 1311 26317 1413 26351
rect 1447 26317 1549 26351
rect 1583 26317 1685 26351
rect 1003 26215 1719 26317
rect 1003 26181 1005 26215
rect 1039 26181 1141 26215
rect 1175 26181 1277 26215
rect 1311 26181 1413 26215
rect 1447 26181 1549 26215
rect 1583 26181 1685 26215
rect 1003 26079 1719 26181
rect 1003 26045 1005 26079
rect 1039 26045 1141 26079
rect 1175 26045 1277 26079
rect 1311 26045 1413 26079
rect 1447 26045 1549 26079
rect 1583 26045 1685 26079
rect 1003 25943 1719 26045
rect 1003 25909 1005 25943
rect 1039 25909 1141 25943
rect 1175 25909 1277 25943
rect 1311 25909 1413 25943
rect 1447 25909 1549 25943
rect 1583 25909 1685 25943
rect 1003 25807 1719 25909
rect 1003 25773 1005 25807
rect 1039 25773 1141 25807
rect 1175 25773 1277 25807
rect 1311 25773 1413 25807
rect 1447 25773 1549 25807
rect 1583 25773 1685 25807
rect 1003 25671 1719 25773
rect 1003 25637 1005 25671
rect 1039 25637 1141 25671
rect 1175 25637 1277 25671
rect 1311 25637 1413 25671
rect 1447 25637 1549 25671
rect 1583 25637 1685 25671
rect 1003 25535 1719 25637
rect 1003 25501 1005 25535
rect 1039 25501 1141 25535
rect 1175 25501 1277 25535
rect 1311 25501 1413 25535
rect 1447 25501 1549 25535
rect 1583 25501 1685 25535
rect 1003 25399 1719 25501
rect 1003 25365 1005 25399
rect 1039 25365 1141 25399
rect 1175 25365 1277 25399
rect 1311 25365 1413 25399
rect 1447 25365 1549 25399
rect 1583 25365 1685 25399
rect 1003 25263 1719 25365
rect 1003 25229 1005 25263
rect 1039 25229 1141 25263
rect 1175 25229 1277 25263
rect 1311 25229 1413 25263
rect 1447 25229 1549 25263
rect 1583 25229 1685 25263
rect 1003 25127 1719 25229
rect 1003 25093 1005 25127
rect 1039 25093 1141 25127
rect 1175 25093 1277 25127
rect 1311 25093 1413 25127
rect 1447 25093 1549 25127
rect 1583 25093 1685 25127
rect 1003 24991 1719 25093
rect 1003 24957 1005 24991
rect 1039 24957 1141 24991
rect 1175 24957 1277 24991
rect 1311 24957 1413 24991
rect 1447 24957 1549 24991
rect 1583 24957 1685 24991
rect 1003 24855 1719 24957
rect 1003 24821 1005 24855
rect 1039 24821 1141 24855
rect 1175 24821 1277 24855
rect 1311 24821 1413 24855
rect 1447 24821 1549 24855
rect 1583 24821 1685 24855
rect 1003 24719 1719 24821
rect 1003 24685 1005 24719
rect 1039 24685 1141 24719
rect 1175 24685 1277 24719
rect 1311 24685 1413 24719
rect 1447 24685 1549 24719
rect 1583 24685 1685 24719
rect 1003 24583 1719 24685
rect 1003 24549 1005 24583
rect 1039 24549 1141 24583
rect 1175 24549 1277 24583
rect 1311 24549 1413 24583
rect 1447 24549 1549 24583
rect 1583 24549 1685 24583
rect 1003 24447 1719 24549
rect 1003 24413 1005 24447
rect 1039 24413 1141 24447
rect 1175 24413 1277 24447
rect 1311 24413 1413 24447
rect 1447 24413 1549 24447
rect 1583 24413 1685 24447
rect 1003 24311 1719 24413
rect 1003 24277 1005 24311
rect 1039 24277 1141 24311
rect 1175 24277 1277 24311
rect 1311 24277 1413 24311
rect 1447 24277 1549 24311
rect 1583 24277 1685 24311
rect 1003 24175 1719 24277
rect 1003 24141 1005 24175
rect 1039 24141 1141 24175
rect 1175 24141 1277 24175
rect 1311 24141 1413 24175
rect 1447 24141 1549 24175
rect 1583 24141 1685 24175
rect 1003 24039 1719 24141
rect 1003 24005 1005 24039
rect 1039 24005 1141 24039
rect 1175 24005 1277 24039
rect 1311 24005 1413 24039
rect 1447 24005 1549 24039
rect 1583 24005 1685 24039
rect 1003 23903 1719 24005
rect 1003 23869 1005 23903
rect 1039 23869 1141 23903
rect 1175 23869 1277 23903
rect 1311 23869 1413 23903
rect 1447 23869 1549 23903
rect 1583 23869 1685 23903
rect 1003 23767 1719 23869
rect 1003 23733 1005 23767
rect 1039 23733 1141 23767
rect 1175 23733 1277 23767
rect 1311 23733 1413 23767
rect 1447 23733 1549 23767
rect 1583 23733 1685 23767
rect 1003 23631 1719 23733
rect 1003 23597 1005 23631
rect 1039 23597 1141 23631
rect 1175 23597 1277 23631
rect 1311 23597 1413 23631
rect 1447 23597 1549 23631
rect 1583 23597 1685 23631
rect 1003 23495 1719 23597
rect 1003 23461 1005 23495
rect 1039 23461 1141 23495
rect 1175 23461 1277 23495
rect 1311 23461 1413 23495
rect 1447 23461 1549 23495
rect 1583 23461 1685 23495
rect 1003 23359 1719 23461
rect 1003 23325 1005 23359
rect 1039 23325 1141 23359
rect 1175 23325 1277 23359
rect 1311 23325 1413 23359
rect 1447 23325 1549 23359
rect 1583 23325 1685 23359
rect 1003 23223 1719 23325
rect 1003 23189 1005 23223
rect 1039 23189 1141 23223
rect 1175 23189 1277 23223
rect 1311 23189 1413 23223
rect 1447 23189 1549 23223
rect 1583 23189 1685 23223
rect 1003 23087 1719 23189
rect 1003 23053 1005 23087
rect 1039 23053 1141 23087
rect 1175 23053 1277 23087
rect 1311 23053 1413 23087
rect 1447 23053 1549 23087
rect 1583 23053 1685 23087
rect 1003 22951 1719 23053
rect 1003 22917 1005 22951
rect 1039 22917 1141 22951
rect 1175 22917 1277 22951
rect 1311 22917 1413 22951
rect 1447 22917 1549 22951
rect 1583 22917 1685 22951
rect 1003 22815 1719 22917
rect 1003 22781 1005 22815
rect 1039 22781 1141 22815
rect 1175 22781 1277 22815
rect 1311 22781 1413 22815
rect 1447 22781 1549 22815
rect 1583 22781 1685 22815
rect 1003 22679 1719 22781
rect 1003 22645 1005 22679
rect 1039 22645 1141 22679
rect 1175 22645 1277 22679
rect 1311 22645 1413 22679
rect 1447 22645 1549 22679
rect 1583 22645 1685 22679
rect 1003 22543 1719 22645
rect 1003 22509 1005 22543
rect 1039 22509 1141 22543
rect 1175 22509 1277 22543
rect 1311 22509 1413 22543
rect 1447 22509 1549 22543
rect 1583 22509 1685 22543
rect 1003 22407 1719 22509
rect 1003 22373 1005 22407
rect 1039 22373 1141 22407
rect 1175 22373 1277 22407
rect 1311 22373 1413 22407
rect 1447 22373 1549 22407
rect 1583 22373 1685 22407
rect 1003 22271 1719 22373
rect 1003 22237 1005 22271
rect 1039 22237 1141 22271
rect 1175 22237 1277 22271
rect 1311 22237 1413 22271
rect 1447 22237 1549 22271
rect 1583 22237 1685 22271
rect 1003 22135 1719 22237
rect 1003 22101 1005 22135
rect 1039 22101 1141 22135
rect 1175 22101 1277 22135
rect 1311 22101 1413 22135
rect 1447 22101 1549 22135
rect 1583 22101 1685 22135
rect 1003 21999 1719 22101
rect 1003 21965 1005 21999
rect 1039 21965 1141 21999
rect 1175 21965 1277 21999
rect 1311 21965 1413 21999
rect 1447 21965 1549 21999
rect 1583 21965 1685 21999
rect 1003 21863 1719 21965
rect 1003 21829 1005 21863
rect 1039 21829 1141 21863
rect 1175 21829 1277 21863
rect 1311 21829 1413 21863
rect 1447 21829 1549 21863
rect 1583 21829 1685 21863
rect 1003 21727 1719 21829
rect 1003 21693 1005 21727
rect 1039 21693 1141 21727
rect 1175 21693 1277 21727
rect 1311 21693 1413 21727
rect 1447 21693 1549 21727
rect 1583 21693 1685 21727
rect 1003 21591 1719 21693
rect 1003 21557 1005 21591
rect 1039 21557 1141 21591
rect 1175 21557 1277 21591
rect 1311 21557 1413 21591
rect 1447 21557 1549 21591
rect 1583 21557 1685 21591
rect 1003 21455 1719 21557
rect 1003 21421 1005 21455
rect 1039 21421 1141 21455
rect 1175 21421 1277 21455
rect 1311 21421 1413 21455
rect 1447 21421 1549 21455
rect 1583 21421 1685 21455
rect 1003 21319 1719 21421
rect 1003 21285 1005 21319
rect 1039 21285 1141 21319
rect 1175 21285 1277 21319
rect 1311 21285 1413 21319
rect 1447 21285 1549 21319
rect 1583 21285 1685 21319
rect 1003 21183 1719 21285
rect 1003 21149 1005 21183
rect 1039 21149 1141 21183
rect 1175 21149 1277 21183
rect 1311 21149 1413 21183
rect 1447 21149 1549 21183
rect 1583 21149 1685 21183
rect 1003 21047 1719 21149
rect 1003 21013 1005 21047
rect 1039 21013 1141 21047
rect 1175 21013 1277 21047
rect 1311 21013 1413 21047
rect 1447 21013 1549 21047
rect 1583 21013 1685 21047
rect 1003 20911 1719 21013
rect 1003 20877 1005 20911
rect 1039 20877 1141 20911
rect 1175 20877 1277 20911
rect 1311 20877 1413 20911
rect 1447 20877 1549 20911
rect 1583 20877 1685 20911
rect 1003 20775 1719 20877
rect 1003 20741 1005 20775
rect 1039 20741 1141 20775
rect 1175 20741 1277 20775
rect 1311 20741 1413 20775
rect 1447 20741 1549 20775
rect 1583 20741 1685 20775
rect 1003 20639 1719 20741
rect 1003 20605 1005 20639
rect 1039 20605 1141 20639
rect 1175 20605 1277 20639
rect 1311 20605 1413 20639
rect 1447 20605 1549 20639
rect 1583 20605 1685 20639
rect 1003 20503 1719 20605
rect 1003 20469 1005 20503
rect 1039 20469 1141 20503
rect 1175 20469 1277 20503
rect 1311 20469 1413 20503
rect 1447 20469 1549 20503
rect 1583 20469 1685 20503
rect 1003 20367 1719 20469
rect 1003 20333 1005 20367
rect 1039 20333 1141 20367
rect 1175 20333 1277 20367
rect 1311 20333 1413 20367
rect 1447 20333 1549 20367
rect 1583 20333 1685 20367
rect 1003 20231 1719 20333
rect 1003 20197 1005 20231
rect 1039 20197 1141 20231
rect 1175 20197 1277 20231
rect 1311 20197 1413 20231
rect 1447 20197 1549 20231
rect 1583 20197 1685 20231
rect 1003 20095 1719 20197
rect 1003 20061 1005 20095
rect 1039 20061 1141 20095
rect 1175 20061 1277 20095
rect 1311 20061 1413 20095
rect 1447 20061 1549 20095
rect 1583 20061 1685 20095
rect 1003 19959 1719 20061
rect 1003 19925 1005 19959
rect 1039 19925 1141 19959
rect 1175 19925 1277 19959
rect 1311 19925 1413 19959
rect 1447 19925 1549 19959
rect 1583 19925 1685 19959
rect 1003 19823 1719 19925
rect 1003 19789 1005 19823
rect 1039 19789 1141 19823
rect 1175 19789 1277 19823
rect 1311 19789 1413 19823
rect 1447 19789 1549 19823
rect 1583 19789 1685 19823
rect 1003 19687 1719 19789
rect 1003 19653 1005 19687
rect 1039 19653 1141 19687
rect 1175 19653 1277 19687
rect 1311 19653 1413 19687
rect 1447 19653 1549 19687
rect 1583 19653 1685 19687
rect 1003 19551 1719 19653
rect 1003 19517 1005 19551
rect 1039 19517 1141 19551
rect 1175 19517 1277 19551
rect 1311 19517 1413 19551
rect 1447 19517 1549 19551
rect 1583 19517 1685 19551
rect 1003 19415 1719 19517
rect 1003 19381 1005 19415
rect 1039 19381 1141 19415
rect 1175 19381 1277 19415
rect 1311 19381 1413 19415
rect 1447 19381 1549 19415
rect 1583 19381 1685 19415
rect 1003 19279 1719 19381
rect 1003 19245 1005 19279
rect 1039 19245 1141 19279
rect 1175 19245 1277 19279
rect 1311 19245 1413 19279
rect 1447 19245 1549 19279
rect 1583 19245 1685 19279
rect 1003 19143 1719 19245
rect 1003 19109 1005 19143
rect 1039 19109 1141 19143
rect 1175 19109 1277 19143
rect 1311 19109 1413 19143
rect 1447 19109 1549 19143
rect 1583 19109 1685 19143
rect 1003 19007 1719 19109
rect 1003 18973 1005 19007
rect 1039 18973 1141 19007
rect 1175 18973 1277 19007
rect 1311 18973 1413 19007
rect 1447 18973 1549 19007
rect 1583 18973 1685 19007
rect 1003 18871 1719 18973
rect 1003 18837 1005 18871
rect 1039 18837 1141 18871
rect 1175 18837 1277 18871
rect 1311 18837 1413 18871
rect 1447 18837 1549 18871
rect 1583 18837 1685 18871
rect 1003 18735 1719 18837
rect 1003 18701 1005 18735
rect 1039 18701 1141 18735
rect 1175 18701 1277 18735
rect 1311 18701 1413 18735
rect 1447 18701 1549 18735
rect 1583 18701 1685 18735
rect 1003 18599 1719 18701
rect 1003 18565 1005 18599
rect 1039 18565 1141 18599
rect 1175 18565 1277 18599
rect 1311 18565 1413 18599
rect 1447 18565 1549 18599
rect 1583 18565 1685 18599
rect 1003 18463 1719 18565
rect 1003 18429 1005 18463
rect 1039 18429 1141 18463
rect 1175 18429 1277 18463
rect 1311 18429 1413 18463
rect 1447 18429 1549 18463
rect 1583 18429 1685 18463
rect 1003 18327 1719 18429
rect 1003 18293 1005 18327
rect 1039 18293 1141 18327
rect 1175 18293 1277 18327
rect 1311 18293 1413 18327
rect 1447 18293 1549 18327
rect 1583 18293 1685 18327
rect 1003 18191 1719 18293
rect 1003 18157 1005 18191
rect 1039 18157 1141 18191
rect 1175 18157 1277 18191
rect 1311 18157 1413 18191
rect 1447 18157 1549 18191
rect 1583 18157 1685 18191
rect 1003 18055 1719 18157
rect 1003 18021 1005 18055
rect 1039 18021 1141 18055
rect 1175 18021 1277 18055
rect 1311 18021 1413 18055
rect 1447 18021 1549 18055
rect 1583 18021 1685 18055
rect 1003 17919 1719 18021
rect 1003 17885 1005 17919
rect 1039 17885 1141 17919
rect 1175 17885 1277 17919
rect 1311 17885 1413 17919
rect 1447 17885 1549 17919
rect 1583 17885 1685 17919
rect 1003 17783 1719 17885
rect 1003 17749 1005 17783
rect 1039 17749 1141 17783
rect 1175 17749 1277 17783
rect 1311 17749 1413 17783
rect 1447 17749 1549 17783
rect 1583 17749 1685 17783
rect 1003 17647 1719 17749
rect 1003 17613 1005 17647
rect 1039 17613 1141 17647
rect 1175 17613 1277 17647
rect 1311 17613 1413 17647
rect 1447 17613 1549 17647
rect 1583 17613 1685 17647
rect 1003 17511 1719 17613
rect 7914 29581 8016 29615
rect 8050 29581 8152 29615
rect 8186 29581 8288 29615
rect 8322 29581 8424 29615
rect 8458 29581 8560 29615
rect 8594 29581 8696 29615
rect 8730 29581 8832 29615
rect 8866 29581 8968 29615
rect 9002 29581 9104 29615
rect 9138 29581 9240 29615
rect 9274 29602 9284 29615
rect 7880 29543 9274 29581
rect 7880 29511 9284 29543
rect 7880 29479 8596 29511
rect 7914 29445 8016 29479
rect 8050 29445 8152 29479
rect 8186 29445 8288 29479
rect 8322 29445 8424 29479
rect 8458 29445 8560 29479
rect 8594 29445 8596 29479
rect 7880 29343 8596 29445
rect 7914 29309 8016 29343
rect 8050 29309 8152 29343
rect 8186 29309 8288 29343
rect 8322 29309 8424 29343
rect 8458 29309 8560 29343
rect 8594 29309 8596 29343
rect 7880 29207 8596 29309
rect 7914 29173 8016 29207
rect 8050 29173 8152 29207
rect 8186 29173 8288 29207
rect 8322 29173 8424 29207
rect 8458 29173 8560 29207
rect 8594 29173 8596 29207
rect 7880 29071 8596 29173
rect 7914 29037 8016 29071
rect 8050 29037 8152 29071
rect 8186 29037 8288 29071
rect 8322 29037 8424 29071
rect 8458 29037 8560 29071
rect 8594 29037 8596 29071
rect 7880 28935 8596 29037
rect 7914 28901 8016 28935
rect 8050 28901 8152 28935
rect 8186 28901 8288 28935
rect 8322 28901 8424 28935
rect 8458 28901 8560 28935
rect 8594 28901 8596 28935
rect 7880 28799 8596 28901
rect 7914 28765 8016 28799
rect 8050 28765 8152 28799
rect 8186 28765 8288 28799
rect 8322 28765 8424 28799
rect 8458 28765 8560 28799
rect 8594 28765 8596 28799
rect 7880 28663 8596 28765
rect 7914 28629 8016 28663
rect 8050 28629 8152 28663
rect 8186 28629 8288 28663
rect 8322 28629 8424 28663
rect 8458 28629 8560 28663
rect 8594 28629 8596 28663
rect 7880 28527 8596 28629
rect 7914 28493 8016 28527
rect 8050 28493 8152 28527
rect 8186 28493 8288 28527
rect 8322 28493 8424 28527
rect 8458 28493 8560 28527
rect 8594 28493 8596 28527
rect 7880 28391 8596 28493
rect 7914 28357 8016 28391
rect 8050 28357 8152 28391
rect 8186 28357 8288 28391
rect 8322 28357 8424 28391
rect 8458 28357 8560 28391
rect 8594 28357 8596 28391
rect 7880 28255 8596 28357
rect 7914 28221 8016 28255
rect 8050 28221 8152 28255
rect 8186 28221 8288 28255
rect 8322 28221 8424 28255
rect 8458 28221 8560 28255
rect 8594 28221 8596 28255
rect 7880 28119 8596 28221
rect 7914 28085 8016 28119
rect 8050 28085 8152 28119
rect 8186 28085 8288 28119
rect 8322 28085 8424 28119
rect 8458 28085 8560 28119
rect 8594 28085 8596 28119
rect 7880 27983 8596 28085
rect 7914 27949 8016 27983
rect 8050 27949 8152 27983
rect 8186 27949 8288 27983
rect 8322 27949 8424 27983
rect 8458 27949 8560 27983
rect 8594 27949 8596 27983
rect 7880 27847 8596 27949
rect 7914 27813 8016 27847
rect 8050 27813 8152 27847
rect 8186 27813 8288 27847
rect 8322 27813 8424 27847
rect 8458 27813 8560 27847
rect 8594 27813 8596 27847
rect 7880 27711 8596 27813
rect 7914 27677 8016 27711
rect 8050 27677 8152 27711
rect 8186 27677 8288 27711
rect 8322 27677 8424 27711
rect 8458 27677 8560 27711
rect 8594 27677 8596 27711
rect 7880 27575 8596 27677
rect 7914 27541 8016 27575
rect 8050 27541 8152 27575
rect 8186 27541 8288 27575
rect 8322 27541 8424 27575
rect 8458 27541 8560 27575
rect 8594 27541 8596 27575
rect 7880 27439 8596 27541
rect 7914 27405 8016 27439
rect 8050 27405 8152 27439
rect 8186 27405 8288 27439
rect 8322 27405 8424 27439
rect 8458 27405 8560 27439
rect 8594 27405 8596 27439
rect 7880 27303 8596 27405
rect 7914 27269 8016 27303
rect 8050 27269 8152 27303
rect 8186 27269 8288 27303
rect 8322 27269 8424 27303
rect 8458 27269 8560 27303
rect 8594 27269 8596 27303
rect 7880 27167 8596 27269
rect 7914 27133 8016 27167
rect 8050 27133 8152 27167
rect 8186 27133 8288 27167
rect 8322 27133 8424 27167
rect 8458 27133 8560 27167
rect 8594 27133 8596 27167
rect 7880 27031 8596 27133
rect 7914 26997 8016 27031
rect 8050 26997 8152 27031
rect 8186 26997 8288 27031
rect 8322 26997 8424 27031
rect 8458 26997 8560 27031
rect 8594 26997 8596 27031
rect 7880 26895 8596 26997
rect 7914 26861 8016 26895
rect 8050 26861 8152 26895
rect 8186 26861 8288 26895
rect 8322 26861 8424 26895
rect 8458 26861 8560 26895
rect 8594 26861 8596 26895
rect 7880 26759 8596 26861
rect 7914 26725 8016 26759
rect 8050 26725 8152 26759
rect 8186 26725 8288 26759
rect 8322 26725 8424 26759
rect 8458 26725 8560 26759
rect 8594 26725 8596 26759
rect 7880 26623 8596 26725
rect 7914 26589 8016 26623
rect 8050 26589 8152 26623
rect 8186 26589 8288 26623
rect 8322 26589 8424 26623
rect 8458 26589 8560 26623
rect 8594 26589 8596 26623
rect 7880 26487 8596 26589
rect 7914 26453 8016 26487
rect 8050 26453 8152 26487
rect 8186 26453 8288 26487
rect 8322 26453 8424 26487
rect 8458 26453 8560 26487
rect 8594 26453 8596 26487
rect 7880 26351 8596 26453
rect 7914 26317 8016 26351
rect 8050 26317 8152 26351
rect 8186 26317 8288 26351
rect 8322 26317 8424 26351
rect 8458 26317 8560 26351
rect 8594 26317 8596 26351
rect 7880 26215 8596 26317
rect 7914 26181 8016 26215
rect 8050 26181 8152 26215
rect 8186 26181 8288 26215
rect 8322 26181 8424 26215
rect 8458 26181 8560 26215
rect 8594 26181 8596 26215
rect 7880 26079 8596 26181
rect 7914 26045 8016 26079
rect 8050 26045 8152 26079
rect 8186 26045 8288 26079
rect 8322 26045 8424 26079
rect 8458 26045 8560 26079
rect 8594 26045 8596 26079
rect 7880 25943 8596 26045
rect 7914 25909 8016 25943
rect 8050 25909 8152 25943
rect 8186 25909 8288 25943
rect 8322 25909 8424 25943
rect 8458 25909 8560 25943
rect 8594 25909 8596 25943
rect 7880 25807 8596 25909
rect 7914 25773 8016 25807
rect 8050 25773 8152 25807
rect 8186 25773 8288 25807
rect 8322 25773 8424 25807
rect 8458 25773 8560 25807
rect 8594 25773 8596 25807
rect 7880 25671 8596 25773
rect 7914 25637 8016 25671
rect 8050 25637 8152 25671
rect 8186 25637 8288 25671
rect 8322 25637 8424 25671
rect 8458 25637 8560 25671
rect 8594 25637 8596 25671
rect 7880 25535 8596 25637
rect 7914 25501 8016 25535
rect 8050 25501 8152 25535
rect 8186 25501 8288 25535
rect 8322 25501 8424 25535
rect 8458 25501 8560 25535
rect 8594 25501 8596 25535
rect 7880 25399 8596 25501
rect 7914 25365 8016 25399
rect 8050 25365 8152 25399
rect 8186 25365 8288 25399
rect 8322 25365 8424 25399
rect 8458 25365 8560 25399
rect 8594 25365 8596 25399
rect 7880 25263 8596 25365
rect 7914 25229 8016 25263
rect 8050 25229 8152 25263
rect 8186 25229 8288 25263
rect 8322 25229 8424 25263
rect 8458 25229 8560 25263
rect 8594 25229 8596 25263
rect 7880 25127 8596 25229
rect 7914 25093 8016 25127
rect 8050 25093 8152 25127
rect 8186 25093 8288 25127
rect 8322 25093 8424 25127
rect 8458 25093 8560 25127
rect 8594 25093 8596 25127
rect 7880 24991 8596 25093
rect 7914 24957 8016 24991
rect 8050 24957 8152 24991
rect 8186 24957 8288 24991
rect 8322 24957 8424 24991
rect 8458 24957 8560 24991
rect 8594 24957 8596 24991
rect 7880 24855 8596 24957
rect 7914 24821 8016 24855
rect 8050 24821 8152 24855
rect 8186 24821 8288 24855
rect 8322 24821 8424 24855
rect 8458 24821 8560 24855
rect 8594 24821 8596 24855
rect 7880 24719 8596 24821
rect 7914 24685 8016 24719
rect 8050 24685 8152 24719
rect 8186 24685 8288 24719
rect 8322 24685 8424 24719
rect 8458 24685 8560 24719
rect 8594 24685 8596 24719
rect 7880 24583 8596 24685
rect 7914 24549 8016 24583
rect 8050 24549 8152 24583
rect 8186 24549 8288 24583
rect 8322 24549 8424 24583
rect 8458 24549 8560 24583
rect 8594 24549 8596 24583
rect 7880 24447 8596 24549
rect 7914 24413 8016 24447
rect 8050 24413 8152 24447
rect 8186 24413 8288 24447
rect 8322 24413 8424 24447
rect 8458 24413 8560 24447
rect 8594 24413 8596 24447
rect 7880 24311 8596 24413
rect 7914 24277 8016 24311
rect 8050 24277 8152 24311
rect 8186 24277 8288 24311
rect 8322 24277 8424 24311
rect 8458 24277 8560 24311
rect 8594 24277 8596 24311
rect 7880 24175 8596 24277
rect 7914 24141 8016 24175
rect 8050 24141 8152 24175
rect 8186 24141 8288 24175
rect 8322 24141 8424 24175
rect 8458 24141 8560 24175
rect 8594 24141 8596 24175
rect 7880 24039 8596 24141
rect 7914 24005 8016 24039
rect 8050 24005 8152 24039
rect 8186 24005 8288 24039
rect 8322 24005 8424 24039
rect 8458 24005 8560 24039
rect 8594 24005 8596 24039
rect 7880 23903 8596 24005
rect 7914 23869 8016 23903
rect 8050 23869 8152 23903
rect 8186 23869 8288 23903
rect 8322 23869 8424 23903
rect 8458 23869 8560 23903
rect 8594 23869 8596 23903
rect 7880 23767 8596 23869
rect 7914 23733 8016 23767
rect 8050 23733 8152 23767
rect 8186 23733 8288 23767
rect 8322 23733 8424 23767
rect 8458 23733 8560 23767
rect 8594 23733 8596 23767
rect 7880 23631 8596 23733
rect 7914 23597 8016 23631
rect 8050 23597 8152 23631
rect 8186 23597 8288 23631
rect 8322 23597 8424 23631
rect 8458 23597 8560 23631
rect 8594 23597 8596 23631
rect 7880 23495 8596 23597
rect 7914 23461 8016 23495
rect 8050 23461 8152 23495
rect 8186 23461 8288 23495
rect 8322 23461 8424 23495
rect 8458 23461 8560 23495
rect 8594 23461 8596 23495
rect 7880 23359 8596 23461
rect 7914 23325 8016 23359
rect 8050 23325 8152 23359
rect 8186 23325 8288 23359
rect 8322 23325 8424 23359
rect 8458 23325 8560 23359
rect 8594 23325 8596 23359
rect 7880 23223 8596 23325
rect 7914 23189 8016 23223
rect 8050 23189 8152 23223
rect 8186 23189 8288 23223
rect 8322 23189 8424 23223
rect 8458 23189 8560 23223
rect 8594 23189 8596 23223
rect 7880 23087 8596 23189
rect 7914 23053 8016 23087
rect 8050 23053 8152 23087
rect 8186 23053 8288 23087
rect 8322 23053 8424 23087
rect 8458 23053 8560 23087
rect 8594 23053 8596 23087
rect 7880 22951 8596 23053
rect 7914 22917 8016 22951
rect 8050 22917 8152 22951
rect 8186 22917 8288 22951
rect 8322 22917 8424 22951
rect 8458 22917 8560 22951
rect 8594 22917 8596 22951
rect 7880 22815 8596 22917
rect 7914 22781 8016 22815
rect 8050 22781 8152 22815
rect 8186 22781 8288 22815
rect 8322 22781 8424 22815
rect 8458 22781 8560 22815
rect 8594 22781 8596 22815
rect 7880 22679 8596 22781
rect 7914 22645 8016 22679
rect 8050 22645 8152 22679
rect 8186 22645 8288 22679
rect 8322 22645 8424 22679
rect 8458 22645 8560 22679
rect 8594 22645 8596 22679
rect 7880 22543 8596 22645
rect 7914 22509 8016 22543
rect 8050 22509 8152 22543
rect 8186 22509 8288 22543
rect 8322 22509 8424 22543
rect 8458 22509 8560 22543
rect 8594 22509 8596 22543
rect 7880 22407 8596 22509
rect 7914 22373 8016 22407
rect 8050 22373 8152 22407
rect 8186 22373 8288 22407
rect 8322 22373 8424 22407
rect 8458 22373 8560 22407
rect 8594 22373 8596 22407
rect 7880 22271 8596 22373
rect 7914 22237 8016 22271
rect 8050 22237 8152 22271
rect 8186 22237 8288 22271
rect 8322 22237 8424 22271
rect 8458 22237 8560 22271
rect 8594 22237 8596 22271
rect 7880 22135 8596 22237
rect 7914 22101 8016 22135
rect 8050 22101 8152 22135
rect 8186 22101 8288 22135
rect 8322 22101 8424 22135
rect 8458 22101 8560 22135
rect 8594 22101 8596 22135
rect 7880 21999 8596 22101
rect 7914 21965 8016 21999
rect 8050 21965 8152 21999
rect 8186 21965 8288 21999
rect 8322 21965 8424 21999
rect 8458 21965 8560 21999
rect 8594 21965 8596 21999
rect 7880 21863 8596 21965
rect 7914 21829 8016 21863
rect 8050 21829 8152 21863
rect 8186 21829 8288 21863
rect 8322 21829 8424 21863
rect 8458 21829 8560 21863
rect 8594 21829 8596 21863
rect 7880 21727 8596 21829
rect 7914 21693 8016 21727
rect 8050 21693 8152 21727
rect 8186 21693 8288 21727
rect 8322 21693 8424 21727
rect 8458 21693 8560 21727
rect 8594 21693 8596 21727
rect 7880 21591 8596 21693
rect 7914 21557 8016 21591
rect 8050 21557 8152 21591
rect 8186 21557 8288 21591
rect 8322 21557 8424 21591
rect 8458 21557 8560 21591
rect 8594 21557 8596 21591
rect 7880 21455 8596 21557
rect 7914 21421 8016 21455
rect 8050 21421 8152 21455
rect 8186 21421 8288 21455
rect 8322 21421 8424 21455
rect 8458 21421 8560 21455
rect 8594 21421 8596 21455
rect 7880 21319 8596 21421
rect 7914 21285 8016 21319
rect 8050 21285 8152 21319
rect 8186 21285 8288 21319
rect 8322 21285 8424 21319
rect 8458 21285 8560 21319
rect 8594 21285 8596 21319
rect 7880 21183 8596 21285
rect 7914 21149 8016 21183
rect 8050 21149 8152 21183
rect 8186 21149 8288 21183
rect 8322 21149 8424 21183
rect 8458 21149 8560 21183
rect 8594 21149 8596 21183
rect 7880 21047 8596 21149
rect 7914 21013 8016 21047
rect 8050 21013 8152 21047
rect 8186 21013 8288 21047
rect 8322 21013 8424 21047
rect 8458 21013 8560 21047
rect 8594 21013 8596 21047
rect 7880 20911 8596 21013
rect 7914 20877 8016 20911
rect 8050 20877 8152 20911
rect 8186 20877 8288 20911
rect 8322 20877 8424 20911
rect 8458 20877 8560 20911
rect 8594 20877 8596 20911
rect 7880 20775 8596 20877
rect 7914 20741 8016 20775
rect 8050 20741 8152 20775
rect 8186 20741 8288 20775
rect 8322 20741 8424 20775
rect 8458 20741 8560 20775
rect 8594 20741 8596 20775
rect 7880 20639 8596 20741
rect 7914 20605 8016 20639
rect 8050 20605 8152 20639
rect 8186 20605 8288 20639
rect 8322 20605 8424 20639
rect 8458 20605 8560 20639
rect 8594 20605 8596 20639
rect 7880 20503 8596 20605
rect 7914 20469 8016 20503
rect 8050 20469 8152 20503
rect 8186 20469 8288 20503
rect 8322 20469 8424 20503
rect 8458 20469 8560 20503
rect 8594 20469 8596 20503
rect 7880 20405 8596 20469
rect 9278 20405 9284 29511
rect 7880 20367 9284 20405
rect 7914 20333 8016 20367
rect 8050 20333 8152 20367
rect 8186 20333 8288 20367
rect 8322 20333 8424 20367
rect 8458 20333 8560 20367
rect 8594 20366 8696 20367
rect 8730 20366 8832 20367
rect 8866 20366 8968 20367
rect 9002 20366 9104 20367
rect 9138 20366 9240 20367
rect 9274 20366 9284 20367
rect 8594 20333 8596 20366
rect 7880 20332 8596 20333
rect 8630 20332 8668 20366
rect 8730 20333 8740 20366
rect 8702 20332 8740 20333
rect 8774 20332 8812 20366
rect 8866 20333 8884 20366
rect 8846 20332 8884 20333
rect 8918 20332 8956 20366
rect 9002 20333 9028 20366
rect 8990 20332 9028 20333
rect 9062 20332 9100 20366
rect 9138 20333 9172 20366
rect 9134 20332 9172 20333
rect 9206 20333 9240 20366
rect 9206 20332 9244 20333
rect 9278 20332 9284 20366
rect 7880 20293 9284 20332
rect 7880 20259 8596 20293
rect 8630 20259 8668 20293
rect 8702 20259 8740 20293
rect 8774 20259 8812 20293
rect 8846 20259 8884 20293
rect 8918 20259 8956 20293
rect 8990 20259 9028 20293
rect 9062 20259 9100 20293
rect 9134 20259 9172 20293
rect 9206 20259 9244 20293
rect 9278 20259 9284 20293
rect 7880 20231 9284 20259
rect 7914 20197 8016 20231
rect 8050 20197 8152 20231
rect 8186 20197 8288 20231
rect 8322 20197 8424 20231
rect 8458 20197 8560 20231
rect 8594 20220 8696 20231
rect 8730 20220 8832 20231
rect 8866 20220 8968 20231
rect 9002 20220 9104 20231
rect 9138 20220 9240 20231
rect 9274 20220 9284 20231
rect 8594 20197 8596 20220
rect 7880 20186 8596 20197
rect 8630 20186 8668 20220
rect 8730 20197 8740 20220
rect 8702 20186 8740 20197
rect 8774 20186 8812 20220
rect 8866 20197 8884 20220
rect 8846 20186 8884 20197
rect 8918 20186 8956 20220
rect 9002 20197 9028 20220
rect 8990 20186 9028 20197
rect 9062 20186 9100 20220
rect 9138 20197 9172 20220
rect 9134 20186 9172 20197
rect 9206 20197 9240 20220
rect 9206 20186 9244 20197
rect 9278 20186 9284 20220
rect 7880 20147 9284 20186
rect 7880 20113 8596 20147
rect 8630 20113 8668 20147
rect 8702 20113 8740 20147
rect 8774 20113 8812 20147
rect 8846 20113 8884 20147
rect 8918 20113 8956 20147
rect 8990 20113 9028 20147
rect 9062 20113 9100 20147
rect 9134 20113 9172 20147
rect 9206 20113 9244 20147
rect 9278 20113 9284 20147
rect 7880 20095 9284 20113
rect 7914 20061 8016 20095
rect 8050 20061 8152 20095
rect 8186 20061 8288 20095
rect 8322 20061 8424 20095
rect 8458 20061 8560 20095
rect 8594 20074 8696 20095
rect 8730 20074 8832 20095
rect 8866 20074 8968 20095
rect 9002 20074 9104 20095
rect 9138 20074 9240 20095
rect 9274 20074 9284 20095
rect 8594 20061 8596 20074
rect 7880 20040 8596 20061
rect 8630 20040 8668 20074
rect 8730 20061 8740 20074
rect 8702 20040 8740 20061
rect 8774 20040 8812 20074
rect 8866 20061 8884 20074
rect 8846 20040 8884 20061
rect 8918 20040 8956 20074
rect 9002 20061 9028 20074
rect 8990 20040 9028 20061
rect 9062 20040 9100 20074
rect 9138 20061 9172 20074
rect 9134 20040 9172 20061
rect 9206 20061 9240 20074
rect 9206 20040 9244 20061
rect 9278 20040 9284 20074
rect 7880 20001 9284 20040
rect 7880 19967 8596 20001
rect 8630 19967 8668 20001
rect 8702 19967 8740 20001
rect 8774 19967 8812 20001
rect 8846 19967 8884 20001
rect 8918 19967 8956 20001
rect 8990 19967 9028 20001
rect 9062 19967 9100 20001
rect 9134 19967 9172 20001
rect 9206 19967 9244 20001
rect 9278 19967 9284 20001
rect 7880 19959 9284 19967
rect 7914 19925 8016 19959
rect 8050 19925 8152 19959
rect 8186 19925 8288 19959
rect 8322 19925 8424 19959
rect 8458 19925 8560 19959
rect 8594 19928 8696 19959
rect 8730 19928 8832 19959
rect 8866 19928 8968 19959
rect 9002 19928 9104 19959
rect 9138 19928 9240 19959
rect 9274 19928 9284 19959
rect 8594 19925 8596 19928
rect 7880 19894 8596 19925
rect 8630 19894 8668 19928
rect 8730 19925 8740 19928
rect 8702 19894 8740 19925
rect 8774 19894 8812 19928
rect 8866 19925 8884 19928
rect 8846 19894 8884 19925
rect 8918 19894 8956 19928
rect 9002 19925 9028 19928
rect 8990 19894 9028 19925
rect 9062 19894 9100 19928
rect 9138 19925 9172 19928
rect 9134 19894 9172 19925
rect 9206 19925 9240 19928
rect 9206 19894 9244 19925
rect 9278 19894 9284 19928
rect 7880 19855 9284 19894
rect 7880 19823 8596 19855
rect 7914 19789 8016 19823
rect 8050 19789 8152 19823
rect 8186 19789 8288 19823
rect 8322 19789 8424 19823
rect 8458 19789 8560 19823
rect 8594 19821 8596 19823
rect 8630 19821 8668 19855
rect 8702 19823 8740 19855
rect 8730 19821 8740 19823
rect 8774 19821 8812 19855
rect 8846 19823 8884 19855
rect 8866 19821 8884 19823
rect 8918 19821 8956 19855
rect 8990 19823 9028 19855
rect 9002 19821 9028 19823
rect 9062 19821 9100 19855
rect 9134 19823 9172 19855
rect 9138 19821 9172 19823
rect 9206 19823 9244 19855
rect 9206 19821 9240 19823
rect 9278 19821 9284 19855
rect 8594 19789 8696 19821
rect 8730 19789 8832 19821
rect 8866 19789 8968 19821
rect 9002 19789 9104 19821
rect 9138 19789 9240 19821
rect 9274 19789 9284 19821
rect 7880 19782 9284 19789
rect 7880 19748 8596 19782
rect 8630 19748 8668 19782
rect 8702 19748 8740 19782
rect 8774 19748 8812 19782
rect 8846 19748 8884 19782
rect 8918 19748 8956 19782
rect 8990 19748 9028 19782
rect 9062 19748 9100 19782
rect 9134 19748 9172 19782
rect 9206 19748 9244 19782
rect 9278 19748 9284 19782
rect 7880 19709 9284 19748
rect 7880 19687 8596 19709
rect 7914 19653 8016 19687
rect 8050 19653 8152 19687
rect 8186 19653 8288 19687
rect 8322 19653 8424 19687
rect 8458 19653 8560 19687
rect 8594 19675 8596 19687
rect 8630 19675 8668 19709
rect 8702 19687 8740 19709
rect 8730 19675 8740 19687
rect 8774 19675 8812 19709
rect 8846 19687 8884 19709
rect 8866 19675 8884 19687
rect 8918 19675 8956 19709
rect 8990 19687 9028 19709
rect 9002 19675 9028 19687
rect 9062 19675 9100 19709
rect 9134 19687 9172 19709
rect 9138 19675 9172 19687
rect 9206 19687 9244 19709
rect 9206 19675 9240 19687
rect 9278 19675 9284 19709
rect 8594 19653 8696 19675
rect 8730 19653 8832 19675
rect 8866 19653 8968 19675
rect 9002 19653 9104 19675
rect 9138 19653 9240 19675
rect 9274 19653 9284 19675
rect 7880 19636 9284 19653
rect 7880 19602 8596 19636
rect 8630 19602 8668 19636
rect 8702 19602 8740 19636
rect 8774 19602 8812 19636
rect 8846 19602 8884 19636
rect 8918 19602 8956 19636
rect 8990 19602 9028 19636
rect 9062 19602 9100 19636
rect 9134 19602 9172 19636
rect 9206 19602 9244 19636
rect 9278 19602 9284 19636
rect 7880 19563 9284 19602
rect 7880 19551 8596 19563
rect 7914 19517 8016 19551
rect 8050 19517 8152 19551
rect 8186 19517 8288 19551
rect 8322 19517 8424 19551
rect 8458 19517 8560 19551
rect 8594 19529 8596 19551
rect 8630 19529 8668 19563
rect 8702 19551 8740 19563
rect 8730 19529 8740 19551
rect 8774 19529 8812 19563
rect 8846 19551 8884 19563
rect 8866 19529 8884 19551
rect 8918 19529 8956 19563
rect 8990 19551 9028 19563
rect 9002 19529 9028 19551
rect 9062 19529 9100 19563
rect 9134 19551 9172 19563
rect 9138 19529 9172 19551
rect 9206 19551 9244 19563
rect 9206 19529 9240 19551
rect 9278 19529 9284 19563
rect 8594 19517 8696 19529
rect 8730 19517 8832 19529
rect 8866 19517 8968 19529
rect 9002 19517 9104 19529
rect 9138 19517 9240 19529
rect 9274 19517 9284 19529
rect 7880 19490 9284 19517
rect 7880 19456 8596 19490
rect 8630 19456 8668 19490
rect 8702 19456 8740 19490
rect 8774 19456 8812 19490
rect 8846 19456 8884 19490
rect 8918 19456 8956 19490
rect 8990 19456 9028 19490
rect 9062 19456 9100 19490
rect 9134 19456 9172 19490
rect 9206 19456 9244 19490
rect 9278 19456 9284 19490
rect 7880 19417 9284 19456
rect 7880 19415 8596 19417
rect 7914 19381 8016 19415
rect 8050 19381 8152 19415
rect 8186 19381 8288 19415
rect 8322 19381 8424 19415
rect 8458 19381 8560 19415
rect 8594 19383 8596 19415
rect 8630 19383 8668 19417
rect 8702 19415 8740 19417
rect 8730 19383 8740 19415
rect 8774 19383 8812 19417
rect 8846 19415 8884 19417
rect 8866 19383 8884 19415
rect 8918 19383 8956 19417
rect 8990 19415 9028 19417
rect 9002 19383 9028 19415
rect 9062 19383 9100 19417
rect 9134 19415 9172 19417
rect 9138 19383 9172 19415
rect 9206 19415 9244 19417
rect 9206 19383 9240 19415
rect 9278 19383 9284 19417
rect 8594 19381 8696 19383
rect 8730 19381 8832 19383
rect 8866 19381 8968 19383
rect 9002 19381 9104 19383
rect 9138 19381 9240 19383
rect 9274 19381 9284 19383
rect 7880 19344 9284 19381
rect 7880 19310 8596 19344
rect 8630 19310 8668 19344
rect 8702 19310 8740 19344
rect 8774 19310 8812 19344
rect 8846 19310 8884 19344
rect 8918 19310 8956 19344
rect 8990 19310 9028 19344
rect 9062 19310 9100 19344
rect 9134 19310 9172 19344
rect 9206 19310 9244 19344
rect 9278 19310 9284 19344
rect 7880 19279 9284 19310
rect 7914 19245 8016 19279
rect 8050 19245 8152 19279
rect 8186 19245 8288 19279
rect 8322 19245 8424 19279
rect 8458 19245 8560 19279
rect 8594 19271 8696 19279
rect 8730 19271 8832 19279
rect 8866 19271 8968 19279
rect 9002 19271 9104 19279
rect 9138 19271 9240 19279
rect 9274 19271 9284 19279
rect 8594 19245 8596 19271
rect 7880 19237 8596 19245
rect 8630 19237 8668 19271
rect 8730 19245 8740 19271
rect 8702 19237 8740 19245
rect 8774 19237 8812 19271
rect 8866 19245 8884 19271
rect 8846 19237 8884 19245
rect 8918 19237 8956 19271
rect 9002 19245 9028 19271
rect 8990 19237 9028 19245
rect 9062 19237 9100 19271
rect 9138 19245 9172 19271
rect 9134 19237 9172 19245
rect 9206 19245 9240 19271
rect 9206 19237 9244 19245
rect 9278 19237 9284 19271
rect 7880 19198 9284 19237
rect 7880 19164 8596 19198
rect 8630 19164 8668 19198
rect 8702 19164 8740 19198
rect 8774 19164 8812 19198
rect 8846 19164 8884 19198
rect 8918 19164 8956 19198
rect 8990 19164 9028 19198
rect 9062 19164 9100 19198
rect 9134 19164 9172 19198
rect 9206 19164 9244 19198
rect 9278 19164 9284 19198
rect 7880 19143 9284 19164
rect 7914 19109 8016 19143
rect 8050 19109 8152 19143
rect 8186 19109 8288 19143
rect 8322 19109 8424 19143
rect 8458 19109 8560 19143
rect 8594 19125 8696 19143
rect 8730 19125 8832 19143
rect 8866 19125 8968 19143
rect 9002 19125 9104 19143
rect 9138 19125 9240 19143
rect 9274 19125 9284 19143
rect 8594 19109 8596 19125
rect 7880 19091 8596 19109
rect 8630 19091 8668 19125
rect 8730 19109 8740 19125
rect 8702 19091 8740 19109
rect 8774 19091 8812 19125
rect 8866 19109 8884 19125
rect 8846 19091 8884 19109
rect 8918 19091 8956 19125
rect 9002 19109 9028 19125
rect 8990 19091 9028 19109
rect 9062 19091 9100 19125
rect 9138 19109 9172 19125
rect 9134 19091 9172 19109
rect 9206 19109 9240 19125
rect 9206 19091 9244 19109
rect 9278 19091 9284 19125
rect 7880 19052 9284 19091
rect 7880 19018 8596 19052
rect 8630 19018 8668 19052
rect 8702 19018 8740 19052
rect 8774 19018 8812 19052
rect 8846 19018 8884 19052
rect 8918 19018 8956 19052
rect 8990 19018 9028 19052
rect 9062 19018 9100 19052
rect 9134 19018 9172 19052
rect 9206 19018 9244 19052
rect 9278 19018 9284 19052
rect 7880 19007 9284 19018
rect 7914 18973 8016 19007
rect 8050 18973 8152 19007
rect 8186 18973 8288 19007
rect 8322 18973 8424 19007
rect 8458 18973 8560 19007
rect 8594 18979 8696 19007
rect 8730 18979 8832 19007
rect 8866 18979 8968 19007
rect 9002 18979 9104 19007
rect 9138 18979 9240 19007
rect 9274 18979 9284 19007
rect 8594 18973 8596 18979
rect 7880 18945 8596 18973
rect 8630 18945 8668 18979
rect 8730 18973 8740 18979
rect 8702 18945 8740 18973
rect 8774 18945 8812 18979
rect 8866 18973 8884 18979
rect 8846 18945 8884 18973
rect 8918 18945 8956 18979
rect 9002 18973 9028 18979
rect 8990 18945 9028 18973
rect 9062 18945 9100 18979
rect 9138 18973 9172 18979
rect 9134 18945 9172 18973
rect 9206 18973 9240 18979
rect 9206 18945 9244 18973
rect 9278 18945 9284 18979
rect 7880 18906 9284 18945
rect 7880 18872 8596 18906
rect 8630 18872 8668 18906
rect 8702 18872 8740 18906
rect 8774 18872 8812 18906
rect 8846 18872 8884 18906
rect 8918 18872 8956 18906
rect 8990 18872 9028 18906
rect 9062 18872 9100 18906
rect 9134 18872 9172 18906
rect 9206 18872 9244 18906
rect 9278 18872 9284 18906
rect 7880 18871 9284 18872
rect 7914 18837 8016 18871
rect 8050 18837 8152 18871
rect 8186 18837 8288 18871
rect 8322 18837 8424 18871
rect 8458 18837 8560 18871
rect 8594 18837 8696 18871
rect 8730 18837 8832 18871
rect 8866 18837 8968 18871
rect 9002 18837 9104 18871
rect 9138 18837 9240 18871
rect 9274 18837 9284 18871
rect 7880 18833 9284 18837
rect 7880 18799 8596 18833
rect 8630 18799 8668 18833
rect 8702 18799 8740 18833
rect 8774 18799 8812 18833
rect 8846 18799 8884 18833
rect 8918 18799 8956 18833
rect 8990 18799 9028 18833
rect 9062 18799 9100 18833
rect 9134 18799 9172 18833
rect 9206 18799 9244 18833
rect 9278 18799 9284 18833
rect 7880 18760 9284 18799
rect 7880 18735 8596 18760
rect 7914 18701 8016 18735
rect 8050 18701 8152 18735
rect 8186 18701 8288 18735
rect 8322 18701 8424 18735
rect 8458 18701 8560 18735
rect 8594 18726 8596 18735
rect 8630 18726 8668 18760
rect 8702 18735 8740 18760
rect 8730 18726 8740 18735
rect 8774 18726 8812 18760
rect 8846 18735 8884 18760
rect 8866 18726 8884 18735
rect 8918 18726 8956 18760
rect 8990 18735 9028 18760
rect 9002 18726 9028 18735
rect 9062 18726 9100 18760
rect 9134 18735 9172 18760
rect 9138 18726 9172 18735
rect 9206 18735 9244 18760
rect 9206 18726 9240 18735
rect 9278 18726 9284 18760
rect 8594 18701 8696 18726
rect 8730 18701 8832 18726
rect 8866 18701 8968 18726
rect 9002 18701 9104 18726
rect 9138 18701 9240 18726
rect 9274 18701 9284 18726
rect 7880 18687 9284 18701
rect 7880 18653 8596 18687
rect 8630 18653 8668 18687
rect 8702 18653 8740 18687
rect 8774 18653 8812 18687
rect 8846 18653 8884 18687
rect 8918 18653 8956 18687
rect 8990 18653 9028 18687
rect 9062 18653 9100 18687
rect 9134 18653 9172 18687
rect 9206 18653 9244 18687
rect 9278 18653 9284 18687
rect 7880 18614 9284 18653
rect 7880 18599 8596 18614
rect 7914 18565 8016 18599
rect 8050 18565 8152 18599
rect 8186 18565 8288 18599
rect 8322 18565 8424 18599
rect 8458 18565 8560 18599
rect 8594 18580 8596 18599
rect 8630 18580 8668 18614
rect 8702 18599 8740 18614
rect 8730 18580 8740 18599
rect 8774 18580 8812 18614
rect 8846 18599 8884 18614
rect 8866 18580 8884 18599
rect 8918 18580 8956 18614
rect 8990 18599 9028 18614
rect 9002 18580 9028 18599
rect 9062 18580 9100 18614
rect 9134 18599 9172 18614
rect 9138 18580 9172 18599
rect 9206 18599 9244 18614
rect 9206 18580 9240 18599
rect 9278 18580 9284 18614
rect 8594 18565 8696 18580
rect 8730 18565 8832 18580
rect 8866 18565 8968 18580
rect 9002 18565 9104 18580
rect 9138 18565 9240 18580
rect 9274 18565 9284 18580
rect 7880 18541 9284 18565
rect 7880 18507 8596 18541
rect 8630 18507 8668 18541
rect 8702 18507 8740 18541
rect 8774 18507 8812 18541
rect 8846 18507 8884 18541
rect 8918 18507 8956 18541
rect 8990 18507 9028 18541
rect 9062 18507 9100 18541
rect 9134 18507 9172 18541
rect 9206 18507 9244 18541
rect 9278 18507 9284 18541
rect 7880 18468 9284 18507
rect 7880 18463 8596 18468
rect 7914 18429 8016 18463
rect 8050 18429 8152 18463
rect 8186 18429 8288 18463
rect 8322 18429 8424 18463
rect 8458 18429 8560 18463
rect 8594 18434 8596 18463
rect 8630 18434 8668 18468
rect 8702 18463 8740 18468
rect 8730 18434 8740 18463
rect 8774 18434 8812 18468
rect 8846 18463 8884 18468
rect 8866 18434 8884 18463
rect 8918 18434 8956 18468
rect 8990 18463 9028 18468
rect 9002 18434 9028 18463
rect 9062 18434 9100 18468
rect 9134 18463 9172 18468
rect 9138 18434 9172 18463
rect 9206 18463 9244 18468
rect 9206 18434 9240 18463
rect 9278 18434 9284 18468
rect 8594 18429 8696 18434
rect 8730 18429 8832 18434
rect 8866 18429 8968 18434
rect 9002 18429 9104 18434
rect 9138 18429 9240 18434
rect 9274 18429 9284 18434
rect 7880 18395 9284 18429
rect 7880 18361 8596 18395
rect 8630 18361 8668 18395
rect 8702 18361 8740 18395
rect 8774 18361 8812 18395
rect 8846 18361 8884 18395
rect 8918 18361 8956 18395
rect 8990 18361 9028 18395
rect 9062 18361 9100 18395
rect 9134 18361 9172 18395
rect 9206 18361 9244 18395
rect 9278 18361 9284 18395
rect 7880 18327 9284 18361
rect 7914 18293 8016 18327
rect 8050 18293 8152 18327
rect 8186 18293 8288 18327
rect 8322 18293 8424 18327
rect 8458 18293 8560 18327
rect 8594 18322 8696 18327
rect 8730 18322 8832 18327
rect 8866 18322 8968 18327
rect 9002 18322 9104 18327
rect 9138 18322 9240 18327
rect 9274 18322 9284 18327
rect 8594 18293 8596 18322
rect 7880 18288 8596 18293
rect 8630 18288 8668 18322
rect 8730 18293 8740 18322
rect 8702 18288 8740 18293
rect 8774 18288 8812 18322
rect 8866 18293 8884 18322
rect 8846 18288 8884 18293
rect 8918 18288 8956 18322
rect 9002 18293 9028 18322
rect 8990 18288 9028 18293
rect 9062 18288 9100 18322
rect 9138 18293 9172 18322
rect 9134 18288 9172 18293
rect 9206 18293 9240 18322
rect 9206 18288 9244 18293
rect 9278 18288 9284 18322
rect 7880 18249 9284 18288
rect 7880 18215 8596 18249
rect 8630 18215 8668 18249
rect 8702 18215 8740 18249
rect 8774 18215 8812 18249
rect 8846 18215 8884 18249
rect 8918 18215 8956 18249
rect 8990 18215 9028 18249
rect 9062 18215 9100 18249
rect 9134 18215 9172 18249
rect 9206 18215 9244 18249
rect 9278 18215 9284 18249
rect 7880 18191 9284 18215
rect 7914 18157 8016 18191
rect 8050 18157 8152 18191
rect 8186 18157 8288 18191
rect 8322 18157 8424 18191
rect 8458 18157 8560 18191
rect 8594 18176 8696 18191
rect 8730 18176 8832 18191
rect 8866 18176 8968 18191
rect 9002 18176 9104 18191
rect 9138 18176 9240 18191
rect 9274 18176 9284 18191
rect 8594 18157 8596 18176
rect 7880 18142 8596 18157
rect 8630 18142 8668 18176
rect 8730 18157 8740 18176
rect 8702 18142 8740 18157
rect 8774 18142 8812 18176
rect 8866 18157 8884 18176
rect 8846 18142 8884 18157
rect 8918 18142 8956 18176
rect 9002 18157 9028 18176
rect 8990 18142 9028 18157
rect 9062 18142 9100 18176
rect 9138 18157 9172 18176
rect 9134 18142 9172 18157
rect 9206 18157 9240 18176
rect 9206 18142 9244 18157
rect 9278 18142 9284 18176
rect 7880 18103 9284 18142
rect 7880 18069 8596 18103
rect 8630 18069 8668 18103
rect 8702 18069 8740 18103
rect 8774 18069 8812 18103
rect 8846 18069 8884 18103
rect 8918 18069 8956 18103
rect 8990 18069 9028 18103
rect 9062 18069 9100 18103
rect 9134 18069 9172 18103
rect 9206 18069 9244 18103
rect 9278 18069 9284 18103
rect 7880 18055 9284 18069
rect 7914 18021 8016 18055
rect 8050 18021 8152 18055
rect 8186 18021 8288 18055
rect 8322 18021 8424 18055
rect 8458 18021 8560 18055
rect 8594 18030 8696 18055
rect 8730 18030 8832 18055
rect 8866 18030 8968 18055
rect 9002 18030 9104 18055
rect 9138 18030 9240 18055
rect 9274 18030 9284 18055
rect 8594 18021 8596 18030
rect 7880 17996 8596 18021
rect 8630 17996 8668 18030
rect 8730 18021 8740 18030
rect 8702 17996 8740 18021
rect 8774 17996 8812 18030
rect 8866 18021 8884 18030
rect 8846 17996 8884 18021
rect 8918 17996 8956 18030
rect 9002 18021 9028 18030
rect 8990 17996 9028 18021
rect 9062 17996 9100 18030
rect 9138 18021 9172 18030
rect 9134 17996 9172 18021
rect 9206 18021 9240 18030
rect 9206 17996 9244 18021
rect 9278 17996 9284 18030
rect 7880 17957 9284 17996
rect 7880 17923 8596 17957
rect 8630 17923 8668 17957
rect 8702 17923 8740 17957
rect 8774 17923 8812 17957
rect 8846 17923 8884 17957
rect 8918 17923 8956 17957
rect 8990 17923 9028 17957
rect 9062 17923 9100 17957
rect 9134 17923 9172 17957
rect 9206 17923 9244 17957
rect 9278 17923 9284 17957
rect 7880 17919 9284 17923
rect 7914 17885 8016 17919
rect 8050 17885 8152 17919
rect 8186 17885 8288 17919
rect 8322 17885 8424 17919
rect 8458 17885 8560 17919
rect 8594 17885 8696 17919
rect 8730 17885 8832 17919
rect 8866 17885 8968 17919
rect 9002 17885 9104 17919
rect 9138 17885 9240 17919
rect 9274 17885 9284 17919
rect 7880 17884 9284 17885
rect 7880 17850 8596 17884
rect 8630 17850 8668 17884
rect 8702 17850 8740 17884
rect 8774 17850 8812 17884
rect 8846 17850 8884 17884
rect 8918 17850 8956 17884
rect 8990 17850 9028 17884
rect 9062 17850 9100 17884
rect 9134 17850 9172 17884
rect 9206 17850 9244 17884
rect 9278 17850 9284 17884
rect 7880 17811 9284 17850
rect 7880 17783 8596 17811
rect 7914 17749 8016 17783
rect 8050 17749 8152 17783
rect 8186 17749 8288 17783
rect 8322 17749 8424 17783
rect 8458 17749 8560 17783
rect 8594 17777 8596 17783
rect 8630 17777 8668 17811
rect 8702 17783 8740 17811
rect 8730 17777 8740 17783
rect 8774 17777 8812 17811
rect 8846 17783 8884 17811
rect 8866 17777 8884 17783
rect 8918 17777 8956 17811
rect 8990 17783 9028 17811
rect 9002 17777 9028 17783
rect 9062 17777 9100 17811
rect 9134 17783 9172 17811
rect 9138 17777 9172 17783
rect 9206 17783 9244 17811
rect 9206 17777 9240 17783
rect 9278 17777 9284 17811
rect 8594 17749 8696 17777
rect 8730 17749 8832 17777
rect 8866 17749 8968 17777
rect 9002 17749 9104 17777
rect 9138 17749 9240 17777
rect 9274 17749 9284 17777
rect 7880 17738 9284 17749
rect 7880 17704 8596 17738
rect 8630 17704 8668 17738
rect 8702 17704 8740 17738
rect 8774 17704 8812 17738
rect 8846 17704 8884 17738
rect 8918 17704 8956 17738
rect 8990 17704 9028 17738
rect 9062 17704 9100 17738
rect 9134 17704 9172 17738
rect 9206 17704 9244 17738
rect 9278 17704 9284 17738
rect 7880 17672 9284 17704
rect 7880 17647 9274 17672
rect 7914 17613 8016 17647
rect 8050 17613 8152 17647
rect 8186 17613 8288 17647
rect 8322 17613 8424 17647
rect 8458 17613 8560 17647
rect 8594 17613 8696 17647
rect 8730 17613 8832 17647
rect 8866 17613 8968 17647
rect 9002 17613 9104 17647
rect 9138 17613 9240 17647
rect 7880 17581 9274 17613
rect 1003 17477 1005 17511
rect 1039 17477 1141 17511
rect 1175 17477 1277 17511
rect 1311 17477 1413 17511
rect 1447 17477 1549 17511
rect 1583 17477 1685 17511
rect 1003 17375 1719 17477
rect 1003 17341 1005 17375
rect 1039 17341 1141 17375
rect 1175 17341 1277 17375
rect 1311 17341 1413 17375
rect 1447 17341 1549 17375
rect 1583 17341 1685 17375
rect 1003 17239 1719 17341
rect 1003 17205 1005 17239
rect 1039 17205 1141 17239
rect 1175 17205 1277 17239
rect 1311 17205 1413 17239
rect 1447 17205 1549 17239
rect 1583 17205 1685 17239
rect 1003 17103 1719 17205
rect 1003 17069 1005 17103
rect 1039 17069 1141 17103
rect 1175 17069 1277 17103
rect 1311 17069 1413 17103
rect 1447 17069 1549 17103
rect 1583 17069 1685 17103
rect 1003 16967 1719 17069
rect 1003 16933 1005 16967
rect 1039 16933 1141 16967
rect 1175 16933 1277 16967
rect 1311 16933 1413 16967
rect 1447 16933 1549 16967
rect 1583 16933 1685 16967
rect 1003 16831 1719 16933
rect 1003 16797 1005 16831
rect 1039 16797 1141 16831
rect 1175 16797 1277 16831
rect 1311 16797 1413 16831
rect 1447 16797 1549 16831
rect 1583 16797 1685 16831
rect 1003 16695 1719 16797
rect 1003 16661 1005 16695
rect 1039 16661 1141 16695
rect 1175 16661 1277 16695
rect 1311 16661 1413 16695
rect 1447 16661 1549 16695
rect 1583 16661 1685 16695
rect 1003 16559 1719 16661
rect 1003 16525 1005 16559
rect 1039 16525 1141 16559
rect 1175 16525 1277 16559
rect 1311 16525 1413 16559
rect 1447 16525 1549 16559
rect 1583 16525 1685 16559
rect 1003 16423 1719 16525
rect 7870 17549 9284 17581
rect 1003 16389 1005 16423
rect 1039 16389 1141 16423
rect 1175 16389 1277 16423
rect 1311 16389 1413 16423
rect 1447 16389 1549 16423
rect 1583 16389 1685 16423
rect 1003 16287 1719 16389
rect 1003 16253 1005 16287
rect 1039 16253 1141 16287
rect 1175 16253 1277 16287
rect 1311 16253 1413 16287
rect 1447 16253 1549 16287
rect 1583 16253 1685 16287
rect 1003 16151 1719 16253
rect 1003 16117 1005 16151
rect 1039 16117 1141 16151
rect 1175 16117 1277 16151
rect 1311 16117 1413 16151
rect 1447 16117 1549 16151
rect 1583 16117 1685 16151
rect 1003 16015 1719 16117
rect 1003 15981 1005 16015
rect 1039 15981 1141 16015
rect 1175 15981 1277 16015
rect 1311 15981 1413 16015
rect 1447 15981 1549 16015
rect 1583 15981 1685 16015
rect 1003 15879 1719 15981
rect 1003 15845 1005 15879
rect 1039 15845 1141 15879
rect 1175 15845 1277 15879
rect 1311 15845 1413 15879
rect 1447 15845 1549 15879
rect 1583 15845 1685 15879
rect 1003 15743 1719 15845
rect 1003 15709 1005 15743
rect 1039 15709 1141 15743
rect 1175 15709 1277 15743
rect 1311 15709 1413 15743
rect 1447 15709 1549 15743
rect 1583 15709 1685 15743
rect 1003 15607 1719 15709
rect 1003 15573 1005 15607
rect 1039 15573 1141 15607
rect 1175 15573 1277 15607
rect 1311 15573 1413 15607
rect 1447 15573 1549 15607
rect 1583 15573 1685 15607
rect 1003 15471 1719 15573
rect 1003 15437 1005 15471
rect 1039 15437 1141 15471
rect 1175 15437 1277 15471
rect 1311 15437 1413 15471
rect 1447 15437 1549 15471
rect 1583 15437 1685 15471
rect 1003 15335 1719 15437
rect 1003 15301 1005 15335
rect 1039 15301 1141 15335
rect 1175 15301 1277 15335
rect 1311 15301 1413 15335
rect 1447 15301 1549 15335
rect 1583 15301 1685 15335
rect 1003 15199 1719 15301
rect 1003 15165 1005 15199
rect 1039 15165 1141 15199
rect 1175 15165 1277 15199
rect 1311 15165 1413 15199
rect 1447 15165 1549 15199
rect 1583 15165 1685 15199
rect 1003 15063 1719 15165
rect 1003 15029 1005 15063
rect 1039 15029 1141 15063
rect 1175 15029 1277 15063
rect 1311 15029 1413 15063
rect 1447 15029 1549 15063
rect 1583 15029 1685 15063
rect 1003 14927 1719 15029
rect 1003 14893 1005 14927
rect 1039 14893 1141 14927
rect 1175 14893 1277 14927
rect 1311 14893 1413 14927
rect 1447 14893 1549 14927
rect 1583 14893 1685 14927
rect 1003 14791 1719 14893
rect 1003 14757 1005 14791
rect 1039 14757 1141 14791
rect 1175 14757 1277 14791
rect 1311 14757 1413 14791
rect 1447 14757 1549 14791
rect 1583 14757 1685 14791
rect 1003 14655 1719 14757
rect 1003 14621 1005 14655
rect 1039 14621 1141 14655
rect 1175 14621 1277 14655
rect 1311 14621 1413 14655
rect 1447 14621 1549 14655
rect 1583 14621 1685 14655
rect 1003 14519 1719 14621
rect 1003 14485 1005 14519
rect 1039 14485 1141 14519
rect 1175 14485 1277 14519
rect 1311 14485 1413 14519
rect 1447 14485 1549 14519
rect 1583 14485 1685 14519
rect 1003 14383 1719 14485
rect 1003 14349 1005 14383
rect 1039 14349 1141 14383
rect 1175 14349 1277 14383
rect 1311 14349 1413 14383
rect 1447 14349 1549 14383
rect 1583 14349 1685 14383
rect 1003 14247 1719 14349
rect 1003 14213 1005 14247
rect 1039 14213 1141 14247
rect 1175 14213 1277 14247
rect 1311 14213 1413 14247
rect 1447 14213 1549 14247
rect 1583 14213 1685 14247
rect 1003 14111 1719 14213
rect 1003 14077 1005 14111
rect 1039 14077 1141 14111
rect 1175 14077 1277 14111
rect 1311 14077 1413 14111
rect 1447 14077 1549 14111
rect 1583 14077 1685 14111
rect 1003 13975 1719 14077
rect 1003 13941 1005 13975
rect 1039 13941 1141 13975
rect 1175 13941 1277 13975
rect 1311 13941 1413 13975
rect 1447 13941 1549 13975
rect 1583 13941 1685 13975
rect 1003 13839 1719 13941
rect 1003 13805 1005 13839
rect 1039 13805 1141 13839
rect 1175 13805 1277 13839
rect 1311 13805 1413 13839
rect 1447 13805 1549 13839
rect 1583 13805 1685 13839
rect 1003 13703 1719 13805
rect 1003 13669 1005 13703
rect 1039 13669 1141 13703
rect 1175 13669 1277 13703
rect 1311 13669 1413 13703
rect 1447 13669 1549 13703
rect 1583 13669 1685 13703
rect 1003 13567 1719 13669
rect 1003 13533 1005 13567
rect 1039 13533 1141 13567
rect 1175 13533 1277 13567
rect 1311 13533 1413 13567
rect 1447 13533 1549 13567
rect 1583 13533 1685 13567
rect 1003 13431 1719 13533
rect 1003 13397 1005 13431
rect 1039 13397 1141 13431
rect 1175 13397 1277 13431
rect 1311 13397 1413 13431
rect 1447 13397 1549 13431
rect 1583 13397 1685 13431
rect 1003 13295 1719 13397
rect 1003 13261 1005 13295
rect 1039 13261 1141 13295
rect 1175 13261 1277 13295
rect 1311 13261 1413 13295
rect 1447 13261 1549 13295
rect 1583 13261 1685 13295
rect 1003 13159 1719 13261
rect 1003 13125 1005 13159
rect 1039 13125 1141 13159
rect 1175 13125 1277 13159
rect 1311 13125 1413 13159
rect 1447 13125 1549 13159
rect 1583 13125 1685 13159
rect 1003 13023 1719 13125
rect 1003 12989 1005 13023
rect 1039 12989 1141 13023
rect 1175 12989 1277 13023
rect 1311 12989 1413 13023
rect 1447 12989 1549 13023
rect 1583 12989 1685 13023
rect 1003 12887 1719 12989
rect 1003 12853 1005 12887
rect 1039 12853 1141 12887
rect 1175 12853 1277 12887
rect 1311 12853 1413 12887
rect 1447 12853 1549 12887
rect 1583 12853 1685 12887
rect 1003 12751 1719 12853
rect 1003 12717 1005 12751
rect 1039 12717 1141 12751
rect 1175 12717 1277 12751
rect 1311 12717 1413 12751
rect 1447 12717 1549 12751
rect 1583 12717 1685 12751
rect 1003 12615 1719 12717
rect 1003 12581 1005 12615
rect 1039 12581 1141 12615
rect 1175 12581 1277 12615
rect 1311 12581 1413 12615
rect 1447 12581 1549 12615
rect 1583 12581 1685 12615
rect 1003 12479 1719 12581
rect 1003 12445 1005 12479
rect 1039 12445 1141 12479
rect 1175 12445 1277 12479
rect 1311 12445 1413 12479
rect 1447 12445 1549 12479
rect 1583 12445 1685 12479
rect 1003 12343 1719 12445
rect 1003 12309 1005 12343
rect 1039 12309 1141 12343
rect 1175 12309 1277 12343
rect 1311 12309 1413 12343
rect 1447 12309 1549 12343
rect 1583 12309 1685 12343
rect 1003 12207 1719 12309
rect 1003 12173 1005 12207
rect 1039 12173 1141 12207
rect 1175 12173 1277 12207
rect 1311 12173 1413 12207
rect 1447 12173 1549 12207
rect 1583 12173 1685 12207
rect 1003 12071 1719 12173
rect 1003 12037 1005 12071
rect 1039 12037 1141 12071
rect 1175 12037 1277 12071
rect 1311 12037 1413 12071
rect 1447 12037 1549 12071
rect 1583 12037 1685 12071
rect 1003 11935 1719 12037
rect 1003 11901 1005 11935
rect 1039 11901 1141 11935
rect 1175 11901 1277 11935
rect 1311 11901 1413 11935
rect 1447 11901 1549 11935
rect 1583 11901 1685 11935
rect 1003 11799 1719 11901
rect 1003 11765 1005 11799
rect 1039 11765 1141 11799
rect 1175 11765 1277 11799
rect 1311 11765 1413 11799
rect 1447 11765 1549 11799
rect 1583 11765 1685 11799
rect 1003 11663 1719 11765
rect 1003 11629 1005 11663
rect 1039 11629 1141 11663
rect 1175 11629 1277 11663
rect 1311 11629 1413 11663
rect 1447 11629 1549 11663
rect 1583 11629 1685 11663
rect 1003 11527 1719 11629
rect 1003 11493 1005 11527
rect 1039 11493 1141 11527
rect 1175 11493 1277 11527
rect 1311 11493 1413 11527
rect 1447 11493 1549 11527
rect 1583 11493 1685 11527
rect 1003 11391 1719 11493
rect 1003 11357 1005 11391
rect 1039 11357 1141 11391
rect 1175 11357 1277 11391
rect 1311 11357 1413 11391
rect 1447 11357 1549 11391
rect 1583 11357 1685 11391
rect 1003 11255 1719 11357
rect 1003 11221 1005 11255
rect 1039 11221 1141 11255
rect 1175 11221 1277 11255
rect 1311 11221 1413 11255
rect 1447 11221 1549 11255
rect 1583 11221 1685 11255
rect 1003 11119 1719 11221
rect 1003 11085 1005 11119
rect 1039 11085 1141 11119
rect 1175 11085 1277 11119
rect 1311 11085 1413 11119
rect 1447 11085 1549 11119
rect 1583 11085 1685 11119
rect 1003 10983 1719 11085
rect 1003 10949 1005 10983
rect 1039 10949 1141 10983
rect 1175 10949 1277 10983
rect 1311 10949 1413 10983
rect 1447 10949 1549 10983
rect 1583 10949 1685 10983
rect 1003 10847 1719 10949
rect 1003 10813 1005 10847
rect 1039 10813 1141 10847
rect 1175 10813 1277 10847
rect 1311 10813 1413 10847
rect 1447 10813 1549 10847
rect 1583 10813 1685 10847
rect 1003 10711 1719 10813
rect 1003 10677 1005 10711
rect 1039 10677 1141 10711
rect 1175 10677 1277 10711
rect 1311 10677 1413 10711
rect 1447 10677 1549 10711
rect 1583 10677 1685 10711
rect 1003 10575 1719 10677
rect 1003 10541 1005 10575
rect 1039 10541 1141 10575
rect 1175 10541 1277 10575
rect 1311 10541 1413 10575
rect 1447 10541 1549 10575
rect 1583 10541 1685 10575
rect 1003 10439 1719 10541
rect 1003 10405 1005 10439
rect 1039 10405 1141 10439
rect 1175 10405 1277 10439
rect 1311 10405 1413 10439
rect 1447 10405 1549 10439
rect 1583 10405 1685 10439
rect 1003 10303 1719 10405
rect 1003 10269 1005 10303
rect 1039 10269 1141 10303
rect 1175 10269 1277 10303
rect 1311 10269 1413 10303
rect 1447 10269 1549 10303
rect 1583 10269 1685 10303
rect 1003 10167 1719 10269
rect 1003 10133 1005 10167
rect 1039 10133 1141 10167
rect 1175 10133 1277 10167
rect 1311 10133 1413 10167
rect 1447 10133 1549 10167
rect 1583 10133 1685 10167
rect 1003 10031 1719 10133
rect 1003 9997 1005 10031
rect 1039 9997 1141 10031
rect 1175 9997 1277 10031
rect 1311 9997 1413 10031
rect 1447 9997 1549 10031
rect 1583 9997 1685 10031
rect 1003 9895 1719 9997
rect 1003 9861 1005 9895
rect 1039 9861 1141 9895
rect 1175 9861 1277 9895
rect 1311 9861 1413 9895
rect 1447 9861 1549 9895
rect 1583 9861 1685 9895
rect 1003 9759 1719 9861
rect 1003 9725 1005 9759
rect 1039 9725 1141 9759
rect 1175 9725 1277 9759
rect 1311 9725 1413 9759
rect 1447 9725 1549 9759
rect 1583 9725 1685 9759
rect 1003 9623 1719 9725
rect 1003 9589 1005 9623
rect 1039 9589 1141 9623
rect 1175 9589 1277 9623
rect 1311 9589 1413 9623
rect 1447 9589 1549 9623
rect 1583 9589 1685 9623
rect 1003 9487 1719 9589
rect 1003 9453 1005 9487
rect 1039 9453 1141 9487
rect 1175 9453 1277 9487
rect 1311 9453 1413 9487
rect 1447 9453 1549 9487
rect 1583 9453 1685 9487
rect 1003 9351 1719 9453
rect 1003 9317 1005 9351
rect 1039 9317 1141 9351
rect 1175 9317 1277 9351
rect 1311 9317 1413 9351
rect 1447 9317 1549 9351
rect 1583 9317 1685 9351
rect 1003 9215 1719 9317
rect 1003 9181 1005 9215
rect 1039 9181 1141 9215
rect 1175 9181 1277 9215
rect 1311 9181 1413 9215
rect 1447 9181 1549 9215
rect 1583 9181 1685 9215
rect 1003 9079 1719 9181
rect 1003 9045 1005 9079
rect 1039 9045 1141 9079
rect 1175 9045 1277 9079
rect 1311 9045 1413 9079
rect 1447 9045 1549 9079
rect 1583 9045 1685 9079
rect 1003 8943 1719 9045
rect 1003 8909 1005 8943
rect 1039 8909 1141 8943
rect 1175 8909 1277 8943
rect 1311 8909 1413 8943
rect 1447 8909 1549 8943
rect 1583 8909 1685 8943
rect 1003 8807 1719 8909
rect 1003 8773 1005 8807
rect 1039 8773 1141 8807
rect 1175 8773 1277 8807
rect 1311 8773 1413 8807
rect 1447 8773 1549 8807
rect 1583 8773 1685 8807
rect 1003 8671 1719 8773
rect 1003 8637 1005 8671
rect 1039 8637 1141 8671
rect 1175 8637 1277 8671
rect 1311 8637 1413 8671
rect 1447 8637 1549 8671
rect 1583 8637 1685 8671
rect 1003 8535 1719 8637
rect 1003 8501 1005 8535
rect 1039 8501 1141 8535
rect 1175 8501 1277 8535
rect 1311 8501 1413 8535
rect 1447 8501 1549 8535
rect 1583 8501 1685 8535
rect 1003 8399 1719 8501
rect 1003 8365 1005 8399
rect 1039 8365 1141 8399
rect 1175 8365 1277 8399
rect 1311 8365 1413 8399
rect 1447 8365 1549 8399
rect 1583 8365 1685 8399
rect 1003 8263 1719 8365
rect 1003 8229 1005 8263
rect 1039 8229 1141 8263
rect 1175 8229 1277 8263
rect 1311 8229 1413 8263
rect 1447 8229 1549 8263
rect 1583 8229 1685 8263
rect 1003 8127 1719 8229
rect 1003 8093 1005 8127
rect 1039 8093 1141 8127
rect 1175 8093 1277 8127
rect 1311 8093 1413 8127
rect 1447 8093 1549 8127
rect 1583 8093 1685 8127
rect 1003 7991 1719 8093
rect 1003 7957 1005 7991
rect 1039 7957 1141 7991
rect 1175 7957 1277 7991
rect 1311 7957 1413 7991
rect 1447 7957 1549 7991
rect 1583 7957 1685 7991
rect 1003 7855 1719 7957
rect 1003 7821 1005 7855
rect 1039 7821 1141 7855
rect 1175 7821 1277 7855
rect 1311 7821 1413 7855
rect 1447 7821 1549 7855
rect 1583 7821 1685 7855
rect 1003 7719 1719 7821
rect 1003 7685 1005 7719
rect 1039 7685 1141 7719
rect 1175 7685 1277 7719
rect 1311 7685 1413 7719
rect 1447 7685 1549 7719
rect 1583 7685 1685 7719
rect 1003 7583 1719 7685
rect 1003 7549 1005 7583
rect 1039 7549 1141 7583
rect 1175 7549 1277 7583
rect 1311 7549 1413 7583
rect 1447 7549 1549 7583
rect 1583 7549 1685 7583
rect 1003 7447 1719 7549
rect 1003 7413 1005 7447
rect 1039 7413 1141 7447
rect 1175 7413 1277 7447
rect 1311 7413 1413 7447
rect 1447 7413 1549 7447
rect 1583 7413 1685 7447
rect 1003 7311 1719 7413
rect 1003 7277 1005 7311
rect 1039 7277 1141 7311
rect 1175 7277 1277 7311
rect 1311 7277 1413 7311
rect 1447 7277 1549 7311
rect 1583 7277 1685 7311
rect 1003 7175 1719 7277
rect 1003 7141 1005 7175
rect 1039 7141 1141 7175
rect 1175 7141 1277 7175
rect 1311 7141 1413 7175
rect 1447 7141 1549 7175
rect 1583 7141 1685 7175
rect 1003 7039 1719 7141
rect 1003 7005 1005 7039
rect 1039 7005 1141 7039
rect 1175 7005 1277 7039
rect 1311 7005 1413 7039
rect 1447 7005 1549 7039
rect 1583 7005 1685 7039
rect 1003 6903 1719 7005
rect 1003 6869 1005 6903
rect 1039 6869 1141 6903
rect 1175 6869 1277 6903
rect 1311 6869 1413 6903
rect 1447 6869 1549 6903
rect 1583 6869 1685 6903
rect 1003 6767 1719 6869
rect 1003 6733 1005 6767
rect 1039 6733 1141 6767
rect 1175 6733 1277 6767
rect 1311 6733 1413 6767
rect 1447 6733 1549 6767
rect 1583 6733 1685 6767
rect 1003 6631 1719 6733
rect 1003 6597 1005 6631
rect 1039 6597 1141 6631
rect 1175 6597 1277 6631
rect 1311 6597 1413 6631
rect 1447 6597 1549 6631
rect 1583 6597 1685 6631
rect 1003 6495 1719 6597
rect 1003 6461 1005 6495
rect 1039 6461 1141 6495
rect 1175 6461 1277 6495
rect 1311 6461 1413 6495
rect 1447 6461 1549 6495
rect 1583 6461 1685 6495
rect 1003 6359 1719 6461
rect 1003 6325 1005 6359
rect 1039 6325 1141 6359
rect 1175 6325 1277 6359
rect 1311 6325 1413 6359
rect 1447 6325 1549 6359
rect 1583 6325 1685 6359
rect 1003 6223 1719 6325
rect 1003 6189 1005 6223
rect 1039 6189 1141 6223
rect 1175 6189 1277 6223
rect 1311 6189 1413 6223
rect 1447 6189 1549 6223
rect 1583 6189 1685 6223
rect 1003 6087 1719 6189
rect 1003 6053 1005 6087
rect 1039 6053 1141 6087
rect 1175 6053 1277 6087
rect 1311 6053 1413 6087
rect 1447 6053 1549 6087
rect 1583 6053 1685 6087
rect 1003 5951 1719 6053
rect 1003 5917 1005 5951
rect 1039 5917 1141 5951
rect 1175 5917 1277 5951
rect 1311 5917 1413 5951
rect 1447 5917 1549 5951
rect 1583 5917 1685 5951
rect 1003 5815 1719 5917
rect 1003 5781 1005 5815
rect 1039 5781 1141 5815
rect 1175 5781 1277 5815
rect 1311 5781 1413 5815
rect 1447 5781 1549 5815
rect 1583 5781 1685 5815
rect 1003 5679 1719 5781
rect 1003 5645 1005 5679
rect 1039 5645 1141 5679
rect 1175 5645 1277 5679
rect 1311 5645 1413 5679
rect 1447 5645 1549 5679
rect 1583 5645 1685 5679
rect 1003 5543 1719 5645
rect 1003 5509 1005 5543
rect 1039 5509 1141 5543
rect 1175 5509 1277 5543
rect 1311 5509 1413 5543
rect 1447 5509 1549 5543
rect 1583 5509 1685 5543
rect 1003 5407 1719 5509
rect 1003 5373 1005 5407
rect 1039 5373 1141 5407
rect 1175 5373 1277 5407
rect 1311 5373 1413 5407
rect 1447 5373 1549 5407
rect 1583 5373 1685 5407
rect 1003 5271 1719 5373
rect 1003 5237 1005 5271
rect 1039 5237 1141 5271
rect 1175 5237 1277 5271
rect 1311 5237 1413 5271
rect 1447 5237 1549 5271
rect 1583 5237 1685 5271
rect 1003 5135 1719 5237
rect 1003 5101 1005 5135
rect 1039 5101 1141 5135
rect 1175 5101 1277 5135
rect 1311 5101 1413 5135
rect 1447 5101 1549 5135
rect 1583 5101 1685 5135
rect 1003 4999 1719 5101
rect 1003 4965 1005 4999
rect 1039 4965 1141 4999
rect 1175 4965 1277 4999
rect 1311 4965 1413 4999
rect 1447 4965 1549 4999
rect 1583 4965 1685 4999
rect 1003 4863 1719 4965
rect 1003 4829 1005 4863
rect 1039 4829 1141 4863
rect 1175 4829 1277 4863
rect 1311 4829 1413 4863
rect 1447 4829 1549 4863
rect 1583 4829 1685 4863
rect 1003 4727 1719 4829
rect 1003 4693 1005 4727
rect 1039 4693 1141 4727
rect 1175 4693 1277 4727
rect 1311 4693 1413 4727
rect 1447 4693 1549 4727
rect 1583 4693 1685 4727
rect 1003 4591 1719 4693
rect 1003 4557 1005 4591
rect 1039 4557 1141 4591
rect 1175 4557 1277 4591
rect 1311 4557 1413 4591
rect 1447 4557 1549 4591
rect 1583 4557 1685 4591
rect 1003 4455 1719 4557
rect 1003 4421 1005 4455
rect 1039 4421 1141 4455
rect 1175 4421 1277 4455
rect 1311 4421 1413 4455
rect 1447 4421 1549 4455
rect 1583 4421 1685 4455
rect 1003 4319 1719 4421
rect 1003 4285 1005 4319
rect 1039 4285 1141 4319
rect 1175 4285 1277 4319
rect 1311 4285 1413 4319
rect 1447 4285 1549 4319
rect 1583 4285 1685 4319
rect 1003 4183 1719 4285
rect 1003 4149 1005 4183
rect 1039 4149 1141 4183
rect 1175 4149 1277 4183
rect 1311 4149 1413 4183
rect 1447 4149 1549 4183
rect 1583 4149 1685 4183
rect 1003 4047 1719 4149
rect 1003 4013 1005 4047
rect 1039 4013 1141 4047
rect 1175 4013 1277 4047
rect 1311 4013 1413 4047
rect 1447 4013 1549 4047
rect 1583 4013 1685 4047
rect 1003 3911 1719 4013
rect 1003 3877 1005 3911
rect 1039 3877 1141 3911
rect 1175 3877 1277 3911
rect 1311 3877 1413 3911
rect 1447 3877 1549 3911
rect 1583 3877 1685 3911
rect 1003 3775 1719 3877
rect 1003 3741 1005 3775
rect 1039 3741 1141 3775
rect 1175 3741 1277 3775
rect 1311 3741 1413 3775
rect 1447 3741 1549 3775
rect 1583 3741 1685 3775
rect 1003 3639 1719 3741
rect 1003 3605 1005 3639
rect 1039 3605 1141 3639
rect 1175 3605 1277 3639
rect 1311 3605 1413 3639
rect 1447 3605 1549 3639
rect 1583 3605 1685 3639
rect 1003 3503 1719 3605
rect 1003 3469 1005 3503
rect 1039 3469 1141 3503
rect 1175 3469 1277 3503
rect 1311 3469 1413 3503
rect 1447 3469 1549 3503
rect 1583 3469 1685 3503
rect 1003 3367 1719 3469
rect 1003 3333 1005 3367
rect 1039 3333 1141 3367
rect 1175 3333 1277 3367
rect 1311 3333 1413 3367
rect 1447 3333 1549 3367
rect 1583 3333 1685 3367
rect 1003 3231 1719 3333
rect 1003 3197 1005 3231
rect 1039 3197 1141 3231
rect 1175 3197 1277 3231
rect 1311 3197 1413 3231
rect 1447 3197 1549 3231
rect 1583 3197 1685 3231
rect 1003 3125 1719 3197
rect 315 3095 1719 3125
rect 315 3086 325 3095
rect 359 3086 461 3095
rect 495 3086 597 3095
rect 631 3086 733 3095
rect 767 3086 869 3095
rect 903 3086 1005 3095
rect 315 3052 321 3086
rect 359 3061 393 3086
rect 355 3052 393 3061
rect 427 3061 461 3086
rect 427 3052 465 3061
rect 499 3052 537 3086
rect 571 3061 597 3086
rect 571 3052 609 3061
rect 643 3052 681 3086
rect 715 3061 733 3086
rect 715 3052 753 3061
rect 787 3052 825 3086
rect 859 3061 869 3086
rect 859 3052 897 3061
rect 931 3052 969 3086
rect 1003 3061 1005 3086
rect 1039 3061 1141 3095
rect 1175 3061 1277 3095
rect 1311 3061 1413 3095
rect 1447 3061 1549 3095
rect 1583 3061 1685 3095
rect 1003 3052 1719 3061
rect 315 3013 1719 3052
rect 315 2979 321 3013
rect 355 2979 393 3013
rect 427 2979 465 3013
rect 499 2979 537 3013
rect 571 2979 609 3013
rect 643 2979 681 3013
rect 715 2979 753 3013
rect 787 2979 825 3013
rect 859 2979 897 3013
rect 931 2979 969 3013
rect 1003 2979 1719 3013
rect 315 2959 1719 2979
rect 315 2940 325 2959
rect 359 2940 461 2959
rect 495 2940 597 2959
rect 631 2940 733 2959
rect 767 2940 869 2959
rect 903 2940 1005 2959
rect 315 2906 321 2940
rect 359 2925 393 2940
rect 355 2906 393 2925
rect 427 2925 461 2940
rect 427 2906 465 2925
rect 499 2906 537 2940
rect 571 2925 597 2940
rect 571 2906 609 2925
rect 643 2906 681 2940
rect 715 2925 733 2940
rect 715 2906 753 2925
rect 787 2906 825 2940
rect 859 2925 869 2940
rect 859 2906 897 2925
rect 931 2906 969 2940
rect 1003 2925 1005 2940
rect 1039 2925 1141 2959
rect 1175 2925 1277 2959
rect 1311 2925 1413 2959
rect 1447 2925 1549 2959
rect 1583 2925 1685 2959
rect 1003 2906 1719 2925
rect 315 2867 1719 2906
rect 315 2833 321 2867
rect 355 2833 393 2867
rect 427 2833 465 2867
rect 499 2833 537 2867
rect 571 2833 609 2867
rect 643 2833 681 2867
rect 715 2833 753 2867
rect 787 2833 825 2867
rect 859 2833 897 2867
rect 931 2833 969 2867
rect 1003 2833 1719 2867
rect 315 2823 1719 2833
rect 315 2794 325 2823
rect 359 2794 461 2823
rect 495 2794 597 2823
rect 631 2794 733 2823
rect 767 2794 869 2823
rect 903 2794 1005 2823
rect 315 2760 321 2794
rect 359 2789 393 2794
rect 355 2760 393 2789
rect 427 2789 461 2794
rect 427 2760 465 2789
rect 499 2760 537 2794
rect 571 2789 597 2794
rect 571 2760 609 2789
rect 643 2760 681 2794
rect 715 2789 733 2794
rect 715 2760 753 2789
rect 787 2760 825 2794
rect 859 2789 869 2794
rect 859 2760 897 2789
rect 931 2760 969 2794
rect 1003 2789 1005 2794
rect 1039 2789 1141 2823
rect 1175 2789 1277 2823
rect 1311 2789 1413 2823
rect 1447 2789 1549 2823
rect 1583 2789 1685 2823
rect 1003 2760 1719 2789
rect 315 2721 1719 2760
rect 315 2687 321 2721
rect 355 2687 393 2721
rect 427 2687 465 2721
rect 499 2687 537 2721
rect 571 2687 609 2721
rect 643 2687 681 2721
rect 715 2687 753 2721
rect 787 2687 825 2721
rect 859 2687 897 2721
rect 931 2687 969 2721
rect 1003 2687 1719 2721
rect 315 2653 325 2687
rect 359 2653 461 2687
rect 495 2653 597 2687
rect 631 2653 733 2687
rect 767 2653 869 2687
rect 903 2653 1005 2687
rect 1039 2653 1141 2687
rect 1175 2653 1277 2687
rect 1311 2653 1413 2687
rect 1447 2653 1549 2687
rect 1583 2653 1685 2687
rect 315 2648 1719 2653
rect 315 2614 321 2648
rect 355 2614 393 2648
rect 427 2614 465 2648
rect 499 2614 537 2648
rect 571 2614 609 2648
rect 643 2614 681 2648
rect 715 2614 753 2648
rect 787 2614 825 2648
rect 859 2614 897 2648
rect 931 2614 969 2648
rect 1003 2614 1719 2648
rect 315 2575 1719 2614
rect 315 2541 321 2575
rect 355 2551 393 2575
rect 359 2541 393 2551
rect 427 2551 465 2575
rect 427 2541 461 2551
rect 499 2541 537 2575
rect 571 2551 609 2575
rect 571 2541 597 2551
rect 643 2541 681 2575
rect 715 2551 753 2575
rect 715 2541 733 2551
rect 787 2541 825 2575
rect 859 2551 897 2575
rect 859 2541 869 2551
rect 931 2541 969 2575
rect 1003 2551 1719 2575
rect 1003 2541 1005 2551
rect 315 2517 325 2541
rect 359 2517 461 2541
rect 495 2517 597 2541
rect 631 2517 733 2541
rect 767 2517 869 2541
rect 903 2517 1005 2541
rect 1039 2517 1141 2551
rect 1175 2517 1277 2551
rect 1311 2517 1413 2551
rect 1447 2517 1549 2551
rect 1583 2517 1685 2551
rect 315 2502 1719 2517
rect 315 2468 321 2502
rect 355 2468 393 2502
rect 427 2468 465 2502
rect 499 2468 537 2502
rect 571 2468 609 2502
rect 643 2468 681 2502
rect 715 2468 753 2502
rect 787 2468 825 2502
rect 859 2468 897 2502
rect 931 2468 969 2502
rect 1003 2468 1719 2502
rect 315 2429 1719 2468
rect 315 2395 321 2429
rect 355 2414 393 2429
rect 359 2395 393 2414
rect 427 2414 465 2429
rect 427 2395 461 2414
rect 499 2395 537 2429
rect 571 2414 609 2429
rect 571 2395 597 2414
rect 643 2395 681 2429
rect 715 2414 753 2429
rect 715 2395 733 2414
rect 787 2395 825 2429
rect 859 2414 897 2429
rect 859 2395 869 2414
rect 931 2395 969 2429
rect 1003 2414 1719 2429
rect 1003 2395 1005 2414
rect 315 2380 325 2395
rect 359 2380 461 2395
rect 495 2380 597 2395
rect 631 2380 733 2395
rect 767 2380 869 2395
rect 903 2380 1005 2395
rect 1039 2380 1141 2414
rect 1175 2380 1277 2414
rect 1311 2380 1413 2414
rect 1447 2380 1549 2414
rect 1583 2380 1685 2414
rect 315 2356 1719 2380
rect 315 2322 321 2356
rect 355 2322 393 2356
rect 427 2322 465 2356
rect 499 2322 537 2356
rect 571 2322 609 2356
rect 643 2322 681 2356
rect 715 2322 753 2356
rect 787 2322 825 2356
rect 859 2322 897 2356
rect 931 2322 969 2356
rect 1003 2322 1719 2356
rect 315 2283 1719 2322
rect 315 2249 321 2283
rect 355 2277 393 2283
rect 359 2249 393 2277
rect 427 2277 465 2283
rect 427 2249 461 2277
rect 499 2249 537 2283
rect 571 2277 609 2283
rect 571 2249 597 2277
rect 643 2249 681 2283
rect 715 2277 753 2283
rect 715 2249 733 2277
rect 787 2249 825 2283
rect 859 2277 897 2283
rect 859 2249 869 2277
rect 931 2249 969 2283
rect 1003 2277 1719 2283
rect 1003 2249 1005 2277
rect 315 2243 325 2249
rect 359 2243 461 2249
rect 495 2243 597 2249
rect 631 2243 733 2249
rect 767 2243 869 2249
rect 903 2243 1005 2249
rect 1039 2243 1141 2277
rect 1175 2243 1277 2277
rect 1311 2243 1413 2277
rect 1447 2243 1549 2277
rect 1583 2243 1685 2277
rect 315 2210 1719 2243
rect 315 2176 321 2210
rect 355 2176 393 2210
rect 427 2176 465 2210
rect 499 2176 537 2210
rect 571 2176 609 2210
rect 643 2176 681 2210
rect 715 2176 753 2210
rect 787 2176 825 2210
rect 859 2176 897 2210
rect 931 2176 969 2210
rect 1003 2176 1719 2210
rect 315 2140 1719 2176
rect 315 2137 325 2140
rect 359 2137 461 2140
rect 495 2137 597 2140
rect 631 2137 733 2140
rect 767 2137 869 2140
rect 903 2137 1005 2140
rect 315 2103 321 2137
rect 359 2106 393 2137
rect 355 2103 393 2106
rect 427 2106 461 2137
rect 427 2103 465 2106
rect 499 2103 537 2137
rect 571 2106 597 2137
rect 571 2103 609 2106
rect 643 2103 681 2137
rect 715 2106 733 2137
rect 715 2103 753 2106
rect 787 2103 825 2137
rect 859 2106 869 2137
rect 859 2103 897 2106
rect 931 2103 969 2137
rect 1003 2106 1005 2137
rect 1039 2106 1141 2140
rect 1175 2106 1277 2140
rect 1311 2106 1413 2140
rect 1447 2106 1549 2140
rect 1583 2106 1685 2140
rect 1003 2103 1719 2106
rect 315 2064 1719 2103
rect 315 2030 321 2064
rect 355 2030 393 2064
rect 427 2030 465 2064
rect 499 2030 537 2064
rect 571 2030 609 2064
rect 643 2030 681 2064
rect 715 2030 753 2064
rect 787 2030 825 2064
rect 859 2030 897 2064
rect 931 2030 969 2064
rect 1003 2030 1719 2064
rect 315 2003 1719 2030
rect 315 1991 325 2003
rect 359 1991 461 2003
rect 495 1991 597 2003
rect 631 1991 733 2003
rect 767 1991 869 2003
rect 903 1991 1005 2003
rect 315 1957 321 1991
rect 359 1969 393 1991
rect 355 1957 393 1969
rect 427 1969 461 1991
rect 427 1957 465 1969
rect 499 1957 537 1991
rect 571 1969 597 1991
rect 571 1957 609 1969
rect 643 1957 681 1991
rect 715 1969 733 1991
rect 715 1957 753 1969
rect 787 1957 825 1991
rect 859 1969 869 1991
rect 859 1957 897 1969
rect 931 1957 969 1991
rect 1003 1969 1005 1991
rect 1039 1969 1141 2003
rect 1175 1969 1277 2003
rect 1311 1969 1413 2003
rect 1447 1969 1549 2003
rect 1583 1969 1685 2003
rect 1003 1957 1719 1969
rect 315 1918 1719 1957
rect 315 1884 321 1918
rect 355 1884 393 1918
rect 427 1884 465 1918
rect 499 1884 537 1918
rect 571 1884 609 1918
rect 643 1884 681 1918
rect 715 1884 753 1918
rect 787 1884 825 1918
rect 859 1884 897 1918
rect 931 1884 969 1918
rect 1003 1884 1719 1918
rect 315 1866 1719 1884
rect 315 1845 325 1866
rect 359 1845 461 1866
rect 495 1845 597 1866
rect 631 1845 733 1866
rect 767 1845 869 1866
rect 903 1845 1005 1866
rect 315 1811 321 1845
rect 359 1832 393 1845
rect 355 1811 393 1832
rect 427 1832 461 1845
rect 427 1811 465 1832
rect 499 1811 537 1845
rect 571 1832 597 1845
rect 571 1811 609 1832
rect 643 1811 681 1845
rect 715 1832 733 1845
rect 715 1811 753 1832
rect 787 1811 825 1845
rect 859 1832 869 1845
rect 859 1811 897 1832
rect 931 1811 969 1845
rect 1003 1832 1005 1845
rect 1039 1832 1141 1866
rect 1175 1832 1277 1866
rect 1311 1832 1413 1866
rect 1447 1832 1549 1866
rect 1583 1832 1685 1866
rect 1003 1811 1719 1832
rect 315 1772 1719 1811
rect 315 1738 321 1772
rect 355 1738 393 1772
rect 427 1738 465 1772
rect 499 1738 537 1772
rect 571 1738 609 1772
rect 643 1738 681 1772
rect 715 1738 753 1772
rect 787 1738 825 1772
rect 859 1738 897 1772
rect 931 1738 969 1772
rect 1003 1738 1719 1772
rect 315 1729 1719 1738
rect 315 1699 325 1729
rect 359 1699 461 1729
rect 495 1699 597 1729
rect 631 1699 733 1729
rect 767 1699 869 1729
rect 903 1699 1005 1729
rect 315 1665 321 1699
rect 359 1695 393 1699
rect 355 1665 393 1695
rect 427 1695 461 1699
rect 427 1665 465 1695
rect 499 1665 537 1699
rect 571 1695 597 1699
rect 571 1665 609 1695
rect 643 1665 681 1699
rect 715 1695 733 1699
rect 715 1665 753 1695
rect 787 1665 825 1699
rect 859 1695 869 1699
rect 859 1665 897 1695
rect 931 1665 969 1699
rect 1003 1695 1005 1699
rect 1039 1695 1141 1729
rect 1175 1695 1277 1729
rect 1311 1695 1413 1729
rect 1447 1695 1549 1729
rect 1583 1695 1685 1729
rect 4998 16472 7559 16478
rect 4998 16438 5080 16472
rect 5114 16438 5139 16472
rect 5190 16438 5207 16472
rect 5266 16438 5275 16472
rect 5342 16438 5343 16472
rect 5377 16438 5385 16472
rect 5445 16438 5462 16472
rect 5513 16438 5547 16472
rect 5606 16438 5615 16472
rect 5678 16438 5683 16472
rect 5750 16438 5751 16472
rect 5785 16438 5788 16472
rect 5853 16438 5860 16472
rect 5921 16438 5932 16472
rect 5989 16438 6004 16472
rect 6057 16438 6076 16472
rect 6125 16438 6148 16472
rect 6193 16438 6220 16472
rect 6261 16438 6292 16472
rect 6329 16438 6363 16472
rect 6398 16438 6431 16472
rect 6470 16438 6499 16472
rect 6542 16438 6567 16472
rect 6614 16438 6635 16472
rect 6686 16438 6703 16472
rect 6758 16438 6771 16472
rect 6830 16438 6839 16472
rect 6902 16438 6907 16472
rect 6974 16438 6975 16472
rect 7009 16438 7012 16472
rect 7077 16438 7084 16472
rect 7145 16438 7156 16472
rect 7213 16438 7228 16472
rect 7281 16438 7301 16472
rect 7349 16438 7374 16472
rect 7417 16438 7447 16472
rect 7485 16438 7559 16472
rect 4998 16432 7559 16438
rect 4998 16404 5044 16432
rect 4998 16366 5004 16404
rect 5038 16366 5044 16404
rect 4998 16336 5044 16366
rect 4998 16293 5004 16336
rect 5038 16293 5044 16336
rect 4998 16268 5044 16293
rect 4998 16220 5004 16268
rect 5038 16220 5044 16268
rect 4998 16200 5044 16220
rect 4998 16147 5004 16200
rect 5038 16147 5044 16200
rect 4998 16132 5044 16147
rect 4998 16074 5004 16132
rect 5038 16074 5044 16132
rect 4998 16064 5044 16074
rect 4998 16001 5004 16064
rect 5038 16001 5044 16064
rect 4998 15996 5044 16001
rect 4998 15894 5004 15996
rect 5038 15894 5044 15996
rect 4998 15889 5044 15894
rect 4998 15826 5004 15889
rect 5038 15826 5044 15889
rect 4998 15816 5044 15826
rect 4998 15758 5004 15816
rect 5038 15758 5044 15816
rect 4998 15743 5044 15758
rect 4998 15690 5004 15743
rect 5038 15690 5044 15743
rect 4998 15670 5044 15690
rect 4998 15622 5004 15670
rect 5038 15622 5044 15670
rect 4998 15597 5044 15622
rect 4998 15554 5004 15597
rect 5038 15554 5044 15597
rect 4998 15524 5044 15554
rect 4998 15486 5004 15524
rect 5038 15486 5044 15524
rect 4998 15452 5044 15486
rect 4998 15417 5004 15452
rect 5038 15417 5044 15452
rect 4998 15384 5044 15417
rect 4998 15344 5004 15384
rect 5038 15344 5044 15384
rect 4998 15316 5044 15344
rect 4998 15271 5004 15316
rect 5038 15271 5044 15316
rect 4998 15248 5044 15271
rect 4998 15198 5004 15248
rect 5038 15198 5044 15248
rect 4998 15180 5044 15198
rect 4998 15125 5004 15180
rect 5038 15125 5044 15180
rect 4998 15112 5044 15125
rect 4998 15052 5004 15112
rect 5038 15052 5044 15112
rect 4998 15044 5044 15052
rect 4998 14979 5004 15044
rect 5038 14979 5044 15044
rect 4998 14976 5044 14979
rect 4998 14942 5004 14976
rect 5038 14942 5044 14976
rect 4998 14940 5044 14942
rect 4998 14874 5004 14940
rect 5038 14874 5044 14940
rect 4998 14867 5044 14874
rect 4998 14806 5004 14867
rect 5038 14806 5044 14867
rect 4998 14795 5044 14806
rect 4998 14738 5004 14795
rect 5038 14738 5044 14795
rect 4998 14723 5044 14738
rect 4998 14670 5004 14723
rect 5038 14670 5044 14723
rect 4998 14651 5044 14670
rect 4998 14602 5004 14651
rect 5038 14602 5044 14651
rect 4998 14579 5044 14602
rect 4998 14534 5004 14579
rect 5038 14534 5044 14579
rect 4998 14507 5044 14534
rect 4998 14466 5004 14507
rect 5038 14466 5044 14507
rect 4998 14435 5044 14466
rect 4998 14398 5004 14435
rect 5038 14398 5044 14435
rect 4998 14364 5044 14398
rect 4998 14329 5004 14364
rect 5038 14329 5044 14364
rect 4998 14296 5044 14329
rect 4998 14257 5004 14296
rect 5038 14257 5044 14296
rect 4998 14228 5044 14257
rect 4998 14185 5004 14228
rect 5038 14185 5044 14228
rect 4998 14160 5044 14185
rect 4998 14113 5004 14160
rect 5038 14113 5044 14160
rect 4998 14092 5044 14113
rect 4998 14041 5004 14092
rect 5038 14041 5044 14092
rect 4998 14024 5044 14041
rect 4998 13969 5004 14024
rect 5038 13969 5044 14024
rect 4998 13956 5044 13969
rect 4998 13897 5004 13956
rect 5038 13897 5044 13956
rect 4998 13888 5044 13897
rect 4998 13825 5004 13888
rect 5038 13825 5044 13888
rect 4998 13820 5044 13825
rect 4998 13753 5004 13820
rect 5038 13753 5044 13820
rect 4998 13752 5044 13753
rect 4998 13718 5004 13752
rect 5038 13718 5044 13752
rect 4998 13715 5044 13718
rect 4998 13650 5004 13715
rect 5038 13650 5044 13715
rect 4998 13643 5044 13650
rect 4998 13582 5004 13643
rect 5038 13582 5044 13643
rect 4998 13571 5044 13582
rect 4998 13514 5004 13571
rect 5038 13514 5044 13571
rect 4998 13499 5044 13514
rect 4998 13446 5004 13499
rect 5038 13446 5044 13499
rect 4998 13427 5044 13446
rect 4998 13378 5004 13427
rect 5038 13378 5044 13427
rect 4998 13355 5044 13378
rect 4998 13310 5004 13355
rect 5038 13310 5044 13355
rect 4998 13283 5044 13310
rect 4998 13242 5004 13283
rect 5038 13242 5044 13283
rect 4998 13211 5044 13242
rect 4998 13174 5004 13211
rect 5038 13174 5044 13211
rect 4998 13140 5044 13174
rect 4998 13105 5004 13140
rect 5038 13105 5044 13140
rect 4998 13072 5044 13105
rect 4998 13033 5004 13072
rect 5038 13033 5044 13072
rect 4998 13004 5044 13033
rect 4998 12961 5004 13004
rect 5038 12961 5044 13004
rect 4998 12936 5044 12961
rect 4998 12889 5004 12936
rect 5038 12889 5044 12936
rect 4998 12868 5044 12889
rect 4998 12817 5004 12868
rect 5038 12817 5044 12868
rect 4998 12800 5044 12817
rect 4998 12745 5004 12800
rect 5038 12745 5044 12800
rect 4998 12732 5044 12745
rect 4998 12673 5004 12732
rect 5038 12673 5044 12732
rect 4998 12664 5044 12673
rect 4998 12601 5004 12664
rect 5038 12601 5044 12664
rect 4998 12596 5044 12601
rect 4998 12529 5004 12596
rect 5038 12529 5044 12596
rect 4998 12528 5044 12529
rect 4998 12494 5004 12528
rect 5038 12494 5044 12528
rect 4998 12491 5044 12494
rect 4998 12426 5004 12491
rect 5038 12426 5044 12491
rect 4998 12419 5044 12426
rect 4998 12358 5004 12419
rect 5038 12358 5044 12419
rect 4998 12347 5044 12358
rect 4998 12290 5004 12347
rect 5038 12290 5044 12347
rect 4998 12275 5044 12290
rect 4998 12222 5004 12275
rect 5038 12222 5044 12275
rect 4998 12203 5044 12222
rect 4998 12154 5004 12203
rect 5038 12154 5044 12203
rect 4998 12131 5044 12154
rect 4998 12086 5004 12131
rect 5038 12086 5044 12131
rect 4998 12059 5044 12086
rect 4998 12018 5004 12059
rect 5038 12018 5044 12059
rect 4998 11987 5044 12018
rect 4998 11950 5004 11987
rect 5038 11950 5044 11987
rect 4998 11916 5044 11950
rect 4998 11881 5004 11916
rect 5038 11881 5044 11916
rect 4998 11848 5044 11881
rect 4998 11809 5004 11848
rect 5038 11809 5044 11848
rect 4998 11780 5044 11809
rect 4998 11737 5004 11780
rect 5038 11737 5044 11780
rect 4998 11712 5044 11737
rect 4998 11665 5004 11712
rect 5038 11665 5044 11712
rect 4998 11644 5044 11665
rect 4998 11593 5004 11644
rect 5038 11593 5044 11644
rect 4998 11576 5044 11593
rect 4998 11521 5004 11576
rect 5038 11521 5044 11576
rect 4998 11508 5044 11521
rect 4998 11449 5004 11508
rect 5038 11449 5044 11508
rect 4998 11440 5044 11449
rect 4998 11377 5004 11440
rect 5038 11377 5044 11440
rect 4998 11372 5044 11377
rect 4998 11305 5004 11372
rect 5038 11305 5044 11372
rect 4998 11304 5044 11305
rect 4998 11270 5004 11304
rect 5038 11270 5044 11304
rect 4998 11267 5044 11270
rect 4998 11202 5004 11267
rect 5038 11202 5044 11267
rect 4998 11195 5044 11202
rect 4998 11134 5004 11195
rect 5038 11134 5044 11195
rect 4998 11123 5044 11134
rect 4998 11066 5004 11123
rect 5038 11066 5044 11123
rect 4998 11051 5044 11066
rect 4998 10998 5004 11051
rect 5038 10998 5044 11051
rect 4998 10979 5044 10998
rect 4998 10930 5004 10979
rect 5038 10930 5044 10979
rect 4998 10907 5044 10930
rect 4998 10862 5004 10907
rect 5038 10862 5044 10907
rect 4998 10835 5044 10862
rect 4998 10794 5004 10835
rect 5038 10794 5044 10835
rect 4998 10763 5044 10794
rect 4998 10726 5004 10763
rect 5038 10726 5044 10763
rect 4998 10692 5044 10726
rect 4998 10657 5004 10692
rect 5038 10657 5044 10692
rect 4998 10624 5044 10657
rect 4998 10585 5004 10624
rect 5038 10585 5044 10624
rect 4998 10556 5044 10585
rect 4998 10513 5004 10556
rect 5038 10513 5044 10556
rect 4998 10488 5044 10513
rect 4998 10441 5004 10488
rect 5038 10441 5044 10488
rect 4998 10420 5044 10441
rect 4998 10369 5004 10420
rect 5038 10369 5044 10420
rect 4998 10352 5044 10369
rect 4998 10297 5004 10352
rect 5038 10297 5044 10352
rect 4998 10284 5044 10297
rect 4998 10225 5004 10284
rect 5038 10225 5044 10284
rect 4998 10216 5044 10225
rect 4998 10153 5004 10216
rect 5038 10153 5044 10216
rect 4998 10148 5044 10153
rect 4998 10081 5004 10148
rect 5038 10081 5044 10148
rect 4998 10080 5044 10081
rect 4998 10046 5004 10080
rect 5038 10046 5044 10080
rect 4998 10043 5044 10046
rect 4998 9978 5004 10043
rect 5038 9978 5044 10043
rect 4998 9971 5044 9978
rect 4998 9910 5004 9971
rect 5038 9910 5044 9971
rect 4998 9899 5044 9910
rect 4998 9842 5004 9899
rect 5038 9842 5044 9899
rect 4998 9827 5044 9842
rect 4998 9774 5004 9827
rect 5038 9774 5044 9827
rect 4998 9755 5044 9774
rect 4998 9706 5004 9755
rect 5038 9706 5044 9755
rect 4998 9683 5044 9706
rect 4998 9638 5004 9683
rect 5038 9638 5044 9683
rect 4998 9611 5044 9638
rect 4998 9570 5004 9611
rect 5038 9570 5044 9611
rect 4998 9539 5044 9570
rect 4998 9502 5004 9539
rect 5038 9502 5044 9539
rect 4998 9468 5044 9502
rect 4998 9433 5004 9468
rect 5038 9433 5044 9468
rect 4998 9400 5044 9433
rect 4998 9361 5004 9400
rect 5038 9361 5044 9400
rect 4998 9332 5044 9361
rect 4998 9289 5004 9332
rect 5038 9289 5044 9332
rect 4998 9264 5044 9289
rect 4998 9217 5004 9264
rect 5038 9217 5044 9264
rect 4998 9196 5044 9217
rect 4998 9145 5004 9196
rect 5038 9145 5044 9196
rect 4998 9128 5044 9145
rect 4998 9073 5004 9128
rect 5038 9073 5044 9128
rect 4998 9060 5044 9073
rect 4998 9001 5004 9060
rect 5038 9001 5044 9060
rect 4998 8992 5044 9001
rect 4998 8929 5004 8992
rect 5038 8929 5044 8992
rect 4998 8924 5044 8929
rect 4998 8857 5004 8924
rect 5038 8857 5044 8924
rect 4998 8856 5044 8857
rect 4998 8822 5004 8856
rect 5038 8822 5044 8856
rect 4998 8819 5044 8822
rect 4998 8754 5004 8819
rect 5038 8754 5044 8819
rect 4998 8747 5044 8754
rect 4998 8686 5004 8747
rect 5038 8686 5044 8747
rect 4998 8675 5044 8686
rect 4998 8618 5004 8675
rect 5038 8618 5044 8675
rect 4998 8603 5044 8618
rect 4998 8550 5004 8603
rect 5038 8550 5044 8603
rect 4998 8531 5044 8550
rect 4998 8482 5004 8531
rect 5038 8482 5044 8531
rect 4998 8459 5044 8482
rect 4998 8414 5004 8459
rect 5038 8414 5044 8459
rect 4998 8387 5044 8414
rect 4998 8346 5004 8387
rect 5038 8346 5044 8387
rect 4998 8315 5044 8346
rect 4998 8278 5004 8315
rect 5038 8278 5044 8315
rect 4998 8244 5044 8278
rect 4998 8209 5004 8244
rect 5038 8209 5044 8244
rect 4998 8176 5044 8209
rect 4998 8137 5004 8176
rect 5038 8137 5044 8176
rect 4998 8108 5044 8137
rect 4998 8065 5004 8108
rect 5038 8065 5044 8108
rect 4998 8040 5044 8065
rect 4998 7993 5004 8040
rect 5038 7993 5044 8040
rect 4998 7972 5044 7993
rect 4998 7921 5004 7972
rect 5038 7921 5044 7972
rect 4998 7904 5044 7921
rect 4998 7849 5004 7904
rect 5038 7849 5044 7904
rect 4998 7836 5044 7849
rect 4998 7777 5004 7836
rect 5038 7777 5044 7836
rect 4998 7768 5044 7777
rect 4998 7705 5004 7768
rect 5038 7705 5044 7768
rect 4998 7700 5044 7705
rect 4998 7633 5004 7700
rect 5038 7633 5044 7700
rect 4998 7632 5044 7633
rect 4998 7598 5004 7632
rect 5038 7598 5044 7632
rect 4998 7595 5044 7598
rect 4998 7530 5004 7595
rect 5038 7530 5044 7595
rect 4998 7523 5044 7530
rect 4998 7462 5004 7523
rect 5038 7462 5044 7523
rect 4998 7451 5044 7462
rect 4998 7394 5004 7451
rect 5038 7394 5044 7451
rect 4998 7379 5044 7394
rect 4998 7326 5004 7379
rect 5038 7326 5044 7379
rect 4998 7307 5044 7326
rect 4998 7258 5004 7307
rect 5038 7258 5044 7307
rect 4998 7235 5044 7258
rect 4998 7190 5004 7235
rect 5038 7190 5044 7235
rect 4998 7163 5044 7190
rect 4998 7122 5004 7163
rect 5038 7122 5044 7163
rect 4998 7091 5044 7122
rect 4998 7054 5004 7091
rect 5038 7054 5044 7091
rect 4998 7020 5044 7054
rect 4998 6985 5004 7020
rect 5038 6985 5044 7020
rect 4998 6952 5044 6985
rect 4998 6913 5004 6952
rect 5038 6913 5044 6952
rect 4998 6884 5044 6913
rect 4998 6841 5004 6884
rect 5038 6841 5044 6884
rect 4998 6816 5044 6841
rect 4998 6769 5004 6816
rect 5038 6769 5044 6816
rect 4998 6748 5044 6769
rect 4998 6697 5004 6748
rect 5038 6697 5044 6748
rect 4998 6680 5044 6697
rect 4998 6625 5004 6680
rect 5038 6625 5044 6680
rect 4998 6612 5044 6625
rect 4998 6553 5004 6612
rect 5038 6553 5044 6612
rect 4998 6544 5044 6553
rect 4998 6481 5004 6544
rect 5038 6481 5044 6544
rect 4998 6476 5044 6481
rect 4998 6409 5004 6476
rect 5038 6409 5044 6476
rect 4998 6408 5044 6409
rect 4998 6374 5004 6408
rect 5038 6374 5044 6408
rect 4998 6371 5044 6374
rect 4998 6306 5004 6371
rect 5038 6306 5044 6371
rect 4998 6299 5044 6306
rect 4998 6238 5004 6299
rect 5038 6238 5044 6299
rect 4998 6227 5044 6238
rect 4998 6170 5004 6227
rect 5038 6170 5044 6227
rect 4998 6155 5044 6170
rect 4998 6102 5004 6155
rect 5038 6102 5044 6155
rect 4998 6083 5044 6102
rect 4998 6034 5004 6083
rect 5038 6034 5044 6083
rect 4998 6011 5044 6034
rect 4998 5966 5004 6011
rect 5038 5966 5044 6011
rect 4998 5939 5044 5966
rect 4998 5898 5004 5939
rect 5038 5898 5044 5939
rect 4998 5867 5044 5898
rect 4998 5830 5004 5867
rect 5038 5830 5044 5867
rect 4998 5796 5044 5830
rect 4998 5761 5004 5796
rect 5038 5761 5044 5796
rect 4998 5728 5044 5761
rect 4998 5689 5004 5728
rect 5038 5689 5044 5728
rect 4998 5660 5044 5689
rect 4998 5617 5004 5660
rect 5038 5617 5044 5660
rect 4998 5592 5044 5617
rect 4998 5545 5004 5592
rect 5038 5545 5044 5592
rect 4998 5524 5044 5545
rect 4998 5473 5004 5524
rect 5038 5473 5044 5524
rect 4998 5456 5044 5473
rect 4998 5401 5004 5456
rect 5038 5401 5044 5456
rect 4998 5388 5044 5401
rect 4998 5329 5004 5388
rect 5038 5329 5044 5388
rect 4998 5320 5044 5329
rect 4998 5257 5004 5320
rect 5038 5257 5044 5320
rect 4998 5252 5044 5257
rect 4998 5185 5004 5252
rect 5038 5185 5044 5252
rect 4998 5184 5044 5185
rect 4998 5150 5004 5184
rect 5038 5150 5044 5184
rect 4998 5147 5044 5150
rect 4998 5082 5004 5147
rect 5038 5082 5044 5147
rect 4998 5075 5044 5082
rect 4998 5014 5004 5075
rect 5038 5014 5044 5075
rect 4998 5003 5044 5014
rect 4998 4946 5004 5003
rect 5038 4946 5044 5003
rect 4998 4931 5044 4946
rect 4998 4878 5004 4931
rect 5038 4878 5044 4931
rect 4998 4859 5044 4878
rect 4998 4810 5004 4859
rect 5038 4810 5044 4859
rect 4998 4787 5044 4810
rect 4998 4742 5004 4787
rect 5038 4742 5044 4787
rect 4998 4715 5044 4742
rect 4998 4674 5004 4715
rect 5038 4674 5044 4715
rect 4998 4643 5044 4674
rect 4998 4606 5004 4643
rect 5038 4606 5044 4643
rect 4998 4572 5044 4606
rect 4998 4537 5004 4572
rect 5038 4537 5044 4572
rect 4998 4504 5044 4537
rect 4998 4465 5004 4504
rect 5038 4465 5044 4504
rect 4998 4436 5044 4465
rect 4998 4393 5004 4436
rect 5038 4393 5044 4436
rect 4998 4368 5044 4393
rect 4998 4321 5004 4368
rect 5038 4321 5044 4368
rect 4998 4300 5044 4321
rect 4998 4249 5004 4300
rect 5038 4249 5044 4300
rect 4998 4232 5044 4249
rect 4998 4177 5004 4232
rect 5038 4177 5044 4232
rect 4998 4164 5044 4177
rect 4998 4105 5004 4164
rect 5038 4105 5044 4164
rect 4998 4096 5044 4105
rect 4998 4033 5004 4096
rect 5038 4033 5044 4096
rect 4998 4028 5044 4033
rect 4998 3961 5004 4028
rect 5038 3961 5044 4028
rect 4998 3960 5044 3961
rect 4998 3926 5004 3960
rect 5038 3926 5044 3960
rect 4998 3923 5044 3926
rect 4998 3858 5004 3923
rect 5038 3858 5044 3923
rect 4998 3851 5044 3858
rect 4998 3790 5004 3851
rect 5038 3790 5044 3851
rect 4998 3779 5044 3790
rect 4998 3722 5004 3779
rect 5038 3722 5044 3779
rect 4998 3707 5044 3722
rect 4998 3654 5004 3707
rect 5038 3654 5044 3707
rect 4998 3635 5044 3654
rect 4998 3586 5004 3635
rect 5038 3586 5044 3635
rect 4998 3563 5044 3586
rect 4998 3518 5004 3563
rect 5038 3518 5044 3563
rect 4998 3491 5044 3518
rect 4998 3450 5004 3491
rect 5038 3450 5044 3491
rect 4998 3419 5044 3450
rect 4998 3382 5004 3419
rect 5038 3382 5044 3419
rect 4998 3348 5044 3382
rect 4998 3313 5004 3348
rect 5038 3313 5044 3348
rect 4998 3280 5044 3313
rect 4998 3241 5004 3280
rect 5038 3241 5044 3280
rect 4998 3212 5044 3241
rect 4998 3169 5004 3212
rect 5038 3169 5044 3212
rect 4998 3144 5044 3169
rect 4998 3097 5004 3144
rect 5038 3097 5044 3144
rect 4998 3076 5044 3097
rect 4998 3025 5004 3076
rect 5038 3025 5044 3076
rect 4998 3008 5044 3025
rect 4998 2953 5004 3008
rect 5038 2953 5044 3008
rect 4998 2940 5044 2953
rect 4998 2881 5004 2940
rect 5038 2881 5044 2940
rect 4998 2872 5044 2881
rect 4998 2809 5004 2872
rect 5038 2809 5044 2872
rect 4998 2804 5044 2809
rect 4998 2737 5004 2804
rect 5038 2737 5044 2804
rect 4998 2736 5044 2737
rect 4998 2702 5004 2736
rect 5038 2702 5044 2736
rect 4998 2699 5044 2702
rect 4998 2634 5004 2699
rect 5038 2634 5044 2699
rect 4998 2627 5044 2634
rect 4998 2566 5004 2627
rect 5038 2566 5044 2627
rect 4998 2555 5044 2566
rect 4998 2498 5004 2555
rect 5038 2498 5044 2555
rect 4998 2483 5044 2498
rect 4998 2430 5004 2483
rect 5038 2430 5044 2483
rect 4998 2411 5044 2430
rect 4998 2362 5004 2411
rect 5038 2362 5044 2411
rect 4998 2339 5044 2362
rect 4998 2294 5004 2339
rect 5038 2294 5044 2339
rect 4998 2267 5044 2294
rect 4998 2226 5004 2267
rect 5038 2226 5044 2267
rect 4998 2195 5044 2226
rect 4998 2158 5004 2195
rect 5038 2158 5044 2195
rect 4998 2124 5044 2158
rect 4998 2089 5004 2124
rect 5038 2089 5044 2124
rect 4998 2056 5044 2089
rect 4998 2017 5004 2056
rect 5038 2017 5044 2056
rect 4998 1988 5044 2017
rect 4998 1945 5004 1988
rect 5038 1945 5044 1988
rect 4998 1907 5044 1945
rect 4998 1873 5004 1907
rect 5038 1873 5044 1907
rect 4998 1855 5044 1873
rect 4998 1801 5004 1855
rect 5038 1801 5044 1855
rect 4998 1769 5044 1801
rect 7513 16400 7559 16432
rect 7513 16349 7519 16400
rect 7553 16349 7559 16400
rect 7513 16328 7559 16349
rect 7513 16281 7519 16328
rect 7553 16281 7559 16328
rect 7513 16256 7559 16281
rect 7513 16213 7519 16256
rect 7553 16213 7559 16256
rect 7513 16184 7559 16213
rect 7513 16145 7519 16184
rect 7553 16145 7559 16184
rect 7513 16112 7559 16145
rect 7513 16077 7519 16112
rect 7553 16077 7559 16112
rect 7513 16043 7559 16077
rect 7513 16006 7519 16043
rect 7553 16006 7559 16043
rect 7513 15975 7559 16006
rect 7513 15934 7519 15975
rect 7553 15934 7559 15975
rect 7513 15907 7559 15934
rect 7513 15862 7519 15907
rect 7553 15862 7559 15907
rect 7513 15839 7559 15862
rect 7513 15790 7519 15839
rect 7553 15790 7559 15839
rect 7513 15771 7559 15790
rect 7513 15718 7519 15771
rect 7553 15718 7559 15771
rect 7513 15703 7559 15718
rect 7513 15646 7519 15703
rect 7553 15646 7559 15703
rect 7513 15635 7559 15646
rect 7513 15574 7519 15635
rect 7553 15574 7559 15635
rect 7513 15567 7559 15574
rect 7513 15502 7519 15567
rect 7553 15502 7559 15567
rect 7513 15499 7559 15502
rect 7513 15465 7519 15499
rect 7553 15465 7559 15499
rect 7513 15464 7559 15465
rect 7513 15397 7519 15464
rect 7553 15397 7559 15464
rect 7513 15392 7559 15397
rect 7513 15329 7519 15392
rect 7553 15329 7559 15392
rect 7513 15320 7559 15329
rect 7513 15261 7519 15320
rect 7553 15261 7559 15320
rect 7513 15248 7559 15261
rect 7513 15193 7519 15248
rect 7553 15193 7559 15248
rect 7513 15176 7559 15193
rect 7513 15125 7519 15176
rect 7553 15125 7559 15176
rect 7513 15104 7559 15125
rect 7513 15057 7519 15104
rect 7553 15057 7559 15104
rect 7513 15032 7559 15057
rect 7513 14989 7519 15032
rect 7553 14989 7559 15032
rect 7513 14960 7559 14989
rect 7513 14921 7519 14960
rect 7553 14921 7559 14960
rect 7513 14888 7559 14921
rect 7513 14853 7519 14888
rect 7553 14853 7559 14888
rect 7513 14819 7559 14853
rect 7513 14782 7519 14819
rect 7553 14782 7559 14819
rect 7513 14751 7559 14782
rect 7513 14710 7519 14751
rect 7553 14710 7559 14751
rect 7513 14683 7559 14710
rect 7513 14638 7519 14683
rect 7553 14638 7559 14683
rect 7513 14615 7559 14638
rect 7513 14566 7519 14615
rect 7553 14566 7559 14615
rect 7513 14547 7559 14566
rect 7513 14494 7519 14547
rect 7553 14494 7559 14547
rect 7513 14479 7559 14494
rect 7513 14422 7519 14479
rect 7553 14422 7559 14479
rect 7513 14411 7559 14422
rect 7513 14350 7519 14411
rect 7553 14350 7559 14411
rect 7513 14343 7559 14350
rect 7513 14278 7519 14343
rect 7553 14278 7559 14343
rect 7513 14275 7559 14278
rect 7513 14241 7519 14275
rect 7553 14241 7559 14275
rect 7513 14240 7559 14241
rect 7513 14173 7519 14240
rect 7553 14173 7559 14240
rect 7513 14168 7559 14173
rect 7513 14105 7519 14168
rect 7553 14105 7559 14168
rect 7513 14096 7559 14105
rect 7513 14037 7519 14096
rect 7553 14037 7559 14096
rect 7513 14024 7559 14037
rect 7513 13969 7519 14024
rect 7553 13969 7559 14024
rect 7513 13952 7559 13969
rect 7513 13901 7519 13952
rect 7553 13901 7559 13952
rect 7513 13880 7559 13901
rect 7513 13833 7519 13880
rect 7553 13833 7559 13880
rect 7513 13808 7559 13833
rect 7513 13765 7519 13808
rect 7553 13765 7559 13808
rect 7513 13736 7559 13765
rect 7513 13697 7519 13736
rect 7553 13697 7559 13736
rect 7513 13664 7559 13697
rect 7513 13629 7519 13664
rect 7553 13629 7559 13664
rect 7513 13595 7559 13629
rect 7513 13558 7519 13595
rect 7553 13558 7559 13595
rect 7513 13527 7559 13558
rect 7513 13486 7519 13527
rect 7553 13486 7559 13527
rect 7513 13459 7559 13486
rect 7513 13414 7519 13459
rect 7553 13414 7559 13459
rect 7513 13391 7559 13414
rect 7513 13342 7519 13391
rect 7553 13342 7559 13391
rect 7513 13323 7559 13342
rect 7513 13270 7519 13323
rect 7553 13270 7559 13323
rect 7513 13255 7559 13270
rect 7513 13198 7519 13255
rect 7553 13198 7559 13255
rect 7513 13187 7559 13198
rect 7513 13126 7519 13187
rect 7553 13126 7559 13187
rect 7513 13119 7559 13126
rect 7513 13054 7519 13119
rect 7553 13054 7559 13119
rect 7513 13051 7559 13054
rect 7513 13017 7519 13051
rect 7553 13017 7559 13051
rect 7513 13016 7559 13017
rect 7513 12949 7519 13016
rect 7553 12949 7559 13016
rect 7513 12944 7559 12949
rect 7513 12881 7519 12944
rect 7553 12881 7559 12944
rect 7513 12872 7559 12881
rect 7513 12813 7519 12872
rect 7553 12813 7559 12872
rect 7513 12800 7559 12813
rect 7513 12745 7519 12800
rect 7553 12745 7559 12800
rect 7513 12728 7559 12745
rect 7513 12677 7519 12728
rect 7553 12677 7559 12728
rect 7513 12656 7559 12677
rect 7513 12609 7519 12656
rect 7553 12609 7559 12656
rect 7513 12584 7559 12609
rect 7513 12541 7519 12584
rect 7553 12541 7559 12584
rect 7513 12512 7559 12541
rect 7513 12473 7519 12512
rect 7553 12473 7559 12512
rect 7513 12440 7559 12473
rect 7513 12405 7519 12440
rect 7553 12405 7559 12440
rect 7513 12371 7559 12405
rect 7513 12334 7519 12371
rect 7553 12334 7559 12371
rect 7513 12303 7559 12334
rect 7513 12262 7519 12303
rect 7553 12262 7559 12303
rect 7513 12235 7559 12262
rect 7513 12190 7519 12235
rect 7553 12190 7559 12235
rect 7513 12167 7559 12190
rect 7513 12118 7519 12167
rect 7553 12118 7559 12167
rect 7513 12099 7559 12118
rect 7513 12046 7519 12099
rect 7553 12046 7559 12099
rect 7513 12031 7559 12046
rect 7513 11974 7519 12031
rect 7553 11974 7559 12031
rect 7513 11963 7559 11974
rect 7513 11902 7519 11963
rect 7553 11902 7559 11963
rect 7513 11895 7559 11902
rect 7513 11830 7519 11895
rect 7553 11830 7559 11895
rect 7513 11827 7559 11830
rect 7513 11793 7519 11827
rect 7553 11793 7559 11827
rect 7513 11792 7559 11793
rect 7513 11725 7519 11792
rect 7553 11725 7559 11792
rect 7513 11720 7559 11725
rect 7513 11657 7519 11720
rect 7553 11657 7559 11720
rect 7513 11648 7559 11657
rect 7513 11589 7519 11648
rect 7553 11589 7559 11648
rect 7513 11576 7559 11589
rect 7513 11521 7519 11576
rect 7553 11521 7559 11576
rect 7513 11504 7559 11521
rect 7513 11453 7519 11504
rect 7553 11453 7559 11504
rect 7513 11432 7559 11453
rect 7513 11385 7519 11432
rect 7553 11385 7559 11432
rect 7513 11360 7559 11385
rect 7513 11317 7519 11360
rect 7553 11317 7559 11360
rect 7513 11288 7559 11317
rect 7513 11249 7519 11288
rect 7553 11249 7559 11288
rect 7513 11216 7559 11249
rect 7513 11181 7519 11216
rect 7553 11181 7559 11216
rect 7513 11147 7559 11181
rect 7513 11110 7519 11147
rect 7553 11110 7559 11147
rect 7513 11079 7559 11110
rect 7513 11038 7519 11079
rect 7553 11038 7559 11079
rect 7513 11011 7559 11038
rect 7513 10966 7519 11011
rect 7553 10966 7559 11011
rect 7513 10943 7559 10966
rect 7513 10894 7519 10943
rect 7553 10894 7559 10943
rect 7513 10875 7559 10894
rect 7513 10822 7519 10875
rect 7553 10822 7559 10875
rect 7513 10807 7559 10822
rect 7513 10750 7519 10807
rect 7553 10750 7559 10807
rect 7513 10739 7559 10750
rect 7513 10678 7519 10739
rect 7553 10678 7559 10739
rect 7513 10671 7559 10678
rect 7513 10606 7519 10671
rect 7553 10606 7559 10671
rect 7513 10603 7559 10606
rect 7513 10569 7519 10603
rect 7553 10569 7559 10603
rect 7513 10568 7559 10569
rect 7513 10501 7519 10568
rect 7553 10501 7559 10568
rect 7513 10496 7559 10501
rect 7513 10433 7519 10496
rect 7553 10433 7559 10496
rect 7513 10424 7559 10433
rect 7513 10365 7519 10424
rect 7553 10365 7559 10424
rect 7513 10352 7559 10365
rect 7513 10297 7519 10352
rect 7553 10297 7559 10352
rect 7513 10280 7559 10297
rect 7513 10229 7519 10280
rect 7553 10229 7559 10280
rect 7513 10208 7559 10229
rect 7513 10161 7519 10208
rect 7553 10161 7559 10208
rect 7513 10136 7559 10161
rect 7513 10093 7519 10136
rect 7553 10093 7559 10136
rect 7513 10064 7559 10093
rect 7513 10025 7519 10064
rect 7553 10025 7559 10064
rect 7513 9992 7559 10025
rect 7513 9957 7519 9992
rect 7553 9957 7559 9992
rect 7513 9923 7559 9957
rect 7513 9886 7519 9923
rect 7553 9886 7559 9923
rect 7513 9855 7559 9886
rect 7513 9814 7519 9855
rect 7553 9814 7559 9855
rect 7513 9787 7559 9814
rect 7513 9742 7519 9787
rect 7553 9742 7559 9787
rect 7513 9719 7559 9742
rect 7513 9670 7519 9719
rect 7553 9670 7559 9719
rect 7513 9651 7559 9670
rect 7513 9598 7519 9651
rect 7553 9598 7559 9651
rect 7513 9583 7559 9598
rect 7513 9526 7519 9583
rect 7553 9526 7559 9583
rect 7513 9515 7559 9526
rect 7513 9454 7519 9515
rect 7553 9454 7559 9515
rect 7513 9447 7559 9454
rect 7513 9382 7519 9447
rect 7553 9382 7559 9447
rect 7513 9379 7559 9382
rect 7513 9345 7519 9379
rect 7553 9345 7559 9379
rect 7513 9344 7559 9345
rect 7513 9277 7519 9344
rect 7553 9277 7559 9344
rect 7513 9272 7559 9277
rect 7513 9209 7519 9272
rect 7553 9209 7559 9272
rect 7513 9200 7559 9209
rect 7513 9141 7519 9200
rect 7553 9141 7559 9200
rect 7513 9128 7559 9141
rect 7513 9073 7519 9128
rect 7553 9073 7559 9128
rect 7513 9056 7559 9073
rect 7513 9005 7519 9056
rect 7553 9005 7559 9056
rect 7513 8984 7559 9005
rect 7513 8937 7519 8984
rect 7553 8937 7559 8984
rect 7513 8912 7559 8937
rect 7513 8869 7519 8912
rect 7553 8869 7559 8912
rect 7513 8840 7559 8869
rect 7513 8801 7519 8840
rect 7553 8801 7559 8840
rect 7513 8768 7559 8801
rect 7513 8733 7519 8768
rect 7553 8733 7559 8768
rect 7513 8699 7559 8733
rect 7513 8662 7519 8699
rect 7553 8662 7559 8699
rect 7513 8631 7559 8662
rect 7513 8590 7519 8631
rect 7553 8590 7559 8631
rect 7513 8563 7559 8590
rect 7513 8518 7519 8563
rect 7553 8518 7559 8563
rect 7513 8495 7559 8518
rect 7513 8446 7519 8495
rect 7553 8446 7559 8495
rect 7513 8427 7559 8446
rect 7513 8374 7519 8427
rect 7553 8374 7559 8427
rect 7513 8359 7559 8374
rect 7513 8302 7519 8359
rect 7553 8302 7559 8359
rect 7513 8291 7559 8302
rect 7513 8230 7519 8291
rect 7553 8230 7559 8291
rect 7513 8223 7559 8230
rect 7513 8158 7519 8223
rect 7553 8158 7559 8223
rect 7513 8155 7559 8158
rect 7513 8121 7519 8155
rect 7553 8121 7559 8155
rect 7513 8120 7559 8121
rect 7513 8053 7519 8120
rect 7553 8053 7559 8120
rect 7513 8048 7559 8053
rect 7513 7985 7519 8048
rect 7553 7985 7559 8048
rect 7513 7976 7559 7985
rect 7513 7917 7519 7976
rect 7553 7917 7559 7976
rect 7513 7904 7559 7917
rect 7513 7849 7519 7904
rect 7553 7849 7559 7904
rect 7513 7832 7559 7849
rect 7513 7781 7519 7832
rect 7553 7781 7559 7832
rect 7513 7760 7559 7781
rect 7513 7713 7519 7760
rect 7553 7713 7559 7760
rect 7513 7688 7559 7713
rect 7513 7645 7519 7688
rect 7553 7645 7559 7688
rect 7513 7616 7559 7645
rect 7513 7577 7519 7616
rect 7553 7577 7559 7616
rect 7513 7544 7559 7577
rect 7513 7509 7519 7544
rect 7553 7509 7559 7544
rect 7513 7475 7559 7509
rect 7513 7438 7519 7475
rect 7553 7438 7559 7475
rect 7513 7407 7559 7438
rect 7513 7366 7519 7407
rect 7553 7366 7559 7407
rect 7513 7339 7559 7366
rect 7513 7294 7519 7339
rect 7553 7294 7559 7339
rect 7513 7271 7559 7294
rect 7513 7222 7519 7271
rect 7553 7222 7559 7271
rect 7513 7203 7559 7222
rect 7513 7150 7519 7203
rect 7553 7150 7559 7203
rect 7513 7135 7559 7150
rect 7513 7078 7519 7135
rect 7553 7078 7559 7135
rect 7513 7067 7559 7078
rect 7513 7006 7519 7067
rect 7553 7006 7559 7067
rect 7513 6999 7559 7006
rect 7513 6934 7519 6999
rect 7553 6934 7559 6999
rect 7513 6931 7559 6934
rect 7513 6897 7519 6931
rect 7553 6897 7559 6931
rect 7513 6896 7559 6897
rect 7513 6829 7519 6896
rect 7553 6829 7559 6896
rect 7513 6824 7559 6829
rect 7513 6761 7519 6824
rect 7553 6761 7559 6824
rect 7513 6752 7559 6761
rect 7513 6693 7519 6752
rect 7553 6693 7559 6752
rect 7513 6680 7559 6693
rect 7513 6625 7519 6680
rect 7553 6625 7559 6680
rect 7513 6608 7559 6625
rect 7513 6557 7519 6608
rect 7553 6557 7559 6608
rect 7513 6536 7559 6557
rect 7513 6489 7519 6536
rect 7553 6489 7559 6536
rect 7513 6464 7559 6489
rect 7513 6421 7519 6464
rect 7553 6421 7559 6464
rect 7513 6392 7559 6421
rect 7513 6353 7519 6392
rect 7553 6353 7559 6392
rect 7513 6320 7559 6353
rect 7513 6285 7519 6320
rect 7553 6285 7559 6320
rect 7513 6251 7559 6285
rect 7513 6214 7519 6251
rect 7553 6214 7559 6251
rect 7513 6183 7559 6214
rect 7513 6142 7519 6183
rect 7553 6142 7559 6183
rect 7513 6115 7559 6142
rect 7513 6070 7519 6115
rect 7553 6070 7559 6115
rect 7513 6047 7559 6070
rect 7513 5998 7519 6047
rect 7553 5998 7559 6047
rect 7513 5979 7559 5998
rect 7513 5926 7519 5979
rect 7553 5926 7559 5979
rect 7513 5911 7559 5926
rect 7513 5854 7519 5911
rect 7553 5854 7559 5911
rect 7513 5843 7559 5854
rect 7513 5782 7519 5843
rect 7553 5782 7559 5843
rect 7513 5775 7559 5782
rect 7513 5710 7519 5775
rect 7553 5710 7559 5775
rect 7513 5707 7559 5710
rect 7513 5673 7519 5707
rect 7553 5673 7559 5707
rect 7513 5672 7559 5673
rect 7513 5605 7519 5672
rect 7553 5605 7559 5672
rect 7513 5600 7559 5605
rect 7513 5537 7519 5600
rect 7553 5537 7559 5600
rect 7513 5528 7559 5537
rect 7513 5469 7519 5528
rect 7553 5469 7559 5528
rect 7513 5456 7559 5469
rect 7513 5401 7519 5456
rect 7553 5401 7559 5456
rect 7513 5384 7559 5401
rect 7513 5333 7519 5384
rect 7553 5333 7559 5384
rect 7513 5312 7559 5333
rect 7513 5265 7519 5312
rect 7553 5265 7559 5312
rect 7513 5240 7559 5265
rect 7513 5197 7519 5240
rect 7553 5197 7559 5240
rect 7513 5168 7559 5197
rect 7513 5129 7519 5168
rect 7553 5129 7559 5168
rect 7513 5096 7559 5129
rect 7513 5061 7519 5096
rect 7553 5061 7559 5096
rect 7513 5027 7559 5061
rect 7513 4990 7519 5027
rect 7553 4990 7559 5027
rect 7513 4959 7559 4990
rect 7513 4918 7519 4959
rect 7553 4918 7559 4959
rect 7513 4891 7559 4918
rect 7513 4846 7519 4891
rect 7553 4846 7559 4891
rect 7513 4823 7559 4846
rect 7513 4774 7519 4823
rect 7553 4774 7559 4823
rect 7513 4755 7559 4774
rect 7513 4702 7519 4755
rect 7553 4702 7559 4755
rect 7513 4687 7559 4702
rect 7513 4630 7519 4687
rect 7553 4630 7559 4687
rect 7513 4619 7559 4630
rect 7513 4558 7519 4619
rect 7553 4558 7559 4619
rect 7513 4551 7559 4558
rect 7513 4486 7519 4551
rect 7553 4486 7559 4551
rect 7513 4483 7559 4486
rect 7513 4449 7519 4483
rect 7553 4449 7559 4483
rect 7513 4448 7559 4449
rect 7513 4381 7519 4448
rect 7553 4381 7559 4448
rect 7513 4376 7559 4381
rect 7513 4313 7519 4376
rect 7553 4313 7559 4376
rect 7513 4304 7559 4313
rect 7513 4245 7519 4304
rect 7553 4245 7559 4304
rect 7513 4232 7559 4245
rect 7513 4177 7519 4232
rect 7553 4177 7559 4232
rect 7513 4160 7559 4177
rect 7513 4109 7519 4160
rect 7553 4109 7559 4160
rect 7513 4088 7559 4109
rect 7513 4041 7519 4088
rect 7553 4041 7559 4088
rect 7513 4016 7559 4041
rect 7513 3973 7519 4016
rect 7553 3973 7559 4016
rect 7513 3944 7559 3973
rect 7513 3905 7519 3944
rect 7553 3905 7559 3944
rect 7513 3872 7559 3905
rect 7513 3837 7519 3872
rect 7553 3837 7559 3872
rect 7513 3803 7559 3837
rect 7513 3766 7519 3803
rect 7553 3766 7559 3803
rect 7513 3735 7559 3766
rect 7513 3694 7519 3735
rect 7553 3694 7559 3735
rect 7513 3667 7559 3694
rect 7513 3622 7519 3667
rect 7553 3622 7559 3667
rect 7513 3599 7559 3622
rect 7513 3550 7519 3599
rect 7553 3550 7559 3599
rect 7513 3531 7559 3550
rect 7513 3478 7519 3531
rect 7553 3478 7559 3531
rect 7513 3463 7559 3478
rect 7513 3406 7519 3463
rect 7553 3406 7559 3463
rect 7513 3395 7559 3406
rect 7513 3334 7519 3395
rect 7553 3334 7559 3395
rect 7513 3327 7559 3334
rect 7513 3261 7519 3327
rect 7553 3261 7559 3327
rect 7513 3259 7559 3261
rect 7513 3225 7519 3259
rect 7553 3225 7559 3259
rect 7513 3222 7559 3225
rect 7513 3157 7519 3222
rect 7553 3157 7559 3222
rect 7513 3149 7559 3157
rect 7513 3089 7519 3149
rect 7553 3089 7559 3149
rect 7513 3076 7559 3089
rect 7513 3021 7519 3076
rect 7553 3021 7559 3076
rect 7513 3003 7559 3021
rect 7513 2953 7519 3003
rect 7553 2953 7559 3003
rect 7513 2930 7559 2953
rect 7513 2885 7519 2930
rect 7553 2885 7559 2930
rect 7513 2857 7559 2885
rect 7513 2817 7519 2857
rect 7553 2817 7559 2857
rect 7513 2784 7559 2817
rect 7513 2749 7519 2784
rect 7553 2749 7559 2784
rect 7513 2715 7559 2749
rect 7513 2677 7519 2715
rect 7553 2677 7559 2715
rect 7513 2647 7559 2677
rect 7513 2604 7519 2647
rect 7553 2604 7559 2647
rect 7513 2579 7559 2604
rect 7513 2531 7519 2579
rect 7553 2531 7559 2579
rect 7513 2511 7559 2531
rect 7513 2458 7519 2511
rect 7553 2458 7559 2511
rect 7513 2443 7559 2458
rect 7513 2385 7519 2443
rect 7553 2385 7559 2443
rect 7513 2375 7559 2385
rect 7513 2312 7519 2375
rect 7553 2312 7559 2375
rect 7513 2307 7559 2312
rect 7513 2205 7519 2307
rect 7553 2205 7559 2307
rect 7513 2200 7559 2205
rect 7513 2137 7519 2200
rect 7553 2137 7559 2200
rect 7513 2127 7559 2137
rect 7513 2069 7519 2127
rect 7553 2069 7559 2127
rect 7513 2054 7559 2069
rect 7513 2001 7519 2054
rect 7553 2001 7559 2054
rect 7513 1981 7559 2001
rect 7513 1933 7519 1981
rect 7553 1933 7559 1981
rect 7513 1908 7559 1933
rect 7513 1865 7519 1908
rect 7553 1865 7559 1908
rect 7513 1835 7559 1865
rect 7513 1797 7519 1835
rect 7553 1797 7559 1835
rect 7513 1769 7559 1797
rect 4998 1763 7559 1769
rect 4998 1729 5072 1763
rect 5110 1729 5140 1763
rect 5185 1729 5208 1763
rect 5259 1729 5276 1763
rect 5333 1729 5344 1763
rect 5407 1729 5412 1763
rect 5446 1729 5447 1763
rect 5514 1729 5521 1763
rect 5582 1729 5595 1763
rect 5650 1729 5669 1763
rect 5718 1729 5743 1763
rect 5786 1729 5817 1763
rect 5854 1729 5888 1763
rect 5925 1729 5956 1763
rect 5999 1729 6024 1763
rect 6073 1729 6092 1763
rect 6147 1729 6160 1763
rect 6221 1729 6228 1763
rect 6295 1729 6296 1763
rect 6330 1729 6335 1763
rect 6398 1729 6409 1763
rect 6466 1729 6483 1763
rect 6534 1729 6557 1763
rect 6602 1729 6631 1763
rect 6670 1729 6704 1763
rect 6739 1729 6772 1763
rect 6813 1729 6840 1763
rect 6887 1729 6908 1763
rect 6961 1729 6976 1763
rect 7035 1729 7044 1763
rect 7109 1729 7112 1763
rect 7146 1729 7149 1763
rect 7214 1729 7223 1763
rect 7282 1729 7297 1763
rect 7350 1729 7371 1763
rect 7418 1729 7445 1763
rect 7479 1729 7559 1763
rect 4998 1723 7559 1729
rect 7870 2395 7876 17549
rect 9278 2395 9284 17549
rect 7870 2380 7880 2395
rect 7914 2380 8016 2395
rect 8050 2380 8152 2395
rect 8186 2380 8288 2395
rect 8322 2380 8424 2395
rect 8458 2380 8560 2395
rect 8594 2380 8696 2395
rect 8730 2380 8832 2395
rect 8866 2380 8968 2395
rect 9002 2380 9104 2395
rect 9138 2380 9240 2395
rect 9274 2380 9284 2395
rect 7870 2356 9284 2380
rect 7870 2322 7876 2356
rect 7910 2322 7948 2356
rect 7982 2322 8020 2356
rect 8054 2322 8092 2356
rect 8126 2322 8164 2356
rect 8198 2322 8236 2356
rect 8270 2322 8308 2356
rect 8342 2322 8380 2356
rect 8414 2322 8452 2356
rect 8486 2322 8524 2356
rect 8558 2322 8596 2356
rect 8630 2322 8668 2356
rect 8702 2322 8740 2356
rect 8774 2322 8812 2356
rect 8846 2322 8884 2356
rect 8918 2322 8956 2356
rect 8990 2322 9028 2356
rect 9062 2322 9100 2356
rect 9134 2322 9172 2356
rect 9206 2322 9244 2356
rect 9278 2322 9284 2356
rect 7870 2283 9284 2322
rect 7870 2249 7876 2283
rect 7910 2277 7948 2283
rect 7914 2249 7948 2277
rect 7982 2277 8020 2283
rect 7982 2249 8016 2277
rect 8054 2249 8092 2283
rect 8126 2277 8164 2283
rect 8126 2249 8152 2277
rect 8198 2249 8236 2283
rect 8270 2277 8308 2283
rect 8270 2249 8288 2277
rect 8342 2249 8380 2283
rect 8414 2277 8452 2283
rect 8414 2249 8424 2277
rect 8486 2249 8524 2283
rect 8558 2277 8596 2283
rect 8558 2249 8560 2277
rect 7870 2243 7880 2249
rect 7914 2243 8016 2249
rect 8050 2243 8152 2249
rect 8186 2243 8288 2249
rect 8322 2243 8424 2249
rect 8458 2243 8560 2249
rect 8594 2249 8596 2277
rect 8630 2249 8668 2283
rect 8702 2277 8740 2283
rect 8730 2249 8740 2277
rect 8774 2249 8812 2283
rect 8846 2277 8884 2283
rect 8866 2249 8884 2277
rect 8918 2249 8956 2283
rect 8990 2277 9028 2283
rect 9002 2249 9028 2277
rect 9062 2249 9100 2283
rect 9134 2277 9172 2283
rect 9138 2249 9172 2277
rect 9206 2277 9244 2283
rect 9206 2249 9240 2277
rect 9278 2249 9284 2283
rect 8594 2243 8696 2249
rect 8730 2243 8832 2249
rect 8866 2243 8968 2249
rect 9002 2243 9104 2249
rect 9138 2243 9240 2249
rect 9274 2243 9284 2249
rect 7870 2210 9284 2243
rect 7870 2176 7876 2210
rect 7910 2176 7948 2210
rect 7982 2176 8020 2210
rect 8054 2176 8092 2210
rect 8126 2176 8164 2210
rect 8198 2176 8236 2210
rect 8270 2176 8308 2210
rect 8342 2176 8380 2210
rect 8414 2176 8452 2210
rect 8486 2176 8524 2210
rect 8558 2176 8596 2210
rect 8630 2176 8668 2210
rect 8702 2176 8740 2210
rect 8774 2176 8812 2210
rect 8846 2176 8884 2210
rect 8918 2176 8956 2210
rect 8990 2176 9028 2210
rect 9062 2176 9100 2210
rect 9134 2176 9172 2210
rect 9206 2176 9244 2210
rect 9278 2176 9284 2210
rect 7870 2140 9284 2176
rect 7870 2137 7880 2140
rect 7914 2137 8016 2140
rect 8050 2137 8152 2140
rect 8186 2137 8288 2140
rect 8322 2137 8424 2140
rect 8458 2137 8560 2140
rect 7870 2103 7876 2137
rect 7914 2106 7948 2137
rect 7910 2103 7948 2106
rect 7982 2106 8016 2137
rect 7982 2103 8020 2106
rect 8054 2103 8092 2137
rect 8126 2106 8152 2137
rect 8126 2103 8164 2106
rect 8198 2103 8236 2137
rect 8270 2106 8288 2137
rect 8270 2103 8308 2106
rect 8342 2103 8380 2137
rect 8414 2106 8424 2137
rect 8414 2103 8452 2106
rect 8486 2103 8524 2137
rect 8558 2106 8560 2137
rect 8594 2137 8696 2140
rect 8730 2137 8832 2140
rect 8866 2137 8968 2140
rect 9002 2137 9104 2140
rect 9138 2137 9240 2140
rect 9274 2137 9284 2140
rect 8594 2106 8596 2137
rect 8558 2103 8596 2106
rect 8630 2103 8668 2137
rect 8730 2106 8740 2137
rect 8702 2103 8740 2106
rect 8774 2103 8812 2137
rect 8866 2106 8884 2137
rect 8846 2103 8884 2106
rect 8918 2103 8956 2137
rect 9002 2106 9028 2137
rect 8990 2103 9028 2106
rect 9062 2103 9100 2137
rect 9138 2106 9172 2137
rect 9134 2103 9172 2106
rect 9206 2106 9240 2137
rect 9206 2103 9244 2106
rect 9278 2103 9284 2137
rect 7870 2064 9284 2103
rect 7870 2030 7876 2064
rect 7910 2030 7948 2064
rect 7982 2030 8020 2064
rect 8054 2030 8092 2064
rect 8126 2030 8164 2064
rect 8198 2030 8236 2064
rect 8270 2030 8308 2064
rect 8342 2030 8380 2064
rect 8414 2030 8452 2064
rect 8486 2030 8524 2064
rect 8558 2030 8596 2064
rect 8630 2030 8668 2064
rect 8702 2030 8740 2064
rect 8774 2030 8812 2064
rect 8846 2030 8884 2064
rect 8918 2030 8956 2064
rect 8990 2030 9028 2064
rect 9062 2030 9100 2064
rect 9134 2030 9172 2064
rect 9206 2030 9244 2064
rect 9278 2030 9284 2064
rect 7870 2003 9284 2030
rect 7870 1991 7880 2003
rect 7914 1991 8016 2003
rect 8050 1991 8152 2003
rect 8186 1991 8288 2003
rect 8322 1991 8424 2003
rect 8458 1991 8560 2003
rect 7870 1957 7876 1991
rect 7914 1969 7948 1991
rect 7910 1957 7948 1969
rect 7982 1969 8016 1991
rect 7982 1957 8020 1969
rect 8054 1957 8092 1991
rect 8126 1969 8152 1991
rect 8126 1957 8164 1969
rect 8198 1957 8236 1991
rect 8270 1969 8288 1991
rect 8270 1957 8308 1969
rect 8342 1957 8380 1991
rect 8414 1969 8424 1991
rect 8414 1957 8452 1969
rect 8486 1957 8524 1991
rect 8558 1969 8560 1991
rect 8594 1991 8696 2003
rect 8730 1991 8832 2003
rect 8866 1991 8968 2003
rect 9002 1991 9104 2003
rect 9138 1991 9240 2003
rect 9274 1991 9284 2003
rect 8594 1969 8596 1991
rect 8558 1957 8596 1969
rect 8630 1957 8668 1991
rect 8730 1969 8740 1991
rect 8702 1957 8740 1969
rect 8774 1957 8812 1991
rect 8866 1969 8884 1991
rect 8846 1957 8884 1969
rect 8918 1957 8956 1991
rect 9002 1969 9028 1991
rect 8990 1957 9028 1969
rect 9062 1957 9100 1991
rect 9138 1969 9172 1991
rect 9134 1957 9172 1969
rect 9206 1969 9240 1991
rect 9206 1957 9244 1969
rect 9278 1957 9284 1991
rect 7870 1918 9284 1957
rect 7870 1884 7876 1918
rect 7910 1884 7948 1918
rect 7982 1884 8020 1918
rect 8054 1884 8092 1918
rect 8126 1884 8164 1918
rect 8198 1884 8236 1918
rect 8270 1884 8308 1918
rect 8342 1884 8380 1918
rect 8414 1884 8452 1918
rect 8486 1884 8524 1918
rect 8558 1884 8596 1918
rect 8630 1884 8668 1918
rect 8702 1884 8740 1918
rect 8774 1884 8812 1918
rect 8846 1884 8884 1918
rect 8918 1884 8956 1918
rect 8990 1884 9028 1918
rect 9062 1884 9100 1918
rect 9134 1884 9172 1918
rect 9206 1884 9244 1918
rect 9278 1884 9284 1918
rect 7870 1866 9284 1884
rect 7870 1845 7880 1866
rect 7914 1845 8016 1866
rect 8050 1845 8152 1866
rect 8186 1845 8288 1866
rect 8322 1845 8424 1866
rect 8458 1845 8560 1866
rect 7870 1811 7876 1845
rect 7914 1832 7948 1845
rect 7910 1811 7948 1832
rect 7982 1832 8016 1845
rect 7982 1811 8020 1832
rect 8054 1811 8092 1845
rect 8126 1832 8152 1845
rect 8126 1811 8164 1832
rect 8198 1811 8236 1845
rect 8270 1832 8288 1845
rect 8270 1811 8308 1832
rect 8342 1811 8380 1845
rect 8414 1832 8424 1845
rect 8414 1811 8452 1832
rect 8486 1811 8524 1845
rect 8558 1832 8560 1845
rect 8594 1845 8696 1866
rect 8730 1845 8832 1866
rect 8866 1845 8968 1866
rect 9002 1845 9104 1866
rect 9138 1845 9240 1866
rect 9274 1845 9284 1866
rect 8594 1832 8596 1845
rect 8558 1811 8596 1832
rect 8630 1811 8668 1845
rect 8730 1832 8740 1845
rect 8702 1811 8740 1832
rect 8774 1811 8812 1845
rect 8866 1832 8884 1845
rect 8846 1811 8884 1832
rect 8918 1811 8956 1845
rect 9002 1832 9028 1845
rect 8990 1811 9028 1832
rect 9062 1811 9100 1845
rect 9138 1832 9172 1845
rect 9134 1811 9172 1832
rect 9206 1832 9240 1845
rect 9206 1811 9244 1832
rect 9278 1811 9284 1845
rect 7870 1772 9284 1811
rect 7870 1738 7876 1772
rect 7910 1738 7948 1772
rect 7982 1738 8020 1772
rect 8054 1738 8092 1772
rect 8126 1738 8164 1772
rect 8198 1738 8236 1772
rect 8270 1738 8308 1772
rect 8342 1738 8380 1772
rect 8414 1738 8452 1772
rect 8486 1738 8524 1772
rect 8558 1738 8596 1772
rect 8630 1738 8668 1772
rect 8702 1738 8740 1772
rect 8774 1738 8812 1772
rect 8846 1738 8884 1772
rect 8918 1738 8956 1772
rect 8990 1738 9028 1772
rect 9062 1738 9100 1772
rect 9134 1738 9172 1772
rect 9206 1738 9244 1772
rect 9278 1738 9284 1772
rect 7870 1729 9284 1738
rect 1003 1665 1719 1695
rect 315 1626 1719 1665
rect 315 1592 321 1626
rect 355 1592 393 1626
rect 427 1592 465 1626
rect 499 1592 537 1626
rect 571 1592 609 1626
rect 643 1592 681 1626
rect 715 1592 753 1626
rect 787 1592 825 1626
rect 859 1592 897 1626
rect 931 1592 969 1626
rect 1003 1592 1719 1626
rect 315 1558 325 1592
rect 359 1558 461 1592
rect 495 1558 597 1592
rect 631 1558 733 1592
rect 767 1558 869 1592
rect 903 1558 1005 1592
rect 1039 1558 1141 1592
rect 1175 1558 1277 1592
rect 1311 1558 1413 1592
rect 1447 1558 1549 1592
rect 1583 1558 1685 1592
rect 315 1553 1719 1558
rect 315 1519 321 1553
rect 355 1519 393 1553
rect 427 1519 465 1553
rect 499 1519 537 1553
rect 571 1519 609 1553
rect 643 1519 681 1553
rect 715 1519 753 1553
rect 787 1519 825 1553
rect 859 1519 897 1553
rect 931 1519 969 1553
rect 1003 1519 1719 1553
rect 315 1480 1719 1519
rect 315 1446 321 1480
rect 355 1455 393 1480
rect 359 1446 393 1455
rect 427 1455 465 1480
rect 427 1446 461 1455
rect 499 1446 537 1480
rect 571 1455 609 1480
rect 571 1446 597 1455
rect 643 1446 681 1480
rect 715 1455 753 1480
rect 715 1446 733 1455
rect 787 1446 825 1480
rect 859 1455 897 1480
rect 859 1446 869 1455
rect 931 1446 969 1480
rect 1003 1455 1719 1480
rect 1003 1446 1005 1455
rect 315 1421 325 1446
rect 359 1421 461 1446
rect 495 1421 597 1446
rect 631 1421 733 1446
rect 767 1421 869 1446
rect 903 1421 1005 1446
rect 1039 1421 1141 1455
rect 1175 1421 1277 1455
rect 1311 1421 1413 1455
rect 1447 1421 1549 1455
rect 1583 1421 1685 1455
rect 315 1407 1719 1421
rect 315 1373 321 1407
rect 355 1373 393 1407
rect 427 1373 465 1407
rect 499 1373 537 1407
rect 571 1373 609 1407
rect 643 1373 681 1407
rect 715 1373 753 1407
rect 787 1373 825 1407
rect 859 1373 897 1407
rect 931 1373 969 1407
rect 1003 1373 1719 1407
rect 315 1334 1719 1373
rect 315 1300 321 1334
rect 355 1318 393 1334
rect 359 1300 393 1318
rect 427 1318 465 1334
rect 427 1300 461 1318
rect 499 1300 537 1334
rect 571 1318 609 1334
rect 571 1300 597 1318
rect 643 1300 681 1334
rect 715 1318 753 1334
rect 715 1300 733 1318
rect 787 1300 825 1334
rect 859 1318 897 1334
rect 859 1300 869 1318
rect 931 1300 969 1334
rect 1003 1318 1719 1334
rect 1003 1300 1005 1318
rect 315 1284 325 1300
rect 359 1284 461 1300
rect 495 1284 597 1300
rect 631 1284 733 1300
rect 767 1284 869 1300
rect 903 1284 1005 1300
rect 1039 1284 1141 1318
rect 1175 1284 1277 1318
rect 1311 1284 1413 1318
rect 1447 1284 1549 1318
rect 1583 1284 1685 1318
rect 315 1261 1719 1284
rect 315 1227 321 1261
rect 355 1227 393 1261
rect 427 1227 465 1261
rect 499 1227 537 1261
rect 571 1227 609 1261
rect 643 1227 681 1261
rect 715 1227 753 1261
rect 787 1227 825 1261
rect 859 1227 897 1261
rect 931 1227 969 1261
rect 1003 1227 1719 1261
rect 315 1188 1719 1227
rect 315 1154 321 1188
rect 355 1181 393 1188
rect 359 1154 393 1181
rect 427 1181 465 1188
rect 427 1154 461 1181
rect 499 1154 537 1188
rect 571 1181 609 1188
rect 571 1154 597 1181
rect 643 1154 681 1188
rect 715 1181 753 1188
rect 715 1154 733 1181
rect 787 1154 825 1188
rect 859 1181 897 1188
rect 859 1154 869 1181
rect 931 1154 969 1188
rect 1003 1181 1719 1188
rect 1003 1154 1005 1181
rect 315 1147 325 1154
rect 359 1147 461 1154
rect 495 1147 597 1154
rect 631 1147 733 1154
rect 767 1147 869 1154
rect 903 1147 1005 1154
rect 1039 1147 1141 1181
rect 1175 1147 1277 1181
rect 1311 1147 1413 1181
rect 1447 1147 1549 1181
rect 1583 1147 1685 1181
rect 315 1115 1719 1147
rect 315 1081 321 1115
rect 355 1081 393 1115
rect 427 1081 465 1115
rect 499 1081 537 1115
rect 571 1081 609 1115
rect 643 1081 681 1115
rect 715 1081 753 1115
rect 787 1081 825 1115
rect 859 1081 897 1115
rect 931 1081 969 1115
rect 1003 1081 1719 1115
rect 315 1044 1719 1081
rect 315 1042 325 1044
rect 359 1042 461 1044
rect 495 1042 597 1044
rect 631 1042 733 1044
rect 767 1042 869 1044
rect 903 1042 1005 1044
rect 315 1008 321 1042
rect 359 1010 393 1042
rect 355 1008 393 1010
rect 427 1010 461 1042
rect 427 1008 465 1010
rect 499 1008 537 1042
rect 571 1010 597 1042
rect 571 1008 609 1010
rect 643 1008 681 1042
rect 715 1010 733 1042
rect 715 1008 753 1010
rect 787 1008 825 1042
rect 859 1010 869 1042
rect 859 1008 897 1010
rect 931 1008 969 1042
rect 1003 1010 1005 1042
rect 1039 1010 1141 1044
rect 1175 1010 1277 1044
rect 1311 1010 1413 1044
rect 1447 1010 1549 1044
rect 1583 1010 1685 1044
rect 1003 1008 1719 1010
rect 315 969 1719 1008
rect 315 935 321 969
rect 355 935 393 969
rect 427 935 465 969
rect 499 935 537 969
rect 571 935 609 969
rect 643 935 681 969
rect 715 935 753 969
rect 787 935 825 969
rect 859 935 897 969
rect 931 935 969 969
rect 1003 935 1719 969
rect 315 907 1719 935
rect 315 896 325 907
rect 359 896 461 907
rect 495 896 597 907
rect 631 896 733 907
rect 767 896 869 907
rect 903 896 1005 907
rect 315 862 321 896
rect 359 873 393 896
rect 355 862 393 873
rect 427 873 461 896
rect 427 862 465 873
rect 499 862 537 896
rect 571 873 597 896
rect 571 862 609 873
rect 643 862 681 896
rect 715 873 733 896
rect 715 862 753 873
rect 787 862 825 896
rect 859 873 869 896
rect 859 862 897 873
rect 931 862 969 896
rect 1003 873 1005 896
rect 1039 873 1141 907
rect 1175 873 1277 907
rect 1311 873 1413 907
rect 1447 873 1549 907
rect 1583 873 1685 907
rect 1003 862 1719 873
rect 315 823 1719 862
rect 315 789 321 823
rect 355 789 393 823
rect 427 789 465 823
rect 499 789 537 823
rect 571 789 609 823
rect 643 789 681 823
rect 715 789 753 823
rect 787 789 825 823
rect 859 789 897 823
rect 931 789 969 823
rect 1003 789 1719 823
rect 315 770 1719 789
rect 315 750 325 770
rect 359 750 461 770
rect 495 750 597 770
rect 631 750 733 770
rect 767 750 869 770
rect 903 750 1005 770
rect 315 716 321 750
rect 359 736 393 750
rect 355 716 393 736
rect 427 736 461 750
rect 427 716 465 736
rect 499 716 537 750
rect 571 736 597 750
rect 571 716 609 736
rect 643 716 681 750
rect 715 736 733 750
rect 715 716 753 736
rect 787 716 825 750
rect 859 736 869 750
rect 859 716 897 736
rect 931 716 969 750
rect 1003 736 1005 750
rect 1039 736 1141 770
rect 1175 736 1277 770
rect 1311 736 1413 770
rect 1447 736 1549 770
rect 1583 736 1685 770
rect 1003 716 1719 736
rect 315 677 1719 716
rect 315 643 321 677
rect 355 643 393 677
rect 427 643 465 677
rect 499 643 537 677
rect 571 643 609 677
rect 643 643 681 677
rect 715 643 753 677
rect 787 643 825 677
rect 859 643 897 677
rect 931 643 969 677
rect 1003 643 1719 677
rect 315 633 1719 643
rect 315 604 325 633
rect 359 604 461 633
rect 495 604 597 633
rect 631 604 733 633
rect 767 604 869 633
rect 903 604 1005 633
rect 315 570 321 604
rect 359 599 393 604
rect 355 570 393 599
rect 427 599 461 604
rect 427 570 465 599
rect 499 570 537 604
rect 571 599 597 604
rect 571 570 609 599
rect 643 570 681 604
rect 715 599 733 604
rect 715 570 753 599
rect 787 570 825 604
rect 859 599 869 604
rect 859 570 897 599
rect 931 570 969 604
rect 1003 599 1005 604
rect 1039 599 1141 633
rect 1175 599 1277 633
rect 1311 599 1413 633
rect 1447 599 1549 633
rect 1583 599 1685 633
rect 1003 570 1719 599
rect 315 531 1719 570
rect 315 497 321 531
rect 355 497 393 531
rect 427 497 465 531
rect 499 497 537 531
rect 571 497 609 531
rect 643 497 681 531
rect 715 497 753 531
rect 787 497 825 531
rect 859 497 897 531
rect 931 497 969 531
rect 1003 497 1719 531
rect 315 496 1719 497
rect 315 462 325 496
rect 359 462 461 496
rect 495 462 597 496
rect 631 462 733 496
rect 767 462 869 496
rect 903 462 1005 496
rect 1039 462 1141 496
rect 1175 462 1277 496
rect 1311 462 1413 496
rect 1447 462 1549 496
rect 1583 462 1685 496
rect 315 458 1719 462
rect 315 424 321 458
rect 355 424 393 458
rect 427 424 465 458
rect 499 424 537 458
rect 571 424 609 458
rect 643 424 681 458
rect 715 424 753 458
rect 787 424 825 458
rect 859 424 897 458
rect 931 424 969 458
rect 1003 424 1719 458
rect 315 385 1719 424
rect 315 351 321 385
rect 355 359 393 385
rect 359 351 393 359
rect 427 359 465 385
rect 427 351 461 359
rect 499 351 537 385
rect 571 359 609 385
rect 571 351 597 359
rect 643 351 681 385
rect 715 359 753 385
rect 715 351 733 359
rect 787 351 825 385
rect 859 359 897 385
rect 859 351 869 359
rect 931 351 969 385
rect 1003 359 1719 385
rect 1003 351 1005 359
rect 315 325 325 351
rect 359 325 461 351
rect 495 325 597 351
rect 631 325 733 351
rect 767 325 869 351
rect 903 325 1005 351
rect 1039 325 1141 359
rect 1175 325 1277 359
rect 1311 325 1413 359
rect 1447 325 1549 359
rect 1583 325 1685 359
rect 315 312 1719 325
rect 315 278 321 312
rect 355 278 393 312
rect 427 278 465 312
rect 499 278 537 312
rect 571 278 609 312
rect 643 278 681 312
rect 715 278 753 312
rect 787 278 825 312
rect 859 278 897 312
rect 931 278 969 312
rect 1003 278 1719 312
rect 315 239 1719 278
rect 315 205 321 239
rect 355 222 393 239
rect 359 205 393 222
rect 427 222 465 239
rect 427 205 461 222
rect 499 205 537 239
rect 571 222 609 239
rect 571 205 597 222
rect 643 205 681 239
rect 715 222 753 239
rect 715 205 733 222
rect 787 205 825 239
rect 859 222 897 239
rect 859 205 869 222
rect 931 205 969 239
rect 1003 222 1719 239
rect 1003 205 1005 222
rect 315 188 325 205
rect 359 188 461 205
rect 495 188 597 205
rect 631 188 733 205
rect 767 188 869 205
rect 903 188 1005 205
rect 1039 188 1141 222
rect 1175 188 1277 222
rect 1311 188 1413 222
rect 1447 188 1549 222
rect 1583 188 1685 222
rect 315 166 1719 188
rect 315 132 321 166
rect 355 132 393 166
rect 427 132 465 166
rect 499 132 537 166
rect 571 132 609 166
rect 643 132 681 166
rect 715 132 753 166
rect 787 132 825 166
rect 859 132 897 166
rect 931 132 969 166
rect 1003 132 1719 166
rect 315 93 1719 132
rect 315 59 321 93
rect 355 85 393 93
rect 359 59 393 85
rect 427 85 465 93
rect 427 59 461 85
rect 499 59 537 93
rect 571 85 609 93
rect 571 59 597 85
rect 643 59 681 93
rect 715 85 753 93
rect 715 59 733 85
rect 787 59 825 93
rect 859 85 897 93
rect 859 59 869 85
rect 931 59 969 93
rect 1003 85 1719 93
rect 1003 59 1005 85
rect 315 51 325 59
rect 359 51 461 59
rect 495 51 597 59
rect 631 51 733 59
rect 767 51 869 59
rect 903 51 1005 59
rect 1039 51 1141 85
rect 1175 51 1277 85
rect 1311 51 1413 85
rect 1447 51 1549 85
rect 1583 51 1685 85
rect 315 27 1719 51
rect 7870 1699 7880 1729
rect 7914 1699 8016 1729
rect 8050 1699 8152 1729
rect 8186 1699 8288 1729
rect 8322 1699 8424 1729
rect 8458 1699 8560 1729
rect 7870 1665 7876 1699
rect 7914 1695 7948 1699
rect 7910 1665 7948 1695
rect 7982 1695 8016 1699
rect 7982 1665 8020 1695
rect 8054 1665 8092 1699
rect 8126 1695 8152 1699
rect 8126 1665 8164 1695
rect 8198 1665 8236 1699
rect 8270 1695 8288 1699
rect 8270 1665 8308 1695
rect 8342 1665 8380 1699
rect 8414 1695 8424 1699
rect 8414 1665 8452 1695
rect 8486 1665 8524 1699
rect 8558 1695 8560 1699
rect 8594 1699 8696 1729
rect 8730 1699 8832 1729
rect 8866 1699 8968 1729
rect 9002 1699 9104 1729
rect 9138 1699 9240 1729
rect 9274 1699 9284 1729
rect 8594 1695 8596 1699
rect 8558 1665 8596 1695
rect 8630 1665 8668 1699
rect 8730 1695 8740 1699
rect 8702 1665 8740 1695
rect 8774 1665 8812 1699
rect 8866 1695 8884 1699
rect 8846 1665 8884 1695
rect 8918 1665 8956 1699
rect 9002 1695 9028 1699
rect 8990 1665 9028 1695
rect 9062 1665 9100 1699
rect 9138 1695 9172 1699
rect 9134 1665 9172 1695
rect 9206 1695 9240 1699
rect 9206 1665 9244 1695
rect 9278 1665 9284 1699
rect 7870 1626 9284 1665
rect 7870 1592 7876 1626
rect 7910 1592 7948 1626
rect 7982 1592 8020 1626
rect 8054 1592 8092 1626
rect 8126 1592 8164 1626
rect 8198 1592 8236 1626
rect 8270 1592 8308 1626
rect 8342 1592 8380 1626
rect 8414 1592 8452 1626
rect 8486 1592 8524 1626
rect 8558 1592 8596 1626
rect 8630 1592 8668 1626
rect 8702 1592 8740 1626
rect 8774 1592 8812 1626
rect 8846 1592 8884 1626
rect 8918 1592 8956 1626
rect 8990 1592 9028 1626
rect 9062 1592 9100 1626
rect 9134 1592 9172 1626
rect 9206 1592 9244 1626
rect 9278 1592 9284 1626
rect 7870 1558 7880 1592
rect 7914 1558 8016 1592
rect 8050 1558 8152 1592
rect 8186 1558 8288 1592
rect 8322 1558 8424 1592
rect 8458 1558 8560 1592
rect 8594 1558 8696 1592
rect 8730 1558 8832 1592
rect 8866 1558 8968 1592
rect 9002 1558 9104 1592
rect 9138 1558 9240 1592
rect 9274 1558 9284 1592
rect 7870 1553 9284 1558
rect 7870 1519 7876 1553
rect 7910 1519 7948 1553
rect 7982 1519 8020 1553
rect 8054 1519 8092 1553
rect 8126 1519 8164 1553
rect 8198 1519 8236 1553
rect 8270 1519 8308 1553
rect 8342 1519 8380 1553
rect 8414 1519 8452 1553
rect 8486 1519 8524 1553
rect 8558 1519 8596 1553
rect 8630 1519 8668 1553
rect 8702 1519 8740 1553
rect 8774 1519 8812 1553
rect 8846 1519 8884 1553
rect 8918 1519 8956 1553
rect 8990 1519 9028 1553
rect 9062 1519 9100 1553
rect 9134 1519 9172 1553
rect 9206 1519 9244 1553
rect 9278 1519 9284 1553
rect 7870 1480 9284 1519
rect 7870 1446 7876 1480
rect 7910 1455 7948 1480
rect 7914 1446 7948 1455
rect 7982 1455 8020 1480
rect 7982 1446 8016 1455
rect 8054 1446 8092 1480
rect 8126 1455 8164 1480
rect 8126 1446 8152 1455
rect 8198 1446 8236 1480
rect 8270 1455 8308 1480
rect 8270 1446 8288 1455
rect 8342 1446 8380 1480
rect 8414 1455 8452 1480
rect 8414 1446 8424 1455
rect 8486 1446 8524 1480
rect 8558 1455 8596 1480
rect 8558 1446 8560 1455
rect 7870 1421 7880 1446
rect 7914 1421 8016 1446
rect 8050 1421 8152 1446
rect 8186 1421 8288 1446
rect 8322 1421 8424 1446
rect 8458 1421 8560 1446
rect 8594 1446 8596 1455
rect 8630 1446 8668 1480
rect 8702 1455 8740 1480
rect 8730 1446 8740 1455
rect 8774 1446 8812 1480
rect 8846 1455 8884 1480
rect 8866 1446 8884 1455
rect 8918 1446 8956 1480
rect 8990 1455 9028 1480
rect 9002 1446 9028 1455
rect 9062 1446 9100 1480
rect 9134 1455 9172 1480
rect 9138 1446 9172 1455
rect 9206 1455 9244 1480
rect 9206 1446 9240 1455
rect 9278 1446 9284 1480
rect 8594 1421 8696 1446
rect 8730 1421 8832 1446
rect 8866 1421 8968 1446
rect 9002 1421 9104 1446
rect 9138 1421 9240 1446
rect 9274 1421 9284 1446
rect 7870 1407 9284 1421
rect 7870 1373 7876 1407
rect 7910 1373 7948 1407
rect 7982 1373 8020 1407
rect 8054 1373 8092 1407
rect 8126 1373 8164 1407
rect 8198 1373 8236 1407
rect 8270 1373 8308 1407
rect 8342 1373 8380 1407
rect 8414 1373 8452 1407
rect 8486 1373 8524 1407
rect 8558 1373 8596 1407
rect 8630 1373 8668 1407
rect 8702 1373 8740 1407
rect 8774 1373 8812 1407
rect 8846 1373 8884 1407
rect 8918 1373 8956 1407
rect 8990 1373 9028 1407
rect 9062 1373 9100 1407
rect 9134 1373 9172 1407
rect 9206 1373 9244 1407
rect 9278 1373 9284 1407
rect 7870 1334 9284 1373
rect 7870 1300 7876 1334
rect 7910 1318 7948 1334
rect 7914 1300 7948 1318
rect 7982 1318 8020 1334
rect 7982 1300 8016 1318
rect 8054 1300 8092 1334
rect 8126 1318 8164 1334
rect 8126 1300 8152 1318
rect 8198 1300 8236 1334
rect 8270 1318 8308 1334
rect 8270 1300 8288 1318
rect 8342 1300 8380 1334
rect 8414 1318 8452 1334
rect 8414 1300 8424 1318
rect 8486 1300 8524 1334
rect 8558 1318 8596 1334
rect 8558 1300 8560 1318
rect 7870 1284 7880 1300
rect 7914 1284 8016 1300
rect 8050 1284 8152 1300
rect 8186 1284 8288 1300
rect 8322 1284 8424 1300
rect 8458 1284 8560 1300
rect 8594 1300 8596 1318
rect 8630 1300 8668 1334
rect 8702 1318 8740 1334
rect 8730 1300 8740 1318
rect 8774 1300 8812 1334
rect 8846 1318 8884 1334
rect 8866 1300 8884 1318
rect 8918 1300 8956 1334
rect 8990 1318 9028 1334
rect 9002 1300 9028 1318
rect 9062 1300 9100 1334
rect 9134 1318 9172 1334
rect 9138 1300 9172 1318
rect 9206 1318 9244 1334
rect 9206 1300 9240 1318
rect 9278 1300 9284 1334
rect 8594 1284 8696 1300
rect 8730 1284 8832 1300
rect 8866 1284 8968 1300
rect 9002 1284 9104 1300
rect 9138 1284 9240 1300
rect 9274 1284 9284 1300
rect 7870 1261 9284 1284
rect 7870 1227 7876 1261
rect 7910 1227 7948 1261
rect 7982 1227 8020 1261
rect 8054 1227 8092 1261
rect 8126 1227 8164 1261
rect 8198 1227 8236 1261
rect 8270 1227 8308 1261
rect 8342 1227 8380 1261
rect 8414 1227 8452 1261
rect 8486 1227 8524 1261
rect 8558 1227 8596 1261
rect 8630 1227 8668 1261
rect 8702 1227 8740 1261
rect 8774 1227 8812 1261
rect 8846 1227 8884 1261
rect 8918 1227 8956 1261
rect 8990 1227 9028 1261
rect 9062 1227 9100 1261
rect 9134 1227 9172 1261
rect 9206 1227 9244 1261
rect 9278 1227 9284 1261
rect 7870 1188 9284 1227
rect 7870 1154 7876 1188
rect 7910 1181 7948 1188
rect 7914 1154 7948 1181
rect 7982 1181 8020 1188
rect 7982 1154 8016 1181
rect 8054 1154 8092 1188
rect 8126 1181 8164 1188
rect 8126 1154 8152 1181
rect 8198 1154 8236 1188
rect 8270 1181 8308 1188
rect 8270 1154 8288 1181
rect 8342 1154 8380 1188
rect 8414 1181 8452 1188
rect 8414 1154 8424 1181
rect 8486 1154 8524 1188
rect 8558 1181 8596 1188
rect 8558 1154 8560 1181
rect 7870 1147 7880 1154
rect 7914 1147 8016 1154
rect 8050 1147 8152 1154
rect 8186 1147 8288 1154
rect 8322 1147 8424 1154
rect 8458 1147 8560 1154
rect 8594 1154 8596 1181
rect 8630 1154 8668 1188
rect 8702 1181 8740 1188
rect 8730 1154 8740 1181
rect 8774 1154 8812 1188
rect 8846 1181 8884 1188
rect 8866 1154 8884 1181
rect 8918 1154 8956 1188
rect 8990 1181 9028 1188
rect 9002 1154 9028 1181
rect 9062 1154 9100 1188
rect 9134 1181 9172 1188
rect 9138 1154 9172 1181
rect 9206 1181 9244 1188
rect 9206 1154 9240 1181
rect 9278 1154 9284 1188
rect 8594 1147 8696 1154
rect 8730 1147 8832 1154
rect 8866 1147 8968 1154
rect 9002 1147 9104 1154
rect 9138 1147 9240 1154
rect 9274 1147 9284 1154
rect 7870 1115 9284 1147
rect 7870 1081 7876 1115
rect 7910 1081 7948 1115
rect 7982 1081 8020 1115
rect 8054 1081 8092 1115
rect 8126 1081 8164 1115
rect 8198 1081 8236 1115
rect 8270 1081 8308 1115
rect 8342 1081 8380 1115
rect 8414 1081 8452 1115
rect 8486 1081 8524 1115
rect 8558 1081 8596 1115
rect 8630 1081 8668 1115
rect 8702 1081 8740 1115
rect 8774 1081 8812 1115
rect 8846 1081 8884 1115
rect 8918 1081 8956 1115
rect 8990 1081 9028 1115
rect 9062 1081 9100 1115
rect 9134 1081 9172 1115
rect 9206 1081 9244 1115
rect 9278 1081 9284 1115
rect 7870 1044 9284 1081
rect 7870 1042 7880 1044
rect 7914 1042 8016 1044
rect 8050 1042 8152 1044
rect 8186 1042 8288 1044
rect 8322 1042 8424 1044
rect 8458 1042 8560 1044
rect 7870 1008 7876 1042
rect 7914 1010 7948 1042
rect 7910 1008 7948 1010
rect 7982 1010 8016 1042
rect 7982 1008 8020 1010
rect 8054 1008 8092 1042
rect 8126 1010 8152 1042
rect 8126 1008 8164 1010
rect 8198 1008 8236 1042
rect 8270 1010 8288 1042
rect 8270 1008 8308 1010
rect 8342 1008 8380 1042
rect 8414 1010 8424 1042
rect 8414 1008 8452 1010
rect 8486 1008 8524 1042
rect 8558 1010 8560 1042
rect 8594 1042 8696 1044
rect 8730 1042 8832 1044
rect 8866 1042 8968 1044
rect 9002 1042 9104 1044
rect 9138 1042 9240 1044
rect 9274 1042 9284 1044
rect 8594 1010 8596 1042
rect 8558 1008 8596 1010
rect 8630 1008 8668 1042
rect 8730 1010 8740 1042
rect 8702 1008 8740 1010
rect 8774 1008 8812 1042
rect 8866 1010 8884 1042
rect 8846 1008 8884 1010
rect 8918 1008 8956 1042
rect 9002 1010 9028 1042
rect 8990 1008 9028 1010
rect 9062 1008 9100 1042
rect 9138 1010 9172 1042
rect 9134 1008 9172 1010
rect 9206 1010 9240 1042
rect 9206 1008 9244 1010
rect 9278 1008 9284 1042
rect 7870 969 9284 1008
rect 7870 935 7876 969
rect 7910 935 7948 969
rect 7982 935 8020 969
rect 8054 935 8092 969
rect 8126 935 8164 969
rect 8198 935 8236 969
rect 8270 935 8308 969
rect 8342 935 8380 969
rect 8414 935 8452 969
rect 8486 935 8524 969
rect 8558 935 8596 969
rect 8630 935 8668 969
rect 8702 935 8740 969
rect 8774 935 8812 969
rect 8846 935 8884 969
rect 8918 935 8956 969
rect 8990 935 9028 969
rect 9062 935 9100 969
rect 9134 935 9172 969
rect 9206 935 9244 969
rect 9278 935 9284 969
rect 7870 907 9284 935
rect 7870 896 7880 907
rect 7914 896 8016 907
rect 8050 896 8152 907
rect 8186 896 8288 907
rect 8322 896 8424 907
rect 8458 896 8560 907
rect 7870 862 7876 896
rect 7914 873 7948 896
rect 7910 862 7948 873
rect 7982 873 8016 896
rect 7982 862 8020 873
rect 8054 862 8092 896
rect 8126 873 8152 896
rect 8126 862 8164 873
rect 8198 862 8236 896
rect 8270 873 8288 896
rect 8270 862 8308 873
rect 8342 862 8380 896
rect 8414 873 8424 896
rect 8414 862 8452 873
rect 8486 862 8524 896
rect 8558 873 8560 896
rect 8594 896 8696 907
rect 8730 896 8832 907
rect 8866 896 8968 907
rect 9002 896 9104 907
rect 9138 896 9240 907
rect 9274 896 9284 907
rect 8594 873 8596 896
rect 8558 862 8596 873
rect 8630 862 8668 896
rect 8730 873 8740 896
rect 8702 862 8740 873
rect 8774 862 8812 896
rect 8866 873 8884 896
rect 8846 862 8884 873
rect 8918 862 8956 896
rect 9002 873 9028 896
rect 8990 862 9028 873
rect 9062 862 9100 896
rect 9138 873 9172 896
rect 9134 862 9172 873
rect 9206 873 9240 896
rect 9206 862 9244 873
rect 9278 862 9284 896
rect 7870 823 9284 862
rect 7870 789 7876 823
rect 7910 789 7948 823
rect 7982 789 8020 823
rect 8054 789 8092 823
rect 8126 789 8164 823
rect 8198 789 8236 823
rect 8270 789 8308 823
rect 8342 789 8380 823
rect 8414 789 8452 823
rect 8486 789 8524 823
rect 8558 789 8596 823
rect 8630 789 8668 823
rect 8702 789 8740 823
rect 8774 789 8812 823
rect 8846 789 8884 823
rect 8918 789 8956 823
rect 8990 789 9028 823
rect 9062 789 9100 823
rect 9134 789 9172 823
rect 9206 789 9244 823
rect 9278 789 9284 823
rect 7870 770 9284 789
rect 7870 750 7880 770
rect 7914 750 8016 770
rect 8050 750 8152 770
rect 8186 750 8288 770
rect 8322 750 8424 770
rect 8458 750 8560 770
rect 7870 716 7876 750
rect 7914 736 7948 750
rect 7910 716 7948 736
rect 7982 736 8016 750
rect 7982 716 8020 736
rect 8054 716 8092 750
rect 8126 736 8152 750
rect 8126 716 8164 736
rect 8198 716 8236 750
rect 8270 736 8288 750
rect 8270 716 8308 736
rect 8342 716 8380 750
rect 8414 736 8424 750
rect 8414 716 8452 736
rect 8486 716 8524 750
rect 8558 736 8560 750
rect 8594 750 8696 770
rect 8730 750 8832 770
rect 8866 750 8968 770
rect 9002 750 9104 770
rect 9138 750 9240 770
rect 9274 750 9284 770
rect 8594 736 8596 750
rect 8558 716 8596 736
rect 8630 716 8668 750
rect 8730 736 8740 750
rect 8702 716 8740 736
rect 8774 716 8812 750
rect 8866 736 8884 750
rect 8846 716 8884 736
rect 8918 716 8956 750
rect 9002 736 9028 750
rect 8990 716 9028 736
rect 9062 716 9100 750
rect 9138 736 9172 750
rect 9134 716 9172 736
rect 9206 736 9240 750
rect 9206 716 9244 736
rect 9278 716 9284 750
rect 7870 677 9284 716
rect 7870 643 7876 677
rect 7910 643 7948 677
rect 7982 643 8020 677
rect 8054 643 8092 677
rect 8126 643 8164 677
rect 8198 643 8236 677
rect 8270 643 8308 677
rect 8342 643 8380 677
rect 8414 643 8452 677
rect 8486 643 8524 677
rect 8558 643 8596 677
rect 8630 643 8668 677
rect 8702 643 8740 677
rect 8774 643 8812 677
rect 8846 643 8884 677
rect 8918 643 8956 677
rect 8990 643 9028 677
rect 9062 643 9100 677
rect 9134 643 9172 677
rect 9206 643 9244 677
rect 9278 643 9284 677
rect 7870 633 9284 643
rect 7870 604 7880 633
rect 7914 604 8016 633
rect 8050 604 8152 633
rect 8186 604 8288 633
rect 8322 604 8424 633
rect 8458 604 8560 633
rect 7870 570 7876 604
rect 7914 599 7948 604
rect 7910 570 7948 599
rect 7982 599 8016 604
rect 7982 570 8020 599
rect 8054 570 8092 604
rect 8126 599 8152 604
rect 8126 570 8164 599
rect 8198 570 8236 604
rect 8270 599 8288 604
rect 8270 570 8308 599
rect 8342 570 8380 604
rect 8414 599 8424 604
rect 8414 570 8452 599
rect 8486 570 8524 604
rect 8558 599 8560 604
rect 8594 604 8696 633
rect 8730 604 8832 633
rect 8866 604 8968 633
rect 9002 604 9104 633
rect 9138 604 9240 633
rect 9274 604 9284 633
rect 8594 599 8596 604
rect 8558 570 8596 599
rect 8630 570 8668 604
rect 8730 599 8740 604
rect 8702 570 8740 599
rect 8774 570 8812 604
rect 8866 599 8884 604
rect 8846 570 8884 599
rect 8918 570 8956 604
rect 9002 599 9028 604
rect 8990 570 9028 599
rect 9062 570 9100 604
rect 9138 599 9172 604
rect 9134 570 9172 599
rect 9206 599 9240 604
rect 9206 570 9244 599
rect 9278 570 9284 604
rect 7870 531 9284 570
rect 7870 497 7876 531
rect 7910 497 7948 531
rect 7982 497 8020 531
rect 8054 497 8092 531
rect 8126 497 8164 531
rect 8198 497 8236 531
rect 8270 497 8308 531
rect 8342 497 8380 531
rect 8414 497 8452 531
rect 8486 497 8524 531
rect 8558 497 8596 531
rect 8630 497 8668 531
rect 8702 497 8740 531
rect 8774 497 8812 531
rect 8846 497 8884 531
rect 8918 497 8956 531
rect 8990 497 9028 531
rect 9062 497 9100 531
rect 9134 497 9172 531
rect 9206 497 9244 531
rect 9278 497 9284 531
rect 7870 496 9284 497
rect 7870 462 7880 496
rect 7914 462 8016 496
rect 8050 462 8152 496
rect 8186 462 8288 496
rect 8322 462 8424 496
rect 8458 462 8560 496
rect 8594 462 8696 496
rect 8730 462 8832 496
rect 8866 462 8968 496
rect 9002 462 9104 496
rect 9138 462 9240 496
rect 9274 462 9284 496
rect 7870 458 9284 462
rect 7870 424 7876 458
rect 7910 424 7948 458
rect 7982 424 8020 458
rect 8054 424 8092 458
rect 8126 424 8164 458
rect 8198 424 8236 458
rect 8270 424 8308 458
rect 8342 424 8380 458
rect 8414 424 8452 458
rect 8486 424 8524 458
rect 8558 424 8596 458
rect 8630 424 8668 458
rect 8702 424 8740 458
rect 8774 424 8812 458
rect 8846 424 8884 458
rect 8918 424 8956 458
rect 8990 424 9028 458
rect 9062 424 9100 458
rect 9134 424 9172 458
rect 9206 424 9244 458
rect 9278 424 9284 458
rect 7870 385 9284 424
rect 7870 351 7876 385
rect 7910 359 7948 385
rect 7914 351 7948 359
rect 7982 359 8020 385
rect 7982 351 8016 359
rect 8054 351 8092 385
rect 8126 359 8164 385
rect 8126 351 8152 359
rect 8198 351 8236 385
rect 8270 359 8308 385
rect 8270 351 8288 359
rect 8342 351 8380 385
rect 8414 359 8452 385
rect 8414 351 8424 359
rect 8486 351 8524 385
rect 8558 359 8596 385
rect 8558 351 8560 359
rect 7870 325 7880 351
rect 7914 325 8016 351
rect 8050 325 8152 351
rect 8186 325 8288 351
rect 8322 325 8424 351
rect 8458 325 8560 351
rect 8594 351 8596 359
rect 8630 351 8668 385
rect 8702 359 8740 385
rect 8730 351 8740 359
rect 8774 351 8812 385
rect 8846 359 8884 385
rect 8866 351 8884 359
rect 8918 351 8956 385
rect 8990 359 9028 385
rect 9002 351 9028 359
rect 9062 351 9100 385
rect 9134 359 9172 385
rect 9138 351 9172 359
rect 9206 359 9244 385
rect 9206 351 9240 359
rect 9278 351 9284 385
rect 8594 325 8696 351
rect 8730 325 8832 351
rect 8866 325 8968 351
rect 9002 325 9104 351
rect 9138 325 9240 351
rect 9274 325 9284 351
rect 7870 312 9284 325
rect 7870 278 7876 312
rect 7910 278 7948 312
rect 7982 278 8020 312
rect 8054 278 8092 312
rect 8126 278 8164 312
rect 8198 278 8236 312
rect 8270 278 8308 312
rect 8342 278 8380 312
rect 8414 278 8452 312
rect 8486 278 8524 312
rect 8558 278 8596 312
rect 8630 278 8668 312
rect 8702 278 8740 312
rect 8774 278 8812 312
rect 8846 278 8884 312
rect 8918 278 8956 312
rect 8990 278 9028 312
rect 9062 278 9100 312
rect 9134 278 9172 312
rect 9206 278 9244 312
rect 9278 278 9284 312
rect 7870 239 9284 278
rect 7870 205 7876 239
rect 7910 222 7948 239
rect 7914 205 7948 222
rect 7982 222 8020 239
rect 7982 205 8016 222
rect 8054 205 8092 239
rect 8126 222 8164 239
rect 8126 205 8152 222
rect 8198 205 8236 239
rect 8270 222 8308 239
rect 8270 205 8288 222
rect 8342 205 8380 239
rect 8414 222 8452 239
rect 8414 205 8424 222
rect 8486 205 8524 239
rect 8558 222 8596 239
rect 8558 205 8560 222
rect 7870 188 7880 205
rect 7914 188 8016 205
rect 8050 188 8152 205
rect 8186 188 8288 205
rect 8322 188 8424 205
rect 8458 188 8560 205
rect 8594 205 8596 222
rect 8630 205 8668 239
rect 8702 222 8740 239
rect 8730 205 8740 222
rect 8774 205 8812 239
rect 8846 222 8884 239
rect 8866 205 8884 222
rect 8918 205 8956 239
rect 8990 222 9028 239
rect 9002 205 9028 222
rect 9062 205 9100 239
rect 9134 222 9172 239
rect 9138 205 9172 222
rect 9206 222 9244 239
rect 9206 205 9240 222
rect 9278 205 9284 239
rect 8594 188 8696 205
rect 8730 188 8832 205
rect 8866 188 8968 205
rect 9002 188 9104 205
rect 9138 188 9240 205
rect 9274 188 9284 205
rect 7870 166 9284 188
rect 7870 132 7876 166
rect 7910 132 7948 166
rect 7982 132 8020 166
rect 8054 132 8092 166
rect 8126 132 8164 166
rect 8198 132 8236 166
rect 8270 132 8308 166
rect 8342 132 8380 166
rect 8414 132 8452 166
rect 8486 132 8524 166
rect 8558 132 8596 166
rect 8630 132 8668 166
rect 8702 132 8740 166
rect 8774 132 8812 166
rect 8846 132 8884 166
rect 8918 132 8956 166
rect 8990 132 9028 166
rect 9062 132 9100 166
rect 9134 132 9172 166
rect 9206 132 9244 166
rect 9278 132 9284 166
rect 7870 93 9284 132
rect 7870 59 7876 93
rect 7910 85 7948 93
rect 7914 59 7948 85
rect 7982 85 8020 93
rect 7982 59 8016 85
rect 8054 59 8092 93
rect 8126 85 8164 93
rect 8126 59 8152 85
rect 8198 59 8236 93
rect 8270 85 8308 93
rect 8270 59 8288 85
rect 8342 59 8380 93
rect 8414 85 8452 93
rect 8414 59 8424 85
rect 8486 59 8524 93
rect 8558 85 8596 93
rect 8558 59 8560 85
rect 7870 51 7880 59
rect 7914 51 8016 59
rect 8050 51 8152 59
rect 8186 51 8288 59
rect 8322 51 8424 59
rect 8458 51 8560 59
rect 8594 59 8596 85
rect 8630 59 8668 93
rect 8702 85 8740 93
rect 8730 59 8740 85
rect 8774 59 8812 93
rect 8846 85 8884 93
rect 8866 59 8884 85
rect 8918 59 8956 93
rect 8990 85 9028 93
rect 9002 59 9028 85
rect 9062 59 9100 93
rect 9134 85 9172 93
rect 9138 59 9172 85
rect 9206 85 9244 93
rect 9206 59 9240 85
rect 9278 59 9284 93
rect 8594 51 8696 59
rect 8730 51 8832 59
rect 8866 51 8968 59
rect 9002 51 9104 59
rect 9138 51 9240 59
rect 9274 51 9284 59
rect 7870 27 9284 51
<< viali >>
rect 321 39917 325 39943
rect 325 39917 359 39943
rect 359 39917 461 39943
rect 461 39917 495 39943
rect 495 39917 597 39943
rect 597 39917 631 39943
rect 631 39917 733 39943
rect 733 39917 767 39943
rect 767 39917 869 39943
rect 869 39917 903 39943
rect 903 39917 1005 39943
rect 1005 39917 1039 39943
rect 1039 39917 1141 39943
rect 1141 39917 1175 39943
rect 1175 39917 1277 39943
rect 1277 39917 1311 39943
rect 1311 39917 1413 39943
rect 1413 39917 1447 39943
rect 1447 39917 1549 39943
rect 1549 39917 1583 39943
rect 1583 39917 1685 39943
rect 1685 39917 1719 39943
rect 1719 39917 1723 39943
rect 321 39815 1723 39917
rect 321 39781 325 39815
rect 325 39781 359 39815
rect 359 39781 461 39815
rect 461 39781 495 39815
rect 495 39781 597 39815
rect 597 39781 631 39815
rect 631 39781 733 39815
rect 733 39781 767 39815
rect 767 39781 869 39815
rect 869 39781 903 39815
rect 903 39781 1005 39815
rect 1005 39781 1039 39815
rect 1039 39781 1141 39815
rect 1141 39781 1175 39815
rect 1175 39781 1277 39815
rect 1277 39781 1311 39815
rect 1311 39781 1413 39815
rect 1413 39781 1447 39815
rect 1447 39781 1549 39815
rect 1549 39781 1583 39815
rect 1583 39781 1685 39815
rect 1685 39781 1719 39815
rect 1719 39781 1723 39815
rect 321 39679 1723 39781
rect 321 39645 325 39679
rect 325 39645 359 39679
rect 359 39645 461 39679
rect 461 39645 495 39679
rect 495 39645 597 39679
rect 597 39645 631 39679
rect 631 39645 733 39679
rect 733 39645 767 39679
rect 767 39645 869 39679
rect 869 39645 903 39679
rect 903 39645 1005 39679
rect 1005 39645 1039 39679
rect 1039 39645 1141 39679
rect 1141 39645 1175 39679
rect 1175 39645 1277 39679
rect 1277 39645 1311 39679
rect 1311 39645 1413 39679
rect 1413 39645 1447 39679
rect 1447 39645 1549 39679
rect 1549 39645 1583 39679
rect 1583 39645 1685 39679
rect 1685 39645 1719 39679
rect 1719 39645 1723 39679
rect 321 39543 1723 39645
rect 321 39509 325 39543
rect 325 39509 359 39543
rect 359 39509 461 39543
rect 461 39509 495 39543
rect 495 39509 597 39543
rect 597 39509 631 39543
rect 631 39509 733 39543
rect 733 39509 767 39543
rect 767 39509 869 39543
rect 869 39509 903 39543
rect 903 39509 1005 39543
rect 1005 39509 1039 39543
rect 1039 39509 1141 39543
rect 1141 39509 1175 39543
rect 1175 39509 1277 39543
rect 1277 39509 1311 39543
rect 1311 39509 1413 39543
rect 1413 39509 1447 39543
rect 1447 39509 1549 39543
rect 1549 39509 1583 39543
rect 1583 39509 1685 39543
rect 1685 39509 1719 39543
rect 1719 39509 1723 39543
rect 321 39407 1723 39509
rect 321 39373 325 39407
rect 325 39373 359 39407
rect 359 39373 461 39407
rect 461 39373 495 39407
rect 495 39373 597 39407
rect 597 39373 631 39407
rect 631 39373 733 39407
rect 733 39373 767 39407
rect 767 39373 869 39407
rect 869 39373 903 39407
rect 903 39373 1005 39407
rect 1005 39373 1039 39407
rect 1039 39373 1141 39407
rect 1141 39373 1175 39407
rect 1175 39373 1277 39407
rect 1277 39373 1311 39407
rect 1311 39373 1413 39407
rect 1413 39373 1447 39407
rect 1447 39373 1549 39407
rect 1549 39373 1583 39407
rect 1583 39373 1685 39407
rect 1685 39373 1719 39407
rect 1719 39373 1723 39407
rect 321 39271 1723 39373
rect 321 39237 325 39271
rect 325 39237 359 39271
rect 359 39237 461 39271
rect 461 39237 495 39271
rect 495 39237 597 39271
rect 597 39237 631 39271
rect 631 39237 733 39271
rect 733 39237 767 39271
rect 767 39237 869 39271
rect 869 39237 903 39271
rect 903 39237 1005 39271
rect 1005 39237 1039 39271
rect 1039 39237 1141 39271
rect 1141 39237 1175 39271
rect 1175 39237 1277 39271
rect 1277 39237 1311 39271
rect 1311 39237 1413 39271
rect 1413 39237 1447 39271
rect 1447 39237 1549 39271
rect 1549 39237 1583 39271
rect 1583 39237 1685 39271
rect 1685 39237 1719 39271
rect 1719 39237 1723 39271
rect 321 39135 1723 39237
rect 321 39101 325 39135
rect 325 39101 359 39135
rect 359 39101 461 39135
rect 461 39101 495 39135
rect 495 39101 597 39135
rect 597 39101 631 39135
rect 631 39101 733 39135
rect 733 39101 767 39135
rect 767 39101 869 39135
rect 869 39101 903 39135
rect 903 39101 1005 39135
rect 1005 39101 1039 39135
rect 1039 39101 1141 39135
rect 1141 39101 1175 39135
rect 1175 39101 1277 39135
rect 1277 39101 1311 39135
rect 1311 39101 1413 39135
rect 1413 39101 1447 39135
rect 1447 39101 1549 39135
rect 1549 39101 1583 39135
rect 1583 39101 1685 39135
rect 1685 39101 1719 39135
rect 1719 39101 1723 39135
rect 321 38999 1723 39101
rect 321 38965 325 38999
rect 325 38965 359 38999
rect 359 38965 461 38999
rect 461 38965 495 38999
rect 495 38965 597 38999
rect 597 38965 631 38999
rect 631 38965 733 38999
rect 733 38965 767 38999
rect 767 38965 869 38999
rect 869 38965 903 38999
rect 903 38965 1005 38999
rect 1005 38965 1039 38999
rect 1039 38965 1141 38999
rect 1141 38965 1175 38999
rect 1175 38965 1277 38999
rect 1277 38965 1311 38999
rect 1311 38965 1413 38999
rect 1413 38965 1447 38999
rect 1447 38965 1549 38999
rect 1549 38965 1583 38999
rect 1583 38965 1685 38999
rect 1685 38965 1719 38999
rect 1719 38965 1723 38999
rect 321 38863 1723 38965
rect 321 38829 325 38863
rect 325 38829 359 38863
rect 359 38829 461 38863
rect 461 38829 495 38863
rect 495 38829 597 38863
rect 597 38829 631 38863
rect 631 38829 733 38863
rect 733 38829 767 38863
rect 767 38829 869 38863
rect 869 38829 903 38863
rect 903 38829 1005 38863
rect 1005 38829 1039 38863
rect 1039 38829 1141 38863
rect 1141 38829 1175 38863
rect 1175 38829 1277 38863
rect 1277 38829 1311 38863
rect 1311 38829 1413 38863
rect 1413 38829 1447 38863
rect 1447 38829 1549 38863
rect 1549 38829 1583 38863
rect 1583 38829 1685 38863
rect 1685 38829 1719 38863
rect 1719 38829 1723 38863
rect 321 38727 1723 38829
rect 321 38693 325 38727
rect 325 38693 359 38727
rect 359 38693 461 38727
rect 461 38693 495 38727
rect 495 38693 597 38727
rect 597 38693 631 38727
rect 631 38693 733 38727
rect 733 38693 767 38727
rect 767 38693 869 38727
rect 869 38693 903 38727
rect 903 38693 1005 38727
rect 1005 38693 1039 38727
rect 1039 38693 1141 38727
rect 1141 38693 1175 38727
rect 1175 38693 1277 38727
rect 1277 38693 1311 38727
rect 1311 38693 1413 38727
rect 1413 38693 1447 38727
rect 1447 38693 1549 38727
rect 1549 38693 1583 38727
rect 1583 38693 1685 38727
rect 1685 38693 1719 38727
rect 1719 38693 1723 38727
rect 321 38591 1723 38693
rect 321 38557 325 38591
rect 325 38557 359 38591
rect 359 38557 461 38591
rect 461 38557 495 38591
rect 495 38557 597 38591
rect 597 38557 631 38591
rect 631 38557 733 38591
rect 733 38557 767 38591
rect 767 38557 869 38591
rect 869 38557 903 38591
rect 903 38557 1005 38591
rect 1005 38557 1039 38591
rect 1039 38557 1141 38591
rect 1141 38557 1175 38591
rect 1175 38557 1277 38591
rect 1277 38557 1311 38591
rect 1311 38557 1413 38591
rect 1413 38557 1447 38591
rect 1447 38557 1549 38591
rect 1549 38557 1583 38591
rect 1583 38557 1685 38591
rect 1685 38557 1719 38591
rect 1719 38557 1723 38591
rect 321 38455 1723 38557
rect 321 38421 325 38455
rect 325 38421 359 38455
rect 359 38421 461 38455
rect 461 38421 495 38455
rect 495 38421 597 38455
rect 597 38421 631 38455
rect 631 38421 733 38455
rect 733 38421 767 38455
rect 767 38421 869 38455
rect 869 38421 903 38455
rect 903 38421 1005 38455
rect 1005 38421 1039 38455
rect 1039 38421 1141 38455
rect 1141 38421 1175 38455
rect 1175 38421 1277 38455
rect 1277 38421 1311 38455
rect 1311 38421 1413 38455
rect 1413 38421 1447 38455
rect 1447 38421 1549 38455
rect 1549 38421 1583 38455
rect 1583 38421 1685 38455
rect 1685 38421 1719 38455
rect 1719 38421 1723 38455
rect 321 38319 1723 38421
rect 321 38285 325 38319
rect 325 38285 359 38319
rect 359 38285 461 38319
rect 461 38285 495 38319
rect 495 38285 597 38319
rect 597 38285 631 38319
rect 631 38285 733 38319
rect 733 38285 767 38319
rect 767 38285 869 38319
rect 869 38285 903 38319
rect 903 38285 1005 38319
rect 1005 38285 1039 38319
rect 1039 38285 1141 38319
rect 1141 38285 1175 38319
rect 1175 38285 1277 38319
rect 1277 38285 1311 38319
rect 1311 38285 1413 38319
rect 1413 38285 1447 38319
rect 1447 38285 1549 38319
rect 1549 38285 1583 38319
rect 1583 38285 1685 38319
rect 1685 38285 1719 38319
rect 1719 38285 1723 38319
rect 321 38183 1723 38285
rect 321 38149 325 38183
rect 325 38149 359 38183
rect 359 38149 461 38183
rect 461 38149 495 38183
rect 495 38149 597 38183
rect 597 38149 631 38183
rect 631 38149 733 38183
rect 733 38149 767 38183
rect 767 38149 869 38183
rect 869 38149 903 38183
rect 903 38149 1005 38183
rect 1005 38149 1039 38183
rect 1039 38149 1141 38183
rect 1141 38149 1175 38183
rect 1175 38149 1277 38183
rect 1277 38149 1311 38183
rect 1311 38149 1413 38183
rect 1413 38149 1447 38183
rect 1447 38149 1549 38183
rect 1549 38149 1583 38183
rect 1583 38149 1685 38183
rect 1685 38149 1719 38183
rect 1719 38149 1723 38183
rect 321 38047 1723 38149
rect 321 38013 325 38047
rect 325 38013 359 38047
rect 359 38013 461 38047
rect 461 38013 495 38047
rect 495 38013 597 38047
rect 597 38013 631 38047
rect 631 38013 733 38047
rect 733 38013 767 38047
rect 767 38013 869 38047
rect 869 38013 903 38047
rect 903 38013 1005 38047
rect 1005 38013 1039 38047
rect 1039 38013 1141 38047
rect 1141 38013 1175 38047
rect 1175 38013 1277 38047
rect 1277 38013 1311 38047
rect 1311 38013 1413 38047
rect 1413 38013 1447 38047
rect 1447 38013 1549 38047
rect 1549 38013 1583 38047
rect 1583 38013 1685 38047
rect 1685 38013 1719 38047
rect 1719 38013 1723 38047
rect 321 37911 1723 38013
rect 321 37877 325 37911
rect 325 37877 359 37911
rect 359 37877 461 37911
rect 461 37877 495 37911
rect 495 37877 597 37911
rect 597 37877 631 37911
rect 631 37877 733 37911
rect 733 37877 767 37911
rect 767 37877 869 37911
rect 869 37877 903 37911
rect 903 37877 1005 37911
rect 1005 37877 1039 37911
rect 1039 37877 1141 37911
rect 1141 37877 1175 37911
rect 1175 37877 1277 37911
rect 1277 37877 1311 37911
rect 1311 37877 1413 37911
rect 1413 37877 1447 37911
rect 1447 37877 1549 37911
rect 1549 37877 1583 37911
rect 1583 37877 1685 37911
rect 1685 37877 1719 37911
rect 1719 37877 1723 37911
rect 321 37775 1723 37877
rect 321 37741 325 37775
rect 325 37741 359 37775
rect 359 37741 461 37775
rect 461 37741 495 37775
rect 495 37741 597 37775
rect 597 37741 631 37775
rect 631 37741 733 37775
rect 733 37741 767 37775
rect 767 37741 869 37775
rect 869 37741 903 37775
rect 903 37741 1005 37775
rect 1005 37741 1039 37775
rect 1039 37741 1141 37775
rect 1141 37741 1175 37775
rect 1175 37741 1277 37775
rect 1277 37741 1311 37775
rect 1311 37741 1413 37775
rect 1413 37741 1447 37775
rect 1447 37741 1549 37775
rect 1549 37741 1583 37775
rect 1583 37741 1685 37775
rect 1685 37741 1719 37775
rect 1719 37741 1723 37775
rect 321 37639 1723 37741
rect 321 37605 325 37639
rect 325 37605 359 37639
rect 359 37605 461 37639
rect 461 37605 495 37639
rect 495 37605 597 37639
rect 597 37605 631 37639
rect 631 37605 733 37639
rect 733 37605 767 37639
rect 767 37605 869 37639
rect 869 37605 903 37639
rect 903 37605 1005 37639
rect 1005 37605 1039 37639
rect 1039 37605 1141 37639
rect 1141 37605 1175 37639
rect 1175 37605 1277 37639
rect 1277 37605 1311 37639
rect 1311 37605 1413 37639
rect 1413 37605 1447 37639
rect 1447 37605 1549 37639
rect 1549 37605 1583 37639
rect 1583 37605 1685 37639
rect 1685 37605 1719 37639
rect 1719 37605 1723 37639
rect 321 37503 1723 37605
rect 321 37469 325 37503
rect 325 37469 359 37503
rect 359 37469 461 37503
rect 461 37469 495 37503
rect 495 37469 597 37503
rect 597 37469 631 37503
rect 631 37469 733 37503
rect 733 37469 767 37503
rect 767 37469 869 37503
rect 869 37469 903 37503
rect 903 37469 1005 37503
rect 1005 37469 1039 37503
rect 1039 37469 1141 37503
rect 1141 37469 1175 37503
rect 1175 37469 1277 37503
rect 1277 37469 1311 37503
rect 1311 37469 1413 37503
rect 1413 37469 1447 37503
rect 1447 37469 1549 37503
rect 1549 37469 1583 37503
rect 1583 37469 1685 37503
rect 1685 37469 1719 37503
rect 1719 37469 1723 37503
rect 321 37367 1723 37469
rect 321 37333 325 37367
rect 325 37333 359 37367
rect 359 37333 461 37367
rect 461 37333 495 37367
rect 495 37333 597 37367
rect 597 37333 631 37367
rect 631 37333 733 37367
rect 733 37333 767 37367
rect 767 37333 869 37367
rect 869 37333 903 37367
rect 903 37333 1005 37367
rect 1005 37333 1039 37367
rect 1039 37333 1141 37367
rect 1141 37333 1175 37367
rect 1175 37333 1277 37367
rect 1277 37333 1311 37367
rect 1311 37333 1413 37367
rect 1413 37333 1447 37367
rect 1447 37333 1549 37367
rect 1549 37333 1583 37367
rect 1583 37333 1685 37367
rect 1685 37333 1719 37367
rect 1719 37333 1723 37367
rect 321 37231 1723 37333
rect 321 37197 325 37231
rect 325 37197 359 37231
rect 359 37197 461 37231
rect 461 37197 495 37231
rect 495 37197 597 37231
rect 597 37197 631 37231
rect 631 37197 733 37231
rect 733 37197 767 37231
rect 767 37197 869 37231
rect 869 37197 903 37231
rect 903 37197 1005 37231
rect 1005 37197 1039 37231
rect 1039 37197 1141 37231
rect 1141 37197 1175 37231
rect 1175 37197 1277 37231
rect 1277 37197 1311 37231
rect 1311 37197 1413 37231
rect 1413 37197 1447 37231
rect 1447 37197 1549 37231
rect 1549 37197 1583 37231
rect 1583 37197 1685 37231
rect 1685 37197 1719 37231
rect 1719 37197 1723 37231
rect 321 37095 1723 37197
rect 321 37061 325 37095
rect 325 37061 359 37095
rect 359 37061 461 37095
rect 461 37061 495 37095
rect 495 37061 597 37095
rect 597 37061 631 37095
rect 631 37061 733 37095
rect 733 37061 767 37095
rect 767 37061 869 37095
rect 869 37061 903 37095
rect 903 37061 1005 37095
rect 1005 37061 1039 37095
rect 1039 37061 1141 37095
rect 1141 37061 1175 37095
rect 1175 37061 1277 37095
rect 1277 37061 1311 37095
rect 1311 37061 1413 37095
rect 1413 37061 1447 37095
rect 1447 37061 1549 37095
rect 1549 37061 1583 37095
rect 1583 37061 1685 37095
rect 1685 37061 1719 37095
rect 1719 37061 1723 37095
rect 321 36959 1723 37061
rect 321 36925 325 36959
rect 325 36925 359 36959
rect 359 36925 461 36959
rect 461 36925 495 36959
rect 495 36925 597 36959
rect 597 36925 631 36959
rect 631 36925 733 36959
rect 733 36925 767 36959
rect 767 36925 869 36959
rect 869 36925 903 36959
rect 903 36925 1005 36959
rect 1005 36925 1039 36959
rect 1039 36925 1141 36959
rect 1141 36925 1175 36959
rect 1175 36925 1277 36959
rect 1277 36925 1311 36959
rect 1311 36925 1413 36959
rect 1413 36925 1447 36959
rect 1447 36925 1549 36959
rect 1549 36925 1583 36959
rect 1583 36925 1685 36959
rect 1685 36925 1719 36959
rect 1719 36925 1723 36959
rect 321 36823 1723 36925
rect 321 36789 325 36823
rect 325 36789 359 36823
rect 359 36789 461 36823
rect 461 36789 495 36823
rect 495 36789 597 36823
rect 597 36789 631 36823
rect 631 36789 733 36823
rect 733 36789 767 36823
rect 767 36789 869 36823
rect 869 36789 903 36823
rect 903 36789 1005 36823
rect 1005 36789 1039 36823
rect 1039 36789 1141 36823
rect 1141 36789 1175 36823
rect 1175 36789 1277 36823
rect 1277 36789 1311 36823
rect 1311 36789 1413 36823
rect 1413 36789 1447 36823
rect 1447 36789 1549 36823
rect 1549 36789 1583 36823
rect 1583 36789 1685 36823
rect 1685 36789 1719 36823
rect 1719 36789 1723 36823
rect 321 36687 1723 36789
rect 321 36653 325 36687
rect 325 36653 359 36687
rect 359 36653 461 36687
rect 461 36653 495 36687
rect 495 36653 597 36687
rect 597 36653 631 36687
rect 631 36653 733 36687
rect 733 36653 767 36687
rect 767 36653 869 36687
rect 869 36653 903 36687
rect 903 36653 1005 36687
rect 1005 36653 1039 36687
rect 1039 36653 1141 36687
rect 1141 36653 1175 36687
rect 1175 36653 1277 36687
rect 1277 36653 1311 36687
rect 1311 36653 1413 36687
rect 1413 36653 1447 36687
rect 1447 36653 1549 36687
rect 1549 36653 1583 36687
rect 1583 36653 1685 36687
rect 1685 36653 1719 36687
rect 1719 36653 1723 36687
rect 321 36551 1723 36653
rect 321 36517 325 36551
rect 325 36517 359 36551
rect 359 36517 461 36551
rect 461 36517 495 36551
rect 495 36517 597 36551
rect 597 36517 631 36551
rect 631 36517 733 36551
rect 733 36517 767 36551
rect 767 36517 869 36551
rect 869 36517 903 36551
rect 903 36517 1005 36551
rect 1005 36517 1039 36551
rect 1039 36517 1141 36551
rect 1141 36517 1175 36551
rect 1175 36517 1277 36551
rect 1277 36517 1311 36551
rect 1311 36517 1413 36551
rect 1413 36517 1447 36551
rect 1447 36517 1549 36551
rect 1549 36517 1583 36551
rect 1583 36517 1685 36551
rect 1685 36517 1719 36551
rect 1719 36517 1723 36551
rect 321 36415 1723 36517
rect 321 36381 325 36415
rect 325 36381 359 36415
rect 359 36381 461 36415
rect 461 36381 495 36415
rect 495 36381 597 36415
rect 597 36381 631 36415
rect 631 36381 733 36415
rect 733 36381 767 36415
rect 767 36381 869 36415
rect 869 36381 903 36415
rect 903 36381 1005 36415
rect 1005 36381 1039 36415
rect 1039 36381 1141 36415
rect 1141 36381 1175 36415
rect 1175 36381 1277 36415
rect 1277 36381 1311 36415
rect 1311 36381 1413 36415
rect 1413 36381 1447 36415
rect 1447 36381 1549 36415
rect 1549 36381 1583 36415
rect 1583 36381 1685 36415
rect 1685 36381 1719 36415
rect 1719 36381 1723 36415
rect 321 36279 1723 36381
rect 321 36245 325 36279
rect 325 36245 359 36279
rect 359 36245 461 36279
rect 461 36245 495 36279
rect 495 36245 597 36279
rect 597 36245 631 36279
rect 631 36245 733 36279
rect 733 36245 767 36279
rect 767 36245 869 36279
rect 869 36245 903 36279
rect 903 36245 1005 36279
rect 1005 36245 1039 36279
rect 1039 36245 1141 36279
rect 1141 36245 1175 36279
rect 1175 36245 1277 36279
rect 1277 36245 1311 36279
rect 1311 36245 1413 36279
rect 1413 36245 1447 36279
rect 1447 36245 1549 36279
rect 1549 36245 1583 36279
rect 1583 36245 1685 36279
rect 1685 36245 1719 36279
rect 1719 36245 1723 36279
rect 321 36143 1723 36245
rect 321 36109 325 36143
rect 325 36109 359 36143
rect 359 36109 461 36143
rect 461 36109 495 36143
rect 495 36109 597 36143
rect 597 36109 631 36143
rect 631 36109 733 36143
rect 733 36109 767 36143
rect 767 36109 869 36143
rect 869 36109 903 36143
rect 903 36109 1005 36143
rect 1005 36109 1039 36143
rect 1039 36109 1141 36143
rect 1141 36109 1175 36143
rect 1175 36109 1277 36143
rect 1277 36109 1311 36143
rect 1311 36109 1413 36143
rect 1413 36109 1447 36143
rect 1447 36109 1549 36143
rect 1549 36109 1583 36143
rect 1583 36109 1685 36143
rect 1685 36109 1719 36143
rect 1719 36109 1723 36143
rect 321 36007 1723 36109
rect 321 35973 325 36007
rect 325 35973 359 36007
rect 359 35973 461 36007
rect 461 35973 495 36007
rect 495 35973 597 36007
rect 597 35973 631 36007
rect 631 35973 733 36007
rect 733 35973 767 36007
rect 767 35973 869 36007
rect 869 35973 903 36007
rect 903 35973 1005 36007
rect 1005 35973 1039 36007
rect 1039 35973 1141 36007
rect 1141 35973 1175 36007
rect 1175 35973 1277 36007
rect 1277 35973 1311 36007
rect 1311 35973 1413 36007
rect 1413 35973 1447 36007
rect 1447 35973 1549 36007
rect 1549 35973 1583 36007
rect 1583 35973 1685 36007
rect 1685 35973 1719 36007
rect 1719 35973 1723 36007
rect 321 35871 1723 35973
rect 321 35837 325 35871
rect 325 35837 359 35871
rect 359 35837 461 35871
rect 461 35837 495 35871
rect 495 35837 597 35871
rect 597 35837 631 35871
rect 631 35837 733 35871
rect 733 35837 767 35871
rect 767 35837 869 35871
rect 869 35837 903 35871
rect 903 35837 1005 35871
rect 1005 35837 1039 35871
rect 1039 35837 1141 35871
rect 1141 35837 1175 35871
rect 1175 35837 1277 35871
rect 1277 35837 1311 35871
rect 1311 35837 1413 35871
rect 1413 35837 1447 35871
rect 1447 35837 1549 35871
rect 1549 35837 1583 35871
rect 1583 35837 1685 35871
rect 1685 35837 1719 35871
rect 1719 35837 1723 35871
rect 321 35735 1723 35837
rect 321 35701 325 35735
rect 325 35701 359 35735
rect 359 35701 461 35735
rect 461 35701 495 35735
rect 495 35701 597 35735
rect 597 35701 631 35735
rect 631 35701 733 35735
rect 733 35701 767 35735
rect 767 35701 869 35735
rect 869 35701 903 35735
rect 903 35701 1005 35735
rect 1005 35701 1039 35735
rect 1039 35701 1141 35735
rect 1141 35701 1175 35735
rect 1175 35701 1277 35735
rect 1277 35701 1311 35735
rect 1311 35701 1413 35735
rect 1413 35701 1447 35735
rect 1447 35701 1549 35735
rect 1549 35701 1583 35735
rect 1583 35701 1685 35735
rect 1685 35701 1719 35735
rect 1719 35701 1723 35735
rect 321 35599 1723 35701
rect 321 35565 325 35599
rect 325 35565 359 35599
rect 359 35565 461 35599
rect 461 35565 495 35599
rect 495 35565 597 35599
rect 597 35565 631 35599
rect 631 35565 733 35599
rect 733 35565 767 35599
rect 767 35565 869 35599
rect 869 35565 903 35599
rect 903 35565 1005 35599
rect 1005 35565 1039 35599
rect 1039 35565 1141 35599
rect 1141 35565 1175 35599
rect 1175 35565 1277 35599
rect 1277 35565 1311 35599
rect 1311 35565 1413 35599
rect 1413 35565 1447 35599
rect 1447 35565 1549 35599
rect 1549 35565 1583 35599
rect 1583 35565 1685 35599
rect 1685 35565 1719 35599
rect 1719 35565 1723 35599
rect 321 35463 1723 35565
rect 321 35429 325 35463
rect 325 35429 359 35463
rect 359 35429 461 35463
rect 461 35429 495 35463
rect 495 35429 597 35463
rect 597 35429 631 35463
rect 631 35429 733 35463
rect 733 35429 767 35463
rect 767 35429 869 35463
rect 869 35429 903 35463
rect 903 35429 1005 35463
rect 1005 35429 1039 35463
rect 1039 35429 1141 35463
rect 1141 35429 1175 35463
rect 1175 35429 1277 35463
rect 1277 35429 1311 35463
rect 1311 35429 1413 35463
rect 1413 35429 1447 35463
rect 1447 35429 1549 35463
rect 1549 35429 1583 35463
rect 1583 35429 1685 35463
rect 1685 35429 1719 35463
rect 1719 35429 1723 35463
rect 321 35327 1723 35429
rect 321 35293 325 35327
rect 325 35293 359 35327
rect 359 35293 461 35327
rect 461 35293 495 35327
rect 495 35293 597 35327
rect 597 35293 631 35327
rect 631 35293 733 35327
rect 733 35293 767 35327
rect 767 35293 869 35327
rect 869 35293 903 35327
rect 903 35293 1005 35327
rect 1005 35293 1039 35327
rect 1039 35293 1141 35327
rect 1141 35293 1175 35327
rect 1175 35293 1277 35327
rect 1277 35293 1311 35327
rect 1311 35293 1413 35327
rect 1413 35293 1447 35327
rect 1447 35293 1549 35327
rect 1549 35293 1583 35327
rect 1583 35293 1685 35327
rect 1685 35293 1719 35327
rect 1719 35293 1723 35327
rect 321 35191 1723 35293
rect 321 35157 325 35191
rect 325 35157 359 35191
rect 359 35157 461 35191
rect 461 35157 495 35191
rect 495 35157 597 35191
rect 597 35157 631 35191
rect 631 35157 733 35191
rect 733 35157 767 35191
rect 767 35157 869 35191
rect 869 35157 903 35191
rect 903 35157 1005 35191
rect 1005 35157 1039 35191
rect 1039 35157 1141 35191
rect 1141 35157 1175 35191
rect 1175 35157 1277 35191
rect 1277 35157 1311 35191
rect 1311 35157 1413 35191
rect 1413 35157 1447 35191
rect 1447 35157 1549 35191
rect 1549 35157 1583 35191
rect 1583 35157 1685 35191
rect 1685 35157 1719 35191
rect 1719 35157 1723 35191
rect 321 35055 1723 35157
rect 321 35021 325 35055
rect 325 35021 359 35055
rect 359 35021 461 35055
rect 461 35021 495 35055
rect 495 35021 597 35055
rect 597 35021 631 35055
rect 631 35021 733 35055
rect 733 35021 767 35055
rect 767 35021 869 35055
rect 869 35021 903 35055
rect 903 35021 1005 35055
rect 1005 35021 1039 35055
rect 1039 35021 1141 35055
rect 1141 35021 1175 35055
rect 1175 35021 1277 35055
rect 1277 35021 1311 35055
rect 1311 35021 1413 35055
rect 1413 35021 1447 35055
rect 1447 35021 1549 35055
rect 1549 35021 1583 35055
rect 1583 35021 1685 35055
rect 1685 35021 1719 35055
rect 1719 35021 1723 35055
rect 321 34919 1723 35021
rect 321 34885 325 34919
rect 325 34885 359 34919
rect 359 34885 461 34919
rect 461 34885 495 34919
rect 495 34885 597 34919
rect 597 34885 631 34919
rect 631 34885 733 34919
rect 733 34885 767 34919
rect 767 34885 869 34919
rect 869 34885 903 34919
rect 903 34885 1005 34919
rect 1005 34885 1039 34919
rect 1039 34885 1141 34919
rect 1141 34885 1175 34919
rect 1175 34885 1277 34919
rect 1277 34885 1311 34919
rect 1311 34885 1413 34919
rect 1413 34885 1447 34919
rect 1447 34885 1549 34919
rect 1549 34885 1583 34919
rect 1583 34885 1685 34919
rect 1685 34885 1719 34919
rect 1719 34885 1723 34919
rect 321 34783 1723 34885
rect 321 34749 325 34783
rect 325 34749 359 34783
rect 359 34749 461 34783
rect 461 34749 495 34783
rect 495 34749 597 34783
rect 597 34749 631 34783
rect 631 34749 733 34783
rect 733 34749 767 34783
rect 767 34749 869 34783
rect 869 34749 903 34783
rect 903 34749 1005 34783
rect 1005 34749 1039 34783
rect 1039 34749 1141 34783
rect 1141 34749 1175 34783
rect 1175 34749 1277 34783
rect 1277 34749 1311 34783
rect 1311 34749 1413 34783
rect 1413 34749 1447 34783
rect 1447 34749 1549 34783
rect 1549 34749 1583 34783
rect 1583 34749 1685 34783
rect 1685 34749 1719 34783
rect 1719 34749 1723 34783
rect 321 34647 1723 34749
rect 321 34613 325 34647
rect 325 34613 359 34647
rect 359 34613 461 34647
rect 461 34613 495 34647
rect 495 34613 597 34647
rect 597 34613 631 34647
rect 631 34613 733 34647
rect 733 34613 767 34647
rect 767 34613 869 34647
rect 869 34613 903 34647
rect 903 34613 1005 34647
rect 1005 34613 1039 34647
rect 1039 34613 1141 34647
rect 1141 34613 1175 34647
rect 1175 34613 1277 34647
rect 1277 34613 1311 34647
rect 1311 34613 1413 34647
rect 1413 34613 1447 34647
rect 1447 34613 1549 34647
rect 1549 34613 1583 34647
rect 1583 34613 1685 34647
rect 1685 34613 1719 34647
rect 1719 34613 1723 34647
rect 321 34511 1723 34613
rect 321 34477 325 34511
rect 325 34477 359 34511
rect 359 34477 461 34511
rect 461 34477 495 34511
rect 495 34477 597 34511
rect 597 34477 631 34511
rect 631 34477 733 34511
rect 733 34477 767 34511
rect 767 34477 869 34511
rect 869 34477 903 34511
rect 903 34477 1005 34511
rect 1005 34477 1039 34511
rect 1039 34477 1141 34511
rect 1141 34477 1175 34511
rect 1175 34477 1277 34511
rect 1277 34477 1311 34511
rect 1311 34477 1413 34511
rect 1413 34477 1447 34511
rect 1447 34477 1549 34511
rect 1549 34477 1583 34511
rect 1583 34477 1685 34511
rect 1685 34477 1719 34511
rect 1719 34477 1723 34511
rect 321 34375 1723 34477
rect 321 34341 325 34375
rect 325 34341 359 34375
rect 359 34341 461 34375
rect 461 34341 495 34375
rect 495 34341 597 34375
rect 597 34341 631 34375
rect 631 34341 733 34375
rect 733 34341 767 34375
rect 767 34341 869 34375
rect 869 34341 903 34375
rect 903 34341 1005 34375
rect 1005 34341 1039 34375
rect 1039 34341 1141 34375
rect 1141 34341 1175 34375
rect 1175 34341 1277 34375
rect 1277 34341 1311 34375
rect 1311 34341 1413 34375
rect 1413 34341 1447 34375
rect 1447 34341 1549 34375
rect 1549 34341 1583 34375
rect 1583 34341 1685 34375
rect 1685 34341 1719 34375
rect 1719 34341 1723 34375
rect 321 34239 1723 34341
rect 321 34205 325 34239
rect 325 34205 359 34239
rect 359 34205 461 34239
rect 461 34205 495 34239
rect 495 34205 597 34239
rect 597 34205 631 34239
rect 631 34205 733 34239
rect 733 34205 767 34239
rect 767 34205 869 34239
rect 869 34205 903 34239
rect 903 34205 1005 34239
rect 1005 34205 1039 34239
rect 1039 34205 1141 34239
rect 1141 34205 1175 34239
rect 1175 34205 1277 34239
rect 1277 34205 1311 34239
rect 1311 34205 1413 34239
rect 1413 34205 1447 34239
rect 1447 34205 1549 34239
rect 1549 34205 1583 34239
rect 1583 34205 1685 34239
rect 1685 34205 1719 34239
rect 1719 34205 1723 34239
rect 321 34103 1723 34205
rect 321 34069 325 34103
rect 325 34069 359 34103
rect 359 34069 461 34103
rect 461 34069 495 34103
rect 495 34069 597 34103
rect 597 34069 631 34103
rect 631 34069 733 34103
rect 733 34069 767 34103
rect 767 34069 869 34103
rect 869 34069 903 34103
rect 903 34069 1005 34103
rect 1005 34069 1039 34103
rect 1039 34069 1141 34103
rect 1141 34069 1175 34103
rect 1175 34069 1277 34103
rect 1277 34069 1311 34103
rect 1311 34069 1413 34103
rect 1413 34069 1447 34103
rect 1447 34069 1549 34103
rect 1549 34069 1583 34103
rect 1583 34069 1685 34103
rect 1685 34069 1719 34103
rect 1719 34069 1723 34103
rect 321 33967 1723 34069
rect 321 33933 325 33967
rect 325 33933 359 33967
rect 359 33933 461 33967
rect 461 33933 495 33967
rect 495 33933 597 33967
rect 597 33933 631 33967
rect 631 33933 733 33967
rect 733 33933 767 33967
rect 767 33933 869 33967
rect 869 33933 903 33967
rect 903 33933 1005 33967
rect 1005 33933 1039 33967
rect 1039 33933 1141 33967
rect 1141 33933 1175 33967
rect 1175 33933 1277 33967
rect 1277 33933 1311 33967
rect 1311 33933 1413 33967
rect 1413 33933 1447 33967
rect 1447 33933 1549 33967
rect 1549 33933 1583 33967
rect 1583 33933 1685 33967
rect 1685 33933 1719 33967
rect 1719 33933 1723 33967
rect 321 33831 1723 33933
rect 321 33797 325 33831
rect 325 33797 359 33831
rect 359 33797 461 33831
rect 461 33797 495 33831
rect 495 33797 597 33831
rect 597 33797 631 33831
rect 631 33797 733 33831
rect 733 33797 767 33831
rect 767 33797 869 33831
rect 869 33797 903 33831
rect 903 33797 1005 33831
rect 1005 33797 1039 33831
rect 1039 33797 1141 33831
rect 1141 33797 1175 33831
rect 1175 33797 1277 33831
rect 1277 33797 1311 33831
rect 1311 33797 1413 33831
rect 1413 33797 1447 33831
rect 1447 33797 1549 33831
rect 1549 33797 1583 33831
rect 1583 33797 1685 33831
rect 1685 33797 1719 33831
rect 1719 33797 1723 33831
rect 321 33695 1723 33797
rect 321 33661 325 33695
rect 325 33661 359 33695
rect 359 33661 461 33695
rect 461 33661 495 33695
rect 495 33661 597 33695
rect 597 33661 631 33695
rect 631 33661 733 33695
rect 733 33661 767 33695
rect 767 33661 869 33695
rect 869 33661 903 33695
rect 903 33661 1005 33695
rect 1005 33661 1039 33695
rect 1039 33661 1141 33695
rect 1141 33661 1175 33695
rect 1175 33661 1277 33695
rect 1277 33661 1311 33695
rect 1311 33661 1413 33695
rect 1413 33661 1447 33695
rect 1447 33661 1549 33695
rect 1549 33661 1583 33695
rect 1583 33661 1685 33695
rect 1685 33661 1719 33695
rect 1719 33661 1723 33695
rect 321 33559 1723 33661
rect 321 33525 325 33559
rect 325 33525 359 33559
rect 359 33525 461 33559
rect 461 33525 495 33559
rect 495 33525 597 33559
rect 597 33525 631 33559
rect 631 33525 733 33559
rect 733 33525 767 33559
rect 767 33525 869 33559
rect 869 33525 903 33559
rect 903 33525 1005 33559
rect 1005 33525 1039 33559
rect 1039 33525 1141 33559
rect 1141 33525 1175 33559
rect 1175 33525 1277 33559
rect 1277 33525 1311 33559
rect 1311 33525 1413 33559
rect 1413 33525 1447 33559
rect 1447 33525 1549 33559
rect 1549 33525 1583 33559
rect 1583 33525 1685 33559
rect 1685 33525 1719 33559
rect 1719 33525 1723 33559
rect 321 33423 1723 33525
rect 321 33389 325 33423
rect 325 33389 359 33423
rect 359 33389 461 33423
rect 461 33389 495 33423
rect 495 33389 597 33423
rect 597 33389 631 33423
rect 631 33389 733 33423
rect 733 33389 767 33423
rect 767 33389 869 33423
rect 869 33389 903 33423
rect 903 33389 1005 33423
rect 1005 33389 1039 33423
rect 1039 33389 1141 33423
rect 1141 33389 1175 33423
rect 1175 33389 1277 33423
rect 1277 33389 1311 33423
rect 1311 33389 1413 33423
rect 1413 33389 1447 33423
rect 1447 33389 1549 33423
rect 1549 33389 1583 33423
rect 1583 33389 1685 33423
rect 1685 33389 1719 33423
rect 1719 33389 1723 33423
rect 321 33357 1723 33389
rect 321 33287 355 33318
rect 321 33284 325 33287
rect 325 33284 355 33287
rect 393 33284 427 33318
rect 465 33287 499 33318
rect 465 33284 495 33287
rect 495 33284 499 33287
rect 537 33284 571 33318
rect 609 33287 643 33318
rect 609 33284 631 33287
rect 631 33284 643 33287
rect 681 33284 715 33318
rect 753 33287 787 33318
rect 753 33284 767 33287
rect 767 33284 787 33287
rect 825 33284 859 33318
rect 897 33287 931 33318
rect 897 33284 903 33287
rect 903 33284 931 33287
rect 969 33284 1003 33318
rect 1041 33284 1075 33318
rect 1113 33287 1147 33318
rect 1113 33284 1141 33287
rect 1141 33284 1147 33287
rect 1185 33284 1219 33318
rect 1257 33287 1291 33318
rect 1257 33284 1277 33287
rect 1277 33284 1291 33287
rect 1329 33284 1363 33318
rect 1401 33287 1435 33318
rect 1401 33284 1413 33287
rect 1413 33284 1435 33287
rect 1473 33284 1507 33318
rect 1545 33287 1579 33318
rect 1545 33284 1549 33287
rect 1549 33284 1579 33287
rect 1617 33284 1651 33318
rect 1689 33287 1723 33318
rect 1689 33284 1719 33287
rect 1719 33284 1723 33287
rect 321 33211 355 33245
rect 393 33211 427 33245
rect 465 33211 499 33245
rect 537 33211 571 33245
rect 609 33211 643 33245
rect 681 33211 715 33245
rect 753 33211 787 33245
rect 825 33211 859 33245
rect 897 33211 931 33245
rect 969 33211 1003 33245
rect 1041 33211 1075 33245
rect 1113 33211 1147 33245
rect 1185 33211 1219 33245
rect 1257 33211 1291 33245
rect 1329 33211 1363 33245
rect 1401 33211 1435 33245
rect 1473 33211 1507 33245
rect 1545 33211 1579 33245
rect 1617 33211 1651 33245
rect 1689 33211 1723 33245
rect 321 33151 355 33172
rect 321 33138 325 33151
rect 325 33138 355 33151
rect 393 33138 427 33172
rect 465 33151 499 33172
rect 465 33138 495 33151
rect 495 33138 499 33151
rect 537 33138 571 33172
rect 609 33151 643 33172
rect 609 33138 631 33151
rect 631 33138 643 33151
rect 681 33138 715 33172
rect 753 33151 787 33172
rect 753 33138 767 33151
rect 767 33138 787 33151
rect 825 33138 859 33172
rect 897 33151 931 33172
rect 897 33138 903 33151
rect 903 33138 931 33151
rect 969 33138 1003 33172
rect 1041 33138 1075 33172
rect 1113 33151 1147 33172
rect 1113 33138 1141 33151
rect 1141 33138 1147 33151
rect 1185 33138 1219 33172
rect 1257 33151 1291 33172
rect 1257 33138 1277 33151
rect 1277 33138 1291 33151
rect 1329 33138 1363 33172
rect 1401 33151 1435 33172
rect 1401 33138 1413 33151
rect 1413 33138 1435 33151
rect 1473 33138 1507 33172
rect 1545 33151 1579 33172
rect 1545 33138 1549 33151
rect 1549 33138 1579 33151
rect 1617 33138 1651 33172
rect 1689 33151 1723 33172
rect 1689 33138 1719 33151
rect 1719 33138 1723 33151
rect 321 33065 355 33099
rect 393 33065 427 33099
rect 465 33065 499 33099
rect 537 33065 571 33099
rect 609 33065 643 33099
rect 681 33065 715 33099
rect 753 33065 787 33099
rect 825 33065 859 33099
rect 897 33065 931 33099
rect 969 33065 1003 33099
rect 1041 33065 1075 33099
rect 1113 33065 1147 33099
rect 1185 33065 1219 33099
rect 1257 33065 1291 33099
rect 1329 33065 1363 33099
rect 1401 33065 1435 33099
rect 1473 33065 1507 33099
rect 1545 33065 1579 33099
rect 1617 33065 1651 33099
rect 1689 33065 1723 33099
rect 321 33015 355 33026
rect 321 32992 325 33015
rect 325 32992 355 33015
rect 393 32992 427 33026
rect 465 33015 499 33026
rect 465 32992 495 33015
rect 495 32992 499 33015
rect 537 32992 571 33026
rect 609 33015 643 33026
rect 609 32992 631 33015
rect 631 32992 643 33015
rect 681 32992 715 33026
rect 753 33015 787 33026
rect 753 32992 767 33015
rect 767 32992 787 33015
rect 825 32992 859 33026
rect 897 33015 931 33026
rect 897 32992 903 33015
rect 903 32992 931 33015
rect 969 32992 1003 33026
rect 1041 32992 1075 33026
rect 1113 33015 1147 33026
rect 1113 32992 1141 33015
rect 1141 32992 1147 33015
rect 1185 32992 1219 33026
rect 1257 33015 1291 33026
rect 1257 32992 1277 33015
rect 1277 32992 1291 33015
rect 1329 32992 1363 33026
rect 1401 33015 1435 33026
rect 1401 32992 1413 33015
rect 1413 32992 1435 33015
rect 1473 32992 1507 33026
rect 1545 33015 1579 33026
rect 1545 32992 1549 33015
rect 1549 32992 1579 33015
rect 1617 32992 1651 33026
rect 1689 33015 1723 33026
rect 1689 32992 1719 33015
rect 1719 32992 1723 33015
rect 321 32919 355 32953
rect 393 32919 427 32953
rect 465 32919 499 32953
rect 537 32919 571 32953
rect 609 32919 643 32953
rect 681 32919 715 32953
rect 753 32919 787 32953
rect 825 32919 859 32953
rect 897 32919 931 32953
rect 969 32919 1003 32953
rect 1041 32919 1075 32953
rect 1113 32919 1147 32953
rect 1185 32919 1219 32953
rect 1257 32919 1291 32953
rect 1329 32919 1363 32953
rect 1401 32919 1435 32953
rect 1473 32919 1507 32953
rect 1545 32919 1579 32953
rect 1617 32919 1651 32953
rect 1689 32919 1723 32953
rect 321 32879 355 32880
rect 321 32846 325 32879
rect 325 32846 355 32879
rect 393 32846 427 32880
rect 465 32879 499 32880
rect 465 32846 495 32879
rect 495 32846 499 32879
rect 537 32846 571 32880
rect 609 32879 643 32880
rect 609 32846 631 32879
rect 631 32846 643 32879
rect 681 32846 715 32880
rect 753 32879 787 32880
rect 753 32846 767 32879
rect 767 32846 787 32879
rect 825 32846 859 32880
rect 897 32879 931 32880
rect 897 32846 903 32879
rect 903 32846 931 32879
rect 969 32846 1003 32880
rect 1041 32846 1075 32880
rect 1113 32879 1147 32880
rect 1113 32846 1141 32879
rect 1141 32846 1147 32879
rect 1185 32846 1219 32880
rect 1257 32879 1291 32880
rect 1257 32846 1277 32879
rect 1277 32846 1291 32879
rect 1329 32846 1363 32880
rect 1401 32879 1435 32880
rect 1401 32846 1413 32879
rect 1413 32846 1435 32879
rect 1473 32846 1507 32880
rect 1545 32879 1579 32880
rect 1545 32846 1549 32879
rect 1549 32846 1579 32879
rect 1617 32846 1651 32880
rect 1689 32879 1723 32880
rect 1689 32846 1719 32879
rect 1719 32846 1723 32879
rect 321 32773 355 32807
rect 393 32773 427 32807
rect 465 32773 499 32807
rect 537 32773 571 32807
rect 609 32773 643 32807
rect 681 32773 715 32807
rect 753 32773 787 32807
rect 825 32773 859 32807
rect 897 32773 931 32807
rect 969 32773 1003 32807
rect 1041 32773 1075 32807
rect 1113 32773 1147 32807
rect 1185 32773 1219 32807
rect 1257 32773 1291 32807
rect 1329 32773 1363 32807
rect 1401 32773 1435 32807
rect 1473 32773 1507 32807
rect 1545 32773 1579 32807
rect 1617 32773 1651 32807
rect 1689 32773 1723 32807
rect 321 32709 325 32734
rect 325 32709 355 32734
rect 321 32700 355 32709
rect 393 32700 427 32734
rect 465 32709 495 32734
rect 495 32709 499 32734
rect 465 32700 499 32709
rect 537 32700 571 32734
rect 609 32709 631 32734
rect 631 32709 643 32734
rect 609 32700 643 32709
rect 681 32700 715 32734
rect 753 32709 767 32734
rect 767 32709 787 32734
rect 753 32700 787 32709
rect 825 32700 859 32734
rect 897 32709 903 32734
rect 903 32709 931 32734
rect 897 32700 931 32709
rect 969 32700 1003 32734
rect 1041 32700 1075 32734
rect 1113 32709 1141 32734
rect 1141 32709 1147 32734
rect 1113 32700 1147 32709
rect 1185 32700 1219 32734
rect 1257 32709 1277 32734
rect 1277 32709 1291 32734
rect 1257 32700 1291 32709
rect 1329 32700 1363 32734
rect 1401 32709 1413 32734
rect 1413 32709 1435 32734
rect 1401 32700 1435 32709
rect 1473 32700 1507 32734
rect 1545 32709 1549 32734
rect 1549 32709 1579 32734
rect 1545 32700 1579 32709
rect 1617 32700 1651 32734
rect 1689 32709 1719 32734
rect 1719 32709 1723 32734
rect 1689 32700 1723 32709
rect 321 32627 355 32661
rect 393 32627 427 32661
rect 465 32627 499 32661
rect 537 32627 571 32661
rect 609 32627 643 32661
rect 681 32627 715 32661
rect 753 32627 787 32661
rect 825 32627 859 32661
rect 897 32627 931 32661
rect 969 32627 1003 32661
rect 1041 32627 1075 32661
rect 1113 32627 1147 32661
rect 1185 32627 1219 32661
rect 1257 32627 1291 32661
rect 1329 32627 1363 32661
rect 1401 32627 1435 32661
rect 1473 32627 1507 32661
rect 1545 32627 1579 32661
rect 1617 32627 1651 32661
rect 1689 32627 1723 32661
rect 321 32573 325 32588
rect 325 32573 355 32588
rect 321 32554 355 32573
rect 393 32554 427 32588
rect 465 32573 495 32588
rect 495 32573 499 32588
rect 465 32554 499 32573
rect 537 32554 571 32588
rect 609 32573 631 32588
rect 631 32573 643 32588
rect 609 32554 643 32573
rect 681 32554 715 32588
rect 753 32573 767 32588
rect 767 32573 787 32588
rect 753 32554 787 32573
rect 825 32554 859 32588
rect 897 32573 903 32588
rect 903 32573 931 32588
rect 897 32554 931 32573
rect 969 32554 1003 32588
rect 1041 32554 1075 32588
rect 1113 32573 1141 32588
rect 1141 32573 1147 32588
rect 1113 32554 1147 32573
rect 1185 32554 1219 32588
rect 1257 32573 1277 32588
rect 1277 32573 1291 32588
rect 1257 32554 1291 32573
rect 1329 32554 1363 32588
rect 1401 32573 1413 32588
rect 1413 32573 1435 32588
rect 1401 32554 1435 32573
rect 1473 32554 1507 32588
rect 1545 32573 1549 32588
rect 1549 32573 1579 32588
rect 1545 32554 1579 32573
rect 1617 32554 1651 32588
rect 1689 32573 1719 32588
rect 1719 32573 1723 32588
rect 1689 32554 1723 32573
rect 321 32481 355 32515
rect 393 32481 427 32515
rect 465 32481 499 32515
rect 537 32481 571 32515
rect 609 32481 643 32515
rect 681 32481 715 32515
rect 753 32481 787 32515
rect 825 32481 859 32515
rect 897 32481 931 32515
rect 969 32481 1003 32515
rect 1041 32481 1075 32515
rect 1113 32481 1147 32515
rect 1185 32481 1219 32515
rect 1257 32481 1291 32515
rect 1329 32481 1363 32515
rect 1401 32481 1435 32515
rect 1473 32481 1507 32515
rect 1545 32481 1579 32515
rect 1617 32481 1651 32515
rect 1689 32481 1723 32515
rect 321 32437 325 32442
rect 325 32437 355 32442
rect 321 32408 355 32437
rect 393 32408 427 32442
rect 465 32437 495 32442
rect 495 32437 499 32442
rect 465 32408 499 32437
rect 537 32408 571 32442
rect 609 32437 631 32442
rect 631 32437 643 32442
rect 609 32408 643 32437
rect 681 32408 715 32442
rect 753 32437 767 32442
rect 767 32437 787 32442
rect 753 32408 787 32437
rect 825 32408 859 32442
rect 897 32437 903 32442
rect 903 32437 931 32442
rect 897 32408 931 32437
rect 969 32408 1003 32442
rect 1041 32408 1075 32442
rect 1113 32437 1141 32442
rect 1141 32437 1147 32442
rect 1113 32408 1147 32437
rect 1185 32408 1219 32442
rect 1257 32437 1277 32442
rect 1277 32437 1291 32442
rect 1257 32408 1291 32437
rect 1329 32408 1363 32442
rect 1401 32437 1413 32442
rect 1413 32437 1435 32442
rect 1401 32408 1435 32437
rect 1473 32408 1507 32442
rect 1545 32437 1549 32442
rect 1549 32437 1579 32442
rect 1545 32408 1579 32437
rect 1617 32408 1651 32442
rect 1689 32437 1719 32442
rect 1719 32437 1723 32442
rect 1689 32408 1723 32437
rect 321 32335 355 32369
rect 393 32335 427 32369
rect 465 32335 499 32369
rect 537 32335 571 32369
rect 609 32335 643 32369
rect 681 32335 715 32369
rect 753 32335 787 32369
rect 825 32335 859 32369
rect 897 32335 931 32369
rect 969 32335 1003 32369
rect 1041 32335 1075 32369
rect 1113 32335 1147 32369
rect 1185 32335 1219 32369
rect 1257 32335 1291 32369
rect 1329 32335 1363 32369
rect 1401 32335 1435 32369
rect 1473 32335 1507 32369
rect 1545 32335 1579 32369
rect 1617 32335 1651 32369
rect 1689 32335 1723 32369
rect 321 32262 355 32296
rect 393 32262 427 32296
rect 465 32262 499 32296
rect 537 32262 571 32296
rect 609 32262 643 32296
rect 681 32262 715 32296
rect 753 32262 787 32296
rect 825 32262 859 32296
rect 897 32262 931 32296
rect 969 32262 1003 32296
rect 1041 32262 1075 32296
rect 1113 32262 1147 32296
rect 1185 32262 1219 32296
rect 1257 32262 1291 32296
rect 1329 32262 1363 32296
rect 1401 32262 1435 32296
rect 1473 32262 1507 32296
rect 1545 32262 1579 32296
rect 1617 32262 1651 32296
rect 1689 32262 1723 32296
rect 321 32199 355 32223
rect 321 32189 325 32199
rect 325 32189 355 32199
rect 393 32189 427 32223
rect 465 32199 499 32223
rect 465 32189 495 32199
rect 495 32189 499 32199
rect 537 32189 571 32223
rect 609 32199 643 32223
rect 609 32189 631 32199
rect 631 32189 643 32199
rect 681 32189 715 32223
rect 753 32199 787 32223
rect 753 32189 767 32199
rect 767 32189 787 32199
rect 825 32189 859 32223
rect 897 32199 931 32223
rect 897 32189 903 32199
rect 903 32189 931 32199
rect 969 32189 1003 32223
rect 1041 32189 1075 32223
rect 1113 32199 1147 32223
rect 1113 32189 1141 32199
rect 1141 32189 1147 32199
rect 1185 32189 1219 32223
rect 1257 32199 1291 32223
rect 1257 32189 1277 32199
rect 1277 32189 1291 32199
rect 1329 32189 1363 32223
rect 1401 32199 1435 32223
rect 1401 32189 1413 32199
rect 1413 32189 1435 32199
rect 1473 32189 1507 32223
rect 1545 32199 1579 32223
rect 1545 32189 1549 32199
rect 1549 32189 1579 32199
rect 1617 32189 1651 32223
rect 1689 32199 1723 32223
rect 1689 32189 1719 32199
rect 1719 32189 1723 32199
rect 321 32116 355 32150
rect 393 32116 427 32150
rect 465 32116 499 32150
rect 537 32116 571 32150
rect 609 32116 643 32150
rect 681 32116 715 32150
rect 753 32116 787 32150
rect 825 32116 859 32150
rect 897 32116 931 32150
rect 969 32116 1003 32150
rect 1041 32116 1075 32150
rect 1113 32116 1147 32150
rect 1185 32116 1219 32150
rect 1257 32116 1291 32150
rect 1329 32116 1363 32150
rect 1401 32116 1435 32150
rect 1473 32116 1507 32150
rect 1545 32116 1579 32150
rect 1617 32116 1651 32150
rect 1689 32116 1723 32150
rect 321 32063 355 32077
rect 321 32043 325 32063
rect 325 32043 355 32063
rect 393 32043 427 32077
rect 465 32063 499 32077
rect 465 32043 495 32063
rect 495 32043 499 32063
rect 537 32043 571 32077
rect 609 32063 643 32077
rect 609 32043 631 32063
rect 631 32043 643 32063
rect 681 32043 715 32077
rect 753 32063 787 32077
rect 753 32043 767 32063
rect 767 32043 787 32063
rect 825 32043 859 32077
rect 897 32063 931 32077
rect 897 32043 903 32063
rect 903 32043 931 32063
rect 969 32043 1003 32077
rect 1041 32043 1075 32077
rect 1113 32063 1147 32077
rect 1113 32043 1141 32063
rect 1141 32043 1147 32063
rect 1185 32043 1219 32077
rect 1257 32063 1291 32077
rect 1257 32043 1277 32063
rect 1277 32043 1291 32063
rect 1329 32043 1363 32077
rect 1401 32063 1435 32077
rect 1401 32043 1413 32063
rect 1413 32043 1435 32063
rect 1473 32043 1507 32077
rect 1545 32063 1579 32077
rect 1545 32043 1549 32063
rect 1549 32043 1579 32063
rect 1617 32043 1651 32077
rect 1689 32063 1723 32077
rect 1689 32043 1719 32063
rect 1719 32043 1723 32063
rect 321 31970 355 32004
rect 393 31970 427 32004
rect 465 31970 499 32004
rect 537 31970 571 32004
rect 609 31970 643 32004
rect 681 31970 715 32004
rect 753 31970 787 32004
rect 825 31970 859 32004
rect 897 31970 931 32004
rect 969 31970 1003 32004
rect 1041 31970 1075 32004
rect 1113 31970 1147 32004
rect 1185 31970 1219 32004
rect 1257 31970 1291 32004
rect 1329 31970 1363 32004
rect 1401 31970 1435 32004
rect 1473 31970 1507 32004
rect 1545 31970 1579 32004
rect 1617 31970 1651 32004
rect 1689 31970 1723 32004
rect 321 31927 355 31931
rect 321 31897 325 31927
rect 325 31897 355 31927
rect 393 31897 427 31931
rect 465 31927 499 31931
rect 465 31897 495 31927
rect 495 31897 499 31927
rect 537 31897 571 31931
rect 609 31927 643 31931
rect 609 31897 631 31927
rect 631 31897 643 31927
rect 681 31897 715 31931
rect 753 31927 787 31931
rect 753 31897 767 31927
rect 767 31897 787 31927
rect 825 31897 859 31931
rect 897 31927 931 31931
rect 897 31897 903 31927
rect 903 31897 931 31927
rect 969 31897 1003 31931
rect 1041 31897 1075 31931
rect 1113 31927 1147 31931
rect 1113 31897 1141 31927
rect 1141 31897 1147 31927
rect 1185 31897 1219 31931
rect 1257 31927 1291 31931
rect 1257 31897 1277 31927
rect 1277 31897 1291 31927
rect 1329 31897 1363 31931
rect 1401 31927 1435 31931
rect 1401 31897 1413 31927
rect 1413 31897 1435 31927
rect 1473 31897 1507 31931
rect 1545 31927 1579 31931
rect 1545 31897 1549 31927
rect 1549 31897 1579 31927
rect 1617 31897 1651 31931
rect 1689 31927 1723 31931
rect 1689 31897 1719 31927
rect 1719 31897 1723 31927
rect 321 31824 355 31858
rect 393 31824 427 31858
rect 465 31824 499 31858
rect 537 31824 571 31858
rect 609 31824 643 31858
rect 681 31824 715 31858
rect 753 31824 787 31858
rect 825 31824 859 31858
rect 897 31824 931 31858
rect 969 31824 1003 31858
rect 1041 31824 1075 31858
rect 1113 31824 1147 31858
rect 1185 31824 1219 31858
rect 1257 31824 1291 31858
rect 1329 31824 1363 31858
rect 1401 31824 1435 31858
rect 1473 31824 1507 31858
rect 1545 31824 1579 31858
rect 1617 31824 1651 31858
rect 1689 31824 1723 31858
rect 321 31757 325 31785
rect 325 31757 355 31785
rect 321 31751 355 31757
rect 393 31751 427 31785
rect 465 31757 495 31785
rect 495 31757 499 31785
rect 465 31751 499 31757
rect 537 31751 571 31785
rect 609 31757 631 31785
rect 631 31757 643 31785
rect 609 31751 643 31757
rect 681 31751 715 31785
rect 753 31757 767 31785
rect 767 31757 787 31785
rect 753 31751 787 31757
rect 825 31751 859 31785
rect 897 31757 903 31785
rect 903 31757 931 31785
rect 897 31751 931 31757
rect 969 31751 1003 31785
rect 1041 31751 1075 31785
rect 1113 31757 1141 31785
rect 1141 31757 1147 31785
rect 1113 31751 1147 31757
rect 1185 31751 1219 31785
rect 1257 31757 1277 31785
rect 1277 31757 1291 31785
rect 1257 31751 1291 31757
rect 1329 31751 1363 31785
rect 1401 31757 1413 31785
rect 1413 31757 1435 31785
rect 1401 31751 1435 31757
rect 1473 31751 1507 31785
rect 1545 31757 1549 31785
rect 1549 31757 1579 31785
rect 1545 31751 1579 31757
rect 1617 31751 1651 31785
rect 1689 31757 1719 31785
rect 1719 31757 1723 31785
rect 1689 31751 1723 31757
rect 321 31678 355 31712
rect 393 31678 427 31712
rect 465 31678 499 31712
rect 537 31678 571 31712
rect 609 31678 643 31712
rect 681 31678 715 31712
rect 753 31678 787 31712
rect 825 31678 859 31712
rect 897 31678 931 31712
rect 969 31678 1003 31712
rect 1041 31678 1075 31712
rect 1113 31678 1147 31712
rect 1185 31678 1219 31712
rect 1257 31678 1291 31712
rect 1329 31678 1363 31712
rect 1401 31678 1435 31712
rect 1473 31678 1507 31712
rect 1545 31678 1579 31712
rect 1617 31678 1651 31712
rect 1689 31678 1723 31712
rect 321 31621 325 31639
rect 325 31621 355 31639
rect 321 31605 355 31621
rect 393 31605 427 31639
rect 465 31621 495 31639
rect 495 31621 499 31639
rect 465 31605 499 31621
rect 537 31605 571 31639
rect 609 31621 631 31639
rect 631 31621 643 31639
rect 609 31605 643 31621
rect 681 31605 715 31639
rect 753 31621 767 31639
rect 767 31621 787 31639
rect 753 31605 787 31621
rect 825 31605 859 31639
rect 897 31621 903 31639
rect 903 31621 931 31639
rect 897 31605 931 31621
rect 969 31605 1003 31639
rect 1041 31605 1075 31639
rect 1113 31621 1141 31639
rect 1141 31621 1147 31639
rect 1113 31605 1147 31621
rect 1185 31605 1219 31639
rect 1257 31621 1277 31639
rect 1277 31621 1291 31639
rect 1257 31605 1291 31621
rect 1329 31605 1363 31639
rect 1401 31621 1413 31639
rect 1413 31621 1435 31639
rect 1401 31605 1435 31621
rect 1473 31605 1507 31639
rect 1545 31621 1549 31639
rect 1549 31621 1579 31639
rect 1545 31605 1579 31621
rect 1617 31605 1651 31639
rect 1689 31621 1719 31639
rect 1719 31621 1723 31639
rect 1689 31605 1723 31621
rect 321 31532 355 31566
rect 393 31532 427 31566
rect 465 31532 499 31566
rect 537 31532 571 31566
rect 609 31532 643 31566
rect 681 31532 715 31566
rect 753 31532 787 31566
rect 825 31532 859 31566
rect 897 31532 931 31566
rect 969 31532 1003 31566
rect 1041 31532 1075 31566
rect 1113 31532 1147 31566
rect 1185 31532 1219 31566
rect 1257 31532 1291 31566
rect 1329 31532 1363 31566
rect 1401 31532 1435 31566
rect 1473 31532 1507 31566
rect 1545 31532 1579 31566
rect 1617 31532 1651 31566
rect 1689 31532 1723 31566
rect 321 31485 325 31493
rect 325 31485 355 31493
rect 321 31459 355 31485
rect 393 31459 427 31493
rect 465 31485 495 31493
rect 495 31485 499 31493
rect 465 31459 499 31485
rect 537 31459 571 31493
rect 609 31485 631 31493
rect 631 31485 643 31493
rect 609 31459 643 31485
rect 681 31459 715 31493
rect 753 31485 767 31493
rect 767 31485 787 31493
rect 753 31459 787 31485
rect 825 31459 859 31493
rect 897 31485 903 31493
rect 903 31485 931 31493
rect 897 31459 931 31485
rect 969 31459 1003 31493
rect 1041 31459 1075 31493
rect 1113 31485 1141 31493
rect 1141 31485 1147 31493
rect 1113 31459 1147 31485
rect 1185 31459 1219 31493
rect 1257 31485 1277 31493
rect 1277 31485 1291 31493
rect 1257 31459 1291 31485
rect 1329 31459 1363 31493
rect 1401 31485 1413 31493
rect 1413 31485 1435 31493
rect 1401 31459 1435 31485
rect 1473 31459 1507 31493
rect 1545 31485 1549 31493
rect 1549 31485 1579 31493
rect 1545 31459 1579 31485
rect 1617 31459 1651 31493
rect 1689 31485 1719 31493
rect 1719 31485 1723 31493
rect 1689 31459 1723 31485
rect 321 31386 355 31420
rect 393 31386 427 31420
rect 465 31386 499 31420
rect 537 31386 571 31420
rect 609 31386 643 31420
rect 681 31386 715 31420
rect 753 31386 787 31420
rect 825 31386 859 31420
rect 897 31386 931 31420
rect 969 31386 1003 31420
rect 1041 31386 1075 31420
rect 1113 31386 1147 31420
rect 1185 31386 1219 31420
rect 1257 31386 1291 31420
rect 1329 31386 1363 31420
rect 1401 31386 1435 31420
rect 1473 31386 1507 31420
rect 1545 31386 1579 31420
rect 1617 31386 1651 31420
rect 1689 31386 1723 31420
rect 321 31313 355 31347
rect 393 31313 427 31347
rect 465 31313 499 31347
rect 537 31313 571 31347
rect 609 31313 643 31347
rect 681 31313 715 31347
rect 753 31313 787 31347
rect 825 31313 859 31347
rect 897 31313 931 31347
rect 969 31313 1003 31347
rect 1041 31313 1075 31347
rect 1113 31313 1147 31347
rect 1185 31313 1219 31347
rect 1257 31313 1291 31347
rect 1329 31313 1363 31347
rect 1401 31313 1435 31347
rect 1473 31313 1507 31347
rect 1545 31313 1579 31347
rect 1617 31313 1651 31347
rect 1689 31313 1723 31347
rect 321 31247 355 31274
rect 321 31240 325 31247
rect 325 31240 355 31247
rect 393 31240 427 31274
rect 465 31247 499 31274
rect 465 31240 495 31247
rect 495 31240 499 31247
rect 537 31240 571 31274
rect 609 31247 643 31274
rect 609 31240 631 31247
rect 631 31240 643 31247
rect 681 31240 715 31274
rect 753 31247 787 31274
rect 753 31240 767 31247
rect 767 31240 787 31247
rect 825 31240 859 31274
rect 897 31247 931 31274
rect 897 31240 903 31247
rect 903 31240 931 31247
rect 969 31240 1003 31274
rect 1041 31240 1075 31274
rect 1113 31247 1147 31274
rect 1113 31240 1141 31247
rect 1141 31240 1147 31247
rect 1185 31240 1219 31274
rect 1257 31247 1291 31274
rect 1257 31240 1277 31247
rect 1277 31240 1291 31247
rect 1329 31240 1363 31274
rect 1401 31247 1435 31274
rect 1401 31240 1413 31247
rect 1413 31240 1435 31247
rect 1473 31240 1507 31274
rect 1545 31247 1579 31274
rect 1545 31240 1549 31247
rect 1549 31240 1579 31247
rect 1617 31240 1651 31274
rect 1689 31247 1723 31274
rect 1689 31240 1719 31247
rect 1719 31240 1723 31247
rect 321 31167 355 31201
rect 393 31167 427 31201
rect 465 31167 499 31201
rect 537 31167 571 31201
rect 609 31167 643 31201
rect 681 31167 715 31201
rect 753 31167 787 31201
rect 825 31167 859 31201
rect 897 31167 931 31201
rect 969 31167 1003 31201
rect 1041 31167 1075 31201
rect 1113 31167 1147 31201
rect 1185 31167 1219 31201
rect 1257 31167 1291 31201
rect 1329 31167 1363 31201
rect 1401 31167 1435 31201
rect 1473 31167 1507 31201
rect 1545 31167 1579 31201
rect 1617 31167 1651 31201
rect 1689 31167 1723 31201
rect 321 31111 355 31128
rect 321 31094 325 31111
rect 325 31094 355 31111
rect 393 31094 427 31128
rect 465 31111 499 31128
rect 465 31094 495 31111
rect 495 31094 499 31111
rect 537 31094 571 31128
rect 609 31111 643 31128
rect 609 31094 631 31111
rect 631 31094 643 31111
rect 681 31094 715 31128
rect 753 31111 787 31128
rect 753 31094 767 31111
rect 767 31094 787 31111
rect 825 31094 859 31128
rect 897 31111 931 31128
rect 897 31094 903 31111
rect 903 31094 931 31111
rect 969 31094 1003 31128
rect 1041 31094 1075 31128
rect 1113 31111 1147 31128
rect 1113 31094 1141 31111
rect 1141 31094 1147 31111
rect 1185 31094 1219 31128
rect 1257 31111 1291 31128
rect 1257 31094 1277 31111
rect 1277 31094 1291 31111
rect 1329 31094 1363 31128
rect 1401 31111 1435 31128
rect 1401 31094 1413 31111
rect 1413 31094 1435 31111
rect 1473 31094 1507 31128
rect 1545 31111 1579 31128
rect 1545 31094 1549 31111
rect 1549 31094 1579 31111
rect 1617 31094 1651 31128
rect 1689 31111 1723 31128
rect 1689 31094 1719 31111
rect 1719 31094 1723 31111
rect 321 31021 355 31055
rect 393 31021 427 31055
rect 465 31021 499 31055
rect 537 31021 571 31055
rect 609 31021 643 31055
rect 681 31021 715 31055
rect 753 31021 787 31055
rect 825 31021 859 31055
rect 897 31021 931 31055
rect 969 31021 1003 31055
rect 1041 31021 1075 31055
rect 1113 31021 1147 31055
rect 1185 31021 1219 31055
rect 1257 31021 1291 31055
rect 1329 31021 1363 31055
rect 1401 31021 1435 31055
rect 1473 31021 1507 31055
rect 1545 31021 1579 31055
rect 1617 31021 1651 31055
rect 1689 31021 1723 31055
rect 321 30975 355 30982
rect 321 30948 325 30975
rect 325 30948 355 30975
rect 393 30948 427 30982
rect 465 30975 499 30982
rect 465 30948 495 30975
rect 495 30948 499 30975
rect 537 30948 571 30982
rect 609 30975 643 30982
rect 609 30948 631 30975
rect 631 30948 643 30975
rect 681 30948 715 30982
rect 753 30975 787 30982
rect 753 30948 767 30975
rect 767 30948 787 30975
rect 825 30948 859 30982
rect 897 30975 931 30982
rect 897 30948 903 30975
rect 903 30948 931 30975
rect 969 30948 1003 30982
rect 1041 30948 1075 30982
rect 1113 30975 1147 30982
rect 1113 30948 1141 30975
rect 1141 30948 1147 30975
rect 1185 30948 1219 30982
rect 1257 30975 1291 30982
rect 1257 30948 1277 30975
rect 1277 30948 1291 30975
rect 1329 30948 1363 30982
rect 1401 30975 1435 30982
rect 1401 30948 1413 30975
rect 1413 30948 1435 30975
rect 1473 30948 1507 30982
rect 1545 30975 1579 30982
rect 1545 30948 1549 30975
rect 1549 30948 1579 30975
rect 1617 30948 1651 30982
rect 1689 30975 1723 30982
rect 1689 30948 1719 30975
rect 1719 30948 1723 30975
rect 321 30875 355 30909
rect 393 30875 427 30909
rect 465 30875 499 30909
rect 537 30875 571 30909
rect 609 30875 643 30909
rect 681 30875 715 30909
rect 753 30875 787 30909
rect 825 30875 859 30909
rect 897 30875 931 30909
rect 969 30875 1003 30909
rect 1041 30875 1075 30909
rect 1113 30875 1147 30909
rect 1185 30875 1219 30909
rect 1257 30875 1291 30909
rect 1329 30875 1363 30909
rect 1401 30875 1435 30909
rect 1473 30875 1507 30909
rect 1545 30875 1579 30909
rect 1617 30875 1651 30909
rect 1689 30875 1723 30909
rect 321 30805 325 30836
rect 325 30805 355 30836
rect 321 30802 355 30805
rect 393 30802 427 30836
rect 465 30805 495 30836
rect 495 30805 499 30836
rect 465 30802 499 30805
rect 537 30802 571 30836
rect 609 30805 631 30836
rect 631 30805 643 30836
rect 609 30802 643 30805
rect 681 30802 715 30836
rect 753 30805 767 30836
rect 767 30805 787 30836
rect 753 30802 787 30805
rect 825 30802 859 30836
rect 897 30805 903 30836
rect 903 30805 931 30836
rect 897 30802 931 30805
rect 969 30802 1003 30836
rect 1041 30802 1075 30836
rect 1113 30805 1141 30836
rect 1141 30805 1147 30836
rect 1113 30802 1147 30805
rect 1185 30802 1219 30836
rect 1257 30805 1277 30836
rect 1277 30805 1291 30836
rect 1257 30802 1291 30805
rect 1329 30802 1363 30836
rect 1401 30805 1413 30836
rect 1413 30805 1435 30836
rect 1401 30802 1435 30805
rect 1473 30802 1507 30836
rect 1545 30805 1549 30836
rect 1549 30805 1579 30836
rect 1545 30802 1579 30805
rect 1617 30802 1651 30836
rect 1689 30805 1719 30836
rect 1719 30805 1723 30836
rect 1689 30802 1723 30805
rect 321 30729 355 30763
rect 393 30729 427 30763
rect 465 30729 499 30763
rect 537 30729 571 30763
rect 609 30729 643 30763
rect 681 30729 715 30763
rect 753 30729 787 30763
rect 825 30729 859 30763
rect 897 30729 931 30763
rect 969 30729 1003 30763
rect 1041 30729 1075 30763
rect 1113 30729 1147 30763
rect 1185 30729 1219 30763
rect 1257 30729 1291 30763
rect 1329 30729 1363 30763
rect 1401 30729 1435 30763
rect 1473 30729 1507 30763
rect 1545 30729 1579 30763
rect 1617 30729 1651 30763
rect 1689 30729 1723 30763
rect 321 30669 325 30690
rect 325 30669 355 30690
rect 321 30656 355 30669
rect 393 30656 427 30690
rect 465 30669 495 30690
rect 495 30669 499 30690
rect 465 30656 499 30669
rect 537 30656 571 30690
rect 609 30669 631 30690
rect 631 30669 643 30690
rect 609 30656 643 30669
rect 681 30656 715 30690
rect 753 30669 767 30690
rect 767 30669 787 30690
rect 753 30656 787 30669
rect 825 30656 859 30690
rect 897 30669 903 30690
rect 903 30669 931 30690
rect 897 30656 931 30669
rect 969 30656 1003 30690
rect 1041 30656 1075 30690
rect 1113 30669 1141 30690
rect 1141 30669 1147 30690
rect 1113 30656 1147 30669
rect 1185 30656 1219 30690
rect 1257 30669 1277 30690
rect 1277 30669 1291 30690
rect 1257 30656 1291 30669
rect 1329 30656 1363 30690
rect 1401 30669 1413 30690
rect 1413 30669 1435 30690
rect 1401 30656 1435 30669
rect 1473 30656 1507 30690
rect 1545 30669 1549 30690
rect 1549 30669 1579 30690
rect 1545 30656 1579 30669
rect 1617 30656 1651 30690
rect 1689 30669 1719 30690
rect 1719 30669 1723 30690
rect 1689 30656 1723 30669
rect 321 30583 355 30617
rect 393 30583 427 30617
rect 465 30583 499 30617
rect 537 30583 571 30617
rect 609 30583 643 30617
rect 681 30583 715 30617
rect 753 30583 787 30617
rect 825 30583 859 30617
rect 897 30583 931 30617
rect 969 30583 1003 30617
rect 1041 30583 1075 30617
rect 1113 30583 1147 30617
rect 1185 30583 1219 30617
rect 1257 30583 1291 30617
rect 1329 30583 1363 30617
rect 1401 30583 1435 30617
rect 1473 30583 1507 30617
rect 1545 30583 1579 30617
rect 1617 30583 1651 30617
rect 1689 30583 1723 30617
rect 321 30533 325 30544
rect 325 30533 355 30544
rect 321 30510 355 30533
rect 393 30510 427 30544
rect 465 30533 495 30544
rect 495 30533 499 30544
rect 465 30510 499 30533
rect 537 30510 571 30544
rect 609 30533 631 30544
rect 631 30533 643 30544
rect 609 30510 643 30533
rect 681 30510 715 30544
rect 753 30533 767 30544
rect 767 30533 787 30544
rect 753 30510 787 30533
rect 825 30510 859 30544
rect 897 30533 903 30544
rect 903 30533 931 30544
rect 897 30510 931 30533
rect 969 30510 1003 30544
rect 1041 30510 1075 30544
rect 1113 30533 1141 30544
rect 1141 30533 1147 30544
rect 1113 30510 1147 30533
rect 1185 30510 1219 30544
rect 1257 30533 1277 30544
rect 1277 30533 1291 30544
rect 1257 30510 1291 30533
rect 1329 30510 1363 30544
rect 1401 30533 1413 30544
rect 1413 30533 1435 30544
rect 1401 30510 1435 30533
rect 1473 30510 1507 30544
rect 1545 30533 1549 30544
rect 1549 30533 1579 30544
rect 1545 30510 1579 30533
rect 1617 30510 1651 30544
rect 1689 30533 1719 30544
rect 1719 30533 1723 30544
rect 1689 30510 1723 30533
rect 321 30437 355 30471
rect 393 30437 427 30471
rect 465 30437 499 30471
rect 537 30437 571 30471
rect 609 30437 643 30471
rect 681 30437 715 30471
rect 753 30437 787 30471
rect 825 30437 859 30471
rect 897 30437 931 30471
rect 969 30437 1003 30471
rect 1041 30437 1075 30471
rect 1113 30437 1147 30471
rect 1185 30437 1219 30471
rect 1257 30437 1291 30471
rect 1329 30437 1363 30471
rect 1401 30437 1435 30471
rect 1473 30437 1507 30471
rect 1545 30437 1579 30471
rect 1617 30437 1651 30471
rect 1689 30437 1723 30471
rect 321 30397 325 30398
rect 325 30397 355 30398
rect 321 30364 355 30397
rect 393 30364 427 30398
rect 465 30397 495 30398
rect 495 30397 499 30398
rect 465 30364 499 30397
rect 537 30364 571 30398
rect 609 30397 631 30398
rect 631 30397 643 30398
rect 609 30364 643 30397
rect 681 30364 715 30398
rect 753 30397 767 30398
rect 767 30397 787 30398
rect 753 30364 787 30397
rect 825 30364 859 30398
rect 897 30397 903 30398
rect 903 30397 931 30398
rect 897 30364 931 30397
rect 969 30364 1003 30398
rect 1041 30364 1075 30398
rect 1113 30397 1141 30398
rect 1141 30397 1147 30398
rect 1113 30364 1147 30397
rect 1185 30364 1219 30398
rect 1257 30397 1277 30398
rect 1277 30397 1291 30398
rect 1257 30364 1291 30397
rect 1329 30364 1363 30398
rect 1401 30397 1413 30398
rect 1413 30397 1435 30398
rect 1401 30364 1435 30397
rect 1473 30364 1507 30398
rect 1545 30397 1549 30398
rect 1549 30397 1579 30398
rect 1545 30364 1579 30397
rect 1617 30364 1651 30398
rect 1689 30397 1719 30398
rect 1719 30397 1723 30398
rect 1689 30364 1723 30397
rect 321 30295 355 30325
rect 321 30291 325 30295
rect 325 30291 355 30295
rect 393 30291 427 30325
rect 465 30295 499 30325
rect 465 30291 495 30295
rect 495 30291 499 30295
rect 537 30291 571 30325
rect 609 30295 643 30325
rect 609 30291 631 30295
rect 631 30291 643 30295
rect 681 30291 715 30325
rect 753 30295 787 30325
rect 753 30291 767 30295
rect 767 30291 787 30295
rect 825 30291 859 30325
rect 897 30295 931 30325
rect 897 30291 903 30295
rect 903 30291 931 30295
rect 969 30291 1003 30325
rect 1041 30291 1075 30325
rect 1113 30295 1147 30325
rect 1113 30291 1141 30295
rect 1141 30291 1147 30295
rect 1185 30291 1219 30325
rect 1257 30295 1291 30325
rect 1257 30291 1277 30295
rect 1277 30291 1291 30295
rect 1329 30291 1363 30325
rect 1401 30295 1435 30325
rect 1401 30291 1413 30295
rect 1413 30291 1435 30295
rect 1473 30291 1507 30325
rect 1545 30295 1579 30325
rect 1545 30291 1549 30295
rect 1549 30291 1579 30295
rect 1617 30291 1651 30325
rect 1689 30295 1723 30325
rect 1689 30291 1719 30295
rect 1719 30291 1723 30295
rect 321 30218 355 30252
rect 393 30218 427 30252
rect 465 30218 499 30252
rect 537 30218 571 30252
rect 609 30218 643 30252
rect 681 30218 715 30252
rect 753 30218 787 30252
rect 825 30218 859 30252
rect 897 30218 931 30252
rect 969 30218 1003 30252
rect 1041 30218 1075 30252
rect 1113 30218 1147 30252
rect 1185 30218 1219 30252
rect 1257 30218 1291 30252
rect 1329 30218 1363 30252
rect 1401 30218 1435 30252
rect 1473 30218 1507 30252
rect 1545 30218 1579 30252
rect 1617 30218 1651 30252
rect 1689 30218 1723 30252
rect 321 30159 355 30179
rect 321 30145 325 30159
rect 325 30145 355 30159
rect 393 30145 427 30179
rect 465 30159 499 30179
rect 465 30145 495 30159
rect 495 30145 499 30159
rect 537 30145 571 30179
rect 609 30159 643 30179
rect 609 30145 631 30159
rect 631 30145 643 30159
rect 681 30145 715 30179
rect 753 30159 787 30179
rect 753 30145 767 30159
rect 767 30145 787 30159
rect 825 30145 859 30179
rect 897 30159 931 30179
rect 897 30145 903 30159
rect 903 30145 931 30159
rect 969 30145 1003 30179
rect 1041 30145 1075 30179
rect 1113 30159 1147 30179
rect 1113 30145 1141 30159
rect 1141 30145 1147 30159
rect 1185 30145 1219 30179
rect 1257 30159 1291 30179
rect 1257 30145 1277 30159
rect 1277 30145 1291 30159
rect 1329 30145 1363 30179
rect 1401 30159 1435 30179
rect 1401 30145 1413 30159
rect 1413 30145 1435 30159
rect 1473 30145 1507 30179
rect 1545 30159 1579 30179
rect 1545 30145 1549 30159
rect 1549 30145 1579 30159
rect 1617 30145 1651 30179
rect 1689 30159 1723 30179
rect 1689 30145 1719 30159
rect 1719 30145 1723 30159
rect 321 30072 355 30106
rect 393 30072 427 30106
rect 465 30072 499 30106
rect 537 30072 571 30106
rect 609 30072 643 30106
rect 681 30072 715 30106
rect 753 30072 787 30106
rect 825 30072 859 30106
rect 897 30072 931 30106
rect 969 30072 1003 30106
rect 1041 30072 1075 30106
rect 1113 30072 1147 30106
rect 1185 30072 1219 30106
rect 1257 30072 1291 30106
rect 1329 30072 1363 30106
rect 1401 30072 1435 30106
rect 1473 30072 1507 30106
rect 1545 30072 1579 30106
rect 1617 30072 1651 30106
rect 1689 30072 1723 30106
rect 321 30023 355 30033
rect 321 29999 325 30023
rect 325 29999 355 30023
rect 393 29999 427 30033
rect 465 30023 499 30033
rect 465 29999 495 30023
rect 495 29999 499 30023
rect 537 29999 571 30033
rect 609 30023 643 30033
rect 609 29999 631 30023
rect 631 29999 643 30023
rect 681 29999 715 30033
rect 753 30023 787 30033
rect 753 29999 767 30023
rect 767 29999 787 30023
rect 825 29999 859 30033
rect 897 30023 931 30033
rect 897 29999 903 30023
rect 903 29999 931 30023
rect 969 29999 1003 30033
rect 1041 29999 1075 30033
rect 1113 30023 1147 30033
rect 1113 29999 1141 30023
rect 1141 29999 1147 30023
rect 1185 29999 1219 30033
rect 1257 30023 1291 30033
rect 1257 29999 1277 30023
rect 1277 29999 1291 30023
rect 1329 29999 1363 30033
rect 1401 30023 1435 30033
rect 1401 29999 1413 30023
rect 1413 29999 1435 30023
rect 1473 29999 1507 30033
rect 1545 30023 1579 30033
rect 1545 29999 1549 30023
rect 1549 29999 1579 30023
rect 1617 29999 1651 30033
rect 1689 30023 1723 30033
rect 1689 29999 1719 30023
rect 1719 29999 1723 30023
rect 321 29926 355 29960
rect 393 29926 427 29960
rect 465 29926 499 29960
rect 537 29926 571 29960
rect 609 29926 643 29960
rect 681 29926 715 29960
rect 753 29926 787 29960
rect 825 29926 859 29960
rect 897 29926 931 29960
rect 969 29926 1003 29960
rect 1041 29926 1075 29960
rect 1113 29926 1147 29960
rect 1185 29926 1219 29960
rect 1257 29926 1291 29960
rect 1329 29926 1363 29960
rect 1401 29926 1435 29960
rect 1473 29926 1507 29960
rect 1545 29926 1579 29960
rect 1617 29926 1651 29960
rect 1689 29926 1723 29960
rect 321 29853 325 29887
rect 325 29853 355 29887
rect 393 29853 427 29887
rect 465 29853 495 29887
rect 495 29853 499 29887
rect 537 29853 571 29887
rect 609 29853 631 29887
rect 631 29853 643 29887
rect 681 29853 715 29887
rect 753 29853 767 29887
rect 767 29853 787 29887
rect 825 29853 859 29887
rect 897 29853 903 29887
rect 903 29853 931 29887
rect 969 29853 1003 29887
rect 1041 29853 1075 29887
rect 1113 29853 1141 29887
rect 1141 29853 1147 29887
rect 1185 29853 1219 29887
rect 1257 29853 1277 29887
rect 1277 29853 1291 29887
rect 1329 29853 1363 29887
rect 1401 29853 1413 29887
rect 1413 29853 1435 29887
rect 1473 29853 1507 29887
rect 1545 29853 1549 29887
rect 1549 29853 1579 29887
rect 1617 29853 1651 29887
rect 1689 29853 1719 29887
rect 1719 29853 1723 29887
rect 321 29780 355 29814
rect 393 29780 427 29814
rect 465 29780 499 29814
rect 537 29780 571 29814
rect 609 29780 643 29814
rect 681 29780 715 29814
rect 753 29780 787 29814
rect 825 29780 859 29814
rect 897 29780 931 29814
rect 969 29780 1003 29814
rect 1041 29780 1075 29814
rect 1113 29780 1147 29814
rect 1185 29780 1219 29814
rect 1257 29780 1291 29814
rect 1329 29780 1363 29814
rect 1401 29780 1435 29814
rect 1473 29780 1507 29814
rect 1545 29780 1579 29814
rect 1617 29780 1651 29814
rect 1689 29780 1723 29814
rect 321 29717 325 29741
rect 325 29717 355 29741
rect 321 29707 355 29717
rect 393 29707 427 29741
rect 465 29717 495 29741
rect 495 29717 499 29741
rect 465 29707 499 29717
rect 537 29707 571 29741
rect 609 29717 631 29741
rect 631 29717 643 29741
rect 609 29707 643 29717
rect 681 29707 715 29741
rect 753 29717 767 29741
rect 767 29717 787 29741
rect 753 29707 787 29717
rect 825 29707 859 29741
rect 897 29717 903 29741
rect 903 29717 931 29741
rect 897 29707 931 29717
rect 969 29707 1003 29741
rect 1041 29707 1075 29741
rect 1113 29717 1141 29741
rect 1141 29717 1147 29741
rect 1113 29707 1147 29717
rect 1185 29707 1219 29741
rect 1257 29717 1277 29741
rect 1277 29717 1291 29741
rect 1257 29707 1291 29717
rect 1329 29707 1363 29741
rect 1401 29717 1413 29741
rect 1413 29717 1435 29741
rect 1401 29707 1435 29717
rect 1473 29707 1507 29741
rect 1545 29717 1549 29741
rect 1549 29717 1579 29741
rect 1545 29707 1579 29717
rect 1617 29707 1651 29741
rect 1689 29717 1719 29741
rect 1719 29717 1723 29741
rect 1689 29707 1723 29717
rect 321 29634 355 29668
rect 393 29634 427 29668
rect 465 29634 499 29668
rect 537 29634 571 29668
rect 609 29634 643 29668
rect 681 29634 715 29668
rect 753 29634 787 29668
rect 825 29634 859 29668
rect 897 29634 931 29668
rect 969 29634 1003 29668
rect 1041 29634 1075 29668
rect 1113 29634 1147 29668
rect 1185 29634 1219 29668
rect 1257 29634 1291 29668
rect 1329 29634 1363 29668
rect 1401 29634 1435 29668
rect 1473 29634 1507 29668
rect 1545 29634 1579 29668
rect 1617 29634 1651 29668
rect 1689 29634 1723 29668
rect 7876 39917 7880 39943
rect 7880 39917 7914 39943
rect 7914 39917 8016 39943
rect 8016 39917 8050 39943
rect 8050 39917 8152 39943
rect 8152 39917 8186 39943
rect 8186 39917 8288 39943
rect 8288 39917 8322 39943
rect 8322 39917 8424 39943
rect 8424 39917 8458 39943
rect 8458 39917 8560 39943
rect 8560 39917 8594 39943
rect 8594 39917 8696 39943
rect 8696 39917 8730 39943
rect 8730 39917 8832 39943
rect 8832 39917 8866 39943
rect 8866 39917 8968 39943
rect 8968 39917 9002 39943
rect 9002 39917 9104 39943
rect 9104 39917 9138 39943
rect 9138 39917 9240 39943
rect 9240 39917 9274 39943
rect 9274 39917 9278 39943
rect 7876 39815 9278 39917
rect 7876 39781 7880 39815
rect 7880 39781 7914 39815
rect 7914 39781 8016 39815
rect 8016 39781 8050 39815
rect 8050 39781 8152 39815
rect 8152 39781 8186 39815
rect 8186 39781 8288 39815
rect 8288 39781 8322 39815
rect 8322 39781 8424 39815
rect 8424 39781 8458 39815
rect 8458 39781 8560 39815
rect 8560 39781 8594 39815
rect 8594 39781 8696 39815
rect 8696 39781 8730 39815
rect 8730 39781 8832 39815
rect 8832 39781 8866 39815
rect 8866 39781 8968 39815
rect 8968 39781 9002 39815
rect 9002 39781 9104 39815
rect 9104 39781 9138 39815
rect 9138 39781 9240 39815
rect 9240 39781 9274 39815
rect 9274 39781 9278 39815
rect 7876 39679 9278 39781
rect 7876 39645 7880 39679
rect 7880 39645 7914 39679
rect 7914 39645 8016 39679
rect 8016 39645 8050 39679
rect 8050 39645 8152 39679
rect 8152 39645 8186 39679
rect 8186 39645 8288 39679
rect 8288 39645 8322 39679
rect 8322 39645 8424 39679
rect 8424 39645 8458 39679
rect 8458 39645 8560 39679
rect 8560 39645 8594 39679
rect 8594 39645 8696 39679
rect 8696 39645 8730 39679
rect 8730 39645 8832 39679
rect 8832 39645 8866 39679
rect 8866 39645 8968 39679
rect 8968 39645 9002 39679
rect 9002 39645 9104 39679
rect 9104 39645 9138 39679
rect 9138 39645 9240 39679
rect 9240 39645 9274 39679
rect 9274 39645 9278 39679
rect 7876 39543 9278 39645
rect 7876 39509 7880 39543
rect 7880 39509 7914 39543
rect 7914 39509 8016 39543
rect 8016 39509 8050 39543
rect 8050 39509 8152 39543
rect 8152 39509 8186 39543
rect 8186 39509 8288 39543
rect 8288 39509 8322 39543
rect 8322 39509 8424 39543
rect 8424 39509 8458 39543
rect 8458 39509 8560 39543
rect 8560 39509 8594 39543
rect 8594 39509 8696 39543
rect 8696 39509 8730 39543
rect 8730 39509 8832 39543
rect 8832 39509 8866 39543
rect 8866 39509 8968 39543
rect 8968 39509 9002 39543
rect 9002 39509 9104 39543
rect 9104 39509 9138 39543
rect 9138 39509 9240 39543
rect 9240 39509 9274 39543
rect 9274 39509 9278 39543
rect 7876 39407 9278 39509
rect 7876 39373 7880 39407
rect 7880 39373 7914 39407
rect 7914 39373 8016 39407
rect 8016 39373 8050 39407
rect 8050 39373 8152 39407
rect 8152 39373 8186 39407
rect 8186 39373 8288 39407
rect 8288 39373 8322 39407
rect 8322 39373 8424 39407
rect 8424 39373 8458 39407
rect 8458 39373 8560 39407
rect 8560 39373 8594 39407
rect 8594 39373 8696 39407
rect 8696 39373 8730 39407
rect 8730 39373 8832 39407
rect 8832 39373 8866 39407
rect 8866 39373 8968 39407
rect 8968 39373 9002 39407
rect 9002 39373 9104 39407
rect 9104 39373 9138 39407
rect 9138 39373 9240 39407
rect 9240 39373 9274 39407
rect 9274 39373 9278 39407
rect 7876 39271 9278 39373
rect 7876 39237 7880 39271
rect 7880 39237 7914 39271
rect 7914 39237 8016 39271
rect 8016 39237 8050 39271
rect 8050 39237 8152 39271
rect 8152 39237 8186 39271
rect 8186 39237 8288 39271
rect 8288 39237 8322 39271
rect 8322 39237 8424 39271
rect 8424 39237 8458 39271
rect 8458 39237 8560 39271
rect 8560 39237 8594 39271
rect 8594 39237 8696 39271
rect 8696 39237 8730 39271
rect 8730 39237 8832 39271
rect 8832 39237 8866 39271
rect 8866 39237 8968 39271
rect 8968 39237 9002 39271
rect 9002 39237 9104 39271
rect 9104 39237 9138 39271
rect 9138 39237 9240 39271
rect 9240 39237 9274 39271
rect 9274 39237 9278 39271
rect 7876 39135 9278 39237
rect 7876 39101 7880 39135
rect 7880 39101 7914 39135
rect 7914 39101 8016 39135
rect 8016 39101 8050 39135
rect 8050 39101 8152 39135
rect 8152 39101 8186 39135
rect 8186 39101 8288 39135
rect 8288 39101 8322 39135
rect 8322 39101 8424 39135
rect 8424 39101 8458 39135
rect 8458 39101 8560 39135
rect 8560 39101 8594 39135
rect 8594 39101 8696 39135
rect 8696 39101 8730 39135
rect 8730 39101 8832 39135
rect 8832 39101 8866 39135
rect 8866 39101 8968 39135
rect 8968 39101 9002 39135
rect 9002 39101 9104 39135
rect 9104 39101 9138 39135
rect 9138 39101 9240 39135
rect 9240 39101 9274 39135
rect 9274 39101 9278 39135
rect 7876 38999 9278 39101
rect 7876 38965 7880 38999
rect 7880 38965 7914 38999
rect 7914 38965 8016 38999
rect 8016 38965 8050 38999
rect 8050 38965 8152 38999
rect 8152 38965 8186 38999
rect 8186 38965 8288 38999
rect 8288 38965 8322 38999
rect 8322 38965 8424 38999
rect 8424 38965 8458 38999
rect 8458 38965 8560 38999
rect 8560 38965 8594 38999
rect 8594 38965 8696 38999
rect 8696 38965 8730 38999
rect 8730 38965 8832 38999
rect 8832 38965 8866 38999
rect 8866 38965 8968 38999
rect 8968 38965 9002 38999
rect 9002 38965 9104 38999
rect 9104 38965 9138 38999
rect 9138 38965 9240 38999
rect 9240 38965 9274 38999
rect 9274 38965 9278 38999
rect 7876 38863 9278 38965
rect 7876 38829 7880 38863
rect 7880 38829 7914 38863
rect 7914 38829 8016 38863
rect 8016 38829 8050 38863
rect 8050 38829 8152 38863
rect 8152 38829 8186 38863
rect 8186 38829 8288 38863
rect 8288 38829 8322 38863
rect 8322 38829 8424 38863
rect 8424 38829 8458 38863
rect 8458 38829 8560 38863
rect 8560 38829 8594 38863
rect 8594 38829 8696 38863
rect 8696 38829 8730 38863
rect 8730 38829 8832 38863
rect 8832 38829 8866 38863
rect 8866 38829 8968 38863
rect 8968 38829 9002 38863
rect 9002 38829 9104 38863
rect 9104 38829 9138 38863
rect 9138 38829 9240 38863
rect 9240 38829 9274 38863
rect 9274 38829 9278 38863
rect 7876 38727 9278 38829
rect 7876 38693 7880 38727
rect 7880 38693 7914 38727
rect 7914 38693 8016 38727
rect 8016 38693 8050 38727
rect 8050 38693 8152 38727
rect 8152 38693 8186 38727
rect 8186 38693 8288 38727
rect 8288 38693 8322 38727
rect 8322 38693 8424 38727
rect 8424 38693 8458 38727
rect 8458 38693 8560 38727
rect 8560 38693 8594 38727
rect 8594 38693 8696 38727
rect 8696 38693 8730 38727
rect 8730 38693 8832 38727
rect 8832 38693 8866 38727
rect 8866 38693 8968 38727
rect 8968 38693 9002 38727
rect 9002 38693 9104 38727
rect 9104 38693 9138 38727
rect 9138 38693 9240 38727
rect 9240 38693 9274 38727
rect 9274 38693 9278 38727
rect 7876 38591 9278 38693
rect 7876 38557 7880 38591
rect 7880 38557 7914 38591
rect 7914 38557 8016 38591
rect 8016 38557 8050 38591
rect 8050 38557 8152 38591
rect 8152 38557 8186 38591
rect 8186 38557 8288 38591
rect 8288 38557 8322 38591
rect 8322 38557 8424 38591
rect 8424 38557 8458 38591
rect 8458 38557 8560 38591
rect 8560 38557 8594 38591
rect 8594 38557 8696 38591
rect 8696 38557 8730 38591
rect 8730 38557 8832 38591
rect 8832 38557 8866 38591
rect 8866 38557 8968 38591
rect 8968 38557 9002 38591
rect 9002 38557 9104 38591
rect 9104 38557 9138 38591
rect 9138 38557 9240 38591
rect 9240 38557 9274 38591
rect 9274 38557 9278 38591
rect 7876 38455 9278 38557
rect 7876 38421 7880 38455
rect 7880 38421 7914 38455
rect 7914 38421 8016 38455
rect 8016 38421 8050 38455
rect 8050 38421 8152 38455
rect 8152 38421 8186 38455
rect 8186 38421 8288 38455
rect 8288 38421 8322 38455
rect 8322 38421 8424 38455
rect 8424 38421 8458 38455
rect 8458 38421 8560 38455
rect 8560 38421 8594 38455
rect 8594 38421 8696 38455
rect 8696 38421 8730 38455
rect 8730 38421 8832 38455
rect 8832 38421 8866 38455
rect 8866 38421 8968 38455
rect 8968 38421 9002 38455
rect 9002 38421 9104 38455
rect 9104 38421 9138 38455
rect 9138 38421 9240 38455
rect 9240 38421 9274 38455
rect 9274 38421 9278 38455
rect 7876 38319 9278 38421
rect 7876 38285 7880 38319
rect 7880 38285 7914 38319
rect 7914 38285 8016 38319
rect 8016 38285 8050 38319
rect 8050 38285 8152 38319
rect 8152 38285 8186 38319
rect 8186 38285 8288 38319
rect 8288 38285 8322 38319
rect 8322 38285 8424 38319
rect 8424 38285 8458 38319
rect 8458 38285 8560 38319
rect 8560 38285 8594 38319
rect 8594 38285 8696 38319
rect 8696 38285 8730 38319
rect 8730 38285 8832 38319
rect 8832 38285 8866 38319
rect 8866 38285 8968 38319
rect 8968 38285 9002 38319
rect 9002 38285 9104 38319
rect 9104 38285 9138 38319
rect 9138 38285 9240 38319
rect 9240 38285 9274 38319
rect 9274 38285 9278 38319
rect 7876 38183 9278 38285
rect 7876 38149 7880 38183
rect 7880 38149 7914 38183
rect 7914 38149 8016 38183
rect 8016 38149 8050 38183
rect 8050 38149 8152 38183
rect 8152 38149 8186 38183
rect 8186 38149 8288 38183
rect 8288 38149 8322 38183
rect 8322 38149 8424 38183
rect 8424 38149 8458 38183
rect 8458 38149 8560 38183
rect 8560 38149 8594 38183
rect 8594 38149 8696 38183
rect 8696 38149 8730 38183
rect 8730 38149 8832 38183
rect 8832 38149 8866 38183
rect 8866 38149 8968 38183
rect 8968 38149 9002 38183
rect 9002 38149 9104 38183
rect 9104 38149 9138 38183
rect 9138 38149 9240 38183
rect 9240 38149 9274 38183
rect 9274 38149 9278 38183
rect 7876 38047 9278 38149
rect 7876 38013 7880 38047
rect 7880 38013 7914 38047
rect 7914 38013 8016 38047
rect 8016 38013 8050 38047
rect 8050 38013 8152 38047
rect 8152 38013 8186 38047
rect 8186 38013 8288 38047
rect 8288 38013 8322 38047
rect 8322 38013 8424 38047
rect 8424 38013 8458 38047
rect 8458 38013 8560 38047
rect 8560 38013 8594 38047
rect 8594 38013 8696 38047
rect 8696 38013 8730 38047
rect 8730 38013 8832 38047
rect 8832 38013 8866 38047
rect 8866 38013 8968 38047
rect 8968 38013 9002 38047
rect 9002 38013 9104 38047
rect 9104 38013 9138 38047
rect 9138 38013 9240 38047
rect 9240 38013 9274 38047
rect 9274 38013 9278 38047
rect 7876 37911 9278 38013
rect 7876 37877 7880 37911
rect 7880 37877 7914 37911
rect 7914 37877 8016 37911
rect 8016 37877 8050 37911
rect 8050 37877 8152 37911
rect 8152 37877 8186 37911
rect 8186 37877 8288 37911
rect 8288 37877 8322 37911
rect 8322 37877 8424 37911
rect 8424 37877 8458 37911
rect 8458 37877 8560 37911
rect 8560 37877 8594 37911
rect 8594 37877 8696 37911
rect 8696 37877 8730 37911
rect 8730 37877 8832 37911
rect 8832 37877 8866 37911
rect 8866 37877 8968 37911
rect 8968 37877 9002 37911
rect 9002 37877 9104 37911
rect 9104 37877 9138 37911
rect 9138 37877 9240 37911
rect 9240 37877 9274 37911
rect 9274 37877 9278 37911
rect 7876 37775 9278 37877
rect 7876 37741 7880 37775
rect 7880 37741 7914 37775
rect 7914 37741 8016 37775
rect 8016 37741 8050 37775
rect 8050 37741 8152 37775
rect 8152 37741 8186 37775
rect 8186 37741 8288 37775
rect 8288 37741 8322 37775
rect 8322 37741 8424 37775
rect 8424 37741 8458 37775
rect 8458 37741 8560 37775
rect 8560 37741 8594 37775
rect 8594 37741 8696 37775
rect 8696 37741 8730 37775
rect 8730 37741 8832 37775
rect 8832 37741 8866 37775
rect 8866 37741 8968 37775
rect 8968 37741 9002 37775
rect 9002 37741 9104 37775
rect 9104 37741 9138 37775
rect 9138 37741 9240 37775
rect 9240 37741 9274 37775
rect 9274 37741 9278 37775
rect 7876 37639 9278 37741
rect 7876 37605 7880 37639
rect 7880 37605 7914 37639
rect 7914 37605 8016 37639
rect 8016 37605 8050 37639
rect 8050 37605 8152 37639
rect 8152 37605 8186 37639
rect 8186 37605 8288 37639
rect 8288 37605 8322 37639
rect 8322 37605 8424 37639
rect 8424 37605 8458 37639
rect 8458 37605 8560 37639
rect 8560 37605 8594 37639
rect 8594 37605 8696 37639
rect 8696 37605 8730 37639
rect 8730 37605 8832 37639
rect 8832 37605 8866 37639
rect 8866 37605 8968 37639
rect 8968 37605 9002 37639
rect 9002 37605 9104 37639
rect 9104 37605 9138 37639
rect 9138 37605 9240 37639
rect 9240 37605 9274 37639
rect 9274 37605 9278 37639
rect 7876 37503 9278 37605
rect 7876 37469 7880 37503
rect 7880 37469 7914 37503
rect 7914 37469 8016 37503
rect 8016 37469 8050 37503
rect 8050 37469 8152 37503
rect 8152 37469 8186 37503
rect 8186 37469 8288 37503
rect 8288 37469 8322 37503
rect 8322 37469 8424 37503
rect 8424 37469 8458 37503
rect 8458 37469 8560 37503
rect 8560 37469 8594 37503
rect 8594 37469 8696 37503
rect 8696 37469 8730 37503
rect 8730 37469 8832 37503
rect 8832 37469 8866 37503
rect 8866 37469 8968 37503
rect 8968 37469 9002 37503
rect 9002 37469 9104 37503
rect 9104 37469 9138 37503
rect 9138 37469 9240 37503
rect 9240 37469 9274 37503
rect 9274 37469 9278 37503
rect 7876 37367 9278 37469
rect 7876 37333 7880 37367
rect 7880 37333 7914 37367
rect 7914 37333 8016 37367
rect 8016 37333 8050 37367
rect 8050 37333 8152 37367
rect 8152 37333 8186 37367
rect 8186 37333 8288 37367
rect 8288 37333 8322 37367
rect 8322 37333 8424 37367
rect 8424 37333 8458 37367
rect 8458 37333 8560 37367
rect 8560 37333 8594 37367
rect 8594 37333 8696 37367
rect 8696 37333 8730 37367
rect 8730 37333 8832 37367
rect 8832 37333 8866 37367
rect 8866 37333 8968 37367
rect 8968 37333 9002 37367
rect 9002 37333 9104 37367
rect 9104 37333 9138 37367
rect 9138 37333 9240 37367
rect 9240 37333 9274 37367
rect 9274 37333 9278 37367
rect 7876 37231 9278 37333
rect 7876 37197 7880 37231
rect 7880 37197 7914 37231
rect 7914 37197 8016 37231
rect 8016 37197 8050 37231
rect 8050 37197 8152 37231
rect 8152 37197 8186 37231
rect 8186 37197 8288 37231
rect 8288 37197 8322 37231
rect 8322 37197 8424 37231
rect 8424 37197 8458 37231
rect 8458 37197 8560 37231
rect 8560 37197 8594 37231
rect 8594 37197 8696 37231
rect 8696 37197 8730 37231
rect 8730 37197 8832 37231
rect 8832 37197 8866 37231
rect 8866 37197 8968 37231
rect 8968 37197 9002 37231
rect 9002 37197 9104 37231
rect 9104 37197 9138 37231
rect 9138 37197 9240 37231
rect 9240 37197 9274 37231
rect 9274 37197 9278 37231
rect 7876 37095 9278 37197
rect 7876 37061 7880 37095
rect 7880 37061 7914 37095
rect 7914 37061 8016 37095
rect 8016 37061 8050 37095
rect 8050 37061 8152 37095
rect 8152 37061 8186 37095
rect 8186 37061 8288 37095
rect 8288 37061 8322 37095
rect 8322 37061 8424 37095
rect 8424 37061 8458 37095
rect 8458 37061 8560 37095
rect 8560 37061 8594 37095
rect 8594 37061 8696 37095
rect 8696 37061 8730 37095
rect 8730 37061 8832 37095
rect 8832 37061 8866 37095
rect 8866 37061 8968 37095
rect 8968 37061 9002 37095
rect 9002 37061 9104 37095
rect 9104 37061 9138 37095
rect 9138 37061 9240 37095
rect 9240 37061 9274 37095
rect 9274 37061 9278 37095
rect 7876 36959 9278 37061
rect 7876 36925 7880 36959
rect 7880 36925 7914 36959
rect 7914 36925 8016 36959
rect 8016 36925 8050 36959
rect 8050 36925 8152 36959
rect 8152 36925 8186 36959
rect 8186 36925 8288 36959
rect 8288 36925 8322 36959
rect 8322 36925 8424 36959
rect 8424 36925 8458 36959
rect 8458 36925 8560 36959
rect 8560 36925 8594 36959
rect 8594 36925 8696 36959
rect 8696 36925 8730 36959
rect 8730 36925 8832 36959
rect 8832 36925 8866 36959
rect 8866 36925 8968 36959
rect 8968 36925 9002 36959
rect 9002 36925 9104 36959
rect 9104 36925 9138 36959
rect 9138 36925 9240 36959
rect 9240 36925 9274 36959
rect 9274 36925 9278 36959
rect 7876 36823 9278 36925
rect 7876 36789 7880 36823
rect 7880 36789 7914 36823
rect 7914 36789 8016 36823
rect 8016 36789 8050 36823
rect 8050 36789 8152 36823
rect 8152 36789 8186 36823
rect 8186 36789 8288 36823
rect 8288 36789 8322 36823
rect 8322 36789 8424 36823
rect 8424 36789 8458 36823
rect 8458 36789 8560 36823
rect 8560 36789 8594 36823
rect 8594 36789 8696 36823
rect 8696 36789 8730 36823
rect 8730 36789 8832 36823
rect 8832 36789 8866 36823
rect 8866 36789 8968 36823
rect 8968 36789 9002 36823
rect 9002 36789 9104 36823
rect 9104 36789 9138 36823
rect 9138 36789 9240 36823
rect 9240 36789 9274 36823
rect 9274 36789 9278 36823
rect 7876 36687 9278 36789
rect 7876 36653 7880 36687
rect 7880 36653 7914 36687
rect 7914 36653 8016 36687
rect 8016 36653 8050 36687
rect 8050 36653 8152 36687
rect 8152 36653 8186 36687
rect 8186 36653 8288 36687
rect 8288 36653 8322 36687
rect 8322 36653 8424 36687
rect 8424 36653 8458 36687
rect 8458 36653 8560 36687
rect 8560 36653 8594 36687
rect 8594 36653 8696 36687
rect 8696 36653 8730 36687
rect 8730 36653 8832 36687
rect 8832 36653 8866 36687
rect 8866 36653 8968 36687
rect 8968 36653 9002 36687
rect 9002 36653 9104 36687
rect 9104 36653 9138 36687
rect 9138 36653 9240 36687
rect 9240 36653 9274 36687
rect 9274 36653 9278 36687
rect 7876 36551 9278 36653
rect 7876 36517 7880 36551
rect 7880 36517 7914 36551
rect 7914 36517 8016 36551
rect 8016 36517 8050 36551
rect 8050 36517 8152 36551
rect 8152 36517 8186 36551
rect 8186 36517 8288 36551
rect 8288 36517 8322 36551
rect 8322 36517 8424 36551
rect 8424 36517 8458 36551
rect 8458 36517 8560 36551
rect 8560 36517 8594 36551
rect 8594 36517 8696 36551
rect 8696 36517 8730 36551
rect 8730 36517 8832 36551
rect 8832 36517 8866 36551
rect 8866 36517 8968 36551
rect 8968 36517 9002 36551
rect 9002 36517 9104 36551
rect 9104 36517 9138 36551
rect 9138 36517 9240 36551
rect 9240 36517 9274 36551
rect 9274 36517 9278 36551
rect 7876 36415 9278 36517
rect 7876 36381 7880 36415
rect 7880 36381 7914 36415
rect 7914 36381 8016 36415
rect 8016 36381 8050 36415
rect 8050 36381 8152 36415
rect 8152 36381 8186 36415
rect 8186 36381 8288 36415
rect 8288 36381 8322 36415
rect 8322 36381 8424 36415
rect 8424 36381 8458 36415
rect 8458 36381 8560 36415
rect 8560 36381 8594 36415
rect 8594 36381 8696 36415
rect 8696 36381 8730 36415
rect 8730 36381 8832 36415
rect 8832 36381 8866 36415
rect 8866 36381 8968 36415
rect 8968 36381 9002 36415
rect 9002 36381 9104 36415
rect 9104 36381 9138 36415
rect 9138 36381 9240 36415
rect 9240 36381 9274 36415
rect 9274 36381 9278 36415
rect 7876 36279 9278 36381
rect 7876 36245 7880 36279
rect 7880 36245 7914 36279
rect 7914 36245 8016 36279
rect 8016 36245 8050 36279
rect 8050 36245 8152 36279
rect 8152 36245 8186 36279
rect 8186 36245 8288 36279
rect 8288 36245 8322 36279
rect 8322 36245 8424 36279
rect 8424 36245 8458 36279
rect 8458 36245 8560 36279
rect 8560 36245 8594 36279
rect 8594 36245 8696 36279
rect 8696 36245 8730 36279
rect 8730 36245 8832 36279
rect 8832 36245 8866 36279
rect 8866 36245 8968 36279
rect 8968 36245 9002 36279
rect 9002 36245 9104 36279
rect 9104 36245 9138 36279
rect 9138 36245 9240 36279
rect 9240 36245 9274 36279
rect 9274 36245 9278 36279
rect 7876 36143 9278 36245
rect 7876 36109 7880 36143
rect 7880 36109 7914 36143
rect 7914 36109 8016 36143
rect 8016 36109 8050 36143
rect 8050 36109 8152 36143
rect 8152 36109 8186 36143
rect 8186 36109 8288 36143
rect 8288 36109 8322 36143
rect 8322 36109 8424 36143
rect 8424 36109 8458 36143
rect 8458 36109 8560 36143
rect 8560 36109 8594 36143
rect 8594 36109 8696 36143
rect 8696 36109 8730 36143
rect 8730 36109 8832 36143
rect 8832 36109 8866 36143
rect 8866 36109 8968 36143
rect 8968 36109 9002 36143
rect 9002 36109 9104 36143
rect 9104 36109 9138 36143
rect 9138 36109 9240 36143
rect 9240 36109 9274 36143
rect 9274 36109 9278 36143
rect 7876 36007 9278 36109
rect 7876 35973 7880 36007
rect 7880 35973 7914 36007
rect 7914 35973 8016 36007
rect 8016 35973 8050 36007
rect 8050 35973 8152 36007
rect 8152 35973 8186 36007
rect 8186 35973 8288 36007
rect 8288 35973 8322 36007
rect 8322 35973 8424 36007
rect 8424 35973 8458 36007
rect 8458 35973 8560 36007
rect 8560 35973 8594 36007
rect 8594 35973 8696 36007
rect 8696 35973 8730 36007
rect 8730 35973 8832 36007
rect 8832 35973 8866 36007
rect 8866 35973 8968 36007
rect 8968 35973 9002 36007
rect 9002 35973 9104 36007
rect 9104 35973 9138 36007
rect 9138 35973 9240 36007
rect 9240 35973 9274 36007
rect 9274 35973 9278 36007
rect 7876 35871 9278 35973
rect 7876 35837 7880 35871
rect 7880 35837 7914 35871
rect 7914 35837 8016 35871
rect 8016 35837 8050 35871
rect 8050 35837 8152 35871
rect 8152 35837 8186 35871
rect 8186 35837 8288 35871
rect 8288 35837 8322 35871
rect 8322 35837 8424 35871
rect 8424 35837 8458 35871
rect 8458 35837 8560 35871
rect 8560 35837 8594 35871
rect 8594 35837 8696 35871
rect 8696 35837 8730 35871
rect 8730 35837 8832 35871
rect 8832 35837 8866 35871
rect 8866 35837 8968 35871
rect 8968 35837 9002 35871
rect 9002 35837 9104 35871
rect 9104 35837 9138 35871
rect 9138 35837 9240 35871
rect 9240 35837 9274 35871
rect 9274 35837 9278 35871
rect 7876 35735 9278 35837
rect 7876 35701 7880 35735
rect 7880 35701 7914 35735
rect 7914 35701 8016 35735
rect 8016 35701 8050 35735
rect 8050 35701 8152 35735
rect 8152 35701 8186 35735
rect 8186 35701 8288 35735
rect 8288 35701 8322 35735
rect 8322 35701 8424 35735
rect 8424 35701 8458 35735
rect 8458 35701 8560 35735
rect 8560 35701 8594 35735
rect 8594 35701 8696 35735
rect 8696 35701 8730 35735
rect 8730 35701 8832 35735
rect 8832 35701 8866 35735
rect 8866 35701 8968 35735
rect 8968 35701 9002 35735
rect 9002 35701 9104 35735
rect 9104 35701 9138 35735
rect 9138 35701 9240 35735
rect 9240 35701 9274 35735
rect 9274 35701 9278 35735
rect 7876 35599 9278 35701
rect 7876 35565 7880 35599
rect 7880 35565 7914 35599
rect 7914 35565 8016 35599
rect 8016 35565 8050 35599
rect 8050 35565 8152 35599
rect 8152 35565 8186 35599
rect 8186 35565 8288 35599
rect 8288 35565 8322 35599
rect 8322 35565 8424 35599
rect 8424 35565 8458 35599
rect 8458 35565 8560 35599
rect 8560 35565 8594 35599
rect 8594 35565 8696 35599
rect 8696 35565 8730 35599
rect 8730 35565 8832 35599
rect 8832 35565 8866 35599
rect 8866 35565 8968 35599
rect 8968 35565 9002 35599
rect 9002 35565 9104 35599
rect 9104 35565 9138 35599
rect 9138 35565 9240 35599
rect 9240 35565 9274 35599
rect 9274 35565 9278 35599
rect 7876 35463 9278 35565
rect 7876 35429 7880 35463
rect 7880 35429 7914 35463
rect 7914 35429 8016 35463
rect 8016 35429 8050 35463
rect 8050 35429 8152 35463
rect 8152 35429 8186 35463
rect 8186 35429 8288 35463
rect 8288 35429 8322 35463
rect 8322 35429 8424 35463
rect 8424 35429 8458 35463
rect 8458 35429 8560 35463
rect 8560 35429 8594 35463
rect 8594 35429 8696 35463
rect 8696 35429 8730 35463
rect 8730 35429 8832 35463
rect 8832 35429 8866 35463
rect 8866 35429 8968 35463
rect 8968 35429 9002 35463
rect 9002 35429 9104 35463
rect 9104 35429 9138 35463
rect 9138 35429 9240 35463
rect 9240 35429 9274 35463
rect 9274 35429 9278 35463
rect 7876 35327 9278 35429
rect 7876 35293 7880 35327
rect 7880 35293 7914 35327
rect 7914 35293 8016 35327
rect 8016 35293 8050 35327
rect 8050 35293 8152 35327
rect 8152 35293 8186 35327
rect 8186 35293 8288 35327
rect 8288 35293 8322 35327
rect 8322 35293 8424 35327
rect 8424 35293 8458 35327
rect 8458 35293 8560 35327
rect 8560 35293 8594 35327
rect 8594 35293 8696 35327
rect 8696 35293 8730 35327
rect 8730 35293 8832 35327
rect 8832 35293 8866 35327
rect 8866 35293 8968 35327
rect 8968 35293 9002 35327
rect 9002 35293 9104 35327
rect 9104 35293 9138 35327
rect 9138 35293 9240 35327
rect 9240 35293 9274 35327
rect 9274 35293 9278 35327
rect 7876 35191 9278 35293
rect 7876 35157 7880 35191
rect 7880 35157 7914 35191
rect 7914 35157 8016 35191
rect 8016 35157 8050 35191
rect 8050 35157 8152 35191
rect 8152 35157 8186 35191
rect 8186 35157 8288 35191
rect 8288 35157 8322 35191
rect 8322 35157 8424 35191
rect 8424 35157 8458 35191
rect 8458 35157 8560 35191
rect 8560 35157 8594 35191
rect 8594 35157 8696 35191
rect 8696 35157 8730 35191
rect 8730 35157 8832 35191
rect 8832 35157 8866 35191
rect 8866 35157 8968 35191
rect 8968 35157 9002 35191
rect 9002 35157 9104 35191
rect 9104 35157 9138 35191
rect 9138 35157 9240 35191
rect 9240 35157 9274 35191
rect 9274 35157 9278 35191
rect 7876 35055 9278 35157
rect 7876 35021 7880 35055
rect 7880 35021 7914 35055
rect 7914 35021 8016 35055
rect 8016 35021 8050 35055
rect 8050 35021 8152 35055
rect 8152 35021 8186 35055
rect 8186 35021 8288 35055
rect 8288 35021 8322 35055
rect 8322 35021 8424 35055
rect 8424 35021 8458 35055
rect 8458 35021 8560 35055
rect 8560 35021 8594 35055
rect 8594 35021 8696 35055
rect 8696 35021 8730 35055
rect 8730 35021 8832 35055
rect 8832 35021 8866 35055
rect 8866 35021 8968 35055
rect 8968 35021 9002 35055
rect 9002 35021 9104 35055
rect 9104 35021 9138 35055
rect 9138 35021 9240 35055
rect 9240 35021 9274 35055
rect 9274 35021 9278 35055
rect 7876 34919 9278 35021
rect 7876 34885 7880 34919
rect 7880 34885 7914 34919
rect 7914 34885 8016 34919
rect 8016 34885 8050 34919
rect 8050 34885 8152 34919
rect 8152 34885 8186 34919
rect 8186 34885 8288 34919
rect 8288 34885 8322 34919
rect 8322 34885 8424 34919
rect 8424 34885 8458 34919
rect 8458 34885 8560 34919
rect 8560 34885 8594 34919
rect 8594 34885 8696 34919
rect 8696 34885 8730 34919
rect 8730 34885 8832 34919
rect 8832 34885 8866 34919
rect 8866 34885 8968 34919
rect 8968 34885 9002 34919
rect 9002 34885 9104 34919
rect 9104 34885 9138 34919
rect 9138 34885 9240 34919
rect 9240 34885 9274 34919
rect 9274 34885 9278 34919
rect 7876 34783 9278 34885
rect 7876 34749 7880 34783
rect 7880 34749 7914 34783
rect 7914 34749 8016 34783
rect 8016 34749 8050 34783
rect 8050 34749 8152 34783
rect 8152 34749 8186 34783
rect 8186 34749 8288 34783
rect 8288 34749 8322 34783
rect 8322 34749 8424 34783
rect 8424 34749 8458 34783
rect 8458 34749 8560 34783
rect 8560 34749 8594 34783
rect 8594 34749 8696 34783
rect 8696 34749 8730 34783
rect 8730 34749 8832 34783
rect 8832 34749 8866 34783
rect 8866 34749 8968 34783
rect 8968 34749 9002 34783
rect 9002 34749 9104 34783
rect 9104 34749 9138 34783
rect 9138 34749 9240 34783
rect 9240 34749 9274 34783
rect 9274 34749 9278 34783
rect 7876 34647 9278 34749
rect 7876 34613 7880 34647
rect 7880 34613 7914 34647
rect 7914 34613 8016 34647
rect 8016 34613 8050 34647
rect 8050 34613 8152 34647
rect 8152 34613 8186 34647
rect 8186 34613 8288 34647
rect 8288 34613 8322 34647
rect 8322 34613 8424 34647
rect 8424 34613 8458 34647
rect 8458 34613 8560 34647
rect 8560 34613 8594 34647
rect 8594 34613 8696 34647
rect 8696 34613 8730 34647
rect 8730 34613 8832 34647
rect 8832 34613 8866 34647
rect 8866 34613 8968 34647
rect 8968 34613 9002 34647
rect 9002 34613 9104 34647
rect 9104 34613 9138 34647
rect 9138 34613 9240 34647
rect 9240 34613 9274 34647
rect 9274 34613 9278 34647
rect 7876 34511 9278 34613
rect 7876 34477 7880 34511
rect 7880 34477 7914 34511
rect 7914 34477 8016 34511
rect 8016 34477 8050 34511
rect 8050 34477 8152 34511
rect 8152 34477 8186 34511
rect 8186 34477 8288 34511
rect 8288 34477 8322 34511
rect 8322 34477 8424 34511
rect 8424 34477 8458 34511
rect 8458 34477 8560 34511
rect 8560 34477 8594 34511
rect 8594 34477 8696 34511
rect 8696 34477 8730 34511
rect 8730 34477 8832 34511
rect 8832 34477 8866 34511
rect 8866 34477 8968 34511
rect 8968 34477 9002 34511
rect 9002 34477 9104 34511
rect 9104 34477 9138 34511
rect 9138 34477 9240 34511
rect 9240 34477 9274 34511
rect 9274 34477 9278 34511
rect 7876 34375 9278 34477
rect 7876 34341 7880 34375
rect 7880 34341 7914 34375
rect 7914 34341 8016 34375
rect 8016 34341 8050 34375
rect 8050 34341 8152 34375
rect 8152 34341 8186 34375
rect 8186 34341 8288 34375
rect 8288 34341 8322 34375
rect 8322 34341 8424 34375
rect 8424 34341 8458 34375
rect 8458 34341 8560 34375
rect 8560 34341 8594 34375
rect 8594 34341 8696 34375
rect 8696 34341 8730 34375
rect 8730 34341 8832 34375
rect 8832 34341 8866 34375
rect 8866 34341 8968 34375
rect 8968 34341 9002 34375
rect 9002 34341 9104 34375
rect 9104 34341 9138 34375
rect 9138 34341 9240 34375
rect 9240 34341 9274 34375
rect 9274 34341 9278 34375
rect 7876 34239 9278 34341
rect 7876 34205 7880 34239
rect 7880 34205 7914 34239
rect 7914 34205 8016 34239
rect 8016 34205 8050 34239
rect 8050 34205 8152 34239
rect 8152 34205 8186 34239
rect 8186 34205 8288 34239
rect 8288 34205 8322 34239
rect 8322 34205 8424 34239
rect 8424 34205 8458 34239
rect 8458 34205 8560 34239
rect 8560 34205 8594 34239
rect 8594 34205 8696 34239
rect 8696 34205 8730 34239
rect 8730 34205 8832 34239
rect 8832 34205 8866 34239
rect 8866 34205 8968 34239
rect 8968 34205 9002 34239
rect 9002 34205 9104 34239
rect 9104 34205 9138 34239
rect 9138 34205 9240 34239
rect 9240 34205 9274 34239
rect 9274 34205 9278 34239
rect 7876 34103 9278 34205
rect 7876 34069 7880 34103
rect 7880 34069 7914 34103
rect 7914 34069 8016 34103
rect 8016 34069 8050 34103
rect 8050 34069 8152 34103
rect 8152 34069 8186 34103
rect 8186 34069 8288 34103
rect 8288 34069 8322 34103
rect 8322 34069 8424 34103
rect 8424 34069 8458 34103
rect 8458 34069 8560 34103
rect 8560 34069 8594 34103
rect 8594 34069 8696 34103
rect 8696 34069 8730 34103
rect 8730 34069 8832 34103
rect 8832 34069 8866 34103
rect 8866 34069 8968 34103
rect 8968 34069 9002 34103
rect 9002 34069 9104 34103
rect 9104 34069 9138 34103
rect 9138 34069 9240 34103
rect 9240 34069 9274 34103
rect 9274 34069 9278 34103
rect 7876 33967 9278 34069
rect 7876 33933 7880 33967
rect 7880 33933 7914 33967
rect 7914 33933 8016 33967
rect 8016 33933 8050 33967
rect 8050 33933 8152 33967
rect 8152 33933 8186 33967
rect 8186 33933 8288 33967
rect 8288 33933 8322 33967
rect 8322 33933 8424 33967
rect 8424 33933 8458 33967
rect 8458 33933 8560 33967
rect 8560 33933 8594 33967
rect 8594 33933 8696 33967
rect 8696 33933 8730 33967
rect 8730 33933 8832 33967
rect 8832 33933 8866 33967
rect 8866 33933 8968 33967
rect 8968 33933 9002 33967
rect 9002 33933 9104 33967
rect 9104 33933 9138 33967
rect 9138 33933 9240 33967
rect 9240 33933 9274 33967
rect 9274 33933 9278 33967
rect 7876 33831 9278 33933
rect 7876 33797 7880 33831
rect 7880 33797 7914 33831
rect 7914 33797 8016 33831
rect 8016 33797 8050 33831
rect 8050 33797 8152 33831
rect 8152 33797 8186 33831
rect 8186 33797 8288 33831
rect 8288 33797 8322 33831
rect 8322 33797 8424 33831
rect 8424 33797 8458 33831
rect 8458 33797 8560 33831
rect 8560 33797 8594 33831
rect 8594 33797 8696 33831
rect 8696 33797 8730 33831
rect 8730 33797 8832 33831
rect 8832 33797 8866 33831
rect 8866 33797 8968 33831
rect 8968 33797 9002 33831
rect 9002 33797 9104 33831
rect 9104 33797 9138 33831
rect 9138 33797 9240 33831
rect 9240 33797 9274 33831
rect 9274 33797 9278 33831
rect 7876 33695 9278 33797
rect 7876 33661 7880 33695
rect 7880 33661 7914 33695
rect 7914 33661 8016 33695
rect 8016 33661 8050 33695
rect 8050 33661 8152 33695
rect 8152 33661 8186 33695
rect 8186 33661 8288 33695
rect 8288 33661 8322 33695
rect 8322 33661 8424 33695
rect 8424 33661 8458 33695
rect 8458 33661 8560 33695
rect 8560 33661 8594 33695
rect 8594 33661 8696 33695
rect 8696 33661 8730 33695
rect 8730 33661 8832 33695
rect 8832 33661 8866 33695
rect 8866 33661 8968 33695
rect 8968 33661 9002 33695
rect 9002 33661 9104 33695
rect 9104 33661 9138 33695
rect 9138 33661 9240 33695
rect 9240 33661 9274 33695
rect 9274 33661 9278 33695
rect 7876 33559 9278 33661
rect 7876 33525 7880 33559
rect 7880 33525 7914 33559
rect 7914 33525 8016 33559
rect 8016 33525 8050 33559
rect 8050 33525 8152 33559
rect 8152 33525 8186 33559
rect 8186 33525 8288 33559
rect 8288 33525 8322 33559
rect 8322 33525 8424 33559
rect 8424 33525 8458 33559
rect 8458 33525 8560 33559
rect 8560 33525 8594 33559
rect 8594 33525 8696 33559
rect 8696 33525 8730 33559
rect 8730 33525 8832 33559
rect 8832 33525 8866 33559
rect 8866 33525 8968 33559
rect 8968 33525 9002 33559
rect 9002 33525 9104 33559
rect 9104 33525 9138 33559
rect 9138 33525 9240 33559
rect 9240 33525 9274 33559
rect 9274 33525 9278 33559
rect 7876 33423 9278 33525
rect 7876 33389 7880 33423
rect 7880 33389 7914 33423
rect 7914 33389 8016 33423
rect 8016 33389 8050 33423
rect 8050 33389 8152 33423
rect 8152 33389 8186 33423
rect 8186 33389 8288 33423
rect 8288 33389 8322 33423
rect 8322 33389 8424 33423
rect 8424 33389 8458 33423
rect 8458 33389 8560 33423
rect 8560 33389 8594 33423
rect 8594 33389 8696 33423
rect 8696 33389 8730 33423
rect 8730 33389 8832 33423
rect 8832 33389 8866 33423
rect 8866 33389 8968 33423
rect 8968 33389 9002 33423
rect 9002 33389 9104 33423
rect 9104 33389 9138 33423
rect 9138 33389 9240 33423
rect 9240 33389 9274 33423
rect 9274 33389 9278 33423
rect 7876 33357 9278 33389
rect 7876 33287 7910 33318
rect 7876 33284 7880 33287
rect 7880 33284 7910 33287
rect 7948 33284 7982 33318
rect 8020 33287 8054 33318
rect 8020 33284 8050 33287
rect 8050 33284 8054 33287
rect 8092 33284 8126 33318
rect 8164 33287 8198 33318
rect 8164 33284 8186 33287
rect 8186 33284 8198 33287
rect 8236 33284 8270 33318
rect 8308 33287 8342 33318
rect 8308 33284 8322 33287
rect 8322 33284 8342 33287
rect 8380 33284 8414 33318
rect 8452 33287 8486 33318
rect 8452 33284 8458 33287
rect 8458 33284 8486 33287
rect 8524 33284 8558 33318
rect 8596 33284 8630 33318
rect 8668 33287 8702 33318
rect 8668 33284 8696 33287
rect 8696 33284 8702 33287
rect 8740 33284 8774 33318
rect 8812 33287 8846 33318
rect 8812 33284 8832 33287
rect 8832 33284 8846 33287
rect 8884 33284 8918 33318
rect 8956 33287 8990 33318
rect 8956 33284 8968 33287
rect 8968 33284 8990 33287
rect 9028 33284 9062 33318
rect 9100 33287 9134 33318
rect 9100 33284 9104 33287
rect 9104 33284 9134 33287
rect 9172 33284 9206 33318
rect 9244 33287 9278 33318
rect 9244 33284 9274 33287
rect 9274 33284 9278 33287
rect 7876 33211 7910 33245
rect 7948 33211 7982 33245
rect 8020 33211 8054 33245
rect 8092 33211 8126 33245
rect 8164 33211 8198 33245
rect 8236 33211 8270 33245
rect 8308 33211 8342 33245
rect 8380 33211 8414 33245
rect 8452 33211 8486 33245
rect 8524 33211 8558 33245
rect 8596 33211 8630 33245
rect 8668 33211 8702 33245
rect 8740 33211 8774 33245
rect 8812 33211 8846 33245
rect 8884 33211 8918 33245
rect 8956 33211 8990 33245
rect 9028 33211 9062 33245
rect 9100 33211 9134 33245
rect 9172 33211 9206 33245
rect 9244 33211 9278 33245
rect 7876 33151 7910 33172
rect 7876 33138 7880 33151
rect 7880 33138 7910 33151
rect 7948 33138 7982 33172
rect 8020 33151 8054 33172
rect 8020 33138 8050 33151
rect 8050 33138 8054 33151
rect 8092 33138 8126 33172
rect 8164 33151 8198 33172
rect 8164 33138 8186 33151
rect 8186 33138 8198 33151
rect 8236 33138 8270 33172
rect 8308 33151 8342 33172
rect 8308 33138 8322 33151
rect 8322 33138 8342 33151
rect 8380 33138 8414 33172
rect 8452 33151 8486 33172
rect 8452 33138 8458 33151
rect 8458 33138 8486 33151
rect 8524 33138 8558 33172
rect 8596 33138 8630 33172
rect 8668 33151 8702 33172
rect 8668 33138 8696 33151
rect 8696 33138 8702 33151
rect 8740 33138 8774 33172
rect 8812 33151 8846 33172
rect 8812 33138 8832 33151
rect 8832 33138 8846 33151
rect 8884 33138 8918 33172
rect 8956 33151 8990 33172
rect 8956 33138 8968 33151
rect 8968 33138 8990 33151
rect 9028 33138 9062 33172
rect 9100 33151 9134 33172
rect 9100 33138 9104 33151
rect 9104 33138 9134 33151
rect 9172 33138 9206 33172
rect 9244 33151 9278 33172
rect 9244 33138 9274 33151
rect 9274 33138 9278 33151
rect 7876 33065 7910 33099
rect 7948 33065 7982 33099
rect 8020 33065 8054 33099
rect 8092 33065 8126 33099
rect 8164 33065 8198 33099
rect 8236 33065 8270 33099
rect 8308 33065 8342 33099
rect 8380 33065 8414 33099
rect 8452 33065 8486 33099
rect 8524 33065 8558 33099
rect 8596 33065 8630 33099
rect 8668 33065 8702 33099
rect 8740 33065 8774 33099
rect 8812 33065 8846 33099
rect 8884 33065 8918 33099
rect 8956 33065 8990 33099
rect 9028 33065 9062 33099
rect 9100 33065 9134 33099
rect 9172 33065 9206 33099
rect 9244 33065 9278 33099
rect 7876 33015 7910 33026
rect 7876 32992 7880 33015
rect 7880 32992 7910 33015
rect 7948 32992 7982 33026
rect 8020 33015 8054 33026
rect 8020 32992 8050 33015
rect 8050 32992 8054 33015
rect 8092 32992 8126 33026
rect 8164 33015 8198 33026
rect 8164 32992 8186 33015
rect 8186 32992 8198 33015
rect 8236 32992 8270 33026
rect 8308 33015 8342 33026
rect 8308 32992 8322 33015
rect 8322 32992 8342 33015
rect 8380 32992 8414 33026
rect 8452 33015 8486 33026
rect 8452 32992 8458 33015
rect 8458 32992 8486 33015
rect 8524 32992 8558 33026
rect 8596 32992 8630 33026
rect 8668 33015 8702 33026
rect 8668 32992 8696 33015
rect 8696 32992 8702 33015
rect 8740 32992 8774 33026
rect 8812 33015 8846 33026
rect 8812 32992 8832 33015
rect 8832 32992 8846 33015
rect 8884 32992 8918 33026
rect 8956 33015 8990 33026
rect 8956 32992 8968 33015
rect 8968 32992 8990 33015
rect 9028 32992 9062 33026
rect 9100 33015 9134 33026
rect 9100 32992 9104 33015
rect 9104 32992 9134 33015
rect 9172 32992 9206 33026
rect 9244 33015 9278 33026
rect 9244 32992 9274 33015
rect 9274 32992 9278 33015
rect 7876 32919 7910 32953
rect 7948 32919 7982 32953
rect 8020 32919 8054 32953
rect 8092 32919 8126 32953
rect 8164 32919 8198 32953
rect 8236 32919 8270 32953
rect 8308 32919 8342 32953
rect 8380 32919 8414 32953
rect 8452 32919 8486 32953
rect 8524 32919 8558 32953
rect 8596 32919 8630 32953
rect 8668 32919 8702 32953
rect 8740 32919 8774 32953
rect 8812 32919 8846 32953
rect 8884 32919 8918 32953
rect 8956 32919 8990 32953
rect 9028 32919 9062 32953
rect 9100 32919 9134 32953
rect 9172 32919 9206 32953
rect 9244 32919 9278 32953
rect 7876 32879 7910 32880
rect 7876 32846 7880 32879
rect 7880 32846 7910 32879
rect 7948 32846 7982 32880
rect 8020 32879 8054 32880
rect 8020 32846 8050 32879
rect 8050 32846 8054 32879
rect 8092 32846 8126 32880
rect 8164 32879 8198 32880
rect 8164 32846 8186 32879
rect 8186 32846 8198 32879
rect 8236 32846 8270 32880
rect 8308 32879 8342 32880
rect 8308 32846 8322 32879
rect 8322 32846 8342 32879
rect 8380 32846 8414 32880
rect 8452 32879 8486 32880
rect 8452 32846 8458 32879
rect 8458 32846 8486 32879
rect 8524 32846 8558 32880
rect 8596 32846 8630 32880
rect 8668 32879 8702 32880
rect 8668 32846 8696 32879
rect 8696 32846 8702 32879
rect 8740 32846 8774 32880
rect 8812 32879 8846 32880
rect 8812 32846 8832 32879
rect 8832 32846 8846 32879
rect 8884 32846 8918 32880
rect 8956 32879 8990 32880
rect 8956 32846 8968 32879
rect 8968 32846 8990 32879
rect 9028 32846 9062 32880
rect 9100 32879 9134 32880
rect 9100 32846 9104 32879
rect 9104 32846 9134 32879
rect 9172 32846 9206 32880
rect 9244 32879 9278 32880
rect 9244 32846 9274 32879
rect 9274 32846 9278 32879
rect 7876 32773 7910 32807
rect 7948 32773 7982 32807
rect 8020 32773 8054 32807
rect 8092 32773 8126 32807
rect 8164 32773 8198 32807
rect 8236 32773 8270 32807
rect 8308 32773 8342 32807
rect 8380 32773 8414 32807
rect 8452 32773 8486 32807
rect 8524 32773 8558 32807
rect 8596 32773 8630 32807
rect 8668 32773 8702 32807
rect 8740 32773 8774 32807
rect 8812 32773 8846 32807
rect 8884 32773 8918 32807
rect 8956 32773 8990 32807
rect 9028 32773 9062 32807
rect 9100 32773 9134 32807
rect 9172 32773 9206 32807
rect 9244 32773 9278 32807
rect 7876 32709 7880 32734
rect 7880 32709 7910 32734
rect 7876 32700 7910 32709
rect 7948 32700 7982 32734
rect 8020 32709 8050 32734
rect 8050 32709 8054 32734
rect 8020 32700 8054 32709
rect 8092 32700 8126 32734
rect 8164 32709 8186 32734
rect 8186 32709 8198 32734
rect 8164 32700 8198 32709
rect 8236 32700 8270 32734
rect 8308 32709 8322 32734
rect 8322 32709 8342 32734
rect 8308 32700 8342 32709
rect 8380 32700 8414 32734
rect 8452 32709 8458 32734
rect 8458 32709 8486 32734
rect 8452 32700 8486 32709
rect 8524 32700 8558 32734
rect 8596 32700 8630 32734
rect 8668 32709 8696 32734
rect 8696 32709 8702 32734
rect 8668 32700 8702 32709
rect 8740 32700 8774 32734
rect 8812 32709 8832 32734
rect 8832 32709 8846 32734
rect 8812 32700 8846 32709
rect 8884 32700 8918 32734
rect 8956 32709 8968 32734
rect 8968 32709 8990 32734
rect 8956 32700 8990 32709
rect 9028 32700 9062 32734
rect 9100 32709 9104 32734
rect 9104 32709 9134 32734
rect 9100 32700 9134 32709
rect 9172 32700 9206 32734
rect 9244 32709 9274 32734
rect 9274 32709 9278 32734
rect 9244 32700 9278 32709
rect 7876 32627 7910 32661
rect 7948 32627 7982 32661
rect 8020 32627 8054 32661
rect 8092 32627 8126 32661
rect 8164 32627 8198 32661
rect 8236 32627 8270 32661
rect 8308 32627 8342 32661
rect 8380 32627 8414 32661
rect 8452 32627 8486 32661
rect 8524 32627 8558 32661
rect 8596 32627 8630 32661
rect 8668 32627 8702 32661
rect 8740 32627 8774 32661
rect 8812 32627 8846 32661
rect 8884 32627 8918 32661
rect 8956 32627 8990 32661
rect 9028 32627 9062 32661
rect 9100 32627 9134 32661
rect 9172 32627 9206 32661
rect 9244 32627 9278 32661
rect 7876 32573 7880 32588
rect 7880 32573 7910 32588
rect 7876 32554 7910 32573
rect 7948 32554 7982 32588
rect 8020 32573 8050 32588
rect 8050 32573 8054 32588
rect 8020 32554 8054 32573
rect 8092 32554 8126 32588
rect 8164 32573 8186 32588
rect 8186 32573 8198 32588
rect 8164 32554 8198 32573
rect 8236 32554 8270 32588
rect 8308 32573 8322 32588
rect 8322 32573 8342 32588
rect 8308 32554 8342 32573
rect 8380 32554 8414 32588
rect 8452 32573 8458 32588
rect 8458 32573 8486 32588
rect 8452 32554 8486 32573
rect 8524 32554 8558 32588
rect 8596 32554 8630 32588
rect 8668 32573 8696 32588
rect 8696 32573 8702 32588
rect 8668 32554 8702 32573
rect 8740 32554 8774 32588
rect 8812 32573 8832 32588
rect 8832 32573 8846 32588
rect 8812 32554 8846 32573
rect 8884 32554 8918 32588
rect 8956 32573 8968 32588
rect 8968 32573 8990 32588
rect 8956 32554 8990 32573
rect 9028 32554 9062 32588
rect 9100 32573 9104 32588
rect 9104 32573 9134 32588
rect 9100 32554 9134 32573
rect 9172 32554 9206 32588
rect 9244 32573 9274 32588
rect 9274 32573 9278 32588
rect 9244 32554 9278 32573
rect 7876 32481 7910 32515
rect 7948 32481 7982 32515
rect 8020 32481 8054 32515
rect 8092 32481 8126 32515
rect 8164 32481 8198 32515
rect 8236 32481 8270 32515
rect 8308 32481 8342 32515
rect 8380 32481 8414 32515
rect 8452 32481 8486 32515
rect 8524 32481 8558 32515
rect 8596 32481 8630 32515
rect 8668 32481 8702 32515
rect 8740 32481 8774 32515
rect 8812 32481 8846 32515
rect 8884 32481 8918 32515
rect 8956 32481 8990 32515
rect 9028 32481 9062 32515
rect 9100 32481 9134 32515
rect 9172 32481 9206 32515
rect 9244 32481 9278 32515
rect 7876 32437 7880 32442
rect 7880 32437 7910 32442
rect 7876 32408 7910 32437
rect 7948 32408 7982 32442
rect 8020 32437 8050 32442
rect 8050 32437 8054 32442
rect 8020 32408 8054 32437
rect 8092 32408 8126 32442
rect 8164 32437 8186 32442
rect 8186 32437 8198 32442
rect 8164 32408 8198 32437
rect 8236 32408 8270 32442
rect 8308 32437 8322 32442
rect 8322 32437 8342 32442
rect 8308 32408 8342 32437
rect 8380 32408 8414 32442
rect 8452 32437 8458 32442
rect 8458 32437 8486 32442
rect 8452 32408 8486 32437
rect 8524 32408 8558 32442
rect 8596 32408 8630 32442
rect 8668 32437 8696 32442
rect 8696 32437 8702 32442
rect 8668 32408 8702 32437
rect 8740 32408 8774 32442
rect 8812 32437 8832 32442
rect 8832 32437 8846 32442
rect 8812 32408 8846 32437
rect 8884 32408 8918 32442
rect 8956 32437 8968 32442
rect 8968 32437 8990 32442
rect 8956 32408 8990 32437
rect 9028 32408 9062 32442
rect 9100 32437 9104 32442
rect 9104 32437 9134 32442
rect 9100 32408 9134 32437
rect 9172 32408 9206 32442
rect 9244 32437 9274 32442
rect 9274 32437 9278 32442
rect 9244 32408 9278 32437
rect 7876 32335 7910 32369
rect 7948 32335 7982 32369
rect 8020 32335 8054 32369
rect 8092 32335 8126 32369
rect 8164 32335 8198 32369
rect 8236 32335 8270 32369
rect 8308 32335 8342 32369
rect 8380 32335 8414 32369
rect 8452 32335 8486 32369
rect 8524 32335 8558 32369
rect 8596 32335 8630 32369
rect 8668 32335 8702 32369
rect 8740 32335 8774 32369
rect 8812 32335 8846 32369
rect 8884 32335 8918 32369
rect 8956 32335 8990 32369
rect 9028 32335 9062 32369
rect 9100 32335 9134 32369
rect 9172 32335 9206 32369
rect 9244 32335 9278 32369
rect 7876 32262 7910 32296
rect 7948 32262 7982 32296
rect 8020 32262 8054 32296
rect 8092 32262 8126 32296
rect 8164 32262 8198 32296
rect 8236 32262 8270 32296
rect 8308 32262 8342 32296
rect 8380 32262 8414 32296
rect 8452 32262 8486 32296
rect 8524 32262 8558 32296
rect 8596 32262 8630 32296
rect 8668 32262 8702 32296
rect 8740 32262 8774 32296
rect 8812 32262 8846 32296
rect 8884 32262 8918 32296
rect 8956 32262 8990 32296
rect 9028 32262 9062 32296
rect 9100 32262 9134 32296
rect 9172 32262 9206 32296
rect 9244 32262 9278 32296
rect 7876 32199 7910 32223
rect 7876 32189 7880 32199
rect 7880 32189 7910 32199
rect 7948 32189 7982 32223
rect 8020 32199 8054 32223
rect 8020 32189 8050 32199
rect 8050 32189 8054 32199
rect 8092 32189 8126 32223
rect 8164 32199 8198 32223
rect 8164 32189 8186 32199
rect 8186 32189 8198 32199
rect 8236 32189 8270 32223
rect 8308 32199 8342 32223
rect 8308 32189 8322 32199
rect 8322 32189 8342 32199
rect 8380 32189 8414 32223
rect 8452 32199 8486 32223
rect 8452 32189 8458 32199
rect 8458 32189 8486 32199
rect 8524 32189 8558 32223
rect 8596 32189 8630 32223
rect 8668 32199 8702 32223
rect 8668 32189 8696 32199
rect 8696 32189 8702 32199
rect 8740 32189 8774 32223
rect 8812 32199 8846 32223
rect 8812 32189 8832 32199
rect 8832 32189 8846 32199
rect 8884 32189 8918 32223
rect 8956 32199 8990 32223
rect 8956 32189 8968 32199
rect 8968 32189 8990 32199
rect 9028 32189 9062 32223
rect 9100 32199 9134 32223
rect 9100 32189 9104 32199
rect 9104 32189 9134 32199
rect 9172 32189 9206 32223
rect 9244 32199 9278 32223
rect 9244 32189 9274 32199
rect 9274 32189 9278 32199
rect 7876 32116 7910 32150
rect 7948 32116 7982 32150
rect 8020 32116 8054 32150
rect 8092 32116 8126 32150
rect 8164 32116 8198 32150
rect 8236 32116 8270 32150
rect 8308 32116 8342 32150
rect 8380 32116 8414 32150
rect 8452 32116 8486 32150
rect 8524 32116 8558 32150
rect 8596 32116 8630 32150
rect 8668 32116 8702 32150
rect 8740 32116 8774 32150
rect 8812 32116 8846 32150
rect 8884 32116 8918 32150
rect 8956 32116 8990 32150
rect 9028 32116 9062 32150
rect 9100 32116 9134 32150
rect 9172 32116 9206 32150
rect 9244 32116 9278 32150
rect 7876 32063 7910 32077
rect 7876 32043 7880 32063
rect 7880 32043 7910 32063
rect 7948 32043 7982 32077
rect 8020 32063 8054 32077
rect 8020 32043 8050 32063
rect 8050 32043 8054 32063
rect 8092 32043 8126 32077
rect 8164 32063 8198 32077
rect 8164 32043 8186 32063
rect 8186 32043 8198 32063
rect 8236 32043 8270 32077
rect 8308 32063 8342 32077
rect 8308 32043 8322 32063
rect 8322 32043 8342 32063
rect 8380 32043 8414 32077
rect 8452 32063 8486 32077
rect 8452 32043 8458 32063
rect 8458 32043 8486 32063
rect 8524 32043 8558 32077
rect 8596 32043 8630 32077
rect 8668 32063 8702 32077
rect 8668 32043 8696 32063
rect 8696 32043 8702 32063
rect 8740 32043 8774 32077
rect 8812 32063 8846 32077
rect 8812 32043 8832 32063
rect 8832 32043 8846 32063
rect 8884 32043 8918 32077
rect 8956 32063 8990 32077
rect 8956 32043 8968 32063
rect 8968 32043 8990 32063
rect 9028 32043 9062 32077
rect 9100 32063 9134 32077
rect 9100 32043 9104 32063
rect 9104 32043 9134 32063
rect 9172 32043 9206 32077
rect 9244 32063 9278 32077
rect 9244 32043 9274 32063
rect 9274 32043 9278 32063
rect 7876 31970 7910 32004
rect 7948 31970 7982 32004
rect 8020 31970 8054 32004
rect 8092 31970 8126 32004
rect 8164 31970 8198 32004
rect 8236 31970 8270 32004
rect 8308 31970 8342 32004
rect 8380 31970 8414 32004
rect 8452 31970 8486 32004
rect 8524 31970 8558 32004
rect 8596 31970 8630 32004
rect 8668 31970 8702 32004
rect 8740 31970 8774 32004
rect 8812 31970 8846 32004
rect 8884 31970 8918 32004
rect 8956 31970 8990 32004
rect 9028 31970 9062 32004
rect 9100 31970 9134 32004
rect 9172 31970 9206 32004
rect 9244 31970 9278 32004
rect 7876 31927 7910 31931
rect 7876 31897 7880 31927
rect 7880 31897 7910 31927
rect 7948 31897 7982 31931
rect 8020 31927 8054 31931
rect 8020 31897 8050 31927
rect 8050 31897 8054 31927
rect 8092 31897 8126 31931
rect 8164 31927 8198 31931
rect 8164 31897 8186 31927
rect 8186 31897 8198 31927
rect 8236 31897 8270 31931
rect 8308 31927 8342 31931
rect 8308 31897 8322 31927
rect 8322 31897 8342 31927
rect 8380 31897 8414 31931
rect 8452 31927 8486 31931
rect 8452 31897 8458 31927
rect 8458 31897 8486 31927
rect 8524 31897 8558 31931
rect 8596 31897 8630 31931
rect 8668 31927 8702 31931
rect 8668 31897 8696 31927
rect 8696 31897 8702 31927
rect 8740 31897 8774 31931
rect 8812 31927 8846 31931
rect 8812 31897 8832 31927
rect 8832 31897 8846 31927
rect 8884 31897 8918 31931
rect 8956 31927 8990 31931
rect 8956 31897 8968 31927
rect 8968 31897 8990 31927
rect 9028 31897 9062 31931
rect 9100 31927 9134 31931
rect 9100 31897 9104 31927
rect 9104 31897 9134 31927
rect 9172 31897 9206 31931
rect 9244 31927 9278 31931
rect 9244 31897 9274 31927
rect 9274 31897 9278 31927
rect 7876 31824 7910 31858
rect 7948 31824 7982 31858
rect 8020 31824 8054 31858
rect 8092 31824 8126 31858
rect 8164 31824 8198 31858
rect 8236 31824 8270 31858
rect 8308 31824 8342 31858
rect 8380 31824 8414 31858
rect 8452 31824 8486 31858
rect 8524 31824 8558 31858
rect 8596 31824 8630 31858
rect 8668 31824 8702 31858
rect 8740 31824 8774 31858
rect 8812 31824 8846 31858
rect 8884 31824 8918 31858
rect 8956 31824 8990 31858
rect 9028 31824 9062 31858
rect 9100 31824 9134 31858
rect 9172 31824 9206 31858
rect 9244 31824 9278 31858
rect 7876 31757 7880 31785
rect 7880 31757 7910 31785
rect 7876 31751 7910 31757
rect 7948 31751 7982 31785
rect 8020 31757 8050 31785
rect 8050 31757 8054 31785
rect 8020 31751 8054 31757
rect 8092 31751 8126 31785
rect 8164 31757 8186 31785
rect 8186 31757 8198 31785
rect 8164 31751 8198 31757
rect 8236 31751 8270 31785
rect 8308 31757 8322 31785
rect 8322 31757 8342 31785
rect 8308 31751 8342 31757
rect 8380 31751 8414 31785
rect 8452 31757 8458 31785
rect 8458 31757 8486 31785
rect 8452 31751 8486 31757
rect 8524 31751 8558 31785
rect 8596 31751 8630 31785
rect 8668 31757 8696 31785
rect 8696 31757 8702 31785
rect 8668 31751 8702 31757
rect 8740 31751 8774 31785
rect 8812 31757 8832 31785
rect 8832 31757 8846 31785
rect 8812 31751 8846 31757
rect 8884 31751 8918 31785
rect 8956 31757 8968 31785
rect 8968 31757 8990 31785
rect 8956 31751 8990 31757
rect 9028 31751 9062 31785
rect 9100 31757 9104 31785
rect 9104 31757 9134 31785
rect 9100 31751 9134 31757
rect 9172 31751 9206 31785
rect 9244 31757 9274 31785
rect 9274 31757 9278 31785
rect 9244 31751 9278 31757
rect 7876 31678 7910 31712
rect 7948 31678 7982 31712
rect 8020 31678 8054 31712
rect 8092 31678 8126 31712
rect 8164 31678 8198 31712
rect 8236 31678 8270 31712
rect 8308 31678 8342 31712
rect 8380 31678 8414 31712
rect 8452 31678 8486 31712
rect 8524 31678 8558 31712
rect 8596 31678 8630 31712
rect 8668 31678 8702 31712
rect 8740 31678 8774 31712
rect 8812 31678 8846 31712
rect 8884 31678 8918 31712
rect 8956 31678 8990 31712
rect 9028 31678 9062 31712
rect 9100 31678 9134 31712
rect 9172 31678 9206 31712
rect 9244 31678 9278 31712
rect 7876 31621 7880 31639
rect 7880 31621 7910 31639
rect 7876 31605 7910 31621
rect 7948 31605 7982 31639
rect 8020 31621 8050 31639
rect 8050 31621 8054 31639
rect 8020 31605 8054 31621
rect 8092 31605 8126 31639
rect 8164 31621 8186 31639
rect 8186 31621 8198 31639
rect 8164 31605 8198 31621
rect 8236 31605 8270 31639
rect 8308 31621 8322 31639
rect 8322 31621 8342 31639
rect 8308 31605 8342 31621
rect 8380 31605 8414 31639
rect 8452 31621 8458 31639
rect 8458 31621 8486 31639
rect 8452 31605 8486 31621
rect 8524 31605 8558 31639
rect 8596 31605 8630 31639
rect 8668 31621 8696 31639
rect 8696 31621 8702 31639
rect 8668 31605 8702 31621
rect 8740 31605 8774 31639
rect 8812 31621 8832 31639
rect 8832 31621 8846 31639
rect 8812 31605 8846 31621
rect 8884 31605 8918 31639
rect 8956 31621 8968 31639
rect 8968 31621 8990 31639
rect 8956 31605 8990 31621
rect 9028 31605 9062 31639
rect 9100 31621 9104 31639
rect 9104 31621 9134 31639
rect 9100 31605 9134 31621
rect 9172 31605 9206 31639
rect 9244 31621 9274 31639
rect 9274 31621 9278 31639
rect 9244 31605 9278 31621
rect 7876 31532 7910 31566
rect 7948 31532 7982 31566
rect 8020 31532 8054 31566
rect 8092 31532 8126 31566
rect 8164 31532 8198 31566
rect 8236 31532 8270 31566
rect 8308 31532 8342 31566
rect 8380 31532 8414 31566
rect 8452 31532 8486 31566
rect 8524 31532 8558 31566
rect 8596 31532 8630 31566
rect 8668 31532 8702 31566
rect 8740 31532 8774 31566
rect 8812 31532 8846 31566
rect 8884 31532 8918 31566
rect 8956 31532 8990 31566
rect 9028 31532 9062 31566
rect 9100 31532 9134 31566
rect 9172 31532 9206 31566
rect 9244 31532 9278 31566
rect 7876 31485 7880 31493
rect 7880 31485 7910 31493
rect 7876 31459 7910 31485
rect 7948 31459 7982 31493
rect 8020 31485 8050 31493
rect 8050 31485 8054 31493
rect 8020 31459 8054 31485
rect 8092 31459 8126 31493
rect 8164 31485 8186 31493
rect 8186 31485 8198 31493
rect 8164 31459 8198 31485
rect 8236 31459 8270 31493
rect 8308 31485 8322 31493
rect 8322 31485 8342 31493
rect 8308 31459 8342 31485
rect 8380 31459 8414 31493
rect 8452 31485 8458 31493
rect 8458 31485 8486 31493
rect 8452 31459 8486 31485
rect 8524 31459 8558 31493
rect 8596 31459 8630 31493
rect 8668 31485 8696 31493
rect 8696 31485 8702 31493
rect 8668 31459 8702 31485
rect 8740 31459 8774 31493
rect 8812 31485 8832 31493
rect 8832 31485 8846 31493
rect 8812 31459 8846 31485
rect 8884 31459 8918 31493
rect 8956 31485 8968 31493
rect 8968 31485 8990 31493
rect 8956 31459 8990 31485
rect 9028 31459 9062 31493
rect 9100 31485 9104 31493
rect 9104 31485 9134 31493
rect 9100 31459 9134 31485
rect 9172 31459 9206 31493
rect 9244 31485 9274 31493
rect 9274 31485 9278 31493
rect 9244 31459 9278 31485
rect 7876 31386 7910 31420
rect 7948 31386 7982 31420
rect 8020 31386 8054 31420
rect 8092 31386 8126 31420
rect 8164 31386 8198 31420
rect 8236 31386 8270 31420
rect 8308 31386 8342 31420
rect 8380 31386 8414 31420
rect 8452 31386 8486 31420
rect 8524 31386 8558 31420
rect 8596 31386 8630 31420
rect 8668 31386 8702 31420
rect 8740 31386 8774 31420
rect 8812 31386 8846 31420
rect 8884 31386 8918 31420
rect 8956 31386 8990 31420
rect 9028 31386 9062 31420
rect 9100 31386 9134 31420
rect 9172 31386 9206 31420
rect 9244 31386 9278 31420
rect 7876 31313 7910 31347
rect 7948 31313 7982 31347
rect 8020 31313 8054 31347
rect 8092 31313 8126 31347
rect 8164 31313 8198 31347
rect 8236 31313 8270 31347
rect 8308 31313 8342 31347
rect 8380 31313 8414 31347
rect 8452 31313 8486 31347
rect 8524 31313 8558 31347
rect 8596 31313 8630 31347
rect 8668 31313 8702 31347
rect 8740 31313 8774 31347
rect 8812 31313 8846 31347
rect 8884 31313 8918 31347
rect 8956 31313 8990 31347
rect 9028 31313 9062 31347
rect 9100 31313 9134 31347
rect 9172 31313 9206 31347
rect 9244 31313 9278 31347
rect 7876 31247 7910 31274
rect 7876 31240 7880 31247
rect 7880 31240 7910 31247
rect 7948 31240 7982 31274
rect 8020 31247 8054 31274
rect 8020 31240 8050 31247
rect 8050 31240 8054 31247
rect 8092 31240 8126 31274
rect 8164 31247 8198 31274
rect 8164 31240 8186 31247
rect 8186 31240 8198 31247
rect 8236 31240 8270 31274
rect 8308 31247 8342 31274
rect 8308 31240 8322 31247
rect 8322 31240 8342 31247
rect 8380 31240 8414 31274
rect 8452 31247 8486 31274
rect 8452 31240 8458 31247
rect 8458 31240 8486 31247
rect 8524 31240 8558 31274
rect 8596 31240 8630 31274
rect 8668 31247 8702 31274
rect 8668 31240 8696 31247
rect 8696 31240 8702 31247
rect 8740 31240 8774 31274
rect 8812 31247 8846 31274
rect 8812 31240 8832 31247
rect 8832 31240 8846 31247
rect 8884 31240 8918 31274
rect 8956 31247 8990 31274
rect 8956 31240 8968 31247
rect 8968 31240 8990 31247
rect 9028 31240 9062 31274
rect 9100 31247 9134 31274
rect 9100 31240 9104 31247
rect 9104 31240 9134 31247
rect 9172 31240 9206 31274
rect 9244 31247 9278 31274
rect 9244 31240 9274 31247
rect 9274 31240 9278 31247
rect 7876 31167 7910 31201
rect 7948 31167 7982 31201
rect 8020 31167 8054 31201
rect 8092 31167 8126 31201
rect 8164 31167 8198 31201
rect 8236 31167 8270 31201
rect 8308 31167 8342 31201
rect 8380 31167 8414 31201
rect 8452 31167 8486 31201
rect 8524 31167 8558 31201
rect 8596 31167 8630 31201
rect 8668 31167 8702 31201
rect 8740 31167 8774 31201
rect 8812 31167 8846 31201
rect 8884 31167 8918 31201
rect 8956 31167 8990 31201
rect 9028 31167 9062 31201
rect 9100 31167 9134 31201
rect 9172 31167 9206 31201
rect 9244 31167 9278 31201
rect 7876 31111 7910 31128
rect 7876 31094 7880 31111
rect 7880 31094 7910 31111
rect 7948 31094 7982 31128
rect 8020 31111 8054 31128
rect 8020 31094 8050 31111
rect 8050 31094 8054 31111
rect 8092 31094 8126 31128
rect 8164 31111 8198 31128
rect 8164 31094 8186 31111
rect 8186 31094 8198 31111
rect 8236 31094 8270 31128
rect 8308 31111 8342 31128
rect 8308 31094 8322 31111
rect 8322 31094 8342 31111
rect 8380 31094 8414 31128
rect 8452 31111 8486 31128
rect 8452 31094 8458 31111
rect 8458 31094 8486 31111
rect 8524 31094 8558 31128
rect 8596 31094 8630 31128
rect 8668 31111 8702 31128
rect 8668 31094 8696 31111
rect 8696 31094 8702 31111
rect 8740 31094 8774 31128
rect 8812 31111 8846 31128
rect 8812 31094 8832 31111
rect 8832 31094 8846 31111
rect 8884 31094 8918 31128
rect 8956 31111 8990 31128
rect 8956 31094 8968 31111
rect 8968 31094 8990 31111
rect 9028 31094 9062 31128
rect 9100 31111 9134 31128
rect 9100 31094 9104 31111
rect 9104 31094 9134 31111
rect 9172 31094 9206 31128
rect 9244 31111 9278 31128
rect 9244 31094 9274 31111
rect 9274 31094 9278 31111
rect 7876 31021 7910 31055
rect 7948 31021 7982 31055
rect 8020 31021 8054 31055
rect 8092 31021 8126 31055
rect 8164 31021 8198 31055
rect 8236 31021 8270 31055
rect 8308 31021 8342 31055
rect 8380 31021 8414 31055
rect 8452 31021 8486 31055
rect 8524 31021 8558 31055
rect 8596 31021 8630 31055
rect 8668 31021 8702 31055
rect 8740 31021 8774 31055
rect 8812 31021 8846 31055
rect 8884 31021 8918 31055
rect 8956 31021 8990 31055
rect 9028 31021 9062 31055
rect 9100 31021 9134 31055
rect 9172 31021 9206 31055
rect 9244 31021 9278 31055
rect 7876 30975 7910 30982
rect 7876 30948 7880 30975
rect 7880 30948 7910 30975
rect 7948 30948 7982 30982
rect 8020 30975 8054 30982
rect 8020 30948 8050 30975
rect 8050 30948 8054 30975
rect 8092 30948 8126 30982
rect 8164 30975 8198 30982
rect 8164 30948 8186 30975
rect 8186 30948 8198 30975
rect 8236 30948 8270 30982
rect 8308 30975 8342 30982
rect 8308 30948 8322 30975
rect 8322 30948 8342 30975
rect 8380 30948 8414 30982
rect 8452 30975 8486 30982
rect 8452 30948 8458 30975
rect 8458 30948 8486 30975
rect 8524 30948 8558 30982
rect 8596 30948 8630 30982
rect 8668 30975 8702 30982
rect 8668 30948 8696 30975
rect 8696 30948 8702 30975
rect 8740 30948 8774 30982
rect 8812 30975 8846 30982
rect 8812 30948 8832 30975
rect 8832 30948 8846 30975
rect 8884 30948 8918 30982
rect 8956 30975 8990 30982
rect 8956 30948 8968 30975
rect 8968 30948 8990 30975
rect 9028 30948 9062 30982
rect 9100 30975 9134 30982
rect 9100 30948 9104 30975
rect 9104 30948 9134 30975
rect 9172 30948 9206 30982
rect 9244 30975 9278 30982
rect 9244 30948 9274 30975
rect 9274 30948 9278 30975
rect 7876 30875 7910 30909
rect 7948 30875 7982 30909
rect 8020 30875 8054 30909
rect 8092 30875 8126 30909
rect 8164 30875 8198 30909
rect 8236 30875 8270 30909
rect 8308 30875 8342 30909
rect 8380 30875 8414 30909
rect 8452 30875 8486 30909
rect 8524 30875 8558 30909
rect 8596 30875 8630 30909
rect 8668 30875 8702 30909
rect 8740 30875 8774 30909
rect 8812 30875 8846 30909
rect 8884 30875 8918 30909
rect 8956 30875 8990 30909
rect 9028 30875 9062 30909
rect 9100 30875 9134 30909
rect 9172 30875 9206 30909
rect 9244 30875 9278 30909
rect 7876 30805 7880 30836
rect 7880 30805 7910 30836
rect 7876 30802 7910 30805
rect 7948 30802 7982 30836
rect 8020 30805 8050 30836
rect 8050 30805 8054 30836
rect 8020 30802 8054 30805
rect 8092 30802 8126 30836
rect 8164 30805 8186 30836
rect 8186 30805 8198 30836
rect 8164 30802 8198 30805
rect 8236 30802 8270 30836
rect 8308 30805 8322 30836
rect 8322 30805 8342 30836
rect 8308 30802 8342 30805
rect 8380 30802 8414 30836
rect 8452 30805 8458 30836
rect 8458 30805 8486 30836
rect 8452 30802 8486 30805
rect 8524 30802 8558 30836
rect 8596 30802 8630 30836
rect 8668 30805 8696 30836
rect 8696 30805 8702 30836
rect 8668 30802 8702 30805
rect 8740 30802 8774 30836
rect 8812 30805 8832 30836
rect 8832 30805 8846 30836
rect 8812 30802 8846 30805
rect 8884 30802 8918 30836
rect 8956 30805 8968 30836
rect 8968 30805 8990 30836
rect 8956 30802 8990 30805
rect 9028 30802 9062 30836
rect 9100 30805 9104 30836
rect 9104 30805 9134 30836
rect 9100 30802 9134 30805
rect 9172 30802 9206 30836
rect 9244 30805 9274 30836
rect 9274 30805 9278 30836
rect 9244 30802 9278 30805
rect 7876 30729 7910 30763
rect 7948 30729 7982 30763
rect 8020 30729 8054 30763
rect 8092 30729 8126 30763
rect 8164 30729 8198 30763
rect 8236 30729 8270 30763
rect 8308 30729 8342 30763
rect 8380 30729 8414 30763
rect 8452 30729 8486 30763
rect 8524 30729 8558 30763
rect 8596 30729 8630 30763
rect 8668 30729 8702 30763
rect 8740 30729 8774 30763
rect 8812 30729 8846 30763
rect 8884 30729 8918 30763
rect 8956 30729 8990 30763
rect 9028 30729 9062 30763
rect 9100 30729 9134 30763
rect 9172 30729 9206 30763
rect 9244 30729 9278 30763
rect 7876 30669 7880 30690
rect 7880 30669 7910 30690
rect 7876 30656 7910 30669
rect 7948 30656 7982 30690
rect 8020 30669 8050 30690
rect 8050 30669 8054 30690
rect 8020 30656 8054 30669
rect 8092 30656 8126 30690
rect 8164 30669 8186 30690
rect 8186 30669 8198 30690
rect 8164 30656 8198 30669
rect 8236 30656 8270 30690
rect 8308 30669 8322 30690
rect 8322 30669 8342 30690
rect 8308 30656 8342 30669
rect 8380 30656 8414 30690
rect 8452 30669 8458 30690
rect 8458 30669 8486 30690
rect 8452 30656 8486 30669
rect 8524 30656 8558 30690
rect 8596 30656 8630 30690
rect 8668 30669 8696 30690
rect 8696 30669 8702 30690
rect 8668 30656 8702 30669
rect 8740 30656 8774 30690
rect 8812 30669 8832 30690
rect 8832 30669 8846 30690
rect 8812 30656 8846 30669
rect 8884 30656 8918 30690
rect 8956 30669 8968 30690
rect 8968 30669 8990 30690
rect 8956 30656 8990 30669
rect 9028 30656 9062 30690
rect 9100 30669 9104 30690
rect 9104 30669 9134 30690
rect 9100 30656 9134 30669
rect 9172 30656 9206 30690
rect 9244 30669 9274 30690
rect 9274 30669 9278 30690
rect 9244 30656 9278 30669
rect 7876 30583 7910 30617
rect 7948 30583 7982 30617
rect 8020 30583 8054 30617
rect 8092 30583 8126 30617
rect 8164 30583 8198 30617
rect 8236 30583 8270 30617
rect 8308 30583 8342 30617
rect 8380 30583 8414 30617
rect 8452 30583 8486 30617
rect 8524 30583 8558 30617
rect 8596 30583 8630 30617
rect 8668 30583 8702 30617
rect 8740 30583 8774 30617
rect 8812 30583 8846 30617
rect 8884 30583 8918 30617
rect 8956 30583 8990 30617
rect 9028 30583 9062 30617
rect 9100 30583 9134 30617
rect 9172 30583 9206 30617
rect 9244 30583 9278 30617
rect 7876 30533 7880 30544
rect 7880 30533 7910 30544
rect 7876 30510 7910 30533
rect 7948 30510 7982 30544
rect 8020 30533 8050 30544
rect 8050 30533 8054 30544
rect 8020 30510 8054 30533
rect 8092 30510 8126 30544
rect 8164 30533 8186 30544
rect 8186 30533 8198 30544
rect 8164 30510 8198 30533
rect 8236 30510 8270 30544
rect 8308 30533 8322 30544
rect 8322 30533 8342 30544
rect 8308 30510 8342 30533
rect 8380 30510 8414 30544
rect 8452 30533 8458 30544
rect 8458 30533 8486 30544
rect 8452 30510 8486 30533
rect 8524 30510 8558 30544
rect 8596 30510 8630 30544
rect 8668 30533 8696 30544
rect 8696 30533 8702 30544
rect 8668 30510 8702 30533
rect 8740 30510 8774 30544
rect 8812 30533 8832 30544
rect 8832 30533 8846 30544
rect 8812 30510 8846 30533
rect 8884 30510 8918 30544
rect 8956 30533 8968 30544
rect 8968 30533 8990 30544
rect 8956 30510 8990 30533
rect 9028 30510 9062 30544
rect 9100 30533 9104 30544
rect 9104 30533 9134 30544
rect 9100 30510 9134 30533
rect 9172 30510 9206 30544
rect 9244 30533 9274 30544
rect 9274 30533 9278 30544
rect 9244 30510 9278 30533
rect 7876 30437 7910 30471
rect 7948 30437 7982 30471
rect 8020 30437 8054 30471
rect 8092 30437 8126 30471
rect 8164 30437 8198 30471
rect 8236 30437 8270 30471
rect 8308 30437 8342 30471
rect 8380 30437 8414 30471
rect 8452 30437 8486 30471
rect 8524 30437 8558 30471
rect 8596 30437 8630 30471
rect 8668 30437 8702 30471
rect 8740 30437 8774 30471
rect 8812 30437 8846 30471
rect 8884 30437 8918 30471
rect 8956 30437 8990 30471
rect 9028 30437 9062 30471
rect 9100 30437 9134 30471
rect 9172 30437 9206 30471
rect 9244 30437 9278 30471
rect 7876 30397 7880 30398
rect 7880 30397 7910 30398
rect 7876 30364 7910 30397
rect 7948 30364 7982 30398
rect 8020 30397 8050 30398
rect 8050 30397 8054 30398
rect 8020 30364 8054 30397
rect 8092 30364 8126 30398
rect 8164 30397 8186 30398
rect 8186 30397 8198 30398
rect 8164 30364 8198 30397
rect 8236 30364 8270 30398
rect 8308 30397 8322 30398
rect 8322 30397 8342 30398
rect 8308 30364 8342 30397
rect 8380 30364 8414 30398
rect 8452 30397 8458 30398
rect 8458 30397 8486 30398
rect 8452 30364 8486 30397
rect 8524 30364 8558 30398
rect 8596 30364 8630 30398
rect 8668 30397 8696 30398
rect 8696 30397 8702 30398
rect 8668 30364 8702 30397
rect 8740 30364 8774 30398
rect 8812 30397 8832 30398
rect 8832 30397 8846 30398
rect 8812 30364 8846 30397
rect 8884 30364 8918 30398
rect 8956 30397 8968 30398
rect 8968 30397 8990 30398
rect 8956 30364 8990 30397
rect 9028 30364 9062 30398
rect 9100 30397 9104 30398
rect 9104 30397 9134 30398
rect 9100 30364 9134 30397
rect 9172 30364 9206 30398
rect 9244 30397 9274 30398
rect 9274 30397 9278 30398
rect 9244 30364 9278 30397
rect 7876 30295 7910 30325
rect 7876 30291 7880 30295
rect 7880 30291 7910 30295
rect 7948 30291 7982 30325
rect 8020 30295 8054 30325
rect 8020 30291 8050 30295
rect 8050 30291 8054 30295
rect 8092 30291 8126 30325
rect 8164 30295 8198 30325
rect 8164 30291 8186 30295
rect 8186 30291 8198 30295
rect 8236 30291 8270 30325
rect 8308 30295 8342 30325
rect 8308 30291 8322 30295
rect 8322 30291 8342 30295
rect 8380 30291 8414 30325
rect 8452 30295 8486 30325
rect 8452 30291 8458 30295
rect 8458 30291 8486 30295
rect 8524 30291 8558 30325
rect 8596 30291 8630 30325
rect 8668 30295 8702 30325
rect 8668 30291 8696 30295
rect 8696 30291 8702 30295
rect 8740 30291 8774 30325
rect 8812 30295 8846 30325
rect 8812 30291 8832 30295
rect 8832 30291 8846 30295
rect 8884 30291 8918 30325
rect 8956 30295 8990 30325
rect 8956 30291 8968 30295
rect 8968 30291 8990 30295
rect 9028 30291 9062 30325
rect 9100 30295 9134 30325
rect 9100 30291 9104 30295
rect 9104 30291 9134 30295
rect 9172 30291 9206 30325
rect 9244 30295 9278 30325
rect 9244 30291 9274 30295
rect 9274 30291 9278 30295
rect 7876 30218 7910 30252
rect 7948 30218 7982 30252
rect 8020 30218 8054 30252
rect 8092 30218 8126 30252
rect 8164 30218 8198 30252
rect 8236 30218 8270 30252
rect 8308 30218 8342 30252
rect 8380 30218 8414 30252
rect 8452 30218 8486 30252
rect 8524 30218 8558 30252
rect 8596 30218 8630 30252
rect 8668 30218 8702 30252
rect 8740 30218 8774 30252
rect 8812 30218 8846 30252
rect 8884 30218 8918 30252
rect 8956 30218 8990 30252
rect 9028 30218 9062 30252
rect 9100 30218 9134 30252
rect 9172 30218 9206 30252
rect 9244 30218 9278 30252
rect 7876 30159 7910 30179
rect 7876 30145 7880 30159
rect 7880 30145 7910 30159
rect 7948 30145 7982 30179
rect 8020 30159 8054 30179
rect 8020 30145 8050 30159
rect 8050 30145 8054 30159
rect 8092 30145 8126 30179
rect 8164 30159 8198 30179
rect 8164 30145 8186 30159
rect 8186 30145 8198 30159
rect 8236 30145 8270 30179
rect 8308 30159 8342 30179
rect 8308 30145 8322 30159
rect 8322 30145 8342 30159
rect 8380 30145 8414 30179
rect 8452 30159 8486 30179
rect 8452 30145 8458 30159
rect 8458 30145 8486 30159
rect 8524 30145 8558 30179
rect 8596 30145 8630 30179
rect 8668 30159 8702 30179
rect 8668 30145 8696 30159
rect 8696 30145 8702 30159
rect 8740 30145 8774 30179
rect 8812 30159 8846 30179
rect 8812 30145 8832 30159
rect 8832 30145 8846 30159
rect 8884 30145 8918 30179
rect 8956 30159 8990 30179
rect 8956 30145 8968 30159
rect 8968 30145 8990 30159
rect 9028 30145 9062 30179
rect 9100 30159 9134 30179
rect 9100 30145 9104 30159
rect 9104 30145 9134 30159
rect 9172 30145 9206 30179
rect 9244 30159 9278 30179
rect 9244 30145 9274 30159
rect 9274 30145 9278 30159
rect 7876 30072 7910 30106
rect 7948 30072 7982 30106
rect 8020 30072 8054 30106
rect 8092 30072 8126 30106
rect 8164 30072 8198 30106
rect 8236 30072 8270 30106
rect 8308 30072 8342 30106
rect 8380 30072 8414 30106
rect 8452 30072 8486 30106
rect 8524 30072 8558 30106
rect 8596 30072 8630 30106
rect 8668 30072 8702 30106
rect 8740 30072 8774 30106
rect 8812 30072 8846 30106
rect 8884 30072 8918 30106
rect 8956 30072 8990 30106
rect 9028 30072 9062 30106
rect 9100 30072 9134 30106
rect 9172 30072 9206 30106
rect 9244 30072 9278 30106
rect 7876 30023 7910 30033
rect 7876 29999 7880 30023
rect 7880 29999 7910 30023
rect 7948 29999 7982 30033
rect 8020 30023 8054 30033
rect 8020 29999 8050 30023
rect 8050 29999 8054 30023
rect 8092 29999 8126 30033
rect 8164 30023 8198 30033
rect 8164 29999 8186 30023
rect 8186 29999 8198 30023
rect 8236 29999 8270 30033
rect 8308 30023 8342 30033
rect 8308 29999 8322 30023
rect 8322 29999 8342 30023
rect 8380 29999 8414 30033
rect 8452 30023 8486 30033
rect 8452 29999 8458 30023
rect 8458 29999 8486 30023
rect 8524 29999 8558 30033
rect 8596 29999 8630 30033
rect 8668 30023 8702 30033
rect 8668 29999 8696 30023
rect 8696 29999 8702 30023
rect 8740 29999 8774 30033
rect 8812 30023 8846 30033
rect 8812 29999 8832 30023
rect 8832 29999 8846 30023
rect 8884 29999 8918 30033
rect 8956 30023 8990 30033
rect 8956 29999 8968 30023
rect 8968 29999 8990 30023
rect 9028 29999 9062 30033
rect 9100 30023 9134 30033
rect 9100 29999 9104 30023
rect 9104 29999 9134 30023
rect 9172 29999 9206 30033
rect 9244 30023 9278 30033
rect 9244 29999 9274 30023
rect 9274 29999 9278 30023
rect 7876 29926 7910 29960
rect 7948 29926 7982 29960
rect 8020 29926 8054 29960
rect 8092 29926 8126 29960
rect 8164 29926 8198 29960
rect 8236 29926 8270 29960
rect 8308 29926 8342 29960
rect 8380 29926 8414 29960
rect 8452 29926 8486 29960
rect 8524 29926 8558 29960
rect 8596 29926 8630 29960
rect 8668 29926 8702 29960
rect 8740 29926 8774 29960
rect 8812 29926 8846 29960
rect 8884 29926 8918 29960
rect 8956 29926 8990 29960
rect 9028 29926 9062 29960
rect 9100 29926 9134 29960
rect 9172 29926 9206 29960
rect 9244 29926 9278 29960
rect 7876 29853 7880 29887
rect 7880 29853 7910 29887
rect 7948 29853 7982 29887
rect 8020 29853 8050 29887
rect 8050 29853 8054 29887
rect 8092 29853 8126 29887
rect 8164 29853 8186 29887
rect 8186 29853 8198 29887
rect 8236 29853 8270 29887
rect 8308 29853 8322 29887
rect 8322 29853 8342 29887
rect 8380 29853 8414 29887
rect 8452 29853 8458 29887
rect 8458 29853 8486 29887
rect 8524 29853 8558 29887
rect 8596 29853 8630 29887
rect 8668 29853 8696 29887
rect 8696 29853 8702 29887
rect 8740 29853 8774 29887
rect 8812 29853 8832 29887
rect 8832 29853 8846 29887
rect 8884 29853 8918 29887
rect 8956 29853 8968 29887
rect 8968 29853 8990 29887
rect 9028 29853 9062 29887
rect 9100 29853 9104 29887
rect 9104 29853 9134 29887
rect 9172 29853 9206 29887
rect 9244 29853 9274 29887
rect 9274 29853 9278 29887
rect 7876 29780 7910 29814
rect 7948 29780 7982 29814
rect 8020 29780 8054 29814
rect 8092 29780 8126 29814
rect 8164 29780 8198 29814
rect 8236 29780 8270 29814
rect 8308 29780 8342 29814
rect 8380 29780 8414 29814
rect 8452 29780 8486 29814
rect 8524 29780 8558 29814
rect 8596 29780 8630 29814
rect 8668 29780 8702 29814
rect 8740 29780 8774 29814
rect 8812 29780 8846 29814
rect 8884 29780 8918 29814
rect 8956 29780 8990 29814
rect 9028 29780 9062 29814
rect 9100 29780 9134 29814
rect 9172 29780 9206 29814
rect 9244 29780 9278 29814
rect 7876 29717 7880 29741
rect 7880 29717 7910 29741
rect 7876 29707 7910 29717
rect 7948 29707 7982 29741
rect 8020 29717 8050 29741
rect 8050 29717 8054 29741
rect 8020 29707 8054 29717
rect 8092 29707 8126 29741
rect 8164 29717 8186 29741
rect 8186 29717 8198 29741
rect 8164 29707 8198 29717
rect 8236 29707 8270 29741
rect 8308 29717 8322 29741
rect 8322 29717 8342 29741
rect 8308 29707 8342 29717
rect 8380 29707 8414 29741
rect 8452 29717 8458 29741
rect 8458 29717 8486 29741
rect 8452 29707 8486 29717
rect 8524 29707 8558 29741
rect 8596 29707 8630 29741
rect 8668 29717 8696 29741
rect 8696 29717 8702 29741
rect 8668 29707 8702 29717
rect 8740 29707 8774 29741
rect 8812 29717 8832 29741
rect 8832 29717 8846 29741
rect 8812 29707 8846 29717
rect 8884 29707 8918 29741
rect 8956 29717 8968 29741
rect 8968 29717 8990 29741
rect 8956 29707 8990 29717
rect 9028 29707 9062 29741
rect 9100 29717 9104 29741
rect 9104 29717 9134 29741
rect 9100 29707 9134 29717
rect 9172 29707 9206 29741
rect 9244 29717 9274 29741
rect 9274 29717 9278 29741
rect 9244 29707 9278 29717
rect 7876 29634 7910 29668
rect 7948 29634 7982 29668
rect 8020 29634 8054 29668
rect 8092 29634 8126 29668
rect 8164 29634 8198 29668
rect 8236 29634 8270 29668
rect 8308 29634 8342 29668
rect 8380 29634 8414 29668
rect 8452 29634 8486 29668
rect 8524 29634 8558 29668
rect 8596 29634 8630 29668
rect 8668 29634 8702 29668
rect 8740 29634 8774 29668
rect 8812 29634 8846 29668
rect 8884 29634 8918 29668
rect 8956 29634 8990 29668
rect 9028 29634 9062 29668
rect 9100 29634 9134 29668
rect 9172 29634 9206 29668
rect 9244 29634 9278 29668
rect 321 29479 1003 29511
rect 321 29445 325 29479
rect 325 29445 359 29479
rect 359 29445 461 29479
rect 461 29445 495 29479
rect 495 29445 597 29479
rect 597 29445 631 29479
rect 631 29445 733 29479
rect 733 29445 767 29479
rect 767 29445 869 29479
rect 869 29445 903 29479
rect 903 29445 1003 29479
rect 321 29343 1003 29445
rect 321 29309 325 29343
rect 325 29309 359 29343
rect 359 29309 461 29343
rect 461 29309 495 29343
rect 495 29309 597 29343
rect 597 29309 631 29343
rect 631 29309 733 29343
rect 733 29309 767 29343
rect 767 29309 869 29343
rect 869 29309 903 29343
rect 903 29309 1003 29343
rect 321 29207 1003 29309
rect 321 29173 325 29207
rect 325 29173 359 29207
rect 359 29173 461 29207
rect 461 29173 495 29207
rect 495 29173 597 29207
rect 597 29173 631 29207
rect 631 29173 733 29207
rect 733 29173 767 29207
rect 767 29173 869 29207
rect 869 29173 903 29207
rect 903 29173 1003 29207
rect 321 29071 1003 29173
rect 321 29037 325 29071
rect 325 29037 359 29071
rect 359 29037 461 29071
rect 461 29037 495 29071
rect 495 29037 597 29071
rect 597 29037 631 29071
rect 631 29037 733 29071
rect 733 29037 767 29071
rect 767 29037 869 29071
rect 869 29037 903 29071
rect 903 29037 1003 29071
rect 321 28935 1003 29037
rect 321 28901 325 28935
rect 325 28901 359 28935
rect 359 28901 461 28935
rect 461 28901 495 28935
rect 495 28901 597 28935
rect 597 28901 631 28935
rect 631 28901 733 28935
rect 733 28901 767 28935
rect 767 28901 869 28935
rect 869 28901 903 28935
rect 903 28901 1003 28935
rect 321 28799 1003 28901
rect 321 28765 325 28799
rect 325 28765 359 28799
rect 359 28765 461 28799
rect 461 28765 495 28799
rect 495 28765 597 28799
rect 597 28765 631 28799
rect 631 28765 733 28799
rect 733 28765 767 28799
rect 767 28765 869 28799
rect 869 28765 903 28799
rect 903 28765 1003 28799
rect 321 28663 1003 28765
rect 321 28629 325 28663
rect 325 28629 359 28663
rect 359 28629 461 28663
rect 461 28629 495 28663
rect 495 28629 597 28663
rect 597 28629 631 28663
rect 631 28629 733 28663
rect 733 28629 767 28663
rect 767 28629 869 28663
rect 869 28629 903 28663
rect 903 28629 1003 28663
rect 321 28527 1003 28629
rect 321 28493 325 28527
rect 325 28493 359 28527
rect 359 28493 461 28527
rect 461 28493 495 28527
rect 495 28493 597 28527
rect 597 28493 631 28527
rect 631 28493 733 28527
rect 733 28493 767 28527
rect 767 28493 869 28527
rect 869 28493 903 28527
rect 903 28493 1003 28527
rect 321 28391 1003 28493
rect 321 28357 325 28391
rect 325 28357 359 28391
rect 359 28357 461 28391
rect 461 28357 495 28391
rect 495 28357 597 28391
rect 597 28357 631 28391
rect 631 28357 733 28391
rect 733 28357 767 28391
rect 767 28357 869 28391
rect 869 28357 903 28391
rect 903 28357 1003 28391
rect 321 28255 1003 28357
rect 321 28221 325 28255
rect 325 28221 359 28255
rect 359 28221 461 28255
rect 461 28221 495 28255
rect 495 28221 597 28255
rect 597 28221 631 28255
rect 631 28221 733 28255
rect 733 28221 767 28255
rect 767 28221 869 28255
rect 869 28221 903 28255
rect 903 28221 1003 28255
rect 321 28119 1003 28221
rect 321 28085 325 28119
rect 325 28085 359 28119
rect 359 28085 461 28119
rect 461 28085 495 28119
rect 495 28085 597 28119
rect 597 28085 631 28119
rect 631 28085 733 28119
rect 733 28085 767 28119
rect 767 28085 869 28119
rect 869 28085 903 28119
rect 903 28085 1003 28119
rect 321 27983 1003 28085
rect 321 27949 325 27983
rect 325 27949 359 27983
rect 359 27949 461 27983
rect 461 27949 495 27983
rect 495 27949 597 27983
rect 597 27949 631 27983
rect 631 27949 733 27983
rect 733 27949 767 27983
rect 767 27949 869 27983
rect 869 27949 903 27983
rect 903 27949 1003 27983
rect 321 27847 1003 27949
rect 321 27813 325 27847
rect 325 27813 359 27847
rect 359 27813 461 27847
rect 461 27813 495 27847
rect 495 27813 597 27847
rect 597 27813 631 27847
rect 631 27813 733 27847
rect 733 27813 767 27847
rect 767 27813 869 27847
rect 869 27813 903 27847
rect 903 27813 1003 27847
rect 321 27711 1003 27813
rect 321 27677 325 27711
rect 325 27677 359 27711
rect 359 27677 461 27711
rect 461 27677 495 27711
rect 495 27677 597 27711
rect 597 27677 631 27711
rect 631 27677 733 27711
rect 733 27677 767 27711
rect 767 27677 869 27711
rect 869 27677 903 27711
rect 903 27677 1003 27711
rect 321 27575 1003 27677
rect 321 27541 325 27575
rect 325 27541 359 27575
rect 359 27541 461 27575
rect 461 27541 495 27575
rect 495 27541 597 27575
rect 597 27541 631 27575
rect 631 27541 733 27575
rect 733 27541 767 27575
rect 767 27541 869 27575
rect 869 27541 903 27575
rect 903 27541 1003 27575
rect 321 27439 1003 27541
rect 321 27405 325 27439
rect 325 27405 359 27439
rect 359 27405 461 27439
rect 461 27405 495 27439
rect 495 27405 597 27439
rect 597 27405 631 27439
rect 631 27405 733 27439
rect 733 27405 767 27439
rect 767 27405 869 27439
rect 869 27405 903 27439
rect 903 27405 1003 27439
rect 321 27303 1003 27405
rect 321 27269 325 27303
rect 325 27269 359 27303
rect 359 27269 461 27303
rect 461 27269 495 27303
rect 495 27269 597 27303
rect 597 27269 631 27303
rect 631 27269 733 27303
rect 733 27269 767 27303
rect 767 27269 869 27303
rect 869 27269 903 27303
rect 903 27269 1003 27303
rect 321 27167 1003 27269
rect 321 27133 325 27167
rect 325 27133 359 27167
rect 359 27133 461 27167
rect 461 27133 495 27167
rect 495 27133 597 27167
rect 597 27133 631 27167
rect 631 27133 733 27167
rect 733 27133 767 27167
rect 767 27133 869 27167
rect 869 27133 903 27167
rect 903 27133 1003 27167
rect 321 27031 1003 27133
rect 321 26997 325 27031
rect 325 26997 359 27031
rect 359 26997 461 27031
rect 461 26997 495 27031
rect 495 26997 597 27031
rect 597 26997 631 27031
rect 631 26997 733 27031
rect 733 26997 767 27031
rect 767 26997 869 27031
rect 869 26997 903 27031
rect 903 26997 1003 27031
rect 321 26895 1003 26997
rect 321 26861 325 26895
rect 325 26861 359 26895
rect 359 26861 461 26895
rect 461 26861 495 26895
rect 495 26861 597 26895
rect 597 26861 631 26895
rect 631 26861 733 26895
rect 733 26861 767 26895
rect 767 26861 869 26895
rect 869 26861 903 26895
rect 903 26861 1003 26895
rect 321 26759 1003 26861
rect 321 26725 325 26759
rect 325 26725 359 26759
rect 359 26725 461 26759
rect 461 26725 495 26759
rect 495 26725 597 26759
rect 597 26725 631 26759
rect 631 26725 733 26759
rect 733 26725 767 26759
rect 767 26725 869 26759
rect 869 26725 903 26759
rect 903 26725 1003 26759
rect 321 26623 1003 26725
rect 321 26589 325 26623
rect 325 26589 359 26623
rect 359 26589 461 26623
rect 461 26589 495 26623
rect 495 26589 597 26623
rect 597 26589 631 26623
rect 631 26589 733 26623
rect 733 26589 767 26623
rect 767 26589 869 26623
rect 869 26589 903 26623
rect 903 26589 1003 26623
rect 321 26487 1003 26589
rect 321 26453 325 26487
rect 325 26453 359 26487
rect 359 26453 461 26487
rect 461 26453 495 26487
rect 495 26453 597 26487
rect 597 26453 631 26487
rect 631 26453 733 26487
rect 733 26453 767 26487
rect 767 26453 869 26487
rect 869 26453 903 26487
rect 903 26453 1003 26487
rect 321 26351 1003 26453
rect 321 26317 325 26351
rect 325 26317 359 26351
rect 359 26317 461 26351
rect 461 26317 495 26351
rect 495 26317 597 26351
rect 597 26317 631 26351
rect 631 26317 733 26351
rect 733 26317 767 26351
rect 767 26317 869 26351
rect 869 26317 903 26351
rect 903 26317 1003 26351
rect 321 26215 1003 26317
rect 321 26181 325 26215
rect 325 26181 359 26215
rect 359 26181 461 26215
rect 461 26181 495 26215
rect 495 26181 597 26215
rect 597 26181 631 26215
rect 631 26181 733 26215
rect 733 26181 767 26215
rect 767 26181 869 26215
rect 869 26181 903 26215
rect 903 26181 1003 26215
rect 321 26079 1003 26181
rect 321 26045 325 26079
rect 325 26045 359 26079
rect 359 26045 461 26079
rect 461 26045 495 26079
rect 495 26045 597 26079
rect 597 26045 631 26079
rect 631 26045 733 26079
rect 733 26045 767 26079
rect 767 26045 869 26079
rect 869 26045 903 26079
rect 903 26045 1003 26079
rect 321 25943 1003 26045
rect 321 25909 325 25943
rect 325 25909 359 25943
rect 359 25909 461 25943
rect 461 25909 495 25943
rect 495 25909 597 25943
rect 597 25909 631 25943
rect 631 25909 733 25943
rect 733 25909 767 25943
rect 767 25909 869 25943
rect 869 25909 903 25943
rect 903 25909 1003 25943
rect 321 25807 1003 25909
rect 321 25773 325 25807
rect 325 25773 359 25807
rect 359 25773 461 25807
rect 461 25773 495 25807
rect 495 25773 597 25807
rect 597 25773 631 25807
rect 631 25773 733 25807
rect 733 25773 767 25807
rect 767 25773 869 25807
rect 869 25773 903 25807
rect 903 25773 1003 25807
rect 321 25671 1003 25773
rect 321 25637 325 25671
rect 325 25637 359 25671
rect 359 25637 461 25671
rect 461 25637 495 25671
rect 495 25637 597 25671
rect 597 25637 631 25671
rect 631 25637 733 25671
rect 733 25637 767 25671
rect 767 25637 869 25671
rect 869 25637 903 25671
rect 903 25637 1003 25671
rect 321 25535 1003 25637
rect 321 25501 325 25535
rect 325 25501 359 25535
rect 359 25501 461 25535
rect 461 25501 495 25535
rect 495 25501 597 25535
rect 597 25501 631 25535
rect 631 25501 733 25535
rect 733 25501 767 25535
rect 767 25501 869 25535
rect 869 25501 903 25535
rect 903 25501 1003 25535
rect 321 25399 1003 25501
rect 321 25365 325 25399
rect 325 25365 359 25399
rect 359 25365 461 25399
rect 461 25365 495 25399
rect 495 25365 597 25399
rect 597 25365 631 25399
rect 631 25365 733 25399
rect 733 25365 767 25399
rect 767 25365 869 25399
rect 869 25365 903 25399
rect 903 25365 1003 25399
rect 321 25263 1003 25365
rect 321 25229 325 25263
rect 325 25229 359 25263
rect 359 25229 461 25263
rect 461 25229 495 25263
rect 495 25229 597 25263
rect 597 25229 631 25263
rect 631 25229 733 25263
rect 733 25229 767 25263
rect 767 25229 869 25263
rect 869 25229 903 25263
rect 903 25229 1003 25263
rect 321 25127 1003 25229
rect 321 25093 325 25127
rect 325 25093 359 25127
rect 359 25093 461 25127
rect 461 25093 495 25127
rect 495 25093 597 25127
rect 597 25093 631 25127
rect 631 25093 733 25127
rect 733 25093 767 25127
rect 767 25093 869 25127
rect 869 25093 903 25127
rect 903 25093 1003 25127
rect 321 24991 1003 25093
rect 321 24957 325 24991
rect 325 24957 359 24991
rect 359 24957 461 24991
rect 461 24957 495 24991
rect 495 24957 597 24991
rect 597 24957 631 24991
rect 631 24957 733 24991
rect 733 24957 767 24991
rect 767 24957 869 24991
rect 869 24957 903 24991
rect 903 24957 1003 24991
rect 321 24855 1003 24957
rect 321 24821 325 24855
rect 325 24821 359 24855
rect 359 24821 461 24855
rect 461 24821 495 24855
rect 495 24821 597 24855
rect 597 24821 631 24855
rect 631 24821 733 24855
rect 733 24821 767 24855
rect 767 24821 869 24855
rect 869 24821 903 24855
rect 903 24821 1003 24855
rect 321 24719 1003 24821
rect 321 24685 325 24719
rect 325 24685 359 24719
rect 359 24685 461 24719
rect 461 24685 495 24719
rect 495 24685 597 24719
rect 597 24685 631 24719
rect 631 24685 733 24719
rect 733 24685 767 24719
rect 767 24685 869 24719
rect 869 24685 903 24719
rect 903 24685 1003 24719
rect 321 24583 1003 24685
rect 321 24549 325 24583
rect 325 24549 359 24583
rect 359 24549 461 24583
rect 461 24549 495 24583
rect 495 24549 597 24583
rect 597 24549 631 24583
rect 631 24549 733 24583
rect 733 24549 767 24583
rect 767 24549 869 24583
rect 869 24549 903 24583
rect 903 24549 1003 24583
rect 321 24447 1003 24549
rect 321 24413 325 24447
rect 325 24413 359 24447
rect 359 24413 461 24447
rect 461 24413 495 24447
rect 495 24413 597 24447
rect 597 24413 631 24447
rect 631 24413 733 24447
rect 733 24413 767 24447
rect 767 24413 869 24447
rect 869 24413 903 24447
rect 903 24413 1003 24447
rect 321 24311 1003 24413
rect 321 24277 325 24311
rect 325 24277 359 24311
rect 359 24277 461 24311
rect 461 24277 495 24311
rect 495 24277 597 24311
rect 597 24277 631 24311
rect 631 24277 733 24311
rect 733 24277 767 24311
rect 767 24277 869 24311
rect 869 24277 903 24311
rect 903 24277 1003 24311
rect 321 24175 1003 24277
rect 321 24141 325 24175
rect 325 24141 359 24175
rect 359 24141 461 24175
rect 461 24141 495 24175
rect 495 24141 597 24175
rect 597 24141 631 24175
rect 631 24141 733 24175
rect 733 24141 767 24175
rect 767 24141 869 24175
rect 869 24141 903 24175
rect 903 24141 1003 24175
rect 321 24039 1003 24141
rect 321 24005 325 24039
rect 325 24005 359 24039
rect 359 24005 461 24039
rect 461 24005 495 24039
rect 495 24005 597 24039
rect 597 24005 631 24039
rect 631 24005 733 24039
rect 733 24005 767 24039
rect 767 24005 869 24039
rect 869 24005 903 24039
rect 903 24005 1003 24039
rect 321 23903 1003 24005
rect 321 23869 325 23903
rect 325 23869 359 23903
rect 359 23869 461 23903
rect 461 23869 495 23903
rect 495 23869 597 23903
rect 597 23869 631 23903
rect 631 23869 733 23903
rect 733 23869 767 23903
rect 767 23869 869 23903
rect 869 23869 903 23903
rect 903 23869 1003 23903
rect 321 23767 1003 23869
rect 321 23733 325 23767
rect 325 23733 359 23767
rect 359 23733 461 23767
rect 461 23733 495 23767
rect 495 23733 597 23767
rect 597 23733 631 23767
rect 631 23733 733 23767
rect 733 23733 767 23767
rect 767 23733 869 23767
rect 869 23733 903 23767
rect 903 23733 1003 23767
rect 321 23631 1003 23733
rect 321 23597 325 23631
rect 325 23597 359 23631
rect 359 23597 461 23631
rect 461 23597 495 23631
rect 495 23597 597 23631
rect 597 23597 631 23631
rect 631 23597 733 23631
rect 733 23597 767 23631
rect 767 23597 869 23631
rect 869 23597 903 23631
rect 903 23597 1003 23631
rect 321 23495 1003 23597
rect 321 23461 325 23495
rect 325 23461 359 23495
rect 359 23461 461 23495
rect 461 23461 495 23495
rect 495 23461 597 23495
rect 597 23461 631 23495
rect 631 23461 733 23495
rect 733 23461 767 23495
rect 767 23461 869 23495
rect 869 23461 903 23495
rect 903 23461 1003 23495
rect 321 23359 1003 23461
rect 321 23325 325 23359
rect 325 23325 359 23359
rect 359 23325 461 23359
rect 461 23325 495 23359
rect 495 23325 597 23359
rect 597 23325 631 23359
rect 631 23325 733 23359
rect 733 23325 767 23359
rect 767 23325 869 23359
rect 869 23325 903 23359
rect 903 23325 1003 23359
rect 321 23223 1003 23325
rect 321 23189 325 23223
rect 325 23189 359 23223
rect 359 23189 461 23223
rect 461 23189 495 23223
rect 495 23189 597 23223
rect 597 23189 631 23223
rect 631 23189 733 23223
rect 733 23189 767 23223
rect 767 23189 869 23223
rect 869 23189 903 23223
rect 903 23189 1003 23223
rect 321 23087 1003 23189
rect 321 23053 325 23087
rect 325 23053 359 23087
rect 359 23053 461 23087
rect 461 23053 495 23087
rect 495 23053 597 23087
rect 597 23053 631 23087
rect 631 23053 733 23087
rect 733 23053 767 23087
rect 767 23053 869 23087
rect 869 23053 903 23087
rect 903 23053 1003 23087
rect 321 22951 1003 23053
rect 321 22917 325 22951
rect 325 22917 359 22951
rect 359 22917 461 22951
rect 461 22917 495 22951
rect 495 22917 597 22951
rect 597 22917 631 22951
rect 631 22917 733 22951
rect 733 22917 767 22951
rect 767 22917 869 22951
rect 869 22917 903 22951
rect 903 22917 1003 22951
rect 321 22815 1003 22917
rect 321 22781 325 22815
rect 325 22781 359 22815
rect 359 22781 461 22815
rect 461 22781 495 22815
rect 495 22781 597 22815
rect 597 22781 631 22815
rect 631 22781 733 22815
rect 733 22781 767 22815
rect 767 22781 869 22815
rect 869 22781 903 22815
rect 903 22781 1003 22815
rect 321 22679 1003 22781
rect 321 22645 325 22679
rect 325 22645 359 22679
rect 359 22645 461 22679
rect 461 22645 495 22679
rect 495 22645 597 22679
rect 597 22645 631 22679
rect 631 22645 733 22679
rect 733 22645 767 22679
rect 767 22645 869 22679
rect 869 22645 903 22679
rect 903 22645 1003 22679
rect 321 22543 1003 22645
rect 321 22509 325 22543
rect 325 22509 359 22543
rect 359 22509 461 22543
rect 461 22509 495 22543
rect 495 22509 597 22543
rect 597 22509 631 22543
rect 631 22509 733 22543
rect 733 22509 767 22543
rect 767 22509 869 22543
rect 869 22509 903 22543
rect 903 22509 1003 22543
rect 321 22407 1003 22509
rect 321 22373 325 22407
rect 325 22373 359 22407
rect 359 22373 461 22407
rect 461 22373 495 22407
rect 495 22373 597 22407
rect 597 22373 631 22407
rect 631 22373 733 22407
rect 733 22373 767 22407
rect 767 22373 869 22407
rect 869 22373 903 22407
rect 903 22373 1003 22407
rect 321 22271 1003 22373
rect 321 22237 325 22271
rect 325 22237 359 22271
rect 359 22237 461 22271
rect 461 22237 495 22271
rect 495 22237 597 22271
rect 597 22237 631 22271
rect 631 22237 733 22271
rect 733 22237 767 22271
rect 767 22237 869 22271
rect 869 22237 903 22271
rect 903 22237 1003 22271
rect 321 22135 1003 22237
rect 321 22101 325 22135
rect 325 22101 359 22135
rect 359 22101 461 22135
rect 461 22101 495 22135
rect 495 22101 597 22135
rect 597 22101 631 22135
rect 631 22101 733 22135
rect 733 22101 767 22135
rect 767 22101 869 22135
rect 869 22101 903 22135
rect 903 22101 1003 22135
rect 321 21999 1003 22101
rect 321 21965 325 21999
rect 325 21965 359 21999
rect 359 21965 461 21999
rect 461 21965 495 21999
rect 495 21965 597 21999
rect 597 21965 631 21999
rect 631 21965 733 21999
rect 733 21965 767 21999
rect 767 21965 869 21999
rect 869 21965 903 21999
rect 903 21965 1003 21999
rect 321 21863 1003 21965
rect 321 21829 325 21863
rect 325 21829 359 21863
rect 359 21829 461 21863
rect 461 21829 495 21863
rect 495 21829 597 21863
rect 597 21829 631 21863
rect 631 21829 733 21863
rect 733 21829 767 21863
rect 767 21829 869 21863
rect 869 21829 903 21863
rect 903 21829 1003 21863
rect 321 21727 1003 21829
rect 321 21693 325 21727
rect 325 21693 359 21727
rect 359 21693 461 21727
rect 461 21693 495 21727
rect 495 21693 597 21727
rect 597 21693 631 21727
rect 631 21693 733 21727
rect 733 21693 767 21727
rect 767 21693 869 21727
rect 869 21693 903 21727
rect 903 21693 1003 21727
rect 321 21591 1003 21693
rect 321 21557 325 21591
rect 325 21557 359 21591
rect 359 21557 461 21591
rect 461 21557 495 21591
rect 495 21557 597 21591
rect 597 21557 631 21591
rect 631 21557 733 21591
rect 733 21557 767 21591
rect 767 21557 869 21591
rect 869 21557 903 21591
rect 903 21557 1003 21591
rect 321 21455 1003 21557
rect 321 21421 325 21455
rect 325 21421 359 21455
rect 359 21421 461 21455
rect 461 21421 495 21455
rect 495 21421 597 21455
rect 597 21421 631 21455
rect 631 21421 733 21455
rect 733 21421 767 21455
rect 767 21421 869 21455
rect 869 21421 903 21455
rect 903 21421 1003 21455
rect 321 21319 1003 21421
rect 321 21285 325 21319
rect 325 21285 359 21319
rect 359 21285 461 21319
rect 461 21285 495 21319
rect 495 21285 597 21319
rect 597 21285 631 21319
rect 631 21285 733 21319
rect 733 21285 767 21319
rect 767 21285 869 21319
rect 869 21285 903 21319
rect 903 21285 1003 21319
rect 321 21183 1003 21285
rect 321 21149 325 21183
rect 325 21149 359 21183
rect 359 21149 461 21183
rect 461 21149 495 21183
rect 495 21149 597 21183
rect 597 21149 631 21183
rect 631 21149 733 21183
rect 733 21149 767 21183
rect 767 21149 869 21183
rect 869 21149 903 21183
rect 903 21149 1003 21183
rect 321 21047 1003 21149
rect 321 21013 325 21047
rect 325 21013 359 21047
rect 359 21013 461 21047
rect 461 21013 495 21047
rect 495 21013 597 21047
rect 597 21013 631 21047
rect 631 21013 733 21047
rect 733 21013 767 21047
rect 767 21013 869 21047
rect 869 21013 903 21047
rect 903 21013 1003 21047
rect 321 20911 1003 21013
rect 321 20877 325 20911
rect 325 20877 359 20911
rect 359 20877 461 20911
rect 461 20877 495 20911
rect 495 20877 597 20911
rect 597 20877 631 20911
rect 631 20877 733 20911
rect 733 20877 767 20911
rect 767 20877 869 20911
rect 869 20877 903 20911
rect 903 20877 1003 20911
rect 321 20775 1003 20877
rect 321 20741 325 20775
rect 325 20741 359 20775
rect 359 20741 461 20775
rect 461 20741 495 20775
rect 495 20741 597 20775
rect 597 20741 631 20775
rect 631 20741 733 20775
rect 733 20741 767 20775
rect 767 20741 869 20775
rect 869 20741 903 20775
rect 903 20741 1003 20775
rect 321 20639 1003 20741
rect 321 20605 325 20639
rect 325 20605 359 20639
rect 359 20605 461 20639
rect 461 20605 495 20639
rect 495 20605 597 20639
rect 597 20605 631 20639
rect 631 20605 733 20639
rect 733 20605 767 20639
rect 767 20605 869 20639
rect 869 20605 903 20639
rect 903 20605 1003 20639
rect 321 20503 1003 20605
rect 321 20469 325 20503
rect 325 20469 359 20503
rect 359 20469 461 20503
rect 461 20469 495 20503
rect 495 20469 597 20503
rect 597 20469 631 20503
rect 631 20469 733 20503
rect 733 20469 767 20503
rect 767 20469 869 20503
rect 869 20469 903 20503
rect 903 20469 1003 20503
rect 321 20367 1003 20469
rect 321 20333 325 20367
rect 325 20333 359 20367
rect 359 20333 461 20367
rect 461 20333 495 20367
rect 495 20333 597 20367
rect 597 20333 631 20367
rect 631 20333 733 20367
rect 733 20333 767 20367
rect 767 20333 869 20367
rect 869 20333 903 20367
rect 903 20333 1003 20367
rect 321 20231 1003 20333
rect 321 20197 325 20231
rect 325 20197 359 20231
rect 359 20197 461 20231
rect 461 20197 495 20231
rect 495 20197 597 20231
rect 597 20197 631 20231
rect 631 20197 733 20231
rect 733 20197 767 20231
rect 767 20197 869 20231
rect 869 20197 903 20231
rect 903 20197 1003 20231
rect 321 20095 1003 20197
rect 321 20061 325 20095
rect 325 20061 359 20095
rect 359 20061 461 20095
rect 461 20061 495 20095
rect 495 20061 597 20095
rect 597 20061 631 20095
rect 631 20061 733 20095
rect 733 20061 767 20095
rect 767 20061 869 20095
rect 869 20061 903 20095
rect 903 20061 1003 20095
rect 321 19959 1003 20061
rect 321 19925 325 19959
rect 325 19925 359 19959
rect 359 19925 461 19959
rect 461 19925 495 19959
rect 495 19925 597 19959
rect 597 19925 631 19959
rect 631 19925 733 19959
rect 733 19925 767 19959
rect 767 19925 869 19959
rect 869 19925 903 19959
rect 903 19925 1003 19959
rect 321 19823 1003 19925
rect 321 19789 325 19823
rect 325 19789 359 19823
rect 359 19789 461 19823
rect 461 19789 495 19823
rect 495 19789 597 19823
rect 597 19789 631 19823
rect 631 19789 733 19823
rect 733 19789 767 19823
rect 767 19789 869 19823
rect 869 19789 903 19823
rect 903 19789 1003 19823
rect 321 19687 1003 19789
rect 321 19653 325 19687
rect 325 19653 359 19687
rect 359 19653 461 19687
rect 461 19653 495 19687
rect 495 19653 597 19687
rect 597 19653 631 19687
rect 631 19653 733 19687
rect 733 19653 767 19687
rect 767 19653 869 19687
rect 869 19653 903 19687
rect 903 19653 1003 19687
rect 321 19551 1003 19653
rect 321 19517 325 19551
rect 325 19517 359 19551
rect 359 19517 461 19551
rect 461 19517 495 19551
rect 495 19517 597 19551
rect 597 19517 631 19551
rect 631 19517 733 19551
rect 733 19517 767 19551
rect 767 19517 869 19551
rect 869 19517 903 19551
rect 903 19517 1003 19551
rect 321 19415 1003 19517
rect 321 19381 325 19415
rect 325 19381 359 19415
rect 359 19381 461 19415
rect 461 19381 495 19415
rect 495 19381 597 19415
rect 597 19381 631 19415
rect 631 19381 733 19415
rect 733 19381 767 19415
rect 767 19381 869 19415
rect 869 19381 903 19415
rect 903 19381 1003 19415
rect 321 19279 1003 19381
rect 321 19245 325 19279
rect 325 19245 359 19279
rect 359 19245 461 19279
rect 461 19245 495 19279
rect 495 19245 597 19279
rect 597 19245 631 19279
rect 631 19245 733 19279
rect 733 19245 767 19279
rect 767 19245 869 19279
rect 869 19245 903 19279
rect 903 19245 1003 19279
rect 321 19143 1003 19245
rect 321 19109 325 19143
rect 325 19109 359 19143
rect 359 19109 461 19143
rect 461 19109 495 19143
rect 495 19109 597 19143
rect 597 19109 631 19143
rect 631 19109 733 19143
rect 733 19109 767 19143
rect 767 19109 869 19143
rect 869 19109 903 19143
rect 903 19109 1003 19143
rect 321 19007 1003 19109
rect 321 18973 325 19007
rect 325 18973 359 19007
rect 359 18973 461 19007
rect 461 18973 495 19007
rect 495 18973 597 19007
rect 597 18973 631 19007
rect 631 18973 733 19007
rect 733 18973 767 19007
rect 767 18973 869 19007
rect 869 18973 903 19007
rect 903 18973 1003 19007
rect 321 18871 1003 18973
rect 321 18837 325 18871
rect 325 18837 359 18871
rect 359 18837 461 18871
rect 461 18837 495 18871
rect 495 18837 597 18871
rect 597 18837 631 18871
rect 631 18837 733 18871
rect 733 18837 767 18871
rect 767 18837 869 18871
rect 869 18837 903 18871
rect 903 18837 1003 18871
rect 321 18735 1003 18837
rect 321 18701 325 18735
rect 325 18701 359 18735
rect 359 18701 461 18735
rect 461 18701 495 18735
rect 495 18701 597 18735
rect 597 18701 631 18735
rect 631 18701 733 18735
rect 733 18701 767 18735
rect 767 18701 869 18735
rect 869 18701 903 18735
rect 903 18701 1003 18735
rect 321 18599 1003 18701
rect 321 18565 325 18599
rect 325 18565 359 18599
rect 359 18565 461 18599
rect 461 18565 495 18599
rect 495 18565 597 18599
rect 597 18565 631 18599
rect 631 18565 733 18599
rect 733 18565 767 18599
rect 767 18565 869 18599
rect 869 18565 903 18599
rect 903 18565 1003 18599
rect 321 18463 1003 18565
rect 321 18429 325 18463
rect 325 18429 359 18463
rect 359 18429 461 18463
rect 461 18429 495 18463
rect 495 18429 597 18463
rect 597 18429 631 18463
rect 631 18429 733 18463
rect 733 18429 767 18463
rect 767 18429 869 18463
rect 869 18429 903 18463
rect 903 18429 1003 18463
rect 321 18327 1003 18429
rect 321 18293 325 18327
rect 325 18293 359 18327
rect 359 18293 461 18327
rect 461 18293 495 18327
rect 495 18293 597 18327
rect 597 18293 631 18327
rect 631 18293 733 18327
rect 733 18293 767 18327
rect 767 18293 869 18327
rect 869 18293 903 18327
rect 903 18293 1003 18327
rect 321 18191 1003 18293
rect 321 18157 325 18191
rect 325 18157 359 18191
rect 359 18157 461 18191
rect 461 18157 495 18191
rect 495 18157 597 18191
rect 597 18157 631 18191
rect 631 18157 733 18191
rect 733 18157 767 18191
rect 767 18157 869 18191
rect 869 18157 903 18191
rect 903 18157 1003 18191
rect 321 18055 1003 18157
rect 321 18021 325 18055
rect 325 18021 359 18055
rect 359 18021 461 18055
rect 461 18021 495 18055
rect 495 18021 597 18055
rect 597 18021 631 18055
rect 631 18021 733 18055
rect 733 18021 767 18055
rect 767 18021 869 18055
rect 869 18021 903 18055
rect 903 18021 1003 18055
rect 321 17919 1003 18021
rect 321 17885 325 17919
rect 325 17885 359 17919
rect 359 17885 461 17919
rect 461 17885 495 17919
rect 495 17885 597 17919
rect 597 17885 631 17919
rect 631 17885 733 17919
rect 733 17885 767 17919
rect 767 17885 869 17919
rect 869 17885 903 17919
rect 903 17885 1003 17919
rect 321 17783 1003 17885
rect 321 17749 325 17783
rect 325 17749 359 17783
rect 359 17749 461 17783
rect 461 17749 495 17783
rect 495 17749 597 17783
rect 597 17749 631 17783
rect 631 17749 733 17783
rect 733 17749 767 17783
rect 767 17749 869 17783
rect 869 17749 903 17783
rect 903 17749 1003 17783
rect 321 17647 1003 17749
rect 321 17613 325 17647
rect 325 17613 359 17647
rect 359 17613 461 17647
rect 461 17613 495 17647
rect 495 17613 597 17647
rect 597 17613 631 17647
rect 631 17613 733 17647
rect 733 17613 767 17647
rect 767 17613 869 17647
rect 869 17613 903 17647
rect 903 17613 1003 17647
rect 321 17511 1003 17613
rect 8596 29479 9278 29511
rect 8596 29445 8696 29479
rect 8696 29445 8730 29479
rect 8730 29445 8832 29479
rect 8832 29445 8866 29479
rect 8866 29445 8968 29479
rect 8968 29445 9002 29479
rect 9002 29445 9104 29479
rect 9104 29445 9138 29479
rect 9138 29445 9240 29479
rect 9240 29445 9274 29479
rect 9274 29445 9278 29479
rect 8596 29343 9278 29445
rect 8596 29309 8696 29343
rect 8696 29309 8730 29343
rect 8730 29309 8832 29343
rect 8832 29309 8866 29343
rect 8866 29309 8968 29343
rect 8968 29309 9002 29343
rect 9002 29309 9104 29343
rect 9104 29309 9138 29343
rect 9138 29309 9240 29343
rect 9240 29309 9274 29343
rect 9274 29309 9278 29343
rect 8596 29207 9278 29309
rect 8596 29173 8696 29207
rect 8696 29173 8730 29207
rect 8730 29173 8832 29207
rect 8832 29173 8866 29207
rect 8866 29173 8968 29207
rect 8968 29173 9002 29207
rect 9002 29173 9104 29207
rect 9104 29173 9138 29207
rect 9138 29173 9240 29207
rect 9240 29173 9274 29207
rect 9274 29173 9278 29207
rect 8596 29071 9278 29173
rect 8596 29037 8696 29071
rect 8696 29037 8730 29071
rect 8730 29037 8832 29071
rect 8832 29037 8866 29071
rect 8866 29037 8968 29071
rect 8968 29037 9002 29071
rect 9002 29037 9104 29071
rect 9104 29037 9138 29071
rect 9138 29037 9240 29071
rect 9240 29037 9274 29071
rect 9274 29037 9278 29071
rect 8596 28935 9278 29037
rect 8596 28901 8696 28935
rect 8696 28901 8730 28935
rect 8730 28901 8832 28935
rect 8832 28901 8866 28935
rect 8866 28901 8968 28935
rect 8968 28901 9002 28935
rect 9002 28901 9104 28935
rect 9104 28901 9138 28935
rect 9138 28901 9240 28935
rect 9240 28901 9274 28935
rect 9274 28901 9278 28935
rect 8596 28799 9278 28901
rect 8596 28765 8696 28799
rect 8696 28765 8730 28799
rect 8730 28765 8832 28799
rect 8832 28765 8866 28799
rect 8866 28765 8968 28799
rect 8968 28765 9002 28799
rect 9002 28765 9104 28799
rect 9104 28765 9138 28799
rect 9138 28765 9240 28799
rect 9240 28765 9274 28799
rect 9274 28765 9278 28799
rect 8596 28663 9278 28765
rect 8596 28629 8696 28663
rect 8696 28629 8730 28663
rect 8730 28629 8832 28663
rect 8832 28629 8866 28663
rect 8866 28629 8968 28663
rect 8968 28629 9002 28663
rect 9002 28629 9104 28663
rect 9104 28629 9138 28663
rect 9138 28629 9240 28663
rect 9240 28629 9274 28663
rect 9274 28629 9278 28663
rect 8596 28527 9278 28629
rect 8596 28493 8696 28527
rect 8696 28493 8730 28527
rect 8730 28493 8832 28527
rect 8832 28493 8866 28527
rect 8866 28493 8968 28527
rect 8968 28493 9002 28527
rect 9002 28493 9104 28527
rect 9104 28493 9138 28527
rect 9138 28493 9240 28527
rect 9240 28493 9274 28527
rect 9274 28493 9278 28527
rect 8596 28391 9278 28493
rect 8596 28357 8696 28391
rect 8696 28357 8730 28391
rect 8730 28357 8832 28391
rect 8832 28357 8866 28391
rect 8866 28357 8968 28391
rect 8968 28357 9002 28391
rect 9002 28357 9104 28391
rect 9104 28357 9138 28391
rect 9138 28357 9240 28391
rect 9240 28357 9274 28391
rect 9274 28357 9278 28391
rect 8596 28255 9278 28357
rect 8596 28221 8696 28255
rect 8696 28221 8730 28255
rect 8730 28221 8832 28255
rect 8832 28221 8866 28255
rect 8866 28221 8968 28255
rect 8968 28221 9002 28255
rect 9002 28221 9104 28255
rect 9104 28221 9138 28255
rect 9138 28221 9240 28255
rect 9240 28221 9274 28255
rect 9274 28221 9278 28255
rect 8596 28119 9278 28221
rect 8596 28085 8696 28119
rect 8696 28085 8730 28119
rect 8730 28085 8832 28119
rect 8832 28085 8866 28119
rect 8866 28085 8968 28119
rect 8968 28085 9002 28119
rect 9002 28085 9104 28119
rect 9104 28085 9138 28119
rect 9138 28085 9240 28119
rect 9240 28085 9274 28119
rect 9274 28085 9278 28119
rect 8596 27983 9278 28085
rect 8596 27949 8696 27983
rect 8696 27949 8730 27983
rect 8730 27949 8832 27983
rect 8832 27949 8866 27983
rect 8866 27949 8968 27983
rect 8968 27949 9002 27983
rect 9002 27949 9104 27983
rect 9104 27949 9138 27983
rect 9138 27949 9240 27983
rect 9240 27949 9274 27983
rect 9274 27949 9278 27983
rect 8596 27847 9278 27949
rect 8596 27813 8696 27847
rect 8696 27813 8730 27847
rect 8730 27813 8832 27847
rect 8832 27813 8866 27847
rect 8866 27813 8968 27847
rect 8968 27813 9002 27847
rect 9002 27813 9104 27847
rect 9104 27813 9138 27847
rect 9138 27813 9240 27847
rect 9240 27813 9274 27847
rect 9274 27813 9278 27847
rect 8596 27711 9278 27813
rect 8596 27677 8696 27711
rect 8696 27677 8730 27711
rect 8730 27677 8832 27711
rect 8832 27677 8866 27711
rect 8866 27677 8968 27711
rect 8968 27677 9002 27711
rect 9002 27677 9104 27711
rect 9104 27677 9138 27711
rect 9138 27677 9240 27711
rect 9240 27677 9274 27711
rect 9274 27677 9278 27711
rect 8596 27575 9278 27677
rect 8596 27541 8696 27575
rect 8696 27541 8730 27575
rect 8730 27541 8832 27575
rect 8832 27541 8866 27575
rect 8866 27541 8968 27575
rect 8968 27541 9002 27575
rect 9002 27541 9104 27575
rect 9104 27541 9138 27575
rect 9138 27541 9240 27575
rect 9240 27541 9274 27575
rect 9274 27541 9278 27575
rect 8596 27439 9278 27541
rect 8596 27405 8696 27439
rect 8696 27405 8730 27439
rect 8730 27405 8832 27439
rect 8832 27405 8866 27439
rect 8866 27405 8968 27439
rect 8968 27405 9002 27439
rect 9002 27405 9104 27439
rect 9104 27405 9138 27439
rect 9138 27405 9240 27439
rect 9240 27405 9274 27439
rect 9274 27405 9278 27439
rect 8596 27303 9278 27405
rect 8596 27269 8696 27303
rect 8696 27269 8730 27303
rect 8730 27269 8832 27303
rect 8832 27269 8866 27303
rect 8866 27269 8968 27303
rect 8968 27269 9002 27303
rect 9002 27269 9104 27303
rect 9104 27269 9138 27303
rect 9138 27269 9240 27303
rect 9240 27269 9274 27303
rect 9274 27269 9278 27303
rect 8596 27167 9278 27269
rect 8596 27133 8696 27167
rect 8696 27133 8730 27167
rect 8730 27133 8832 27167
rect 8832 27133 8866 27167
rect 8866 27133 8968 27167
rect 8968 27133 9002 27167
rect 9002 27133 9104 27167
rect 9104 27133 9138 27167
rect 9138 27133 9240 27167
rect 9240 27133 9274 27167
rect 9274 27133 9278 27167
rect 8596 27031 9278 27133
rect 8596 26997 8696 27031
rect 8696 26997 8730 27031
rect 8730 26997 8832 27031
rect 8832 26997 8866 27031
rect 8866 26997 8968 27031
rect 8968 26997 9002 27031
rect 9002 26997 9104 27031
rect 9104 26997 9138 27031
rect 9138 26997 9240 27031
rect 9240 26997 9274 27031
rect 9274 26997 9278 27031
rect 8596 26895 9278 26997
rect 8596 26861 8696 26895
rect 8696 26861 8730 26895
rect 8730 26861 8832 26895
rect 8832 26861 8866 26895
rect 8866 26861 8968 26895
rect 8968 26861 9002 26895
rect 9002 26861 9104 26895
rect 9104 26861 9138 26895
rect 9138 26861 9240 26895
rect 9240 26861 9274 26895
rect 9274 26861 9278 26895
rect 8596 26759 9278 26861
rect 8596 26725 8696 26759
rect 8696 26725 8730 26759
rect 8730 26725 8832 26759
rect 8832 26725 8866 26759
rect 8866 26725 8968 26759
rect 8968 26725 9002 26759
rect 9002 26725 9104 26759
rect 9104 26725 9138 26759
rect 9138 26725 9240 26759
rect 9240 26725 9274 26759
rect 9274 26725 9278 26759
rect 8596 26623 9278 26725
rect 8596 26589 8696 26623
rect 8696 26589 8730 26623
rect 8730 26589 8832 26623
rect 8832 26589 8866 26623
rect 8866 26589 8968 26623
rect 8968 26589 9002 26623
rect 9002 26589 9104 26623
rect 9104 26589 9138 26623
rect 9138 26589 9240 26623
rect 9240 26589 9274 26623
rect 9274 26589 9278 26623
rect 8596 26487 9278 26589
rect 8596 26453 8696 26487
rect 8696 26453 8730 26487
rect 8730 26453 8832 26487
rect 8832 26453 8866 26487
rect 8866 26453 8968 26487
rect 8968 26453 9002 26487
rect 9002 26453 9104 26487
rect 9104 26453 9138 26487
rect 9138 26453 9240 26487
rect 9240 26453 9274 26487
rect 9274 26453 9278 26487
rect 8596 26351 9278 26453
rect 8596 26317 8696 26351
rect 8696 26317 8730 26351
rect 8730 26317 8832 26351
rect 8832 26317 8866 26351
rect 8866 26317 8968 26351
rect 8968 26317 9002 26351
rect 9002 26317 9104 26351
rect 9104 26317 9138 26351
rect 9138 26317 9240 26351
rect 9240 26317 9274 26351
rect 9274 26317 9278 26351
rect 8596 26215 9278 26317
rect 8596 26181 8696 26215
rect 8696 26181 8730 26215
rect 8730 26181 8832 26215
rect 8832 26181 8866 26215
rect 8866 26181 8968 26215
rect 8968 26181 9002 26215
rect 9002 26181 9104 26215
rect 9104 26181 9138 26215
rect 9138 26181 9240 26215
rect 9240 26181 9274 26215
rect 9274 26181 9278 26215
rect 8596 26079 9278 26181
rect 8596 26045 8696 26079
rect 8696 26045 8730 26079
rect 8730 26045 8832 26079
rect 8832 26045 8866 26079
rect 8866 26045 8968 26079
rect 8968 26045 9002 26079
rect 9002 26045 9104 26079
rect 9104 26045 9138 26079
rect 9138 26045 9240 26079
rect 9240 26045 9274 26079
rect 9274 26045 9278 26079
rect 8596 25943 9278 26045
rect 8596 25909 8696 25943
rect 8696 25909 8730 25943
rect 8730 25909 8832 25943
rect 8832 25909 8866 25943
rect 8866 25909 8968 25943
rect 8968 25909 9002 25943
rect 9002 25909 9104 25943
rect 9104 25909 9138 25943
rect 9138 25909 9240 25943
rect 9240 25909 9274 25943
rect 9274 25909 9278 25943
rect 8596 25807 9278 25909
rect 8596 25773 8696 25807
rect 8696 25773 8730 25807
rect 8730 25773 8832 25807
rect 8832 25773 8866 25807
rect 8866 25773 8968 25807
rect 8968 25773 9002 25807
rect 9002 25773 9104 25807
rect 9104 25773 9138 25807
rect 9138 25773 9240 25807
rect 9240 25773 9274 25807
rect 9274 25773 9278 25807
rect 8596 25671 9278 25773
rect 8596 25637 8696 25671
rect 8696 25637 8730 25671
rect 8730 25637 8832 25671
rect 8832 25637 8866 25671
rect 8866 25637 8968 25671
rect 8968 25637 9002 25671
rect 9002 25637 9104 25671
rect 9104 25637 9138 25671
rect 9138 25637 9240 25671
rect 9240 25637 9274 25671
rect 9274 25637 9278 25671
rect 8596 25535 9278 25637
rect 8596 25501 8696 25535
rect 8696 25501 8730 25535
rect 8730 25501 8832 25535
rect 8832 25501 8866 25535
rect 8866 25501 8968 25535
rect 8968 25501 9002 25535
rect 9002 25501 9104 25535
rect 9104 25501 9138 25535
rect 9138 25501 9240 25535
rect 9240 25501 9274 25535
rect 9274 25501 9278 25535
rect 8596 25399 9278 25501
rect 8596 25365 8696 25399
rect 8696 25365 8730 25399
rect 8730 25365 8832 25399
rect 8832 25365 8866 25399
rect 8866 25365 8968 25399
rect 8968 25365 9002 25399
rect 9002 25365 9104 25399
rect 9104 25365 9138 25399
rect 9138 25365 9240 25399
rect 9240 25365 9274 25399
rect 9274 25365 9278 25399
rect 8596 25263 9278 25365
rect 8596 25229 8696 25263
rect 8696 25229 8730 25263
rect 8730 25229 8832 25263
rect 8832 25229 8866 25263
rect 8866 25229 8968 25263
rect 8968 25229 9002 25263
rect 9002 25229 9104 25263
rect 9104 25229 9138 25263
rect 9138 25229 9240 25263
rect 9240 25229 9274 25263
rect 9274 25229 9278 25263
rect 8596 25127 9278 25229
rect 8596 25093 8696 25127
rect 8696 25093 8730 25127
rect 8730 25093 8832 25127
rect 8832 25093 8866 25127
rect 8866 25093 8968 25127
rect 8968 25093 9002 25127
rect 9002 25093 9104 25127
rect 9104 25093 9138 25127
rect 9138 25093 9240 25127
rect 9240 25093 9274 25127
rect 9274 25093 9278 25127
rect 8596 24991 9278 25093
rect 8596 24957 8696 24991
rect 8696 24957 8730 24991
rect 8730 24957 8832 24991
rect 8832 24957 8866 24991
rect 8866 24957 8968 24991
rect 8968 24957 9002 24991
rect 9002 24957 9104 24991
rect 9104 24957 9138 24991
rect 9138 24957 9240 24991
rect 9240 24957 9274 24991
rect 9274 24957 9278 24991
rect 8596 24855 9278 24957
rect 8596 24821 8696 24855
rect 8696 24821 8730 24855
rect 8730 24821 8832 24855
rect 8832 24821 8866 24855
rect 8866 24821 8968 24855
rect 8968 24821 9002 24855
rect 9002 24821 9104 24855
rect 9104 24821 9138 24855
rect 9138 24821 9240 24855
rect 9240 24821 9274 24855
rect 9274 24821 9278 24855
rect 8596 24719 9278 24821
rect 8596 24685 8696 24719
rect 8696 24685 8730 24719
rect 8730 24685 8832 24719
rect 8832 24685 8866 24719
rect 8866 24685 8968 24719
rect 8968 24685 9002 24719
rect 9002 24685 9104 24719
rect 9104 24685 9138 24719
rect 9138 24685 9240 24719
rect 9240 24685 9274 24719
rect 9274 24685 9278 24719
rect 8596 24583 9278 24685
rect 8596 24549 8696 24583
rect 8696 24549 8730 24583
rect 8730 24549 8832 24583
rect 8832 24549 8866 24583
rect 8866 24549 8968 24583
rect 8968 24549 9002 24583
rect 9002 24549 9104 24583
rect 9104 24549 9138 24583
rect 9138 24549 9240 24583
rect 9240 24549 9274 24583
rect 9274 24549 9278 24583
rect 8596 24447 9278 24549
rect 8596 24413 8696 24447
rect 8696 24413 8730 24447
rect 8730 24413 8832 24447
rect 8832 24413 8866 24447
rect 8866 24413 8968 24447
rect 8968 24413 9002 24447
rect 9002 24413 9104 24447
rect 9104 24413 9138 24447
rect 9138 24413 9240 24447
rect 9240 24413 9274 24447
rect 9274 24413 9278 24447
rect 8596 24311 9278 24413
rect 8596 24277 8696 24311
rect 8696 24277 8730 24311
rect 8730 24277 8832 24311
rect 8832 24277 8866 24311
rect 8866 24277 8968 24311
rect 8968 24277 9002 24311
rect 9002 24277 9104 24311
rect 9104 24277 9138 24311
rect 9138 24277 9240 24311
rect 9240 24277 9274 24311
rect 9274 24277 9278 24311
rect 8596 24175 9278 24277
rect 8596 24141 8696 24175
rect 8696 24141 8730 24175
rect 8730 24141 8832 24175
rect 8832 24141 8866 24175
rect 8866 24141 8968 24175
rect 8968 24141 9002 24175
rect 9002 24141 9104 24175
rect 9104 24141 9138 24175
rect 9138 24141 9240 24175
rect 9240 24141 9274 24175
rect 9274 24141 9278 24175
rect 8596 24039 9278 24141
rect 8596 24005 8696 24039
rect 8696 24005 8730 24039
rect 8730 24005 8832 24039
rect 8832 24005 8866 24039
rect 8866 24005 8968 24039
rect 8968 24005 9002 24039
rect 9002 24005 9104 24039
rect 9104 24005 9138 24039
rect 9138 24005 9240 24039
rect 9240 24005 9274 24039
rect 9274 24005 9278 24039
rect 8596 23903 9278 24005
rect 8596 23869 8696 23903
rect 8696 23869 8730 23903
rect 8730 23869 8832 23903
rect 8832 23869 8866 23903
rect 8866 23869 8968 23903
rect 8968 23869 9002 23903
rect 9002 23869 9104 23903
rect 9104 23869 9138 23903
rect 9138 23869 9240 23903
rect 9240 23869 9274 23903
rect 9274 23869 9278 23903
rect 8596 23767 9278 23869
rect 8596 23733 8696 23767
rect 8696 23733 8730 23767
rect 8730 23733 8832 23767
rect 8832 23733 8866 23767
rect 8866 23733 8968 23767
rect 8968 23733 9002 23767
rect 9002 23733 9104 23767
rect 9104 23733 9138 23767
rect 9138 23733 9240 23767
rect 9240 23733 9274 23767
rect 9274 23733 9278 23767
rect 8596 23631 9278 23733
rect 8596 23597 8696 23631
rect 8696 23597 8730 23631
rect 8730 23597 8832 23631
rect 8832 23597 8866 23631
rect 8866 23597 8968 23631
rect 8968 23597 9002 23631
rect 9002 23597 9104 23631
rect 9104 23597 9138 23631
rect 9138 23597 9240 23631
rect 9240 23597 9274 23631
rect 9274 23597 9278 23631
rect 8596 23495 9278 23597
rect 8596 23461 8696 23495
rect 8696 23461 8730 23495
rect 8730 23461 8832 23495
rect 8832 23461 8866 23495
rect 8866 23461 8968 23495
rect 8968 23461 9002 23495
rect 9002 23461 9104 23495
rect 9104 23461 9138 23495
rect 9138 23461 9240 23495
rect 9240 23461 9274 23495
rect 9274 23461 9278 23495
rect 8596 23359 9278 23461
rect 8596 23325 8696 23359
rect 8696 23325 8730 23359
rect 8730 23325 8832 23359
rect 8832 23325 8866 23359
rect 8866 23325 8968 23359
rect 8968 23325 9002 23359
rect 9002 23325 9104 23359
rect 9104 23325 9138 23359
rect 9138 23325 9240 23359
rect 9240 23325 9274 23359
rect 9274 23325 9278 23359
rect 8596 23223 9278 23325
rect 8596 23189 8696 23223
rect 8696 23189 8730 23223
rect 8730 23189 8832 23223
rect 8832 23189 8866 23223
rect 8866 23189 8968 23223
rect 8968 23189 9002 23223
rect 9002 23189 9104 23223
rect 9104 23189 9138 23223
rect 9138 23189 9240 23223
rect 9240 23189 9274 23223
rect 9274 23189 9278 23223
rect 8596 23087 9278 23189
rect 8596 23053 8696 23087
rect 8696 23053 8730 23087
rect 8730 23053 8832 23087
rect 8832 23053 8866 23087
rect 8866 23053 8968 23087
rect 8968 23053 9002 23087
rect 9002 23053 9104 23087
rect 9104 23053 9138 23087
rect 9138 23053 9240 23087
rect 9240 23053 9274 23087
rect 9274 23053 9278 23087
rect 8596 22951 9278 23053
rect 8596 22917 8696 22951
rect 8696 22917 8730 22951
rect 8730 22917 8832 22951
rect 8832 22917 8866 22951
rect 8866 22917 8968 22951
rect 8968 22917 9002 22951
rect 9002 22917 9104 22951
rect 9104 22917 9138 22951
rect 9138 22917 9240 22951
rect 9240 22917 9274 22951
rect 9274 22917 9278 22951
rect 8596 22815 9278 22917
rect 8596 22781 8696 22815
rect 8696 22781 8730 22815
rect 8730 22781 8832 22815
rect 8832 22781 8866 22815
rect 8866 22781 8968 22815
rect 8968 22781 9002 22815
rect 9002 22781 9104 22815
rect 9104 22781 9138 22815
rect 9138 22781 9240 22815
rect 9240 22781 9274 22815
rect 9274 22781 9278 22815
rect 8596 22679 9278 22781
rect 8596 22645 8696 22679
rect 8696 22645 8730 22679
rect 8730 22645 8832 22679
rect 8832 22645 8866 22679
rect 8866 22645 8968 22679
rect 8968 22645 9002 22679
rect 9002 22645 9104 22679
rect 9104 22645 9138 22679
rect 9138 22645 9240 22679
rect 9240 22645 9274 22679
rect 9274 22645 9278 22679
rect 8596 22543 9278 22645
rect 8596 22509 8696 22543
rect 8696 22509 8730 22543
rect 8730 22509 8832 22543
rect 8832 22509 8866 22543
rect 8866 22509 8968 22543
rect 8968 22509 9002 22543
rect 9002 22509 9104 22543
rect 9104 22509 9138 22543
rect 9138 22509 9240 22543
rect 9240 22509 9274 22543
rect 9274 22509 9278 22543
rect 8596 22407 9278 22509
rect 8596 22373 8696 22407
rect 8696 22373 8730 22407
rect 8730 22373 8832 22407
rect 8832 22373 8866 22407
rect 8866 22373 8968 22407
rect 8968 22373 9002 22407
rect 9002 22373 9104 22407
rect 9104 22373 9138 22407
rect 9138 22373 9240 22407
rect 9240 22373 9274 22407
rect 9274 22373 9278 22407
rect 8596 22271 9278 22373
rect 8596 22237 8696 22271
rect 8696 22237 8730 22271
rect 8730 22237 8832 22271
rect 8832 22237 8866 22271
rect 8866 22237 8968 22271
rect 8968 22237 9002 22271
rect 9002 22237 9104 22271
rect 9104 22237 9138 22271
rect 9138 22237 9240 22271
rect 9240 22237 9274 22271
rect 9274 22237 9278 22271
rect 8596 22135 9278 22237
rect 8596 22101 8696 22135
rect 8696 22101 8730 22135
rect 8730 22101 8832 22135
rect 8832 22101 8866 22135
rect 8866 22101 8968 22135
rect 8968 22101 9002 22135
rect 9002 22101 9104 22135
rect 9104 22101 9138 22135
rect 9138 22101 9240 22135
rect 9240 22101 9274 22135
rect 9274 22101 9278 22135
rect 8596 21999 9278 22101
rect 8596 21965 8696 21999
rect 8696 21965 8730 21999
rect 8730 21965 8832 21999
rect 8832 21965 8866 21999
rect 8866 21965 8968 21999
rect 8968 21965 9002 21999
rect 9002 21965 9104 21999
rect 9104 21965 9138 21999
rect 9138 21965 9240 21999
rect 9240 21965 9274 21999
rect 9274 21965 9278 21999
rect 8596 21863 9278 21965
rect 8596 21829 8696 21863
rect 8696 21829 8730 21863
rect 8730 21829 8832 21863
rect 8832 21829 8866 21863
rect 8866 21829 8968 21863
rect 8968 21829 9002 21863
rect 9002 21829 9104 21863
rect 9104 21829 9138 21863
rect 9138 21829 9240 21863
rect 9240 21829 9274 21863
rect 9274 21829 9278 21863
rect 8596 21727 9278 21829
rect 8596 21693 8696 21727
rect 8696 21693 8730 21727
rect 8730 21693 8832 21727
rect 8832 21693 8866 21727
rect 8866 21693 8968 21727
rect 8968 21693 9002 21727
rect 9002 21693 9104 21727
rect 9104 21693 9138 21727
rect 9138 21693 9240 21727
rect 9240 21693 9274 21727
rect 9274 21693 9278 21727
rect 8596 21591 9278 21693
rect 8596 21557 8696 21591
rect 8696 21557 8730 21591
rect 8730 21557 8832 21591
rect 8832 21557 8866 21591
rect 8866 21557 8968 21591
rect 8968 21557 9002 21591
rect 9002 21557 9104 21591
rect 9104 21557 9138 21591
rect 9138 21557 9240 21591
rect 9240 21557 9274 21591
rect 9274 21557 9278 21591
rect 8596 21455 9278 21557
rect 8596 21421 8696 21455
rect 8696 21421 8730 21455
rect 8730 21421 8832 21455
rect 8832 21421 8866 21455
rect 8866 21421 8968 21455
rect 8968 21421 9002 21455
rect 9002 21421 9104 21455
rect 9104 21421 9138 21455
rect 9138 21421 9240 21455
rect 9240 21421 9274 21455
rect 9274 21421 9278 21455
rect 8596 21319 9278 21421
rect 8596 21285 8696 21319
rect 8696 21285 8730 21319
rect 8730 21285 8832 21319
rect 8832 21285 8866 21319
rect 8866 21285 8968 21319
rect 8968 21285 9002 21319
rect 9002 21285 9104 21319
rect 9104 21285 9138 21319
rect 9138 21285 9240 21319
rect 9240 21285 9274 21319
rect 9274 21285 9278 21319
rect 8596 21183 9278 21285
rect 8596 21149 8696 21183
rect 8696 21149 8730 21183
rect 8730 21149 8832 21183
rect 8832 21149 8866 21183
rect 8866 21149 8968 21183
rect 8968 21149 9002 21183
rect 9002 21149 9104 21183
rect 9104 21149 9138 21183
rect 9138 21149 9240 21183
rect 9240 21149 9274 21183
rect 9274 21149 9278 21183
rect 8596 21047 9278 21149
rect 8596 21013 8696 21047
rect 8696 21013 8730 21047
rect 8730 21013 8832 21047
rect 8832 21013 8866 21047
rect 8866 21013 8968 21047
rect 8968 21013 9002 21047
rect 9002 21013 9104 21047
rect 9104 21013 9138 21047
rect 9138 21013 9240 21047
rect 9240 21013 9274 21047
rect 9274 21013 9278 21047
rect 8596 20911 9278 21013
rect 8596 20877 8696 20911
rect 8696 20877 8730 20911
rect 8730 20877 8832 20911
rect 8832 20877 8866 20911
rect 8866 20877 8968 20911
rect 8968 20877 9002 20911
rect 9002 20877 9104 20911
rect 9104 20877 9138 20911
rect 9138 20877 9240 20911
rect 9240 20877 9274 20911
rect 9274 20877 9278 20911
rect 8596 20775 9278 20877
rect 8596 20741 8696 20775
rect 8696 20741 8730 20775
rect 8730 20741 8832 20775
rect 8832 20741 8866 20775
rect 8866 20741 8968 20775
rect 8968 20741 9002 20775
rect 9002 20741 9104 20775
rect 9104 20741 9138 20775
rect 9138 20741 9240 20775
rect 9240 20741 9274 20775
rect 9274 20741 9278 20775
rect 8596 20639 9278 20741
rect 8596 20605 8696 20639
rect 8696 20605 8730 20639
rect 8730 20605 8832 20639
rect 8832 20605 8866 20639
rect 8866 20605 8968 20639
rect 8968 20605 9002 20639
rect 9002 20605 9104 20639
rect 9104 20605 9138 20639
rect 9138 20605 9240 20639
rect 9240 20605 9274 20639
rect 9274 20605 9278 20639
rect 8596 20503 9278 20605
rect 8596 20469 8696 20503
rect 8696 20469 8730 20503
rect 8730 20469 8832 20503
rect 8832 20469 8866 20503
rect 8866 20469 8968 20503
rect 8968 20469 9002 20503
rect 9002 20469 9104 20503
rect 9104 20469 9138 20503
rect 9138 20469 9240 20503
rect 9240 20469 9274 20503
rect 9274 20469 9278 20503
rect 8596 20405 9278 20469
rect 8596 20332 8630 20366
rect 8668 20333 8696 20366
rect 8696 20333 8702 20366
rect 8668 20332 8702 20333
rect 8740 20332 8774 20366
rect 8812 20333 8832 20366
rect 8832 20333 8846 20366
rect 8812 20332 8846 20333
rect 8884 20332 8918 20366
rect 8956 20333 8968 20366
rect 8968 20333 8990 20366
rect 8956 20332 8990 20333
rect 9028 20332 9062 20366
rect 9100 20333 9104 20366
rect 9104 20333 9134 20366
rect 9100 20332 9134 20333
rect 9172 20332 9206 20366
rect 9244 20333 9274 20366
rect 9274 20333 9278 20366
rect 9244 20332 9278 20333
rect 8596 20259 8630 20293
rect 8668 20259 8702 20293
rect 8740 20259 8774 20293
rect 8812 20259 8846 20293
rect 8884 20259 8918 20293
rect 8956 20259 8990 20293
rect 9028 20259 9062 20293
rect 9100 20259 9134 20293
rect 9172 20259 9206 20293
rect 9244 20259 9278 20293
rect 8596 20186 8630 20220
rect 8668 20197 8696 20220
rect 8696 20197 8702 20220
rect 8668 20186 8702 20197
rect 8740 20186 8774 20220
rect 8812 20197 8832 20220
rect 8832 20197 8846 20220
rect 8812 20186 8846 20197
rect 8884 20186 8918 20220
rect 8956 20197 8968 20220
rect 8968 20197 8990 20220
rect 8956 20186 8990 20197
rect 9028 20186 9062 20220
rect 9100 20197 9104 20220
rect 9104 20197 9134 20220
rect 9100 20186 9134 20197
rect 9172 20186 9206 20220
rect 9244 20197 9274 20220
rect 9274 20197 9278 20220
rect 9244 20186 9278 20197
rect 8596 20113 8630 20147
rect 8668 20113 8702 20147
rect 8740 20113 8774 20147
rect 8812 20113 8846 20147
rect 8884 20113 8918 20147
rect 8956 20113 8990 20147
rect 9028 20113 9062 20147
rect 9100 20113 9134 20147
rect 9172 20113 9206 20147
rect 9244 20113 9278 20147
rect 8596 20040 8630 20074
rect 8668 20061 8696 20074
rect 8696 20061 8702 20074
rect 8668 20040 8702 20061
rect 8740 20040 8774 20074
rect 8812 20061 8832 20074
rect 8832 20061 8846 20074
rect 8812 20040 8846 20061
rect 8884 20040 8918 20074
rect 8956 20061 8968 20074
rect 8968 20061 8990 20074
rect 8956 20040 8990 20061
rect 9028 20040 9062 20074
rect 9100 20061 9104 20074
rect 9104 20061 9134 20074
rect 9100 20040 9134 20061
rect 9172 20040 9206 20074
rect 9244 20061 9274 20074
rect 9274 20061 9278 20074
rect 9244 20040 9278 20061
rect 8596 19967 8630 20001
rect 8668 19967 8702 20001
rect 8740 19967 8774 20001
rect 8812 19967 8846 20001
rect 8884 19967 8918 20001
rect 8956 19967 8990 20001
rect 9028 19967 9062 20001
rect 9100 19967 9134 20001
rect 9172 19967 9206 20001
rect 9244 19967 9278 20001
rect 8596 19894 8630 19928
rect 8668 19925 8696 19928
rect 8696 19925 8702 19928
rect 8668 19894 8702 19925
rect 8740 19894 8774 19928
rect 8812 19925 8832 19928
rect 8832 19925 8846 19928
rect 8812 19894 8846 19925
rect 8884 19894 8918 19928
rect 8956 19925 8968 19928
rect 8968 19925 8990 19928
rect 8956 19894 8990 19925
rect 9028 19894 9062 19928
rect 9100 19925 9104 19928
rect 9104 19925 9134 19928
rect 9100 19894 9134 19925
rect 9172 19894 9206 19928
rect 9244 19925 9274 19928
rect 9274 19925 9278 19928
rect 9244 19894 9278 19925
rect 8596 19821 8630 19855
rect 8668 19823 8702 19855
rect 8668 19821 8696 19823
rect 8696 19821 8702 19823
rect 8740 19821 8774 19855
rect 8812 19823 8846 19855
rect 8812 19821 8832 19823
rect 8832 19821 8846 19823
rect 8884 19821 8918 19855
rect 8956 19823 8990 19855
rect 8956 19821 8968 19823
rect 8968 19821 8990 19823
rect 9028 19821 9062 19855
rect 9100 19823 9134 19855
rect 9100 19821 9104 19823
rect 9104 19821 9134 19823
rect 9172 19821 9206 19855
rect 9244 19823 9278 19855
rect 9244 19821 9274 19823
rect 9274 19821 9278 19823
rect 8596 19748 8630 19782
rect 8668 19748 8702 19782
rect 8740 19748 8774 19782
rect 8812 19748 8846 19782
rect 8884 19748 8918 19782
rect 8956 19748 8990 19782
rect 9028 19748 9062 19782
rect 9100 19748 9134 19782
rect 9172 19748 9206 19782
rect 9244 19748 9278 19782
rect 8596 19675 8630 19709
rect 8668 19687 8702 19709
rect 8668 19675 8696 19687
rect 8696 19675 8702 19687
rect 8740 19675 8774 19709
rect 8812 19687 8846 19709
rect 8812 19675 8832 19687
rect 8832 19675 8846 19687
rect 8884 19675 8918 19709
rect 8956 19687 8990 19709
rect 8956 19675 8968 19687
rect 8968 19675 8990 19687
rect 9028 19675 9062 19709
rect 9100 19687 9134 19709
rect 9100 19675 9104 19687
rect 9104 19675 9134 19687
rect 9172 19675 9206 19709
rect 9244 19687 9278 19709
rect 9244 19675 9274 19687
rect 9274 19675 9278 19687
rect 8596 19602 8630 19636
rect 8668 19602 8702 19636
rect 8740 19602 8774 19636
rect 8812 19602 8846 19636
rect 8884 19602 8918 19636
rect 8956 19602 8990 19636
rect 9028 19602 9062 19636
rect 9100 19602 9134 19636
rect 9172 19602 9206 19636
rect 9244 19602 9278 19636
rect 8596 19529 8630 19563
rect 8668 19551 8702 19563
rect 8668 19529 8696 19551
rect 8696 19529 8702 19551
rect 8740 19529 8774 19563
rect 8812 19551 8846 19563
rect 8812 19529 8832 19551
rect 8832 19529 8846 19551
rect 8884 19529 8918 19563
rect 8956 19551 8990 19563
rect 8956 19529 8968 19551
rect 8968 19529 8990 19551
rect 9028 19529 9062 19563
rect 9100 19551 9134 19563
rect 9100 19529 9104 19551
rect 9104 19529 9134 19551
rect 9172 19529 9206 19563
rect 9244 19551 9278 19563
rect 9244 19529 9274 19551
rect 9274 19529 9278 19551
rect 8596 19456 8630 19490
rect 8668 19456 8702 19490
rect 8740 19456 8774 19490
rect 8812 19456 8846 19490
rect 8884 19456 8918 19490
rect 8956 19456 8990 19490
rect 9028 19456 9062 19490
rect 9100 19456 9134 19490
rect 9172 19456 9206 19490
rect 9244 19456 9278 19490
rect 8596 19383 8630 19417
rect 8668 19415 8702 19417
rect 8668 19383 8696 19415
rect 8696 19383 8702 19415
rect 8740 19383 8774 19417
rect 8812 19415 8846 19417
rect 8812 19383 8832 19415
rect 8832 19383 8846 19415
rect 8884 19383 8918 19417
rect 8956 19415 8990 19417
rect 8956 19383 8968 19415
rect 8968 19383 8990 19415
rect 9028 19383 9062 19417
rect 9100 19415 9134 19417
rect 9100 19383 9104 19415
rect 9104 19383 9134 19415
rect 9172 19383 9206 19417
rect 9244 19415 9278 19417
rect 9244 19383 9274 19415
rect 9274 19383 9278 19415
rect 8596 19310 8630 19344
rect 8668 19310 8702 19344
rect 8740 19310 8774 19344
rect 8812 19310 8846 19344
rect 8884 19310 8918 19344
rect 8956 19310 8990 19344
rect 9028 19310 9062 19344
rect 9100 19310 9134 19344
rect 9172 19310 9206 19344
rect 9244 19310 9278 19344
rect 8596 19237 8630 19271
rect 8668 19245 8696 19271
rect 8696 19245 8702 19271
rect 8668 19237 8702 19245
rect 8740 19237 8774 19271
rect 8812 19245 8832 19271
rect 8832 19245 8846 19271
rect 8812 19237 8846 19245
rect 8884 19237 8918 19271
rect 8956 19245 8968 19271
rect 8968 19245 8990 19271
rect 8956 19237 8990 19245
rect 9028 19237 9062 19271
rect 9100 19245 9104 19271
rect 9104 19245 9134 19271
rect 9100 19237 9134 19245
rect 9172 19237 9206 19271
rect 9244 19245 9274 19271
rect 9274 19245 9278 19271
rect 9244 19237 9278 19245
rect 8596 19164 8630 19198
rect 8668 19164 8702 19198
rect 8740 19164 8774 19198
rect 8812 19164 8846 19198
rect 8884 19164 8918 19198
rect 8956 19164 8990 19198
rect 9028 19164 9062 19198
rect 9100 19164 9134 19198
rect 9172 19164 9206 19198
rect 9244 19164 9278 19198
rect 8596 19091 8630 19125
rect 8668 19109 8696 19125
rect 8696 19109 8702 19125
rect 8668 19091 8702 19109
rect 8740 19091 8774 19125
rect 8812 19109 8832 19125
rect 8832 19109 8846 19125
rect 8812 19091 8846 19109
rect 8884 19091 8918 19125
rect 8956 19109 8968 19125
rect 8968 19109 8990 19125
rect 8956 19091 8990 19109
rect 9028 19091 9062 19125
rect 9100 19109 9104 19125
rect 9104 19109 9134 19125
rect 9100 19091 9134 19109
rect 9172 19091 9206 19125
rect 9244 19109 9274 19125
rect 9274 19109 9278 19125
rect 9244 19091 9278 19109
rect 8596 19018 8630 19052
rect 8668 19018 8702 19052
rect 8740 19018 8774 19052
rect 8812 19018 8846 19052
rect 8884 19018 8918 19052
rect 8956 19018 8990 19052
rect 9028 19018 9062 19052
rect 9100 19018 9134 19052
rect 9172 19018 9206 19052
rect 9244 19018 9278 19052
rect 8596 18945 8630 18979
rect 8668 18973 8696 18979
rect 8696 18973 8702 18979
rect 8668 18945 8702 18973
rect 8740 18945 8774 18979
rect 8812 18973 8832 18979
rect 8832 18973 8846 18979
rect 8812 18945 8846 18973
rect 8884 18945 8918 18979
rect 8956 18973 8968 18979
rect 8968 18973 8990 18979
rect 8956 18945 8990 18973
rect 9028 18945 9062 18979
rect 9100 18973 9104 18979
rect 9104 18973 9134 18979
rect 9100 18945 9134 18973
rect 9172 18945 9206 18979
rect 9244 18973 9274 18979
rect 9274 18973 9278 18979
rect 9244 18945 9278 18973
rect 8596 18872 8630 18906
rect 8668 18872 8702 18906
rect 8740 18872 8774 18906
rect 8812 18872 8846 18906
rect 8884 18872 8918 18906
rect 8956 18872 8990 18906
rect 9028 18872 9062 18906
rect 9100 18872 9134 18906
rect 9172 18872 9206 18906
rect 9244 18872 9278 18906
rect 8596 18799 8630 18833
rect 8668 18799 8702 18833
rect 8740 18799 8774 18833
rect 8812 18799 8846 18833
rect 8884 18799 8918 18833
rect 8956 18799 8990 18833
rect 9028 18799 9062 18833
rect 9100 18799 9134 18833
rect 9172 18799 9206 18833
rect 9244 18799 9278 18833
rect 8596 18726 8630 18760
rect 8668 18735 8702 18760
rect 8668 18726 8696 18735
rect 8696 18726 8702 18735
rect 8740 18726 8774 18760
rect 8812 18735 8846 18760
rect 8812 18726 8832 18735
rect 8832 18726 8846 18735
rect 8884 18726 8918 18760
rect 8956 18735 8990 18760
rect 8956 18726 8968 18735
rect 8968 18726 8990 18735
rect 9028 18726 9062 18760
rect 9100 18735 9134 18760
rect 9100 18726 9104 18735
rect 9104 18726 9134 18735
rect 9172 18726 9206 18760
rect 9244 18735 9278 18760
rect 9244 18726 9274 18735
rect 9274 18726 9278 18735
rect 8596 18653 8630 18687
rect 8668 18653 8702 18687
rect 8740 18653 8774 18687
rect 8812 18653 8846 18687
rect 8884 18653 8918 18687
rect 8956 18653 8990 18687
rect 9028 18653 9062 18687
rect 9100 18653 9134 18687
rect 9172 18653 9206 18687
rect 9244 18653 9278 18687
rect 8596 18580 8630 18614
rect 8668 18599 8702 18614
rect 8668 18580 8696 18599
rect 8696 18580 8702 18599
rect 8740 18580 8774 18614
rect 8812 18599 8846 18614
rect 8812 18580 8832 18599
rect 8832 18580 8846 18599
rect 8884 18580 8918 18614
rect 8956 18599 8990 18614
rect 8956 18580 8968 18599
rect 8968 18580 8990 18599
rect 9028 18580 9062 18614
rect 9100 18599 9134 18614
rect 9100 18580 9104 18599
rect 9104 18580 9134 18599
rect 9172 18580 9206 18614
rect 9244 18599 9278 18614
rect 9244 18580 9274 18599
rect 9274 18580 9278 18599
rect 8596 18507 8630 18541
rect 8668 18507 8702 18541
rect 8740 18507 8774 18541
rect 8812 18507 8846 18541
rect 8884 18507 8918 18541
rect 8956 18507 8990 18541
rect 9028 18507 9062 18541
rect 9100 18507 9134 18541
rect 9172 18507 9206 18541
rect 9244 18507 9278 18541
rect 8596 18434 8630 18468
rect 8668 18463 8702 18468
rect 8668 18434 8696 18463
rect 8696 18434 8702 18463
rect 8740 18434 8774 18468
rect 8812 18463 8846 18468
rect 8812 18434 8832 18463
rect 8832 18434 8846 18463
rect 8884 18434 8918 18468
rect 8956 18463 8990 18468
rect 8956 18434 8968 18463
rect 8968 18434 8990 18463
rect 9028 18434 9062 18468
rect 9100 18463 9134 18468
rect 9100 18434 9104 18463
rect 9104 18434 9134 18463
rect 9172 18434 9206 18468
rect 9244 18463 9278 18468
rect 9244 18434 9274 18463
rect 9274 18434 9278 18463
rect 8596 18361 8630 18395
rect 8668 18361 8702 18395
rect 8740 18361 8774 18395
rect 8812 18361 8846 18395
rect 8884 18361 8918 18395
rect 8956 18361 8990 18395
rect 9028 18361 9062 18395
rect 9100 18361 9134 18395
rect 9172 18361 9206 18395
rect 9244 18361 9278 18395
rect 8596 18288 8630 18322
rect 8668 18293 8696 18322
rect 8696 18293 8702 18322
rect 8668 18288 8702 18293
rect 8740 18288 8774 18322
rect 8812 18293 8832 18322
rect 8832 18293 8846 18322
rect 8812 18288 8846 18293
rect 8884 18288 8918 18322
rect 8956 18293 8968 18322
rect 8968 18293 8990 18322
rect 8956 18288 8990 18293
rect 9028 18288 9062 18322
rect 9100 18293 9104 18322
rect 9104 18293 9134 18322
rect 9100 18288 9134 18293
rect 9172 18288 9206 18322
rect 9244 18293 9274 18322
rect 9274 18293 9278 18322
rect 9244 18288 9278 18293
rect 8596 18215 8630 18249
rect 8668 18215 8702 18249
rect 8740 18215 8774 18249
rect 8812 18215 8846 18249
rect 8884 18215 8918 18249
rect 8956 18215 8990 18249
rect 9028 18215 9062 18249
rect 9100 18215 9134 18249
rect 9172 18215 9206 18249
rect 9244 18215 9278 18249
rect 8596 18142 8630 18176
rect 8668 18157 8696 18176
rect 8696 18157 8702 18176
rect 8668 18142 8702 18157
rect 8740 18142 8774 18176
rect 8812 18157 8832 18176
rect 8832 18157 8846 18176
rect 8812 18142 8846 18157
rect 8884 18142 8918 18176
rect 8956 18157 8968 18176
rect 8968 18157 8990 18176
rect 8956 18142 8990 18157
rect 9028 18142 9062 18176
rect 9100 18157 9104 18176
rect 9104 18157 9134 18176
rect 9100 18142 9134 18157
rect 9172 18142 9206 18176
rect 9244 18157 9274 18176
rect 9274 18157 9278 18176
rect 9244 18142 9278 18157
rect 8596 18069 8630 18103
rect 8668 18069 8702 18103
rect 8740 18069 8774 18103
rect 8812 18069 8846 18103
rect 8884 18069 8918 18103
rect 8956 18069 8990 18103
rect 9028 18069 9062 18103
rect 9100 18069 9134 18103
rect 9172 18069 9206 18103
rect 9244 18069 9278 18103
rect 8596 17996 8630 18030
rect 8668 18021 8696 18030
rect 8696 18021 8702 18030
rect 8668 17996 8702 18021
rect 8740 17996 8774 18030
rect 8812 18021 8832 18030
rect 8832 18021 8846 18030
rect 8812 17996 8846 18021
rect 8884 17996 8918 18030
rect 8956 18021 8968 18030
rect 8968 18021 8990 18030
rect 8956 17996 8990 18021
rect 9028 17996 9062 18030
rect 9100 18021 9104 18030
rect 9104 18021 9134 18030
rect 9100 17996 9134 18021
rect 9172 17996 9206 18030
rect 9244 18021 9274 18030
rect 9274 18021 9278 18030
rect 9244 17996 9278 18021
rect 8596 17923 8630 17957
rect 8668 17923 8702 17957
rect 8740 17923 8774 17957
rect 8812 17923 8846 17957
rect 8884 17923 8918 17957
rect 8956 17923 8990 17957
rect 9028 17923 9062 17957
rect 9100 17923 9134 17957
rect 9172 17923 9206 17957
rect 9244 17923 9278 17957
rect 8596 17850 8630 17884
rect 8668 17850 8702 17884
rect 8740 17850 8774 17884
rect 8812 17850 8846 17884
rect 8884 17850 8918 17884
rect 8956 17850 8990 17884
rect 9028 17850 9062 17884
rect 9100 17850 9134 17884
rect 9172 17850 9206 17884
rect 9244 17850 9278 17884
rect 8596 17777 8630 17811
rect 8668 17783 8702 17811
rect 8668 17777 8696 17783
rect 8696 17777 8702 17783
rect 8740 17777 8774 17811
rect 8812 17783 8846 17811
rect 8812 17777 8832 17783
rect 8832 17777 8846 17783
rect 8884 17777 8918 17811
rect 8956 17783 8990 17811
rect 8956 17777 8968 17783
rect 8968 17777 8990 17783
rect 9028 17777 9062 17811
rect 9100 17783 9134 17811
rect 9100 17777 9104 17783
rect 9104 17777 9134 17783
rect 9172 17777 9206 17811
rect 9244 17783 9278 17811
rect 9244 17777 9274 17783
rect 9274 17777 9278 17783
rect 8596 17704 8630 17738
rect 8668 17704 8702 17738
rect 8740 17704 8774 17738
rect 8812 17704 8846 17738
rect 8884 17704 8918 17738
rect 8956 17704 8990 17738
rect 9028 17704 9062 17738
rect 9100 17704 9134 17738
rect 9172 17704 9206 17738
rect 9244 17704 9278 17738
rect 321 17477 325 17511
rect 325 17477 359 17511
rect 359 17477 461 17511
rect 461 17477 495 17511
rect 495 17477 597 17511
rect 597 17477 631 17511
rect 631 17477 733 17511
rect 733 17477 767 17511
rect 767 17477 869 17511
rect 869 17477 903 17511
rect 903 17477 1003 17511
rect 321 17375 1003 17477
rect 321 17341 325 17375
rect 325 17341 359 17375
rect 359 17341 461 17375
rect 461 17341 495 17375
rect 495 17341 597 17375
rect 597 17341 631 17375
rect 631 17341 733 17375
rect 733 17341 767 17375
rect 767 17341 869 17375
rect 869 17341 903 17375
rect 903 17341 1003 17375
rect 321 17239 1003 17341
rect 321 17205 325 17239
rect 325 17205 359 17239
rect 359 17205 461 17239
rect 461 17205 495 17239
rect 495 17205 597 17239
rect 597 17205 631 17239
rect 631 17205 733 17239
rect 733 17205 767 17239
rect 767 17205 869 17239
rect 869 17205 903 17239
rect 903 17205 1003 17239
rect 321 17103 1003 17205
rect 321 17069 325 17103
rect 325 17069 359 17103
rect 359 17069 461 17103
rect 461 17069 495 17103
rect 495 17069 597 17103
rect 597 17069 631 17103
rect 631 17069 733 17103
rect 733 17069 767 17103
rect 767 17069 869 17103
rect 869 17069 903 17103
rect 903 17069 1003 17103
rect 321 16967 1003 17069
rect 321 16933 325 16967
rect 325 16933 359 16967
rect 359 16933 461 16967
rect 461 16933 495 16967
rect 495 16933 597 16967
rect 597 16933 631 16967
rect 631 16933 733 16967
rect 733 16933 767 16967
rect 767 16933 869 16967
rect 869 16933 903 16967
rect 903 16933 1003 16967
rect 321 16831 1003 16933
rect 321 16797 325 16831
rect 325 16797 359 16831
rect 359 16797 461 16831
rect 461 16797 495 16831
rect 495 16797 597 16831
rect 597 16797 631 16831
rect 631 16797 733 16831
rect 733 16797 767 16831
rect 767 16797 869 16831
rect 869 16797 903 16831
rect 903 16797 1003 16831
rect 321 16695 1003 16797
rect 321 16661 325 16695
rect 325 16661 359 16695
rect 359 16661 461 16695
rect 461 16661 495 16695
rect 495 16661 597 16695
rect 597 16661 631 16695
rect 631 16661 733 16695
rect 733 16661 767 16695
rect 767 16661 869 16695
rect 869 16661 903 16695
rect 903 16661 1003 16695
rect 321 16559 1003 16661
rect 321 16525 325 16559
rect 325 16525 359 16559
rect 359 16525 461 16559
rect 461 16525 495 16559
rect 495 16525 597 16559
rect 597 16525 631 16559
rect 631 16525 733 16559
rect 733 16525 767 16559
rect 767 16525 869 16559
rect 869 16525 903 16559
rect 903 16525 1003 16559
rect 321 16423 1003 16525
rect 321 16389 325 16423
rect 325 16389 359 16423
rect 359 16389 461 16423
rect 461 16389 495 16423
rect 495 16389 597 16423
rect 597 16389 631 16423
rect 631 16389 733 16423
rect 733 16389 767 16423
rect 767 16389 869 16423
rect 869 16389 903 16423
rect 903 16389 1003 16423
rect 321 16287 1003 16389
rect 321 16253 325 16287
rect 325 16253 359 16287
rect 359 16253 461 16287
rect 461 16253 495 16287
rect 495 16253 597 16287
rect 597 16253 631 16287
rect 631 16253 733 16287
rect 733 16253 767 16287
rect 767 16253 869 16287
rect 869 16253 903 16287
rect 903 16253 1003 16287
rect 321 16151 1003 16253
rect 321 16117 325 16151
rect 325 16117 359 16151
rect 359 16117 461 16151
rect 461 16117 495 16151
rect 495 16117 597 16151
rect 597 16117 631 16151
rect 631 16117 733 16151
rect 733 16117 767 16151
rect 767 16117 869 16151
rect 869 16117 903 16151
rect 903 16117 1003 16151
rect 321 16015 1003 16117
rect 321 15981 325 16015
rect 325 15981 359 16015
rect 359 15981 461 16015
rect 461 15981 495 16015
rect 495 15981 597 16015
rect 597 15981 631 16015
rect 631 15981 733 16015
rect 733 15981 767 16015
rect 767 15981 869 16015
rect 869 15981 903 16015
rect 903 15981 1003 16015
rect 321 15879 1003 15981
rect 321 15845 325 15879
rect 325 15845 359 15879
rect 359 15845 461 15879
rect 461 15845 495 15879
rect 495 15845 597 15879
rect 597 15845 631 15879
rect 631 15845 733 15879
rect 733 15845 767 15879
rect 767 15845 869 15879
rect 869 15845 903 15879
rect 903 15845 1003 15879
rect 321 15743 1003 15845
rect 321 15709 325 15743
rect 325 15709 359 15743
rect 359 15709 461 15743
rect 461 15709 495 15743
rect 495 15709 597 15743
rect 597 15709 631 15743
rect 631 15709 733 15743
rect 733 15709 767 15743
rect 767 15709 869 15743
rect 869 15709 903 15743
rect 903 15709 1003 15743
rect 321 15607 1003 15709
rect 321 15573 325 15607
rect 325 15573 359 15607
rect 359 15573 461 15607
rect 461 15573 495 15607
rect 495 15573 597 15607
rect 597 15573 631 15607
rect 631 15573 733 15607
rect 733 15573 767 15607
rect 767 15573 869 15607
rect 869 15573 903 15607
rect 903 15573 1003 15607
rect 321 15471 1003 15573
rect 321 15437 325 15471
rect 325 15437 359 15471
rect 359 15437 461 15471
rect 461 15437 495 15471
rect 495 15437 597 15471
rect 597 15437 631 15471
rect 631 15437 733 15471
rect 733 15437 767 15471
rect 767 15437 869 15471
rect 869 15437 903 15471
rect 903 15437 1003 15471
rect 321 15335 1003 15437
rect 321 15301 325 15335
rect 325 15301 359 15335
rect 359 15301 461 15335
rect 461 15301 495 15335
rect 495 15301 597 15335
rect 597 15301 631 15335
rect 631 15301 733 15335
rect 733 15301 767 15335
rect 767 15301 869 15335
rect 869 15301 903 15335
rect 903 15301 1003 15335
rect 321 15199 1003 15301
rect 321 15165 325 15199
rect 325 15165 359 15199
rect 359 15165 461 15199
rect 461 15165 495 15199
rect 495 15165 597 15199
rect 597 15165 631 15199
rect 631 15165 733 15199
rect 733 15165 767 15199
rect 767 15165 869 15199
rect 869 15165 903 15199
rect 903 15165 1003 15199
rect 321 15063 1003 15165
rect 321 15029 325 15063
rect 325 15029 359 15063
rect 359 15029 461 15063
rect 461 15029 495 15063
rect 495 15029 597 15063
rect 597 15029 631 15063
rect 631 15029 733 15063
rect 733 15029 767 15063
rect 767 15029 869 15063
rect 869 15029 903 15063
rect 903 15029 1003 15063
rect 321 14927 1003 15029
rect 321 14893 325 14927
rect 325 14893 359 14927
rect 359 14893 461 14927
rect 461 14893 495 14927
rect 495 14893 597 14927
rect 597 14893 631 14927
rect 631 14893 733 14927
rect 733 14893 767 14927
rect 767 14893 869 14927
rect 869 14893 903 14927
rect 903 14893 1003 14927
rect 321 14791 1003 14893
rect 321 14757 325 14791
rect 325 14757 359 14791
rect 359 14757 461 14791
rect 461 14757 495 14791
rect 495 14757 597 14791
rect 597 14757 631 14791
rect 631 14757 733 14791
rect 733 14757 767 14791
rect 767 14757 869 14791
rect 869 14757 903 14791
rect 903 14757 1003 14791
rect 321 14655 1003 14757
rect 321 14621 325 14655
rect 325 14621 359 14655
rect 359 14621 461 14655
rect 461 14621 495 14655
rect 495 14621 597 14655
rect 597 14621 631 14655
rect 631 14621 733 14655
rect 733 14621 767 14655
rect 767 14621 869 14655
rect 869 14621 903 14655
rect 903 14621 1003 14655
rect 321 14519 1003 14621
rect 321 14485 325 14519
rect 325 14485 359 14519
rect 359 14485 461 14519
rect 461 14485 495 14519
rect 495 14485 597 14519
rect 597 14485 631 14519
rect 631 14485 733 14519
rect 733 14485 767 14519
rect 767 14485 869 14519
rect 869 14485 903 14519
rect 903 14485 1003 14519
rect 321 14383 1003 14485
rect 321 14349 325 14383
rect 325 14349 359 14383
rect 359 14349 461 14383
rect 461 14349 495 14383
rect 495 14349 597 14383
rect 597 14349 631 14383
rect 631 14349 733 14383
rect 733 14349 767 14383
rect 767 14349 869 14383
rect 869 14349 903 14383
rect 903 14349 1003 14383
rect 321 14247 1003 14349
rect 321 14213 325 14247
rect 325 14213 359 14247
rect 359 14213 461 14247
rect 461 14213 495 14247
rect 495 14213 597 14247
rect 597 14213 631 14247
rect 631 14213 733 14247
rect 733 14213 767 14247
rect 767 14213 869 14247
rect 869 14213 903 14247
rect 903 14213 1003 14247
rect 321 14111 1003 14213
rect 321 14077 325 14111
rect 325 14077 359 14111
rect 359 14077 461 14111
rect 461 14077 495 14111
rect 495 14077 597 14111
rect 597 14077 631 14111
rect 631 14077 733 14111
rect 733 14077 767 14111
rect 767 14077 869 14111
rect 869 14077 903 14111
rect 903 14077 1003 14111
rect 321 13975 1003 14077
rect 321 13941 325 13975
rect 325 13941 359 13975
rect 359 13941 461 13975
rect 461 13941 495 13975
rect 495 13941 597 13975
rect 597 13941 631 13975
rect 631 13941 733 13975
rect 733 13941 767 13975
rect 767 13941 869 13975
rect 869 13941 903 13975
rect 903 13941 1003 13975
rect 321 13839 1003 13941
rect 321 13805 325 13839
rect 325 13805 359 13839
rect 359 13805 461 13839
rect 461 13805 495 13839
rect 495 13805 597 13839
rect 597 13805 631 13839
rect 631 13805 733 13839
rect 733 13805 767 13839
rect 767 13805 869 13839
rect 869 13805 903 13839
rect 903 13805 1003 13839
rect 321 13703 1003 13805
rect 321 13669 325 13703
rect 325 13669 359 13703
rect 359 13669 461 13703
rect 461 13669 495 13703
rect 495 13669 597 13703
rect 597 13669 631 13703
rect 631 13669 733 13703
rect 733 13669 767 13703
rect 767 13669 869 13703
rect 869 13669 903 13703
rect 903 13669 1003 13703
rect 321 13567 1003 13669
rect 321 13533 325 13567
rect 325 13533 359 13567
rect 359 13533 461 13567
rect 461 13533 495 13567
rect 495 13533 597 13567
rect 597 13533 631 13567
rect 631 13533 733 13567
rect 733 13533 767 13567
rect 767 13533 869 13567
rect 869 13533 903 13567
rect 903 13533 1003 13567
rect 321 13431 1003 13533
rect 321 13397 325 13431
rect 325 13397 359 13431
rect 359 13397 461 13431
rect 461 13397 495 13431
rect 495 13397 597 13431
rect 597 13397 631 13431
rect 631 13397 733 13431
rect 733 13397 767 13431
rect 767 13397 869 13431
rect 869 13397 903 13431
rect 903 13397 1003 13431
rect 321 13295 1003 13397
rect 321 13261 325 13295
rect 325 13261 359 13295
rect 359 13261 461 13295
rect 461 13261 495 13295
rect 495 13261 597 13295
rect 597 13261 631 13295
rect 631 13261 733 13295
rect 733 13261 767 13295
rect 767 13261 869 13295
rect 869 13261 903 13295
rect 903 13261 1003 13295
rect 321 13159 1003 13261
rect 321 13125 325 13159
rect 325 13125 359 13159
rect 359 13125 461 13159
rect 461 13125 495 13159
rect 495 13125 597 13159
rect 597 13125 631 13159
rect 631 13125 733 13159
rect 733 13125 767 13159
rect 767 13125 869 13159
rect 869 13125 903 13159
rect 903 13125 1003 13159
rect 321 13023 1003 13125
rect 321 12989 325 13023
rect 325 12989 359 13023
rect 359 12989 461 13023
rect 461 12989 495 13023
rect 495 12989 597 13023
rect 597 12989 631 13023
rect 631 12989 733 13023
rect 733 12989 767 13023
rect 767 12989 869 13023
rect 869 12989 903 13023
rect 903 12989 1003 13023
rect 321 12887 1003 12989
rect 321 12853 325 12887
rect 325 12853 359 12887
rect 359 12853 461 12887
rect 461 12853 495 12887
rect 495 12853 597 12887
rect 597 12853 631 12887
rect 631 12853 733 12887
rect 733 12853 767 12887
rect 767 12853 869 12887
rect 869 12853 903 12887
rect 903 12853 1003 12887
rect 321 12751 1003 12853
rect 321 12717 325 12751
rect 325 12717 359 12751
rect 359 12717 461 12751
rect 461 12717 495 12751
rect 495 12717 597 12751
rect 597 12717 631 12751
rect 631 12717 733 12751
rect 733 12717 767 12751
rect 767 12717 869 12751
rect 869 12717 903 12751
rect 903 12717 1003 12751
rect 321 12615 1003 12717
rect 321 12581 325 12615
rect 325 12581 359 12615
rect 359 12581 461 12615
rect 461 12581 495 12615
rect 495 12581 597 12615
rect 597 12581 631 12615
rect 631 12581 733 12615
rect 733 12581 767 12615
rect 767 12581 869 12615
rect 869 12581 903 12615
rect 903 12581 1003 12615
rect 321 12479 1003 12581
rect 321 12445 325 12479
rect 325 12445 359 12479
rect 359 12445 461 12479
rect 461 12445 495 12479
rect 495 12445 597 12479
rect 597 12445 631 12479
rect 631 12445 733 12479
rect 733 12445 767 12479
rect 767 12445 869 12479
rect 869 12445 903 12479
rect 903 12445 1003 12479
rect 321 12343 1003 12445
rect 321 12309 325 12343
rect 325 12309 359 12343
rect 359 12309 461 12343
rect 461 12309 495 12343
rect 495 12309 597 12343
rect 597 12309 631 12343
rect 631 12309 733 12343
rect 733 12309 767 12343
rect 767 12309 869 12343
rect 869 12309 903 12343
rect 903 12309 1003 12343
rect 321 12207 1003 12309
rect 321 12173 325 12207
rect 325 12173 359 12207
rect 359 12173 461 12207
rect 461 12173 495 12207
rect 495 12173 597 12207
rect 597 12173 631 12207
rect 631 12173 733 12207
rect 733 12173 767 12207
rect 767 12173 869 12207
rect 869 12173 903 12207
rect 903 12173 1003 12207
rect 321 12071 1003 12173
rect 321 12037 325 12071
rect 325 12037 359 12071
rect 359 12037 461 12071
rect 461 12037 495 12071
rect 495 12037 597 12071
rect 597 12037 631 12071
rect 631 12037 733 12071
rect 733 12037 767 12071
rect 767 12037 869 12071
rect 869 12037 903 12071
rect 903 12037 1003 12071
rect 321 11935 1003 12037
rect 321 11901 325 11935
rect 325 11901 359 11935
rect 359 11901 461 11935
rect 461 11901 495 11935
rect 495 11901 597 11935
rect 597 11901 631 11935
rect 631 11901 733 11935
rect 733 11901 767 11935
rect 767 11901 869 11935
rect 869 11901 903 11935
rect 903 11901 1003 11935
rect 321 11799 1003 11901
rect 321 11765 325 11799
rect 325 11765 359 11799
rect 359 11765 461 11799
rect 461 11765 495 11799
rect 495 11765 597 11799
rect 597 11765 631 11799
rect 631 11765 733 11799
rect 733 11765 767 11799
rect 767 11765 869 11799
rect 869 11765 903 11799
rect 903 11765 1003 11799
rect 321 11663 1003 11765
rect 321 11629 325 11663
rect 325 11629 359 11663
rect 359 11629 461 11663
rect 461 11629 495 11663
rect 495 11629 597 11663
rect 597 11629 631 11663
rect 631 11629 733 11663
rect 733 11629 767 11663
rect 767 11629 869 11663
rect 869 11629 903 11663
rect 903 11629 1003 11663
rect 321 11527 1003 11629
rect 321 11493 325 11527
rect 325 11493 359 11527
rect 359 11493 461 11527
rect 461 11493 495 11527
rect 495 11493 597 11527
rect 597 11493 631 11527
rect 631 11493 733 11527
rect 733 11493 767 11527
rect 767 11493 869 11527
rect 869 11493 903 11527
rect 903 11493 1003 11527
rect 321 11391 1003 11493
rect 321 11357 325 11391
rect 325 11357 359 11391
rect 359 11357 461 11391
rect 461 11357 495 11391
rect 495 11357 597 11391
rect 597 11357 631 11391
rect 631 11357 733 11391
rect 733 11357 767 11391
rect 767 11357 869 11391
rect 869 11357 903 11391
rect 903 11357 1003 11391
rect 321 11255 1003 11357
rect 321 11221 325 11255
rect 325 11221 359 11255
rect 359 11221 461 11255
rect 461 11221 495 11255
rect 495 11221 597 11255
rect 597 11221 631 11255
rect 631 11221 733 11255
rect 733 11221 767 11255
rect 767 11221 869 11255
rect 869 11221 903 11255
rect 903 11221 1003 11255
rect 321 11119 1003 11221
rect 321 11085 325 11119
rect 325 11085 359 11119
rect 359 11085 461 11119
rect 461 11085 495 11119
rect 495 11085 597 11119
rect 597 11085 631 11119
rect 631 11085 733 11119
rect 733 11085 767 11119
rect 767 11085 869 11119
rect 869 11085 903 11119
rect 903 11085 1003 11119
rect 321 10983 1003 11085
rect 321 10949 325 10983
rect 325 10949 359 10983
rect 359 10949 461 10983
rect 461 10949 495 10983
rect 495 10949 597 10983
rect 597 10949 631 10983
rect 631 10949 733 10983
rect 733 10949 767 10983
rect 767 10949 869 10983
rect 869 10949 903 10983
rect 903 10949 1003 10983
rect 321 10847 1003 10949
rect 321 10813 325 10847
rect 325 10813 359 10847
rect 359 10813 461 10847
rect 461 10813 495 10847
rect 495 10813 597 10847
rect 597 10813 631 10847
rect 631 10813 733 10847
rect 733 10813 767 10847
rect 767 10813 869 10847
rect 869 10813 903 10847
rect 903 10813 1003 10847
rect 321 10711 1003 10813
rect 321 10677 325 10711
rect 325 10677 359 10711
rect 359 10677 461 10711
rect 461 10677 495 10711
rect 495 10677 597 10711
rect 597 10677 631 10711
rect 631 10677 733 10711
rect 733 10677 767 10711
rect 767 10677 869 10711
rect 869 10677 903 10711
rect 903 10677 1003 10711
rect 321 10575 1003 10677
rect 321 10541 325 10575
rect 325 10541 359 10575
rect 359 10541 461 10575
rect 461 10541 495 10575
rect 495 10541 597 10575
rect 597 10541 631 10575
rect 631 10541 733 10575
rect 733 10541 767 10575
rect 767 10541 869 10575
rect 869 10541 903 10575
rect 903 10541 1003 10575
rect 321 10439 1003 10541
rect 321 10405 325 10439
rect 325 10405 359 10439
rect 359 10405 461 10439
rect 461 10405 495 10439
rect 495 10405 597 10439
rect 597 10405 631 10439
rect 631 10405 733 10439
rect 733 10405 767 10439
rect 767 10405 869 10439
rect 869 10405 903 10439
rect 903 10405 1003 10439
rect 321 10303 1003 10405
rect 321 10269 325 10303
rect 325 10269 359 10303
rect 359 10269 461 10303
rect 461 10269 495 10303
rect 495 10269 597 10303
rect 597 10269 631 10303
rect 631 10269 733 10303
rect 733 10269 767 10303
rect 767 10269 869 10303
rect 869 10269 903 10303
rect 903 10269 1003 10303
rect 321 10167 1003 10269
rect 321 10133 325 10167
rect 325 10133 359 10167
rect 359 10133 461 10167
rect 461 10133 495 10167
rect 495 10133 597 10167
rect 597 10133 631 10167
rect 631 10133 733 10167
rect 733 10133 767 10167
rect 767 10133 869 10167
rect 869 10133 903 10167
rect 903 10133 1003 10167
rect 321 10031 1003 10133
rect 321 9997 325 10031
rect 325 9997 359 10031
rect 359 9997 461 10031
rect 461 9997 495 10031
rect 495 9997 597 10031
rect 597 9997 631 10031
rect 631 9997 733 10031
rect 733 9997 767 10031
rect 767 9997 869 10031
rect 869 9997 903 10031
rect 903 9997 1003 10031
rect 321 9895 1003 9997
rect 321 9861 325 9895
rect 325 9861 359 9895
rect 359 9861 461 9895
rect 461 9861 495 9895
rect 495 9861 597 9895
rect 597 9861 631 9895
rect 631 9861 733 9895
rect 733 9861 767 9895
rect 767 9861 869 9895
rect 869 9861 903 9895
rect 903 9861 1003 9895
rect 321 9759 1003 9861
rect 321 9725 325 9759
rect 325 9725 359 9759
rect 359 9725 461 9759
rect 461 9725 495 9759
rect 495 9725 597 9759
rect 597 9725 631 9759
rect 631 9725 733 9759
rect 733 9725 767 9759
rect 767 9725 869 9759
rect 869 9725 903 9759
rect 903 9725 1003 9759
rect 321 9623 1003 9725
rect 321 9589 325 9623
rect 325 9589 359 9623
rect 359 9589 461 9623
rect 461 9589 495 9623
rect 495 9589 597 9623
rect 597 9589 631 9623
rect 631 9589 733 9623
rect 733 9589 767 9623
rect 767 9589 869 9623
rect 869 9589 903 9623
rect 903 9589 1003 9623
rect 321 9487 1003 9589
rect 321 9453 325 9487
rect 325 9453 359 9487
rect 359 9453 461 9487
rect 461 9453 495 9487
rect 495 9453 597 9487
rect 597 9453 631 9487
rect 631 9453 733 9487
rect 733 9453 767 9487
rect 767 9453 869 9487
rect 869 9453 903 9487
rect 903 9453 1003 9487
rect 321 9351 1003 9453
rect 321 9317 325 9351
rect 325 9317 359 9351
rect 359 9317 461 9351
rect 461 9317 495 9351
rect 495 9317 597 9351
rect 597 9317 631 9351
rect 631 9317 733 9351
rect 733 9317 767 9351
rect 767 9317 869 9351
rect 869 9317 903 9351
rect 903 9317 1003 9351
rect 321 9215 1003 9317
rect 321 9181 325 9215
rect 325 9181 359 9215
rect 359 9181 461 9215
rect 461 9181 495 9215
rect 495 9181 597 9215
rect 597 9181 631 9215
rect 631 9181 733 9215
rect 733 9181 767 9215
rect 767 9181 869 9215
rect 869 9181 903 9215
rect 903 9181 1003 9215
rect 321 9079 1003 9181
rect 321 9045 325 9079
rect 325 9045 359 9079
rect 359 9045 461 9079
rect 461 9045 495 9079
rect 495 9045 597 9079
rect 597 9045 631 9079
rect 631 9045 733 9079
rect 733 9045 767 9079
rect 767 9045 869 9079
rect 869 9045 903 9079
rect 903 9045 1003 9079
rect 321 8943 1003 9045
rect 321 8909 325 8943
rect 325 8909 359 8943
rect 359 8909 461 8943
rect 461 8909 495 8943
rect 495 8909 597 8943
rect 597 8909 631 8943
rect 631 8909 733 8943
rect 733 8909 767 8943
rect 767 8909 869 8943
rect 869 8909 903 8943
rect 903 8909 1003 8943
rect 321 8807 1003 8909
rect 321 8773 325 8807
rect 325 8773 359 8807
rect 359 8773 461 8807
rect 461 8773 495 8807
rect 495 8773 597 8807
rect 597 8773 631 8807
rect 631 8773 733 8807
rect 733 8773 767 8807
rect 767 8773 869 8807
rect 869 8773 903 8807
rect 903 8773 1003 8807
rect 321 8671 1003 8773
rect 321 8637 325 8671
rect 325 8637 359 8671
rect 359 8637 461 8671
rect 461 8637 495 8671
rect 495 8637 597 8671
rect 597 8637 631 8671
rect 631 8637 733 8671
rect 733 8637 767 8671
rect 767 8637 869 8671
rect 869 8637 903 8671
rect 903 8637 1003 8671
rect 321 8535 1003 8637
rect 321 8501 325 8535
rect 325 8501 359 8535
rect 359 8501 461 8535
rect 461 8501 495 8535
rect 495 8501 597 8535
rect 597 8501 631 8535
rect 631 8501 733 8535
rect 733 8501 767 8535
rect 767 8501 869 8535
rect 869 8501 903 8535
rect 903 8501 1003 8535
rect 321 8399 1003 8501
rect 321 8365 325 8399
rect 325 8365 359 8399
rect 359 8365 461 8399
rect 461 8365 495 8399
rect 495 8365 597 8399
rect 597 8365 631 8399
rect 631 8365 733 8399
rect 733 8365 767 8399
rect 767 8365 869 8399
rect 869 8365 903 8399
rect 903 8365 1003 8399
rect 321 8263 1003 8365
rect 321 8229 325 8263
rect 325 8229 359 8263
rect 359 8229 461 8263
rect 461 8229 495 8263
rect 495 8229 597 8263
rect 597 8229 631 8263
rect 631 8229 733 8263
rect 733 8229 767 8263
rect 767 8229 869 8263
rect 869 8229 903 8263
rect 903 8229 1003 8263
rect 321 8127 1003 8229
rect 321 8093 325 8127
rect 325 8093 359 8127
rect 359 8093 461 8127
rect 461 8093 495 8127
rect 495 8093 597 8127
rect 597 8093 631 8127
rect 631 8093 733 8127
rect 733 8093 767 8127
rect 767 8093 869 8127
rect 869 8093 903 8127
rect 903 8093 1003 8127
rect 321 7991 1003 8093
rect 321 7957 325 7991
rect 325 7957 359 7991
rect 359 7957 461 7991
rect 461 7957 495 7991
rect 495 7957 597 7991
rect 597 7957 631 7991
rect 631 7957 733 7991
rect 733 7957 767 7991
rect 767 7957 869 7991
rect 869 7957 903 7991
rect 903 7957 1003 7991
rect 321 7855 1003 7957
rect 321 7821 325 7855
rect 325 7821 359 7855
rect 359 7821 461 7855
rect 461 7821 495 7855
rect 495 7821 597 7855
rect 597 7821 631 7855
rect 631 7821 733 7855
rect 733 7821 767 7855
rect 767 7821 869 7855
rect 869 7821 903 7855
rect 903 7821 1003 7855
rect 321 7719 1003 7821
rect 321 7685 325 7719
rect 325 7685 359 7719
rect 359 7685 461 7719
rect 461 7685 495 7719
rect 495 7685 597 7719
rect 597 7685 631 7719
rect 631 7685 733 7719
rect 733 7685 767 7719
rect 767 7685 869 7719
rect 869 7685 903 7719
rect 903 7685 1003 7719
rect 321 7583 1003 7685
rect 321 7549 325 7583
rect 325 7549 359 7583
rect 359 7549 461 7583
rect 461 7549 495 7583
rect 495 7549 597 7583
rect 597 7549 631 7583
rect 631 7549 733 7583
rect 733 7549 767 7583
rect 767 7549 869 7583
rect 869 7549 903 7583
rect 903 7549 1003 7583
rect 321 7447 1003 7549
rect 321 7413 325 7447
rect 325 7413 359 7447
rect 359 7413 461 7447
rect 461 7413 495 7447
rect 495 7413 597 7447
rect 597 7413 631 7447
rect 631 7413 733 7447
rect 733 7413 767 7447
rect 767 7413 869 7447
rect 869 7413 903 7447
rect 903 7413 1003 7447
rect 321 7311 1003 7413
rect 321 7277 325 7311
rect 325 7277 359 7311
rect 359 7277 461 7311
rect 461 7277 495 7311
rect 495 7277 597 7311
rect 597 7277 631 7311
rect 631 7277 733 7311
rect 733 7277 767 7311
rect 767 7277 869 7311
rect 869 7277 903 7311
rect 903 7277 1003 7311
rect 321 7175 1003 7277
rect 321 7141 325 7175
rect 325 7141 359 7175
rect 359 7141 461 7175
rect 461 7141 495 7175
rect 495 7141 597 7175
rect 597 7141 631 7175
rect 631 7141 733 7175
rect 733 7141 767 7175
rect 767 7141 869 7175
rect 869 7141 903 7175
rect 903 7141 1003 7175
rect 321 7039 1003 7141
rect 321 7005 325 7039
rect 325 7005 359 7039
rect 359 7005 461 7039
rect 461 7005 495 7039
rect 495 7005 597 7039
rect 597 7005 631 7039
rect 631 7005 733 7039
rect 733 7005 767 7039
rect 767 7005 869 7039
rect 869 7005 903 7039
rect 903 7005 1003 7039
rect 321 6903 1003 7005
rect 321 6869 325 6903
rect 325 6869 359 6903
rect 359 6869 461 6903
rect 461 6869 495 6903
rect 495 6869 597 6903
rect 597 6869 631 6903
rect 631 6869 733 6903
rect 733 6869 767 6903
rect 767 6869 869 6903
rect 869 6869 903 6903
rect 903 6869 1003 6903
rect 321 6767 1003 6869
rect 321 6733 325 6767
rect 325 6733 359 6767
rect 359 6733 461 6767
rect 461 6733 495 6767
rect 495 6733 597 6767
rect 597 6733 631 6767
rect 631 6733 733 6767
rect 733 6733 767 6767
rect 767 6733 869 6767
rect 869 6733 903 6767
rect 903 6733 1003 6767
rect 321 6631 1003 6733
rect 321 6597 325 6631
rect 325 6597 359 6631
rect 359 6597 461 6631
rect 461 6597 495 6631
rect 495 6597 597 6631
rect 597 6597 631 6631
rect 631 6597 733 6631
rect 733 6597 767 6631
rect 767 6597 869 6631
rect 869 6597 903 6631
rect 903 6597 1003 6631
rect 321 6495 1003 6597
rect 321 6461 325 6495
rect 325 6461 359 6495
rect 359 6461 461 6495
rect 461 6461 495 6495
rect 495 6461 597 6495
rect 597 6461 631 6495
rect 631 6461 733 6495
rect 733 6461 767 6495
rect 767 6461 869 6495
rect 869 6461 903 6495
rect 903 6461 1003 6495
rect 321 6359 1003 6461
rect 321 6325 325 6359
rect 325 6325 359 6359
rect 359 6325 461 6359
rect 461 6325 495 6359
rect 495 6325 597 6359
rect 597 6325 631 6359
rect 631 6325 733 6359
rect 733 6325 767 6359
rect 767 6325 869 6359
rect 869 6325 903 6359
rect 903 6325 1003 6359
rect 321 6223 1003 6325
rect 321 6189 325 6223
rect 325 6189 359 6223
rect 359 6189 461 6223
rect 461 6189 495 6223
rect 495 6189 597 6223
rect 597 6189 631 6223
rect 631 6189 733 6223
rect 733 6189 767 6223
rect 767 6189 869 6223
rect 869 6189 903 6223
rect 903 6189 1003 6223
rect 321 6087 1003 6189
rect 321 6053 325 6087
rect 325 6053 359 6087
rect 359 6053 461 6087
rect 461 6053 495 6087
rect 495 6053 597 6087
rect 597 6053 631 6087
rect 631 6053 733 6087
rect 733 6053 767 6087
rect 767 6053 869 6087
rect 869 6053 903 6087
rect 903 6053 1003 6087
rect 321 5951 1003 6053
rect 321 5917 325 5951
rect 325 5917 359 5951
rect 359 5917 461 5951
rect 461 5917 495 5951
rect 495 5917 597 5951
rect 597 5917 631 5951
rect 631 5917 733 5951
rect 733 5917 767 5951
rect 767 5917 869 5951
rect 869 5917 903 5951
rect 903 5917 1003 5951
rect 321 5815 1003 5917
rect 321 5781 325 5815
rect 325 5781 359 5815
rect 359 5781 461 5815
rect 461 5781 495 5815
rect 495 5781 597 5815
rect 597 5781 631 5815
rect 631 5781 733 5815
rect 733 5781 767 5815
rect 767 5781 869 5815
rect 869 5781 903 5815
rect 903 5781 1003 5815
rect 321 5679 1003 5781
rect 321 5645 325 5679
rect 325 5645 359 5679
rect 359 5645 461 5679
rect 461 5645 495 5679
rect 495 5645 597 5679
rect 597 5645 631 5679
rect 631 5645 733 5679
rect 733 5645 767 5679
rect 767 5645 869 5679
rect 869 5645 903 5679
rect 903 5645 1003 5679
rect 321 5543 1003 5645
rect 321 5509 325 5543
rect 325 5509 359 5543
rect 359 5509 461 5543
rect 461 5509 495 5543
rect 495 5509 597 5543
rect 597 5509 631 5543
rect 631 5509 733 5543
rect 733 5509 767 5543
rect 767 5509 869 5543
rect 869 5509 903 5543
rect 903 5509 1003 5543
rect 321 5407 1003 5509
rect 321 5373 325 5407
rect 325 5373 359 5407
rect 359 5373 461 5407
rect 461 5373 495 5407
rect 495 5373 597 5407
rect 597 5373 631 5407
rect 631 5373 733 5407
rect 733 5373 767 5407
rect 767 5373 869 5407
rect 869 5373 903 5407
rect 903 5373 1003 5407
rect 321 5271 1003 5373
rect 321 5237 325 5271
rect 325 5237 359 5271
rect 359 5237 461 5271
rect 461 5237 495 5271
rect 495 5237 597 5271
rect 597 5237 631 5271
rect 631 5237 733 5271
rect 733 5237 767 5271
rect 767 5237 869 5271
rect 869 5237 903 5271
rect 903 5237 1003 5271
rect 321 5135 1003 5237
rect 321 5101 325 5135
rect 325 5101 359 5135
rect 359 5101 461 5135
rect 461 5101 495 5135
rect 495 5101 597 5135
rect 597 5101 631 5135
rect 631 5101 733 5135
rect 733 5101 767 5135
rect 767 5101 869 5135
rect 869 5101 903 5135
rect 903 5101 1003 5135
rect 321 4999 1003 5101
rect 321 4965 325 4999
rect 325 4965 359 4999
rect 359 4965 461 4999
rect 461 4965 495 4999
rect 495 4965 597 4999
rect 597 4965 631 4999
rect 631 4965 733 4999
rect 733 4965 767 4999
rect 767 4965 869 4999
rect 869 4965 903 4999
rect 903 4965 1003 4999
rect 321 4863 1003 4965
rect 321 4829 325 4863
rect 325 4829 359 4863
rect 359 4829 461 4863
rect 461 4829 495 4863
rect 495 4829 597 4863
rect 597 4829 631 4863
rect 631 4829 733 4863
rect 733 4829 767 4863
rect 767 4829 869 4863
rect 869 4829 903 4863
rect 903 4829 1003 4863
rect 321 4727 1003 4829
rect 321 4693 325 4727
rect 325 4693 359 4727
rect 359 4693 461 4727
rect 461 4693 495 4727
rect 495 4693 597 4727
rect 597 4693 631 4727
rect 631 4693 733 4727
rect 733 4693 767 4727
rect 767 4693 869 4727
rect 869 4693 903 4727
rect 903 4693 1003 4727
rect 321 4591 1003 4693
rect 321 4557 325 4591
rect 325 4557 359 4591
rect 359 4557 461 4591
rect 461 4557 495 4591
rect 495 4557 597 4591
rect 597 4557 631 4591
rect 631 4557 733 4591
rect 733 4557 767 4591
rect 767 4557 869 4591
rect 869 4557 903 4591
rect 903 4557 1003 4591
rect 321 4455 1003 4557
rect 321 4421 325 4455
rect 325 4421 359 4455
rect 359 4421 461 4455
rect 461 4421 495 4455
rect 495 4421 597 4455
rect 597 4421 631 4455
rect 631 4421 733 4455
rect 733 4421 767 4455
rect 767 4421 869 4455
rect 869 4421 903 4455
rect 903 4421 1003 4455
rect 321 4319 1003 4421
rect 321 4285 325 4319
rect 325 4285 359 4319
rect 359 4285 461 4319
rect 461 4285 495 4319
rect 495 4285 597 4319
rect 597 4285 631 4319
rect 631 4285 733 4319
rect 733 4285 767 4319
rect 767 4285 869 4319
rect 869 4285 903 4319
rect 903 4285 1003 4319
rect 321 4183 1003 4285
rect 321 4149 325 4183
rect 325 4149 359 4183
rect 359 4149 461 4183
rect 461 4149 495 4183
rect 495 4149 597 4183
rect 597 4149 631 4183
rect 631 4149 733 4183
rect 733 4149 767 4183
rect 767 4149 869 4183
rect 869 4149 903 4183
rect 903 4149 1003 4183
rect 321 4047 1003 4149
rect 321 4013 325 4047
rect 325 4013 359 4047
rect 359 4013 461 4047
rect 461 4013 495 4047
rect 495 4013 597 4047
rect 597 4013 631 4047
rect 631 4013 733 4047
rect 733 4013 767 4047
rect 767 4013 869 4047
rect 869 4013 903 4047
rect 903 4013 1003 4047
rect 321 3911 1003 4013
rect 321 3877 325 3911
rect 325 3877 359 3911
rect 359 3877 461 3911
rect 461 3877 495 3911
rect 495 3877 597 3911
rect 597 3877 631 3911
rect 631 3877 733 3911
rect 733 3877 767 3911
rect 767 3877 869 3911
rect 869 3877 903 3911
rect 903 3877 1003 3911
rect 321 3775 1003 3877
rect 321 3741 325 3775
rect 325 3741 359 3775
rect 359 3741 461 3775
rect 461 3741 495 3775
rect 495 3741 597 3775
rect 597 3741 631 3775
rect 631 3741 733 3775
rect 733 3741 767 3775
rect 767 3741 869 3775
rect 869 3741 903 3775
rect 903 3741 1003 3775
rect 321 3639 1003 3741
rect 321 3605 325 3639
rect 325 3605 359 3639
rect 359 3605 461 3639
rect 461 3605 495 3639
rect 495 3605 597 3639
rect 597 3605 631 3639
rect 631 3605 733 3639
rect 733 3605 767 3639
rect 767 3605 869 3639
rect 869 3605 903 3639
rect 903 3605 1003 3639
rect 321 3503 1003 3605
rect 321 3469 325 3503
rect 325 3469 359 3503
rect 359 3469 461 3503
rect 461 3469 495 3503
rect 495 3469 597 3503
rect 597 3469 631 3503
rect 631 3469 733 3503
rect 733 3469 767 3503
rect 767 3469 869 3503
rect 869 3469 903 3503
rect 903 3469 1003 3503
rect 321 3367 1003 3469
rect 321 3333 325 3367
rect 325 3333 359 3367
rect 359 3333 461 3367
rect 461 3333 495 3367
rect 495 3333 597 3367
rect 597 3333 631 3367
rect 631 3333 733 3367
rect 733 3333 767 3367
rect 767 3333 869 3367
rect 869 3333 903 3367
rect 903 3333 1003 3367
rect 321 3231 1003 3333
rect 321 3197 325 3231
rect 325 3197 359 3231
rect 359 3197 461 3231
rect 461 3197 495 3231
rect 495 3197 597 3231
rect 597 3197 631 3231
rect 631 3197 733 3231
rect 733 3197 767 3231
rect 767 3197 869 3231
rect 869 3197 903 3231
rect 903 3197 1003 3231
rect 321 3125 1003 3197
rect 321 3061 325 3086
rect 325 3061 355 3086
rect 321 3052 355 3061
rect 393 3052 427 3086
rect 465 3061 495 3086
rect 495 3061 499 3086
rect 465 3052 499 3061
rect 537 3052 571 3086
rect 609 3061 631 3086
rect 631 3061 643 3086
rect 609 3052 643 3061
rect 681 3052 715 3086
rect 753 3061 767 3086
rect 767 3061 787 3086
rect 753 3052 787 3061
rect 825 3052 859 3086
rect 897 3061 903 3086
rect 903 3061 931 3086
rect 897 3052 931 3061
rect 969 3052 1003 3086
rect 321 2979 355 3013
rect 393 2979 427 3013
rect 465 2979 499 3013
rect 537 2979 571 3013
rect 609 2979 643 3013
rect 681 2979 715 3013
rect 753 2979 787 3013
rect 825 2979 859 3013
rect 897 2979 931 3013
rect 969 2979 1003 3013
rect 321 2925 325 2940
rect 325 2925 355 2940
rect 321 2906 355 2925
rect 393 2906 427 2940
rect 465 2925 495 2940
rect 495 2925 499 2940
rect 465 2906 499 2925
rect 537 2906 571 2940
rect 609 2925 631 2940
rect 631 2925 643 2940
rect 609 2906 643 2925
rect 681 2906 715 2940
rect 753 2925 767 2940
rect 767 2925 787 2940
rect 753 2906 787 2925
rect 825 2906 859 2940
rect 897 2925 903 2940
rect 903 2925 931 2940
rect 897 2906 931 2925
rect 969 2906 1003 2940
rect 321 2833 355 2867
rect 393 2833 427 2867
rect 465 2833 499 2867
rect 537 2833 571 2867
rect 609 2833 643 2867
rect 681 2833 715 2867
rect 753 2833 787 2867
rect 825 2833 859 2867
rect 897 2833 931 2867
rect 969 2833 1003 2867
rect 321 2789 325 2794
rect 325 2789 355 2794
rect 321 2760 355 2789
rect 393 2760 427 2794
rect 465 2789 495 2794
rect 495 2789 499 2794
rect 465 2760 499 2789
rect 537 2760 571 2794
rect 609 2789 631 2794
rect 631 2789 643 2794
rect 609 2760 643 2789
rect 681 2760 715 2794
rect 753 2789 767 2794
rect 767 2789 787 2794
rect 753 2760 787 2789
rect 825 2760 859 2794
rect 897 2789 903 2794
rect 903 2789 931 2794
rect 897 2760 931 2789
rect 969 2760 1003 2794
rect 321 2687 355 2721
rect 393 2687 427 2721
rect 465 2687 499 2721
rect 537 2687 571 2721
rect 609 2687 643 2721
rect 681 2687 715 2721
rect 753 2687 787 2721
rect 825 2687 859 2721
rect 897 2687 931 2721
rect 969 2687 1003 2721
rect 321 2614 355 2648
rect 393 2614 427 2648
rect 465 2614 499 2648
rect 537 2614 571 2648
rect 609 2614 643 2648
rect 681 2614 715 2648
rect 753 2614 787 2648
rect 825 2614 859 2648
rect 897 2614 931 2648
rect 969 2614 1003 2648
rect 321 2551 355 2575
rect 321 2541 325 2551
rect 325 2541 355 2551
rect 393 2541 427 2575
rect 465 2551 499 2575
rect 465 2541 495 2551
rect 495 2541 499 2551
rect 537 2541 571 2575
rect 609 2551 643 2575
rect 609 2541 631 2551
rect 631 2541 643 2551
rect 681 2541 715 2575
rect 753 2551 787 2575
rect 753 2541 767 2551
rect 767 2541 787 2551
rect 825 2541 859 2575
rect 897 2551 931 2575
rect 897 2541 903 2551
rect 903 2541 931 2551
rect 969 2541 1003 2575
rect 321 2468 355 2502
rect 393 2468 427 2502
rect 465 2468 499 2502
rect 537 2468 571 2502
rect 609 2468 643 2502
rect 681 2468 715 2502
rect 753 2468 787 2502
rect 825 2468 859 2502
rect 897 2468 931 2502
rect 969 2468 1003 2502
rect 321 2414 355 2429
rect 321 2395 325 2414
rect 325 2395 355 2414
rect 393 2395 427 2429
rect 465 2414 499 2429
rect 465 2395 495 2414
rect 495 2395 499 2414
rect 537 2395 571 2429
rect 609 2414 643 2429
rect 609 2395 631 2414
rect 631 2395 643 2414
rect 681 2395 715 2429
rect 753 2414 787 2429
rect 753 2395 767 2414
rect 767 2395 787 2414
rect 825 2395 859 2429
rect 897 2414 931 2429
rect 897 2395 903 2414
rect 903 2395 931 2414
rect 969 2395 1003 2429
rect 321 2322 355 2356
rect 393 2322 427 2356
rect 465 2322 499 2356
rect 537 2322 571 2356
rect 609 2322 643 2356
rect 681 2322 715 2356
rect 753 2322 787 2356
rect 825 2322 859 2356
rect 897 2322 931 2356
rect 969 2322 1003 2356
rect 321 2277 355 2283
rect 321 2249 325 2277
rect 325 2249 355 2277
rect 393 2249 427 2283
rect 465 2277 499 2283
rect 465 2249 495 2277
rect 495 2249 499 2277
rect 537 2249 571 2283
rect 609 2277 643 2283
rect 609 2249 631 2277
rect 631 2249 643 2277
rect 681 2249 715 2283
rect 753 2277 787 2283
rect 753 2249 767 2277
rect 767 2249 787 2277
rect 825 2249 859 2283
rect 897 2277 931 2283
rect 897 2249 903 2277
rect 903 2249 931 2277
rect 969 2249 1003 2283
rect 321 2176 355 2210
rect 393 2176 427 2210
rect 465 2176 499 2210
rect 537 2176 571 2210
rect 609 2176 643 2210
rect 681 2176 715 2210
rect 753 2176 787 2210
rect 825 2176 859 2210
rect 897 2176 931 2210
rect 969 2176 1003 2210
rect 321 2106 325 2137
rect 325 2106 355 2137
rect 321 2103 355 2106
rect 393 2103 427 2137
rect 465 2106 495 2137
rect 495 2106 499 2137
rect 465 2103 499 2106
rect 537 2103 571 2137
rect 609 2106 631 2137
rect 631 2106 643 2137
rect 609 2103 643 2106
rect 681 2103 715 2137
rect 753 2106 767 2137
rect 767 2106 787 2137
rect 753 2103 787 2106
rect 825 2103 859 2137
rect 897 2106 903 2137
rect 903 2106 931 2137
rect 897 2103 931 2106
rect 969 2103 1003 2137
rect 321 2030 355 2064
rect 393 2030 427 2064
rect 465 2030 499 2064
rect 537 2030 571 2064
rect 609 2030 643 2064
rect 681 2030 715 2064
rect 753 2030 787 2064
rect 825 2030 859 2064
rect 897 2030 931 2064
rect 969 2030 1003 2064
rect 321 1969 325 1991
rect 325 1969 355 1991
rect 321 1957 355 1969
rect 393 1957 427 1991
rect 465 1969 495 1991
rect 495 1969 499 1991
rect 465 1957 499 1969
rect 537 1957 571 1991
rect 609 1969 631 1991
rect 631 1969 643 1991
rect 609 1957 643 1969
rect 681 1957 715 1991
rect 753 1969 767 1991
rect 767 1969 787 1991
rect 753 1957 787 1969
rect 825 1957 859 1991
rect 897 1969 903 1991
rect 903 1969 931 1991
rect 897 1957 931 1969
rect 969 1957 1003 1991
rect 321 1884 355 1918
rect 393 1884 427 1918
rect 465 1884 499 1918
rect 537 1884 571 1918
rect 609 1884 643 1918
rect 681 1884 715 1918
rect 753 1884 787 1918
rect 825 1884 859 1918
rect 897 1884 931 1918
rect 969 1884 1003 1918
rect 321 1832 325 1845
rect 325 1832 355 1845
rect 321 1811 355 1832
rect 393 1811 427 1845
rect 465 1832 495 1845
rect 495 1832 499 1845
rect 465 1811 499 1832
rect 537 1811 571 1845
rect 609 1832 631 1845
rect 631 1832 643 1845
rect 609 1811 643 1832
rect 681 1811 715 1845
rect 753 1832 767 1845
rect 767 1832 787 1845
rect 753 1811 787 1832
rect 825 1811 859 1845
rect 897 1832 903 1845
rect 903 1832 931 1845
rect 897 1811 931 1832
rect 969 1811 1003 1845
rect 321 1738 355 1772
rect 393 1738 427 1772
rect 465 1738 499 1772
rect 537 1738 571 1772
rect 609 1738 643 1772
rect 681 1738 715 1772
rect 753 1738 787 1772
rect 825 1738 859 1772
rect 897 1738 931 1772
rect 969 1738 1003 1772
rect 321 1695 325 1699
rect 325 1695 355 1699
rect 321 1665 355 1695
rect 393 1665 427 1699
rect 465 1695 495 1699
rect 495 1695 499 1699
rect 465 1665 499 1695
rect 537 1665 571 1699
rect 609 1695 631 1699
rect 631 1695 643 1699
rect 609 1665 643 1695
rect 681 1665 715 1699
rect 753 1695 767 1699
rect 767 1695 787 1699
rect 753 1665 787 1695
rect 825 1665 859 1699
rect 897 1695 903 1699
rect 903 1695 931 1699
rect 897 1665 931 1695
rect 969 1665 1003 1699
rect 5080 16438 5114 16472
rect 5156 16438 5173 16472
rect 5173 16438 5190 16472
rect 5232 16438 5241 16472
rect 5241 16438 5266 16472
rect 5308 16438 5309 16472
rect 5309 16438 5342 16472
rect 5385 16438 5411 16472
rect 5411 16438 5419 16472
rect 5462 16438 5479 16472
rect 5479 16438 5496 16472
rect 5572 16438 5581 16472
rect 5581 16438 5606 16472
rect 5644 16438 5649 16472
rect 5649 16438 5678 16472
rect 5716 16438 5717 16472
rect 5717 16438 5750 16472
rect 5788 16438 5819 16472
rect 5819 16438 5822 16472
rect 5860 16438 5887 16472
rect 5887 16438 5894 16472
rect 5932 16438 5955 16472
rect 5955 16438 5966 16472
rect 6004 16438 6023 16472
rect 6023 16438 6038 16472
rect 6076 16438 6091 16472
rect 6091 16438 6110 16472
rect 6148 16438 6159 16472
rect 6159 16438 6182 16472
rect 6220 16438 6227 16472
rect 6227 16438 6254 16472
rect 6292 16438 6295 16472
rect 6295 16438 6326 16472
rect 6364 16438 6397 16472
rect 6397 16438 6398 16472
rect 6436 16438 6465 16472
rect 6465 16438 6470 16472
rect 6508 16438 6533 16472
rect 6533 16438 6542 16472
rect 6580 16438 6601 16472
rect 6601 16438 6614 16472
rect 6652 16438 6669 16472
rect 6669 16438 6686 16472
rect 6724 16438 6737 16472
rect 6737 16438 6758 16472
rect 6796 16438 6805 16472
rect 6805 16438 6830 16472
rect 6868 16438 6873 16472
rect 6873 16438 6902 16472
rect 6940 16438 6941 16472
rect 6941 16438 6974 16472
rect 7012 16438 7043 16472
rect 7043 16438 7046 16472
rect 7084 16438 7111 16472
rect 7111 16438 7118 16472
rect 7156 16438 7179 16472
rect 7179 16438 7190 16472
rect 7228 16438 7247 16472
rect 7247 16438 7262 16472
rect 7301 16438 7315 16472
rect 7315 16438 7335 16472
rect 7374 16438 7383 16472
rect 7383 16438 7408 16472
rect 7447 16438 7451 16472
rect 7451 16438 7481 16472
rect 5004 16370 5038 16400
rect 5004 16366 5038 16370
rect 5004 16302 5038 16327
rect 5004 16293 5038 16302
rect 5004 16234 5038 16254
rect 5004 16220 5038 16234
rect 5004 16166 5038 16181
rect 5004 16147 5038 16166
rect 5004 16098 5038 16108
rect 5004 16074 5038 16098
rect 5004 16030 5038 16035
rect 5004 16001 5038 16030
rect 5004 15928 5038 15962
rect 5004 15860 5038 15889
rect 5004 15855 5038 15860
rect 5004 15792 5038 15816
rect 5004 15782 5038 15792
rect 5004 15724 5038 15743
rect 5004 15709 5038 15724
rect 5004 15656 5038 15670
rect 5004 15636 5038 15656
rect 5004 15588 5038 15597
rect 5004 15563 5038 15588
rect 5004 15520 5038 15524
rect 5004 15490 5038 15520
rect 5004 15418 5038 15451
rect 5004 15417 5038 15418
rect 5004 15350 5038 15378
rect 5004 15344 5038 15350
rect 5004 15282 5038 15305
rect 5004 15271 5038 15282
rect 5004 15214 5038 15232
rect 5004 15198 5038 15214
rect 5004 15146 5038 15159
rect 5004 15125 5038 15146
rect 5004 15078 5038 15086
rect 5004 15052 5038 15078
rect 5004 15010 5038 15013
rect 5004 14979 5038 15010
rect 5004 14908 5038 14940
rect 5004 14906 5038 14908
rect 5004 14840 5038 14867
rect 5004 14833 5038 14840
rect 5004 14772 5038 14795
rect 5004 14761 5038 14772
rect 5004 14704 5038 14723
rect 5004 14689 5038 14704
rect 5004 14636 5038 14651
rect 5004 14617 5038 14636
rect 5004 14568 5038 14579
rect 5004 14545 5038 14568
rect 5004 14500 5038 14507
rect 5004 14473 5038 14500
rect 5004 14432 5038 14435
rect 5004 14401 5038 14432
rect 5004 14330 5038 14363
rect 5004 14329 5038 14330
rect 5004 14262 5038 14291
rect 5004 14257 5038 14262
rect 5004 14194 5038 14219
rect 5004 14185 5038 14194
rect 5004 14126 5038 14147
rect 5004 14113 5038 14126
rect 5004 14058 5038 14075
rect 5004 14041 5038 14058
rect 5004 13990 5038 14003
rect 5004 13969 5038 13990
rect 5004 13922 5038 13931
rect 5004 13897 5038 13922
rect 5004 13854 5038 13859
rect 5004 13825 5038 13854
rect 5004 13786 5038 13787
rect 5004 13753 5038 13786
rect 5004 13684 5038 13715
rect 5004 13681 5038 13684
rect 5004 13616 5038 13643
rect 5004 13609 5038 13616
rect 5004 13548 5038 13571
rect 5004 13537 5038 13548
rect 5004 13480 5038 13499
rect 5004 13465 5038 13480
rect 5004 13412 5038 13427
rect 5004 13393 5038 13412
rect 5004 13344 5038 13355
rect 5004 13321 5038 13344
rect 5004 13276 5038 13283
rect 5004 13249 5038 13276
rect 5004 13208 5038 13211
rect 5004 13177 5038 13208
rect 5004 13106 5038 13139
rect 5004 13105 5038 13106
rect 5004 13038 5038 13067
rect 5004 13033 5038 13038
rect 5004 12970 5038 12995
rect 5004 12961 5038 12970
rect 5004 12902 5038 12923
rect 5004 12889 5038 12902
rect 5004 12834 5038 12851
rect 5004 12817 5038 12834
rect 5004 12766 5038 12779
rect 5004 12745 5038 12766
rect 5004 12698 5038 12707
rect 5004 12673 5038 12698
rect 5004 12630 5038 12635
rect 5004 12601 5038 12630
rect 5004 12562 5038 12563
rect 5004 12529 5038 12562
rect 5004 12460 5038 12491
rect 5004 12457 5038 12460
rect 5004 12392 5038 12419
rect 5004 12385 5038 12392
rect 5004 12324 5038 12347
rect 5004 12313 5038 12324
rect 5004 12256 5038 12275
rect 5004 12241 5038 12256
rect 5004 12188 5038 12203
rect 5004 12169 5038 12188
rect 5004 12120 5038 12131
rect 5004 12097 5038 12120
rect 5004 12052 5038 12059
rect 5004 12025 5038 12052
rect 5004 11984 5038 11987
rect 5004 11953 5038 11984
rect 5004 11882 5038 11915
rect 5004 11881 5038 11882
rect 5004 11814 5038 11843
rect 5004 11809 5038 11814
rect 5004 11746 5038 11771
rect 5004 11737 5038 11746
rect 5004 11678 5038 11699
rect 5004 11665 5038 11678
rect 5004 11610 5038 11627
rect 5004 11593 5038 11610
rect 5004 11542 5038 11555
rect 5004 11521 5038 11542
rect 5004 11474 5038 11483
rect 5004 11449 5038 11474
rect 5004 11406 5038 11411
rect 5004 11377 5038 11406
rect 5004 11338 5038 11339
rect 5004 11305 5038 11338
rect 5004 11236 5038 11267
rect 5004 11233 5038 11236
rect 5004 11168 5038 11195
rect 5004 11161 5038 11168
rect 5004 11100 5038 11123
rect 5004 11089 5038 11100
rect 5004 11032 5038 11051
rect 5004 11017 5038 11032
rect 5004 10964 5038 10979
rect 5004 10945 5038 10964
rect 5004 10896 5038 10907
rect 5004 10873 5038 10896
rect 5004 10828 5038 10835
rect 5004 10801 5038 10828
rect 5004 10760 5038 10763
rect 5004 10729 5038 10760
rect 5004 10658 5038 10691
rect 5004 10657 5038 10658
rect 5004 10590 5038 10619
rect 5004 10585 5038 10590
rect 5004 10522 5038 10547
rect 5004 10513 5038 10522
rect 5004 10454 5038 10475
rect 5004 10441 5038 10454
rect 5004 10386 5038 10403
rect 5004 10369 5038 10386
rect 5004 10318 5038 10331
rect 5004 10297 5038 10318
rect 5004 10250 5038 10259
rect 5004 10225 5038 10250
rect 5004 10182 5038 10187
rect 5004 10153 5038 10182
rect 5004 10114 5038 10115
rect 5004 10081 5038 10114
rect 5004 10012 5038 10043
rect 5004 10009 5038 10012
rect 5004 9944 5038 9971
rect 5004 9937 5038 9944
rect 5004 9876 5038 9899
rect 5004 9865 5038 9876
rect 5004 9808 5038 9827
rect 5004 9793 5038 9808
rect 5004 9740 5038 9755
rect 5004 9721 5038 9740
rect 5004 9672 5038 9683
rect 5004 9649 5038 9672
rect 5004 9604 5038 9611
rect 5004 9577 5038 9604
rect 5004 9536 5038 9539
rect 5004 9505 5038 9536
rect 5004 9434 5038 9467
rect 5004 9433 5038 9434
rect 5004 9366 5038 9395
rect 5004 9361 5038 9366
rect 5004 9298 5038 9323
rect 5004 9289 5038 9298
rect 5004 9230 5038 9251
rect 5004 9217 5038 9230
rect 5004 9162 5038 9179
rect 5004 9145 5038 9162
rect 5004 9094 5038 9107
rect 5004 9073 5038 9094
rect 5004 9026 5038 9035
rect 5004 9001 5038 9026
rect 5004 8958 5038 8963
rect 5004 8929 5038 8958
rect 5004 8890 5038 8891
rect 5004 8857 5038 8890
rect 5004 8788 5038 8819
rect 5004 8785 5038 8788
rect 5004 8720 5038 8747
rect 5004 8713 5038 8720
rect 5004 8652 5038 8675
rect 5004 8641 5038 8652
rect 5004 8584 5038 8603
rect 5004 8569 5038 8584
rect 5004 8516 5038 8531
rect 5004 8497 5038 8516
rect 5004 8448 5038 8459
rect 5004 8425 5038 8448
rect 5004 8380 5038 8387
rect 5004 8353 5038 8380
rect 5004 8312 5038 8315
rect 5004 8281 5038 8312
rect 5004 8210 5038 8243
rect 5004 8209 5038 8210
rect 5004 8142 5038 8171
rect 5004 8137 5038 8142
rect 5004 8074 5038 8099
rect 5004 8065 5038 8074
rect 5004 8006 5038 8027
rect 5004 7993 5038 8006
rect 5004 7938 5038 7955
rect 5004 7921 5038 7938
rect 5004 7870 5038 7883
rect 5004 7849 5038 7870
rect 5004 7802 5038 7811
rect 5004 7777 5038 7802
rect 5004 7734 5038 7739
rect 5004 7705 5038 7734
rect 5004 7666 5038 7667
rect 5004 7633 5038 7666
rect 5004 7564 5038 7595
rect 5004 7561 5038 7564
rect 5004 7496 5038 7523
rect 5004 7489 5038 7496
rect 5004 7428 5038 7451
rect 5004 7417 5038 7428
rect 5004 7360 5038 7379
rect 5004 7345 5038 7360
rect 5004 7292 5038 7307
rect 5004 7273 5038 7292
rect 5004 7224 5038 7235
rect 5004 7201 5038 7224
rect 5004 7156 5038 7163
rect 5004 7129 5038 7156
rect 5004 7088 5038 7091
rect 5004 7057 5038 7088
rect 5004 6986 5038 7019
rect 5004 6985 5038 6986
rect 5004 6918 5038 6947
rect 5004 6913 5038 6918
rect 5004 6850 5038 6875
rect 5004 6841 5038 6850
rect 5004 6782 5038 6803
rect 5004 6769 5038 6782
rect 5004 6714 5038 6731
rect 5004 6697 5038 6714
rect 5004 6646 5038 6659
rect 5004 6625 5038 6646
rect 5004 6578 5038 6587
rect 5004 6553 5038 6578
rect 5004 6510 5038 6515
rect 5004 6481 5038 6510
rect 5004 6442 5038 6443
rect 5004 6409 5038 6442
rect 5004 6340 5038 6371
rect 5004 6337 5038 6340
rect 5004 6272 5038 6299
rect 5004 6265 5038 6272
rect 5004 6204 5038 6227
rect 5004 6193 5038 6204
rect 5004 6136 5038 6155
rect 5004 6121 5038 6136
rect 5004 6068 5038 6083
rect 5004 6049 5038 6068
rect 5004 6000 5038 6011
rect 5004 5977 5038 6000
rect 5004 5932 5038 5939
rect 5004 5905 5038 5932
rect 5004 5864 5038 5867
rect 5004 5833 5038 5864
rect 5004 5762 5038 5795
rect 5004 5761 5038 5762
rect 5004 5694 5038 5723
rect 5004 5689 5038 5694
rect 5004 5626 5038 5651
rect 5004 5617 5038 5626
rect 5004 5558 5038 5579
rect 5004 5545 5038 5558
rect 5004 5490 5038 5507
rect 5004 5473 5038 5490
rect 5004 5422 5038 5435
rect 5004 5401 5038 5422
rect 5004 5354 5038 5363
rect 5004 5329 5038 5354
rect 5004 5286 5038 5291
rect 5004 5257 5038 5286
rect 5004 5218 5038 5219
rect 5004 5185 5038 5218
rect 5004 5116 5038 5147
rect 5004 5113 5038 5116
rect 5004 5048 5038 5075
rect 5004 5041 5038 5048
rect 5004 4980 5038 5003
rect 5004 4969 5038 4980
rect 5004 4912 5038 4931
rect 5004 4897 5038 4912
rect 5004 4844 5038 4859
rect 5004 4825 5038 4844
rect 5004 4776 5038 4787
rect 5004 4753 5038 4776
rect 5004 4708 5038 4715
rect 5004 4681 5038 4708
rect 5004 4640 5038 4643
rect 5004 4609 5038 4640
rect 5004 4538 5038 4571
rect 5004 4537 5038 4538
rect 5004 4470 5038 4499
rect 5004 4465 5038 4470
rect 5004 4402 5038 4427
rect 5004 4393 5038 4402
rect 5004 4334 5038 4355
rect 5004 4321 5038 4334
rect 5004 4266 5038 4283
rect 5004 4249 5038 4266
rect 5004 4198 5038 4211
rect 5004 4177 5038 4198
rect 5004 4130 5038 4139
rect 5004 4105 5038 4130
rect 5004 4062 5038 4067
rect 5004 4033 5038 4062
rect 5004 3994 5038 3995
rect 5004 3961 5038 3994
rect 5004 3892 5038 3923
rect 5004 3889 5038 3892
rect 5004 3824 5038 3851
rect 5004 3817 5038 3824
rect 5004 3756 5038 3779
rect 5004 3745 5038 3756
rect 5004 3688 5038 3707
rect 5004 3673 5038 3688
rect 5004 3620 5038 3635
rect 5004 3601 5038 3620
rect 5004 3552 5038 3563
rect 5004 3529 5038 3552
rect 5004 3484 5038 3491
rect 5004 3457 5038 3484
rect 5004 3416 5038 3419
rect 5004 3385 5038 3416
rect 5004 3314 5038 3347
rect 5004 3313 5038 3314
rect 5004 3246 5038 3275
rect 5004 3241 5038 3246
rect 5004 3178 5038 3203
rect 5004 3169 5038 3178
rect 5004 3110 5038 3131
rect 5004 3097 5038 3110
rect 5004 3042 5038 3059
rect 5004 3025 5038 3042
rect 5004 2974 5038 2987
rect 5004 2953 5038 2974
rect 5004 2906 5038 2915
rect 5004 2881 5038 2906
rect 5004 2838 5038 2843
rect 5004 2809 5038 2838
rect 5004 2770 5038 2771
rect 5004 2737 5038 2770
rect 5004 2668 5038 2699
rect 5004 2665 5038 2668
rect 5004 2600 5038 2627
rect 5004 2593 5038 2600
rect 5004 2532 5038 2555
rect 5004 2521 5038 2532
rect 5004 2464 5038 2483
rect 5004 2449 5038 2464
rect 5004 2396 5038 2411
rect 5004 2377 5038 2396
rect 5004 2328 5038 2339
rect 5004 2305 5038 2328
rect 5004 2260 5038 2267
rect 5004 2233 5038 2260
rect 5004 2192 5038 2195
rect 5004 2161 5038 2192
rect 5004 2090 5038 2123
rect 5004 2089 5038 2090
rect 5004 2022 5038 2051
rect 5004 2017 5038 2022
rect 5004 1954 5038 1979
rect 5004 1945 5038 1954
rect 5004 1873 5038 1907
rect 5004 1821 5038 1835
rect 5004 1801 5038 1821
rect 7519 16383 7553 16400
rect 7519 16366 7553 16383
rect 7519 16315 7553 16328
rect 7519 16294 7553 16315
rect 7519 16247 7553 16256
rect 7519 16222 7553 16247
rect 7519 16179 7553 16184
rect 7519 16150 7553 16179
rect 7519 16111 7553 16112
rect 7519 16078 7553 16111
rect 7519 16009 7553 16040
rect 7519 16006 7553 16009
rect 7519 15941 7553 15968
rect 7519 15934 7553 15941
rect 7519 15873 7553 15896
rect 7519 15862 7553 15873
rect 7519 15805 7553 15824
rect 7519 15790 7553 15805
rect 7519 15737 7553 15752
rect 7519 15718 7553 15737
rect 7519 15669 7553 15680
rect 7519 15646 7553 15669
rect 7519 15601 7553 15608
rect 7519 15574 7553 15601
rect 7519 15533 7553 15536
rect 7519 15502 7553 15533
rect 7519 15431 7553 15464
rect 7519 15430 7553 15431
rect 7519 15363 7553 15392
rect 7519 15358 7553 15363
rect 7519 15295 7553 15320
rect 7519 15286 7553 15295
rect 7519 15227 7553 15248
rect 7519 15214 7553 15227
rect 7519 15159 7553 15176
rect 7519 15142 7553 15159
rect 7519 15091 7553 15104
rect 7519 15070 7553 15091
rect 7519 15023 7553 15032
rect 7519 14998 7553 15023
rect 7519 14955 7553 14960
rect 7519 14926 7553 14955
rect 7519 14887 7553 14888
rect 7519 14854 7553 14887
rect 7519 14785 7553 14816
rect 7519 14782 7553 14785
rect 7519 14717 7553 14744
rect 7519 14710 7553 14717
rect 7519 14649 7553 14672
rect 7519 14638 7553 14649
rect 7519 14581 7553 14600
rect 7519 14566 7553 14581
rect 7519 14513 7553 14528
rect 7519 14494 7553 14513
rect 7519 14445 7553 14456
rect 7519 14422 7553 14445
rect 7519 14377 7553 14384
rect 7519 14350 7553 14377
rect 7519 14309 7553 14312
rect 7519 14278 7553 14309
rect 7519 14207 7553 14240
rect 7519 14206 7553 14207
rect 7519 14139 7553 14168
rect 7519 14134 7553 14139
rect 7519 14071 7553 14096
rect 7519 14062 7553 14071
rect 7519 14003 7553 14024
rect 7519 13990 7553 14003
rect 7519 13935 7553 13952
rect 7519 13918 7553 13935
rect 7519 13867 7553 13880
rect 7519 13846 7553 13867
rect 7519 13799 7553 13808
rect 7519 13774 7553 13799
rect 7519 13731 7553 13736
rect 7519 13702 7553 13731
rect 7519 13663 7553 13664
rect 7519 13630 7553 13663
rect 7519 13561 7553 13592
rect 7519 13558 7553 13561
rect 7519 13493 7553 13520
rect 7519 13486 7553 13493
rect 7519 13425 7553 13448
rect 7519 13414 7553 13425
rect 7519 13357 7553 13376
rect 7519 13342 7553 13357
rect 7519 13289 7553 13304
rect 7519 13270 7553 13289
rect 7519 13221 7553 13232
rect 7519 13198 7553 13221
rect 7519 13153 7553 13160
rect 7519 13126 7553 13153
rect 7519 13085 7553 13088
rect 7519 13054 7553 13085
rect 7519 12983 7553 13016
rect 7519 12982 7553 12983
rect 7519 12915 7553 12944
rect 7519 12910 7553 12915
rect 7519 12847 7553 12872
rect 7519 12838 7553 12847
rect 7519 12779 7553 12800
rect 7519 12766 7553 12779
rect 7519 12711 7553 12728
rect 7519 12694 7553 12711
rect 7519 12643 7553 12656
rect 7519 12622 7553 12643
rect 7519 12575 7553 12584
rect 7519 12550 7553 12575
rect 7519 12507 7553 12512
rect 7519 12478 7553 12507
rect 7519 12439 7553 12440
rect 7519 12406 7553 12439
rect 7519 12337 7553 12368
rect 7519 12334 7553 12337
rect 7519 12269 7553 12296
rect 7519 12262 7553 12269
rect 7519 12201 7553 12224
rect 7519 12190 7553 12201
rect 7519 12133 7553 12152
rect 7519 12118 7553 12133
rect 7519 12065 7553 12080
rect 7519 12046 7553 12065
rect 7519 11997 7553 12008
rect 7519 11974 7553 11997
rect 7519 11929 7553 11936
rect 7519 11902 7553 11929
rect 7519 11861 7553 11864
rect 7519 11830 7553 11861
rect 7519 11759 7553 11792
rect 7519 11758 7553 11759
rect 7519 11691 7553 11720
rect 7519 11686 7553 11691
rect 7519 11623 7553 11648
rect 7519 11614 7553 11623
rect 7519 11555 7553 11576
rect 7519 11542 7553 11555
rect 7519 11487 7553 11504
rect 7519 11470 7553 11487
rect 7519 11419 7553 11432
rect 7519 11398 7553 11419
rect 7519 11351 7553 11360
rect 7519 11326 7553 11351
rect 7519 11283 7553 11288
rect 7519 11254 7553 11283
rect 7519 11215 7553 11216
rect 7519 11182 7553 11215
rect 7519 11113 7553 11144
rect 7519 11110 7553 11113
rect 7519 11045 7553 11072
rect 7519 11038 7553 11045
rect 7519 10977 7553 11000
rect 7519 10966 7553 10977
rect 7519 10909 7553 10928
rect 7519 10894 7553 10909
rect 7519 10841 7553 10856
rect 7519 10822 7553 10841
rect 7519 10773 7553 10784
rect 7519 10750 7553 10773
rect 7519 10705 7553 10712
rect 7519 10678 7553 10705
rect 7519 10637 7553 10640
rect 7519 10606 7553 10637
rect 7519 10535 7553 10568
rect 7519 10534 7553 10535
rect 7519 10467 7553 10496
rect 7519 10462 7553 10467
rect 7519 10399 7553 10424
rect 7519 10390 7553 10399
rect 7519 10331 7553 10352
rect 7519 10318 7553 10331
rect 7519 10263 7553 10280
rect 7519 10246 7553 10263
rect 7519 10195 7553 10208
rect 7519 10174 7553 10195
rect 7519 10127 7553 10136
rect 7519 10102 7553 10127
rect 7519 10059 7553 10064
rect 7519 10030 7553 10059
rect 7519 9991 7553 9992
rect 7519 9958 7553 9991
rect 7519 9889 7553 9920
rect 7519 9886 7553 9889
rect 7519 9821 7553 9848
rect 7519 9814 7553 9821
rect 7519 9753 7553 9776
rect 7519 9742 7553 9753
rect 7519 9685 7553 9704
rect 7519 9670 7553 9685
rect 7519 9617 7553 9632
rect 7519 9598 7553 9617
rect 7519 9549 7553 9560
rect 7519 9526 7553 9549
rect 7519 9481 7553 9488
rect 7519 9454 7553 9481
rect 7519 9413 7553 9416
rect 7519 9382 7553 9413
rect 7519 9311 7553 9344
rect 7519 9310 7553 9311
rect 7519 9243 7553 9272
rect 7519 9238 7553 9243
rect 7519 9175 7553 9200
rect 7519 9166 7553 9175
rect 7519 9107 7553 9128
rect 7519 9094 7553 9107
rect 7519 9039 7553 9056
rect 7519 9022 7553 9039
rect 7519 8971 7553 8984
rect 7519 8950 7553 8971
rect 7519 8903 7553 8912
rect 7519 8878 7553 8903
rect 7519 8835 7553 8840
rect 7519 8806 7553 8835
rect 7519 8767 7553 8768
rect 7519 8734 7553 8767
rect 7519 8665 7553 8696
rect 7519 8662 7553 8665
rect 7519 8597 7553 8624
rect 7519 8590 7553 8597
rect 7519 8529 7553 8552
rect 7519 8518 7553 8529
rect 7519 8461 7553 8480
rect 7519 8446 7553 8461
rect 7519 8393 7553 8408
rect 7519 8374 7553 8393
rect 7519 8325 7553 8336
rect 7519 8302 7553 8325
rect 7519 8257 7553 8264
rect 7519 8230 7553 8257
rect 7519 8189 7553 8192
rect 7519 8158 7553 8189
rect 7519 8087 7553 8120
rect 7519 8086 7553 8087
rect 7519 8019 7553 8048
rect 7519 8014 7553 8019
rect 7519 7951 7553 7976
rect 7519 7942 7553 7951
rect 7519 7883 7553 7904
rect 7519 7870 7553 7883
rect 7519 7815 7553 7832
rect 7519 7798 7553 7815
rect 7519 7747 7553 7760
rect 7519 7726 7553 7747
rect 7519 7679 7553 7688
rect 7519 7654 7553 7679
rect 7519 7611 7553 7616
rect 7519 7582 7553 7611
rect 7519 7543 7553 7544
rect 7519 7510 7553 7543
rect 7519 7441 7553 7472
rect 7519 7438 7553 7441
rect 7519 7373 7553 7400
rect 7519 7366 7553 7373
rect 7519 7305 7553 7328
rect 7519 7294 7553 7305
rect 7519 7237 7553 7256
rect 7519 7222 7553 7237
rect 7519 7169 7553 7184
rect 7519 7150 7553 7169
rect 7519 7101 7553 7112
rect 7519 7078 7553 7101
rect 7519 7033 7553 7040
rect 7519 7006 7553 7033
rect 7519 6965 7553 6968
rect 7519 6934 7553 6965
rect 7519 6863 7553 6896
rect 7519 6862 7553 6863
rect 7519 6795 7553 6824
rect 7519 6790 7553 6795
rect 7519 6727 7553 6752
rect 7519 6718 7553 6727
rect 7519 6659 7553 6680
rect 7519 6646 7553 6659
rect 7519 6591 7553 6608
rect 7519 6574 7553 6591
rect 7519 6523 7553 6536
rect 7519 6502 7553 6523
rect 7519 6455 7553 6464
rect 7519 6430 7553 6455
rect 7519 6387 7553 6392
rect 7519 6358 7553 6387
rect 7519 6319 7553 6320
rect 7519 6286 7553 6319
rect 7519 6217 7553 6248
rect 7519 6214 7553 6217
rect 7519 6149 7553 6176
rect 7519 6142 7553 6149
rect 7519 6081 7553 6104
rect 7519 6070 7553 6081
rect 7519 6013 7553 6032
rect 7519 5998 7553 6013
rect 7519 5945 7553 5960
rect 7519 5926 7553 5945
rect 7519 5877 7553 5888
rect 7519 5854 7553 5877
rect 7519 5809 7553 5816
rect 7519 5782 7553 5809
rect 7519 5741 7553 5744
rect 7519 5710 7553 5741
rect 7519 5639 7553 5672
rect 7519 5638 7553 5639
rect 7519 5571 7553 5600
rect 7519 5566 7553 5571
rect 7519 5503 7553 5528
rect 7519 5494 7553 5503
rect 7519 5435 7553 5456
rect 7519 5422 7553 5435
rect 7519 5367 7553 5384
rect 7519 5350 7553 5367
rect 7519 5299 7553 5312
rect 7519 5278 7553 5299
rect 7519 5231 7553 5240
rect 7519 5206 7553 5231
rect 7519 5163 7553 5168
rect 7519 5134 7553 5163
rect 7519 5095 7553 5096
rect 7519 5062 7553 5095
rect 7519 4993 7553 5024
rect 7519 4990 7553 4993
rect 7519 4925 7553 4952
rect 7519 4918 7553 4925
rect 7519 4857 7553 4880
rect 7519 4846 7553 4857
rect 7519 4789 7553 4808
rect 7519 4774 7553 4789
rect 7519 4721 7553 4736
rect 7519 4702 7553 4721
rect 7519 4653 7553 4664
rect 7519 4630 7553 4653
rect 7519 4585 7553 4592
rect 7519 4558 7553 4585
rect 7519 4517 7553 4520
rect 7519 4486 7553 4517
rect 7519 4415 7553 4448
rect 7519 4414 7553 4415
rect 7519 4347 7553 4376
rect 7519 4342 7553 4347
rect 7519 4279 7553 4304
rect 7519 4270 7553 4279
rect 7519 4211 7553 4232
rect 7519 4198 7553 4211
rect 7519 4143 7553 4160
rect 7519 4126 7553 4143
rect 7519 4075 7553 4088
rect 7519 4054 7553 4075
rect 7519 4007 7553 4016
rect 7519 3982 7553 4007
rect 7519 3939 7553 3944
rect 7519 3910 7553 3939
rect 7519 3871 7553 3872
rect 7519 3838 7553 3871
rect 7519 3769 7553 3800
rect 7519 3766 7553 3769
rect 7519 3701 7553 3728
rect 7519 3694 7553 3701
rect 7519 3633 7553 3656
rect 7519 3622 7553 3633
rect 7519 3565 7553 3584
rect 7519 3550 7553 3565
rect 7519 3497 7553 3512
rect 7519 3478 7553 3497
rect 7519 3429 7553 3440
rect 7519 3406 7553 3429
rect 7519 3361 7553 3368
rect 7519 3334 7553 3361
rect 7519 3293 7553 3295
rect 7519 3261 7553 3293
rect 7519 3191 7553 3222
rect 7519 3188 7553 3191
rect 7519 3123 7553 3149
rect 7519 3115 7553 3123
rect 7519 3055 7553 3076
rect 7519 3042 7553 3055
rect 7519 2987 7553 3003
rect 7519 2969 7553 2987
rect 7519 2919 7553 2930
rect 7519 2896 7553 2919
rect 7519 2851 7553 2857
rect 7519 2823 7553 2851
rect 7519 2783 7553 2784
rect 7519 2750 7553 2783
rect 7519 2681 7553 2711
rect 7519 2677 7553 2681
rect 7519 2613 7553 2638
rect 7519 2604 7553 2613
rect 7519 2545 7553 2565
rect 7519 2531 7553 2545
rect 7519 2477 7553 2492
rect 7519 2458 7553 2477
rect 7519 2409 7553 2419
rect 7519 2385 7553 2409
rect 7519 2341 7553 2346
rect 7519 2312 7553 2341
rect 7519 2239 7553 2273
rect 7519 2171 7553 2200
rect 7519 2166 7553 2171
rect 7519 2103 7553 2127
rect 7519 2093 7553 2103
rect 7519 2035 7553 2054
rect 7519 2020 7553 2035
rect 7519 1967 7553 1981
rect 7519 1947 7553 1967
rect 7519 1899 7553 1908
rect 7519 1874 7553 1899
rect 7519 1831 7553 1835
rect 7519 1801 7553 1831
rect 5076 1729 5106 1763
rect 5106 1729 5110 1763
rect 5151 1729 5174 1763
rect 5174 1729 5185 1763
rect 5225 1729 5242 1763
rect 5242 1729 5259 1763
rect 5299 1729 5310 1763
rect 5310 1729 5333 1763
rect 5373 1729 5378 1763
rect 5378 1729 5407 1763
rect 5447 1729 5480 1763
rect 5480 1729 5481 1763
rect 5521 1729 5548 1763
rect 5548 1729 5555 1763
rect 5595 1729 5616 1763
rect 5616 1729 5629 1763
rect 5669 1729 5684 1763
rect 5684 1729 5703 1763
rect 5743 1729 5752 1763
rect 5752 1729 5777 1763
rect 5817 1729 5820 1763
rect 5820 1729 5851 1763
rect 5891 1729 5922 1763
rect 5922 1729 5925 1763
rect 5965 1729 5990 1763
rect 5990 1729 5999 1763
rect 6039 1729 6058 1763
rect 6058 1729 6073 1763
rect 6113 1729 6126 1763
rect 6126 1729 6147 1763
rect 6187 1729 6194 1763
rect 6194 1729 6221 1763
rect 6261 1729 6262 1763
rect 6262 1729 6295 1763
rect 6335 1729 6364 1763
rect 6364 1729 6369 1763
rect 6409 1729 6432 1763
rect 6432 1729 6443 1763
rect 6483 1729 6500 1763
rect 6500 1729 6517 1763
rect 6557 1729 6568 1763
rect 6568 1729 6591 1763
rect 6631 1729 6636 1763
rect 6636 1729 6665 1763
rect 6705 1729 6738 1763
rect 6738 1729 6739 1763
rect 6779 1729 6806 1763
rect 6806 1729 6813 1763
rect 6853 1729 6874 1763
rect 6874 1729 6887 1763
rect 6927 1729 6942 1763
rect 6942 1729 6961 1763
rect 7001 1729 7010 1763
rect 7010 1729 7035 1763
rect 7075 1729 7078 1763
rect 7078 1729 7109 1763
rect 7149 1729 7180 1763
rect 7180 1729 7183 1763
rect 7223 1729 7248 1763
rect 7248 1729 7257 1763
rect 7297 1729 7316 1763
rect 7316 1729 7331 1763
rect 7371 1729 7384 1763
rect 7384 1729 7405 1763
rect 7445 1729 7479 1763
rect 7876 17511 9278 17549
rect 7876 17477 7880 17511
rect 7880 17477 7914 17511
rect 7914 17477 8016 17511
rect 8016 17477 8050 17511
rect 8050 17477 8152 17511
rect 8152 17477 8186 17511
rect 8186 17477 8288 17511
rect 8288 17477 8322 17511
rect 8322 17477 8424 17511
rect 8424 17477 8458 17511
rect 8458 17477 8560 17511
rect 8560 17477 8594 17511
rect 8594 17477 8696 17511
rect 8696 17477 8730 17511
rect 8730 17477 8832 17511
rect 8832 17477 8866 17511
rect 8866 17477 8968 17511
rect 8968 17477 9002 17511
rect 9002 17477 9104 17511
rect 9104 17477 9138 17511
rect 9138 17477 9240 17511
rect 9240 17477 9274 17511
rect 9274 17477 9278 17511
rect 7876 17375 9278 17477
rect 7876 17341 7880 17375
rect 7880 17341 7914 17375
rect 7914 17341 8016 17375
rect 8016 17341 8050 17375
rect 8050 17341 8152 17375
rect 8152 17341 8186 17375
rect 8186 17341 8288 17375
rect 8288 17341 8322 17375
rect 8322 17341 8424 17375
rect 8424 17341 8458 17375
rect 8458 17341 8560 17375
rect 8560 17341 8594 17375
rect 8594 17341 8696 17375
rect 8696 17341 8730 17375
rect 8730 17341 8832 17375
rect 8832 17341 8866 17375
rect 8866 17341 8968 17375
rect 8968 17341 9002 17375
rect 9002 17341 9104 17375
rect 9104 17341 9138 17375
rect 9138 17341 9240 17375
rect 9240 17341 9274 17375
rect 9274 17341 9278 17375
rect 7876 17239 9278 17341
rect 7876 17205 7880 17239
rect 7880 17205 7914 17239
rect 7914 17205 8016 17239
rect 8016 17205 8050 17239
rect 8050 17205 8152 17239
rect 8152 17205 8186 17239
rect 8186 17205 8288 17239
rect 8288 17205 8322 17239
rect 8322 17205 8424 17239
rect 8424 17205 8458 17239
rect 8458 17205 8560 17239
rect 8560 17205 8594 17239
rect 8594 17205 8696 17239
rect 8696 17205 8730 17239
rect 8730 17205 8832 17239
rect 8832 17205 8866 17239
rect 8866 17205 8968 17239
rect 8968 17205 9002 17239
rect 9002 17205 9104 17239
rect 9104 17205 9138 17239
rect 9138 17205 9240 17239
rect 9240 17205 9274 17239
rect 9274 17205 9278 17239
rect 7876 17103 9278 17205
rect 7876 17069 7880 17103
rect 7880 17069 7914 17103
rect 7914 17069 8016 17103
rect 8016 17069 8050 17103
rect 8050 17069 8152 17103
rect 8152 17069 8186 17103
rect 8186 17069 8288 17103
rect 8288 17069 8322 17103
rect 8322 17069 8424 17103
rect 8424 17069 8458 17103
rect 8458 17069 8560 17103
rect 8560 17069 8594 17103
rect 8594 17069 8696 17103
rect 8696 17069 8730 17103
rect 8730 17069 8832 17103
rect 8832 17069 8866 17103
rect 8866 17069 8968 17103
rect 8968 17069 9002 17103
rect 9002 17069 9104 17103
rect 9104 17069 9138 17103
rect 9138 17069 9240 17103
rect 9240 17069 9274 17103
rect 9274 17069 9278 17103
rect 7876 16967 9278 17069
rect 7876 16933 7880 16967
rect 7880 16933 7914 16967
rect 7914 16933 8016 16967
rect 8016 16933 8050 16967
rect 8050 16933 8152 16967
rect 8152 16933 8186 16967
rect 8186 16933 8288 16967
rect 8288 16933 8322 16967
rect 8322 16933 8424 16967
rect 8424 16933 8458 16967
rect 8458 16933 8560 16967
rect 8560 16933 8594 16967
rect 8594 16933 8696 16967
rect 8696 16933 8730 16967
rect 8730 16933 8832 16967
rect 8832 16933 8866 16967
rect 8866 16933 8968 16967
rect 8968 16933 9002 16967
rect 9002 16933 9104 16967
rect 9104 16933 9138 16967
rect 9138 16933 9240 16967
rect 9240 16933 9274 16967
rect 9274 16933 9278 16967
rect 7876 16831 9278 16933
rect 7876 16797 7880 16831
rect 7880 16797 7914 16831
rect 7914 16797 8016 16831
rect 8016 16797 8050 16831
rect 8050 16797 8152 16831
rect 8152 16797 8186 16831
rect 8186 16797 8288 16831
rect 8288 16797 8322 16831
rect 8322 16797 8424 16831
rect 8424 16797 8458 16831
rect 8458 16797 8560 16831
rect 8560 16797 8594 16831
rect 8594 16797 8696 16831
rect 8696 16797 8730 16831
rect 8730 16797 8832 16831
rect 8832 16797 8866 16831
rect 8866 16797 8968 16831
rect 8968 16797 9002 16831
rect 9002 16797 9104 16831
rect 9104 16797 9138 16831
rect 9138 16797 9240 16831
rect 9240 16797 9274 16831
rect 9274 16797 9278 16831
rect 7876 16695 9278 16797
rect 7876 16661 7880 16695
rect 7880 16661 7914 16695
rect 7914 16661 8016 16695
rect 8016 16661 8050 16695
rect 8050 16661 8152 16695
rect 8152 16661 8186 16695
rect 8186 16661 8288 16695
rect 8288 16661 8322 16695
rect 8322 16661 8424 16695
rect 8424 16661 8458 16695
rect 8458 16661 8560 16695
rect 8560 16661 8594 16695
rect 8594 16661 8696 16695
rect 8696 16661 8730 16695
rect 8730 16661 8832 16695
rect 8832 16661 8866 16695
rect 8866 16661 8968 16695
rect 8968 16661 9002 16695
rect 9002 16661 9104 16695
rect 9104 16661 9138 16695
rect 9138 16661 9240 16695
rect 9240 16661 9274 16695
rect 9274 16661 9278 16695
rect 7876 16559 9278 16661
rect 7876 16525 7880 16559
rect 7880 16525 7914 16559
rect 7914 16525 8016 16559
rect 8016 16525 8050 16559
rect 8050 16525 8152 16559
rect 8152 16525 8186 16559
rect 8186 16525 8288 16559
rect 8288 16525 8322 16559
rect 8322 16525 8424 16559
rect 8424 16525 8458 16559
rect 8458 16525 8560 16559
rect 8560 16525 8594 16559
rect 8594 16525 8696 16559
rect 8696 16525 8730 16559
rect 8730 16525 8832 16559
rect 8832 16525 8866 16559
rect 8866 16525 8968 16559
rect 8968 16525 9002 16559
rect 9002 16525 9104 16559
rect 9104 16525 9138 16559
rect 9138 16525 9240 16559
rect 9240 16525 9274 16559
rect 9274 16525 9278 16559
rect 7876 16423 9278 16525
rect 7876 16389 7880 16423
rect 7880 16389 7914 16423
rect 7914 16389 8016 16423
rect 8016 16389 8050 16423
rect 8050 16389 8152 16423
rect 8152 16389 8186 16423
rect 8186 16389 8288 16423
rect 8288 16389 8322 16423
rect 8322 16389 8424 16423
rect 8424 16389 8458 16423
rect 8458 16389 8560 16423
rect 8560 16389 8594 16423
rect 8594 16389 8696 16423
rect 8696 16389 8730 16423
rect 8730 16389 8832 16423
rect 8832 16389 8866 16423
rect 8866 16389 8968 16423
rect 8968 16389 9002 16423
rect 9002 16389 9104 16423
rect 9104 16389 9138 16423
rect 9138 16389 9240 16423
rect 9240 16389 9274 16423
rect 9274 16389 9278 16423
rect 7876 16287 9278 16389
rect 7876 16253 7880 16287
rect 7880 16253 7914 16287
rect 7914 16253 8016 16287
rect 8016 16253 8050 16287
rect 8050 16253 8152 16287
rect 8152 16253 8186 16287
rect 8186 16253 8288 16287
rect 8288 16253 8322 16287
rect 8322 16253 8424 16287
rect 8424 16253 8458 16287
rect 8458 16253 8560 16287
rect 8560 16253 8594 16287
rect 8594 16253 8696 16287
rect 8696 16253 8730 16287
rect 8730 16253 8832 16287
rect 8832 16253 8866 16287
rect 8866 16253 8968 16287
rect 8968 16253 9002 16287
rect 9002 16253 9104 16287
rect 9104 16253 9138 16287
rect 9138 16253 9240 16287
rect 9240 16253 9274 16287
rect 9274 16253 9278 16287
rect 7876 16151 9278 16253
rect 7876 16117 7880 16151
rect 7880 16117 7914 16151
rect 7914 16117 8016 16151
rect 8016 16117 8050 16151
rect 8050 16117 8152 16151
rect 8152 16117 8186 16151
rect 8186 16117 8288 16151
rect 8288 16117 8322 16151
rect 8322 16117 8424 16151
rect 8424 16117 8458 16151
rect 8458 16117 8560 16151
rect 8560 16117 8594 16151
rect 8594 16117 8696 16151
rect 8696 16117 8730 16151
rect 8730 16117 8832 16151
rect 8832 16117 8866 16151
rect 8866 16117 8968 16151
rect 8968 16117 9002 16151
rect 9002 16117 9104 16151
rect 9104 16117 9138 16151
rect 9138 16117 9240 16151
rect 9240 16117 9274 16151
rect 9274 16117 9278 16151
rect 7876 16015 9278 16117
rect 7876 15981 7880 16015
rect 7880 15981 7914 16015
rect 7914 15981 8016 16015
rect 8016 15981 8050 16015
rect 8050 15981 8152 16015
rect 8152 15981 8186 16015
rect 8186 15981 8288 16015
rect 8288 15981 8322 16015
rect 8322 15981 8424 16015
rect 8424 15981 8458 16015
rect 8458 15981 8560 16015
rect 8560 15981 8594 16015
rect 8594 15981 8696 16015
rect 8696 15981 8730 16015
rect 8730 15981 8832 16015
rect 8832 15981 8866 16015
rect 8866 15981 8968 16015
rect 8968 15981 9002 16015
rect 9002 15981 9104 16015
rect 9104 15981 9138 16015
rect 9138 15981 9240 16015
rect 9240 15981 9274 16015
rect 9274 15981 9278 16015
rect 7876 15879 9278 15981
rect 7876 15845 7880 15879
rect 7880 15845 7914 15879
rect 7914 15845 8016 15879
rect 8016 15845 8050 15879
rect 8050 15845 8152 15879
rect 8152 15845 8186 15879
rect 8186 15845 8288 15879
rect 8288 15845 8322 15879
rect 8322 15845 8424 15879
rect 8424 15845 8458 15879
rect 8458 15845 8560 15879
rect 8560 15845 8594 15879
rect 8594 15845 8696 15879
rect 8696 15845 8730 15879
rect 8730 15845 8832 15879
rect 8832 15845 8866 15879
rect 8866 15845 8968 15879
rect 8968 15845 9002 15879
rect 9002 15845 9104 15879
rect 9104 15845 9138 15879
rect 9138 15845 9240 15879
rect 9240 15845 9274 15879
rect 9274 15845 9278 15879
rect 7876 15743 9278 15845
rect 7876 15709 7880 15743
rect 7880 15709 7914 15743
rect 7914 15709 8016 15743
rect 8016 15709 8050 15743
rect 8050 15709 8152 15743
rect 8152 15709 8186 15743
rect 8186 15709 8288 15743
rect 8288 15709 8322 15743
rect 8322 15709 8424 15743
rect 8424 15709 8458 15743
rect 8458 15709 8560 15743
rect 8560 15709 8594 15743
rect 8594 15709 8696 15743
rect 8696 15709 8730 15743
rect 8730 15709 8832 15743
rect 8832 15709 8866 15743
rect 8866 15709 8968 15743
rect 8968 15709 9002 15743
rect 9002 15709 9104 15743
rect 9104 15709 9138 15743
rect 9138 15709 9240 15743
rect 9240 15709 9274 15743
rect 9274 15709 9278 15743
rect 7876 15607 9278 15709
rect 7876 15573 7880 15607
rect 7880 15573 7914 15607
rect 7914 15573 8016 15607
rect 8016 15573 8050 15607
rect 8050 15573 8152 15607
rect 8152 15573 8186 15607
rect 8186 15573 8288 15607
rect 8288 15573 8322 15607
rect 8322 15573 8424 15607
rect 8424 15573 8458 15607
rect 8458 15573 8560 15607
rect 8560 15573 8594 15607
rect 8594 15573 8696 15607
rect 8696 15573 8730 15607
rect 8730 15573 8832 15607
rect 8832 15573 8866 15607
rect 8866 15573 8968 15607
rect 8968 15573 9002 15607
rect 9002 15573 9104 15607
rect 9104 15573 9138 15607
rect 9138 15573 9240 15607
rect 9240 15573 9274 15607
rect 9274 15573 9278 15607
rect 7876 15471 9278 15573
rect 7876 15437 7880 15471
rect 7880 15437 7914 15471
rect 7914 15437 8016 15471
rect 8016 15437 8050 15471
rect 8050 15437 8152 15471
rect 8152 15437 8186 15471
rect 8186 15437 8288 15471
rect 8288 15437 8322 15471
rect 8322 15437 8424 15471
rect 8424 15437 8458 15471
rect 8458 15437 8560 15471
rect 8560 15437 8594 15471
rect 8594 15437 8696 15471
rect 8696 15437 8730 15471
rect 8730 15437 8832 15471
rect 8832 15437 8866 15471
rect 8866 15437 8968 15471
rect 8968 15437 9002 15471
rect 9002 15437 9104 15471
rect 9104 15437 9138 15471
rect 9138 15437 9240 15471
rect 9240 15437 9274 15471
rect 9274 15437 9278 15471
rect 7876 15335 9278 15437
rect 7876 15301 7880 15335
rect 7880 15301 7914 15335
rect 7914 15301 8016 15335
rect 8016 15301 8050 15335
rect 8050 15301 8152 15335
rect 8152 15301 8186 15335
rect 8186 15301 8288 15335
rect 8288 15301 8322 15335
rect 8322 15301 8424 15335
rect 8424 15301 8458 15335
rect 8458 15301 8560 15335
rect 8560 15301 8594 15335
rect 8594 15301 8696 15335
rect 8696 15301 8730 15335
rect 8730 15301 8832 15335
rect 8832 15301 8866 15335
rect 8866 15301 8968 15335
rect 8968 15301 9002 15335
rect 9002 15301 9104 15335
rect 9104 15301 9138 15335
rect 9138 15301 9240 15335
rect 9240 15301 9274 15335
rect 9274 15301 9278 15335
rect 7876 15199 9278 15301
rect 7876 15165 7880 15199
rect 7880 15165 7914 15199
rect 7914 15165 8016 15199
rect 8016 15165 8050 15199
rect 8050 15165 8152 15199
rect 8152 15165 8186 15199
rect 8186 15165 8288 15199
rect 8288 15165 8322 15199
rect 8322 15165 8424 15199
rect 8424 15165 8458 15199
rect 8458 15165 8560 15199
rect 8560 15165 8594 15199
rect 8594 15165 8696 15199
rect 8696 15165 8730 15199
rect 8730 15165 8832 15199
rect 8832 15165 8866 15199
rect 8866 15165 8968 15199
rect 8968 15165 9002 15199
rect 9002 15165 9104 15199
rect 9104 15165 9138 15199
rect 9138 15165 9240 15199
rect 9240 15165 9274 15199
rect 9274 15165 9278 15199
rect 7876 15063 9278 15165
rect 7876 15029 7880 15063
rect 7880 15029 7914 15063
rect 7914 15029 8016 15063
rect 8016 15029 8050 15063
rect 8050 15029 8152 15063
rect 8152 15029 8186 15063
rect 8186 15029 8288 15063
rect 8288 15029 8322 15063
rect 8322 15029 8424 15063
rect 8424 15029 8458 15063
rect 8458 15029 8560 15063
rect 8560 15029 8594 15063
rect 8594 15029 8696 15063
rect 8696 15029 8730 15063
rect 8730 15029 8832 15063
rect 8832 15029 8866 15063
rect 8866 15029 8968 15063
rect 8968 15029 9002 15063
rect 9002 15029 9104 15063
rect 9104 15029 9138 15063
rect 9138 15029 9240 15063
rect 9240 15029 9274 15063
rect 9274 15029 9278 15063
rect 7876 14927 9278 15029
rect 7876 14893 7880 14927
rect 7880 14893 7914 14927
rect 7914 14893 8016 14927
rect 8016 14893 8050 14927
rect 8050 14893 8152 14927
rect 8152 14893 8186 14927
rect 8186 14893 8288 14927
rect 8288 14893 8322 14927
rect 8322 14893 8424 14927
rect 8424 14893 8458 14927
rect 8458 14893 8560 14927
rect 8560 14893 8594 14927
rect 8594 14893 8696 14927
rect 8696 14893 8730 14927
rect 8730 14893 8832 14927
rect 8832 14893 8866 14927
rect 8866 14893 8968 14927
rect 8968 14893 9002 14927
rect 9002 14893 9104 14927
rect 9104 14893 9138 14927
rect 9138 14893 9240 14927
rect 9240 14893 9274 14927
rect 9274 14893 9278 14927
rect 7876 14791 9278 14893
rect 7876 14757 7880 14791
rect 7880 14757 7914 14791
rect 7914 14757 8016 14791
rect 8016 14757 8050 14791
rect 8050 14757 8152 14791
rect 8152 14757 8186 14791
rect 8186 14757 8288 14791
rect 8288 14757 8322 14791
rect 8322 14757 8424 14791
rect 8424 14757 8458 14791
rect 8458 14757 8560 14791
rect 8560 14757 8594 14791
rect 8594 14757 8696 14791
rect 8696 14757 8730 14791
rect 8730 14757 8832 14791
rect 8832 14757 8866 14791
rect 8866 14757 8968 14791
rect 8968 14757 9002 14791
rect 9002 14757 9104 14791
rect 9104 14757 9138 14791
rect 9138 14757 9240 14791
rect 9240 14757 9274 14791
rect 9274 14757 9278 14791
rect 7876 14655 9278 14757
rect 7876 14621 7880 14655
rect 7880 14621 7914 14655
rect 7914 14621 8016 14655
rect 8016 14621 8050 14655
rect 8050 14621 8152 14655
rect 8152 14621 8186 14655
rect 8186 14621 8288 14655
rect 8288 14621 8322 14655
rect 8322 14621 8424 14655
rect 8424 14621 8458 14655
rect 8458 14621 8560 14655
rect 8560 14621 8594 14655
rect 8594 14621 8696 14655
rect 8696 14621 8730 14655
rect 8730 14621 8832 14655
rect 8832 14621 8866 14655
rect 8866 14621 8968 14655
rect 8968 14621 9002 14655
rect 9002 14621 9104 14655
rect 9104 14621 9138 14655
rect 9138 14621 9240 14655
rect 9240 14621 9274 14655
rect 9274 14621 9278 14655
rect 7876 14519 9278 14621
rect 7876 14485 7880 14519
rect 7880 14485 7914 14519
rect 7914 14485 8016 14519
rect 8016 14485 8050 14519
rect 8050 14485 8152 14519
rect 8152 14485 8186 14519
rect 8186 14485 8288 14519
rect 8288 14485 8322 14519
rect 8322 14485 8424 14519
rect 8424 14485 8458 14519
rect 8458 14485 8560 14519
rect 8560 14485 8594 14519
rect 8594 14485 8696 14519
rect 8696 14485 8730 14519
rect 8730 14485 8832 14519
rect 8832 14485 8866 14519
rect 8866 14485 8968 14519
rect 8968 14485 9002 14519
rect 9002 14485 9104 14519
rect 9104 14485 9138 14519
rect 9138 14485 9240 14519
rect 9240 14485 9274 14519
rect 9274 14485 9278 14519
rect 7876 14383 9278 14485
rect 7876 14349 7880 14383
rect 7880 14349 7914 14383
rect 7914 14349 8016 14383
rect 8016 14349 8050 14383
rect 8050 14349 8152 14383
rect 8152 14349 8186 14383
rect 8186 14349 8288 14383
rect 8288 14349 8322 14383
rect 8322 14349 8424 14383
rect 8424 14349 8458 14383
rect 8458 14349 8560 14383
rect 8560 14349 8594 14383
rect 8594 14349 8696 14383
rect 8696 14349 8730 14383
rect 8730 14349 8832 14383
rect 8832 14349 8866 14383
rect 8866 14349 8968 14383
rect 8968 14349 9002 14383
rect 9002 14349 9104 14383
rect 9104 14349 9138 14383
rect 9138 14349 9240 14383
rect 9240 14349 9274 14383
rect 9274 14349 9278 14383
rect 7876 14247 9278 14349
rect 7876 14213 7880 14247
rect 7880 14213 7914 14247
rect 7914 14213 8016 14247
rect 8016 14213 8050 14247
rect 8050 14213 8152 14247
rect 8152 14213 8186 14247
rect 8186 14213 8288 14247
rect 8288 14213 8322 14247
rect 8322 14213 8424 14247
rect 8424 14213 8458 14247
rect 8458 14213 8560 14247
rect 8560 14213 8594 14247
rect 8594 14213 8696 14247
rect 8696 14213 8730 14247
rect 8730 14213 8832 14247
rect 8832 14213 8866 14247
rect 8866 14213 8968 14247
rect 8968 14213 9002 14247
rect 9002 14213 9104 14247
rect 9104 14213 9138 14247
rect 9138 14213 9240 14247
rect 9240 14213 9274 14247
rect 9274 14213 9278 14247
rect 7876 14111 9278 14213
rect 7876 14077 7880 14111
rect 7880 14077 7914 14111
rect 7914 14077 8016 14111
rect 8016 14077 8050 14111
rect 8050 14077 8152 14111
rect 8152 14077 8186 14111
rect 8186 14077 8288 14111
rect 8288 14077 8322 14111
rect 8322 14077 8424 14111
rect 8424 14077 8458 14111
rect 8458 14077 8560 14111
rect 8560 14077 8594 14111
rect 8594 14077 8696 14111
rect 8696 14077 8730 14111
rect 8730 14077 8832 14111
rect 8832 14077 8866 14111
rect 8866 14077 8968 14111
rect 8968 14077 9002 14111
rect 9002 14077 9104 14111
rect 9104 14077 9138 14111
rect 9138 14077 9240 14111
rect 9240 14077 9274 14111
rect 9274 14077 9278 14111
rect 7876 13975 9278 14077
rect 7876 13941 7880 13975
rect 7880 13941 7914 13975
rect 7914 13941 8016 13975
rect 8016 13941 8050 13975
rect 8050 13941 8152 13975
rect 8152 13941 8186 13975
rect 8186 13941 8288 13975
rect 8288 13941 8322 13975
rect 8322 13941 8424 13975
rect 8424 13941 8458 13975
rect 8458 13941 8560 13975
rect 8560 13941 8594 13975
rect 8594 13941 8696 13975
rect 8696 13941 8730 13975
rect 8730 13941 8832 13975
rect 8832 13941 8866 13975
rect 8866 13941 8968 13975
rect 8968 13941 9002 13975
rect 9002 13941 9104 13975
rect 9104 13941 9138 13975
rect 9138 13941 9240 13975
rect 9240 13941 9274 13975
rect 9274 13941 9278 13975
rect 7876 13839 9278 13941
rect 7876 13805 7880 13839
rect 7880 13805 7914 13839
rect 7914 13805 8016 13839
rect 8016 13805 8050 13839
rect 8050 13805 8152 13839
rect 8152 13805 8186 13839
rect 8186 13805 8288 13839
rect 8288 13805 8322 13839
rect 8322 13805 8424 13839
rect 8424 13805 8458 13839
rect 8458 13805 8560 13839
rect 8560 13805 8594 13839
rect 8594 13805 8696 13839
rect 8696 13805 8730 13839
rect 8730 13805 8832 13839
rect 8832 13805 8866 13839
rect 8866 13805 8968 13839
rect 8968 13805 9002 13839
rect 9002 13805 9104 13839
rect 9104 13805 9138 13839
rect 9138 13805 9240 13839
rect 9240 13805 9274 13839
rect 9274 13805 9278 13839
rect 7876 13703 9278 13805
rect 7876 13669 7880 13703
rect 7880 13669 7914 13703
rect 7914 13669 8016 13703
rect 8016 13669 8050 13703
rect 8050 13669 8152 13703
rect 8152 13669 8186 13703
rect 8186 13669 8288 13703
rect 8288 13669 8322 13703
rect 8322 13669 8424 13703
rect 8424 13669 8458 13703
rect 8458 13669 8560 13703
rect 8560 13669 8594 13703
rect 8594 13669 8696 13703
rect 8696 13669 8730 13703
rect 8730 13669 8832 13703
rect 8832 13669 8866 13703
rect 8866 13669 8968 13703
rect 8968 13669 9002 13703
rect 9002 13669 9104 13703
rect 9104 13669 9138 13703
rect 9138 13669 9240 13703
rect 9240 13669 9274 13703
rect 9274 13669 9278 13703
rect 7876 13567 9278 13669
rect 7876 13533 7880 13567
rect 7880 13533 7914 13567
rect 7914 13533 8016 13567
rect 8016 13533 8050 13567
rect 8050 13533 8152 13567
rect 8152 13533 8186 13567
rect 8186 13533 8288 13567
rect 8288 13533 8322 13567
rect 8322 13533 8424 13567
rect 8424 13533 8458 13567
rect 8458 13533 8560 13567
rect 8560 13533 8594 13567
rect 8594 13533 8696 13567
rect 8696 13533 8730 13567
rect 8730 13533 8832 13567
rect 8832 13533 8866 13567
rect 8866 13533 8968 13567
rect 8968 13533 9002 13567
rect 9002 13533 9104 13567
rect 9104 13533 9138 13567
rect 9138 13533 9240 13567
rect 9240 13533 9274 13567
rect 9274 13533 9278 13567
rect 7876 13431 9278 13533
rect 7876 13397 7880 13431
rect 7880 13397 7914 13431
rect 7914 13397 8016 13431
rect 8016 13397 8050 13431
rect 8050 13397 8152 13431
rect 8152 13397 8186 13431
rect 8186 13397 8288 13431
rect 8288 13397 8322 13431
rect 8322 13397 8424 13431
rect 8424 13397 8458 13431
rect 8458 13397 8560 13431
rect 8560 13397 8594 13431
rect 8594 13397 8696 13431
rect 8696 13397 8730 13431
rect 8730 13397 8832 13431
rect 8832 13397 8866 13431
rect 8866 13397 8968 13431
rect 8968 13397 9002 13431
rect 9002 13397 9104 13431
rect 9104 13397 9138 13431
rect 9138 13397 9240 13431
rect 9240 13397 9274 13431
rect 9274 13397 9278 13431
rect 7876 13295 9278 13397
rect 7876 13261 7880 13295
rect 7880 13261 7914 13295
rect 7914 13261 8016 13295
rect 8016 13261 8050 13295
rect 8050 13261 8152 13295
rect 8152 13261 8186 13295
rect 8186 13261 8288 13295
rect 8288 13261 8322 13295
rect 8322 13261 8424 13295
rect 8424 13261 8458 13295
rect 8458 13261 8560 13295
rect 8560 13261 8594 13295
rect 8594 13261 8696 13295
rect 8696 13261 8730 13295
rect 8730 13261 8832 13295
rect 8832 13261 8866 13295
rect 8866 13261 8968 13295
rect 8968 13261 9002 13295
rect 9002 13261 9104 13295
rect 9104 13261 9138 13295
rect 9138 13261 9240 13295
rect 9240 13261 9274 13295
rect 9274 13261 9278 13295
rect 7876 13159 9278 13261
rect 7876 13125 7880 13159
rect 7880 13125 7914 13159
rect 7914 13125 8016 13159
rect 8016 13125 8050 13159
rect 8050 13125 8152 13159
rect 8152 13125 8186 13159
rect 8186 13125 8288 13159
rect 8288 13125 8322 13159
rect 8322 13125 8424 13159
rect 8424 13125 8458 13159
rect 8458 13125 8560 13159
rect 8560 13125 8594 13159
rect 8594 13125 8696 13159
rect 8696 13125 8730 13159
rect 8730 13125 8832 13159
rect 8832 13125 8866 13159
rect 8866 13125 8968 13159
rect 8968 13125 9002 13159
rect 9002 13125 9104 13159
rect 9104 13125 9138 13159
rect 9138 13125 9240 13159
rect 9240 13125 9274 13159
rect 9274 13125 9278 13159
rect 7876 13023 9278 13125
rect 7876 12989 7880 13023
rect 7880 12989 7914 13023
rect 7914 12989 8016 13023
rect 8016 12989 8050 13023
rect 8050 12989 8152 13023
rect 8152 12989 8186 13023
rect 8186 12989 8288 13023
rect 8288 12989 8322 13023
rect 8322 12989 8424 13023
rect 8424 12989 8458 13023
rect 8458 12989 8560 13023
rect 8560 12989 8594 13023
rect 8594 12989 8696 13023
rect 8696 12989 8730 13023
rect 8730 12989 8832 13023
rect 8832 12989 8866 13023
rect 8866 12989 8968 13023
rect 8968 12989 9002 13023
rect 9002 12989 9104 13023
rect 9104 12989 9138 13023
rect 9138 12989 9240 13023
rect 9240 12989 9274 13023
rect 9274 12989 9278 13023
rect 7876 12887 9278 12989
rect 7876 12853 7880 12887
rect 7880 12853 7914 12887
rect 7914 12853 8016 12887
rect 8016 12853 8050 12887
rect 8050 12853 8152 12887
rect 8152 12853 8186 12887
rect 8186 12853 8288 12887
rect 8288 12853 8322 12887
rect 8322 12853 8424 12887
rect 8424 12853 8458 12887
rect 8458 12853 8560 12887
rect 8560 12853 8594 12887
rect 8594 12853 8696 12887
rect 8696 12853 8730 12887
rect 8730 12853 8832 12887
rect 8832 12853 8866 12887
rect 8866 12853 8968 12887
rect 8968 12853 9002 12887
rect 9002 12853 9104 12887
rect 9104 12853 9138 12887
rect 9138 12853 9240 12887
rect 9240 12853 9274 12887
rect 9274 12853 9278 12887
rect 7876 12751 9278 12853
rect 7876 12717 7880 12751
rect 7880 12717 7914 12751
rect 7914 12717 8016 12751
rect 8016 12717 8050 12751
rect 8050 12717 8152 12751
rect 8152 12717 8186 12751
rect 8186 12717 8288 12751
rect 8288 12717 8322 12751
rect 8322 12717 8424 12751
rect 8424 12717 8458 12751
rect 8458 12717 8560 12751
rect 8560 12717 8594 12751
rect 8594 12717 8696 12751
rect 8696 12717 8730 12751
rect 8730 12717 8832 12751
rect 8832 12717 8866 12751
rect 8866 12717 8968 12751
rect 8968 12717 9002 12751
rect 9002 12717 9104 12751
rect 9104 12717 9138 12751
rect 9138 12717 9240 12751
rect 9240 12717 9274 12751
rect 9274 12717 9278 12751
rect 7876 12615 9278 12717
rect 7876 12581 7880 12615
rect 7880 12581 7914 12615
rect 7914 12581 8016 12615
rect 8016 12581 8050 12615
rect 8050 12581 8152 12615
rect 8152 12581 8186 12615
rect 8186 12581 8288 12615
rect 8288 12581 8322 12615
rect 8322 12581 8424 12615
rect 8424 12581 8458 12615
rect 8458 12581 8560 12615
rect 8560 12581 8594 12615
rect 8594 12581 8696 12615
rect 8696 12581 8730 12615
rect 8730 12581 8832 12615
rect 8832 12581 8866 12615
rect 8866 12581 8968 12615
rect 8968 12581 9002 12615
rect 9002 12581 9104 12615
rect 9104 12581 9138 12615
rect 9138 12581 9240 12615
rect 9240 12581 9274 12615
rect 9274 12581 9278 12615
rect 7876 12479 9278 12581
rect 7876 12445 7880 12479
rect 7880 12445 7914 12479
rect 7914 12445 8016 12479
rect 8016 12445 8050 12479
rect 8050 12445 8152 12479
rect 8152 12445 8186 12479
rect 8186 12445 8288 12479
rect 8288 12445 8322 12479
rect 8322 12445 8424 12479
rect 8424 12445 8458 12479
rect 8458 12445 8560 12479
rect 8560 12445 8594 12479
rect 8594 12445 8696 12479
rect 8696 12445 8730 12479
rect 8730 12445 8832 12479
rect 8832 12445 8866 12479
rect 8866 12445 8968 12479
rect 8968 12445 9002 12479
rect 9002 12445 9104 12479
rect 9104 12445 9138 12479
rect 9138 12445 9240 12479
rect 9240 12445 9274 12479
rect 9274 12445 9278 12479
rect 7876 12343 9278 12445
rect 7876 12309 7880 12343
rect 7880 12309 7914 12343
rect 7914 12309 8016 12343
rect 8016 12309 8050 12343
rect 8050 12309 8152 12343
rect 8152 12309 8186 12343
rect 8186 12309 8288 12343
rect 8288 12309 8322 12343
rect 8322 12309 8424 12343
rect 8424 12309 8458 12343
rect 8458 12309 8560 12343
rect 8560 12309 8594 12343
rect 8594 12309 8696 12343
rect 8696 12309 8730 12343
rect 8730 12309 8832 12343
rect 8832 12309 8866 12343
rect 8866 12309 8968 12343
rect 8968 12309 9002 12343
rect 9002 12309 9104 12343
rect 9104 12309 9138 12343
rect 9138 12309 9240 12343
rect 9240 12309 9274 12343
rect 9274 12309 9278 12343
rect 7876 12207 9278 12309
rect 7876 12173 7880 12207
rect 7880 12173 7914 12207
rect 7914 12173 8016 12207
rect 8016 12173 8050 12207
rect 8050 12173 8152 12207
rect 8152 12173 8186 12207
rect 8186 12173 8288 12207
rect 8288 12173 8322 12207
rect 8322 12173 8424 12207
rect 8424 12173 8458 12207
rect 8458 12173 8560 12207
rect 8560 12173 8594 12207
rect 8594 12173 8696 12207
rect 8696 12173 8730 12207
rect 8730 12173 8832 12207
rect 8832 12173 8866 12207
rect 8866 12173 8968 12207
rect 8968 12173 9002 12207
rect 9002 12173 9104 12207
rect 9104 12173 9138 12207
rect 9138 12173 9240 12207
rect 9240 12173 9274 12207
rect 9274 12173 9278 12207
rect 7876 12071 9278 12173
rect 7876 12037 7880 12071
rect 7880 12037 7914 12071
rect 7914 12037 8016 12071
rect 8016 12037 8050 12071
rect 8050 12037 8152 12071
rect 8152 12037 8186 12071
rect 8186 12037 8288 12071
rect 8288 12037 8322 12071
rect 8322 12037 8424 12071
rect 8424 12037 8458 12071
rect 8458 12037 8560 12071
rect 8560 12037 8594 12071
rect 8594 12037 8696 12071
rect 8696 12037 8730 12071
rect 8730 12037 8832 12071
rect 8832 12037 8866 12071
rect 8866 12037 8968 12071
rect 8968 12037 9002 12071
rect 9002 12037 9104 12071
rect 9104 12037 9138 12071
rect 9138 12037 9240 12071
rect 9240 12037 9274 12071
rect 9274 12037 9278 12071
rect 7876 11935 9278 12037
rect 7876 11901 7880 11935
rect 7880 11901 7914 11935
rect 7914 11901 8016 11935
rect 8016 11901 8050 11935
rect 8050 11901 8152 11935
rect 8152 11901 8186 11935
rect 8186 11901 8288 11935
rect 8288 11901 8322 11935
rect 8322 11901 8424 11935
rect 8424 11901 8458 11935
rect 8458 11901 8560 11935
rect 8560 11901 8594 11935
rect 8594 11901 8696 11935
rect 8696 11901 8730 11935
rect 8730 11901 8832 11935
rect 8832 11901 8866 11935
rect 8866 11901 8968 11935
rect 8968 11901 9002 11935
rect 9002 11901 9104 11935
rect 9104 11901 9138 11935
rect 9138 11901 9240 11935
rect 9240 11901 9274 11935
rect 9274 11901 9278 11935
rect 7876 11799 9278 11901
rect 7876 11765 7880 11799
rect 7880 11765 7914 11799
rect 7914 11765 8016 11799
rect 8016 11765 8050 11799
rect 8050 11765 8152 11799
rect 8152 11765 8186 11799
rect 8186 11765 8288 11799
rect 8288 11765 8322 11799
rect 8322 11765 8424 11799
rect 8424 11765 8458 11799
rect 8458 11765 8560 11799
rect 8560 11765 8594 11799
rect 8594 11765 8696 11799
rect 8696 11765 8730 11799
rect 8730 11765 8832 11799
rect 8832 11765 8866 11799
rect 8866 11765 8968 11799
rect 8968 11765 9002 11799
rect 9002 11765 9104 11799
rect 9104 11765 9138 11799
rect 9138 11765 9240 11799
rect 9240 11765 9274 11799
rect 9274 11765 9278 11799
rect 7876 11663 9278 11765
rect 7876 11629 7880 11663
rect 7880 11629 7914 11663
rect 7914 11629 8016 11663
rect 8016 11629 8050 11663
rect 8050 11629 8152 11663
rect 8152 11629 8186 11663
rect 8186 11629 8288 11663
rect 8288 11629 8322 11663
rect 8322 11629 8424 11663
rect 8424 11629 8458 11663
rect 8458 11629 8560 11663
rect 8560 11629 8594 11663
rect 8594 11629 8696 11663
rect 8696 11629 8730 11663
rect 8730 11629 8832 11663
rect 8832 11629 8866 11663
rect 8866 11629 8968 11663
rect 8968 11629 9002 11663
rect 9002 11629 9104 11663
rect 9104 11629 9138 11663
rect 9138 11629 9240 11663
rect 9240 11629 9274 11663
rect 9274 11629 9278 11663
rect 7876 11527 9278 11629
rect 7876 11493 7880 11527
rect 7880 11493 7914 11527
rect 7914 11493 8016 11527
rect 8016 11493 8050 11527
rect 8050 11493 8152 11527
rect 8152 11493 8186 11527
rect 8186 11493 8288 11527
rect 8288 11493 8322 11527
rect 8322 11493 8424 11527
rect 8424 11493 8458 11527
rect 8458 11493 8560 11527
rect 8560 11493 8594 11527
rect 8594 11493 8696 11527
rect 8696 11493 8730 11527
rect 8730 11493 8832 11527
rect 8832 11493 8866 11527
rect 8866 11493 8968 11527
rect 8968 11493 9002 11527
rect 9002 11493 9104 11527
rect 9104 11493 9138 11527
rect 9138 11493 9240 11527
rect 9240 11493 9274 11527
rect 9274 11493 9278 11527
rect 7876 11391 9278 11493
rect 7876 11357 7880 11391
rect 7880 11357 7914 11391
rect 7914 11357 8016 11391
rect 8016 11357 8050 11391
rect 8050 11357 8152 11391
rect 8152 11357 8186 11391
rect 8186 11357 8288 11391
rect 8288 11357 8322 11391
rect 8322 11357 8424 11391
rect 8424 11357 8458 11391
rect 8458 11357 8560 11391
rect 8560 11357 8594 11391
rect 8594 11357 8696 11391
rect 8696 11357 8730 11391
rect 8730 11357 8832 11391
rect 8832 11357 8866 11391
rect 8866 11357 8968 11391
rect 8968 11357 9002 11391
rect 9002 11357 9104 11391
rect 9104 11357 9138 11391
rect 9138 11357 9240 11391
rect 9240 11357 9274 11391
rect 9274 11357 9278 11391
rect 7876 11255 9278 11357
rect 7876 11221 7880 11255
rect 7880 11221 7914 11255
rect 7914 11221 8016 11255
rect 8016 11221 8050 11255
rect 8050 11221 8152 11255
rect 8152 11221 8186 11255
rect 8186 11221 8288 11255
rect 8288 11221 8322 11255
rect 8322 11221 8424 11255
rect 8424 11221 8458 11255
rect 8458 11221 8560 11255
rect 8560 11221 8594 11255
rect 8594 11221 8696 11255
rect 8696 11221 8730 11255
rect 8730 11221 8832 11255
rect 8832 11221 8866 11255
rect 8866 11221 8968 11255
rect 8968 11221 9002 11255
rect 9002 11221 9104 11255
rect 9104 11221 9138 11255
rect 9138 11221 9240 11255
rect 9240 11221 9274 11255
rect 9274 11221 9278 11255
rect 7876 11119 9278 11221
rect 7876 11085 7880 11119
rect 7880 11085 7914 11119
rect 7914 11085 8016 11119
rect 8016 11085 8050 11119
rect 8050 11085 8152 11119
rect 8152 11085 8186 11119
rect 8186 11085 8288 11119
rect 8288 11085 8322 11119
rect 8322 11085 8424 11119
rect 8424 11085 8458 11119
rect 8458 11085 8560 11119
rect 8560 11085 8594 11119
rect 8594 11085 8696 11119
rect 8696 11085 8730 11119
rect 8730 11085 8832 11119
rect 8832 11085 8866 11119
rect 8866 11085 8968 11119
rect 8968 11085 9002 11119
rect 9002 11085 9104 11119
rect 9104 11085 9138 11119
rect 9138 11085 9240 11119
rect 9240 11085 9274 11119
rect 9274 11085 9278 11119
rect 7876 10983 9278 11085
rect 7876 10949 7880 10983
rect 7880 10949 7914 10983
rect 7914 10949 8016 10983
rect 8016 10949 8050 10983
rect 8050 10949 8152 10983
rect 8152 10949 8186 10983
rect 8186 10949 8288 10983
rect 8288 10949 8322 10983
rect 8322 10949 8424 10983
rect 8424 10949 8458 10983
rect 8458 10949 8560 10983
rect 8560 10949 8594 10983
rect 8594 10949 8696 10983
rect 8696 10949 8730 10983
rect 8730 10949 8832 10983
rect 8832 10949 8866 10983
rect 8866 10949 8968 10983
rect 8968 10949 9002 10983
rect 9002 10949 9104 10983
rect 9104 10949 9138 10983
rect 9138 10949 9240 10983
rect 9240 10949 9274 10983
rect 9274 10949 9278 10983
rect 7876 10847 9278 10949
rect 7876 10813 7880 10847
rect 7880 10813 7914 10847
rect 7914 10813 8016 10847
rect 8016 10813 8050 10847
rect 8050 10813 8152 10847
rect 8152 10813 8186 10847
rect 8186 10813 8288 10847
rect 8288 10813 8322 10847
rect 8322 10813 8424 10847
rect 8424 10813 8458 10847
rect 8458 10813 8560 10847
rect 8560 10813 8594 10847
rect 8594 10813 8696 10847
rect 8696 10813 8730 10847
rect 8730 10813 8832 10847
rect 8832 10813 8866 10847
rect 8866 10813 8968 10847
rect 8968 10813 9002 10847
rect 9002 10813 9104 10847
rect 9104 10813 9138 10847
rect 9138 10813 9240 10847
rect 9240 10813 9274 10847
rect 9274 10813 9278 10847
rect 7876 10711 9278 10813
rect 7876 10677 7880 10711
rect 7880 10677 7914 10711
rect 7914 10677 8016 10711
rect 8016 10677 8050 10711
rect 8050 10677 8152 10711
rect 8152 10677 8186 10711
rect 8186 10677 8288 10711
rect 8288 10677 8322 10711
rect 8322 10677 8424 10711
rect 8424 10677 8458 10711
rect 8458 10677 8560 10711
rect 8560 10677 8594 10711
rect 8594 10677 8696 10711
rect 8696 10677 8730 10711
rect 8730 10677 8832 10711
rect 8832 10677 8866 10711
rect 8866 10677 8968 10711
rect 8968 10677 9002 10711
rect 9002 10677 9104 10711
rect 9104 10677 9138 10711
rect 9138 10677 9240 10711
rect 9240 10677 9274 10711
rect 9274 10677 9278 10711
rect 7876 10575 9278 10677
rect 7876 10541 7880 10575
rect 7880 10541 7914 10575
rect 7914 10541 8016 10575
rect 8016 10541 8050 10575
rect 8050 10541 8152 10575
rect 8152 10541 8186 10575
rect 8186 10541 8288 10575
rect 8288 10541 8322 10575
rect 8322 10541 8424 10575
rect 8424 10541 8458 10575
rect 8458 10541 8560 10575
rect 8560 10541 8594 10575
rect 8594 10541 8696 10575
rect 8696 10541 8730 10575
rect 8730 10541 8832 10575
rect 8832 10541 8866 10575
rect 8866 10541 8968 10575
rect 8968 10541 9002 10575
rect 9002 10541 9104 10575
rect 9104 10541 9138 10575
rect 9138 10541 9240 10575
rect 9240 10541 9274 10575
rect 9274 10541 9278 10575
rect 7876 10439 9278 10541
rect 7876 10405 7880 10439
rect 7880 10405 7914 10439
rect 7914 10405 8016 10439
rect 8016 10405 8050 10439
rect 8050 10405 8152 10439
rect 8152 10405 8186 10439
rect 8186 10405 8288 10439
rect 8288 10405 8322 10439
rect 8322 10405 8424 10439
rect 8424 10405 8458 10439
rect 8458 10405 8560 10439
rect 8560 10405 8594 10439
rect 8594 10405 8696 10439
rect 8696 10405 8730 10439
rect 8730 10405 8832 10439
rect 8832 10405 8866 10439
rect 8866 10405 8968 10439
rect 8968 10405 9002 10439
rect 9002 10405 9104 10439
rect 9104 10405 9138 10439
rect 9138 10405 9240 10439
rect 9240 10405 9274 10439
rect 9274 10405 9278 10439
rect 7876 10303 9278 10405
rect 7876 10269 7880 10303
rect 7880 10269 7914 10303
rect 7914 10269 8016 10303
rect 8016 10269 8050 10303
rect 8050 10269 8152 10303
rect 8152 10269 8186 10303
rect 8186 10269 8288 10303
rect 8288 10269 8322 10303
rect 8322 10269 8424 10303
rect 8424 10269 8458 10303
rect 8458 10269 8560 10303
rect 8560 10269 8594 10303
rect 8594 10269 8696 10303
rect 8696 10269 8730 10303
rect 8730 10269 8832 10303
rect 8832 10269 8866 10303
rect 8866 10269 8968 10303
rect 8968 10269 9002 10303
rect 9002 10269 9104 10303
rect 9104 10269 9138 10303
rect 9138 10269 9240 10303
rect 9240 10269 9274 10303
rect 9274 10269 9278 10303
rect 7876 10167 9278 10269
rect 7876 10133 7880 10167
rect 7880 10133 7914 10167
rect 7914 10133 8016 10167
rect 8016 10133 8050 10167
rect 8050 10133 8152 10167
rect 8152 10133 8186 10167
rect 8186 10133 8288 10167
rect 8288 10133 8322 10167
rect 8322 10133 8424 10167
rect 8424 10133 8458 10167
rect 8458 10133 8560 10167
rect 8560 10133 8594 10167
rect 8594 10133 8696 10167
rect 8696 10133 8730 10167
rect 8730 10133 8832 10167
rect 8832 10133 8866 10167
rect 8866 10133 8968 10167
rect 8968 10133 9002 10167
rect 9002 10133 9104 10167
rect 9104 10133 9138 10167
rect 9138 10133 9240 10167
rect 9240 10133 9274 10167
rect 9274 10133 9278 10167
rect 7876 10031 9278 10133
rect 7876 9997 7880 10031
rect 7880 9997 7914 10031
rect 7914 9997 8016 10031
rect 8016 9997 8050 10031
rect 8050 9997 8152 10031
rect 8152 9997 8186 10031
rect 8186 9997 8288 10031
rect 8288 9997 8322 10031
rect 8322 9997 8424 10031
rect 8424 9997 8458 10031
rect 8458 9997 8560 10031
rect 8560 9997 8594 10031
rect 8594 9997 8696 10031
rect 8696 9997 8730 10031
rect 8730 9997 8832 10031
rect 8832 9997 8866 10031
rect 8866 9997 8968 10031
rect 8968 9997 9002 10031
rect 9002 9997 9104 10031
rect 9104 9997 9138 10031
rect 9138 9997 9240 10031
rect 9240 9997 9274 10031
rect 9274 9997 9278 10031
rect 7876 9895 9278 9997
rect 7876 9861 7880 9895
rect 7880 9861 7914 9895
rect 7914 9861 8016 9895
rect 8016 9861 8050 9895
rect 8050 9861 8152 9895
rect 8152 9861 8186 9895
rect 8186 9861 8288 9895
rect 8288 9861 8322 9895
rect 8322 9861 8424 9895
rect 8424 9861 8458 9895
rect 8458 9861 8560 9895
rect 8560 9861 8594 9895
rect 8594 9861 8696 9895
rect 8696 9861 8730 9895
rect 8730 9861 8832 9895
rect 8832 9861 8866 9895
rect 8866 9861 8968 9895
rect 8968 9861 9002 9895
rect 9002 9861 9104 9895
rect 9104 9861 9138 9895
rect 9138 9861 9240 9895
rect 9240 9861 9274 9895
rect 9274 9861 9278 9895
rect 7876 9759 9278 9861
rect 7876 9725 7880 9759
rect 7880 9725 7914 9759
rect 7914 9725 8016 9759
rect 8016 9725 8050 9759
rect 8050 9725 8152 9759
rect 8152 9725 8186 9759
rect 8186 9725 8288 9759
rect 8288 9725 8322 9759
rect 8322 9725 8424 9759
rect 8424 9725 8458 9759
rect 8458 9725 8560 9759
rect 8560 9725 8594 9759
rect 8594 9725 8696 9759
rect 8696 9725 8730 9759
rect 8730 9725 8832 9759
rect 8832 9725 8866 9759
rect 8866 9725 8968 9759
rect 8968 9725 9002 9759
rect 9002 9725 9104 9759
rect 9104 9725 9138 9759
rect 9138 9725 9240 9759
rect 9240 9725 9274 9759
rect 9274 9725 9278 9759
rect 7876 9623 9278 9725
rect 7876 9589 7880 9623
rect 7880 9589 7914 9623
rect 7914 9589 8016 9623
rect 8016 9589 8050 9623
rect 8050 9589 8152 9623
rect 8152 9589 8186 9623
rect 8186 9589 8288 9623
rect 8288 9589 8322 9623
rect 8322 9589 8424 9623
rect 8424 9589 8458 9623
rect 8458 9589 8560 9623
rect 8560 9589 8594 9623
rect 8594 9589 8696 9623
rect 8696 9589 8730 9623
rect 8730 9589 8832 9623
rect 8832 9589 8866 9623
rect 8866 9589 8968 9623
rect 8968 9589 9002 9623
rect 9002 9589 9104 9623
rect 9104 9589 9138 9623
rect 9138 9589 9240 9623
rect 9240 9589 9274 9623
rect 9274 9589 9278 9623
rect 7876 9487 9278 9589
rect 7876 9453 7880 9487
rect 7880 9453 7914 9487
rect 7914 9453 8016 9487
rect 8016 9453 8050 9487
rect 8050 9453 8152 9487
rect 8152 9453 8186 9487
rect 8186 9453 8288 9487
rect 8288 9453 8322 9487
rect 8322 9453 8424 9487
rect 8424 9453 8458 9487
rect 8458 9453 8560 9487
rect 8560 9453 8594 9487
rect 8594 9453 8696 9487
rect 8696 9453 8730 9487
rect 8730 9453 8832 9487
rect 8832 9453 8866 9487
rect 8866 9453 8968 9487
rect 8968 9453 9002 9487
rect 9002 9453 9104 9487
rect 9104 9453 9138 9487
rect 9138 9453 9240 9487
rect 9240 9453 9274 9487
rect 9274 9453 9278 9487
rect 7876 9351 9278 9453
rect 7876 9317 7880 9351
rect 7880 9317 7914 9351
rect 7914 9317 8016 9351
rect 8016 9317 8050 9351
rect 8050 9317 8152 9351
rect 8152 9317 8186 9351
rect 8186 9317 8288 9351
rect 8288 9317 8322 9351
rect 8322 9317 8424 9351
rect 8424 9317 8458 9351
rect 8458 9317 8560 9351
rect 8560 9317 8594 9351
rect 8594 9317 8696 9351
rect 8696 9317 8730 9351
rect 8730 9317 8832 9351
rect 8832 9317 8866 9351
rect 8866 9317 8968 9351
rect 8968 9317 9002 9351
rect 9002 9317 9104 9351
rect 9104 9317 9138 9351
rect 9138 9317 9240 9351
rect 9240 9317 9274 9351
rect 9274 9317 9278 9351
rect 7876 9215 9278 9317
rect 7876 9181 7880 9215
rect 7880 9181 7914 9215
rect 7914 9181 8016 9215
rect 8016 9181 8050 9215
rect 8050 9181 8152 9215
rect 8152 9181 8186 9215
rect 8186 9181 8288 9215
rect 8288 9181 8322 9215
rect 8322 9181 8424 9215
rect 8424 9181 8458 9215
rect 8458 9181 8560 9215
rect 8560 9181 8594 9215
rect 8594 9181 8696 9215
rect 8696 9181 8730 9215
rect 8730 9181 8832 9215
rect 8832 9181 8866 9215
rect 8866 9181 8968 9215
rect 8968 9181 9002 9215
rect 9002 9181 9104 9215
rect 9104 9181 9138 9215
rect 9138 9181 9240 9215
rect 9240 9181 9274 9215
rect 9274 9181 9278 9215
rect 7876 9079 9278 9181
rect 7876 9045 7880 9079
rect 7880 9045 7914 9079
rect 7914 9045 8016 9079
rect 8016 9045 8050 9079
rect 8050 9045 8152 9079
rect 8152 9045 8186 9079
rect 8186 9045 8288 9079
rect 8288 9045 8322 9079
rect 8322 9045 8424 9079
rect 8424 9045 8458 9079
rect 8458 9045 8560 9079
rect 8560 9045 8594 9079
rect 8594 9045 8696 9079
rect 8696 9045 8730 9079
rect 8730 9045 8832 9079
rect 8832 9045 8866 9079
rect 8866 9045 8968 9079
rect 8968 9045 9002 9079
rect 9002 9045 9104 9079
rect 9104 9045 9138 9079
rect 9138 9045 9240 9079
rect 9240 9045 9274 9079
rect 9274 9045 9278 9079
rect 7876 8943 9278 9045
rect 7876 8909 7880 8943
rect 7880 8909 7914 8943
rect 7914 8909 8016 8943
rect 8016 8909 8050 8943
rect 8050 8909 8152 8943
rect 8152 8909 8186 8943
rect 8186 8909 8288 8943
rect 8288 8909 8322 8943
rect 8322 8909 8424 8943
rect 8424 8909 8458 8943
rect 8458 8909 8560 8943
rect 8560 8909 8594 8943
rect 8594 8909 8696 8943
rect 8696 8909 8730 8943
rect 8730 8909 8832 8943
rect 8832 8909 8866 8943
rect 8866 8909 8968 8943
rect 8968 8909 9002 8943
rect 9002 8909 9104 8943
rect 9104 8909 9138 8943
rect 9138 8909 9240 8943
rect 9240 8909 9274 8943
rect 9274 8909 9278 8943
rect 7876 8807 9278 8909
rect 7876 8773 7880 8807
rect 7880 8773 7914 8807
rect 7914 8773 8016 8807
rect 8016 8773 8050 8807
rect 8050 8773 8152 8807
rect 8152 8773 8186 8807
rect 8186 8773 8288 8807
rect 8288 8773 8322 8807
rect 8322 8773 8424 8807
rect 8424 8773 8458 8807
rect 8458 8773 8560 8807
rect 8560 8773 8594 8807
rect 8594 8773 8696 8807
rect 8696 8773 8730 8807
rect 8730 8773 8832 8807
rect 8832 8773 8866 8807
rect 8866 8773 8968 8807
rect 8968 8773 9002 8807
rect 9002 8773 9104 8807
rect 9104 8773 9138 8807
rect 9138 8773 9240 8807
rect 9240 8773 9274 8807
rect 9274 8773 9278 8807
rect 7876 8671 9278 8773
rect 7876 8637 7880 8671
rect 7880 8637 7914 8671
rect 7914 8637 8016 8671
rect 8016 8637 8050 8671
rect 8050 8637 8152 8671
rect 8152 8637 8186 8671
rect 8186 8637 8288 8671
rect 8288 8637 8322 8671
rect 8322 8637 8424 8671
rect 8424 8637 8458 8671
rect 8458 8637 8560 8671
rect 8560 8637 8594 8671
rect 8594 8637 8696 8671
rect 8696 8637 8730 8671
rect 8730 8637 8832 8671
rect 8832 8637 8866 8671
rect 8866 8637 8968 8671
rect 8968 8637 9002 8671
rect 9002 8637 9104 8671
rect 9104 8637 9138 8671
rect 9138 8637 9240 8671
rect 9240 8637 9274 8671
rect 9274 8637 9278 8671
rect 7876 8535 9278 8637
rect 7876 8501 7880 8535
rect 7880 8501 7914 8535
rect 7914 8501 8016 8535
rect 8016 8501 8050 8535
rect 8050 8501 8152 8535
rect 8152 8501 8186 8535
rect 8186 8501 8288 8535
rect 8288 8501 8322 8535
rect 8322 8501 8424 8535
rect 8424 8501 8458 8535
rect 8458 8501 8560 8535
rect 8560 8501 8594 8535
rect 8594 8501 8696 8535
rect 8696 8501 8730 8535
rect 8730 8501 8832 8535
rect 8832 8501 8866 8535
rect 8866 8501 8968 8535
rect 8968 8501 9002 8535
rect 9002 8501 9104 8535
rect 9104 8501 9138 8535
rect 9138 8501 9240 8535
rect 9240 8501 9274 8535
rect 9274 8501 9278 8535
rect 7876 8399 9278 8501
rect 7876 8365 7880 8399
rect 7880 8365 7914 8399
rect 7914 8365 8016 8399
rect 8016 8365 8050 8399
rect 8050 8365 8152 8399
rect 8152 8365 8186 8399
rect 8186 8365 8288 8399
rect 8288 8365 8322 8399
rect 8322 8365 8424 8399
rect 8424 8365 8458 8399
rect 8458 8365 8560 8399
rect 8560 8365 8594 8399
rect 8594 8365 8696 8399
rect 8696 8365 8730 8399
rect 8730 8365 8832 8399
rect 8832 8365 8866 8399
rect 8866 8365 8968 8399
rect 8968 8365 9002 8399
rect 9002 8365 9104 8399
rect 9104 8365 9138 8399
rect 9138 8365 9240 8399
rect 9240 8365 9274 8399
rect 9274 8365 9278 8399
rect 7876 8263 9278 8365
rect 7876 8229 7880 8263
rect 7880 8229 7914 8263
rect 7914 8229 8016 8263
rect 8016 8229 8050 8263
rect 8050 8229 8152 8263
rect 8152 8229 8186 8263
rect 8186 8229 8288 8263
rect 8288 8229 8322 8263
rect 8322 8229 8424 8263
rect 8424 8229 8458 8263
rect 8458 8229 8560 8263
rect 8560 8229 8594 8263
rect 8594 8229 8696 8263
rect 8696 8229 8730 8263
rect 8730 8229 8832 8263
rect 8832 8229 8866 8263
rect 8866 8229 8968 8263
rect 8968 8229 9002 8263
rect 9002 8229 9104 8263
rect 9104 8229 9138 8263
rect 9138 8229 9240 8263
rect 9240 8229 9274 8263
rect 9274 8229 9278 8263
rect 7876 8127 9278 8229
rect 7876 8093 7880 8127
rect 7880 8093 7914 8127
rect 7914 8093 8016 8127
rect 8016 8093 8050 8127
rect 8050 8093 8152 8127
rect 8152 8093 8186 8127
rect 8186 8093 8288 8127
rect 8288 8093 8322 8127
rect 8322 8093 8424 8127
rect 8424 8093 8458 8127
rect 8458 8093 8560 8127
rect 8560 8093 8594 8127
rect 8594 8093 8696 8127
rect 8696 8093 8730 8127
rect 8730 8093 8832 8127
rect 8832 8093 8866 8127
rect 8866 8093 8968 8127
rect 8968 8093 9002 8127
rect 9002 8093 9104 8127
rect 9104 8093 9138 8127
rect 9138 8093 9240 8127
rect 9240 8093 9274 8127
rect 9274 8093 9278 8127
rect 7876 7991 9278 8093
rect 7876 7957 7880 7991
rect 7880 7957 7914 7991
rect 7914 7957 8016 7991
rect 8016 7957 8050 7991
rect 8050 7957 8152 7991
rect 8152 7957 8186 7991
rect 8186 7957 8288 7991
rect 8288 7957 8322 7991
rect 8322 7957 8424 7991
rect 8424 7957 8458 7991
rect 8458 7957 8560 7991
rect 8560 7957 8594 7991
rect 8594 7957 8696 7991
rect 8696 7957 8730 7991
rect 8730 7957 8832 7991
rect 8832 7957 8866 7991
rect 8866 7957 8968 7991
rect 8968 7957 9002 7991
rect 9002 7957 9104 7991
rect 9104 7957 9138 7991
rect 9138 7957 9240 7991
rect 9240 7957 9274 7991
rect 9274 7957 9278 7991
rect 7876 7855 9278 7957
rect 7876 7821 7880 7855
rect 7880 7821 7914 7855
rect 7914 7821 8016 7855
rect 8016 7821 8050 7855
rect 8050 7821 8152 7855
rect 8152 7821 8186 7855
rect 8186 7821 8288 7855
rect 8288 7821 8322 7855
rect 8322 7821 8424 7855
rect 8424 7821 8458 7855
rect 8458 7821 8560 7855
rect 8560 7821 8594 7855
rect 8594 7821 8696 7855
rect 8696 7821 8730 7855
rect 8730 7821 8832 7855
rect 8832 7821 8866 7855
rect 8866 7821 8968 7855
rect 8968 7821 9002 7855
rect 9002 7821 9104 7855
rect 9104 7821 9138 7855
rect 9138 7821 9240 7855
rect 9240 7821 9274 7855
rect 9274 7821 9278 7855
rect 7876 7719 9278 7821
rect 7876 7685 7880 7719
rect 7880 7685 7914 7719
rect 7914 7685 8016 7719
rect 8016 7685 8050 7719
rect 8050 7685 8152 7719
rect 8152 7685 8186 7719
rect 8186 7685 8288 7719
rect 8288 7685 8322 7719
rect 8322 7685 8424 7719
rect 8424 7685 8458 7719
rect 8458 7685 8560 7719
rect 8560 7685 8594 7719
rect 8594 7685 8696 7719
rect 8696 7685 8730 7719
rect 8730 7685 8832 7719
rect 8832 7685 8866 7719
rect 8866 7685 8968 7719
rect 8968 7685 9002 7719
rect 9002 7685 9104 7719
rect 9104 7685 9138 7719
rect 9138 7685 9240 7719
rect 9240 7685 9274 7719
rect 9274 7685 9278 7719
rect 7876 7583 9278 7685
rect 7876 7549 7880 7583
rect 7880 7549 7914 7583
rect 7914 7549 8016 7583
rect 8016 7549 8050 7583
rect 8050 7549 8152 7583
rect 8152 7549 8186 7583
rect 8186 7549 8288 7583
rect 8288 7549 8322 7583
rect 8322 7549 8424 7583
rect 8424 7549 8458 7583
rect 8458 7549 8560 7583
rect 8560 7549 8594 7583
rect 8594 7549 8696 7583
rect 8696 7549 8730 7583
rect 8730 7549 8832 7583
rect 8832 7549 8866 7583
rect 8866 7549 8968 7583
rect 8968 7549 9002 7583
rect 9002 7549 9104 7583
rect 9104 7549 9138 7583
rect 9138 7549 9240 7583
rect 9240 7549 9274 7583
rect 9274 7549 9278 7583
rect 7876 7447 9278 7549
rect 7876 7413 7880 7447
rect 7880 7413 7914 7447
rect 7914 7413 8016 7447
rect 8016 7413 8050 7447
rect 8050 7413 8152 7447
rect 8152 7413 8186 7447
rect 8186 7413 8288 7447
rect 8288 7413 8322 7447
rect 8322 7413 8424 7447
rect 8424 7413 8458 7447
rect 8458 7413 8560 7447
rect 8560 7413 8594 7447
rect 8594 7413 8696 7447
rect 8696 7413 8730 7447
rect 8730 7413 8832 7447
rect 8832 7413 8866 7447
rect 8866 7413 8968 7447
rect 8968 7413 9002 7447
rect 9002 7413 9104 7447
rect 9104 7413 9138 7447
rect 9138 7413 9240 7447
rect 9240 7413 9274 7447
rect 9274 7413 9278 7447
rect 7876 7311 9278 7413
rect 7876 7277 7880 7311
rect 7880 7277 7914 7311
rect 7914 7277 8016 7311
rect 8016 7277 8050 7311
rect 8050 7277 8152 7311
rect 8152 7277 8186 7311
rect 8186 7277 8288 7311
rect 8288 7277 8322 7311
rect 8322 7277 8424 7311
rect 8424 7277 8458 7311
rect 8458 7277 8560 7311
rect 8560 7277 8594 7311
rect 8594 7277 8696 7311
rect 8696 7277 8730 7311
rect 8730 7277 8832 7311
rect 8832 7277 8866 7311
rect 8866 7277 8968 7311
rect 8968 7277 9002 7311
rect 9002 7277 9104 7311
rect 9104 7277 9138 7311
rect 9138 7277 9240 7311
rect 9240 7277 9274 7311
rect 9274 7277 9278 7311
rect 7876 7175 9278 7277
rect 7876 7141 7880 7175
rect 7880 7141 7914 7175
rect 7914 7141 8016 7175
rect 8016 7141 8050 7175
rect 8050 7141 8152 7175
rect 8152 7141 8186 7175
rect 8186 7141 8288 7175
rect 8288 7141 8322 7175
rect 8322 7141 8424 7175
rect 8424 7141 8458 7175
rect 8458 7141 8560 7175
rect 8560 7141 8594 7175
rect 8594 7141 8696 7175
rect 8696 7141 8730 7175
rect 8730 7141 8832 7175
rect 8832 7141 8866 7175
rect 8866 7141 8968 7175
rect 8968 7141 9002 7175
rect 9002 7141 9104 7175
rect 9104 7141 9138 7175
rect 9138 7141 9240 7175
rect 9240 7141 9274 7175
rect 9274 7141 9278 7175
rect 7876 7039 9278 7141
rect 7876 7005 7880 7039
rect 7880 7005 7914 7039
rect 7914 7005 8016 7039
rect 8016 7005 8050 7039
rect 8050 7005 8152 7039
rect 8152 7005 8186 7039
rect 8186 7005 8288 7039
rect 8288 7005 8322 7039
rect 8322 7005 8424 7039
rect 8424 7005 8458 7039
rect 8458 7005 8560 7039
rect 8560 7005 8594 7039
rect 8594 7005 8696 7039
rect 8696 7005 8730 7039
rect 8730 7005 8832 7039
rect 8832 7005 8866 7039
rect 8866 7005 8968 7039
rect 8968 7005 9002 7039
rect 9002 7005 9104 7039
rect 9104 7005 9138 7039
rect 9138 7005 9240 7039
rect 9240 7005 9274 7039
rect 9274 7005 9278 7039
rect 7876 6903 9278 7005
rect 7876 6869 7880 6903
rect 7880 6869 7914 6903
rect 7914 6869 8016 6903
rect 8016 6869 8050 6903
rect 8050 6869 8152 6903
rect 8152 6869 8186 6903
rect 8186 6869 8288 6903
rect 8288 6869 8322 6903
rect 8322 6869 8424 6903
rect 8424 6869 8458 6903
rect 8458 6869 8560 6903
rect 8560 6869 8594 6903
rect 8594 6869 8696 6903
rect 8696 6869 8730 6903
rect 8730 6869 8832 6903
rect 8832 6869 8866 6903
rect 8866 6869 8968 6903
rect 8968 6869 9002 6903
rect 9002 6869 9104 6903
rect 9104 6869 9138 6903
rect 9138 6869 9240 6903
rect 9240 6869 9274 6903
rect 9274 6869 9278 6903
rect 7876 6767 9278 6869
rect 7876 6733 7880 6767
rect 7880 6733 7914 6767
rect 7914 6733 8016 6767
rect 8016 6733 8050 6767
rect 8050 6733 8152 6767
rect 8152 6733 8186 6767
rect 8186 6733 8288 6767
rect 8288 6733 8322 6767
rect 8322 6733 8424 6767
rect 8424 6733 8458 6767
rect 8458 6733 8560 6767
rect 8560 6733 8594 6767
rect 8594 6733 8696 6767
rect 8696 6733 8730 6767
rect 8730 6733 8832 6767
rect 8832 6733 8866 6767
rect 8866 6733 8968 6767
rect 8968 6733 9002 6767
rect 9002 6733 9104 6767
rect 9104 6733 9138 6767
rect 9138 6733 9240 6767
rect 9240 6733 9274 6767
rect 9274 6733 9278 6767
rect 7876 6631 9278 6733
rect 7876 6597 7880 6631
rect 7880 6597 7914 6631
rect 7914 6597 8016 6631
rect 8016 6597 8050 6631
rect 8050 6597 8152 6631
rect 8152 6597 8186 6631
rect 8186 6597 8288 6631
rect 8288 6597 8322 6631
rect 8322 6597 8424 6631
rect 8424 6597 8458 6631
rect 8458 6597 8560 6631
rect 8560 6597 8594 6631
rect 8594 6597 8696 6631
rect 8696 6597 8730 6631
rect 8730 6597 8832 6631
rect 8832 6597 8866 6631
rect 8866 6597 8968 6631
rect 8968 6597 9002 6631
rect 9002 6597 9104 6631
rect 9104 6597 9138 6631
rect 9138 6597 9240 6631
rect 9240 6597 9274 6631
rect 9274 6597 9278 6631
rect 7876 6495 9278 6597
rect 7876 6461 7880 6495
rect 7880 6461 7914 6495
rect 7914 6461 8016 6495
rect 8016 6461 8050 6495
rect 8050 6461 8152 6495
rect 8152 6461 8186 6495
rect 8186 6461 8288 6495
rect 8288 6461 8322 6495
rect 8322 6461 8424 6495
rect 8424 6461 8458 6495
rect 8458 6461 8560 6495
rect 8560 6461 8594 6495
rect 8594 6461 8696 6495
rect 8696 6461 8730 6495
rect 8730 6461 8832 6495
rect 8832 6461 8866 6495
rect 8866 6461 8968 6495
rect 8968 6461 9002 6495
rect 9002 6461 9104 6495
rect 9104 6461 9138 6495
rect 9138 6461 9240 6495
rect 9240 6461 9274 6495
rect 9274 6461 9278 6495
rect 7876 6359 9278 6461
rect 7876 6325 7880 6359
rect 7880 6325 7914 6359
rect 7914 6325 8016 6359
rect 8016 6325 8050 6359
rect 8050 6325 8152 6359
rect 8152 6325 8186 6359
rect 8186 6325 8288 6359
rect 8288 6325 8322 6359
rect 8322 6325 8424 6359
rect 8424 6325 8458 6359
rect 8458 6325 8560 6359
rect 8560 6325 8594 6359
rect 8594 6325 8696 6359
rect 8696 6325 8730 6359
rect 8730 6325 8832 6359
rect 8832 6325 8866 6359
rect 8866 6325 8968 6359
rect 8968 6325 9002 6359
rect 9002 6325 9104 6359
rect 9104 6325 9138 6359
rect 9138 6325 9240 6359
rect 9240 6325 9274 6359
rect 9274 6325 9278 6359
rect 7876 6223 9278 6325
rect 7876 6189 7880 6223
rect 7880 6189 7914 6223
rect 7914 6189 8016 6223
rect 8016 6189 8050 6223
rect 8050 6189 8152 6223
rect 8152 6189 8186 6223
rect 8186 6189 8288 6223
rect 8288 6189 8322 6223
rect 8322 6189 8424 6223
rect 8424 6189 8458 6223
rect 8458 6189 8560 6223
rect 8560 6189 8594 6223
rect 8594 6189 8696 6223
rect 8696 6189 8730 6223
rect 8730 6189 8832 6223
rect 8832 6189 8866 6223
rect 8866 6189 8968 6223
rect 8968 6189 9002 6223
rect 9002 6189 9104 6223
rect 9104 6189 9138 6223
rect 9138 6189 9240 6223
rect 9240 6189 9274 6223
rect 9274 6189 9278 6223
rect 7876 6087 9278 6189
rect 7876 6053 7880 6087
rect 7880 6053 7914 6087
rect 7914 6053 8016 6087
rect 8016 6053 8050 6087
rect 8050 6053 8152 6087
rect 8152 6053 8186 6087
rect 8186 6053 8288 6087
rect 8288 6053 8322 6087
rect 8322 6053 8424 6087
rect 8424 6053 8458 6087
rect 8458 6053 8560 6087
rect 8560 6053 8594 6087
rect 8594 6053 8696 6087
rect 8696 6053 8730 6087
rect 8730 6053 8832 6087
rect 8832 6053 8866 6087
rect 8866 6053 8968 6087
rect 8968 6053 9002 6087
rect 9002 6053 9104 6087
rect 9104 6053 9138 6087
rect 9138 6053 9240 6087
rect 9240 6053 9274 6087
rect 9274 6053 9278 6087
rect 7876 5951 9278 6053
rect 7876 5917 7880 5951
rect 7880 5917 7914 5951
rect 7914 5917 8016 5951
rect 8016 5917 8050 5951
rect 8050 5917 8152 5951
rect 8152 5917 8186 5951
rect 8186 5917 8288 5951
rect 8288 5917 8322 5951
rect 8322 5917 8424 5951
rect 8424 5917 8458 5951
rect 8458 5917 8560 5951
rect 8560 5917 8594 5951
rect 8594 5917 8696 5951
rect 8696 5917 8730 5951
rect 8730 5917 8832 5951
rect 8832 5917 8866 5951
rect 8866 5917 8968 5951
rect 8968 5917 9002 5951
rect 9002 5917 9104 5951
rect 9104 5917 9138 5951
rect 9138 5917 9240 5951
rect 9240 5917 9274 5951
rect 9274 5917 9278 5951
rect 7876 5815 9278 5917
rect 7876 5781 7880 5815
rect 7880 5781 7914 5815
rect 7914 5781 8016 5815
rect 8016 5781 8050 5815
rect 8050 5781 8152 5815
rect 8152 5781 8186 5815
rect 8186 5781 8288 5815
rect 8288 5781 8322 5815
rect 8322 5781 8424 5815
rect 8424 5781 8458 5815
rect 8458 5781 8560 5815
rect 8560 5781 8594 5815
rect 8594 5781 8696 5815
rect 8696 5781 8730 5815
rect 8730 5781 8832 5815
rect 8832 5781 8866 5815
rect 8866 5781 8968 5815
rect 8968 5781 9002 5815
rect 9002 5781 9104 5815
rect 9104 5781 9138 5815
rect 9138 5781 9240 5815
rect 9240 5781 9274 5815
rect 9274 5781 9278 5815
rect 7876 5679 9278 5781
rect 7876 5645 7880 5679
rect 7880 5645 7914 5679
rect 7914 5645 8016 5679
rect 8016 5645 8050 5679
rect 8050 5645 8152 5679
rect 8152 5645 8186 5679
rect 8186 5645 8288 5679
rect 8288 5645 8322 5679
rect 8322 5645 8424 5679
rect 8424 5645 8458 5679
rect 8458 5645 8560 5679
rect 8560 5645 8594 5679
rect 8594 5645 8696 5679
rect 8696 5645 8730 5679
rect 8730 5645 8832 5679
rect 8832 5645 8866 5679
rect 8866 5645 8968 5679
rect 8968 5645 9002 5679
rect 9002 5645 9104 5679
rect 9104 5645 9138 5679
rect 9138 5645 9240 5679
rect 9240 5645 9274 5679
rect 9274 5645 9278 5679
rect 7876 5543 9278 5645
rect 7876 5509 7880 5543
rect 7880 5509 7914 5543
rect 7914 5509 8016 5543
rect 8016 5509 8050 5543
rect 8050 5509 8152 5543
rect 8152 5509 8186 5543
rect 8186 5509 8288 5543
rect 8288 5509 8322 5543
rect 8322 5509 8424 5543
rect 8424 5509 8458 5543
rect 8458 5509 8560 5543
rect 8560 5509 8594 5543
rect 8594 5509 8696 5543
rect 8696 5509 8730 5543
rect 8730 5509 8832 5543
rect 8832 5509 8866 5543
rect 8866 5509 8968 5543
rect 8968 5509 9002 5543
rect 9002 5509 9104 5543
rect 9104 5509 9138 5543
rect 9138 5509 9240 5543
rect 9240 5509 9274 5543
rect 9274 5509 9278 5543
rect 7876 5407 9278 5509
rect 7876 5373 7880 5407
rect 7880 5373 7914 5407
rect 7914 5373 8016 5407
rect 8016 5373 8050 5407
rect 8050 5373 8152 5407
rect 8152 5373 8186 5407
rect 8186 5373 8288 5407
rect 8288 5373 8322 5407
rect 8322 5373 8424 5407
rect 8424 5373 8458 5407
rect 8458 5373 8560 5407
rect 8560 5373 8594 5407
rect 8594 5373 8696 5407
rect 8696 5373 8730 5407
rect 8730 5373 8832 5407
rect 8832 5373 8866 5407
rect 8866 5373 8968 5407
rect 8968 5373 9002 5407
rect 9002 5373 9104 5407
rect 9104 5373 9138 5407
rect 9138 5373 9240 5407
rect 9240 5373 9274 5407
rect 9274 5373 9278 5407
rect 7876 5271 9278 5373
rect 7876 5237 7880 5271
rect 7880 5237 7914 5271
rect 7914 5237 8016 5271
rect 8016 5237 8050 5271
rect 8050 5237 8152 5271
rect 8152 5237 8186 5271
rect 8186 5237 8288 5271
rect 8288 5237 8322 5271
rect 8322 5237 8424 5271
rect 8424 5237 8458 5271
rect 8458 5237 8560 5271
rect 8560 5237 8594 5271
rect 8594 5237 8696 5271
rect 8696 5237 8730 5271
rect 8730 5237 8832 5271
rect 8832 5237 8866 5271
rect 8866 5237 8968 5271
rect 8968 5237 9002 5271
rect 9002 5237 9104 5271
rect 9104 5237 9138 5271
rect 9138 5237 9240 5271
rect 9240 5237 9274 5271
rect 9274 5237 9278 5271
rect 7876 5135 9278 5237
rect 7876 5101 7880 5135
rect 7880 5101 7914 5135
rect 7914 5101 8016 5135
rect 8016 5101 8050 5135
rect 8050 5101 8152 5135
rect 8152 5101 8186 5135
rect 8186 5101 8288 5135
rect 8288 5101 8322 5135
rect 8322 5101 8424 5135
rect 8424 5101 8458 5135
rect 8458 5101 8560 5135
rect 8560 5101 8594 5135
rect 8594 5101 8696 5135
rect 8696 5101 8730 5135
rect 8730 5101 8832 5135
rect 8832 5101 8866 5135
rect 8866 5101 8968 5135
rect 8968 5101 9002 5135
rect 9002 5101 9104 5135
rect 9104 5101 9138 5135
rect 9138 5101 9240 5135
rect 9240 5101 9274 5135
rect 9274 5101 9278 5135
rect 7876 4999 9278 5101
rect 7876 4965 7880 4999
rect 7880 4965 7914 4999
rect 7914 4965 8016 4999
rect 8016 4965 8050 4999
rect 8050 4965 8152 4999
rect 8152 4965 8186 4999
rect 8186 4965 8288 4999
rect 8288 4965 8322 4999
rect 8322 4965 8424 4999
rect 8424 4965 8458 4999
rect 8458 4965 8560 4999
rect 8560 4965 8594 4999
rect 8594 4965 8696 4999
rect 8696 4965 8730 4999
rect 8730 4965 8832 4999
rect 8832 4965 8866 4999
rect 8866 4965 8968 4999
rect 8968 4965 9002 4999
rect 9002 4965 9104 4999
rect 9104 4965 9138 4999
rect 9138 4965 9240 4999
rect 9240 4965 9274 4999
rect 9274 4965 9278 4999
rect 7876 4863 9278 4965
rect 7876 4829 7880 4863
rect 7880 4829 7914 4863
rect 7914 4829 8016 4863
rect 8016 4829 8050 4863
rect 8050 4829 8152 4863
rect 8152 4829 8186 4863
rect 8186 4829 8288 4863
rect 8288 4829 8322 4863
rect 8322 4829 8424 4863
rect 8424 4829 8458 4863
rect 8458 4829 8560 4863
rect 8560 4829 8594 4863
rect 8594 4829 8696 4863
rect 8696 4829 8730 4863
rect 8730 4829 8832 4863
rect 8832 4829 8866 4863
rect 8866 4829 8968 4863
rect 8968 4829 9002 4863
rect 9002 4829 9104 4863
rect 9104 4829 9138 4863
rect 9138 4829 9240 4863
rect 9240 4829 9274 4863
rect 9274 4829 9278 4863
rect 7876 4727 9278 4829
rect 7876 4693 7880 4727
rect 7880 4693 7914 4727
rect 7914 4693 8016 4727
rect 8016 4693 8050 4727
rect 8050 4693 8152 4727
rect 8152 4693 8186 4727
rect 8186 4693 8288 4727
rect 8288 4693 8322 4727
rect 8322 4693 8424 4727
rect 8424 4693 8458 4727
rect 8458 4693 8560 4727
rect 8560 4693 8594 4727
rect 8594 4693 8696 4727
rect 8696 4693 8730 4727
rect 8730 4693 8832 4727
rect 8832 4693 8866 4727
rect 8866 4693 8968 4727
rect 8968 4693 9002 4727
rect 9002 4693 9104 4727
rect 9104 4693 9138 4727
rect 9138 4693 9240 4727
rect 9240 4693 9274 4727
rect 9274 4693 9278 4727
rect 7876 4591 9278 4693
rect 7876 4557 7880 4591
rect 7880 4557 7914 4591
rect 7914 4557 8016 4591
rect 8016 4557 8050 4591
rect 8050 4557 8152 4591
rect 8152 4557 8186 4591
rect 8186 4557 8288 4591
rect 8288 4557 8322 4591
rect 8322 4557 8424 4591
rect 8424 4557 8458 4591
rect 8458 4557 8560 4591
rect 8560 4557 8594 4591
rect 8594 4557 8696 4591
rect 8696 4557 8730 4591
rect 8730 4557 8832 4591
rect 8832 4557 8866 4591
rect 8866 4557 8968 4591
rect 8968 4557 9002 4591
rect 9002 4557 9104 4591
rect 9104 4557 9138 4591
rect 9138 4557 9240 4591
rect 9240 4557 9274 4591
rect 9274 4557 9278 4591
rect 7876 4455 9278 4557
rect 7876 4421 7880 4455
rect 7880 4421 7914 4455
rect 7914 4421 8016 4455
rect 8016 4421 8050 4455
rect 8050 4421 8152 4455
rect 8152 4421 8186 4455
rect 8186 4421 8288 4455
rect 8288 4421 8322 4455
rect 8322 4421 8424 4455
rect 8424 4421 8458 4455
rect 8458 4421 8560 4455
rect 8560 4421 8594 4455
rect 8594 4421 8696 4455
rect 8696 4421 8730 4455
rect 8730 4421 8832 4455
rect 8832 4421 8866 4455
rect 8866 4421 8968 4455
rect 8968 4421 9002 4455
rect 9002 4421 9104 4455
rect 9104 4421 9138 4455
rect 9138 4421 9240 4455
rect 9240 4421 9274 4455
rect 9274 4421 9278 4455
rect 7876 4319 9278 4421
rect 7876 4285 7880 4319
rect 7880 4285 7914 4319
rect 7914 4285 8016 4319
rect 8016 4285 8050 4319
rect 8050 4285 8152 4319
rect 8152 4285 8186 4319
rect 8186 4285 8288 4319
rect 8288 4285 8322 4319
rect 8322 4285 8424 4319
rect 8424 4285 8458 4319
rect 8458 4285 8560 4319
rect 8560 4285 8594 4319
rect 8594 4285 8696 4319
rect 8696 4285 8730 4319
rect 8730 4285 8832 4319
rect 8832 4285 8866 4319
rect 8866 4285 8968 4319
rect 8968 4285 9002 4319
rect 9002 4285 9104 4319
rect 9104 4285 9138 4319
rect 9138 4285 9240 4319
rect 9240 4285 9274 4319
rect 9274 4285 9278 4319
rect 7876 4183 9278 4285
rect 7876 4149 7880 4183
rect 7880 4149 7914 4183
rect 7914 4149 8016 4183
rect 8016 4149 8050 4183
rect 8050 4149 8152 4183
rect 8152 4149 8186 4183
rect 8186 4149 8288 4183
rect 8288 4149 8322 4183
rect 8322 4149 8424 4183
rect 8424 4149 8458 4183
rect 8458 4149 8560 4183
rect 8560 4149 8594 4183
rect 8594 4149 8696 4183
rect 8696 4149 8730 4183
rect 8730 4149 8832 4183
rect 8832 4149 8866 4183
rect 8866 4149 8968 4183
rect 8968 4149 9002 4183
rect 9002 4149 9104 4183
rect 9104 4149 9138 4183
rect 9138 4149 9240 4183
rect 9240 4149 9274 4183
rect 9274 4149 9278 4183
rect 7876 4047 9278 4149
rect 7876 4013 7880 4047
rect 7880 4013 7914 4047
rect 7914 4013 8016 4047
rect 8016 4013 8050 4047
rect 8050 4013 8152 4047
rect 8152 4013 8186 4047
rect 8186 4013 8288 4047
rect 8288 4013 8322 4047
rect 8322 4013 8424 4047
rect 8424 4013 8458 4047
rect 8458 4013 8560 4047
rect 8560 4013 8594 4047
rect 8594 4013 8696 4047
rect 8696 4013 8730 4047
rect 8730 4013 8832 4047
rect 8832 4013 8866 4047
rect 8866 4013 8968 4047
rect 8968 4013 9002 4047
rect 9002 4013 9104 4047
rect 9104 4013 9138 4047
rect 9138 4013 9240 4047
rect 9240 4013 9274 4047
rect 9274 4013 9278 4047
rect 7876 3911 9278 4013
rect 7876 3877 7880 3911
rect 7880 3877 7914 3911
rect 7914 3877 8016 3911
rect 8016 3877 8050 3911
rect 8050 3877 8152 3911
rect 8152 3877 8186 3911
rect 8186 3877 8288 3911
rect 8288 3877 8322 3911
rect 8322 3877 8424 3911
rect 8424 3877 8458 3911
rect 8458 3877 8560 3911
rect 8560 3877 8594 3911
rect 8594 3877 8696 3911
rect 8696 3877 8730 3911
rect 8730 3877 8832 3911
rect 8832 3877 8866 3911
rect 8866 3877 8968 3911
rect 8968 3877 9002 3911
rect 9002 3877 9104 3911
rect 9104 3877 9138 3911
rect 9138 3877 9240 3911
rect 9240 3877 9274 3911
rect 9274 3877 9278 3911
rect 7876 3775 9278 3877
rect 7876 3741 7880 3775
rect 7880 3741 7914 3775
rect 7914 3741 8016 3775
rect 8016 3741 8050 3775
rect 8050 3741 8152 3775
rect 8152 3741 8186 3775
rect 8186 3741 8288 3775
rect 8288 3741 8322 3775
rect 8322 3741 8424 3775
rect 8424 3741 8458 3775
rect 8458 3741 8560 3775
rect 8560 3741 8594 3775
rect 8594 3741 8696 3775
rect 8696 3741 8730 3775
rect 8730 3741 8832 3775
rect 8832 3741 8866 3775
rect 8866 3741 8968 3775
rect 8968 3741 9002 3775
rect 9002 3741 9104 3775
rect 9104 3741 9138 3775
rect 9138 3741 9240 3775
rect 9240 3741 9274 3775
rect 9274 3741 9278 3775
rect 7876 3639 9278 3741
rect 7876 3605 7880 3639
rect 7880 3605 7914 3639
rect 7914 3605 8016 3639
rect 8016 3605 8050 3639
rect 8050 3605 8152 3639
rect 8152 3605 8186 3639
rect 8186 3605 8288 3639
rect 8288 3605 8322 3639
rect 8322 3605 8424 3639
rect 8424 3605 8458 3639
rect 8458 3605 8560 3639
rect 8560 3605 8594 3639
rect 8594 3605 8696 3639
rect 8696 3605 8730 3639
rect 8730 3605 8832 3639
rect 8832 3605 8866 3639
rect 8866 3605 8968 3639
rect 8968 3605 9002 3639
rect 9002 3605 9104 3639
rect 9104 3605 9138 3639
rect 9138 3605 9240 3639
rect 9240 3605 9274 3639
rect 9274 3605 9278 3639
rect 7876 3503 9278 3605
rect 7876 3469 7880 3503
rect 7880 3469 7914 3503
rect 7914 3469 8016 3503
rect 8016 3469 8050 3503
rect 8050 3469 8152 3503
rect 8152 3469 8186 3503
rect 8186 3469 8288 3503
rect 8288 3469 8322 3503
rect 8322 3469 8424 3503
rect 8424 3469 8458 3503
rect 8458 3469 8560 3503
rect 8560 3469 8594 3503
rect 8594 3469 8696 3503
rect 8696 3469 8730 3503
rect 8730 3469 8832 3503
rect 8832 3469 8866 3503
rect 8866 3469 8968 3503
rect 8968 3469 9002 3503
rect 9002 3469 9104 3503
rect 9104 3469 9138 3503
rect 9138 3469 9240 3503
rect 9240 3469 9274 3503
rect 9274 3469 9278 3503
rect 7876 3367 9278 3469
rect 7876 3333 7880 3367
rect 7880 3333 7914 3367
rect 7914 3333 8016 3367
rect 8016 3333 8050 3367
rect 8050 3333 8152 3367
rect 8152 3333 8186 3367
rect 8186 3333 8288 3367
rect 8288 3333 8322 3367
rect 8322 3333 8424 3367
rect 8424 3333 8458 3367
rect 8458 3333 8560 3367
rect 8560 3333 8594 3367
rect 8594 3333 8696 3367
rect 8696 3333 8730 3367
rect 8730 3333 8832 3367
rect 8832 3333 8866 3367
rect 8866 3333 8968 3367
rect 8968 3333 9002 3367
rect 9002 3333 9104 3367
rect 9104 3333 9138 3367
rect 9138 3333 9240 3367
rect 9240 3333 9274 3367
rect 9274 3333 9278 3367
rect 7876 3231 9278 3333
rect 7876 3197 7880 3231
rect 7880 3197 7914 3231
rect 7914 3197 8016 3231
rect 8016 3197 8050 3231
rect 8050 3197 8152 3231
rect 8152 3197 8186 3231
rect 8186 3197 8288 3231
rect 8288 3197 8322 3231
rect 8322 3197 8424 3231
rect 8424 3197 8458 3231
rect 8458 3197 8560 3231
rect 8560 3197 8594 3231
rect 8594 3197 8696 3231
rect 8696 3197 8730 3231
rect 8730 3197 8832 3231
rect 8832 3197 8866 3231
rect 8866 3197 8968 3231
rect 8968 3197 9002 3231
rect 9002 3197 9104 3231
rect 9104 3197 9138 3231
rect 9138 3197 9240 3231
rect 9240 3197 9274 3231
rect 9274 3197 9278 3231
rect 7876 3095 9278 3197
rect 7876 3061 7880 3095
rect 7880 3061 7914 3095
rect 7914 3061 8016 3095
rect 8016 3061 8050 3095
rect 8050 3061 8152 3095
rect 8152 3061 8186 3095
rect 8186 3061 8288 3095
rect 8288 3061 8322 3095
rect 8322 3061 8424 3095
rect 8424 3061 8458 3095
rect 8458 3061 8560 3095
rect 8560 3061 8594 3095
rect 8594 3061 8696 3095
rect 8696 3061 8730 3095
rect 8730 3061 8832 3095
rect 8832 3061 8866 3095
rect 8866 3061 8968 3095
rect 8968 3061 9002 3095
rect 9002 3061 9104 3095
rect 9104 3061 9138 3095
rect 9138 3061 9240 3095
rect 9240 3061 9274 3095
rect 9274 3061 9278 3095
rect 7876 2959 9278 3061
rect 7876 2925 7880 2959
rect 7880 2925 7914 2959
rect 7914 2925 8016 2959
rect 8016 2925 8050 2959
rect 8050 2925 8152 2959
rect 8152 2925 8186 2959
rect 8186 2925 8288 2959
rect 8288 2925 8322 2959
rect 8322 2925 8424 2959
rect 8424 2925 8458 2959
rect 8458 2925 8560 2959
rect 8560 2925 8594 2959
rect 8594 2925 8696 2959
rect 8696 2925 8730 2959
rect 8730 2925 8832 2959
rect 8832 2925 8866 2959
rect 8866 2925 8968 2959
rect 8968 2925 9002 2959
rect 9002 2925 9104 2959
rect 9104 2925 9138 2959
rect 9138 2925 9240 2959
rect 9240 2925 9274 2959
rect 9274 2925 9278 2959
rect 7876 2823 9278 2925
rect 7876 2789 7880 2823
rect 7880 2789 7914 2823
rect 7914 2789 8016 2823
rect 8016 2789 8050 2823
rect 8050 2789 8152 2823
rect 8152 2789 8186 2823
rect 8186 2789 8288 2823
rect 8288 2789 8322 2823
rect 8322 2789 8424 2823
rect 8424 2789 8458 2823
rect 8458 2789 8560 2823
rect 8560 2789 8594 2823
rect 8594 2789 8696 2823
rect 8696 2789 8730 2823
rect 8730 2789 8832 2823
rect 8832 2789 8866 2823
rect 8866 2789 8968 2823
rect 8968 2789 9002 2823
rect 9002 2789 9104 2823
rect 9104 2789 9138 2823
rect 9138 2789 9240 2823
rect 9240 2789 9274 2823
rect 9274 2789 9278 2823
rect 7876 2687 9278 2789
rect 7876 2653 7880 2687
rect 7880 2653 7914 2687
rect 7914 2653 8016 2687
rect 8016 2653 8050 2687
rect 8050 2653 8152 2687
rect 8152 2653 8186 2687
rect 8186 2653 8288 2687
rect 8288 2653 8322 2687
rect 8322 2653 8424 2687
rect 8424 2653 8458 2687
rect 8458 2653 8560 2687
rect 8560 2653 8594 2687
rect 8594 2653 8696 2687
rect 8696 2653 8730 2687
rect 8730 2653 8832 2687
rect 8832 2653 8866 2687
rect 8866 2653 8968 2687
rect 8968 2653 9002 2687
rect 9002 2653 9104 2687
rect 9104 2653 9138 2687
rect 9138 2653 9240 2687
rect 9240 2653 9274 2687
rect 9274 2653 9278 2687
rect 7876 2551 9278 2653
rect 7876 2517 7880 2551
rect 7880 2517 7914 2551
rect 7914 2517 8016 2551
rect 8016 2517 8050 2551
rect 8050 2517 8152 2551
rect 8152 2517 8186 2551
rect 8186 2517 8288 2551
rect 8288 2517 8322 2551
rect 8322 2517 8424 2551
rect 8424 2517 8458 2551
rect 8458 2517 8560 2551
rect 8560 2517 8594 2551
rect 8594 2517 8696 2551
rect 8696 2517 8730 2551
rect 8730 2517 8832 2551
rect 8832 2517 8866 2551
rect 8866 2517 8968 2551
rect 8968 2517 9002 2551
rect 9002 2517 9104 2551
rect 9104 2517 9138 2551
rect 9138 2517 9240 2551
rect 9240 2517 9274 2551
rect 9274 2517 9278 2551
rect 7876 2414 9278 2517
rect 7876 2395 7880 2414
rect 7880 2395 7914 2414
rect 7914 2395 8016 2414
rect 8016 2395 8050 2414
rect 8050 2395 8152 2414
rect 8152 2395 8186 2414
rect 8186 2395 8288 2414
rect 8288 2395 8322 2414
rect 8322 2395 8424 2414
rect 8424 2395 8458 2414
rect 8458 2395 8560 2414
rect 8560 2395 8594 2414
rect 8594 2395 8696 2414
rect 8696 2395 8730 2414
rect 8730 2395 8832 2414
rect 8832 2395 8866 2414
rect 8866 2395 8968 2414
rect 8968 2395 9002 2414
rect 9002 2395 9104 2414
rect 9104 2395 9138 2414
rect 9138 2395 9240 2414
rect 9240 2395 9274 2414
rect 9274 2395 9278 2414
rect 7876 2322 7910 2356
rect 7948 2322 7982 2356
rect 8020 2322 8054 2356
rect 8092 2322 8126 2356
rect 8164 2322 8198 2356
rect 8236 2322 8270 2356
rect 8308 2322 8342 2356
rect 8380 2322 8414 2356
rect 8452 2322 8486 2356
rect 8524 2322 8558 2356
rect 8596 2322 8630 2356
rect 8668 2322 8702 2356
rect 8740 2322 8774 2356
rect 8812 2322 8846 2356
rect 8884 2322 8918 2356
rect 8956 2322 8990 2356
rect 9028 2322 9062 2356
rect 9100 2322 9134 2356
rect 9172 2322 9206 2356
rect 9244 2322 9278 2356
rect 7876 2277 7910 2283
rect 7876 2249 7880 2277
rect 7880 2249 7910 2277
rect 7948 2249 7982 2283
rect 8020 2277 8054 2283
rect 8020 2249 8050 2277
rect 8050 2249 8054 2277
rect 8092 2249 8126 2283
rect 8164 2277 8198 2283
rect 8164 2249 8186 2277
rect 8186 2249 8198 2277
rect 8236 2249 8270 2283
rect 8308 2277 8342 2283
rect 8308 2249 8322 2277
rect 8322 2249 8342 2277
rect 8380 2249 8414 2283
rect 8452 2277 8486 2283
rect 8452 2249 8458 2277
rect 8458 2249 8486 2277
rect 8524 2249 8558 2283
rect 8596 2249 8630 2283
rect 8668 2277 8702 2283
rect 8668 2249 8696 2277
rect 8696 2249 8702 2277
rect 8740 2249 8774 2283
rect 8812 2277 8846 2283
rect 8812 2249 8832 2277
rect 8832 2249 8846 2277
rect 8884 2249 8918 2283
rect 8956 2277 8990 2283
rect 8956 2249 8968 2277
rect 8968 2249 8990 2277
rect 9028 2249 9062 2283
rect 9100 2277 9134 2283
rect 9100 2249 9104 2277
rect 9104 2249 9134 2277
rect 9172 2249 9206 2283
rect 9244 2277 9278 2283
rect 9244 2249 9274 2277
rect 9274 2249 9278 2277
rect 7876 2176 7910 2210
rect 7948 2176 7982 2210
rect 8020 2176 8054 2210
rect 8092 2176 8126 2210
rect 8164 2176 8198 2210
rect 8236 2176 8270 2210
rect 8308 2176 8342 2210
rect 8380 2176 8414 2210
rect 8452 2176 8486 2210
rect 8524 2176 8558 2210
rect 8596 2176 8630 2210
rect 8668 2176 8702 2210
rect 8740 2176 8774 2210
rect 8812 2176 8846 2210
rect 8884 2176 8918 2210
rect 8956 2176 8990 2210
rect 9028 2176 9062 2210
rect 9100 2176 9134 2210
rect 9172 2176 9206 2210
rect 9244 2176 9278 2210
rect 7876 2106 7880 2137
rect 7880 2106 7910 2137
rect 7876 2103 7910 2106
rect 7948 2103 7982 2137
rect 8020 2106 8050 2137
rect 8050 2106 8054 2137
rect 8020 2103 8054 2106
rect 8092 2103 8126 2137
rect 8164 2106 8186 2137
rect 8186 2106 8198 2137
rect 8164 2103 8198 2106
rect 8236 2103 8270 2137
rect 8308 2106 8322 2137
rect 8322 2106 8342 2137
rect 8308 2103 8342 2106
rect 8380 2103 8414 2137
rect 8452 2106 8458 2137
rect 8458 2106 8486 2137
rect 8452 2103 8486 2106
rect 8524 2103 8558 2137
rect 8596 2103 8630 2137
rect 8668 2106 8696 2137
rect 8696 2106 8702 2137
rect 8668 2103 8702 2106
rect 8740 2103 8774 2137
rect 8812 2106 8832 2137
rect 8832 2106 8846 2137
rect 8812 2103 8846 2106
rect 8884 2103 8918 2137
rect 8956 2106 8968 2137
rect 8968 2106 8990 2137
rect 8956 2103 8990 2106
rect 9028 2103 9062 2137
rect 9100 2106 9104 2137
rect 9104 2106 9134 2137
rect 9100 2103 9134 2106
rect 9172 2103 9206 2137
rect 9244 2106 9274 2137
rect 9274 2106 9278 2137
rect 9244 2103 9278 2106
rect 7876 2030 7910 2064
rect 7948 2030 7982 2064
rect 8020 2030 8054 2064
rect 8092 2030 8126 2064
rect 8164 2030 8198 2064
rect 8236 2030 8270 2064
rect 8308 2030 8342 2064
rect 8380 2030 8414 2064
rect 8452 2030 8486 2064
rect 8524 2030 8558 2064
rect 8596 2030 8630 2064
rect 8668 2030 8702 2064
rect 8740 2030 8774 2064
rect 8812 2030 8846 2064
rect 8884 2030 8918 2064
rect 8956 2030 8990 2064
rect 9028 2030 9062 2064
rect 9100 2030 9134 2064
rect 9172 2030 9206 2064
rect 9244 2030 9278 2064
rect 7876 1969 7880 1991
rect 7880 1969 7910 1991
rect 7876 1957 7910 1969
rect 7948 1957 7982 1991
rect 8020 1969 8050 1991
rect 8050 1969 8054 1991
rect 8020 1957 8054 1969
rect 8092 1957 8126 1991
rect 8164 1969 8186 1991
rect 8186 1969 8198 1991
rect 8164 1957 8198 1969
rect 8236 1957 8270 1991
rect 8308 1969 8322 1991
rect 8322 1969 8342 1991
rect 8308 1957 8342 1969
rect 8380 1957 8414 1991
rect 8452 1969 8458 1991
rect 8458 1969 8486 1991
rect 8452 1957 8486 1969
rect 8524 1957 8558 1991
rect 8596 1957 8630 1991
rect 8668 1969 8696 1991
rect 8696 1969 8702 1991
rect 8668 1957 8702 1969
rect 8740 1957 8774 1991
rect 8812 1969 8832 1991
rect 8832 1969 8846 1991
rect 8812 1957 8846 1969
rect 8884 1957 8918 1991
rect 8956 1969 8968 1991
rect 8968 1969 8990 1991
rect 8956 1957 8990 1969
rect 9028 1957 9062 1991
rect 9100 1969 9104 1991
rect 9104 1969 9134 1991
rect 9100 1957 9134 1969
rect 9172 1957 9206 1991
rect 9244 1969 9274 1991
rect 9274 1969 9278 1991
rect 9244 1957 9278 1969
rect 7876 1884 7910 1918
rect 7948 1884 7982 1918
rect 8020 1884 8054 1918
rect 8092 1884 8126 1918
rect 8164 1884 8198 1918
rect 8236 1884 8270 1918
rect 8308 1884 8342 1918
rect 8380 1884 8414 1918
rect 8452 1884 8486 1918
rect 8524 1884 8558 1918
rect 8596 1884 8630 1918
rect 8668 1884 8702 1918
rect 8740 1884 8774 1918
rect 8812 1884 8846 1918
rect 8884 1884 8918 1918
rect 8956 1884 8990 1918
rect 9028 1884 9062 1918
rect 9100 1884 9134 1918
rect 9172 1884 9206 1918
rect 9244 1884 9278 1918
rect 7876 1832 7880 1845
rect 7880 1832 7910 1845
rect 7876 1811 7910 1832
rect 7948 1811 7982 1845
rect 8020 1832 8050 1845
rect 8050 1832 8054 1845
rect 8020 1811 8054 1832
rect 8092 1811 8126 1845
rect 8164 1832 8186 1845
rect 8186 1832 8198 1845
rect 8164 1811 8198 1832
rect 8236 1811 8270 1845
rect 8308 1832 8322 1845
rect 8322 1832 8342 1845
rect 8308 1811 8342 1832
rect 8380 1811 8414 1845
rect 8452 1832 8458 1845
rect 8458 1832 8486 1845
rect 8452 1811 8486 1832
rect 8524 1811 8558 1845
rect 8596 1811 8630 1845
rect 8668 1832 8696 1845
rect 8696 1832 8702 1845
rect 8668 1811 8702 1832
rect 8740 1811 8774 1845
rect 8812 1832 8832 1845
rect 8832 1832 8846 1845
rect 8812 1811 8846 1832
rect 8884 1811 8918 1845
rect 8956 1832 8968 1845
rect 8968 1832 8990 1845
rect 8956 1811 8990 1832
rect 9028 1811 9062 1845
rect 9100 1832 9104 1845
rect 9104 1832 9134 1845
rect 9100 1811 9134 1832
rect 9172 1811 9206 1845
rect 9244 1832 9274 1845
rect 9274 1832 9278 1845
rect 9244 1811 9278 1832
rect 7876 1738 7910 1772
rect 7948 1738 7982 1772
rect 8020 1738 8054 1772
rect 8092 1738 8126 1772
rect 8164 1738 8198 1772
rect 8236 1738 8270 1772
rect 8308 1738 8342 1772
rect 8380 1738 8414 1772
rect 8452 1738 8486 1772
rect 8524 1738 8558 1772
rect 8596 1738 8630 1772
rect 8668 1738 8702 1772
rect 8740 1738 8774 1772
rect 8812 1738 8846 1772
rect 8884 1738 8918 1772
rect 8956 1738 8990 1772
rect 9028 1738 9062 1772
rect 9100 1738 9134 1772
rect 9172 1738 9206 1772
rect 9244 1738 9278 1772
rect 321 1592 355 1626
rect 393 1592 427 1626
rect 465 1592 499 1626
rect 537 1592 571 1626
rect 609 1592 643 1626
rect 681 1592 715 1626
rect 753 1592 787 1626
rect 825 1592 859 1626
rect 897 1592 931 1626
rect 969 1592 1003 1626
rect 321 1519 355 1553
rect 393 1519 427 1553
rect 465 1519 499 1553
rect 537 1519 571 1553
rect 609 1519 643 1553
rect 681 1519 715 1553
rect 753 1519 787 1553
rect 825 1519 859 1553
rect 897 1519 931 1553
rect 969 1519 1003 1553
rect 321 1455 355 1480
rect 321 1446 325 1455
rect 325 1446 355 1455
rect 393 1446 427 1480
rect 465 1455 499 1480
rect 465 1446 495 1455
rect 495 1446 499 1455
rect 537 1446 571 1480
rect 609 1455 643 1480
rect 609 1446 631 1455
rect 631 1446 643 1455
rect 681 1446 715 1480
rect 753 1455 787 1480
rect 753 1446 767 1455
rect 767 1446 787 1455
rect 825 1446 859 1480
rect 897 1455 931 1480
rect 897 1446 903 1455
rect 903 1446 931 1455
rect 969 1446 1003 1480
rect 321 1373 355 1407
rect 393 1373 427 1407
rect 465 1373 499 1407
rect 537 1373 571 1407
rect 609 1373 643 1407
rect 681 1373 715 1407
rect 753 1373 787 1407
rect 825 1373 859 1407
rect 897 1373 931 1407
rect 969 1373 1003 1407
rect 321 1318 355 1334
rect 321 1300 325 1318
rect 325 1300 355 1318
rect 393 1300 427 1334
rect 465 1318 499 1334
rect 465 1300 495 1318
rect 495 1300 499 1318
rect 537 1300 571 1334
rect 609 1318 643 1334
rect 609 1300 631 1318
rect 631 1300 643 1318
rect 681 1300 715 1334
rect 753 1318 787 1334
rect 753 1300 767 1318
rect 767 1300 787 1318
rect 825 1300 859 1334
rect 897 1318 931 1334
rect 897 1300 903 1318
rect 903 1300 931 1318
rect 969 1300 1003 1334
rect 321 1227 355 1261
rect 393 1227 427 1261
rect 465 1227 499 1261
rect 537 1227 571 1261
rect 609 1227 643 1261
rect 681 1227 715 1261
rect 753 1227 787 1261
rect 825 1227 859 1261
rect 897 1227 931 1261
rect 969 1227 1003 1261
rect 321 1181 355 1188
rect 321 1154 325 1181
rect 325 1154 355 1181
rect 393 1154 427 1188
rect 465 1181 499 1188
rect 465 1154 495 1181
rect 495 1154 499 1181
rect 537 1154 571 1188
rect 609 1181 643 1188
rect 609 1154 631 1181
rect 631 1154 643 1181
rect 681 1154 715 1188
rect 753 1181 787 1188
rect 753 1154 767 1181
rect 767 1154 787 1181
rect 825 1154 859 1188
rect 897 1181 931 1188
rect 897 1154 903 1181
rect 903 1154 931 1181
rect 969 1154 1003 1188
rect 321 1081 355 1115
rect 393 1081 427 1115
rect 465 1081 499 1115
rect 537 1081 571 1115
rect 609 1081 643 1115
rect 681 1081 715 1115
rect 753 1081 787 1115
rect 825 1081 859 1115
rect 897 1081 931 1115
rect 969 1081 1003 1115
rect 321 1010 325 1042
rect 325 1010 355 1042
rect 321 1008 355 1010
rect 393 1008 427 1042
rect 465 1010 495 1042
rect 495 1010 499 1042
rect 465 1008 499 1010
rect 537 1008 571 1042
rect 609 1010 631 1042
rect 631 1010 643 1042
rect 609 1008 643 1010
rect 681 1008 715 1042
rect 753 1010 767 1042
rect 767 1010 787 1042
rect 753 1008 787 1010
rect 825 1008 859 1042
rect 897 1010 903 1042
rect 903 1010 931 1042
rect 897 1008 931 1010
rect 969 1008 1003 1042
rect 321 935 355 969
rect 393 935 427 969
rect 465 935 499 969
rect 537 935 571 969
rect 609 935 643 969
rect 681 935 715 969
rect 753 935 787 969
rect 825 935 859 969
rect 897 935 931 969
rect 969 935 1003 969
rect 321 873 325 896
rect 325 873 355 896
rect 321 862 355 873
rect 393 862 427 896
rect 465 873 495 896
rect 495 873 499 896
rect 465 862 499 873
rect 537 862 571 896
rect 609 873 631 896
rect 631 873 643 896
rect 609 862 643 873
rect 681 862 715 896
rect 753 873 767 896
rect 767 873 787 896
rect 753 862 787 873
rect 825 862 859 896
rect 897 873 903 896
rect 903 873 931 896
rect 897 862 931 873
rect 969 862 1003 896
rect 321 789 355 823
rect 393 789 427 823
rect 465 789 499 823
rect 537 789 571 823
rect 609 789 643 823
rect 681 789 715 823
rect 753 789 787 823
rect 825 789 859 823
rect 897 789 931 823
rect 969 789 1003 823
rect 321 736 325 750
rect 325 736 355 750
rect 321 716 355 736
rect 393 716 427 750
rect 465 736 495 750
rect 495 736 499 750
rect 465 716 499 736
rect 537 716 571 750
rect 609 736 631 750
rect 631 736 643 750
rect 609 716 643 736
rect 681 716 715 750
rect 753 736 767 750
rect 767 736 787 750
rect 753 716 787 736
rect 825 716 859 750
rect 897 736 903 750
rect 903 736 931 750
rect 897 716 931 736
rect 969 716 1003 750
rect 321 643 355 677
rect 393 643 427 677
rect 465 643 499 677
rect 537 643 571 677
rect 609 643 643 677
rect 681 643 715 677
rect 753 643 787 677
rect 825 643 859 677
rect 897 643 931 677
rect 969 643 1003 677
rect 321 599 325 604
rect 325 599 355 604
rect 321 570 355 599
rect 393 570 427 604
rect 465 599 495 604
rect 495 599 499 604
rect 465 570 499 599
rect 537 570 571 604
rect 609 599 631 604
rect 631 599 643 604
rect 609 570 643 599
rect 681 570 715 604
rect 753 599 767 604
rect 767 599 787 604
rect 753 570 787 599
rect 825 570 859 604
rect 897 599 903 604
rect 903 599 931 604
rect 897 570 931 599
rect 969 570 1003 604
rect 321 497 355 531
rect 393 497 427 531
rect 465 497 499 531
rect 537 497 571 531
rect 609 497 643 531
rect 681 497 715 531
rect 753 497 787 531
rect 825 497 859 531
rect 897 497 931 531
rect 969 497 1003 531
rect 321 424 355 458
rect 393 424 427 458
rect 465 424 499 458
rect 537 424 571 458
rect 609 424 643 458
rect 681 424 715 458
rect 753 424 787 458
rect 825 424 859 458
rect 897 424 931 458
rect 969 424 1003 458
rect 321 359 355 385
rect 321 351 325 359
rect 325 351 355 359
rect 393 351 427 385
rect 465 359 499 385
rect 465 351 495 359
rect 495 351 499 359
rect 537 351 571 385
rect 609 359 643 385
rect 609 351 631 359
rect 631 351 643 359
rect 681 351 715 385
rect 753 359 787 385
rect 753 351 767 359
rect 767 351 787 359
rect 825 351 859 385
rect 897 359 931 385
rect 897 351 903 359
rect 903 351 931 359
rect 969 351 1003 385
rect 321 278 355 312
rect 393 278 427 312
rect 465 278 499 312
rect 537 278 571 312
rect 609 278 643 312
rect 681 278 715 312
rect 753 278 787 312
rect 825 278 859 312
rect 897 278 931 312
rect 969 278 1003 312
rect 321 222 355 239
rect 321 205 325 222
rect 325 205 355 222
rect 393 205 427 239
rect 465 222 499 239
rect 465 205 495 222
rect 495 205 499 222
rect 537 205 571 239
rect 609 222 643 239
rect 609 205 631 222
rect 631 205 643 222
rect 681 205 715 239
rect 753 222 787 239
rect 753 205 767 222
rect 767 205 787 222
rect 825 205 859 239
rect 897 222 931 239
rect 897 205 903 222
rect 903 205 931 222
rect 969 205 1003 239
rect 321 132 355 166
rect 393 132 427 166
rect 465 132 499 166
rect 537 132 571 166
rect 609 132 643 166
rect 681 132 715 166
rect 753 132 787 166
rect 825 132 859 166
rect 897 132 931 166
rect 969 132 1003 166
rect 321 85 355 93
rect 321 59 325 85
rect 325 59 355 85
rect 393 59 427 93
rect 465 85 499 93
rect 465 59 495 85
rect 495 59 499 85
rect 537 59 571 93
rect 609 85 643 93
rect 609 59 631 85
rect 631 59 643 85
rect 681 59 715 93
rect 753 85 787 93
rect 753 59 767 85
rect 767 59 787 85
rect 825 59 859 93
rect 897 85 931 93
rect 897 59 903 85
rect 903 59 931 85
rect 969 59 1003 93
rect 7876 1695 7880 1699
rect 7880 1695 7910 1699
rect 7876 1665 7910 1695
rect 7948 1665 7982 1699
rect 8020 1695 8050 1699
rect 8050 1695 8054 1699
rect 8020 1665 8054 1695
rect 8092 1665 8126 1699
rect 8164 1695 8186 1699
rect 8186 1695 8198 1699
rect 8164 1665 8198 1695
rect 8236 1665 8270 1699
rect 8308 1695 8322 1699
rect 8322 1695 8342 1699
rect 8308 1665 8342 1695
rect 8380 1665 8414 1699
rect 8452 1695 8458 1699
rect 8458 1695 8486 1699
rect 8452 1665 8486 1695
rect 8524 1665 8558 1699
rect 8596 1665 8630 1699
rect 8668 1695 8696 1699
rect 8696 1695 8702 1699
rect 8668 1665 8702 1695
rect 8740 1665 8774 1699
rect 8812 1695 8832 1699
rect 8832 1695 8846 1699
rect 8812 1665 8846 1695
rect 8884 1665 8918 1699
rect 8956 1695 8968 1699
rect 8968 1695 8990 1699
rect 8956 1665 8990 1695
rect 9028 1665 9062 1699
rect 9100 1695 9104 1699
rect 9104 1695 9134 1699
rect 9100 1665 9134 1695
rect 9172 1665 9206 1699
rect 9244 1695 9274 1699
rect 9274 1695 9278 1699
rect 9244 1665 9278 1695
rect 7876 1592 7910 1626
rect 7948 1592 7982 1626
rect 8020 1592 8054 1626
rect 8092 1592 8126 1626
rect 8164 1592 8198 1626
rect 8236 1592 8270 1626
rect 8308 1592 8342 1626
rect 8380 1592 8414 1626
rect 8452 1592 8486 1626
rect 8524 1592 8558 1626
rect 8596 1592 8630 1626
rect 8668 1592 8702 1626
rect 8740 1592 8774 1626
rect 8812 1592 8846 1626
rect 8884 1592 8918 1626
rect 8956 1592 8990 1626
rect 9028 1592 9062 1626
rect 9100 1592 9134 1626
rect 9172 1592 9206 1626
rect 9244 1592 9278 1626
rect 7876 1519 7910 1553
rect 7948 1519 7982 1553
rect 8020 1519 8054 1553
rect 8092 1519 8126 1553
rect 8164 1519 8198 1553
rect 8236 1519 8270 1553
rect 8308 1519 8342 1553
rect 8380 1519 8414 1553
rect 8452 1519 8486 1553
rect 8524 1519 8558 1553
rect 8596 1519 8630 1553
rect 8668 1519 8702 1553
rect 8740 1519 8774 1553
rect 8812 1519 8846 1553
rect 8884 1519 8918 1553
rect 8956 1519 8990 1553
rect 9028 1519 9062 1553
rect 9100 1519 9134 1553
rect 9172 1519 9206 1553
rect 9244 1519 9278 1553
rect 7876 1455 7910 1480
rect 7876 1446 7880 1455
rect 7880 1446 7910 1455
rect 7948 1446 7982 1480
rect 8020 1455 8054 1480
rect 8020 1446 8050 1455
rect 8050 1446 8054 1455
rect 8092 1446 8126 1480
rect 8164 1455 8198 1480
rect 8164 1446 8186 1455
rect 8186 1446 8198 1455
rect 8236 1446 8270 1480
rect 8308 1455 8342 1480
rect 8308 1446 8322 1455
rect 8322 1446 8342 1455
rect 8380 1446 8414 1480
rect 8452 1455 8486 1480
rect 8452 1446 8458 1455
rect 8458 1446 8486 1455
rect 8524 1446 8558 1480
rect 8596 1446 8630 1480
rect 8668 1455 8702 1480
rect 8668 1446 8696 1455
rect 8696 1446 8702 1455
rect 8740 1446 8774 1480
rect 8812 1455 8846 1480
rect 8812 1446 8832 1455
rect 8832 1446 8846 1455
rect 8884 1446 8918 1480
rect 8956 1455 8990 1480
rect 8956 1446 8968 1455
rect 8968 1446 8990 1455
rect 9028 1446 9062 1480
rect 9100 1455 9134 1480
rect 9100 1446 9104 1455
rect 9104 1446 9134 1455
rect 9172 1446 9206 1480
rect 9244 1455 9278 1480
rect 9244 1446 9274 1455
rect 9274 1446 9278 1455
rect 7876 1373 7910 1407
rect 7948 1373 7982 1407
rect 8020 1373 8054 1407
rect 8092 1373 8126 1407
rect 8164 1373 8198 1407
rect 8236 1373 8270 1407
rect 8308 1373 8342 1407
rect 8380 1373 8414 1407
rect 8452 1373 8486 1407
rect 8524 1373 8558 1407
rect 8596 1373 8630 1407
rect 8668 1373 8702 1407
rect 8740 1373 8774 1407
rect 8812 1373 8846 1407
rect 8884 1373 8918 1407
rect 8956 1373 8990 1407
rect 9028 1373 9062 1407
rect 9100 1373 9134 1407
rect 9172 1373 9206 1407
rect 9244 1373 9278 1407
rect 7876 1318 7910 1334
rect 7876 1300 7880 1318
rect 7880 1300 7910 1318
rect 7948 1300 7982 1334
rect 8020 1318 8054 1334
rect 8020 1300 8050 1318
rect 8050 1300 8054 1318
rect 8092 1300 8126 1334
rect 8164 1318 8198 1334
rect 8164 1300 8186 1318
rect 8186 1300 8198 1318
rect 8236 1300 8270 1334
rect 8308 1318 8342 1334
rect 8308 1300 8322 1318
rect 8322 1300 8342 1318
rect 8380 1300 8414 1334
rect 8452 1318 8486 1334
rect 8452 1300 8458 1318
rect 8458 1300 8486 1318
rect 8524 1300 8558 1334
rect 8596 1300 8630 1334
rect 8668 1318 8702 1334
rect 8668 1300 8696 1318
rect 8696 1300 8702 1318
rect 8740 1300 8774 1334
rect 8812 1318 8846 1334
rect 8812 1300 8832 1318
rect 8832 1300 8846 1318
rect 8884 1300 8918 1334
rect 8956 1318 8990 1334
rect 8956 1300 8968 1318
rect 8968 1300 8990 1318
rect 9028 1300 9062 1334
rect 9100 1318 9134 1334
rect 9100 1300 9104 1318
rect 9104 1300 9134 1318
rect 9172 1300 9206 1334
rect 9244 1318 9278 1334
rect 9244 1300 9274 1318
rect 9274 1300 9278 1318
rect 7876 1227 7910 1261
rect 7948 1227 7982 1261
rect 8020 1227 8054 1261
rect 8092 1227 8126 1261
rect 8164 1227 8198 1261
rect 8236 1227 8270 1261
rect 8308 1227 8342 1261
rect 8380 1227 8414 1261
rect 8452 1227 8486 1261
rect 8524 1227 8558 1261
rect 8596 1227 8630 1261
rect 8668 1227 8702 1261
rect 8740 1227 8774 1261
rect 8812 1227 8846 1261
rect 8884 1227 8918 1261
rect 8956 1227 8990 1261
rect 9028 1227 9062 1261
rect 9100 1227 9134 1261
rect 9172 1227 9206 1261
rect 9244 1227 9278 1261
rect 7876 1181 7910 1188
rect 7876 1154 7880 1181
rect 7880 1154 7910 1181
rect 7948 1154 7982 1188
rect 8020 1181 8054 1188
rect 8020 1154 8050 1181
rect 8050 1154 8054 1181
rect 8092 1154 8126 1188
rect 8164 1181 8198 1188
rect 8164 1154 8186 1181
rect 8186 1154 8198 1181
rect 8236 1154 8270 1188
rect 8308 1181 8342 1188
rect 8308 1154 8322 1181
rect 8322 1154 8342 1181
rect 8380 1154 8414 1188
rect 8452 1181 8486 1188
rect 8452 1154 8458 1181
rect 8458 1154 8486 1181
rect 8524 1154 8558 1188
rect 8596 1154 8630 1188
rect 8668 1181 8702 1188
rect 8668 1154 8696 1181
rect 8696 1154 8702 1181
rect 8740 1154 8774 1188
rect 8812 1181 8846 1188
rect 8812 1154 8832 1181
rect 8832 1154 8846 1181
rect 8884 1154 8918 1188
rect 8956 1181 8990 1188
rect 8956 1154 8968 1181
rect 8968 1154 8990 1181
rect 9028 1154 9062 1188
rect 9100 1181 9134 1188
rect 9100 1154 9104 1181
rect 9104 1154 9134 1181
rect 9172 1154 9206 1188
rect 9244 1181 9278 1188
rect 9244 1154 9274 1181
rect 9274 1154 9278 1181
rect 7876 1081 7910 1115
rect 7948 1081 7982 1115
rect 8020 1081 8054 1115
rect 8092 1081 8126 1115
rect 8164 1081 8198 1115
rect 8236 1081 8270 1115
rect 8308 1081 8342 1115
rect 8380 1081 8414 1115
rect 8452 1081 8486 1115
rect 8524 1081 8558 1115
rect 8596 1081 8630 1115
rect 8668 1081 8702 1115
rect 8740 1081 8774 1115
rect 8812 1081 8846 1115
rect 8884 1081 8918 1115
rect 8956 1081 8990 1115
rect 9028 1081 9062 1115
rect 9100 1081 9134 1115
rect 9172 1081 9206 1115
rect 9244 1081 9278 1115
rect 7876 1010 7880 1042
rect 7880 1010 7910 1042
rect 7876 1008 7910 1010
rect 7948 1008 7982 1042
rect 8020 1010 8050 1042
rect 8050 1010 8054 1042
rect 8020 1008 8054 1010
rect 8092 1008 8126 1042
rect 8164 1010 8186 1042
rect 8186 1010 8198 1042
rect 8164 1008 8198 1010
rect 8236 1008 8270 1042
rect 8308 1010 8322 1042
rect 8322 1010 8342 1042
rect 8308 1008 8342 1010
rect 8380 1008 8414 1042
rect 8452 1010 8458 1042
rect 8458 1010 8486 1042
rect 8452 1008 8486 1010
rect 8524 1008 8558 1042
rect 8596 1008 8630 1042
rect 8668 1010 8696 1042
rect 8696 1010 8702 1042
rect 8668 1008 8702 1010
rect 8740 1008 8774 1042
rect 8812 1010 8832 1042
rect 8832 1010 8846 1042
rect 8812 1008 8846 1010
rect 8884 1008 8918 1042
rect 8956 1010 8968 1042
rect 8968 1010 8990 1042
rect 8956 1008 8990 1010
rect 9028 1008 9062 1042
rect 9100 1010 9104 1042
rect 9104 1010 9134 1042
rect 9100 1008 9134 1010
rect 9172 1008 9206 1042
rect 9244 1010 9274 1042
rect 9274 1010 9278 1042
rect 9244 1008 9278 1010
rect 7876 935 7910 969
rect 7948 935 7982 969
rect 8020 935 8054 969
rect 8092 935 8126 969
rect 8164 935 8198 969
rect 8236 935 8270 969
rect 8308 935 8342 969
rect 8380 935 8414 969
rect 8452 935 8486 969
rect 8524 935 8558 969
rect 8596 935 8630 969
rect 8668 935 8702 969
rect 8740 935 8774 969
rect 8812 935 8846 969
rect 8884 935 8918 969
rect 8956 935 8990 969
rect 9028 935 9062 969
rect 9100 935 9134 969
rect 9172 935 9206 969
rect 9244 935 9278 969
rect 7876 873 7880 896
rect 7880 873 7910 896
rect 7876 862 7910 873
rect 7948 862 7982 896
rect 8020 873 8050 896
rect 8050 873 8054 896
rect 8020 862 8054 873
rect 8092 862 8126 896
rect 8164 873 8186 896
rect 8186 873 8198 896
rect 8164 862 8198 873
rect 8236 862 8270 896
rect 8308 873 8322 896
rect 8322 873 8342 896
rect 8308 862 8342 873
rect 8380 862 8414 896
rect 8452 873 8458 896
rect 8458 873 8486 896
rect 8452 862 8486 873
rect 8524 862 8558 896
rect 8596 862 8630 896
rect 8668 873 8696 896
rect 8696 873 8702 896
rect 8668 862 8702 873
rect 8740 862 8774 896
rect 8812 873 8832 896
rect 8832 873 8846 896
rect 8812 862 8846 873
rect 8884 862 8918 896
rect 8956 873 8968 896
rect 8968 873 8990 896
rect 8956 862 8990 873
rect 9028 862 9062 896
rect 9100 873 9104 896
rect 9104 873 9134 896
rect 9100 862 9134 873
rect 9172 862 9206 896
rect 9244 873 9274 896
rect 9274 873 9278 896
rect 9244 862 9278 873
rect 7876 789 7910 823
rect 7948 789 7982 823
rect 8020 789 8054 823
rect 8092 789 8126 823
rect 8164 789 8198 823
rect 8236 789 8270 823
rect 8308 789 8342 823
rect 8380 789 8414 823
rect 8452 789 8486 823
rect 8524 789 8558 823
rect 8596 789 8630 823
rect 8668 789 8702 823
rect 8740 789 8774 823
rect 8812 789 8846 823
rect 8884 789 8918 823
rect 8956 789 8990 823
rect 9028 789 9062 823
rect 9100 789 9134 823
rect 9172 789 9206 823
rect 9244 789 9278 823
rect 7876 736 7880 750
rect 7880 736 7910 750
rect 7876 716 7910 736
rect 7948 716 7982 750
rect 8020 736 8050 750
rect 8050 736 8054 750
rect 8020 716 8054 736
rect 8092 716 8126 750
rect 8164 736 8186 750
rect 8186 736 8198 750
rect 8164 716 8198 736
rect 8236 716 8270 750
rect 8308 736 8322 750
rect 8322 736 8342 750
rect 8308 716 8342 736
rect 8380 716 8414 750
rect 8452 736 8458 750
rect 8458 736 8486 750
rect 8452 716 8486 736
rect 8524 716 8558 750
rect 8596 716 8630 750
rect 8668 736 8696 750
rect 8696 736 8702 750
rect 8668 716 8702 736
rect 8740 716 8774 750
rect 8812 736 8832 750
rect 8832 736 8846 750
rect 8812 716 8846 736
rect 8884 716 8918 750
rect 8956 736 8968 750
rect 8968 736 8990 750
rect 8956 716 8990 736
rect 9028 716 9062 750
rect 9100 736 9104 750
rect 9104 736 9134 750
rect 9100 716 9134 736
rect 9172 716 9206 750
rect 9244 736 9274 750
rect 9274 736 9278 750
rect 9244 716 9278 736
rect 7876 643 7910 677
rect 7948 643 7982 677
rect 8020 643 8054 677
rect 8092 643 8126 677
rect 8164 643 8198 677
rect 8236 643 8270 677
rect 8308 643 8342 677
rect 8380 643 8414 677
rect 8452 643 8486 677
rect 8524 643 8558 677
rect 8596 643 8630 677
rect 8668 643 8702 677
rect 8740 643 8774 677
rect 8812 643 8846 677
rect 8884 643 8918 677
rect 8956 643 8990 677
rect 9028 643 9062 677
rect 9100 643 9134 677
rect 9172 643 9206 677
rect 9244 643 9278 677
rect 7876 599 7880 604
rect 7880 599 7910 604
rect 7876 570 7910 599
rect 7948 570 7982 604
rect 8020 599 8050 604
rect 8050 599 8054 604
rect 8020 570 8054 599
rect 8092 570 8126 604
rect 8164 599 8186 604
rect 8186 599 8198 604
rect 8164 570 8198 599
rect 8236 570 8270 604
rect 8308 599 8322 604
rect 8322 599 8342 604
rect 8308 570 8342 599
rect 8380 570 8414 604
rect 8452 599 8458 604
rect 8458 599 8486 604
rect 8452 570 8486 599
rect 8524 570 8558 604
rect 8596 570 8630 604
rect 8668 599 8696 604
rect 8696 599 8702 604
rect 8668 570 8702 599
rect 8740 570 8774 604
rect 8812 599 8832 604
rect 8832 599 8846 604
rect 8812 570 8846 599
rect 8884 570 8918 604
rect 8956 599 8968 604
rect 8968 599 8990 604
rect 8956 570 8990 599
rect 9028 570 9062 604
rect 9100 599 9104 604
rect 9104 599 9134 604
rect 9100 570 9134 599
rect 9172 570 9206 604
rect 9244 599 9274 604
rect 9274 599 9278 604
rect 9244 570 9278 599
rect 7876 497 7910 531
rect 7948 497 7982 531
rect 8020 497 8054 531
rect 8092 497 8126 531
rect 8164 497 8198 531
rect 8236 497 8270 531
rect 8308 497 8342 531
rect 8380 497 8414 531
rect 8452 497 8486 531
rect 8524 497 8558 531
rect 8596 497 8630 531
rect 8668 497 8702 531
rect 8740 497 8774 531
rect 8812 497 8846 531
rect 8884 497 8918 531
rect 8956 497 8990 531
rect 9028 497 9062 531
rect 9100 497 9134 531
rect 9172 497 9206 531
rect 9244 497 9278 531
rect 7876 424 7910 458
rect 7948 424 7982 458
rect 8020 424 8054 458
rect 8092 424 8126 458
rect 8164 424 8198 458
rect 8236 424 8270 458
rect 8308 424 8342 458
rect 8380 424 8414 458
rect 8452 424 8486 458
rect 8524 424 8558 458
rect 8596 424 8630 458
rect 8668 424 8702 458
rect 8740 424 8774 458
rect 8812 424 8846 458
rect 8884 424 8918 458
rect 8956 424 8990 458
rect 9028 424 9062 458
rect 9100 424 9134 458
rect 9172 424 9206 458
rect 9244 424 9278 458
rect 7876 359 7910 385
rect 7876 351 7880 359
rect 7880 351 7910 359
rect 7948 351 7982 385
rect 8020 359 8054 385
rect 8020 351 8050 359
rect 8050 351 8054 359
rect 8092 351 8126 385
rect 8164 359 8198 385
rect 8164 351 8186 359
rect 8186 351 8198 359
rect 8236 351 8270 385
rect 8308 359 8342 385
rect 8308 351 8322 359
rect 8322 351 8342 359
rect 8380 351 8414 385
rect 8452 359 8486 385
rect 8452 351 8458 359
rect 8458 351 8486 359
rect 8524 351 8558 385
rect 8596 351 8630 385
rect 8668 359 8702 385
rect 8668 351 8696 359
rect 8696 351 8702 359
rect 8740 351 8774 385
rect 8812 359 8846 385
rect 8812 351 8832 359
rect 8832 351 8846 359
rect 8884 351 8918 385
rect 8956 359 8990 385
rect 8956 351 8968 359
rect 8968 351 8990 359
rect 9028 351 9062 385
rect 9100 359 9134 385
rect 9100 351 9104 359
rect 9104 351 9134 359
rect 9172 351 9206 385
rect 9244 359 9278 385
rect 9244 351 9274 359
rect 9274 351 9278 359
rect 7876 278 7910 312
rect 7948 278 7982 312
rect 8020 278 8054 312
rect 8092 278 8126 312
rect 8164 278 8198 312
rect 8236 278 8270 312
rect 8308 278 8342 312
rect 8380 278 8414 312
rect 8452 278 8486 312
rect 8524 278 8558 312
rect 8596 278 8630 312
rect 8668 278 8702 312
rect 8740 278 8774 312
rect 8812 278 8846 312
rect 8884 278 8918 312
rect 8956 278 8990 312
rect 9028 278 9062 312
rect 9100 278 9134 312
rect 9172 278 9206 312
rect 9244 278 9278 312
rect 7876 222 7910 239
rect 7876 205 7880 222
rect 7880 205 7910 222
rect 7948 205 7982 239
rect 8020 222 8054 239
rect 8020 205 8050 222
rect 8050 205 8054 222
rect 8092 205 8126 239
rect 8164 222 8198 239
rect 8164 205 8186 222
rect 8186 205 8198 222
rect 8236 205 8270 239
rect 8308 222 8342 239
rect 8308 205 8322 222
rect 8322 205 8342 222
rect 8380 205 8414 239
rect 8452 222 8486 239
rect 8452 205 8458 222
rect 8458 205 8486 222
rect 8524 205 8558 239
rect 8596 205 8630 239
rect 8668 222 8702 239
rect 8668 205 8696 222
rect 8696 205 8702 222
rect 8740 205 8774 239
rect 8812 222 8846 239
rect 8812 205 8832 222
rect 8832 205 8846 222
rect 8884 205 8918 239
rect 8956 222 8990 239
rect 8956 205 8968 222
rect 8968 205 8990 222
rect 9028 205 9062 239
rect 9100 222 9134 239
rect 9100 205 9104 222
rect 9104 205 9134 222
rect 9172 205 9206 239
rect 9244 222 9278 239
rect 9244 205 9274 222
rect 9274 205 9278 222
rect 7876 132 7910 166
rect 7948 132 7982 166
rect 8020 132 8054 166
rect 8092 132 8126 166
rect 8164 132 8198 166
rect 8236 132 8270 166
rect 8308 132 8342 166
rect 8380 132 8414 166
rect 8452 132 8486 166
rect 8524 132 8558 166
rect 8596 132 8630 166
rect 8668 132 8702 166
rect 8740 132 8774 166
rect 8812 132 8846 166
rect 8884 132 8918 166
rect 8956 132 8990 166
rect 9028 132 9062 166
rect 9100 132 9134 166
rect 9172 132 9206 166
rect 9244 132 9278 166
rect 7876 85 7910 93
rect 7876 59 7880 85
rect 7880 59 7910 85
rect 7948 59 7982 93
rect 8020 85 8054 93
rect 8020 59 8050 85
rect 8050 59 8054 85
rect 8092 59 8126 93
rect 8164 85 8198 93
rect 8164 59 8186 85
rect 8186 59 8198 85
rect 8236 59 8270 93
rect 8308 85 8342 93
rect 8308 59 8322 85
rect 8322 59 8342 85
rect 8380 59 8414 93
rect 8452 85 8486 93
rect 8452 59 8458 85
rect 8458 59 8486 85
rect 8524 59 8558 93
rect 8596 59 8630 93
rect 8668 85 8702 93
rect 8668 59 8696 85
rect 8696 59 8702 85
rect 8740 59 8774 93
rect 8812 85 8846 93
rect 8812 59 8832 85
rect 8832 59 8846 85
rect 8884 59 8918 93
rect 8956 85 8990 93
rect 8956 59 8968 85
rect 8968 59 8990 85
rect 9028 59 9062 93
rect 9100 85 9134 93
rect 9100 59 9104 85
rect 9104 59 9134 85
rect 9172 59 9206 93
rect 9244 85 9278 93
rect 9244 59 9274 85
rect 9274 59 9278 85
<< metal1 >>
rect 315 39943 1729 39975
rect 315 33357 321 39943
rect 1723 33357 1729 39943
rect 315 33318 1729 33357
rect 315 33284 321 33318
rect 355 33284 393 33318
rect 427 33284 465 33318
rect 499 33284 537 33318
rect 571 33284 609 33318
rect 643 33284 681 33318
rect 715 33284 753 33318
rect 787 33284 825 33318
rect 859 33284 897 33318
rect 931 33284 969 33318
rect 1003 33284 1041 33318
rect 1075 33284 1113 33318
rect 1147 33284 1185 33318
rect 1219 33284 1257 33318
rect 1291 33284 1329 33318
rect 1363 33284 1401 33318
rect 1435 33284 1473 33318
rect 1507 33284 1545 33318
rect 1579 33284 1617 33318
rect 1651 33284 1689 33318
rect 1723 33284 1729 33318
rect 315 33245 1729 33284
rect 315 33211 321 33245
rect 355 33211 393 33245
rect 427 33211 465 33245
rect 499 33211 537 33245
rect 571 33211 609 33245
rect 643 33211 681 33245
rect 715 33211 753 33245
rect 787 33211 825 33245
rect 859 33211 897 33245
rect 931 33211 969 33245
rect 1003 33211 1041 33245
rect 1075 33211 1113 33245
rect 1147 33211 1185 33245
rect 1219 33211 1257 33245
rect 1291 33211 1329 33245
rect 1363 33211 1401 33245
rect 1435 33211 1473 33245
rect 1507 33211 1545 33245
rect 1579 33211 1617 33245
rect 1651 33211 1689 33245
rect 1723 33211 1729 33245
rect 315 33172 1729 33211
rect 315 33138 321 33172
rect 355 33138 393 33172
rect 427 33138 465 33172
rect 499 33138 537 33172
rect 571 33138 609 33172
rect 643 33138 681 33172
rect 715 33138 753 33172
rect 787 33138 825 33172
rect 859 33138 897 33172
rect 931 33138 969 33172
rect 1003 33138 1041 33172
rect 1075 33138 1113 33172
rect 1147 33138 1185 33172
rect 1219 33138 1257 33172
rect 1291 33138 1329 33172
rect 1363 33138 1401 33172
rect 1435 33138 1473 33172
rect 1507 33138 1545 33172
rect 1579 33138 1617 33172
rect 1651 33138 1689 33172
rect 1723 33138 1729 33172
rect 315 33099 1729 33138
rect 315 33065 321 33099
rect 355 33065 393 33099
rect 427 33065 465 33099
rect 499 33065 537 33099
rect 571 33065 609 33099
rect 643 33065 681 33099
rect 715 33065 753 33099
rect 787 33065 825 33099
rect 859 33065 897 33099
rect 931 33065 969 33099
rect 1003 33065 1041 33099
rect 1075 33065 1113 33099
rect 1147 33065 1185 33099
rect 1219 33065 1257 33099
rect 1291 33065 1329 33099
rect 1363 33065 1401 33099
rect 1435 33065 1473 33099
rect 1507 33065 1545 33099
rect 1579 33065 1617 33099
rect 1651 33065 1689 33099
rect 1723 33065 1729 33099
rect 315 33026 1729 33065
rect 315 32992 321 33026
rect 355 32992 393 33026
rect 427 32992 465 33026
rect 499 32992 537 33026
rect 571 32992 609 33026
rect 643 32992 681 33026
rect 715 32992 753 33026
rect 787 32992 825 33026
rect 859 32992 897 33026
rect 931 32992 969 33026
rect 1003 32992 1041 33026
rect 1075 32992 1113 33026
rect 1147 32992 1185 33026
rect 1219 32992 1257 33026
rect 1291 32992 1329 33026
rect 1363 32992 1401 33026
rect 1435 32992 1473 33026
rect 1507 32992 1545 33026
rect 1579 32992 1617 33026
rect 1651 32992 1689 33026
rect 1723 32992 1729 33026
rect 315 32953 1729 32992
rect 315 32919 321 32953
rect 355 32919 393 32953
rect 427 32919 465 32953
rect 499 32919 537 32953
rect 571 32919 609 32953
rect 643 32919 681 32953
rect 715 32919 753 32953
rect 787 32919 825 32953
rect 859 32919 897 32953
rect 931 32919 969 32953
rect 1003 32919 1041 32953
rect 1075 32919 1113 32953
rect 1147 32919 1185 32953
rect 1219 32919 1257 32953
rect 1291 32919 1329 32953
rect 1363 32919 1401 32953
rect 1435 32919 1473 32953
rect 1507 32919 1545 32953
rect 1579 32919 1617 32953
rect 1651 32919 1689 32953
rect 1723 32919 1729 32953
rect 315 32880 1729 32919
rect 315 32846 321 32880
rect 355 32846 393 32880
rect 427 32846 465 32880
rect 499 32846 537 32880
rect 571 32846 609 32880
rect 643 32846 681 32880
rect 715 32846 753 32880
rect 787 32846 825 32880
rect 859 32846 897 32880
rect 931 32846 969 32880
rect 1003 32846 1041 32880
rect 1075 32846 1113 32880
rect 1147 32846 1185 32880
rect 1219 32846 1257 32880
rect 1291 32846 1329 32880
rect 1363 32846 1401 32880
rect 1435 32846 1473 32880
rect 1507 32846 1545 32880
rect 1579 32846 1617 32880
rect 1651 32846 1689 32880
rect 1723 32846 1729 32880
rect 315 32807 1729 32846
rect 315 32773 321 32807
rect 355 32773 393 32807
rect 427 32773 465 32807
rect 499 32773 537 32807
rect 571 32773 609 32807
rect 643 32773 681 32807
rect 715 32773 753 32807
rect 787 32773 825 32807
rect 859 32773 897 32807
rect 931 32773 969 32807
rect 1003 32773 1041 32807
rect 1075 32773 1113 32807
rect 1147 32773 1185 32807
rect 1219 32773 1257 32807
rect 1291 32773 1329 32807
rect 1363 32773 1401 32807
rect 1435 32773 1473 32807
rect 1507 32773 1545 32807
rect 1579 32773 1617 32807
rect 1651 32773 1689 32807
rect 1723 32773 1729 32807
rect 315 32734 1729 32773
rect 315 32700 321 32734
rect 355 32700 393 32734
rect 427 32700 465 32734
rect 499 32700 537 32734
rect 571 32700 609 32734
rect 643 32700 681 32734
rect 715 32700 753 32734
rect 787 32700 825 32734
rect 859 32700 897 32734
rect 931 32700 969 32734
rect 1003 32700 1041 32734
rect 1075 32700 1113 32734
rect 1147 32700 1185 32734
rect 1219 32700 1257 32734
rect 1291 32700 1329 32734
rect 1363 32700 1401 32734
rect 1435 32700 1473 32734
rect 1507 32700 1545 32734
rect 1579 32700 1617 32734
rect 1651 32700 1689 32734
rect 1723 32700 1729 32734
rect 315 32661 1729 32700
rect 315 32627 321 32661
rect 355 32627 393 32661
rect 427 32627 465 32661
rect 499 32627 537 32661
rect 571 32627 609 32661
rect 643 32627 681 32661
rect 715 32627 753 32661
rect 787 32627 825 32661
rect 859 32627 897 32661
rect 931 32627 969 32661
rect 1003 32627 1041 32661
rect 1075 32627 1113 32661
rect 1147 32627 1185 32661
rect 1219 32627 1257 32661
rect 1291 32627 1329 32661
rect 1363 32627 1401 32661
rect 1435 32627 1473 32661
rect 1507 32627 1545 32661
rect 1579 32627 1617 32661
rect 1651 32627 1689 32661
rect 1723 32627 1729 32661
rect 315 32588 1729 32627
rect 315 32554 321 32588
rect 355 32554 393 32588
rect 427 32554 465 32588
rect 499 32554 537 32588
rect 571 32554 609 32588
rect 643 32554 681 32588
rect 715 32554 753 32588
rect 787 32554 825 32588
rect 859 32554 897 32588
rect 931 32554 969 32588
rect 1003 32554 1041 32588
rect 1075 32554 1113 32588
rect 1147 32554 1185 32588
rect 1219 32554 1257 32588
rect 1291 32554 1329 32588
rect 1363 32554 1401 32588
rect 1435 32554 1473 32588
rect 1507 32554 1545 32588
rect 1579 32554 1617 32588
rect 1651 32554 1689 32588
rect 1723 32554 1729 32588
rect 315 32515 1729 32554
rect 315 32481 321 32515
rect 355 32481 393 32515
rect 427 32481 465 32515
rect 499 32481 537 32515
rect 571 32481 609 32515
rect 643 32481 681 32515
rect 715 32481 753 32515
rect 787 32481 825 32515
rect 859 32481 897 32515
rect 931 32481 969 32515
rect 1003 32481 1041 32515
rect 1075 32481 1113 32515
rect 1147 32481 1185 32515
rect 1219 32481 1257 32515
rect 1291 32481 1329 32515
rect 1363 32481 1401 32515
rect 1435 32481 1473 32515
rect 1507 32481 1545 32515
rect 1579 32481 1617 32515
rect 1651 32481 1689 32515
rect 1723 32481 1729 32515
rect 315 32442 1729 32481
rect 315 32408 321 32442
rect 355 32408 393 32442
rect 427 32408 465 32442
rect 499 32408 537 32442
rect 571 32408 609 32442
rect 643 32408 681 32442
rect 715 32408 753 32442
rect 787 32408 825 32442
rect 859 32408 897 32442
rect 931 32408 969 32442
rect 1003 32408 1041 32442
rect 1075 32408 1113 32442
rect 1147 32408 1185 32442
rect 1219 32408 1257 32442
rect 1291 32408 1329 32442
rect 1363 32408 1401 32442
rect 1435 32408 1473 32442
rect 1507 32408 1545 32442
rect 1579 32408 1617 32442
rect 1651 32408 1689 32442
rect 1723 32408 1729 32442
rect 315 32369 1729 32408
rect 315 32335 321 32369
rect 355 32335 393 32369
rect 427 32335 465 32369
rect 499 32335 537 32369
rect 571 32335 609 32369
rect 643 32335 681 32369
rect 715 32335 753 32369
rect 787 32335 825 32369
rect 859 32335 897 32369
rect 931 32335 969 32369
rect 1003 32335 1041 32369
rect 1075 32335 1113 32369
rect 1147 32335 1185 32369
rect 1219 32335 1257 32369
rect 1291 32335 1329 32369
rect 1363 32335 1401 32369
rect 1435 32335 1473 32369
rect 1507 32335 1545 32369
rect 1579 32335 1617 32369
rect 1651 32335 1689 32369
rect 1723 32335 1729 32369
rect 315 32296 1729 32335
rect 315 32262 321 32296
rect 355 32262 393 32296
rect 427 32262 465 32296
rect 499 32262 537 32296
rect 571 32262 609 32296
rect 643 32262 681 32296
rect 715 32262 753 32296
rect 787 32262 825 32296
rect 859 32262 897 32296
rect 931 32262 969 32296
rect 1003 32262 1041 32296
rect 1075 32262 1113 32296
rect 1147 32262 1185 32296
rect 1219 32262 1257 32296
rect 1291 32262 1329 32296
rect 1363 32262 1401 32296
rect 1435 32262 1473 32296
rect 1507 32262 1545 32296
rect 1579 32262 1617 32296
rect 1651 32262 1689 32296
rect 1723 32262 1729 32296
rect 315 32223 1729 32262
rect 315 32189 321 32223
rect 355 32189 393 32223
rect 427 32189 465 32223
rect 499 32189 537 32223
rect 571 32189 609 32223
rect 643 32189 681 32223
rect 715 32189 753 32223
rect 787 32189 825 32223
rect 859 32189 897 32223
rect 931 32189 969 32223
rect 1003 32189 1041 32223
rect 1075 32189 1113 32223
rect 1147 32189 1185 32223
rect 1219 32189 1257 32223
rect 1291 32189 1329 32223
rect 1363 32189 1401 32223
rect 1435 32189 1473 32223
rect 1507 32189 1545 32223
rect 1579 32189 1617 32223
rect 1651 32189 1689 32223
rect 1723 32189 1729 32223
rect 315 32150 1729 32189
rect 315 32116 321 32150
rect 355 32116 393 32150
rect 427 32116 465 32150
rect 499 32116 537 32150
rect 571 32116 609 32150
rect 643 32116 681 32150
rect 715 32116 753 32150
rect 787 32116 825 32150
rect 859 32116 897 32150
rect 931 32116 969 32150
rect 1003 32116 1041 32150
rect 1075 32116 1113 32150
rect 1147 32116 1185 32150
rect 1219 32116 1257 32150
rect 1291 32116 1329 32150
rect 1363 32116 1401 32150
rect 1435 32116 1473 32150
rect 1507 32116 1545 32150
rect 1579 32116 1617 32150
rect 1651 32116 1689 32150
rect 1723 32116 1729 32150
rect 315 32077 1729 32116
rect 315 32043 321 32077
rect 355 32043 393 32077
rect 427 32043 465 32077
rect 499 32043 537 32077
rect 571 32043 609 32077
rect 643 32043 681 32077
rect 715 32043 753 32077
rect 787 32043 825 32077
rect 859 32043 897 32077
rect 931 32043 969 32077
rect 1003 32043 1041 32077
rect 1075 32043 1113 32077
rect 1147 32043 1185 32077
rect 1219 32043 1257 32077
rect 1291 32043 1329 32077
rect 1363 32043 1401 32077
rect 1435 32043 1473 32077
rect 1507 32043 1545 32077
rect 1579 32043 1617 32077
rect 1651 32043 1689 32077
rect 1723 32043 1729 32077
rect 315 32004 1729 32043
rect 315 31970 321 32004
rect 355 31970 393 32004
rect 427 31970 465 32004
rect 499 31970 537 32004
rect 571 31970 609 32004
rect 643 31970 681 32004
rect 715 31970 753 32004
rect 787 31970 825 32004
rect 859 31970 897 32004
rect 931 31970 969 32004
rect 1003 31970 1041 32004
rect 1075 31970 1113 32004
rect 1147 31970 1185 32004
rect 1219 31970 1257 32004
rect 1291 31970 1329 32004
rect 1363 31970 1401 32004
rect 1435 31970 1473 32004
rect 1507 31970 1545 32004
rect 1579 31970 1617 32004
rect 1651 31970 1689 32004
rect 1723 31970 1729 32004
rect 315 31931 1729 31970
rect 315 31897 321 31931
rect 355 31897 393 31931
rect 427 31897 465 31931
rect 499 31897 537 31931
rect 571 31897 609 31931
rect 643 31897 681 31931
rect 715 31897 753 31931
rect 787 31897 825 31931
rect 859 31897 897 31931
rect 931 31897 969 31931
rect 1003 31897 1041 31931
rect 1075 31897 1113 31931
rect 1147 31897 1185 31931
rect 1219 31897 1257 31931
rect 1291 31897 1329 31931
rect 1363 31897 1401 31931
rect 1435 31897 1473 31931
rect 1507 31897 1545 31931
rect 1579 31897 1617 31931
rect 1651 31897 1689 31931
rect 1723 31897 1729 31931
rect 315 31858 1729 31897
rect 315 31824 321 31858
rect 355 31824 393 31858
rect 427 31824 465 31858
rect 499 31824 537 31858
rect 571 31824 609 31858
rect 643 31824 681 31858
rect 715 31824 753 31858
rect 787 31824 825 31858
rect 859 31824 897 31858
rect 931 31824 969 31858
rect 1003 31824 1041 31858
rect 1075 31824 1113 31858
rect 1147 31824 1185 31858
rect 1219 31824 1257 31858
rect 1291 31824 1329 31858
rect 1363 31824 1401 31858
rect 1435 31824 1473 31858
rect 1507 31824 1545 31858
rect 1579 31824 1617 31858
rect 1651 31824 1689 31858
rect 1723 31824 1729 31858
rect 315 31785 1729 31824
rect 315 31751 321 31785
rect 355 31751 393 31785
rect 427 31751 465 31785
rect 499 31751 537 31785
rect 571 31751 609 31785
rect 643 31751 681 31785
rect 715 31751 753 31785
rect 787 31751 825 31785
rect 859 31751 897 31785
rect 931 31751 969 31785
rect 1003 31751 1041 31785
rect 1075 31751 1113 31785
rect 1147 31751 1185 31785
rect 1219 31751 1257 31785
rect 1291 31751 1329 31785
rect 1363 31751 1401 31785
rect 1435 31751 1473 31785
rect 1507 31751 1545 31785
rect 1579 31751 1617 31785
rect 1651 31751 1689 31785
rect 1723 31751 1729 31785
rect 315 31712 1729 31751
rect 315 31678 321 31712
rect 355 31678 393 31712
rect 427 31678 465 31712
rect 499 31678 537 31712
rect 571 31678 609 31712
rect 643 31678 681 31712
rect 715 31678 753 31712
rect 787 31678 825 31712
rect 859 31678 897 31712
rect 931 31678 969 31712
rect 1003 31678 1041 31712
rect 1075 31678 1113 31712
rect 1147 31678 1185 31712
rect 1219 31678 1257 31712
rect 1291 31678 1329 31712
rect 1363 31678 1401 31712
rect 1435 31678 1473 31712
rect 1507 31678 1545 31712
rect 1579 31678 1617 31712
rect 1651 31678 1689 31712
rect 1723 31678 1729 31712
rect 315 31639 1729 31678
rect 315 31605 321 31639
rect 355 31605 393 31639
rect 427 31605 465 31639
rect 499 31605 537 31639
rect 571 31605 609 31639
rect 643 31605 681 31639
rect 715 31605 753 31639
rect 787 31605 825 31639
rect 859 31605 897 31639
rect 931 31605 969 31639
rect 1003 31605 1041 31639
rect 1075 31605 1113 31639
rect 1147 31605 1185 31639
rect 1219 31605 1257 31639
rect 1291 31605 1329 31639
rect 1363 31605 1401 31639
rect 1435 31605 1473 31639
rect 1507 31605 1545 31639
rect 1579 31605 1617 31639
rect 1651 31605 1689 31639
rect 1723 31605 1729 31639
rect 315 31566 1729 31605
rect 315 31532 321 31566
rect 355 31532 393 31566
rect 427 31532 465 31566
rect 499 31532 537 31566
rect 571 31532 609 31566
rect 643 31532 681 31566
rect 715 31532 753 31566
rect 787 31532 825 31566
rect 859 31532 897 31566
rect 931 31532 969 31566
rect 1003 31532 1041 31566
rect 1075 31532 1113 31566
rect 1147 31532 1185 31566
rect 1219 31532 1257 31566
rect 1291 31532 1329 31566
rect 1363 31532 1401 31566
rect 1435 31532 1473 31566
rect 1507 31532 1545 31566
rect 1579 31532 1617 31566
rect 1651 31532 1689 31566
rect 1723 31532 1729 31566
rect 315 31493 1729 31532
rect 315 31459 321 31493
rect 355 31459 393 31493
rect 427 31459 465 31493
rect 499 31459 537 31493
rect 571 31459 609 31493
rect 643 31459 681 31493
rect 715 31459 753 31493
rect 787 31459 825 31493
rect 859 31459 897 31493
rect 931 31459 969 31493
rect 1003 31459 1041 31493
rect 1075 31459 1113 31493
rect 1147 31459 1185 31493
rect 1219 31459 1257 31493
rect 1291 31459 1329 31493
rect 1363 31459 1401 31493
rect 1435 31459 1473 31493
rect 1507 31459 1545 31493
rect 1579 31459 1617 31493
rect 1651 31459 1689 31493
rect 1723 31459 1729 31493
rect 315 31420 1729 31459
rect 315 31386 321 31420
rect 355 31386 393 31420
rect 427 31386 465 31420
rect 499 31386 537 31420
rect 571 31386 609 31420
rect 643 31386 681 31420
rect 715 31386 753 31420
rect 787 31386 825 31420
rect 859 31386 897 31420
rect 931 31386 969 31420
rect 1003 31386 1041 31420
rect 1075 31386 1113 31420
rect 1147 31386 1185 31420
rect 1219 31386 1257 31420
rect 1291 31386 1329 31420
rect 1363 31386 1401 31420
rect 1435 31386 1473 31420
rect 1507 31386 1545 31420
rect 1579 31386 1617 31420
rect 1651 31386 1689 31420
rect 1723 31386 1729 31420
rect 315 31347 1729 31386
rect 315 31313 321 31347
rect 355 31313 393 31347
rect 427 31313 465 31347
rect 499 31313 537 31347
rect 571 31313 609 31347
rect 643 31313 681 31347
rect 715 31313 753 31347
rect 787 31313 825 31347
rect 859 31313 897 31347
rect 931 31313 969 31347
rect 1003 31313 1041 31347
rect 1075 31313 1113 31347
rect 1147 31313 1185 31347
rect 1219 31313 1257 31347
rect 1291 31313 1329 31347
rect 1363 31313 1401 31347
rect 1435 31313 1473 31347
rect 1507 31313 1545 31347
rect 1579 31313 1617 31347
rect 1651 31313 1689 31347
rect 1723 31313 1729 31347
rect 315 31274 1729 31313
rect 315 31240 321 31274
rect 355 31240 393 31274
rect 427 31240 465 31274
rect 499 31240 537 31274
rect 571 31240 609 31274
rect 643 31240 681 31274
rect 715 31240 753 31274
rect 787 31240 825 31274
rect 859 31240 897 31274
rect 931 31240 969 31274
rect 1003 31240 1041 31274
rect 1075 31240 1113 31274
rect 1147 31240 1185 31274
rect 1219 31240 1257 31274
rect 1291 31240 1329 31274
rect 1363 31240 1401 31274
rect 1435 31240 1473 31274
rect 1507 31240 1545 31274
rect 1579 31240 1617 31274
rect 1651 31240 1689 31274
rect 1723 31240 1729 31274
rect 315 31201 1729 31240
rect 315 31167 321 31201
rect 355 31167 393 31201
rect 427 31167 465 31201
rect 499 31167 537 31201
rect 571 31167 609 31201
rect 643 31167 681 31201
rect 715 31167 753 31201
rect 787 31167 825 31201
rect 859 31167 897 31201
rect 931 31167 969 31201
rect 1003 31167 1041 31201
rect 1075 31167 1113 31201
rect 1147 31167 1185 31201
rect 1219 31167 1257 31201
rect 1291 31167 1329 31201
rect 1363 31167 1401 31201
rect 1435 31167 1473 31201
rect 1507 31167 1545 31201
rect 1579 31167 1617 31201
rect 1651 31167 1689 31201
rect 1723 31167 1729 31201
rect 315 31128 1729 31167
rect 315 31094 321 31128
rect 355 31094 393 31128
rect 427 31094 465 31128
rect 499 31094 537 31128
rect 571 31094 609 31128
rect 643 31094 681 31128
rect 715 31094 753 31128
rect 787 31094 825 31128
rect 859 31094 897 31128
rect 931 31094 969 31128
rect 1003 31094 1041 31128
rect 1075 31094 1113 31128
rect 1147 31094 1185 31128
rect 1219 31094 1257 31128
rect 1291 31094 1329 31128
rect 1363 31094 1401 31128
rect 1435 31094 1473 31128
rect 1507 31094 1545 31128
rect 1579 31094 1617 31128
rect 1651 31094 1689 31128
rect 1723 31094 1729 31128
rect 315 31055 1729 31094
rect 315 31021 321 31055
rect 355 31021 393 31055
rect 427 31021 465 31055
rect 499 31021 537 31055
rect 571 31021 609 31055
rect 643 31021 681 31055
rect 715 31021 753 31055
rect 787 31021 825 31055
rect 859 31021 897 31055
rect 931 31021 969 31055
rect 1003 31021 1041 31055
rect 1075 31021 1113 31055
rect 1147 31021 1185 31055
rect 1219 31021 1257 31055
rect 1291 31021 1329 31055
rect 1363 31021 1401 31055
rect 1435 31021 1473 31055
rect 1507 31021 1545 31055
rect 1579 31021 1617 31055
rect 1651 31021 1689 31055
rect 1723 31021 1729 31055
rect 315 30982 1729 31021
rect 315 30948 321 30982
rect 355 30948 393 30982
rect 427 30948 465 30982
rect 499 30948 537 30982
rect 571 30948 609 30982
rect 643 30948 681 30982
rect 715 30948 753 30982
rect 787 30948 825 30982
rect 859 30948 897 30982
rect 931 30948 969 30982
rect 1003 30948 1041 30982
rect 1075 30948 1113 30982
rect 1147 30948 1185 30982
rect 1219 30948 1257 30982
rect 1291 30948 1329 30982
rect 1363 30948 1401 30982
rect 1435 30948 1473 30982
rect 1507 30948 1545 30982
rect 1579 30948 1617 30982
rect 1651 30948 1689 30982
rect 1723 30948 1729 30982
rect 315 30909 1729 30948
rect 315 30875 321 30909
rect 355 30875 393 30909
rect 427 30875 465 30909
rect 499 30875 537 30909
rect 571 30875 609 30909
rect 643 30875 681 30909
rect 715 30875 753 30909
rect 787 30875 825 30909
rect 859 30875 897 30909
rect 931 30875 969 30909
rect 1003 30875 1041 30909
rect 1075 30875 1113 30909
rect 1147 30875 1185 30909
rect 1219 30875 1257 30909
rect 1291 30875 1329 30909
rect 1363 30875 1401 30909
rect 1435 30875 1473 30909
rect 1507 30875 1545 30909
rect 1579 30875 1617 30909
rect 1651 30875 1689 30909
rect 1723 30875 1729 30909
rect 315 30836 1729 30875
rect 315 30802 321 30836
rect 355 30802 393 30836
rect 427 30802 465 30836
rect 499 30802 537 30836
rect 571 30802 609 30836
rect 643 30802 681 30836
rect 715 30802 753 30836
rect 787 30802 825 30836
rect 859 30802 897 30836
rect 931 30802 969 30836
rect 1003 30802 1041 30836
rect 1075 30802 1113 30836
rect 1147 30802 1185 30836
rect 1219 30802 1257 30836
rect 1291 30802 1329 30836
rect 1363 30802 1401 30836
rect 1435 30802 1473 30836
rect 1507 30802 1545 30836
rect 1579 30802 1617 30836
rect 1651 30802 1689 30836
rect 1723 30802 1729 30836
rect 315 30763 1729 30802
rect 315 30729 321 30763
rect 355 30729 393 30763
rect 427 30729 465 30763
rect 499 30729 537 30763
rect 571 30729 609 30763
rect 643 30729 681 30763
rect 715 30729 753 30763
rect 787 30729 825 30763
rect 859 30729 897 30763
rect 931 30729 969 30763
rect 1003 30729 1041 30763
rect 1075 30729 1113 30763
rect 1147 30729 1185 30763
rect 1219 30729 1257 30763
rect 1291 30729 1329 30763
rect 1363 30729 1401 30763
rect 1435 30729 1473 30763
rect 1507 30729 1545 30763
rect 1579 30729 1617 30763
rect 1651 30729 1689 30763
rect 1723 30729 1729 30763
rect 315 30690 1729 30729
rect 315 30656 321 30690
rect 355 30656 393 30690
rect 427 30656 465 30690
rect 499 30656 537 30690
rect 571 30656 609 30690
rect 643 30656 681 30690
rect 715 30656 753 30690
rect 787 30656 825 30690
rect 859 30656 897 30690
rect 931 30656 969 30690
rect 1003 30656 1041 30690
rect 1075 30656 1113 30690
rect 1147 30656 1185 30690
rect 1219 30656 1257 30690
rect 1291 30656 1329 30690
rect 1363 30656 1401 30690
rect 1435 30656 1473 30690
rect 1507 30656 1545 30690
rect 1579 30656 1617 30690
rect 1651 30656 1689 30690
rect 1723 30656 1729 30690
rect 315 30617 1729 30656
rect 315 30583 321 30617
rect 355 30583 393 30617
rect 427 30583 465 30617
rect 499 30583 537 30617
rect 571 30583 609 30617
rect 643 30583 681 30617
rect 715 30583 753 30617
rect 787 30583 825 30617
rect 859 30583 897 30617
rect 931 30583 969 30617
rect 1003 30583 1041 30617
rect 1075 30583 1113 30617
rect 1147 30583 1185 30617
rect 1219 30583 1257 30617
rect 1291 30583 1329 30617
rect 1363 30583 1401 30617
rect 1435 30583 1473 30617
rect 1507 30583 1545 30617
rect 1579 30583 1617 30617
rect 1651 30583 1689 30617
rect 1723 30583 1729 30617
rect 315 30544 1729 30583
rect 315 30510 321 30544
rect 355 30510 393 30544
rect 427 30510 465 30544
rect 499 30510 537 30544
rect 571 30510 609 30544
rect 643 30510 681 30544
rect 715 30510 753 30544
rect 787 30510 825 30544
rect 859 30510 897 30544
rect 931 30510 969 30544
rect 1003 30510 1041 30544
rect 1075 30510 1113 30544
rect 1147 30510 1185 30544
rect 1219 30510 1257 30544
rect 1291 30510 1329 30544
rect 1363 30510 1401 30544
rect 1435 30510 1473 30544
rect 1507 30510 1545 30544
rect 1579 30510 1617 30544
rect 1651 30510 1689 30544
rect 1723 30510 1729 30544
rect 315 30471 1729 30510
rect 315 30437 321 30471
rect 355 30437 393 30471
rect 427 30437 465 30471
rect 499 30437 537 30471
rect 571 30437 609 30471
rect 643 30437 681 30471
rect 715 30437 753 30471
rect 787 30437 825 30471
rect 859 30437 897 30471
rect 931 30437 969 30471
rect 1003 30437 1041 30471
rect 1075 30437 1113 30471
rect 1147 30437 1185 30471
rect 1219 30437 1257 30471
rect 1291 30437 1329 30471
rect 1363 30437 1401 30471
rect 1435 30437 1473 30471
rect 1507 30437 1545 30471
rect 1579 30437 1617 30471
rect 1651 30437 1689 30471
rect 1723 30437 1729 30471
rect 315 30398 1729 30437
rect 315 30364 321 30398
rect 355 30364 393 30398
rect 427 30364 465 30398
rect 499 30364 537 30398
rect 571 30364 609 30398
rect 643 30364 681 30398
rect 715 30364 753 30398
rect 787 30364 825 30398
rect 859 30364 897 30398
rect 931 30364 969 30398
rect 1003 30364 1041 30398
rect 1075 30364 1113 30398
rect 1147 30364 1185 30398
rect 1219 30364 1257 30398
rect 1291 30364 1329 30398
rect 1363 30364 1401 30398
rect 1435 30364 1473 30398
rect 1507 30364 1545 30398
rect 1579 30364 1617 30398
rect 1651 30364 1689 30398
rect 1723 30364 1729 30398
rect 315 30325 1729 30364
rect 315 30291 321 30325
rect 355 30291 393 30325
rect 427 30291 465 30325
rect 499 30291 537 30325
rect 571 30291 609 30325
rect 643 30291 681 30325
rect 715 30291 753 30325
rect 787 30291 825 30325
rect 859 30291 897 30325
rect 931 30291 969 30325
rect 1003 30291 1041 30325
rect 1075 30291 1113 30325
rect 1147 30291 1185 30325
rect 1219 30291 1257 30325
rect 1291 30291 1329 30325
rect 1363 30291 1401 30325
rect 1435 30291 1473 30325
rect 1507 30291 1545 30325
rect 1579 30291 1617 30325
rect 1651 30291 1689 30325
rect 1723 30291 1729 30325
rect 315 30252 1729 30291
rect 315 30218 321 30252
rect 355 30218 393 30252
rect 427 30218 465 30252
rect 499 30218 537 30252
rect 571 30218 609 30252
rect 643 30218 681 30252
rect 715 30218 753 30252
rect 787 30218 825 30252
rect 859 30218 897 30252
rect 931 30218 969 30252
rect 1003 30218 1041 30252
rect 1075 30218 1113 30252
rect 1147 30218 1185 30252
rect 1219 30218 1257 30252
rect 1291 30218 1329 30252
rect 1363 30218 1401 30252
rect 1435 30218 1473 30252
rect 1507 30218 1545 30252
rect 1579 30218 1617 30252
rect 1651 30218 1689 30252
rect 1723 30218 1729 30252
rect 315 30179 1729 30218
rect 315 30145 321 30179
rect 355 30145 393 30179
rect 427 30145 465 30179
rect 499 30145 537 30179
rect 571 30145 609 30179
rect 643 30145 681 30179
rect 715 30145 753 30179
rect 787 30145 825 30179
rect 859 30145 897 30179
rect 931 30145 969 30179
rect 1003 30145 1041 30179
rect 1075 30145 1113 30179
rect 1147 30145 1185 30179
rect 1219 30145 1257 30179
rect 1291 30145 1329 30179
rect 1363 30145 1401 30179
rect 1435 30145 1473 30179
rect 1507 30145 1545 30179
rect 1579 30145 1617 30179
rect 1651 30145 1689 30179
rect 1723 30145 1729 30179
rect 315 30106 1729 30145
rect 315 30072 321 30106
rect 355 30072 393 30106
rect 427 30072 465 30106
rect 499 30072 537 30106
rect 571 30072 609 30106
rect 643 30072 681 30106
rect 715 30072 753 30106
rect 787 30072 825 30106
rect 859 30072 897 30106
rect 931 30072 969 30106
rect 1003 30072 1041 30106
rect 1075 30072 1113 30106
rect 1147 30072 1185 30106
rect 1219 30072 1257 30106
rect 1291 30072 1329 30106
rect 1363 30072 1401 30106
rect 1435 30072 1473 30106
rect 1507 30072 1545 30106
rect 1579 30072 1617 30106
rect 1651 30072 1689 30106
rect 1723 30072 1729 30106
rect 315 30033 1729 30072
rect 315 29999 321 30033
rect 355 29999 393 30033
rect 427 29999 465 30033
rect 499 29999 537 30033
rect 571 29999 609 30033
rect 643 29999 681 30033
rect 715 29999 753 30033
rect 787 29999 825 30033
rect 859 29999 897 30033
rect 931 29999 969 30033
rect 1003 29999 1041 30033
rect 1075 29999 1113 30033
rect 1147 29999 1185 30033
rect 1219 29999 1257 30033
rect 1291 29999 1329 30033
rect 1363 29999 1401 30033
rect 1435 29999 1473 30033
rect 1507 29999 1545 30033
rect 1579 29999 1617 30033
rect 1651 29999 1689 30033
rect 1723 29999 1729 30033
rect 315 29960 1729 29999
rect 315 29926 321 29960
rect 355 29926 393 29960
rect 427 29926 465 29960
rect 499 29926 537 29960
rect 571 29926 609 29960
rect 643 29926 681 29960
rect 715 29926 753 29960
rect 787 29926 825 29960
rect 859 29926 897 29960
rect 931 29926 969 29960
rect 1003 29926 1041 29960
rect 1075 29926 1113 29960
rect 1147 29926 1185 29960
rect 1219 29926 1257 29960
rect 1291 29926 1329 29960
rect 1363 29926 1401 29960
rect 1435 29926 1473 29960
rect 1507 29926 1545 29960
rect 1579 29926 1617 29960
rect 1651 29926 1689 29960
rect 1723 29926 1729 29960
rect 315 29887 1729 29926
rect 315 29853 321 29887
rect 355 29853 393 29887
rect 427 29853 465 29887
rect 499 29853 537 29887
rect 571 29853 609 29887
rect 643 29853 681 29887
rect 715 29853 753 29887
rect 787 29853 825 29887
rect 859 29853 897 29887
rect 931 29853 969 29887
rect 1003 29853 1041 29887
rect 1075 29853 1113 29887
rect 1147 29853 1185 29887
rect 1219 29853 1257 29887
rect 1291 29853 1329 29887
rect 1363 29853 1401 29887
rect 1435 29853 1473 29887
rect 1507 29853 1545 29887
rect 1579 29853 1617 29887
rect 1651 29853 1689 29887
rect 1723 29853 1729 29887
rect 315 29814 1729 29853
rect 315 29780 321 29814
rect 355 29780 393 29814
rect 427 29780 465 29814
rect 499 29780 537 29814
rect 571 29780 609 29814
rect 643 29780 681 29814
rect 715 29780 753 29814
rect 787 29780 825 29814
rect 859 29780 897 29814
rect 931 29780 969 29814
rect 1003 29780 1041 29814
rect 1075 29780 1113 29814
rect 1147 29780 1185 29814
rect 1219 29780 1257 29814
rect 1291 29780 1329 29814
rect 1363 29780 1401 29814
rect 1435 29780 1473 29814
rect 1507 29780 1545 29814
rect 1579 29780 1617 29814
rect 1651 29780 1689 29814
rect 1723 29780 1729 29814
rect 315 29741 1729 29780
rect 315 29707 321 29741
rect 355 29707 393 29741
rect 427 29707 465 29741
rect 499 29707 537 29741
rect 571 29707 609 29741
rect 643 29707 681 29741
rect 715 29707 753 29741
rect 787 29707 825 29741
rect 859 29707 897 29741
rect 931 29707 969 29741
rect 1003 29707 1041 29741
rect 1075 29707 1113 29741
rect 1147 29707 1185 29741
rect 1219 29707 1257 29741
rect 1291 29707 1329 29741
rect 1363 29707 1401 29741
rect 1435 29707 1473 29741
rect 1507 29707 1545 29741
rect 1579 29707 1617 29741
rect 1651 29707 1689 29741
rect 1723 29707 1729 29741
rect 315 29668 1729 29707
rect 315 29634 321 29668
rect 355 29634 393 29668
rect 427 29634 465 29668
rect 499 29634 537 29668
rect 571 29634 609 29668
rect 643 29634 681 29668
rect 715 29634 753 29668
rect 787 29634 825 29668
rect 859 29634 897 29668
rect 931 29634 969 29668
rect 1003 29634 1041 29668
rect 1075 29634 1113 29668
rect 1147 29634 1185 29668
rect 1219 29634 1257 29668
rect 1291 29634 1329 29668
rect 1363 29634 1401 29668
rect 1435 29634 1473 29668
rect 1507 29634 1545 29668
rect 1579 29634 1617 29668
rect 1651 29634 1689 29668
rect 1723 29634 1729 29668
rect 315 29602 1729 29634
rect 7870 39943 9284 39975
rect 7870 33357 7876 39943
rect 9278 33357 9284 39943
rect 7870 33318 9284 33357
rect 7870 33284 7876 33318
rect 7910 33284 7948 33318
rect 7982 33284 8020 33318
rect 8054 33284 8092 33318
rect 8126 33284 8164 33318
rect 8198 33284 8236 33318
rect 8270 33284 8308 33318
rect 8342 33284 8380 33318
rect 8414 33284 8452 33318
rect 8486 33284 8524 33318
rect 8558 33284 8596 33318
rect 8630 33284 8668 33318
rect 8702 33284 8740 33318
rect 8774 33284 8812 33318
rect 8846 33284 8884 33318
rect 8918 33284 8956 33318
rect 8990 33284 9028 33318
rect 9062 33284 9100 33318
rect 9134 33284 9172 33318
rect 9206 33284 9244 33318
rect 9278 33284 9284 33318
rect 7870 33245 9284 33284
rect 7870 33211 7876 33245
rect 7910 33211 7948 33245
rect 7982 33211 8020 33245
rect 8054 33211 8092 33245
rect 8126 33211 8164 33245
rect 8198 33211 8236 33245
rect 8270 33211 8308 33245
rect 8342 33211 8380 33245
rect 8414 33211 8452 33245
rect 8486 33211 8524 33245
rect 8558 33211 8596 33245
rect 8630 33211 8668 33245
rect 8702 33211 8740 33245
rect 8774 33211 8812 33245
rect 8846 33211 8884 33245
rect 8918 33211 8956 33245
rect 8990 33211 9028 33245
rect 9062 33211 9100 33245
rect 9134 33211 9172 33245
rect 9206 33211 9244 33245
rect 9278 33211 9284 33245
rect 7870 33172 9284 33211
rect 7870 33138 7876 33172
rect 7910 33138 7948 33172
rect 7982 33138 8020 33172
rect 8054 33138 8092 33172
rect 8126 33138 8164 33172
rect 8198 33138 8236 33172
rect 8270 33138 8308 33172
rect 8342 33138 8380 33172
rect 8414 33138 8452 33172
rect 8486 33138 8524 33172
rect 8558 33138 8596 33172
rect 8630 33138 8668 33172
rect 8702 33138 8740 33172
rect 8774 33138 8812 33172
rect 8846 33138 8884 33172
rect 8918 33138 8956 33172
rect 8990 33138 9028 33172
rect 9062 33138 9100 33172
rect 9134 33138 9172 33172
rect 9206 33138 9244 33172
rect 9278 33138 9284 33172
rect 7870 33099 9284 33138
rect 7870 33065 7876 33099
rect 7910 33065 7948 33099
rect 7982 33065 8020 33099
rect 8054 33065 8092 33099
rect 8126 33065 8164 33099
rect 8198 33065 8236 33099
rect 8270 33065 8308 33099
rect 8342 33065 8380 33099
rect 8414 33065 8452 33099
rect 8486 33065 8524 33099
rect 8558 33065 8596 33099
rect 8630 33065 8668 33099
rect 8702 33065 8740 33099
rect 8774 33065 8812 33099
rect 8846 33065 8884 33099
rect 8918 33065 8956 33099
rect 8990 33065 9028 33099
rect 9062 33065 9100 33099
rect 9134 33065 9172 33099
rect 9206 33065 9244 33099
rect 9278 33065 9284 33099
rect 7870 33026 9284 33065
rect 7870 32992 7876 33026
rect 7910 32992 7948 33026
rect 7982 32992 8020 33026
rect 8054 32992 8092 33026
rect 8126 32992 8164 33026
rect 8198 32992 8236 33026
rect 8270 32992 8308 33026
rect 8342 32992 8380 33026
rect 8414 32992 8452 33026
rect 8486 32992 8524 33026
rect 8558 32992 8596 33026
rect 8630 32992 8668 33026
rect 8702 32992 8740 33026
rect 8774 32992 8812 33026
rect 8846 32992 8884 33026
rect 8918 32992 8956 33026
rect 8990 32992 9028 33026
rect 9062 32992 9100 33026
rect 9134 32992 9172 33026
rect 9206 32992 9244 33026
rect 9278 32992 9284 33026
rect 7870 32953 9284 32992
rect 7870 32919 7876 32953
rect 7910 32919 7948 32953
rect 7982 32919 8020 32953
rect 8054 32919 8092 32953
rect 8126 32919 8164 32953
rect 8198 32919 8236 32953
rect 8270 32919 8308 32953
rect 8342 32919 8380 32953
rect 8414 32919 8452 32953
rect 8486 32919 8524 32953
rect 8558 32919 8596 32953
rect 8630 32919 8668 32953
rect 8702 32919 8740 32953
rect 8774 32919 8812 32953
rect 8846 32919 8884 32953
rect 8918 32919 8956 32953
rect 8990 32919 9028 32953
rect 9062 32919 9100 32953
rect 9134 32919 9172 32953
rect 9206 32919 9244 32953
rect 9278 32919 9284 32953
rect 7870 32880 9284 32919
rect 7870 32846 7876 32880
rect 7910 32846 7948 32880
rect 7982 32846 8020 32880
rect 8054 32846 8092 32880
rect 8126 32846 8164 32880
rect 8198 32846 8236 32880
rect 8270 32846 8308 32880
rect 8342 32846 8380 32880
rect 8414 32846 8452 32880
rect 8486 32846 8524 32880
rect 8558 32846 8596 32880
rect 8630 32846 8668 32880
rect 8702 32846 8740 32880
rect 8774 32846 8812 32880
rect 8846 32846 8884 32880
rect 8918 32846 8956 32880
rect 8990 32846 9028 32880
rect 9062 32846 9100 32880
rect 9134 32846 9172 32880
rect 9206 32846 9244 32880
rect 9278 32846 9284 32880
rect 7870 32807 9284 32846
rect 7870 32773 7876 32807
rect 7910 32773 7948 32807
rect 7982 32773 8020 32807
rect 8054 32773 8092 32807
rect 8126 32773 8164 32807
rect 8198 32773 8236 32807
rect 8270 32773 8308 32807
rect 8342 32773 8380 32807
rect 8414 32773 8452 32807
rect 8486 32773 8524 32807
rect 8558 32773 8596 32807
rect 8630 32773 8668 32807
rect 8702 32773 8740 32807
rect 8774 32773 8812 32807
rect 8846 32773 8884 32807
rect 8918 32773 8956 32807
rect 8990 32773 9028 32807
rect 9062 32773 9100 32807
rect 9134 32773 9172 32807
rect 9206 32773 9244 32807
rect 9278 32773 9284 32807
rect 7870 32734 9284 32773
rect 7870 32700 7876 32734
rect 7910 32700 7948 32734
rect 7982 32700 8020 32734
rect 8054 32700 8092 32734
rect 8126 32700 8164 32734
rect 8198 32700 8236 32734
rect 8270 32700 8308 32734
rect 8342 32700 8380 32734
rect 8414 32700 8452 32734
rect 8486 32700 8524 32734
rect 8558 32700 8596 32734
rect 8630 32700 8668 32734
rect 8702 32700 8740 32734
rect 8774 32700 8812 32734
rect 8846 32700 8884 32734
rect 8918 32700 8956 32734
rect 8990 32700 9028 32734
rect 9062 32700 9100 32734
rect 9134 32700 9172 32734
rect 9206 32700 9244 32734
rect 9278 32700 9284 32734
rect 7870 32661 9284 32700
rect 7870 32627 7876 32661
rect 7910 32627 7948 32661
rect 7982 32627 8020 32661
rect 8054 32627 8092 32661
rect 8126 32627 8164 32661
rect 8198 32627 8236 32661
rect 8270 32627 8308 32661
rect 8342 32627 8380 32661
rect 8414 32627 8452 32661
rect 8486 32627 8524 32661
rect 8558 32627 8596 32661
rect 8630 32627 8668 32661
rect 8702 32627 8740 32661
rect 8774 32627 8812 32661
rect 8846 32627 8884 32661
rect 8918 32627 8956 32661
rect 8990 32627 9028 32661
rect 9062 32627 9100 32661
rect 9134 32627 9172 32661
rect 9206 32627 9244 32661
rect 9278 32627 9284 32661
rect 7870 32588 9284 32627
rect 7870 32554 7876 32588
rect 7910 32554 7948 32588
rect 7982 32554 8020 32588
rect 8054 32554 8092 32588
rect 8126 32554 8164 32588
rect 8198 32554 8236 32588
rect 8270 32554 8308 32588
rect 8342 32554 8380 32588
rect 8414 32554 8452 32588
rect 8486 32554 8524 32588
rect 8558 32554 8596 32588
rect 8630 32554 8668 32588
rect 8702 32554 8740 32588
rect 8774 32554 8812 32588
rect 8846 32554 8884 32588
rect 8918 32554 8956 32588
rect 8990 32554 9028 32588
rect 9062 32554 9100 32588
rect 9134 32554 9172 32588
rect 9206 32554 9244 32588
rect 9278 32554 9284 32588
rect 7870 32515 9284 32554
rect 7870 32481 7876 32515
rect 7910 32481 7948 32515
rect 7982 32481 8020 32515
rect 8054 32481 8092 32515
rect 8126 32481 8164 32515
rect 8198 32481 8236 32515
rect 8270 32481 8308 32515
rect 8342 32481 8380 32515
rect 8414 32481 8452 32515
rect 8486 32481 8524 32515
rect 8558 32481 8596 32515
rect 8630 32481 8668 32515
rect 8702 32481 8740 32515
rect 8774 32481 8812 32515
rect 8846 32481 8884 32515
rect 8918 32481 8956 32515
rect 8990 32481 9028 32515
rect 9062 32481 9100 32515
rect 9134 32481 9172 32515
rect 9206 32481 9244 32515
rect 9278 32481 9284 32515
rect 7870 32442 9284 32481
rect 7870 32408 7876 32442
rect 7910 32408 7948 32442
rect 7982 32408 8020 32442
rect 8054 32408 8092 32442
rect 8126 32408 8164 32442
rect 8198 32408 8236 32442
rect 8270 32408 8308 32442
rect 8342 32408 8380 32442
rect 8414 32408 8452 32442
rect 8486 32408 8524 32442
rect 8558 32408 8596 32442
rect 8630 32408 8668 32442
rect 8702 32408 8740 32442
rect 8774 32408 8812 32442
rect 8846 32408 8884 32442
rect 8918 32408 8956 32442
rect 8990 32408 9028 32442
rect 9062 32408 9100 32442
rect 9134 32408 9172 32442
rect 9206 32408 9244 32442
rect 9278 32408 9284 32442
rect 7870 32369 9284 32408
rect 7870 32335 7876 32369
rect 7910 32335 7948 32369
rect 7982 32335 8020 32369
rect 8054 32335 8092 32369
rect 8126 32335 8164 32369
rect 8198 32335 8236 32369
rect 8270 32335 8308 32369
rect 8342 32335 8380 32369
rect 8414 32335 8452 32369
rect 8486 32335 8524 32369
rect 8558 32335 8596 32369
rect 8630 32335 8668 32369
rect 8702 32335 8740 32369
rect 8774 32335 8812 32369
rect 8846 32335 8884 32369
rect 8918 32335 8956 32369
rect 8990 32335 9028 32369
rect 9062 32335 9100 32369
rect 9134 32335 9172 32369
rect 9206 32335 9244 32369
rect 9278 32335 9284 32369
rect 7870 32296 9284 32335
rect 7870 32262 7876 32296
rect 7910 32262 7948 32296
rect 7982 32262 8020 32296
rect 8054 32262 8092 32296
rect 8126 32262 8164 32296
rect 8198 32262 8236 32296
rect 8270 32262 8308 32296
rect 8342 32262 8380 32296
rect 8414 32262 8452 32296
rect 8486 32262 8524 32296
rect 8558 32262 8596 32296
rect 8630 32262 8668 32296
rect 8702 32262 8740 32296
rect 8774 32262 8812 32296
rect 8846 32262 8884 32296
rect 8918 32262 8956 32296
rect 8990 32262 9028 32296
rect 9062 32262 9100 32296
rect 9134 32262 9172 32296
rect 9206 32262 9244 32296
rect 9278 32262 9284 32296
rect 7870 32223 9284 32262
rect 7870 32189 7876 32223
rect 7910 32189 7948 32223
rect 7982 32189 8020 32223
rect 8054 32189 8092 32223
rect 8126 32189 8164 32223
rect 8198 32189 8236 32223
rect 8270 32189 8308 32223
rect 8342 32189 8380 32223
rect 8414 32189 8452 32223
rect 8486 32189 8524 32223
rect 8558 32189 8596 32223
rect 8630 32189 8668 32223
rect 8702 32189 8740 32223
rect 8774 32189 8812 32223
rect 8846 32189 8884 32223
rect 8918 32189 8956 32223
rect 8990 32189 9028 32223
rect 9062 32189 9100 32223
rect 9134 32189 9172 32223
rect 9206 32189 9244 32223
rect 9278 32189 9284 32223
rect 7870 32150 9284 32189
rect 7870 32116 7876 32150
rect 7910 32116 7948 32150
rect 7982 32116 8020 32150
rect 8054 32116 8092 32150
rect 8126 32116 8164 32150
rect 8198 32116 8236 32150
rect 8270 32116 8308 32150
rect 8342 32116 8380 32150
rect 8414 32116 8452 32150
rect 8486 32116 8524 32150
rect 8558 32116 8596 32150
rect 8630 32116 8668 32150
rect 8702 32116 8740 32150
rect 8774 32116 8812 32150
rect 8846 32116 8884 32150
rect 8918 32116 8956 32150
rect 8990 32116 9028 32150
rect 9062 32116 9100 32150
rect 9134 32116 9172 32150
rect 9206 32116 9244 32150
rect 9278 32116 9284 32150
rect 7870 32077 9284 32116
rect 7870 32043 7876 32077
rect 7910 32043 7948 32077
rect 7982 32043 8020 32077
rect 8054 32043 8092 32077
rect 8126 32043 8164 32077
rect 8198 32043 8236 32077
rect 8270 32043 8308 32077
rect 8342 32043 8380 32077
rect 8414 32043 8452 32077
rect 8486 32043 8524 32077
rect 8558 32043 8596 32077
rect 8630 32043 8668 32077
rect 8702 32043 8740 32077
rect 8774 32043 8812 32077
rect 8846 32043 8884 32077
rect 8918 32043 8956 32077
rect 8990 32043 9028 32077
rect 9062 32043 9100 32077
rect 9134 32043 9172 32077
rect 9206 32043 9244 32077
rect 9278 32043 9284 32077
rect 7870 32004 9284 32043
rect 7870 31970 7876 32004
rect 7910 31970 7948 32004
rect 7982 31970 8020 32004
rect 8054 31970 8092 32004
rect 8126 31970 8164 32004
rect 8198 31970 8236 32004
rect 8270 31970 8308 32004
rect 8342 31970 8380 32004
rect 8414 31970 8452 32004
rect 8486 31970 8524 32004
rect 8558 31970 8596 32004
rect 8630 31970 8668 32004
rect 8702 31970 8740 32004
rect 8774 31970 8812 32004
rect 8846 31970 8884 32004
rect 8918 31970 8956 32004
rect 8990 31970 9028 32004
rect 9062 31970 9100 32004
rect 9134 31970 9172 32004
rect 9206 31970 9244 32004
rect 9278 31970 9284 32004
rect 7870 31931 9284 31970
rect 7870 31897 7876 31931
rect 7910 31897 7948 31931
rect 7982 31897 8020 31931
rect 8054 31897 8092 31931
rect 8126 31897 8164 31931
rect 8198 31897 8236 31931
rect 8270 31897 8308 31931
rect 8342 31897 8380 31931
rect 8414 31897 8452 31931
rect 8486 31897 8524 31931
rect 8558 31897 8596 31931
rect 8630 31897 8668 31931
rect 8702 31897 8740 31931
rect 8774 31897 8812 31931
rect 8846 31897 8884 31931
rect 8918 31897 8956 31931
rect 8990 31897 9028 31931
rect 9062 31897 9100 31931
rect 9134 31897 9172 31931
rect 9206 31897 9244 31931
rect 9278 31897 9284 31931
rect 7870 31858 9284 31897
rect 7870 31824 7876 31858
rect 7910 31824 7948 31858
rect 7982 31824 8020 31858
rect 8054 31824 8092 31858
rect 8126 31824 8164 31858
rect 8198 31824 8236 31858
rect 8270 31824 8308 31858
rect 8342 31824 8380 31858
rect 8414 31824 8452 31858
rect 8486 31824 8524 31858
rect 8558 31824 8596 31858
rect 8630 31824 8668 31858
rect 8702 31824 8740 31858
rect 8774 31824 8812 31858
rect 8846 31824 8884 31858
rect 8918 31824 8956 31858
rect 8990 31824 9028 31858
rect 9062 31824 9100 31858
rect 9134 31824 9172 31858
rect 9206 31824 9244 31858
rect 9278 31824 9284 31858
rect 7870 31785 9284 31824
rect 7870 31751 7876 31785
rect 7910 31751 7948 31785
rect 7982 31751 8020 31785
rect 8054 31751 8092 31785
rect 8126 31751 8164 31785
rect 8198 31751 8236 31785
rect 8270 31751 8308 31785
rect 8342 31751 8380 31785
rect 8414 31751 8452 31785
rect 8486 31751 8524 31785
rect 8558 31751 8596 31785
rect 8630 31751 8668 31785
rect 8702 31751 8740 31785
rect 8774 31751 8812 31785
rect 8846 31751 8884 31785
rect 8918 31751 8956 31785
rect 8990 31751 9028 31785
rect 9062 31751 9100 31785
rect 9134 31751 9172 31785
rect 9206 31751 9244 31785
rect 9278 31751 9284 31785
rect 7870 31712 9284 31751
rect 7870 31678 7876 31712
rect 7910 31678 7948 31712
rect 7982 31678 8020 31712
rect 8054 31678 8092 31712
rect 8126 31678 8164 31712
rect 8198 31678 8236 31712
rect 8270 31678 8308 31712
rect 8342 31678 8380 31712
rect 8414 31678 8452 31712
rect 8486 31678 8524 31712
rect 8558 31678 8596 31712
rect 8630 31678 8668 31712
rect 8702 31678 8740 31712
rect 8774 31678 8812 31712
rect 8846 31678 8884 31712
rect 8918 31678 8956 31712
rect 8990 31678 9028 31712
rect 9062 31678 9100 31712
rect 9134 31678 9172 31712
rect 9206 31678 9244 31712
rect 9278 31678 9284 31712
rect 7870 31639 9284 31678
rect 7870 31605 7876 31639
rect 7910 31605 7948 31639
rect 7982 31605 8020 31639
rect 8054 31605 8092 31639
rect 8126 31605 8164 31639
rect 8198 31605 8236 31639
rect 8270 31605 8308 31639
rect 8342 31605 8380 31639
rect 8414 31605 8452 31639
rect 8486 31605 8524 31639
rect 8558 31605 8596 31639
rect 8630 31605 8668 31639
rect 8702 31605 8740 31639
rect 8774 31605 8812 31639
rect 8846 31605 8884 31639
rect 8918 31605 8956 31639
rect 8990 31605 9028 31639
rect 9062 31605 9100 31639
rect 9134 31605 9172 31639
rect 9206 31605 9244 31639
rect 9278 31605 9284 31639
rect 7870 31566 9284 31605
rect 7870 31532 7876 31566
rect 7910 31532 7948 31566
rect 7982 31532 8020 31566
rect 8054 31532 8092 31566
rect 8126 31532 8164 31566
rect 8198 31532 8236 31566
rect 8270 31532 8308 31566
rect 8342 31532 8380 31566
rect 8414 31532 8452 31566
rect 8486 31532 8524 31566
rect 8558 31532 8596 31566
rect 8630 31532 8668 31566
rect 8702 31532 8740 31566
rect 8774 31532 8812 31566
rect 8846 31532 8884 31566
rect 8918 31532 8956 31566
rect 8990 31532 9028 31566
rect 9062 31532 9100 31566
rect 9134 31532 9172 31566
rect 9206 31532 9244 31566
rect 9278 31532 9284 31566
rect 7870 31493 9284 31532
rect 7870 31459 7876 31493
rect 7910 31459 7948 31493
rect 7982 31459 8020 31493
rect 8054 31459 8092 31493
rect 8126 31459 8164 31493
rect 8198 31459 8236 31493
rect 8270 31459 8308 31493
rect 8342 31459 8380 31493
rect 8414 31459 8452 31493
rect 8486 31459 8524 31493
rect 8558 31459 8596 31493
rect 8630 31459 8668 31493
rect 8702 31459 8740 31493
rect 8774 31459 8812 31493
rect 8846 31459 8884 31493
rect 8918 31459 8956 31493
rect 8990 31459 9028 31493
rect 9062 31459 9100 31493
rect 9134 31459 9172 31493
rect 9206 31459 9244 31493
rect 9278 31459 9284 31493
rect 7870 31420 9284 31459
rect 7870 31386 7876 31420
rect 7910 31386 7948 31420
rect 7982 31386 8020 31420
rect 8054 31386 8092 31420
rect 8126 31386 8164 31420
rect 8198 31386 8236 31420
rect 8270 31386 8308 31420
rect 8342 31386 8380 31420
rect 8414 31386 8452 31420
rect 8486 31386 8524 31420
rect 8558 31386 8596 31420
rect 8630 31386 8668 31420
rect 8702 31386 8740 31420
rect 8774 31386 8812 31420
rect 8846 31386 8884 31420
rect 8918 31386 8956 31420
rect 8990 31386 9028 31420
rect 9062 31386 9100 31420
rect 9134 31386 9172 31420
rect 9206 31386 9244 31420
rect 9278 31386 9284 31420
rect 7870 31347 9284 31386
rect 7870 31313 7876 31347
rect 7910 31313 7948 31347
rect 7982 31313 8020 31347
rect 8054 31313 8092 31347
rect 8126 31313 8164 31347
rect 8198 31313 8236 31347
rect 8270 31313 8308 31347
rect 8342 31313 8380 31347
rect 8414 31313 8452 31347
rect 8486 31313 8524 31347
rect 8558 31313 8596 31347
rect 8630 31313 8668 31347
rect 8702 31313 8740 31347
rect 8774 31313 8812 31347
rect 8846 31313 8884 31347
rect 8918 31313 8956 31347
rect 8990 31313 9028 31347
rect 9062 31313 9100 31347
rect 9134 31313 9172 31347
rect 9206 31313 9244 31347
rect 9278 31313 9284 31347
rect 7870 31274 9284 31313
rect 7870 31240 7876 31274
rect 7910 31240 7948 31274
rect 7982 31240 8020 31274
rect 8054 31240 8092 31274
rect 8126 31240 8164 31274
rect 8198 31240 8236 31274
rect 8270 31240 8308 31274
rect 8342 31240 8380 31274
rect 8414 31240 8452 31274
rect 8486 31240 8524 31274
rect 8558 31240 8596 31274
rect 8630 31240 8668 31274
rect 8702 31240 8740 31274
rect 8774 31240 8812 31274
rect 8846 31240 8884 31274
rect 8918 31240 8956 31274
rect 8990 31240 9028 31274
rect 9062 31240 9100 31274
rect 9134 31240 9172 31274
rect 9206 31240 9244 31274
rect 9278 31240 9284 31274
rect 7870 31201 9284 31240
rect 7870 31167 7876 31201
rect 7910 31167 7948 31201
rect 7982 31167 8020 31201
rect 8054 31167 8092 31201
rect 8126 31167 8164 31201
rect 8198 31167 8236 31201
rect 8270 31167 8308 31201
rect 8342 31167 8380 31201
rect 8414 31167 8452 31201
rect 8486 31167 8524 31201
rect 8558 31167 8596 31201
rect 8630 31167 8668 31201
rect 8702 31167 8740 31201
rect 8774 31167 8812 31201
rect 8846 31167 8884 31201
rect 8918 31167 8956 31201
rect 8990 31167 9028 31201
rect 9062 31167 9100 31201
rect 9134 31167 9172 31201
rect 9206 31167 9244 31201
rect 9278 31167 9284 31201
rect 7870 31128 9284 31167
rect 7870 31094 7876 31128
rect 7910 31094 7948 31128
rect 7982 31094 8020 31128
rect 8054 31094 8092 31128
rect 8126 31094 8164 31128
rect 8198 31094 8236 31128
rect 8270 31094 8308 31128
rect 8342 31094 8380 31128
rect 8414 31094 8452 31128
rect 8486 31094 8524 31128
rect 8558 31094 8596 31128
rect 8630 31094 8668 31128
rect 8702 31094 8740 31128
rect 8774 31094 8812 31128
rect 8846 31094 8884 31128
rect 8918 31094 8956 31128
rect 8990 31094 9028 31128
rect 9062 31094 9100 31128
rect 9134 31094 9172 31128
rect 9206 31094 9244 31128
rect 9278 31094 9284 31128
rect 7870 31055 9284 31094
rect 7870 31021 7876 31055
rect 7910 31021 7948 31055
rect 7982 31021 8020 31055
rect 8054 31021 8092 31055
rect 8126 31021 8164 31055
rect 8198 31021 8236 31055
rect 8270 31021 8308 31055
rect 8342 31021 8380 31055
rect 8414 31021 8452 31055
rect 8486 31021 8524 31055
rect 8558 31021 8596 31055
rect 8630 31021 8668 31055
rect 8702 31021 8740 31055
rect 8774 31021 8812 31055
rect 8846 31021 8884 31055
rect 8918 31021 8956 31055
rect 8990 31021 9028 31055
rect 9062 31021 9100 31055
rect 9134 31021 9172 31055
rect 9206 31021 9244 31055
rect 9278 31021 9284 31055
rect 7870 30982 9284 31021
rect 7870 30948 7876 30982
rect 7910 30948 7948 30982
rect 7982 30948 8020 30982
rect 8054 30948 8092 30982
rect 8126 30948 8164 30982
rect 8198 30948 8236 30982
rect 8270 30948 8308 30982
rect 8342 30948 8380 30982
rect 8414 30948 8452 30982
rect 8486 30948 8524 30982
rect 8558 30948 8596 30982
rect 8630 30948 8668 30982
rect 8702 30948 8740 30982
rect 8774 30948 8812 30982
rect 8846 30948 8884 30982
rect 8918 30948 8956 30982
rect 8990 30948 9028 30982
rect 9062 30948 9100 30982
rect 9134 30948 9172 30982
rect 9206 30948 9244 30982
rect 9278 30948 9284 30982
rect 7870 30909 9284 30948
rect 7870 30875 7876 30909
rect 7910 30875 7948 30909
rect 7982 30875 8020 30909
rect 8054 30875 8092 30909
rect 8126 30875 8164 30909
rect 8198 30875 8236 30909
rect 8270 30875 8308 30909
rect 8342 30875 8380 30909
rect 8414 30875 8452 30909
rect 8486 30875 8524 30909
rect 8558 30875 8596 30909
rect 8630 30875 8668 30909
rect 8702 30875 8740 30909
rect 8774 30875 8812 30909
rect 8846 30875 8884 30909
rect 8918 30875 8956 30909
rect 8990 30875 9028 30909
rect 9062 30875 9100 30909
rect 9134 30875 9172 30909
rect 9206 30875 9244 30909
rect 9278 30875 9284 30909
rect 7870 30836 9284 30875
rect 7870 30802 7876 30836
rect 7910 30802 7948 30836
rect 7982 30802 8020 30836
rect 8054 30802 8092 30836
rect 8126 30802 8164 30836
rect 8198 30802 8236 30836
rect 8270 30802 8308 30836
rect 8342 30802 8380 30836
rect 8414 30802 8452 30836
rect 8486 30802 8524 30836
rect 8558 30802 8596 30836
rect 8630 30802 8668 30836
rect 8702 30802 8740 30836
rect 8774 30802 8812 30836
rect 8846 30802 8884 30836
rect 8918 30802 8956 30836
rect 8990 30802 9028 30836
rect 9062 30802 9100 30836
rect 9134 30802 9172 30836
rect 9206 30802 9244 30836
rect 9278 30802 9284 30836
rect 7870 30763 9284 30802
rect 7870 30729 7876 30763
rect 7910 30729 7948 30763
rect 7982 30729 8020 30763
rect 8054 30729 8092 30763
rect 8126 30729 8164 30763
rect 8198 30729 8236 30763
rect 8270 30729 8308 30763
rect 8342 30729 8380 30763
rect 8414 30729 8452 30763
rect 8486 30729 8524 30763
rect 8558 30729 8596 30763
rect 8630 30729 8668 30763
rect 8702 30729 8740 30763
rect 8774 30729 8812 30763
rect 8846 30729 8884 30763
rect 8918 30729 8956 30763
rect 8990 30729 9028 30763
rect 9062 30729 9100 30763
rect 9134 30729 9172 30763
rect 9206 30729 9244 30763
rect 9278 30729 9284 30763
rect 7870 30690 9284 30729
rect 7870 30656 7876 30690
rect 7910 30656 7948 30690
rect 7982 30656 8020 30690
rect 8054 30656 8092 30690
rect 8126 30656 8164 30690
rect 8198 30656 8236 30690
rect 8270 30656 8308 30690
rect 8342 30656 8380 30690
rect 8414 30656 8452 30690
rect 8486 30656 8524 30690
rect 8558 30656 8596 30690
rect 8630 30656 8668 30690
rect 8702 30656 8740 30690
rect 8774 30656 8812 30690
rect 8846 30656 8884 30690
rect 8918 30656 8956 30690
rect 8990 30656 9028 30690
rect 9062 30656 9100 30690
rect 9134 30656 9172 30690
rect 9206 30656 9244 30690
rect 9278 30656 9284 30690
rect 7870 30617 9284 30656
rect 7870 30583 7876 30617
rect 7910 30583 7948 30617
rect 7982 30583 8020 30617
rect 8054 30583 8092 30617
rect 8126 30583 8164 30617
rect 8198 30583 8236 30617
rect 8270 30583 8308 30617
rect 8342 30583 8380 30617
rect 8414 30583 8452 30617
rect 8486 30583 8524 30617
rect 8558 30583 8596 30617
rect 8630 30583 8668 30617
rect 8702 30583 8740 30617
rect 8774 30583 8812 30617
rect 8846 30583 8884 30617
rect 8918 30583 8956 30617
rect 8990 30583 9028 30617
rect 9062 30583 9100 30617
rect 9134 30583 9172 30617
rect 9206 30583 9244 30617
rect 9278 30583 9284 30617
rect 7870 30544 9284 30583
rect 7870 30510 7876 30544
rect 7910 30510 7948 30544
rect 7982 30510 8020 30544
rect 8054 30510 8092 30544
rect 8126 30510 8164 30544
rect 8198 30510 8236 30544
rect 8270 30510 8308 30544
rect 8342 30510 8380 30544
rect 8414 30510 8452 30544
rect 8486 30510 8524 30544
rect 8558 30510 8596 30544
rect 8630 30510 8668 30544
rect 8702 30510 8740 30544
rect 8774 30510 8812 30544
rect 8846 30510 8884 30544
rect 8918 30510 8956 30544
rect 8990 30510 9028 30544
rect 9062 30510 9100 30544
rect 9134 30510 9172 30544
rect 9206 30510 9244 30544
rect 9278 30510 9284 30544
rect 7870 30471 9284 30510
rect 7870 30437 7876 30471
rect 7910 30437 7948 30471
rect 7982 30437 8020 30471
rect 8054 30437 8092 30471
rect 8126 30437 8164 30471
rect 8198 30437 8236 30471
rect 8270 30437 8308 30471
rect 8342 30437 8380 30471
rect 8414 30437 8452 30471
rect 8486 30437 8524 30471
rect 8558 30437 8596 30471
rect 8630 30437 8668 30471
rect 8702 30437 8740 30471
rect 8774 30437 8812 30471
rect 8846 30437 8884 30471
rect 8918 30437 8956 30471
rect 8990 30437 9028 30471
rect 9062 30437 9100 30471
rect 9134 30437 9172 30471
rect 9206 30437 9244 30471
rect 9278 30437 9284 30471
rect 7870 30398 9284 30437
rect 7870 30364 7876 30398
rect 7910 30364 7948 30398
rect 7982 30364 8020 30398
rect 8054 30364 8092 30398
rect 8126 30364 8164 30398
rect 8198 30364 8236 30398
rect 8270 30364 8308 30398
rect 8342 30364 8380 30398
rect 8414 30364 8452 30398
rect 8486 30364 8524 30398
rect 8558 30364 8596 30398
rect 8630 30364 8668 30398
rect 8702 30364 8740 30398
rect 8774 30364 8812 30398
rect 8846 30364 8884 30398
rect 8918 30364 8956 30398
rect 8990 30364 9028 30398
rect 9062 30364 9100 30398
rect 9134 30364 9172 30398
rect 9206 30364 9244 30398
rect 9278 30364 9284 30398
rect 7870 30325 9284 30364
rect 7870 30291 7876 30325
rect 7910 30291 7948 30325
rect 7982 30291 8020 30325
rect 8054 30291 8092 30325
rect 8126 30291 8164 30325
rect 8198 30291 8236 30325
rect 8270 30291 8308 30325
rect 8342 30291 8380 30325
rect 8414 30291 8452 30325
rect 8486 30291 8524 30325
rect 8558 30291 8596 30325
rect 8630 30291 8668 30325
rect 8702 30291 8740 30325
rect 8774 30291 8812 30325
rect 8846 30291 8884 30325
rect 8918 30291 8956 30325
rect 8990 30291 9028 30325
rect 9062 30291 9100 30325
rect 9134 30291 9172 30325
rect 9206 30291 9244 30325
rect 9278 30291 9284 30325
rect 7870 30252 9284 30291
rect 7870 30218 7876 30252
rect 7910 30218 7948 30252
rect 7982 30218 8020 30252
rect 8054 30218 8092 30252
rect 8126 30218 8164 30252
rect 8198 30218 8236 30252
rect 8270 30218 8308 30252
rect 8342 30218 8380 30252
rect 8414 30218 8452 30252
rect 8486 30218 8524 30252
rect 8558 30218 8596 30252
rect 8630 30218 8668 30252
rect 8702 30218 8740 30252
rect 8774 30218 8812 30252
rect 8846 30218 8884 30252
rect 8918 30218 8956 30252
rect 8990 30218 9028 30252
rect 9062 30218 9100 30252
rect 9134 30218 9172 30252
rect 9206 30218 9244 30252
rect 9278 30218 9284 30252
rect 7870 30179 9284 30218
rect 7870 30145 7876 30179
rect 7910 30145 7948 30179
rect 7982 30145 8020 30179
rect 8054 30145 8092 30179
rect 8126 30145 8164 30179
rect 8198 30145 8236 30179
rect 8270 30145 8308 30179
rect 8342 30145 8380 30179
rect 8414 30145 8452 30179
rect 8486 30145 8524 30179
rect 8558 30145 8596 30179
rect 8630 30145 8668 30179
rect 8702 30145 8740 30179
rect 8774 30145 8812 30179
rect 8846 30145 8884 30179
rect 8918 30145 8956 30179
rect 8990 30145 9028 30179
rect 9062 30145 9100 30179
rect 9134 30145 9172 30179
rect 9206 30145 9244 30179
rect 9278 30145 9284 30179
rect 7870 30106 9284 30145
rect 7870 30072 7876 30106
rect 7910 30072 7948 30106
rect 7982 30072 8020 30106
rect 8054 30072 8092 30106
rect 8126 30072 8164 30106
rect 8198 30072 8236 30106
rect 8270 30072 8308 30106
rect 8342 30072 8380 30106
rect 8414 30072 8452 30106
rect 8486 30072 8524 30106
rect 8558 30072 8596 30106
rect 8630 30072 8668 30106
rect 8702 30072 8740 30106
rect 8774 30072 8812 30106
rect 8846 30072 8884 30106
rect 8918 30072 8956 30106
rect 8990 30072 9028 30106
rect 9062 30072 9100 30106
rect 9134 30072 9172 30106
rect 9206 30072 9244 30106
rect 9278 30072 9284 30106
rect 7870 30033 9284 30072
rect 7870 29999 7876 30033
rect 7910 29999 7948 30033
rect 7982 29999 8020 30033
rect 8054 29999 8092 30033
rect 8126 29999 8164 30033
rect 8198 29999 8236 30033
rect 8270 29999 8308 30033
rect 8342 29999 8380 30033
rect 8414 29999 8452 30033
rect 8486 29999 8524 30033
rect 8558 29999 8596 30033
rect 8630 29999 8668 30033
rect 8702 29999 8740 30033
rect 8774 29999 8812 30033
rect 8846 29999 8884 30033
rect 8918 29999 8956 30033
rect 8990 29999 9028 30033
rect 9062 29999 9100 30033
rect 9134 29999 9172 30033
rect 9206 29999 9244 30033
rect 9278 29999 9284 30033
rect 7870 29960 9284 29999
rect 7870 29926 7876 29960
rect 7910 29926 7948 29960
rect 7982 29926 8020 29960
rect 8054 29926 8092 29960
rect 8126 29926 8164 29960
rect 8198 29926 8236 29960
rect 8270 29926 8308 29960
rect 8342 29926 8380 29960
rect 8414 29926 8452 29960
rect 8486 29926 8524 29960
rect 8558 29926 8596 29960
rect 8630 29926 8668 29960
rect 8702 29926 8740 29960
rect 8774 29926 8812 29960
rect 8846 29926 8884 29960
rect 8918 29926 8956 29960
rect 8990 29926 9028 29960
rect 9062 29926 9100 29960
rect 9134 29926 9172 29960
rect 9206 29926 9244 29960
rect 9278 29926 9284 29960
rect 7870 29887 9284 29926
rect 7870 29853 7876 29887
rect 7910 29853 7948 29887
rect 7982 29853 8020 29887
rect 8054 29853 8092 29887
rect 8126 29853 8164 29887
rect 8198 29853 8236 29887
rect 8270 29853 8308 29887
rect 8342 29853 8380 29887
rect 8414 29853 8452 29887
rect 8486 29853 8524 29887
rect 8558 29853 8596 29887
rect 8630 29853 8668 29887
rect 8702 29853 8740 29887
rect 8774 29853 8812 29887
rect 8846 29853 8884 29887
rect 8918 29853 8956 29887
rect 8990 29853 9028 29887
rect 9062 29853 9100 29887
rect 9134 29853 9172 29887
rect 9206 29853 9244 29887
rect 9278 29853 9284 29887
rect 7870 29814 9284 29853
rect 7870 29780 7876 29814
rect 7910 29780 7948 29814
rect 7982 29780 8020 29814
rect 8054 29780 8092 29814
rect 8126 29780 8164 29814
rect 8198 29780 8236 29814
rect 8270 29780 8308 29814
rect 8342 29780 8380 29814
rect 8414 29780 8452 29814
rect 8486 29780 8524 29814
rect 8558 29780 8596 29814
rect 8630 29780 8668 29814
rect 8702 29780 8740 29814
rect 8774 29780 8812 29814
rect 8846 29780 8884 29814
rect 8918 29780 8956 29814
rect 8990 29780 9028 29814
rect 9062 29780 9100 29814
rect 9134 29780 9172 29814
rect 9206 29780 9244 29814
rect 9278 29780 9284 29814
rect 7870 29741 9284 29780
rect 7870 29707 7876 29741
rect 7910 29707 7948 29741
rect 7982 29707 8020 29741
rect 8054 29707 8092 29741
rect 8126 29707 8164 29741
rect 8198 29707 8236 29741
rect 8270 29707 8308 29741
rect 8342 29707 8380 29741
rect 8414 29707 8452 29741
rect 8486 29707 8524 29741
rect 8558 29707 8596 29741
rect 8630 29707 8668 29741
rect 8702 29707 8740 29741
rect 8774 29707 8812 29741
rect 8846 29707 8884 29741
rect 8918 29707 8956 29741
rect 8990 29707 9028 29741
rect 9062 29707 9100 29741
rect 9134 29707 9172 29741
rect 9206 29707 9244 29741
rect 9278 29707 9284 29741
rect 7870 29668 9284 29707
rect 7870 29634 7876 29668
rect 7910 29634 7948 29668
rect 7982 29634 8020 29668
rect 8054 29634 8092 29668
rect 8126 29634 8164 29668
rect 8198 29634 8236 29668
rect 8270 29634 8308 29668
rect 8342 29634 8380 29668
rect 8414 29634 8452 29668
rect 8486 29634 8524 29668
rect 8558 29634 8596 29668
rect 8630 29634 8668 29668
rect 8702 29634 8740 29668
rect 8774 29634 8812 29668
rect 8846 29634 8884 29668
rect 8918 29634 8956 29668
rect 8990 29634 9028 29668
rect 9062 29634 9100 29668
rect 9134 29634 9172 29668
rect 9206 29634 9244 29668
rect 9278 29634 9284 29668
rect 7870 29602 9284 29634
rect 315 29511 1233 29602
tri 1233 29511 1324 29602 nw
tri 8275 29511 8366 29602 ne
rect 8366 29511 9284 29602
rect 315 9241 321 29511
rect 1003 29403 1125 29511
tri 1125 29403 1233 29511 nw
tri 8366 29403 8474 29511 ne
rect 8474 29403 8596 29511
rect 1003 29351 1073 29403
tri 1073 29351 1125 29403 nw
tri 1385 29351 1437 29403 se
rect 1437 29351 3808 29403
rect 3860 29351 3872 29403
rect 3924 29351 3930 29403
rect 5220 29351 5226 29403
rect 5278 29351 5290 29403
rect 5342 29351 7974 29403
tri 7974 29351 8026 29403 sw
tri 8474 29351 8526 29403 ne
rect 8526 29351 8596 29403
rect 1003 29319 1041 29351
tri 1041 29319 1073 29351 nw
tri 1363 29329 1385 29351 se
rect 1385 29329 1437 29351
tri 1437 29329 1459 29351 nw
tri 7952 29332 7971 29351 ne
rect 7971 29332 8026 29351
tri 8026 29332 8045 29351 sw
tri 8526 29332 8545 29351 ne
rect 8545 29332 8596 29351
tri 7971 29329 7974 29332 ne
rect 7974 29329 8045 29332
tri 8045 29329 8048 29332 sw
tri 8545 29329 8548 29332 ne
rect 8548 29329 8596 29332
tri 1353 29319 1363 29329 se
rect 1363 29319 1427 29329
tri 1427 29319 1437 29329 nw
tri 7974 29319 7984 29329 ne
rect 7984 29319 8048 29329
tri 8048 29319 8058 29329 sw
tri 8548 29319 8558 29329 ne
rect 8558 29319 8596 29329
rect 315 9175 321 9189
rect 315 9109 321 9123
rect 315 9043 321 9057
rect 315 8977 321 8991
rect 315 8911 321 8925
rect 315 8844 321 8859
rect 315 8777 321 8792
rect 315 8710 321 8725
rect 315 8643 321 8658
rect 315 8576 321 8591
rect 315 8509 321 8524
rect 315 8442 321 8457
rect 315 8375 321 8390
rect 315 3125 321 8323
rect 1003 3125 1009 29319
tri 1009 29287 1041 29319 nw
tri 1321 29287 1353 29319 se
rect 1353 29291 1399 29319
tri 1399 29291 1427 29319 nw
tri 1445 29291 1473 29319 se
rect 1473 29291 3938 29319
rect 1353 29287 1375 29291
tri 1301 29267 1321 29287 se
rect 1321 29267 1375 29287
tri 1375 29267 1399 29291 nw
tri 1421 29267 1445 29291 se
rect 1445 29267 3938 29291
rect 3990 29267 4002 29319
rect 4054 29267 4060 29319
rect 5319 29267 5325 29319
rect 5377 29267 5389 29319
rect 5441 29296 7938 29319
tri 7938 29296 7961 29319 sw
tri 7984 29296 8007 29319 ne
rect 8007 29296 8058 29319
tri 8058 29296 8081 29319 sw
tri 8558 29296 8581 29319 ne
rect 8581 29296 8596 29319
rect 5441 29287 7961 29296
tri 7961 29287 7970 29296 sw
tri 8007 29287 8016 29296 ne
rect 8016 29287 8081 29296
tri 8081 29287 8090 29296 sw
tri 8581 29287 8590 29296 ne
rect 5441 29283 7970 29287
tri 7970 29283 7974 29287 sw
tri 8016 29283 8020 29287 ne
rect 8020 29283 8090 29287
rect 5441 29267 7974 29283
tri 7974 29267 7990 29283 sw
tri 8020 29267 8036 29283 ne
rect 8036 29267 8090 29283
tri 8090 29267 8110 29287 sw
tri 1289 29255 1301 29267 se
rect 1301 29255 1363 29267
tri 1363 29255 1375 29267 nw
tri 1409 29255 1421 29267 se
rect 1421 29255 1473 29267
tri 1269 29235 1289 29255 se
rect 1289 29245 1353 29255
tri 1353 29245 1363 29255 nw
tri 1399 29245 1409 29255 se
rect 1409 29245 1473 29255
tri 1473 29245 1495 29267 nw
tri 7916 29245 7938 29267 ne
rect 7938 29258 7990 29267
tri 7990 29258 7999 29267 sw
tri 8036 29258 8045 29267 ne
rect 8045 29258 8110 29267
tri 8110 29258 8119 29267 sw
rect 7938 29245 7999 29258
rect 1289 29235 1343 29245
tri 1343 29235 1353 29245 nw
tri 1389 29235 1399 29245 se
rect 1399 29235 1463 29245
tri 1463 29235 1473 29245 nw
tri 7938 29235 7948 29245 ne
rect 7948 29235 7999 29245
tri 7999 29235 8022 29258 sw
tri 8045 29235 8068 29258 ne
rect 8068 29235 8119 29258
tri 8119 29235 8142 29258 sw
tri 1217 29183 1269 29235 se
rect 1269 29217 1325 29235
tri 1325 29217 1343 29235 nw
tri 1371 29217 1389 29235 se
rect 1389 29217 1427 29235
rect 1269 29183 1291 29217
tri 1291 29183 1325 29217 nw
tri 1337 29183 1371 29217 se
rect 1371 29199 1427 29217
tri 1427 29199 1463 29235 nw
tri 1473 29199 1509 29235 se
rect 1509 29199 4045 29235
rect 1371 29183 1411 29199
tri 1411 29183 1427 29199 nw
tri 1457 29183 1473 29199 se
rect 1473 29183 4045 29199
rect 4097 29183 4109 29235
rect 4161 29183 4167 29235
rect 5425 29183 5431 29235
rect 5483 29183 5495 29235
rect 5547 29232 7902 29235
tri 7902 29232 7905 29235 sw
tri 7948 29232 7951 29235 ne
rect 7951 29232 8022 29235
rect 5547 29222 7905 29232
tri 7905 29222 7915 29232 sw
tri 7951 29222 7961 29232 ne
rect 7961 29222 8022 29232
tri 8022 29222 8035 29235 sw
tri 8068 29222 8081 29235 ne
rect 8081 29222 8142 29235
tri 8142 29222 8155 29235 sw
rect 5547 29186 7915 29222
tri 7915 29186 7951 29222 sw
tri 7961 29186 7997 29222 ne
rect 7997 29212 8035 29222
tri 8035 29212 8045 29222 sw
tri 8081 29212 8091 29222 ne
rect 8091 29212 8155 29222
rect 7997 29186 8045 29212
rect 5547 29183 7951 29186
tri 7951 29183 7954 29186 sw
tri 7997 29183 8000 29186 ne
rect 8000 29184 8045 29186
tri 8045 29184 8073 29212 sw
tri 8091 29184 8119 29212 ne
rect 8119 29184 8155 29212
tri 8155 29184 8193 29222 sw
rect 8000 29183 8073 29184
tri 8073 29183 8074 29184 sw
tri 8119 29183 8120 29184 ne
rect 8120 29183 8193 29184
tri 8193 29183 8194 29184 sw
tri 1215 29181 1217 29183 se
rect 1217 29181 1289 29183
tri 1289 29181 1291 29183 nw
tri 1335 29181 1337 29183 se
rect 1337 29181 1409 29183
tri 1409 29181 1411 29183 nw
tri 1455 29181 1457 29183 se
rect 1457 29181 1509 29183
tri 1185 29151 1215 29181 se
rect 1215 29171 1279 29181
tri 1279 29171 1289 29181 nw
tri 1325 29171 1335 29181 se
rect 1335 29171 1399 29181
tri 1399 29171 1409 29181 nw
tri 1445 29171 1455 29181 se
rect 1455 29171 1509 29181
rect 1215 29151 1259 29171
tri 1259 29151 1279 29171 nw
tri 1315 29161 1325 29171 se
rect 1325 29161 1389 29171
tri 1389 29161 1399 29171 nw
tri 1435 29161 1445 29171 se
rect 1445 29161 1509 29171
tri 1509 29161 1531 29183 nw
tri 7880 29161 7902 29183 ne
rect 7902 29161 7954 29183
tri 7954 29161 7976 29183 sw
tri 8000 29161 8022 29183 ne
rect 8022 29161 8074 29183
tri 1305 29151 1315 29161 se
rect 1315 29151 1379 29161
tri 1379 29151 1389 29161 nw
tri 1425 29151 1435 29161 se
rect 1435 29151 1499 29161
tri 1499 29151 1509 29161 nw
tri 7902 29151 7912 29161 ne
rect 7912 29158 7976 29161
tri 7976 29158 7979 29161 sw
tri 8022 29158 8025 29161 ne
rect 8025 29158 8074 29161
rect 7912 29151 7979 29158
tri 7979 29151 7986 29158 sw
tri 8025 29151 8032 29158 ne
rect 8032 29151 8074 29158
tri 8074 29151 8106 29183 sw
tri 8120 29151 8152 29183 ne
rect 8152 29151 8194 29183
tri 8194 29151 8226 29183 sw
tri 1144 29110 1185 29151 se
rect 1185 29143 1251 29151
tri 1251 29143 1259 29151 nw
tri 1297 29143 1305 29151 se
rect 1305 29143 1353 29151
rect 1185 29110 1218 29143
tri 1218 29110 1251 29143 nw
tri 1264 29110 1297 29143 se
rect 1297 29125 1353 29143
tri 1353 29125 1379 29151 nw
tri 1399 29125 1425 29151 se
rect 1425 29125 1463 29151
rect 1297 29110 1338 29125
tri 1338 29110 1353 29125 nw
tri 1384 29110 1399 29125 se
rect 1399 29115 1463 29125
tri 1463 29115 1499 29151 nw
tri 1509 29115 1545 29151 se
rect 1545 29115 4151 29151
rect 1399 29110 1447 29115
rect 1144 29099 1207 29110
tri 1207 29099 1218 29110 nw
tri 1253 29099 1264 29110 se
rect 1264 29099 1327 29110
tri 1327 29099 1338 29110 nw
tri 1373 29099 1384 29110 se
rect 1384 29099 1447 29110
tri 1447 29099 1463 29115 nw
tri 1493 29099 1509 29115 se
rect 1509 29099 4151 29115
rect 4203 29099 4215 29151
rect 4267 29099 4273 29151
rect 5532 29099 5538 29151
rect 5590 29099 5602 29151
rect 5654 29150 7866 29151
tri 7866 29150 7867 29151 sw
tri 7912 29150 7913 29151 ne
rect 7913 29150 7986 29151
tri 7986 29150 7987 29151 sw
tri 8032 29150 8033 29151 ne
rect 8033 29150 8106 29151
tri 8106 29150 8107 29151 sw
tri 8152 29150 8153 29151 ne
rect 8153 29150 8226 29151
tri 8226 29150 8227 29151 sw
rect 5654 29137 7867 29150
tri 7867 29137 7880 29150 sw
tri 7913 29137 7926 29150 ne
rect 7926 29148 7987 29150
tri 7987 29148 7989 29150 sw
tri 8033 29148 8035 29150 ne
rect 8035 29148 8107 29150
tri 8107 29148 8109 29150 sw
tri 8153 29148 8155 29150 ne
rect 8155 29148 8227 29150
tri 8227 29148 8229 29150 sw
rect 7926 29137 7989 29148
rect 5654 29112 7880 29137
tri 7880 29112 7905 29137 sw
tri 7926 29112 7951 29137 ne
rect 7951 29112 7989 29137
tri 7989 29112 8025 29148 sw
tri 8035 29112 8071 29148 ne
rect 8071 29138 8109 29148
tri 8109 29138 8119 29148 sw
tri 8155 29138 8165 29148 ne
rect 8165 29138 8229 29148
rect 8071 29112 8119 29138
rect 5654 29099 7905 29112
tri 7905 29099 7918 29112 sw
tri 7951 29099 7964 29112 ne
rect 7964 29099 8025 29112
tri 8025 29099 8038 29112 sw
tri 8071 29099 8084 29112 ne
rect 8084 29110 8119 29112
tri 8119 29110 8147 29138 sw
tri 8165 29110 8193 29138 ne
rect 8193 29110 8229 29138
tri 8229 29110 8267 29148 sw
rect 8084 29099 8147 29110
tri 8147 29099 8158 29110 sw
tri 8193 29099 8204 29110 ne
rect 8204 29099 8267 29110
rect 1144 7572 1196 29099
tri 1196 29088 1207 29099 nw
tri 1251 29097 1253 29099 se
rect 1253 29097 1325 29099
tri 1325 29097 1327 29099 nw
tri 1371 29097 1373 29099 se
rect 1373 29097 1435 29099
tri 1242 29088 1251 29097 se
rect 1251 29088 1316 29097
tri 1316 29088 1325 29097 nw
tri 1362 29088 1371 29097 se
rect 1371 29088 1435 29097
tri 1241 29087 1242 29088 se
rect 1242 29087 1315 29088
tri 1315 29087 1316 29088 nw
tri 1361 29087 1362 29088 se
rect 1362 29087 1435 29088
tri 1435 29087 1447 29099 nw
tri 1481 29087 1493 29099 se
rect 1493 29087 1545 29099
tri 1231 29077 1241 29087 se
rect 1241 29077 1305 29087
tri 1305 29077 1315 29087 nw
tri 1351 29077 1361 29087 se
rect 1361 29077 1425 29087
tri 1425 29077 1435 29087 nw
tri 1471 29077 1481 29087 se
rect 1481 29077 1545 29087
tri 1545 29077 1567 29099 nw
tri 7844 29077 7866 29099 ne
rect 7866 29077 7918 29099
tri 7918 29077 7940 29099 sw
tri 7964 29077 7986 29099 ne
rect 7986 29084 8038 29099
tri 8038 29084 8053 29099 sw
tri 8084 29084 8099 29099 ne
rect 8099 29084 8158 29099
rect 7986 29077 8053 29084
tri 8053 29077 8060 29084 sw
tri 8099 29077 8106 29084 ne
rect 8106 29077 8158 29084
tri 8158 29077 8180 29099 sw
tri 8204 29088 8215 29099 ne
rect 1144 7508 1196 7520
rect 1144 7450 1196 7456
tri 1228 29074 1231 29077 se
rect 1231 29074 1302 29077
tri 1302 29074 1305 29077 nw
tri 1348 29074 1351 29077 se
rect 1351 29074 1415 29077
rect 1228 29067 1295 29074
tri 1295 29067 1302 29074 nw
tri 1341 29067 1348 29074 se
rect 1348 29067 1415 29074
tri 1415 29067 1425 29077 nw
tri 1461 29067 1471 29077 se
rect 1471 29067 1535 29077
tri 1535 29067 1545 29077 nw
tri 7866 29076 7867 29077 ne
rect 7867 29076 7940 29077
tri 7940 29076 7941 29077 sw
tri 7986 29076 7987 29077 ne
rect 7987 29076 8060 29077
tri 8060 29076 8061 29077 sw
tri 8106 29076 8107 29077 ne
rect 8107 29076 8180 29077
tri 8180 29076 8181 29077 sw
tri 7867 29067 7876 29076 ne
rect 7876 29067 7941 29076
tri 7941 29067 7950 29076 sw
tri 7987 29067 7996 29076 ne
rect 7996 29074 8061 29076
tri 8061 29074 8063 29076 sw
tri 8107 29074 8109 29076 ne
rect 8109 29074 8181 29076
tri 8181 29074 8183 29076 sw
rect 7996 29067 8063 29074
tri 8063 29067 8070 29074 sw
tri 8109 29067 8116 29074 ne
rect 8116 29067 8183 29074
rect 1228 6750 1280 29067
tri 1280 29052 1295 29067 nw
tri 1326 29052 1341 29067 se
rect 1341 29052 1389 29067
tri 1312 29038 1326 29052 se
rect 1326 29041 1389 29052
tri 1389 29041 1415 29067 nw
tri 1435 29041 1461 29067 se
rect 1461 29041 1507 29067
rect 1326 29038 1386 29041
tri 1386 29038 1389 29041 nw
tri 1432 29038 1435 29041 se
rect 1435 29039 1507 29041
tri 1507 29039 1535 29067 nw
tri 1553 29039 1581 29067 se
rect 1581 29039 4250 29067
rect 1435 29038 1483 29039
rect 1312 10688 1364 29038
tri 1364 29016 1386 29038 nw
tri 1410 29016 1432 29038 se
rect 1432 29016 1483 29038
tri 1409 29015 1410 29016 se
rect 1410 29015 1483 29016
tri 1483 29015 1507 29039 nw
tri 1529 29015 1553 29039 se
rect 1553 29015 4250 29039
rect 4302 29015 4314 29067
rect 4366 29015 4372 29067
rect 5662 29015 5668 29067
rect 5720 29015 5732 29067
rect 5784 29040 7830 29067
tri 7830 29040 7857 29067 sw
tri 7876 29040 7903 29067 ne
rect 7903 29066 7950 29067
tri 7950 29066 7951 29067 sw
tri 7996 29066 7997 29067 ne
rect 7997 29066 8070 29067
rect 7903 29040 7951 29066
rect 5784 29015 7857 29040
tri 7857 29015 7882 29040 sw
tri 7903 29015 7928 29040 ne
rect 7928 29038 7951 29040
tri 7951 29038 7979 29066 sw
tri 7997 29038 8025 29066 ne
rect 8025 29052 8070 29066
tri 8070 29052 8085 29067 sw
tri 8116 29052 8131 29067 ne
rect 8025 29038 8085 29052
tri 8085 29038 8099 29052 sw
rect 7928 29015 7979 29038
tri 7979 29015 8002 29038 sw
tri 8025 29016 8047 29038 ne
tri 1397 29003 1409 29015 se
rect 1409 29003 1471 29015
tri 1471 29003 1483 29015 nw
tri 1517 29003 1529 29015 se
rect 1529 29003 1591 29015
tri 1591 29003 1603 29015 nw
tri 7808 29003 7820 29015 ne
rect 7820 29012 7882 29015
tri 7882 29012 7885 29015 sw
tri 7928 29012 7931 29015 ne
rect 7931 29012 8002 29015
rect 7820 29003 7885 29012
tri 7885 29003 7894 29012 sw
tri 7931 29003 7940 29012 ne
rect 7940 29003 8002 29012
tri 8002 29003 8014 29015 sw
rect 1312 10624 1364 10636
rect 1312 10566 1364 10572
tri 1396 29002 1397 29003 se
rect 1397 29002 1470 29003
tri 1470 29002 1471 29003 nw
tri 1516 29002 1517 29003 se
rect 1517 29002 1590 29003
tri 1590 29002 1591 29003 nw
tri 7820 29002 7821 29003 ne
rect 7821 29002 7894 29003
tri 7894 29002 7895 29003 sw
tri 7940 29002 7941 29003 ne
rect 7941 29002 8014 29003
tri 8014 29002 8015 29003 sw
rect 1228 6686 1280 6698
rect 1228 6628 1280 6634
rect 1312 10249 1364 10255
rect 1312 10185 1364 10197
rect 315 3086 1009 3125
rect 315 3052 321 3086
rect 355 3052 393 3086
rect 427 3052 465 3086
rect 499 3052 537 3086
rect 571 3052 609 3086
rect 643 3052 681 3086
rect 715 3052 753 3086
rect 787 3052 825 3086
rect 859 3052 897 3086
rect 931 3052 969 3086
rect 1003 3052 1009 3086
rect 315 3013 1009 3052
rect 315 2979 321 3013
rect 355 2979 393 3013
rect 427 2979 465 3013
rect 499 2979 537 3013
rect 571 2979 609 3013
rect 643 2979 681 3013
rect 715 2979 753 3013
rect 787 2979 825 3013
rect 859 2979 897 3013
rect 931 2979 969 3013
rect 1003 2979 1009 3013
rect 315 2940 1009 2979
rect 315 2906 321 2940
rect 355 2906 393 2940
rect 427 2906 465 2940
rect 499 2906 537 2940
rect 571 2906 609 2940
rect 643 2906 681 2940
rect 715 2906 753 2940
rect 787 2906 825 2940
rect 859 2906 897 2940
rect 931 2906 969 2940
rect 1003 2906 1009 2940
rect 315 2867 1009 2906
rect 315 2833 321 2867
rect 355 2833 393 2867
rect 427 2833 465 2867
rect 499 2833 537 2867
rect 571 2833 609 2867
rect 643 2833 681 2867
rect 715 2833 753 2867
rect 787 2833 825 2867
rect 859 2833 897 2867
rect 931 2833 969 2867
rect 1003 2833 1009 2867
rect 315 2794 1009 2833
rect 315 2760 321 2794
rect 355 2760 393 2794
rect 427 2760 465 2794
rect 499 2760 537 2794
rect 571 2760 609 2794
rect 643 2760 681 2794
rect 715 2760 753 2794
rect 787 2760 825 2794
rect 859 2760 897 2794
rect 931 2760 969 2794
rect 1003 2760 1009 2794
rect 315 2721 1009 2760
rect 315 2687 321 2721
rect 355 2687 393 2721
rect 427 2687 465 2721
rect 499 2687 537 2721
rect 571 2687 609 2721
rect 643 2687 681 2721
rect 715 2687 753 2721
rect 787 2687 825 2721
rect 859 2687 897 2721
rect 931 2687 969 2721
rect 1003 2687 1009 2721
rect 315 2648 1009 2687
rect 315 2614 321 2648
rect 355 2614 393 2648
rect 427 2614 465 2648
rect 499 2614 537 2648
rect 571 2614 609 2648
rect 643 2614 681 2648
rect 715 2614 753 2648
rect 787 2614 825 2648
rect 859 2614 897 2648
rect 931 2614 969 2648
rect 1003 2614 1009 2648
rect 315 2575 1009 2614
rect 315 2541 321 2575
rect 355 2541 393 2575
rect 427 2541 465 2575
rect 499 2541 537 2575
rect 571 2541 609 2575
rect 643 2541 681 2575
rect 715 2541 753 2575
rect 787 2541 825 2575
rect 859 2541 897 2575
rect 931 2541 969 2575
rect 1003 2541 1009 2575
rect 315 2502 1009 2541
rect 315 2468 321 2502
rect 355 2468 393 2502
rect 427 2468 465 2502
rect 499 2468 537 2502
rect 571 2468 609 2502
rect 643 2468 681 2502
rect 715 2468 753 2502
rect 787 2468 825 2502
rect 859 2468 897 2502
rect 931 2468 969 2502
rect 1003 2468 1009 2502
rect 315 2429 1009 2468
rect 315 2395 321 2429
rect 355 2395 393 2429
rect 427 2395 465 2429
rect 499 2395 537 2429
rect 571 2395 609 2429
rect 643 2395 681 2429
rect 715 2395 753 2429
rect 787 2395 825 2429
rect 859 2395 897 2429
rect 931 2395 969 2429
rect 1003 2395 1009 2429
rect 315 2356 1009 2395
rect 315 2322 321 2356
rect 355 2322 393 2356
rect 427 2322 465 2356
rect 499 2322 537 2356
rect 571 2322 609 2356
rect 643 2322 681 2356
rect 715 2322 753 2356
rect 787 2322 825 2356
rect 859 2322 897 2356
rect 931 2322 969 2356
rect 1003 2322 1009 2356
rect 315 2283 1009 2322
rect 315 2249 321 2283
rect 355 2249 393 2283
rect 427 2249 465 2283
rect 499 2249 537 2283
rect 571 2249 609 2283
rect 643 2249 681 2283
rect 715 2249 753 2283
rect 787 2249 825 2283
rect 859 2249 897 2283
rect 931 2249 969 2283
rect 1003 2249 1009 2283
rect 315 2210 1009 2249
rect 315 2176 321 2210
rect 355 2176 393 2210
rect 427 2176 465 2210
rect 499 2176 537 2210
rect 571 2176 609 2210
rect 643 2176 681 2210
rect 715 2176 753 2210
rect 787 2176 825 2210
rect 859 2176 897 2210
rect 931 2176 969 2210
rect 1003 2176 1009 2210
rect 315 2137 1009 2176
rect 315 2103 321 2137
rect 355 2103 393 2137
rect 427 2103 465 2137
rect 499 2103 537 2137
rect 571 2103 609 2137
rect 643 2103 681 2137
rect 715 2103 753 2137
rect 787 2103 825 2137
rect 859 2103 897 2137
rect 931 2103 969 2137
rect 1003 2103 1009 2137
rect 315 2064 1009 2103
rect 315 2030 321 2064
rect 355 2030 393 2064
rect 427 2030 465 2064
rect 499 2030 537 2064
rect 571 2030 609 2064
rect 643 2030 681 2064
rect 715 2030 753 2064
rect 787 2030 825 2064
rect 859 2030 897 2064
rect 931 2030 969 2064
rect 1003 2030 1009 2064
rect 315 1991 1009 2030
rect 315 1957 321 1991
rect 355 1957 393 1991
rect 427 1957 465 1991
rect 499 1957 537 1991
rect 571 1957 609 1991
rect 643 1957 681 1991
rect 715 1957 753 1991
rect 787 1957 825 1991
rect 859 1957 897 1991
rect 931 1957 969 1991
rect 1003 1957 1009 1991
rect 315 1918 1009 1957
rect 315 1884 321 1918
rect 355 1884 393 1918
rect 427 1884 465 1918
rect 499 1884 537 1918
rect 571 1884 609 1918
rect 643 1884 681 1918
rect 715 1884 753 1918
rect 787 1884 825 1918
rect 859 1884 897 1918
rect 931 1884 969 1918
rect 1003 1884 1009 1918
rect 315 1845 1009 1884
rect 315 1811 321 1845
rect 355 1811 393 1845
rect 427 1811 465 1845
rect 499 1811 537 1845
rect 571 1811 609 1845
rect 643 1811 681 1845
rect 715 1811 753 1845
rect 787 1811 825 1845
rect 859 1811 897 1845
rect 931 1811 969 1845
rect 1003 1811 1009 1845
rect 315 1772 1009 1811
rect 315 1738 321 1772
rect 355 1738 393 1772
rect 427 1738 465 1772
rect 499 1738 537 1772
rect 571 1738 609 1772
rect 643 1738 681 1772
rect 715 1738 753 1772
rect 787 1738 825 1772
rect 859 1738 897 1772
rect 931 1738 969 1772
rect 1003 1738 1009 1772
rect 315 1699 1009 1738
rect 315 1665 321 1699
rect 355 1665 393 1699
rect 427 1665 465 1699
rect 499 1665 537 1699
rect 571 1665 609 1699
rect 643 1665 681 1699
rect 715 1665 753 1699
rect 787 1665 825 1699
rect 859 1665 897 1699
rect 931 1665 969 1699
rect 1003 1665 1009 1699
rect 315 1626 1009 1665
rect 315 1592 321 1626
rect 355 1592 393 1626
rect 427 1592 465 1626
rect 499 1592 537 1626
rect 571 1592 609 1626
rect 643 1592 681 1626
rect 715 1592 753 1626
rect 787 1592 825 1626
rect 859 1592 897 1626
rect 931 1592 969 1626
rect 1003 1592 1009 1626
rect 315 1553 1009 1592
rect 315 1519 321 1553
rect 355 1519 393 1553
rect 427 1519 465 1553
rect 499 1519 537 1553
rect 571 1519 609 1553
rect 643 1519 681 1553
rect 715 1519 753 1553
rect 787 1519 825 1553
rect 859 1519 897 1553
rect 931 1519 969 1553
rect 1003 1519 1009 1553
rect 315 1480 1009 1519
rect 315 1446 321 1480
rect 355 1446 393 1480
rect 427 1446 465 1480
rect 499 1446 537 1480
rect 571 1446 609 1480
rect 643 1446 681 1480
rect 715 1446 753 1480
rect 787 1446 825 1480
rect 859 1446 897 1480
rect 931 1446 969 1480
rect 1003 1446 1009 1480
rect 315 1407 1009 1446
rect 315 1373 321 1407
rect 355 1373 393 1407
rect 427 1373 465 1407
rect 499 1373 537 1407
rect 571 1373 609 1407
rect 643 1373 681 1407
rect 715 1373 753 1407
rect 787 1373 825 1407
rect 859 1373 897 1407
rect 931 1373 969 1407
rect 1003 1373 1009 1407
rect 315 1334 1009 1373
rect 315 1300 321 1334
rect 355 1300 393 1334
rect 427 1300 465 1334
rect 499 1300 537 1334
rect 571 1300 609 1334
rect 643 1300 681 1334
rect 715 1300 753 1334
rect 787 1300 825 1334
rect 859 1300 897 1334
rect 931 1300 969 1334
rect 1003 1300 1009 1334
rect 315 1261 1009 1300
rect 315 1227 321 1261
rect 355 1227 393 1261
rect 427 1227 465 1261
rect 499 1227 537 1261
rect 571 1227 609 1261
rect 643 1227 681 1261
rect 715 1227 753 1261
rect 787 1227 825 1261
rect 859 1227 897 1261
rect 931 1227 969 1261
rect 1003 1227 1009 1261
rect 315 1188 1009 1227
rect 315 1154 321 1188
rect 355 1154 393 1188
rect 427 1154 465 1188
rect 499 1154 537 1188
rect 571 1154 609 1188
rect 643 1154 681 1188
rect 715 1154 753 1188
rect 787 1154 825 1188
rect 859 1154 897 1188
rect 931 1154 969 1188
rect 1003 1154 1009 1188
rect 315 1115 1009 1154
rect 315 1081 321 1115
rect 355 1081 393 1115
rect 427 1081 465 1115
rect 499 1081 537 1115
rect 571 1081 609 1115
rect 643 1081 681 1115
rect 715 1081 753 1115
rect 787 1081 825 1115
rect 859 1081 897 1115
rect 931 1081 969 1115
rect 1003 1081 1009 1115
rect 315 1042 1009 1081
rect 315 1008 321 1042
rect 355 1008 393 1042
rect 427 1008 465 1042
rect 499 1008 537 1042
rect 571 1008 609 1042
rect 643 1008 681 1042
rect 715 1008 753 1042
rect 787 1008 825 1042
rect 859 1008 897 1042
rect 931 1008 969 1042
rect 1003 1008 1009 1042
rect 315 969 1009 1008
rect 315 935 321 969
rect 355 935 393 969
rect 427 935 465 969
rect 499 935 537 969
rect 571 935 609 969
rect 643 935 681 969
rect 715 935 753 969
rect 787 935 825 969
rect 859 935 897 969
rect 931 935 969 969
rect 1003 935 1009 969
rect 315 896 1009 935
rect 315 862 321 896
rect 355 862 393 896
rect 427 862 465 896
rect 499 862 537 896
rect 571 862 609 896
rect 643 862 681 896
rect 715 862 753 896
rect 787 862 825 896
rect 859 862 897 896
rect 931 862 969 896
rect 1003 862 1009 896
rect 315 823 1009 862
rect 315 789 321 823
rect 355 789 393 823
rect 427 789 465 823
rect 499 789 537 823
rect 571 789 609 823
rect 643 789 681 823
rect 715 789 753 823
rect 787 789 825 823
rect 859 789 897 823
rect 931 789 969 823
rect 1003 789 1009 823
rect 315 750 1009 789
rect 315 716 321 750
rect 355 716 393 750
rect 427 716 465 750
rect 499 716 537 750
rect 571 716 609 750
rect 643 716 681 750
rect 715 716 753 750
rect 787 716 825 750
rect 859 716 897 750
rect 931 716 969 750
rect 1003 716 1009 750
rect 315 677 1009 716
rect 315 643 321 677
rect 355 643 393 677
rect 427 643 465 677
rect 499 643 537 677
rect 571 643 609 677
rect 643 643 681 677
rect 715 643 753 677
rect 787 643 825 677
rect 859 643 897 677
rect 931 643 969 677
rect 1003 643 1009 677
rect 315 604 1009 643
rect 315 570 321 604
rect 355 570 393 604
rect 427 570 465 604
rect 499 570 537 604
rect 571 570 609 604
rect 643 570 681 604
rect 715 570 753 604
rect 787 570 825 604
rect 859 570 897 604
rect 931 570 969 604
rect 1003 570 1009 604
rect 315 531 1009 570
rect 315 497 321 531
rect 355 497 393 531
rect 427 497 465 531
rect 499 497 537 531
rect 571 497 609 531
rect 643 497 681 531
rect 715 497 753 531
rect 787 497 825 531
rect 859 497 897 531
rect 931 497 969 531
rect 1003 497 1009 531
rect 315 458 1009 497
rect 315 424 321 458
rect 355 424 393 458
rect 427 424 465 458
rect 499 424 537 458
rect 571 424 609 458
rect 643 424 681 458
rect 715 424 753 458
rect 787 424 825 458
rect 859 424 897 458
rect 931 424 969 458
rect 1003 424 1009 458
rect 315 385 1009 424
rect 315 351 321 385
rect 355 351 393 385
rect 427 351 465 385
rect 499 351 537 385
rect 571 351 609 385
rect 643 351 681 385
rect 715 351 753 385
rect 787 351 825 385
rect 859 351 897 385
rect 931 351 969 385
rect 1003 351 1009 385
rect 315 312 1009 351
rect 315 278 321 312
rect 355 278 393 312
rect 427 278 465 312
rect 499 278 537 312
rect 571 278 609 312
rect 643 278 681 312
rect 715 278 753 312
rect 787 278 825 312
rect 859 278 897 312
rect 931 278 969 312
rect 1003 278 1009 312
rect 315 239 1009 278
rect 315 205 321 239
rect 355 205 393 239
rect 427 205 465 239
rect 499 205 537 239
rect 571 205 609 239
rect 643 205 681 239
rect 715 205 753 239
rect 787 205 825 239
rect 859 205 897 239
rect 931 205 969 239
rect 1003 205 1009 239
rect 315 166 1009 205
rect 315 132 321 166
rect 355 132 393 166
rect 427 132 465 166
rect 499 132 537 166
rect 571 132 609 166
rect 643 132 681 166
rect 715 132 753 166
rect 787 132 825 166
rect 859 132 897 166
rect 931 132 969 166
rect 1003 132 1009 166
rect 315 93 1009 132
rect 315 59 321 93
rect 355 59 393 93
rect 427 59 465 93
rect 499 59 537 93
rect 571 59 609 93
rect 643 59 681 93
rect 715 59 753 93
rect 787 59 825 93
rect 859 59 897 93
rect 931 59 969 93
rect 1003 59 1009 93
rect 315 27 1009 59
rect 1312 122 1364 10133
rect 1396 3958 1448 29002
tri 1448 28980 1470 29002 nw
tri 1507 28993 1516 29002 se
rect 1516 28993 1581 29002
tri 1581 28993 1590 29002 nw
tri 7821 28993 7830 29002 ne
rect 7830 28993 7895 29002
tri 1494 28980 1507 28993 se
rect 1507 28980 1568 28993
tri 1568 28980 1581 28993 nw
tri 7830 28980 7843 28993 ne
rect 7843 28980 7895 28993
tri 7895 28980 7917 29002 sw
tri 7941 28980 7963 29002 ne
tri 1480 28966 1494 28980 se
rect 1494 28966 1554 28980
tri 1554 28966 1568 28980 nw
tri 7843 28966 7857 28980 ne
rect 7857 28966 7917 28980
tri 7917 28966 7931 28980 sw
rect 1480 9790 1532 28966
tri 1532 28944 1554 28966 nw
tri 7857 28944 7879 28966 ne
rect 4627 22783 5045 22789
rect 4679 22731 5045 22783
rect 4627 22693 5045 22731
rect 4679 22641 5045 22693
rect 4627 22603 5045 22641
rect 4679 22551 5045 22603
rect 4627 22545 5045 22551
rect 4998 18602 5004 18654
rect 5056 18602 5072 18654
rect 5124 18602 5140 18654
rect 5192 18602 5198 18654
rect 4998 18588 5198 18602
rect 4998 18536 5004 18588
rect 5056 18536 5072 18588
rect 5124 18536 5140 18588
rect 5192 18536 5198 18588
tri 7869 18395 7879 18405 se
rect 7879 18395 7931 28966
tri 7843 18369 7869 18395 se
rect 7869 18383 7931 18395
rect 7869 18369 7917 18383
tri 7917 18369 7931 18383 nw
tri 7835 18361 7843 18369 se
rect 7843 18361 7909 18369
tri 7909 18361 7917 18369 nw
tri 7955 18361 7963 18369 se
rect 7963 18361 8015 29002
tri 7805 18331 7835 18361 se
rect 7835 18337 7885 18361
tri 7885 18337 7909 18361 nw
tri 7931 18337 7955 18361 se
rect 7955 18347 8015 18361
rect 7955 18337 8001 18347
rect 7835 18331 7879 18337
tri 7879 18331 7885 18337 nw
tri 7925 18331 7931 18337 se
rect 7931 18333 8001 18337
tri 8001 18333 8015 18347 nw
rect 7931 18331 7990 18333
tri 7796 18322 7805 18331 se
rect 7805 18322 7870 18331
tri 7870 18322 7879 18331 nw
tri 7916 18322 7925 18331 se
rect 7925 18322 7990 18331
tri 7990 18322 8001 18333 nw
tri 8036 18322 8047 18333 se
rect 8047 18322 8099 29038
tri 7769 18295 7796 18322 se
rect 7796 18295 7843 18322
tri 7843 18295 7870 18322 nw
tri 7889 18295 7916 18322 se
rect 7916 18305 7973 18322
tri 7973 18305 7990 18322 nw
tri 8019 18305 8036 18322 se
rect 8036 18311 8099 18322
rect 8036 18305 8085 18311
rect 7916 18295 7963 18305
tri 7963 18295 7973 18305 nw
tri 8011 18297 8019 18305 se
rect 8019 18297 8085 18305
tri 8085 18297 8099 18311 nw
tri 8009 18295 8011 18297 se
rect 8011 18295 8083 18297
tri 8083 18295 8085 18297 nw
tri 8129 18295 8131 18297 se
rect 8131 18295 8183 29067
tri 7762 18288 7769 18295 se
rect 7769 18288 7836 18295
tri 7836 18288 7843 18295 nw
tri 7882 18288 7889 18295 se
rect 7889 18288 7956 18295
tri 7956 18288 7963 18295 nw
tri 8002 18288 8009 18295 se
rect 8009 18288 8076 18295
tri 8076 18288 8083 18295 nw
tri 8122 18288 8129 18295 se
rect 8129 18288 8183 18295
tri 7731 18257 7762 18288 se
rect 7762 18285 7833 18288
tri 7833 18285 7836 18288 nw
tri 7879 18285 7882 18288 se
rect 7882 18285 7927 18288
rect 7762 18257 7805 18285
tri 7805 18257 7833 18285 nw
tri 7851 18257 7879 18285 se
rect 7879 18259 7927 18285
tri 7927 18259 7956 18288 nw
tri 7973 18259 8002 18288 se
rect 8002 18265 8053 18288
tri 8053 18265 8076 18288 nw
tri 8099 18265 8122 18288 se
rect 8122 18275 8183 18288
rect 8122 18265 8169 18275
rect 8002 18259 8047 18265
tri 8047 18259 8053 18265 nw
tri 8093 18259 8099 18265 se
rect 8099 18261 8169 18265
tri 8169 18261 8183 18275 nw
rect 8099 18259 8157 18261
rect 7879 18257 7917 18259
tri 7723 18249 7731 18257 se
rect 7731 18249 7797 18257
tri 7797 18249 7805 18257 nw
tri 7843 18249 7851 18257 se
rect 7851 18249 7917 18257
tri 7917 18249 7927 18259 nw
tri 7963 18249 7973 18259 se
rect 7973 18249 8037 18259
tri 8037 18249 8047 18259 nw
tri 8083 18249 8093 18259 se
rect 8093 18249 8157 18259
tri 8157 18249 8169 18261 nw
tri 8203 18249 8215 18261 se
rect 8215 18249 8267 29099
tri 7695 18221 7723 18249 se
rect 7723 18221 7769 18249
tri 7769 18221 7797 18249 nw
tri 7815 18221 7843 18249 se
rect 7843 18231 7899 18249
tri 7899 18231 7917 18249 nw
tri 7945 18231 7963 18249 se
rect 7963 18231 8011 18249
rect 7843 18221 7889 18231
tri 7889 18221 7899 18231 nw
tri 7937 18223 7945 18231 se
rect 7945 18223 8011 18231
tri 8011 18223 8037 18249 nw
tri 8057 18223 8083 18249 se
rect 8083 18233 8141 18249
tri 8141 18233 8157 18249 nw
tri 8187 18233 8203 18249 se
rect 8203 18239 8267 18249
rect 8203 18233 8243 18239
rect 8083 18223 8131 18233
tri 8131 18223 8141 18233 nw
tri 8177 18223 8187 18233 se
rect 8187 18223 8243 18233
tri 7935 18221 7937 18223 se
rect 7937 18221 8009 18223
tri 8009 18221 8011 18223 nw
tri 8055 18221 8057 18223 se
rect 8057 18221 8123 18223
tri 7689 18215 7695 18221 se
rect 7695 18215 7763 18221
tri 7763 18215 7769 18221 nw
tri 7809 18215 7815 18221 se
rect 7815 18215 7883 18221
tri 7883 18215 7889 18221 nw
tri 7929 18215 7935 18221 se
rect 7935 18215 8003 18221
tri 8003 18215 8009 18221 nw
tri 8049 18215 8055 18221 se
rect 8055 18215 8123 18221
tri 8123 18215 8131 18223 nw
tri 8169 18215 8177 18223 se
rect 8177 18215 8243 18223
tri 8243 18215 8267 18239 nw
rect 8590 20405 8596 29296
rect 9278 20405 9284 29511
rect 8590 20366 9284 20405
rect 8590 20332 8596 20366
rect 8630 20332 8668 20366
rect 8702 20332 8740 20366
rect 8774 20332 8812 20366
rect 8846 20332 8884 20366
rect 8918 20332 8956 20366
rect 8990 20332 9028 20366
rect 9062 20332 9100 20366
rect 9134 20332 9172 20366
rect 9206 20332 9244 20366
rect 9278 20332 9284 20366
rect 8590 20293 9284 20332
rect 8590 20259 8596 20293
rect 8630 20259 8668 20293
rect 8702 20259 8740 20293
rect 8774 20259 8812 20293
rect 8846 20259 8884 20293
rect 8918 20259 8956 20293
rect 8990 20259 9028 20293
rect 9062 20259 9100 20293
rect 9134 20259 9172 20293
rect 9206 20259 9244 20293
rect 9278 20259 9284 20293
rect 8590 20220 9284 20259
rect 8590 20186 8596 20220
rect 8630 20186 8668 20220
rect 8702 20186 8740 20220
rect 8774 20186 8812 20220
rect 8846 20186 8884 20220
rect 8918 20186 8956 20220
rect 8990 20186 9028 20220
rect 9062 20186 9100 20220
rect 9134 20186 9172 20220
rect 9206 20186 9244 20220
rect 9278 20186 9284 20220
rect 8590 20147 9284 20186
rect 8590 20113 8596 20147
rect 8630 20113 8668 20147
rect 8702 20113 8740 20147
rect 8774 20113 8812 20147
rect 8846 20113 8884 20147
rect 8918 20113 8956 20147
rect 8990 20113 9028 20147
rect 9062 20113 9100 20147
rect 9134 20113 9172 20147
rect 9206 20113 9244 20147
rect 9278 20113 9284 20147
rect 8590 20074 9284 20113
rect 8590 20040 8596 20074
rect 8630 20040 8668 20074
rect 8702 20040 8740 20074
rect 8774 20040 8812 20074
rect 8846 20040 8884 20074
rect 8918 20040 8956 20074
rect 8990 20040 9028 20074
rect 9062 20040 9100 20074
rect 9134 20040 9172 20074
rect 9206 20040 9244 20074
rect 9278 20040 9284 20074
rect 8590 20001 9284 20040
rect 8590 19967 8596 20001
rect 8630 19967 8668 20001
rect 8702 19967 8740 20001
rect 8774 19967 8812 20001
rect 8846 19967 8884 20001
rect 8918 19967 8956 20001
rect 8990 19967 9028 20001
rect 9062 19967 9100 20001
rect 9134 19967 9172 20001
rect 9206 19967 9244 20001
rect 9278 19967 9284 20001
rect 8590 19928 9284 19967
rect 8590 19894 8596 19928
rect 8630 19894 8668 19928
rect 8702 19894 8740 19928
rect 8774 19894 8812 19928
rect 8846 19894 8884 19928
rect 8918 19894 8956 19928
rect 8990 19894 9028 19928
rect 9062 19894 9100 19928
rect 9134 19894 9172 19928
rect 9206 19894 9244 19928
rect 9278 19894 9284 19928
rect 8590 19855 9284 19894
rect 8590 19821 8596 19855
rect 8630 19821 8668 19855
rect 8702 19821 8740 19855
rect 8774 19821 8812 19855
rect 8846 19821 8884 19855
rect 8918 19821 8956 19855
rect 8990 19821 9028 19855
rect 9062 19821 9100 19855
rect 9134 19821 9172 19855
rect 9206 19821 9244 19855
rect 9278 19821 9284 19855
rect 8590 19782 9284 19821
rect 8590 19748 8596 19782
rect 8630 19748 8668 19782
rect 8702 19748 8740 19782
rect 8774 19748 8812 19782
rect 8846 19748 8884 19782
rect 8918 19748 8956 19782
rect 8990 19748 9028 19782
rect 9062 19748 9100 19782
rect 9134 19748 9172 19782
rect 9206 19748 9244 19782
rect 9278 19748 9284 19782
rect 8590 19709 9284 19748
rect 8590 19675 8596 19709
rect 8630 19675 8668 19709
rect 8702 19675 8740 19709
rect 8774 19675 8812 19709
rect 8846 19675 8884 19709
rect 8918 19675 8956 19709
rect 8990 19675 9028 19709
rect 9062 19675 9100 19709
rect 9134 19675 9172 19709
rect 9206 19675 9244 19709
rect 9278 19675 9284 19709
rect 8590 19636 9284 19675
rect 8590 19602 8596 19636
rect 8630 19602 8668 19636
rect 8702 19602 8740 19636
rect 8774 19602 8812 19636
rect 8846 19602 8884 19636
rect 8918 19602 8956 19636
rect 8990 19602 9028 19636
rect 9062 19602 9100 19636
rect 9134 19602 9172 19636
rect 9206 19602 9244 19636
rect 9278 19602 9284 19636
rect 8590 19563 9284 19602
rect 8590 19529 8596 19563
rect 8630 19529 8668 19563
rect 8702 19529 8740 19563
rect 8774 19529 8812 19563
rect 8846 19529 8884 19563
rect 8918 19529 8956 19563
rect 8990 19529 9028 19563
rect 9062 19529 9100 19563
rect 9134 19529 9172 19563
rect 9206 19529 9244 19563
rect 9278 19529 9284 19563
rect 8590 19490 9284 19529
rect 8590 19456 8596 19490
rect 8630 19456 8668 19490
rect 8702 19456 8740 19490
rect 8774 19456 8812 19490
rect 8846 19456 8884 19490
rect 8918 19456 8956 19490
rect 8990 19456 9028 19490
rect 9062 19456 9100 19490
rect 9134 19456 9172 19490
rect 9206 19456 9244 19490
rect 9278 19456 9284 19490
rect 8590 19417 9284 19456
rect 8590 19383 8596 19417
rect 8630 19383 8668 19417
rect 8702 19383 8740 19417
rect 8774 19383 8812 19417
rect 8846 19383 8884 19417
rect 8918 19383 8956 19417
rect 8990 19383 9028 19417
rect 9062 19383 9100 19417
rect 9134 19383 9172 19417
rect 9206 19383 9244 19417
rect 9278 19383 9284 19417
rect 8590 19344 9284 19383
rect 8590 19310 8596 19344
rect 8630 19310 8668 19344
rect 8702 19310 8740 19344
rect 8774 19310 8812 19344
rect 8846 19310 8884 19344
rect 8918 19310 8956 19344
rect 8990 19310 9028 19344
rect 9062 19310 9100 19344
rect 9134 19310 9172 19344
rect 9206 19310 9244 19344
rect 9278 19310 9284 19344
rect 8590 19271 9284 19310
rect 8590 19237 8596 19271
rect 8630 19237 8668 19271
rect 8702 19237 8740 19271
rect 8774 19237 8812 19271
rect 8846 19237 8884 19271
rect 8918 19237 8956 19271
rect 8990 19237 9028 19271
rect 9062 19237 9100 19271
rect 9134 19237 9172 19271
rect 9206 19237 9244 19271
rect 9278 19237 9284 19271
rect 8590 19198 9284 19237
rect 8590 19164 8596 19198
rect 8630 19164 8668 19198
rect 8702 19164 8740 19198
rect 8774 19164 8812 19198
rect 8846 19164 8884 19198
rect 8918 19164 8956 19198
rect 8990 19164 9028 19198
rect 9062 19164 9100 19198
rect 9134 19164 9172 19198
rect 9206 19164 9244 19198
rect 9278 19164 9284 19198
rect 8590 19125 9284 19164
rect 8590 19091 8596 19125
rect 8630 19091 8668 19125
rect 8702 19091 8740 19125
rect 8774 19091 8812 19125
rect 8846 19091 8884 19125
rect 8918 19091 8956 19125
rect 8990 19091 9028 19125
rect 9062 19091 9100 19125
rect 9134 19091 9172 19125
rect 9206 19091 9244 19125
rect 9278 19091 9284 19125
rect 8590 19052 9284 19091
rect 8590 19018 8596 19052
rect 8630 19018 8668 19052
rect 8702 19018 8740 19052
rect 8774 19018 8812 19052
rect 8846 19018 8884 19052
rect 8918 19018 8956 19052
rect 8990 19018 9028 19052
rect 9062 19018 9100 19052
rect 9134 19018 9172 19052
rect 9206 19018 9244 19052
rect 9278 19018 9284 19052
rect 8590 18979 9284 19018
rect 8590 18945 8596 18979
rect 8630 18945 8668 18979
rect 8702 18945 8740 18979
rect 8774 18945 8812 18979
rect 8846 18945 8884 18979
rect 8918 18945 8956 18979
rect 8990 18945 9028 18979
rect 9062 18945 9100 18979
rect 9134 18945 9172 18979
rect 9206 18945 9244 18979
rect 9278 18945 9284 18979
rect 8590 18906 9284 18945
rect 8590 18872 8596 18906
rect 8630 18872 8668 18906
rect 8702 18872 8740 18906
rect 8774 18872 8812 18906
rect 8846 18872 8884 18906
rect 8918 18872 8956 18906
rect 8990 18872 9028 18906
rect 9062 18872 9100 18906
rect 9134 18872 9172 18906
rect 9206 18872 9244 18906
rect 9278 18872 9284 18906
rect 8590 18833 9284 18872
rect 8590 18799 8596 18833
rect 8630 18799 8668 18833
rect 8702 18799 8740 18833
rect 8774 18799 8812 18833
rect 8846 18799 8884 18833
rect 8918 18799 8956 18833
rect 8990 18799 9028 18833
rect 9062 18799 9100 18833
rect 9134 18799 9172 18833
rect 9206 18799 9244 18833
rect 9278 18799 9284 18833
rect 8590 18760 9284 18799
rect 8590 18726 8596 18760
rect 8630 18726 8668 18760
rect 8702 18726 8740 18760
rect 8774 18726 8812 18760
rect 8846 18726 8884 18760
rect 8918 18726 8956 18760
rect 8990 18726 9028 18760
rect 9062 18726 9100 18760
rect 9134 18726 9172 18760
rect 9206 18726 9244 18760
rect 9278 18726 9284 18760
rect 8590 18687 9284 18726
rect 8590 18653 8596 18687
rect 8630 18653 8668 18687
rect 8702 18653 8740 18687
rect 8774 18653 8812 18687
rect 8846 18653 8884 18687
rect 8918 18653 8956 18687
rect 8990 18653 9028 18687
rect 9062 18653 9100 18687
rect 9134 18653 9172 18687
rect 9206 18653 9244 18687
rect 9278 18653 9284 18687
rect 8590 18614 9284 18653
rect 8590 18580 8596 18614
rect 8630 18580 8668 18614
rect 8702 18580 8740 18614
rect 8774 18580 8812 18614
rect 8846 18580 8884 18614
rect 8918 18580 8956 18614
rect 8990 18580 9028 18614
rect 9062 18580 9100 18614
rect 9134 18580 9172 18614
rect 9206 18580 9244 18614
rect 9278 18580 9284 18614
rect 8590 18541 9284 18580
rect 8590 18507 8596 18541
rect 8630 18507 8668 18541
rect 8702 18507 8740 18541
rect 8774 18507 8812 18541
rect 8846 18507 8884 18541
rect 8918 18507 8956 18541
rect 8990 18507 9028 18541
rect 9062 18507 9100 18541
rect 9134 18507 9172 18541
rect 9206 18507 9244 18541
rect 9278 18507 9284 18541
rect 8590 18468 9284 18507
rect 8590 18434 8596 18468
rect 8630 18434 8668 18468
rect 8702 18434 8740 18468
rect 8774 18434 8812 18468
rect 8846 18434 8884 18468
rect 8918 18434 8956 18468
rect 8990 18434 9028 18468
rect 9062 18434 9100 18468
rect 9134 18434 9172 18468
rect 9206 18434 9244 18468
rect 9278 18434 9284 18468
rect 8590 18395 9284 18434
rect 8590 18361 8596 18395
rect 8630 18361 8668 18395
rect 8702 18361 8740 18395
rect 8774 18361 8812 18395
rect 8846 18361 8884 18395
rect 8918 18361 8956 18395
rect 8990 18361 9028 18395
rect 9062 18361 9100 18395
rect 9134 18361 9172 18395
rect 9206 18361 9244 18395
rect 9278 18361 9284 18395
rect 8590 18322 9284 18361
rect 8590 18288 8596 18322
rect 8630 18288 8668 18322
rect 8702 18288 8740 18322
rect 8774 18288 8812 18322
rect 8846 18288 8884 18322
rect 8918 18288 8956 18322
rect 8990 18288 9028 18322
rect 9062 18288 9100 18322
rect 9134 18288 9172 18322
rect 9206 18288 9244 18322
rect 9278 18288 9284 18322
rect 8590 18249 9284 18288
rect 8590 18215 8596 18249
rect 8630 18215 8668 18249
rect 8702 18215 8740 18249
rect 8774 18215 8812 18249
rect 8846 18215 8884 18249
rect 8918 18215 8956 18249
rect 8990 18215 9028 18249
rect 9062 18215 9100 18249
rect 9134 18215 9172 18249
rect 9206 18215 9244 18249
rect 9278 18215 9284 18249
tri 7680 18206 7689 18215 se
rect 7689 18211 7759 18215
tri 7759 18211 7763 18215 nw
tri 7805 18211 7809 18215 se
rect 7809 18211 7853 18215
rect 7689 18206 7754 18211
tri 7754 18206 7759 18211 nw
tri 7800 18206 7805 18211 se
rect 7805 18206 7853 18211
tri 1900 18176 1930 18206 se
rect 1930 18176 7724 18206
tri 7724 18176 7754 18206 nw
tri 7770 18176 7800 18206 se
rect 7800 18185 7853 18206
tri 7853 18185 7883 18215 nw
tri 7899 18185 7929 18215 se
rect 7929 18213 8001 18215
tri 8001 18213 8003 18215 nw
tri 8047 18213 8049 18215 se
rect 8049 18213 8095 18215
rect 7929 18185 7973 18213
tri 7973 18185 8001 18213 nw
tri 8019 18185 8047 18213 se
rect 8047 18187 8095 18213
tri 8095 18187 8123 18215 nw
tri 8141 18187 8169 18215 se
rect 8169 18187 8215 18215
tri 8215 18187 8243 18215 nw
rect 8047 18185 8084 18187
rect 7800 18176 7844 18185
tri 7844 18176 7853 18185 nw
tri 7890 18176 7899 18185 se
rect 7899 18176 7964 18185
tri 7964 18176 7973 18185 nw
tri 8010 18176 8019 18185 se
rect 8019 18176 8084 18185
tri 8084 18176 8095 18187 nw
tri 8130 18176 8141 18187 se
rect 8141 18176 8204 18187
tri 8204 18176 8215 18187 nw
rect 8590 18176 9284 18215
tri 1871 18147 1900 18176 se
rect 1900 18160 7708 18176
tri 7708 18160 7724 18176 nw
tri 7754 18160 7770 18176 se
rect 7770 18160 7825 18176
rect 1900 18154 7702 18160
tri 7702 18154 7708 18160 nw
tri 7748 18154 7754 18160 se
rect 7754 18157 7825 18160
tri 7825 18157 7844 18176 nw
tri 7871 18157 7890 18176 se
rect 7890 18157 7937 18176
rect 7754 18154 7815 18157
rect 1900 18147 1945 18154
tri 1945 18147 1952 18154 nw
tri 7741 18147 7748 18154 se
rect 7748 18147 7815 18154
tri 7815 18147 7825 18157 nw
tri 7863 18149 7871 18157 se
rect 7871 18149 7937 18157
tri 7937 18149 7964 18176 nw
tri 7983 18149 8010 18176 se
rect 8010 18159 8067 18176
tri 8067 18159 8084 18176 nw
tri 8113 18159 8130 18176 se
rect 8130 18159 8170 18176
rect 8010 18149 8057 18159
tri 8057 18149 8067 18159 nw
tri 8103 18149 8113 18159 se
rect 8113 18149 8170 18159
tri 7861 18147 7863 18149 se
rect 7863 18147 7935 18149
tri 7935 18147 7937 18149 nw
tri 7981 18147 7983 18149 se
rect 7983 18147 8050 18149
tri 1866 18142 1871 18147 se
rect 1871 18142 1940 18147
tri 1940 18142 1945 18147 nw
tri 7736 18142 7741 18147 se
rect 7741 18142 7810 18147
tri 7810 18142 7815 18147 nw
tri 7856 18142 7861 18147 se
rect 7861 18142 7930 18147
tri 7930 18142 7935 18147 nw
tri 7976 18142 7981 18147 se
rect 7981 18142 8050 18147
tri 8050 18142 8057 18149 nw
tri 8096 18142 8103 18149 se
rect 8103 18142 8170 18149
tri 8170 18142 8204 18176 nw
rect 8590 18142 8596 18176
rect 8630 18142 8668 18176
rect 8702 18142 8740 18176
rect 8774 18142 8812 18176
rect 8846 18142 8884 18176
rect 8918 18142 8956 18176
rect 8990 18142 9028 18176
rect 9062 18142 9100 18176
rect 9134 18142 9172 18176
rect 9206 18142 9244 18176
rect 9278 18142 9284 18176
tri 1856 18132 1866 18142 se
rect 1866 18132 1930 18142
tri 1930 18132 1940 18142 nw
tri 7726 18132 7736 18142 se
rect 7736 18132 7790 18142
tri 1846 18122 1856 18132 se
rect 1856 18122 1920 18132
tri 1920 18122 1930 18132 nw
tri 7716 18122 7726 18132 se
rect 7726 18122 7790 18132
tri 7790 18122 7810 18142 nw
tri 7836 18122 7856 18142 se
rect 7856 18139 7927 18142
tri 7927 18139 7930 18142 nw
tri 7973 18139 7976 18142 se
rect 7976 18139 8021 18142
rect 7856 18122 7910 18139
tri 7910 18122 7927 18139 nw
tri 7956 18122 7973 18139 se
rect 7973 18122 8021 18139
tri 1827 18103 1846 18122 se
rect 1846 18103 1901 18122
tri 1901 18103 1920 18122 nw
tri 1947 18103 1966 18122 se
rect 1966 18111 7779 18122
tri 7779 18111 7790 18122 nw
tri 7825 18111 7836 18122 se
rect 7836 18111 7899 18122
tri 7899 18111 7910 18122 nw
tri 7945 18111 7956 18122 se
rect 7956 18113 8021 18122
tri 8021 18113 8050 18142 nw
tri 8067 18113 8096 18142 se
rect 8096 18113 8141 18142
tri 8141 18113 8170 18142 nw
rect 7956 18111 8011 18113
rect 1966 18103 7771 18111
tri 7771 18103 7779 18111 nw
tri 7817 18103 7825 18111 se
rect 7825 18103 7891 18111
tri 7891 18103 7899 18111 nw
tri 7937 18103 7945 18111 se
rect 7945 18103 8011 18111
tri 8011 18103 8021 18113 nw
tri 8057 18103 8067 18113 se
rect 8067 18103 8131 18113
tri 8131 18103 8141 18113 nw
rect 8590 18103 9284 18142
tri 1793 18069 1827 18103 se
rect 1827 18086 1884 18103
tri 1884 18086 1901 18103 nw
tri 1930 18086 1947 18103 se
rect 1947 18086 7752 18103
rect 1827 18069 1867 18086
tri 1867 18069 1884 18086 nw
tri 1913 18069 1930 18086 se
rect 1930 18084 7752 18086
tri 7752 18084 7771 18103 nw
tri 7798 18084 7817 18103 se
rect 7817 18084 7863 18103
rect 1930 18070 7738 18084
tri 7738 18070 7752 18084 nw
tri 7789 18075 7798 18084 se
rect 7798 18075 7863 18084
tri 7863 18075 7891 18103 nw
tri 7909 18075 7937 18103 se
rect 7937 18085 7993 18103
tri 7993 18085 8011 18103 nw
tri 8039 18085 8057 18103 se
rect 8057 18085 8097 18103
rect 7937 18075 7983 18085
tri 7983 18075 7993 18085 nw
tri 8029 18075 8039 18085 se
rect 8039 18075 8097 18085
tri 7784 18070 7789 18075 se
rect 7789 18070 7858 18075
tri 7858 18070 7863 18075 nw
tri 7904 18070 7909 18075 se
rect 7909 18070 7977 18075
rect 1930 18069 1987 18070
tri 1987 18069 1988 18070 nw
tri 7783 18069 7784 18070 se
rect 7784 18069 7857 18070
tri 7857 18069 7858 18070 nw
tri 7903 18069 7904 18070 se
rect 7904 18069 7977 18070
tri 7977 18069 7983 18075 nw
tri 8023 18069 8029 18075 se
rect 8029 18069 8097 18075
tri 8097 18069 8131 18103 nw
rect 8590 18069 8596 18103
rect 8630 18069 8668 18103
rect 8702 18069 8740 18103
rect 8774 18069 8812 18103
rect 8846 18069 8884 18103
rect 8918 18069 8956 18103
rect 8990 18069 9028 18103
rect 9062 18069 9100 18103
rect 9134 18069 9172 18103
rect 9206 18069 9244 18103
rect 9278 18069 9284 18103
tri 1782 18058 1793 18069 se
rect 1793 18058 1856 18069
tri 1856 18058 1867 18069 nw
tri 1902 18058 1913 18069 se
rect 1913 18058 1966 18069
tri 1772 18048 1782 18058 se
rect 1782 18048 1846 18058
tri 1846 18048 1856 18058 nw
tri 1892 18048 1902 18058 se
rect 1902 18048 1966 18058
tri 1966 18048 1987 18069 nw
tri 7762 18048 7783 18069 se
rect 7783 18065 7853 18069
tri 7853 18065 7857 18069 nw
tri 7899 18065 7903 18069 se
rect 7903 18065 7947 18069
rect 7783 18048 7836 18065
tri 7836 18048 7853 18065 nw
tri 7882 18048 7899 18065 se
rect 7899 18048 7947 18065
tri 1754 18030 1772 18048 se
rect 1772 18030 1828 18048
tri 1828 18030 1846 18048 nw
tri 1874 18030 1892 18048 se
rect 1892 18038 1956 18048
tri 1956 18038 1966 18048 nw
tri 7752 18038 7762 18048 se
rect 7762 18038 7826 18048
tri 7826 18038 7836 18048 nw
tri 7872 18038 7882 18048 se
rect 7882 18039 7947 18048
tri 7947 18039 7977 18069 nw
tri 7993 18039 8023 18069 se
rect 8023 18039 8067 18069
tri 8067 18039 8097 18069 nw
rect 7882 18038 7938 18039
rect 1892 18030 1948 18038
tri 1948 18030 1956 18038 nw
tri 1994 18030 2002 18038 se
rect 2002 18030 7818 18038
tri 7818 18030 7826 18038 nw
tri 7864 18030 7872 18038 se
rect 7872 18030 7938 18038
tri 7938 18030 7947 18039 nw
tri 7984 18030 7993 18039 se
rect 7993 18030 8058 18039
tri 8058 18030 8067 18039 nw
rect 8590 18030 9284 18069
tri 1720 17996 1754 18030 se
rect 1754 18012 1810 18030
tri 1810 18012 1828 18030 nw
tri 1856 18012 1874 18030 se
rect 1874 18012 1928 18030
rect 1754 17996 1794 18012
tri 1794 17996 1810 18012 nw
tri 1840 17996 1856 18012 se
rect 1856 18010 1928 18012
tri 1928 18010 1948 18030 nw
tri 1974 18010 1994 18030 se
rect 1994 18010 7789 18030
rect 1856 17996 1914 18010
tri 1914 17996 1928 18010 nw
tri 1965 18001 1974 18010 se
rect 1974 18001 7789 18010
tri 7789 18001 7818 18030 nw
tri 7835 18001 7864 18030 se
rect 7864 18011 7919 18030
tri 7919 18011 7938 18030 nw
tri 7965 18011 7984 18030 se
rect 7984 18011 8024 18030
rect 7864 18001 7909 18011
tri 7909 18001 7919 18011 nw
tri 7955 18001 7965 18011 se
rect 7965 18001 8024 18011
tri 1960 17996 1965 18001 se
rect 1965 17996 7784 18001
tri 7784 17996 7789 18001 nw
tri 7830 17996 7835 18001 se
rect 7835 17996 7904 18001
tri 7904 17996 7909 18001 nw
tri 7950 17996 7955 18001 se
rect 7955 17996 8024 18001
tri 8024 17996 8058 18030 nw
rect 8590 17996 8596 18030
rect 8630 17996 8668 18030
rect 8702 17996 8740 18030
rect 8774 17996 8812 18030
rect 8846 17996 8884 18030
rect 8918 17996 8956 18030
rect 8990 17996 9028 18030
rect 9062 17996 9100 18030
rect 9134 17996 9172 18030
rect 9206 17996 9244 18030
rect 9278 17996 9284 18030
tri 1708 17984 1720 17996 se
rect 1720 17984 1782 17996
tri 1782 17984 1794 17996 nw
tri 1828 17984 1840 17996 se
rect 1840 17984 1892 17996
tri 1698 17974 1708 17984 se
rect 1708 17974 1772 17984
tri 1772 17974 1782 17984 nw
tri 1818 17974 1828 17984 se
rect 1828 17974 1892 17984
tri 1892 17974 1914 17996 nw
tri 1938 17974 1960 17996 se
rect 1960 17992 7780 17996
tri 7780 17992 7784 17996 nw
tri 7826 17992 7830 17996 se
rect 7830 17992 7873 17996
rect 1960 17986 7774 17992
tri 7774 17986 7780 17992 nw
tri 7820 17986 7826 17992 se
rect 7826 17986 7873 17992
rect 1960 17974 2012 17986
tri 2012 17974 2024 17986 nw
tri 7808 17974 7820 17986 se
rect 7820 17974 7873 17986
tri 1681 17957 1698 17974 se
rect 1698 17957 1755 17974
tri 1755 17957 1772 17974 nw
tri 1801 17957 1818 17974 se
rect 1818 17964 1882 17974
tri 1882 17964 1892 17974 nw
tri 1928 17964 1938 17974 se
rect 1938 17964 2002 17974
tri 2002 17964 2012 17974 nw
tri 7798 17964 7808 17974 se
rect 7808 17965 7873 17974
tri 7873 17965 7904 17996 nw
tri 7919 17965 7950 17996 se
rect 7950 17965 7993 17996
tri 7993 17965 8024 17996 nw
rect 7808 17964 7865 17965
rect 1818 17957 1875 17964
tri 1875 17957 1882 17964 nw
tri 1921 17957 1928 17964 se
rect 1928 17957 1995 17964
tri 1995 17957 2002 17964 nw
tri 7791 17957 7798 17964 se
rect 7798 17957 7865 17964
tri 7865 17957 7873 17965 nw
tri 7911 17957 7919 17965 se
rect 7919 17957 7985 17965
tri 7985 17957 7993 17965 nw
rect 8590 17957 9284 17996
tri 1647 17923 1681 17957 se
rect 1681 17938 1736 17957
tri 1736 17938 1755 17957 nw
tri 1782 17938 1801 17957 se
rect 1801 17938 1854 17957
rect 1681 17923 1721 17938
tri 1721 17923 1736 17938 nw
tri 1767 17923 1782 17938 se
rect 1782 17936 1854 17938
tri 1854 17936 1875 17957 nw
tri 1918 17954 1921 17957 se
rect 1921 17954 1992 17957
tri 1992 17954 1995 17957 nw
tri 7788 17954 7791 17957 se
rect 7791 17954 7862 17957
tri 7862 17954 7865 17957 nw
tri 7908 17954 7911 17957 se
rect 7911 17954 7951 17957
tri 1900 17936 1918 17954 se
rect 1918 17936 1961 17954
rect 1782 17923 1841 17936
tri 1841 17923 1854 17936 nw
tri 1887 17923 1900 17936 se
rect 1900 17923 1961 17936
tri 1961 17923 1992 17954 nw
tri 2007 17923 2038 17954 se
rect 2038 17937 7845 17954
tri 7845 17937 7862 17954 nw
tri 7891 17937 7908 17954 se
rect 7908 17937 7951 17954
rect 2038 17923 7831 17937
tri 7831 17923 7845 17937 nw
tri 7877 17923 7891 17937 se
rect 7891 17923 7951 17937
tri 7951 17923 7985 17957 nw
rect 8590 17923 8596 17957
rect 8630 17923 8668 17957
rect 8702 17923 8740 17957
rect 8774 17923 8812 17957
rect 8846 17923 8884 17957
rect 8918 17923 8956 17957
rect 8990 17923 9028 17957
rect 9062 17923 9100 17957
rect 9134 17923 9172 17957
rect 9206 17923 9244 17957
rect 9278 17923 9284 17957
tri 1634 17910 1647 17923 se
rect 1647 17910 1708 17923
tri 1708 17910 1721 17923 nw
tri 1754 17910 1767 17923 se
rect 1767 17910 1818 17923
tri 1624 17900 1634 17910 se
rect 1634 17900 1698 17910
tri 1698 17900 1708 17910 nw
tri 1744 17900 1754 17910 se
rect 1754 17900 1818 17910
tri 1818 17900 1841 17923 nw
tri 1864 17900 1887 17923 se
rect 1887 17918 1956 17923
tri 1956 17918 1961 17923 nw
tri 2002 17918 2007 17923 se
rect 2007 17918 7810 17923
rect 1887 17900 1938 17918
tri 1938 17900 1956 17918 nw
tri 1984 17900 2002 17918 se
rect 2002 17902 7810 17918
tri 7810 17902 7831 17923 nw
tri 7856 17902 7877 17923 se
rect 7877 17902 7924 17923
rect 2002 17900 2054 17902
tri 1608 17884 1624 17900 se
rect 1624 17884 1682 17900
tri 1682 17884 1698 17900 nw
tri 1728 17884 1744 17900 se
rect 1744 17890 1808 17900
tri 1808 17890 1818 17900 nw
tri 1860 17896 1864 17900 se
rect 1864 17896 1934 17900
tri 1934 17896 1938 17900 nw
tri 1980 17896 1984 17900 se
rect 1984 17896 2054 17900
tri 2054 17896 2060 17902 nw
tri 7850 17896 7856 17902 se
rect 7856 17896 7924 17902
tri 7924 17896 7951 17923 nw
tri 1854 17890 1860 17896 se
rect 1860 17890 1928 17896
tri 1928 17890 1934 17896 nw
tri 1974 17890 1980 17896 se
rect 1980 17890 2042 17896
rect 1744 17884 1802 17890
tri 1802 17884 1808 17890 nw
tri 1848 17884 1854 17890 se
rect 1854 17884 1922 17890
tri 1922 17884 1928 17890 nw
tri 1968 17884 1974 17890 se
rect 1974 17884 2042 17890
tri 2042 17884 2054 17896 nw
tri 7845 17891 7850 17896 se
rect 7850 17891 7919 17896
tri 7919 17891 7924 17896 nw
tri 8585 17891 8590 17896 se
rect 8590 17891 9284 17923
tri 7838 17884 7845 17891 se
rect 7845 17884 7912 17891
tri 7912 17884 7919 17891 nw
tri 8578 17884 8585 17891 se
rect 8585 17884 9284 17891
tri 1574 17850 1608 17884 se
rect 1608 17864 1662 17884
tri 1662 17864 1682 17884 nw
tri 1708 17864 1728 17884 se
rect 1728 17864 1780 17884
rect 1608 17850 1648 17864
tri 1648 17850 1662 17864 nw
tri 1694 17850 1708 17864 se
rect 1708 17862 1780 17864
tri 1780 17862 1802 17884 nw
tri 1844 17880 1848 17884 se
rect 1848 17880 1918 17884
tri 1918 17880 1922 17884 nw
tri 1964 17880 1968 17884 se
rect 1968 17880 2038 17884
tri 2038 17880 2042 17884 nw
tri 7834 17880 7838 17884 se
rect 7838 17880 7898 17884
tri 1826 17862 1844 17880 se
rect 1844 17862 1888 17880
rect 1708 17850 1768 17862
tri 1768 17850 1780 17862 nw
tri 1814 17850 1826 17862 se
rect 1826 17850 1888 17862
tri 1888 17850 1918 17880 nw
tri 1934 17850 1964 17880 se
rect 1964 17870 2028 17880
tri 2028 17870 2038 17880 nw
tri 7824 17870 7834 17880 se
rect 7834 17870 7898 17880
tri 7898 17870 7912 17884 nw
tri 8564 17870 8578 17884 se
rect 8578 17870 8596 17884
rect 1964 17850 2008 17870
tri 2008 17850 2028 17870 nw
tri 2054 17850 2074 17870 se
rect 2074 17850 7878 17870
tri 7878 17850 7898 17870 nw
tri 8544 17850 8564 17870 se
rect 8564 17850 8596 17870
rect 8630 17850 8668 17884
rect 8702 17850 8740 17884
rect 8774 17850 8812 17884
rect 8846 17850 8884 17884
rect 8918 17850 8956 17884
rect 8990 17850 9028 17884
rect 9062 17850 9100 17884
rect 9134 17850 9172 17884
rect 9206 17850 9244 17884
rect 9278 17850 9284 17884
tri 1564 17840 1574 17850 se
rect 1574 17840 1638 17850
tri 1638 17840 1648 17850 nw
tri 1684 17840 1694 17850 se
rect 1694 17840 1744 17850
rect 1564 17826 1624 17840
tri 1624 17826 1638 17840 nw
tri 1670 17826 1684 17840 se
rect 1684 17826 1744 17840
tri 1744 17826 1768 17850 nw
tri 1790 17826 1814 17850 se
rect 1814 17844 1882 17850
tri 1882 17844 1888 17850 nw
tri 1928 17844 1934 17850 se
rect 1934 17844 2000 17850
rect 1814 17826 1864 17844
tri 1864 17826 1882 17844 nw
tri 1910 17826 1928 17844 se
rect 1928 17842 2000 17844
tri 2000 17842 2008 17850 nw
tri 2046 17842 2054 17850 se
rect 2054 17842 7854 17850
rect 1928 17826 1984 17842
tri 1984 17826 2000 17842 nw
tri 2030 17826 2046 17842 se
rect 2046 17826 7854 17842
tri 7854 17826 7878 17850 nw
tri 8520 17826 8544 17850 se
rect 8544 17826 9284 17850
rect 1564 14838 1616 17826
tri 1616 17818 1624 17826 nw
tri 1662 17818 1670 17826 se
rect 1670 17818 1734 17826
tri 1655 17811 1662 17818 se
rect 1662 17816 1734 17818
tri 1734 17816 1744 17826 nw
tri 1780 17816 1790 17826 se
rect 1790 17816 1854 17826
tri 1854 17816 1864 17826 nw
tri 1900 17816 1910 17826 se
rect 1910 17816 1969 17826
rect 1662 17814 1732 17816
tri 1732 17814 1734 17816 nw
tri 1778 17814 1780 17816 se
rect 1780 17814 1849 17816
rect 1662 17811 1729 17814
tri 1729 17811 1732 17814 nw
tri 1775 17811 1778 17814 se
rect 1778 17811 1849 17814
tri 1849 17811 1854 17816 nw
tri 1895 17811 1900 17816 se
rect 1900 17811 1969 17816
tri 1969 17811 1984 17826 nw
tri 2015 17811 2030 17826 se
rect 2030 17818 7846 17826
tri 7846 17818 7854 17826 nw
tri 8512 17818 8520 17826 se
rect 8520 17818 9284 17826
rect 2030 17811 2089 17818
tri 2089 17811 2096 17818 nw
tri 8505 17811 8512 17818 se
rect 8512 17811 9284 17818
tri 1648 17804 1655 17811 se
rect 1655 17804 1722 17811
tri 1722 17804 1729 17811 nw
tri 1770 17806 1775 17811 se
rect 1775 17806 1844 17811
tri 1844 17806 1849 17811 nw
tri 1890 17806 1895 17811 se
rect 1895 17806 1964 17811
tri 1964 17806 1969 17811 nw
tri 2010 17806 2015 17811 se
rect 2015 17806 2082 17811
tri 1768 17804 1770 17806 se
rect 1770 17804 1842 17806
tri 1842 17804 1844 17806 nw
tri 1888 17804 1890 17806 se
rect 1890 17804 1962 17806
tri 1962 17804 1964 17806 nw
tri 2008 17804 2010 17806 se
rect 2010 17804 2082 17806
tri 2082 17804 2089 17811 nw
tri 8498 17804 8505 17811 se
rect 8505 17804 8596 17811
rect 1648 15736 1700 17804
tri 1700 17782 1722 17804 nw
tri 1746 17782 1768 17804 se
rect 1768 17782 1820 17804
tri 1820 17782 1842 17804 nw
tri 1866 17782 1888 17804 se
rect 1888 17796 1954 17804
tri 1954 17796 1962 17804 nw
tri 2000 17796 2008 17804 se
rect 2008 17796 2074 17804
tri 2074 17796 2082 17804 nw
tri 8490 17796 8498 17804 se
rect 8498 17796 8596 17804
rect 1888 17782 1940 17796
tri 1940 17782 1954 17796 nw
tri 1986 17782 2000 17796 se
rect 2000 17782 2060 17796
tri 2060 17782 2074 17796 nw
tri 8476 17782 8490 17796 se
rect 8490 17782 8596 17796
tri 1741 17777 1746 17782 se
rect 1746 17777 1815 17782
tri 1815 17777 1820 17782 nw
tri 1861 17777 1866 17782 se
rect 1866 17777 1935 17782
tri 1935 17777 1940 17782 nw
tri 1981 17777 1986 17782 se
rect 1986 17777 2055 17782
tri 2055 17777 2060 17782 nw
tri 8471 17777 8476 17782 se
rect 8476 17777 8596 17782
rect 8630 17777 8668 17811
rect 8702 17777 8740 17811
rect 8774 17777 8812 17811
rect 8846 17777 8884 17811
rect 8918 17777 8956 17811
rect 8990 17777 9028 17811
rect 9062 17777 9100 17811
rect 9134 17777 9172 17811
rect 9206 17777 9244 17811
rect 9278 17777 9284 17811
rect 1648 15672 1700 15684
rect 1648 15614 1700 15620
tri 1732 17768 1741 17777 se
rect 1741 17770 1808 17777
tri 1808 17770 1815 17777 nw
tri 1854 17770 1861 17777 se
rect 1861 17770 1926 17777
rect 1741 17768 1806 17770
tri 1806 17768 1808 17770 nw
tri 1852 17768 1854 17770 se
rect 1854 17768 1926 17770
tri 1926 17768 1935 17777 nw
tri 1972 17768 1981 17777 se
rect 1981 17768 2016 17777
rect 1564 14774 1616 14786
rect 1564 14716 1616 14722
rect 1648 15297 1700 15303
rect 1648 15233 1700 15245
rect 1480 9726 1532 9738
rect 1480 9638 1532 9674
rect 1396 3894 1448 3906
rect 1396 3836 1448 3842
rect 1312 58 1364 70
rect 1312 0 1364 6
rect 1648 122 1700 15181
rect 1732 11798 1784 17768
tri 1784 17746 1806 17768 nw
tri 1830 17746 1852 17768 se
rect 1852 17746 1896 17768
tri 1822 17738 1830 17746 se
rect 1830 17738 1896 17746
tri 1896 17738 1926 17768 nw
tri 1942 17738 1972 17768 se
rect 1972 17738 2016 17768
tri 2016 17738 2055 17777 nw
tri 8432 17738 8471 17777 se
rect 8471 17738 9284 17777
rect 1732 11734 1784 11746
rect 1732 11676 1784 11682
tri 1816 17732 1822 17738 se
rect 1822 17732 1890 17738
tri 1890 17732 1896 17738 nw
tri 1936 17732 1942 17738 se
rect 1942 17732 2000 17738
rect 1816 5640 1868 17732
tri 1868 17710 1890 17732 nw
tri 1926 17722 1936 17732 se
rect 1936 17722 2000 17732
tri 2000 17722 2016 17738 nw
tri 8416 17722 8432 17738 se
rect 8432 17722 8596 17738
tri 1914 17710 1926 17722 se
rect 1926 17710 1982 17722
tri 1908 17704 1914 17710 se
rect 1914 17704 1982 17710
tri 1982 17704 2000 17722 nw
tri 8398 17704 8416 17722 se
rect 8416 17704 8596 17722
rect 8630 17704 8668 17738
rect 8702 17704 8740 17738
rect 8774 17704 8812 17738
rect 8846 17704 8884 17738
rect 8918 17704 8956 17738
rect 8990 17704 9028 17738
rect 9062 17704 9100 17738
rect 9134 17704 9172 17738
rect 9206 17704 9244 17738
rect 9278 17704 9284 17738
tri 1900 17696 1908 17704 se
rect 1908 17696 1974 17704
tri 1974 17696 1982 17704 nw
tri 8390 17696 8398 17704 se
rect 8398 17696 9284 17704
rect 1900 12620 1952 17696
tri 1952 17674 1974 17696 nw
tri 8368 17674 8390 17696 se
rect 8390 17674 9284 17696
tri 8275 17581 8368 17674 se
rect 8368 17581 9284 17674
rect 7870 17549 9284 17581
rect 4998 16429 5004 16481
rect 5056 16429 5072 16481
rect 5124 16429 5140 16481
rect 5192 16472 7559 16481
rect 5192 16438 5232 16472
rect 5266 16438 5308 16472
rect 5342 16438 5385 16472
rect 5419 16438 5462 16472
rect 5496 16438 5572 16472
rect 5606 16438 5644 16472
rect 5678 16438 5716 16472
rect 5750 16438 5788 16472
rect 5822 16438 5860 16472
rect 5894 16438 5932 16472
rect 5966 16438 6004 16472
rect 6038 16438 6076 16472
rect 6110 16438 6148 16472
rect 6182 16438 6220 16472
rect 6254 16438 6292 16472
rect 6326 16438 6364 16472
rect 6398 16438 6436 16472
rect 6470 16438 6508 16472
rect 6542 16438 6580 16472
rect 6614 16438 6652 16472
rect 6686 16438 6724 16472
rect 6758 16438 6796 16472
rect 6830 16438 6868 16472
rect 6902 16438 6940 16472
rect 6974 16438 7012 16472
rect 7046 16438 7084 16472
rect 7118 16438 7156 16472
rect 7190 16438 7228 16472
rect 7262 16438 7301 16472
rect 7335 16438 7374 16472
rect 7408 16438 7447 16472
rect 7481 16438 7559 16472
rect 5192 16429 7559 16438
rect 4998 16400 5049 16429
tri 5049 16400 5078 16429 nw
tri 7479 16400 7508 16429 ne
rect 7508 16400 7559 16429
rect 4998 16366 5004 16400
rect 5038 16366 5044 16400
tri 5044 16395 5049 16400 nw
tri 7508 16395 7513 16400 ne
rect 4998 16327 5044 16366
rect 4998 16293 5004 16327
rect 5038 16293 5044 16327
rect 4998 16254 5044 16293
rect 4998 16220 5004 16254
rect 5038 16220 5044 16254
rect 4998 16181 5044 16220
rect 4998 16147 5004 16181
rect 5038 16147 5044 16181
rect 4998 16108 5044 16147
rect 4998 16074 5004 16108
rect 5038 16074 5044 16108
rect 4998 16035 5044 16074
rect 4998 16001 5004 16035
rect 5038 16001 5044 16035
rect 4998 15962 5044 16001
rect 4998 15928 5004 15962
rect 5038 15928 5044 15962
rect 4998 15889 5044 15928
rect 4998 15855 5004 15889
rect 5038 15855 5044 15889
rect 7513 16366 7519 16400
rect 7553 16366 7559 16400
rect 7513 16328 7559 16366
rect 7513 16294 7519 16328
rect 7553 16294 7559 16328
rect 7513 16256 7559 16294
rect 7513 16222 7519 16256
rect 7553 16222 7559 16256
rect 7513 16184 7559 16222
rect 7513 16150 7519 16184
rect 7553 16150 7559 16184
rect 7513 16112 7559 16150
rect 7513 16078 7519 16112
rect 7553 16078 7559 16112
rect 7513 16040 7559 16078
rect 7513 16006 7519 16040
rect 7553 16006 7559 16040
rect 7513 15968 7559 16006
rect 7513 15934 7519 15968
rect 7553 15934 7559 15968
rect 7513 15896 7559 15934
rect 4998 15816 5044 15855
rect 4998 15782 5004 15816
rect 5038 15782 5044 15816
rect 4998 15743 5044 15782
rect 4998 15709 5004 15743
rect 5038 15709 5044 15743
rect 4998 15670 5044 15709
rect 7044 15872 7212 15878
rect 7096 15820 7160 15872
rect 7044 15805 7212 15820
rect 7096 15753 7160 15805
rect 7044 15737 7212 15753
rect 7096 15685 7160 15737
rect 7044 15679 7212 15685
rect 7513 15862 7519 15896
rect 7553 15862 7559 15896
rect 7513 15824 7559 15862
rect 7513 15790 7519 15824
rect 7553 15790 7559 15824
rect 7513 15752 7559 15790
rect 7513 15718 7519 15752
rect 7553 15718 7559 15752
rect 7513 15680 7559 15718
rect 4998 15636 5004 15670
rect 5038 15636 5044 15670
rect 4998 15597 5044 15636
rect 1900 12556 1952 12568
rect 1900 12498 1952 12504
rect 2083 15509 2483 15531
rect 4416 15514 4422 15566
rect 4474 15514 4490 15566
rect 4542 15514 4558 15566
rect 4610 15514 4616 15566
rect 2083 15457 2089 15509
rect 2141 15457 2173 15509
rect 2225 15457 2257 15509
rect 2309 15457 2341 15509
rect 2393 15457 2425 15509
rect 2477 15457 2483 15509
rect 2083 15419 2483 15457
rect 2083 15367 2089 15419
rect 2141 15367 2173 15419
rect 2225 15367 2257 15419
rect 2309 15367 2341 15419
rect 2393 15367 2425 15419
rect 2477 15367 2483 15419
rect 2876 15457 2882 15509
rect 2934 15457 2995 15509
rect 3047 15457 3107 15509
rect 3159 15457 3165 15509
rect 2876 15419 3165 15457
rect 4416 15482 4616 15514
rect 4416 15430 4422 15482
rect 4474 15430 4490 15482
rect 4542 15430 4558 15482
rect 4610 15430 4616 15482
rect 4998 15563 5004 15597
rect 5038 15563 5044 15597
rect 4998 15524 5044 15563
rect 4998 15490 5004 15524
rect 5038 15490 5044 15524
rect 4998 15451 5044 15490
rect 2876 15367 2882 15419
rect 2934 15367 2995 15419
rect 3047 15367 3107 15419
rect 3159 15367 3165 15419
rect 4998 15417 5004 15451
rect 5038 15417 5044 15451
rect 4998 15378 5044 15417
rect 1816 5576 1868 5588
rect 1816 5518 1868 5524
rect 1900 12239 1952 12245
rect 1900 12175 1952 12187
rect 1648 58 1700 70
rect 1648 0 1700 6
rect 1900 122 1952 12123
rect 2083 11975 2483 15367
rect 4998 15344 5004 15378
rect 5038 15344 5044 15378
rect 4998 15305 5044 15344
rect 4998 15271 5004 15305
rect 5038 15271 5044 15305
rect 4998 15232 5044 15271
rect 4998 15198 5004 15232
rect 5038 15198 5044 15232
rect 4998 15159 5044 15198
rect 4998 15125 5004 15159
rect 5038 15125 5044 15159
rect 4998 15086 5044 15125
rect 4998 15052 5004 15086
rect 5038 15052 5044 15086
rect 4998 15013 5044 15052
rect 4998 14979 5004 15013
rect 5038 14979 5044 15013
rect 4998 14940 5044 14979
rect 4998 14906 5004 14940
rect 5038 14906 5044 14940
rect 4998 14867 5044 14906
rect 4998 14833 5004 14867
rect 5038 14833 5044 14867
rect 4998 14795 5044 14833
rect 4998 14761 5004 14795
rect 5038 14761 5044 14795
rect 4998 14723 5044 14761
rect 4998 14689 5004 14723
rect 5038 14689 5044 14723
rect 3877 14678 4077 14684
rect 3929 14626 3951 14678
rect 4003 14626 4025 14678
rect 3877 14610 4077 14626
rect 3929 14558 3951 14610
rect 4003 14558 4025 14610
rect 3877 14542 4077 14558
rect 3929 14490 3951 14542
rect 4003 14490 4025 14542
rect 3877 14484 4077 14490
rect 4998 14651 5044 14689
rect 4998 14617 5004 14651
rect 5038 14617 5044 14651
rect 4998 14579 5044 14617
rect 4998 14545 5004 14579
rect 5038 14545 5044 14579
rect 4998 14507 5044 14545
rect 4998 14473 5004 14507
rect 5038 14473 5044 14507
rect 4998 14435 5044 14473
rect 4416 14371 4422 14423
rect 4474 14371 4490 14423
rect 4542 14371 4558 14423
rect 4610 14371 4616 14423
rect 4416 14339 4616 14371
rect 4416 14287 4422 14339
rect 4474 14287 4490 14339
rect 4542 14287 4558 14339
rect 4610 14287 4616 14339
rect 4998 14401 5004 14435
rect 5038 14401 5044 14435
rect 4998 14363 5044 14401
rect 4998 14329 5004 14363
rect 5038 14329 5044 14363
rect 4998 14291 5044 14329
rect 4998 14257 5004 14291
rect 5038 14257 5044 14291
rect 4998 14219 5044 14257
rect 4998 14185 5004 14219
rect 5038 14185 5044 14219
rect 4998 14147 5044 14185
rect 7513 15646 7519 15680
rect 7553 15646 7559 15680
rect 7513 15608 7559 15646
rect 7513 15574 7519 15608
rect 7553 15574 7559 15608
rect 7513 15536 7559 15574
rect 7513 15502 7519 15536
rect 7553 15502 7559 15536
rect 7513 15464 7559 15502
rect 7513 15430 7519 15464
rect 7553 15430 7559 15464
rect 7513 15392 7559 15430
rect 7513 15358 7519 15392
rect 7553 15358 7559 15392
rect 7513 15320 7559 15358
rect 7513 15286 7519 15320
rect 7553 15286 7559 15320
rect 7513 15248 7559 15286
rect 7513 15214 7519 15248
rect 7553 15214 7559 15248
rect 7513 15176 7559 15214
rect 7513 15142 7519 15176
rect 7553 15142 7559 15176
rect 7513 15104 7559 15142
rect 7513 15070 7519 15104
rect 7553 15070 7559 15104
rect 7513 15032 7559 15070
rect 7513 14998 7519 15032
rect 7553 14998 7559 15032
rect 7513 14960 7559 14998
rect 7513 14926 7519 14960
rect 7553 14926 7559 14960
rect 7513 14888 7559 14926
rect 7513 14854 7519 14888
rect 7553 14854 7559 14888
rect 7513 14816 7559 14854
rect 7513 14782 7519 14816
rect 7553 14782 7559 14816
rect 7513 14744 7559 14782
rect 7513 14710 7519 14744
rect 7553 14710 7559 14744
rect 7513 14672 7559 14710
rect 7513 14638 7519 14672
rect 7553 14638 7559 14672
rect 7513 14600 7559 14638
rect 7513 14566 7519 14600
rect 7553 14566 7559 14600
rect 7513 14528 7559 14566
rect 7513 14494 7519 14528
rect 7553 14494 7559 14528
rect 7513 14456 7559 14494
rect 7513 14422 7519 14456
rect 7553 14422 7559 14456
rect 7513 14384 7559 14422
rect 7513 14350 7519 14384
rect 7553 14350 7559 14384
rect 7513 14312 7559 14350
rect 7513 14278 7519 14312
rect 7553 14278 7559 14312
rect 7513 14240 7559 14278
rect 7513 14206 7519 14240
rect 7553 14206 7559 14240
rect 7513 14168 7559 14206
rect 4998 14113 5004 14147
rect 5038 14113 5044 14147
rect 4998 14075 5044 14113
rect 4998 14041 5004 14075
rect 5038 14041 5044 14075
rect 4998 14003 5044 14041
rect 4998 13969 5004 14003
rect 5038 13969 5044 14003
rect 4998 13931 5044 13969
rect 7044 14153 7212 14159
rect 7096 14101 7160 14153
rect 7044 14086 7212 14101
rect 7096 14034 7160 14086
rect 7044 14018 7212 14034
rect 7096 13966 7160 14018
rect 7044 13960 7212 13966
rect 7513 14134 7519 14168
rect 7553 14134 7559 14168
rect 7513 14096 7559 14134
rect 7513 14062 7519 14096
rect 7553 14062 7559 14096
rect 7513 14024 7559 14062
rect 7513 13990 7519 14024
rect 7553 13990 7559 14024
rect 4998 13897 5004 13931
rect 5038 13897 5044 13931
rect 4998 13859 5044 13897
rect 4998 13825 5004 13859
rect 5038 13825 5044 13859
rect 2917 13789 3024 13795
rect 2917 13737 2944 13789
rect 2996 13737 3024 13789
rect 2917 13721 3024 13737
rect 2917 13669 2944 13721
rect 2996 13669 3024 13721
rect 2917 13653 3024 13669
rect 2917 13601 2944 13653
rect 2996 13601 3024 13653
rect 2917 13595 3024 13601
rect 3877 13462 4077 13822
rect 4998 13787 5044 13825
rect 4416 13042 4616 13784
rect 4656 13544 4708 13775
rect 4736 13544 4788 13775
rect 4998 13753 5004 13787
rect 5038 13753 5044 13787
rect 4998 13715 5044 13753
rect 4998 13681 5004 13715
rect 5038 13681 5044 13715
rect 4998 13643 5044 13681
rect 4998 13609 5004 13643
rect 5038 13609 5044 13643
rect 4998 13571 5044 13609
rect 4416 12990 4422 13042
rect 4474 12990 4490 13042
rect 4542 12990 4558 13042
rect 4610 12990 4616 13042
rect 4416 12958 4616 12990
rect 4416 12906 4422 12958
rect 4474 12906 4490 12958
rect 4542 12906 4558 12958
rect 4610 12906 4616 12958
rect 3877 12852 4077 12858
rect 3929 12800 3951 12852
rect 4003 12800 4025 12852
rect 3877 12784 4077 12800
rect 3929 12732 3951 12784
rect 4003 12732 4025 12784
rect 3877 12716 4077 12732
rect 3929 12664 3951 12716
rect 4003 12664 4025 12716
rect 3877 12658 4077 12664
rect 2083 11923 2089 11975
rect 2141 11923 2173 11975
rect 2225 11923 2257 11975
rect 2309 11923 2341 11975
rect 2393 11923 2425 11975
rect 2477 11923 2483 11975
rect 2083 11885 2483 11923
rect 2083 11833 2089 11885
rect 2141 11833 2173 11885
rect 2225 11833 2257 11885
rect 2309 11833 2341 11885
rect 2393 11833 2425 11885
rect 2477 11833 2483 11885
rect 2876 11923 2882 11975
rect 2934 11923 2995 11975
rect 3047 11923 3107 11975
rect 3159 11923 3165 11975
rect 2876 11885 3165 11923
rect 2876 11833 2882 11885
rect 2934 11833 2995 11885
rect 3047 11833 3107 11885
rect 3159 11833 3165 11885
rect 4416 11909 4616 12906
rect 4416 11857 4422 11909
rect 4474 11857 4490 11909
rect 4542 11857 4558 11909
rect 4610 11857 4616 11909
rect 2083 10461 2483 11833
rect 4416 11825 4616 11857
rect 4416 11773 4422 11825
rect 4474 11773 4490 11825
rect 4542 11773 4558 11825
rect 4610 11773 4616 11825
rect 4416 11461 4616 11773
rect 4416 11409 4433 11461
rect 4485 11409 4558 11461
rect 4610 11409 4616 11461
rect 4416 11377 4616 11409
rect 4416 11325 4433 11377
rect 4485 11325 4558 11377
rect 4610 11325 4616 11377
rect 2917 11223 3024 11272
rect 2917 11216 3051 11223
tri 3051 11216 3058 11223 nw
rect 2917 11195 3030 11216
tri 3030 11195 3051 11216 nw
rect 2917 11089 3024 11195
tri 3024 11189 3030 11195 nw
tri 3024 11089 3040 11105 sw
rect 2917 11072 3040 11089
tri 3040 11072 3057 11089 sw
rect 2917 11071 3057 11072
tri 3057 11071 3058 11072 sw
rect 2917 11040 3024 11071
rect 3877 10982 4077 11315
rect 4416 10511 4616 11325
rect 4998 13537 5004 13571
rect 5038 13537 5044 13571
rect 4998 13499 5044 13537
rect 4998 13465 5004 13499
rect 5038 13465 5044 13499
rect 4998 13427 5044 13465
rect 7513 13952 7559 13990
rect 7513 13918 7519 13952
rect 7553 13918 7559 13952
rect 7513 13880 7559 13918
rect 7513 13846 7519 13880
rect 7553 13846 7559 13880
rect 7513 13808 7559 13846
rect 7513 13774 7519 13808
rect 7553 13774 7559 13808
rect 7513 13736 7559 13774
rect 7513 13702 7519 13736
rect 7553 13702 7559 13736
rect 7513 13664 7559 13702
rect 7513 13630 7519 13664
rect 7553 13630 7559 13664
rect 7513 13592 7559 13630
rect 7513 13558 7519 13592
rect 7553 13558 7559 13592
rect 7513 13520 7559 13558
rect 7513 13486 7519 13520
rect 7553 13486 7559 13520
rect 7513 13448 7559 13486
rect 4998 13393 5004 13427
rect 5038 13393 5044 13427
rect 4998 13355 5044 13393
rect 4998 13321 5004 13355
rect 5038 13321 5044 13355
rect 4998 13283 5044 13321
rect 4998 13249 5004 13283
rect 5038 13249 5044 13283
rect 4998 13211 5044 13249
rect 7044 13431 7212 13437
rect 7096 13379 7160 13431
rect 7044 13364 7212 13379
rect 7096 13312 7160 13364
rect 7044 13296 7212 13312
rect 7096 13244 7160 13296
rect 7044 13238 7212 13244
rect 7513 13414 7519 13448
rect 7553 13414 7559 13448
rect 7513 13376 7559 13414
rect 7513 13342 7519 13376
rect 7553 13342 7559 13376
rect 7513 13304 7559 13342
rect 7513 13270 7519 13304
rect 7553 13270 7559 13304
rect 4998 13177 5004 13211
rect 5038 13177 5044 13211
rect 4998 13139 5044 13177
rect 4998 13105 5004 13139
rect 5038 13105 5044 13139
rect 4998 13067 5044 13105
rect 4998 13033 5004 13067
rect 5038 13033 5044 13067
rect 4998 12995 5044 13033
rect 4998 12961 5004 12995
rect 5038 12961 5044 12995
rect 4998 12923 5044 12961
rect 4998 12889 5004 12923
rect 5038 12889 5044 12923
rect 4998 12851 5044 12889
rect 4998 12817 5004 12851
rect 5038 12817 5044 12851
rect 4998 12779 5044 12817
rect 4998 12745 5004 12779
rect 5038 12745 5044 12779
rect 4998 12707 5044 12745
rect 4998 12673 5004 12707
rect 5038 12673 5044 12707
rect 4998 12635 5044 12673
rect 4998 12601 5004 12635
rect 5038 12601 5044 12635
rect 4998 12563 5044 12601
rect 4998 12529 5004 12563
rect 5038 12529 5044 12563
rect 4998 12491 5044 12529
rect 4998 12457 5004 12491
rect 5038 12457 5044 12491
rect 4998 12419 5044 12457
rect 4998 12385 5004 12419
rect 5038 12385 5044 12419
rect 4998 12347 5044 12385
rect 4998 12313 5004 12347
rect 5038 12313 5044 12347
rect 4998 12275 5044 12313
rect 4998 12241 5004 12275
rect 5038 12241 5044 12275
rect 4998 12203 5044 12241
rect 4998 12169 5004 12203
rect 5038 12169 5044 12203
rect 4998 12131 5044 12169
rect 4998 12097 5004 12131
rect 5038 12097 5044 12131
rect 4998 12059 5044 12097
rect 4998 12025 5004 12059
rect 5038 12025 5044 12059
rect 4998 11987 5044 12025
rect 4998 11953 5004 11987
rect 5038 11953 5044 11987
rect 4998 11915 5044 11953
rect 4998 11881 5004 11915
rect 5038 11881 5044 11915
rect 4998 11843 5044 11881
rect 4998 11809 5004 11843
rect 5038 11809 5044 11843
rect 4998 11771 5044 11809
rect 4998 11737 5004 11771
rect 5038 11737 5044 11771
rect 4998 11699 5044 11737
rect 4998 11665 5004 11699
rect 5038 11665 5044 11699
rect 4998 11627 5044 11665
rect 7513 13232 7559 13270
rect 7513 13198 7519 13232
rect 7553 13198 7559 13232
rect 7513 13160 7559 13198
rect 7513 13126 7519 13160
rect 7553 13126 7559 13160
rect 7513 13088 7559 13126
rect 7513 13054 7519 13088
rect 7553 13054 7559 13088
rect 7513 13016 7559 13054
rect 7513 12982 7519 13016
rect 7553 12982 7559 13016
rect 7513 12944 7559 12982
rect 7513 12910 7519 12944
rect 7553 12910 7559 12944
rect 7513 12872 7559 12910
rect 7513 12838 7519 12872
rect 7553 12838 7559 12872
rect 7513 12800 7559 12838
rect 7513 12766 7519 12800
rect 7553 12766 7559 12800
rect 7513 12728 7559 12766
rect 7513 12694 7519 12728
rect 7553 12694 7559 12728
rect 7513 12656 7559 12694
rect 7513 12622 7519 12656
rect 7553 12622 7559 12656
rect 7513 12584 7559 12622
rect 7513 12550 7519 12584
rect 7553 12550 7559 12584
rect 7513 12512 7559 12550
rect 7513 12478 7519 12512
rect 7553 12478 7559 12512
rect 7513 12440 7559 12478
rect 7513 12406 7519 12440
rect 7553 12406 7559 12440
rect 7513 12368 7559 12406
rect 7513 12334 7519 12368
rect 7553 12334 7559 12368
rect 7513 12296 7559 12334
rect 7513 12262 7519 12296
rect 7553 12262 7559 12296
rect 7513 12224 7559 12262
rect 7513 12190 7519 12224
rect 7553 12190 7559 12224
rect 7513 12152 7559 12190
rect 7513 12118 7519 12152
rect 7553 12118 7559 12152
rect 7513 12080 7559 12118
rect 7513 12046 7519 12080
rect 7553 12046 7559 12080
rect 7513 12008 7559 12046
rect 7513 11974 7519 12008
rect 7553 11974 7559 12008
rect 7513 11936 7559 11974
rect 7513 11902 7519 11936
rect 7553 11902 7559 11936
rect 7513 11864 7559 11902
rect 7513 11830 7519 11864
rect 7553 11830 7559 11864
rect 7513 11792 7559 11830
rect 7513 11758 7519 11792
rect 7553 11758 7559 11792
rect 7513 11720 7559 11758
rect 7513 11686 7519 11720
rect 7553 11686 7559 11720
rect 7513 11648 7559 11686
rect 4998 11593 5004 11627
rect 5038 11593 5044 11627
rect 4998 11555 5044 11593
rect 4998 11521 5004 11555
rect 5038 11521 5044 11555
rect 4998 11483 5044 11521
rect 4998 11449 5004 11483
rect 5038 11449 5044 11483
rect 4998 11411 5044 11449
rect 7044 11632 7212 11638
rect 7096 11580 7160 11632
rect 7044 11565 7212 11580
rect 7096 11513 7160 11565
rect 7044 11497 7212 11513
rect 7096 11445 7160 11497
rect 7044 11439 7212 11445
rect 7513 11614 7519 11648
rect 7553 11614 7559 11648
rect 7513 11576 7559 11614
rect 7513 11542 7519 11576
rect 7553 11542 7559 11576
rect 7513 11504 7559 11542
rect 7513 11470 7519 11504
rect 7553 11470 7559 11504
rect 4998 11377 5004 11411
rect 5038 11377 5044 11411
rect 4998 11339 5044 11377
rect 4998 11305 5004 11339
rect 5038 11305 5044 11339
rect 4998 11267 5044 11305
rect 4656 11035 4708 11266
rect 4736 11035 4788 11266
rect 4998 11233 5004 11267
rect 5038 11233 5044 11267
rect 4998 11195 5044 11233
rect 4998 11161 5004 11195
rect 5038 11161 5044 11195
rect 4998 11123 5044 11161
rect 4998 11089 5004 11123
rect 5038 11089 5044 11123
rect 4998 11051 5044 11089
rect 2083 10409 2089 10461
rect 2141 10409 2173 10461
rect 2225 10409 2257 10461
rect 2309 10409 2341 10461
rect 2393 10409 2425 10461
rect 2477 10409 2483 10461
rect 2083 10371 2483 10409
rect 2083 10319 2089 10371
rect 2141 10319 2173 10371
rect 2225 10319 2257 10371
rect 2309 10319 2341 10371
rect 2393 10319 2425 10371
rect 2477 10319 2483 10371
rect 2876 10409 2882 10461
rect 2934 10409 2995 10461
rect 3047 10409 3107 10461
rect 3159 10409 3165 10461
rect 2876 10371 3165 10409
rect 2876 10319 2882 10371
rect 2934 10319 2995 10371
rect 3047 10319 3107 10371
rect 3159 10319 3165 10371
rect 4416 10459 4422 10511
rect 4474 10459 4490 10511
rect 4542 10459 4558 10511
rect 4610 10459 4616 10511
rect 4416 10427 4616 10459
rect 4416 10375 4422 10427
rect 4474 10375 4490 10427
rect 4542 10375 4558 10427
rect 4610 10375 4616 10427
rect 2083 9241 2483 10319
rect 3877 9630 4077 9636
rect 3929 9578 3951 9630
rect 4003 9578 4025 9630
rect 3877 9562 4077 9578
rect 3929 9510 3951 9562
rect 4003 9510 4025 9562
rect 3877 9494 4077 9510
rect 3929 9442 3951 9494
rect 4003 9442 4025 9494
rect 3877 9436 4077 9442
rect 2083 9189 2085 9241
rect 2137 9189 2171 9241
rect 2223 9189 2257 9241
rect 2309 9189 2343 9241
rect 2395 9189 2429 9241
rect 2481 9189 2483 9241
rect 2083 9160 2483 9189
rect 2083 9108 2085 9160
rect 2137 9108 2171 9160
rect 2223 9108 2257 9160
rect 2309 9108 2343 9160
rect 2395 9108 2429 9160
rect 2481 9108 2483 9160
rect 2083 9079 2483 9108
rect 2083 9027 2085 9079
rect 2137 9027 2171 9079
rect 2223 9027 2257 9079
rect 2309 9027 2343 9079
rect 2395 9027 2429 9079
rect 2481 9027 2483 9079
rect 2083 8997 2483 9027
rect 2083 8945 2085 8997
rect 2137 8945 2171 8997
rect 2223 8945 2257 8997
rect 2309 8945 2343 8997
rect 2395 8945 2429 8997
rect 2481 8945 2483 8997
rect 2083 8915 2483 8945
rect 2083 8863 2085 8915
rect 2137 8863 2171 8915
rect 2223 8863 2257 8915
rect 2309 8863 2343 8915
rect 2395 8863 2429 8915
rect 2481 8863 2483 8915
rect 2083 8833 2483 8863
rect 2083 8781 2085 8833
rect 2137 8781 2171 8833
rect 2223 8781 2257 8833
rect 2309 8781 2343 8833
rect 2395 8781 2429 8833
rect 2481 8781 2483 8833
rect 4416 9389 4616 10375
rect 4416 9337 4422 9389
rect 4474 9337 4490 9389
rect 4542 9337 4558 9389
rect 4610 9337 4616 9389
rect 4416 9305 4616 9337
rect 4416 9253 4422 9305
rect 4474 9253 4490 9305
rect 4542 9253 4558 9305
rect 4610 9253 4616 9305
rect 2083 6927 2483 8781
rect 2917 8710 3024 8783
rect 2917 8658 2944 8710
rect 2996 8658 3024 8710
rect 2917 8642 3024 8658
rect 2917 8590 2944 8642
rect 2996 8590 3024 8642
rect 2917 8583 3024 8590
rect 2917 8574 3023 8583
rect 2917 8522 2944 8574
rect 2996 8522 3023 8574
rect 2917 8516 3023 8522
rect 3877 8450 4077 8810
rect 4416 8002 4616 9253
rect 4998 11017 5004 11051
rect 5038 11017 5044 11051
rect 4998 10979 5044 11017
rect 4998 10945 5004 10979
rect 5038 10945 5044 10979
rect 7513 11432 7559 11470
rect 7513 11398 7519 11432
rect 7553 11398 7559 11432
rect 7513 11360 7559 11398
rect 7513 11326 7519 11360
rect 7553 11326 7559 11360
rect 7513 11288 7559 11326
rect 7513 11254 7519 11288
rect 7553 11254 7559 11288
rect 7513 11216 7559 11254
rect 7513 11182 7519 11216
rect 7553 11182 7559 11216
rect 7513 11144 7559 11182
rect 7513 11110 7519 11144
rect 7553 11110 7559 11144
rect 7513 11072 7559 11110
rect 7513 11038 7519 11072
rect 7553 11038 7559 11072
rect 7513 11000 7559 11038
rect 7513 10966 7519 11000
rect 7553 10966 7559 11000
rect 4998 10907 5044 10945
rect 4998 10873 5004 10907
rect 5038 10873 5044 10907
rect 4998 10835 5044 10873
rect 4998 10801 5004 10835
rect 5038 10801 5044 10835
rect 4998 10763 5044 10801
rect 4998 10729 5004 10763
rect 5038 10729 5044 10763
rect 7044 10944 7212 10950
rect 7096 10892 7160 10944
rect 7044 10877 7212 10892
rect 7096 10825 7160 10877
rect 7044 10809 7212 10825
rect 7096 10757 7160 10809
rect 7044 10751 7212 10757
rect 7513 10928 7559 10966
rect 7513 10894 7519 10928
rect 7553 10894 7559 10928
rect 7513 10856 7559 10894
rect 7513 10822 7519 10856
rect 7553 10822 7559 10856
rect 7513 10784 7559 10822
rect 4998 10691 5044 10729
rect 4998 10657 5004 10691
rect 5038 10657 5044 10691
rect 4998 10619 5044 10657
rect 4998 10585 5004 10619
rect 5038 10585 5044 10619
rect 4998 10547 5044 10585
rect 4998 10513 5004 10547
rect 5038 10513 5044 10547
rect 4998 10475 5044 10513
rect 4998 10441 5004 10475
rect 5038 10441 5044 10475
rect 4998 10403 5044 10441
rect 4998 10369 5004 10403
rect 5038 10369 5044 10403
rect 4998 10331 5044 10369
rect 4998 10297 5004 10331
rect 5038 10297 5044 10331
rect 4998 10259 5044 10297
rect 4998 10225 5004 10259
rect 5038 10225 5044 10259
rect 4998 10187 5044 10225
rect 4998 10153 5004 10187
rect 5038 10153 5044 10187
rect 4998 10115 5044 10153
rect 4998 10081 5004 10115
rect 5038 10081 5044 10115
rect 4998 10043 5044 10081
rect 4998 10009 5004 10043
rect 5038 10009 5044 10043
rect 4998 9971 5044 10009
rect 4998 9937 5004 9971
rect 5038 9937 5044 9971
rect 4998 9899 5044 9937
rect 4998 9865 5004 9899
rect 5038 9865 5044 9899
rect 4998 9827 5044 9865
rect 4998 9793 5004 9827
rect 5038 9793 5044 9827
rect 4998 9755 5044 9793
rect 4998 9721 5004 9755
rect 5038 9721 5044 9755
rect 4998 9683 5044 9721
rect 4998 9649 5004 9683
rect 5038 9649 5044 9683
rect 4998 9611 5044 9649
rect 4998 9577 5004 9611
rect 5038 9577 5044 9611
rect 4998 9539 5044 9577
rect 4998 9505 5004 9539
rect 5038 9505 5044 9539
rect 4998 9467 5044 9505
rect 4998 9433 5004 9467
rect 5038 9433 5044 9467
rect 4998 9395 5044 9433
rect 4998 9361 5004 9395
rect 5038 9361 5044 9395
rect 4998 9323 5044 9361
rect 4998 9289 5004 9323
rect 5038 9289 5044 9323
rect 4998 9251 5044 9289
rect 4998 9217 5004 9251
rect 5038 9217 5044 9251
rect 4998 9179 5044 9217
rect 7513 10750 7519 10784
rect 7553 10750 7559 10784
rect 7513 10712 7559 10750
rect 7513 10678 7519 10712
rect 7553 10678 7559 10712
rect 7513 10640 7559 10678
rect 7513 10606 7519 10640
rect 7553 10606 7559 10640
rect 7513 10568 7559 10606
rect 7513 10534 7519 10568
rect 7553 10534 7559 10568
rect 7513 10496 7559 10534
rect 7513 10462 7519 10496
rect 7553 10462 7559 10496
rect 7513 10424 7559 10462
rect 7513 10390 7519 10424
rect 7553 10390 7559 10424
rect 7513 10352 7559 10390
rect 7513 10318 7519 10352
rect 7553 10318 7559 10352
rect 7513 10280 7559 10318
rect 7513 10246 7519 10280
rect 7553 10246 7559 10280
rect 7513 10208 7559 10246
rect 7513 10174 7519 10208
rect 7553 10174 7559 10208
rect 7513 10136 7559 10174
rect 7513 10102 7519 10136
rect 7553 10102 7559 10136
rect 7513 10064 7559 10102
rect 7513 10030 7519 10064
rect 7553 10030 7559 10064
rect 7513 9992 7559 10030
rect 7513 9958 7519 9992
rect 7553 9958 7559 9992
rect 7513 9920 7559 9958
rect 7513 9886 7519 9920
rect 7553 9886 7559 9920
rect 7513 9848 7559 9886
rect 7513 9814 7519 9848
rect 7553 9814 7559 9848
rect 7513 9776 7559 9814
rect 7513 9742 7519 9776
rect 7553 9742 7559 9776
rect 7513 9704 7559 9742
rect 7513 9670 7519 9704
rect 7553 9670 7559 9704
rect 7513 9632 7559 9670
rect 7513 9598 7519 9632
rect 7553 9598 7559 9632
rect 7513 9560 7559 9598
rect 7513 9526 7519 9560
rect 7553 9526 7559 9560
rect 7513 9488 7559 9526
rect 7513 9454 7519 9488
rect 7553 9454 7559 9488
rect 7513 9416 7559 9454
rect 7513 9382 7519 9416
rect 7553 9382 7559 9416
rect 7513 9344 7559 9382
rect 7513 9310 7519 9344
rect 7553 9310 7559 9344
rect 7513 9272 7559 9310
rect 7513 9238 7519 9272
rect 7553 9238 7559 9272
rect 4998 9145 5004 9179
rect 5038 9145 5044 9179
rect 4998 9107 5044 9145
rect 4998 9073 5004 9107
rect 5038 9073 5044 9107
rect 4998 9035 5044 9073
rect 4998 9001 5004 9035
rect 5038 9001 5044 9035
rect 7044 9198 7212 9204
rect 7096 9146 7160 9198
rect 7044 9131 7212 9146
rect 7096 9079 7160 9131
rect 7044 9063 7212 9079
rect 7096 9011 7160 9063
rect 7044 9005 7212 9011
rect 7513 9200 7559 9238
rect 7513 9166 7519 9200
rect 7553 9166 7559 9200
rect 7513 9128 7559 9166
rect 7513 9094 7519 9128
rect 7553 9094 7559 9128
rect 7513 9056 7559 9094
rect 7513 9022 7519 9056
rect 7553 9022 7559 9056
rect 4998 8963 5044 9001
rect 4998 8929 5004 8963
rect 5038 8929 5044 8963
rect 4998 8891 5044 8929
rect 4998 8857 5004 8891
rect 5038 8857 5044 8891
rect 4998 8819 5044 8857
rect 4998 8785 5004 8819
rect 5038 8785 5044 8819
rect 4998 8747 5044 8785
rect 4656 8513 4708 8744
rect 4736 8513 4788 8744
rect 4998 8713 5004 8747
rect 5038 8713 5044 8747
rect 4998 8675 5044 8713
rect 4998 8641 5004 8675
rect 5038 8641 5044 8675
rect 4998 8603 5044 8641
rect 4998 8569 5004 8603
rect 5038 8569 5044 8603
rect 4998 8531 5044 8569
rect 4416 7950 4422 8002
rect 4474 7950 4490 8002
rect 4542 7950 4558 8002
rect 4610 7950 4616 8002
rect 4416 7918 4616 7950
rect 4416 7866 4422 7918
rect 4474 7866 4490 7918
rect 4542 7866 4558 7918
rect 4610 7866 4616 7918
rect 3877 7804 4077 7810
rect 3929 7752 3951 7804
rect 4003 7752 4025 7804
rect 3877 7736 4077 7752
rect 3929 7684 3951 7736
rect 4003 7684 4025 7736
rect 3877 7668 4077 7684
rect 3929 7616 3951 7668
rect 4003 7616 4025 7668
rect 3877 7610 4077 7616
rect 2083 6875 2089 6927
rect 2141 6875 2173 6927
rect 2225 6875 2257 6927
rect 2309 6875 2341 6927
rect 2393 6875 2425 6927
rect 2477 6875 2483 6927
rect 2083 6837 2483 6875
rect 2083 6785 2089 6837
rect 2141 6785 2173 6837
rect 2225 6785 2257 6837
rect 2309 6785 2341 6837
rect 2393 6785 2425 6837
rect 2477 6785 2483 6837
rect 2083 5413 2483 6785
rect 2083 5361 2089 5413
rect 2141 5361 2173 5413
rect 2225 5361 2257 5413
rect 2309 5361 2341 5413
rect 2393 5361 2425 5413
rect 2477 5361 2483 5413
rect 2083 5323 2483 5361
rect 2083 5271 2089 5323
rect 2141 5271 2173 5323
rect 2225 5271 2257 5323
rect 2309 5271 2341 5323
rect 2393 5271 2425 5323
rect 2477 5271 2483 5323
rect 2656 7191 2708 7197
rect 2656 7127 2708 7139
rect 1900 58 1952 70
rect 1900 0 1952 6
rect 2152 5201 2204 5207
rect 2152 5137 2204 5149
rect 2152 122 2204 5085
rect 2152 58 2204 70
rect 2152 0 2204 6
rect 2404 4399 2456 4405
rect 2404 4335 2456 4347
rect 2404 122 2456 4283
rect 2404 58 2456 70
rect 2404 0 2456 6
rect 2656 122 2708 7075
rect 2876 6875 2882 6927
rect 2934 6875 2995 6927
rect 3047 6875 3107 6927
rect 3159 6875 3165 6927
rect 2876 6837 3165 6875
rect 2876 6785 2882 6837
rect 2934 6785 2995 6837
rect 3047 6785 3107 6837
rect 3159 6785 3165 6837
rect 4416 6880 4616 7866
rect 4416 6828 4422 6880
rect 4474 6828 4490 6880
rect 4542 6828 4558 6880
rect 4610 6828 4616 6880
rect 4416 6796 4616 6828
rect 4416 6744 4422 6796
rect 4474 6744 4490 6796
rect 4542 6744 4558 6796
rect 4610 6744 4616 6796
rect 2917 6175 3024 6197
rect 2917 6155 3038 6175
tri 3038 6155 3058 6175 nw
rect 2917 6049 3024 6155
tri 3024 6141 3038 6155 nw
tri 3024 6049 3032 6057 sw
rect 2917 6032 3032 6049
tri 3032 6032 3049 6049 sw
rect 2917 6023 3049 6032
tri 3049 6023 3058 6032 sw
rect 2917 5997 3024 6023
rect 3877 5950 4077 6220
rect 4416 5486 4616 6744
rect 4998 8497 5004 8531
rect 5038 8497 5044 8531
rect 4998 8459 5044 8497
rect 4998 8425 5004 8459
rect 5038 8425 5044 8459
rect 7513 8984 7559 9022
rect 7513 8950 7519 8984
rect 7553 8950 7559 8984
rect 7513 8912 7559 8950
rect 7513 8878 7519 8912
rect 7553 8878 7559 8912
rect 7513 8840 7559 8878
rect 7513 8806 7519 8840
rect 7553 8806 7559 8840
rect 7513 8768 7559 8806
rect 7513 8734 7519 8768
rect 7553 8734 7559 8768
rect 7513 8696 7559 8734
rect 7513 8662 7519 8696
rect 7553 8662 7559 8696
rect 7513 8624 7559 8662
rect 7513 8590 7519 8624
rect 7553 8590 7559 8624
rect 7513 8552 7559 8590
rect 7513 8518 7519 8552
rect 7553 8518 7559 8552
rect 7513 8480 7559 8518
rect 7513 8446 7519 8480
rect 7553 8446 7559 8480
rect 4998 8387 5044 8425
rect 4998 8353 5004 8387
rect 5038 8353 5044 8387
rect 4998 8315 5044 8353
rect 4998 8281 5004 8315
rect 5038 8281 5044 8315
rect 4998 8243 5044 8281
rect 4998 8209 5004 8243
rect 5038 8209 5044 8243
rect 7044 8429 7212 8435
rect 7096 8377 7160 8429
rect 7044 8362 7212 8377
rect 7096 8310 7160 8362
rect 7044 8294 7212 8310
rect 7096 8242 7160 8294
rect 7044 8236 7212 8242
rect 7513 8408 7559 8446
rect 7513 8374 7519 8408
rect 7553 8374 7559 8408
rect 7513 8336 7559 8374
rect 7513 8302 7519 8336
rect 7553 8302 7559 8336
rect 7513 8264 7559 8302
rect 4998 8171 5044 8209
rect 4998 8137 5004 8171
rect 5038 8137 5044 8171
rect 4998 8099 5044 8137
rect 4998 8065 5004 8099
rect 5038 8065 5044 8099
rect 4998 8027 5044 8065
rect 4998 7993 5004 8027
rect 5038 7993 5044 8027
rect 4998 7955 5044 7993
rect 4998 7921 5004 7955
rect 5038 7921 5044 7955
rect 4998 7883 5044 7921
rect 4998 7849 5004 7883
rect 5038 7849 5044 7883
rect 4998 7811 5044 7849
rect 4998 7777 5004 7811
rect 5038 7777 5044 7811
rect 4998 7739 5044 7777
rect 4998 7705 5004 7739
rect 5038 7705 5044 7739
rect 4998 7667 5044 7705
rect 4998 7633 5004 7667
rect 5038 7633 5044 7667
rect 4998 7595 5044 7633
rect 4998 7561 5004 7595
rect 5038 7561 5044 7595
rect 4998 7523 5044 7561
rect 4998 7489 5004 7523
rect 5038 7489 5044 7523
rect 4998 7451 5044 7489
rect 4998 7417 5004 7451
rect 5038 7417 5044 7451
rect 4998 7379 5044 7417
rect 4998 7345 5004 7379
rect 5038 7345 5044 7379
rect 4998 7307 5044 7345
rect 4998 7273 5004 7307
rect 5038 7273 5044 7307
rect 4998 7235 5044 7273
rect 4998 7201 5004 7235
rect 5038 7201 5044 7235
rect 4998 7163 5044 7201
rect 4998 7129 5004 7163
rect 5038 7129 5044 7163
rect 4998 7091 5044 7129
rect 4998 7057 5004 7091
rect 5038 7057 5044 7091
rect 4998 7019 5044 7057
rect 4998 6985 5004 7019
rect 5038 6985 5044 7019
rect 4998 6947 5044 6985
rect 4998 6913 5004 6947
rect 5038 6913 5044 6947
rect 4998 6875 5044 6913
rect 4998 6841 5004 6875
rect 5038 6841 5044 6875
rect 4998 6803 5044 6841
rect 4998 6769 5004 6803
rect 5038 6769 5044 6803
rect 4998 6731 5044 6769
rect 4998 6697 5004 6731
rect 5038 6697 5044 6731
rect 7513 8230 7519 8264
rect 7553 8230 7559 8264
rect 7513 8192 7559 8230
rect 7513 8158 7519 8192
rect 7553 8158 7559 8192
rect 7513 8120 7559 8158
rect 7513 8086 7519 8120
rect 7553 8086 7559 8120
rect 7513 8048 7559 8086
rect 7513 8014 7519 8048
rect 7553 8014 7559 8048
rect 7513 7976 7559 8014
rect 7513 7942 7519 7976
rect 7553 7942 7559 7976
rect 7513 7904 7559 7942
rect 7513 7870 7519 7904
rect 7553 7870 7559 7904
rect 7513 7832 7559 7870
rect 7513 7798 7519 7832
rect 7553 7798 7559 7832
rect 7513 7760 7559 7798
rect 7513 7726 7519 7760
rect 7553 7726 7559 7760
rect 7513 7688 7559 7726
rect 7513 7654 7519 7688
rect 7553 7654 7559 7688
rect 7513 7616 7559 7654
rect 7513 7582 7519 7616
rect 7553 7582 7559 7616
rect 7513 7544 7559 7582
rect 7513 7510 7519 7544
rect 7553 7510 7559 7544
rect 7513 7472 7559 7510
rect 7513 7438 7519 7472
rect 7553 7438 7559 7472
rect 7513 7400 7559 7438
rect 7513 7366 7519 7400
rect 7553 7366 7559 7400
rect 7513 7328 7559 7366
rect 7513 7294 7519 7328
rect 7553 7294 7559 7328
rect 7513 7256 7559 7294
rect 7513 7222 7519 7256
rect 7553 7222 7559 7256
rect 7513 7184 7559 7222
rect 7513 7150 7519 7184
rect 7553 7150 7559 7184
rect 7513 7112 7559 7150
rect 7513 7078 7519 7112
rect 7553 7078 7559 7112
rect 7513 7040 7559 7078
rect 7513 7006 7519 7040
rect 7553 7006 7559 7040
rect 7513 6968 7559 7006
rect 7513 6934 7519 6968
rect 7553 6934 7559 6968
rect 7513 6896 7559 6934
rect 7513 6862 7519 6896
rect 7553 6862 7559 6896
rect 7513 6824 7559 6862
rect 7513 6790 7519 6824
rect 7553 6790 7559 6824
rect 7513 6752 7559 6790
rect 7513 6718 7519 6752
rect 7553 6718 7559 6752
rect 4998 6659 5044 6697
rect 4998 6625 5004 6659
rect 5038 6625 5044 6659
rect 4998 6587 5044 6625
rect 4998 6553 5004 6587
rect 5038 6553 5044 6587
rect 4998 6515 5044 6553
rect 4998 6481 5004 6515
rect 5038 6481 5044 6515
rect 7044 6697 7212 6703
rect 7096 6645 7160 6697
rect 7044 6630 7212 6645
rect 7096 6578 7160 6630
rect 7044 6562 7212 6578
rect 7096 6510 7160 6562
rect 7044 6504 7212 6510
rect 7513 6680 7559 6718
rect 7513 6646 7519 6680
rect 7553 6646 7559 6680
rect 7513 6608 7559 6646
rect 7513 6574 7519 6608
rect 7553 6574 7559 6608
rect 7513 6536 7559 6574
rect 4998 6443 5044 6481
rect 4998 6409 5004 6443
rect 5038 6409 5044 6443
rect 4998 6371 5044 6409
rect 4998 6337 5004 6371
rect 5038 6337 5044 6371
rect 4998 6299 5044 6337
rect 4998 6265 5004 6299
rect 5038 6265 5044 6299
rect 4998 6227 5044 6265
rect 4656 5990 4708 6221
rect 4736 5990 4788 6221
rect 4998 6193 5004 6227
rect 5038 6193 5044 6227
rect 4998 6155 5044 6193
rect 4998 6121 5004 6155
rect 5038 6121 5044 6155
rect 4998 6083 5044 6121
rect 4998 6049 5004 6083
rect 5038 6049 5044 6083
rect 4998 6011 5044 6049
rect 4416 5434 4422 5486
rect 4474 5434 4490 5486
rect 4542 5434 4558 5486
rect 4610 5434 4616 5486
rect 2876 5361 2882 5413
rect 2934 5361 2995 5413
rect 3047 5361 3107 5413
rect 3159 5361 3165 5413
rect 2876 5323 3165 5361
rect 2876 5271 2882 5323
rect 2934 5271 2995 5323
rect 3047 5271 3107 5323
rect 3159 5271 3165 5323
rect 4416 5402 4616 5434
rect 4416 5350 4422 5402
rect 4474 5350 4490 5402
rect 4542 5350 4558 5402
rect 4610 5350 4616 5402
rect 2876 4083 2882 4135
rect 2934 4083 2995 4135
rect 3047 4083 3107 4135
rect 3159 4083 3165 4135
rect 2876 4045 3165 4083
rect 2876 3993 2882 4045
rect 2934 3993 2995 4045
rect 3047 3993 3107 4045
rect 3159 3993 3165 4045
rect 4416 4058 4616 5350
rect 4998 5977 5004 6011
rect 5038 5977 5044 6011
rect 4998 5939 5044 5977
rect 4998 5905 5004 5939
rect 5038 5905 5044 5939
rect 7513 6502 7519 6536
rect 7553 6502 7559 6536
rect 7513 6464 7559 6502
rect 7513 6430 7519 6464
rect 7553 6430 7559 6464
rect 7513 6392 7559 6430
rect 7513 6358 7519 6392
rect 7553 6358 7559 6392
rect 7513 6320 7559 6358
rect 7513 6286 7519 6320
rect 7553 6286 7559 6320
rect 7513 6248 7559 6286
rect 7513 6214 7519 6248
rect 7553 6214 7559 6248
rect 7513 6176 7559 6214
rect 7513 6142 7519 6176
rect 7553 6142 7559 6176
rect 7513 6104 7559 6142
rect 7513 6070 7519 6104
rect 7553 6070 7559 6104
rect 7513 6032 7559 6070
rect 7513 5998 7519 6032
rect 7553 5998 7559 6032
rect 7513 5960 7559 5998
rect 7513 5926 7519 5960
rect 7553 5926 7559 5960
rect 4998 5867 5044 5905
rect 4998 5833 5004 5867
rect 5038 5833 5044 5867
rect 4998 5795 5044 5833
rect 4998 5761 5004 5795
rect 5038 5761 5044 5795
rect 4998 5723 5044 5761
rect 4998 5689 5004 5723
rect 5038 5689 5044 5723
rect 7044 5910 7212 5916
rect 7096 5858 7160 5910
rect 7044 5843 7212 5858
rect 7096 5791 7160 5843
rect 7044 5775 7212 5791
rect 7096 5723 7160 5775
rect 7044 5717 7212 5723
rect 7513 5888 7559 5926
rect 7513 5854 7519 5888
rect 7553 5854 7559 5888
rect 7513 5816 7559 5854
rect 7513 5782 7519 5816
rect 7553 5782 7559 5816
rect 7513 5744 7559 5782
rect 4998 5651 5044 5689
rect 4998 5617 5004 5651
rect 5038 5617 5044 5651
rect 4998 5579 5044 5617
rect 4998 5545 5004 5579
rect 5038 5545 5044 5579
rect 4998 5507 5044 5545
rect 4998 5473 5004 5507
rect 5038 5473 5044 5507
rect 4998 5435 5044 5473
rect 4998 5401 5004 5435
rect 5038 5401 5044 5435
rect 4998 5363 5044 5401
rect 4998 5329 5004 5363
rect 5038 5329 5044 5363
rect 4998 5291 5044 5329
rect 4998 5257 5004 5291
rect 5038 5257 5044 5291
rect 4998 5219 5044 5257
rect 4998 5185 5004 5219
rect 5038 5185 5044 5219
rect 4998 5147 5044 5185
rect 4998 5113 5004 5147
rect 5038 5113 5044 5147
rect 4998 5075 5044 5113
rect 4998 5041 5004 5075
rect 5038 5041 5044 5075
rect 4998 5003 5044 5041
rect 4998 4969 5004 5003
rect 5038 4969 5044 5003
rect 4998 4931 5044 4969
rect 4998 4897 5004 4931
rect 5038 4897 5044 4931
rect 4998 4859 5044 4897
rect 7513 5710 7519 5744
rect 7553 5710 7559 5744
rect 7513 5672 7559 5710
rect 7513 5638 7519 5672
rect 7553 5638 7559 5672
rect 7513 5600 7559 5638
rect 7513 5566 7519 5600
rect 7553 5566 7559 5600
rect 7513 5528 7559 5566
rect 7513 5494 7519 5528
rect 7553 5494 7559 5528
rect 7513 5456 7559 5494
rect 7513 5422 7519 5456
rect 7553 5422 7559 5456
rect 7513 5384 7559 5422
rect 7513 5350 7519 5384
rect 7553 5350 7559 5384
rect 7513 5312 7559 5350
rect 7513 5278 7519 5312
rect 7553 5278 7559 5312
rect 7513 5240 7559 5278
rect 7513 5206 7519 5240
rect 7553 5206 7559 5240
rect 7513 5168 7559 5206
rect 7513 5134 7519 5168
rect 7553 5134 7559 5168
rect 7513 5096 7559 5134
rect 7513 5062 7519 5096
rect 7553 5062 7559 5096
rect 7513 5024 7559 5062
rect 7513 4990 7519 5024
rect 7553 4990 7559 5024
rect 7513 4952 7559 4990
rect 7513 4918 7519 4952
rect 7553 4918 7559 4952
rect 7513 4880 7559 4918
rect 4998 4825 5004 4859
rect 5038 4825 5044 4859
rect 4656 4557 4708 4788
rect 4736 4557 4788 4788
rect 4998 4787 5044 4825
rect 4998 4753 5004 4787
rect 5038 4753 5044 4787
rect 4998 4715 5044 4753
rect 4998 4681 5004 4715
rect 5038 4681 5044 4715
rect 4998 4643 5044 4681
rect 7044 4861 7212 4867
rect 7096 4809 7160 4861
rect 7044 4794 7212 4809
rect 7096 4742 7160 4794
rect 7044 4726 7212 4742
rect 7096 4674 7160 4726
rect 7044 4668 7212 4674
rect 7513 4846 7519 4880
rect 7553 4846 7559 4880
rect 7513 4808 7559 4846
rect 7513 4774 7519 4808
rect 7553 4774 7559 4808
rect 7513 4736 7559 4774
rect 7513 4702 7519 4736
rect 7553 4702 7559 4736
rect 4998 4609 5004 4643
rect 5038 4609 5044 4643
rect 4998 4571 5044 4609
rect 4416 4006 4422 4058
rect 4474 4006 4490 4058
rect 4542 4006 4558 4058
rect 4610 4006 4616 4058
rect 4416 3974 4616 4006
rect 4416 3922 4422 3974
rect 4474 3922 4490 3974
rect 4542 3922 4558 3974
rect 4610 3922 4616 3974
rect 2917 3383 3024 3387
rect 2917 3368 3043 3383
tri 3043 3368 3058 3383 nw
rect 2917 3311 3024 3368
tri 3024 3349 3043 3368 nw
rect 2917 3259 2944 3311
rect 2996 3259 3024 3311
rect 2917 3243 3024 3259
rect 2917 3191 2944 3243
rect 2996 3191 3024 3243
rect 2917 3175 3024 3191
rect 2917 3123 2944 3175
rect 2996 3123 3024 3175
rect 2917 3117 3024 3123
rect 3877 3311 4077 3463
rect 3929 3259 3951 3311
rect 4003 3259 4025 3311
rect 3877 3243 4077 3259
rect 3929 3191 3951 3243
rect 4003 3191 4025 3243
rect 3877 3175 4077 3191
rect 3929 3123 3951 3175
rect 4003 3123 4025 3175
rect 3877 3117 4077 3123
rect 4416 3316 4616 3922
rect 4998 4537 5004 4571
rect 5038 4537 5044 4571
rect 4998 4499 5044 4537
rect 4998 4465 5004 4499
rect 5038 4465 5044 4499
rect 4998 4427 5044 4465
rect 4998 4393 5004 4427
rect 5038 4393 5044 4427
rect 4998 4355 5044 4393
rect 4998 4321 5004 4355
rect 5038 4321 5044 4355
rect 4998 4283 5044 4321
rect 4998 4249 5004 4283
rect 5038 4249 5044 4283
rect 4998 4211 5044 4249
rect 4998 4177 5004 4211
rect 5038 4177 5044 4211
rect 4998 4139 5044 4177
rect 4998 4105 5004 4139
rect 5038 4105 5044 4139
rect 4998 4067 5044 4105
rect 4998 4033 5004 4067
rect 5038 4033 5044 4067
rect 4998 3995 5044 4033
rect 4998 3961 5004 3995
rect 5038 3961 5044 3995
rect 4998 3923 5044 3961
rect 4998 3889 5004 3923
rect 5038 3889 5044 3923
rect 4998 3851 5044 3889
rect 4998 3817 5004 3851
rect 5038 3817 5044 3851
rect 4998 3779 5044 3817
rect 4998 3745 5004 3779
rect 5038 3745 5044 3779
rect 4998 3707 5044 3745
rect 7513 4664 7559 4702
rect 7513 4630 7519 4664
rect 7553 4630 7559 4664
rect 7513 4592 7559 4630
rect 7513 4558 7519 4592
rect 7553 4558 7559 4592
rect 7513 4520 7559 4558
rect 7513 4486 7519 4520
rect 7553 4486 7559 4520
rect 7513 4448 7559 4486
rect 7513 4414 7519 4448
rect 7553 4414 7559 4448
rect 7513 4376 7559 4414
rect 7513 4342 7519 4376
rect 7553 4342 7559 4376
rect 7513 4304 7559 4342
rect 7513 4270 7519 4304
rect 7553 4270 7559 4304
rect 7513 4232 7559 4270
rect 7513 4198 7519 4232
rect 7553 4198 7559 4232
rect 7513 4160 7559 4198
rect 7513 4126 7519 4160
rect 7553 4126 7559 4160
rect 7513 4088 7559 4126
rect 7513 4054 7519 4088
rect 7553 4054 7559 4088
rect 7513 4016 7559 4054
rect 7513 3982 7519 4016
rect 7553 3982 7559 4016
rect 7513 3944 7559 3982
rect 7513 3910 7519 3944
rect 7553 3910 7559 3944
rect 7513 3872 7559 3910
rect 7513 3838 7519 3872
rect 7553 3838 7559 3872
rect 7513 3800 7559 3838
rect 7513 3766 7519 3800
rect 7553 3766 7559 3800
rect 4998 3673 5004 3707
rect 5038 3673 5044 3707
rect 4998 3635 5044 3673
rect 4998 3601 5004 3635
rect 5038 3601 5044 3635
rect 4998 3563 5044 3601
rect 4998 3529 5004 3563
rect 5038 3529 5044 3563
rect 7044 3725 7212 3731
rect 7096 3673 7160 3725
rect 7044 3658 7212 3673
rect 7096 3606 7160 3658
rect 7044 3590 7212 3606
rect 7096 3538 7160 3590
rect 7044 3532 7212 3538
rect 7513 3728 7559 3766
rect 7513 3694 7519 3728
rect 7553 3694 7559 3728
rect 7513 3656 7559 3694
rect 7513 3622 7519 3656
rect 7553 3622 7559 3656
rect 7513 3584 7559 3622
rect 7513 3550 7519 3584
rect 7553 3550 7559 3584
rect 4998 3491 5044 3529
rect 4998 3457 5004 3491
rect 5038 3457 5044 3491
rect 4998 3419 5044 3457
rect 4468 3264 4490 3316
rect 4542 3264 4564 3316
rect 4416 3188 4616 3264
rect 4468 3136 4490 3188
rect 4542 3136 4564 3188
rect 4416 3060 4616 3136
rect 4468 3008 4490 3060
rect 4542 3008 4564 3060
rect 4416 2932 4616 3008
rect 4468 2880 4490 2932
rect 4542 2880 4564 2932
rect 4656 3044 4708 3408
rect 4736 3281 4788 3408
rect 4736 3217 4788 3229
rect 4736 3159 4788 3165
rect 4998 3385 5004 3419
rect 5038 3385 5044 3419
rect 4998 3347 5044 3385
rect 4998 3313 5004 3347
rect 5038 3313 5044 3347
rect 4998 3275 5044 3313
rect 4998 3241 5004 3275
rect 5038 3241 5044 3275
rect 4998 3203 5044 3241
rect 7513 3512 7559 3550
rect 7513 3478 7519 3512
rect 7553 3478 7559 3512
rect 7513 3440 7559 3478
rect 7513 3406 7519 3440
rect 7553 3406 7559 3440
rect 7513 3368 7559 3406
rect 7513 3334 7519 3368
rect 7553 3334 7559 3368
rect 7513 3295 7559 3334
rect 7513 3261 7519 3295
rect 7553 3261 7559 3295
rect 7513 3222 7559 3261
rect 4998 3169 5004 3203
rect 5038 3169 5044 3203
rect 4656 2980 4708 2992
rect 4656 2922 4708 2928
rect 4998 3131 5044 3169
rect 4998 3097 5004 3131
rect 5038 3097 5044 3131
rect 4998 3059 5044 3097
rect 4998 3025 5004 3059
rect 5038 3025 5044 3059
rect 4998 2987 5044 3025
rect 7044 3215 7212 3221
rect 7096 3163 7160 3215
rect 7044 3148 7212 3163
rect 7096 3096 7160 3148
rect 7044 3080 7212 3096
rect 7096 3028 7160 3080
rect 7044 3022 7212 3028
rect 7513 3188 7519 3222
rect 7553 3188 7559 3222
rect 7513 3149 7559 3188
rect 7513 3115 7519 3149
rect 7553 3115 7559 3149
rect 7513 3076 7559 3115
rect 7513 3042 7519 3076
rect 7553 3042 7559 3076
rect 7513 3003 7559 3042
rect 4998 2953 5004 2987
rect 5038 2953 5044 2987
rect 4416 2804 4616 2880
rect 4468 2752 4490 2804
rect 4542 2752 4564 2804
rect 4416 2676 4616 2752
rect 4468 2624 4490 2676
rect 4542 2624 4564 2676
rect 4416 2547 4616 2624
rect 4468 2495 4490 2547
rect 4542 2495 4564 2547
rect 4416 2418 4616 2495
rect 4468 2366 4490 2418
rect 4542 2366 4564 2418
rect 4416 2360 4616 2366
rect 4998 2915 5044 2953
rect 4998 2881 5004 2915
rect 5038 2881 5044 2915
rect 4998 2843 5044 2881
rect 6079 2988 6131 2994
rect 6079 2924 6131 2936
rect 4998 2809 5004 2843
rect 5038 2809 5044 2843
rect 6076 2872 6079 2880
rect 4998 2771 5044 2809
rect 4998 2737 5004 2771
rect 5038 2737 5044 2771
rect 4998 2699 5044 2737
rect 5989 2827 6041 2833
rect 5989 2763 6041 2775
rect 5989 2705 6041 2711
rect 4998 2665 5004 2699
rect 5038 2665 5044 2699
rect 4998 2627 5044 2665
rect 4998 2593 5004 2627
rect 5038 2593 5044 2627
rect 4998 2555 5044 2593
rect 4998 2521 5004 2555
rect 5038 2521 5044 2555
rect 4998 2483 5044 2521
rect 4998 2449 5004 2483
rect 5038 2449 5044 2483
rect 4998 2411 5044 2449
rect 4998 2377 5004 2411
rect 5038 2377 5044 2411
rect 4998 2339 5044 2377
rect 4998 2305 5004 2339
rect 5038 2305 5044 2339
rect 4998 2267 5044 2305
rect 4998 2233 5004 2267
rect 5038 2233 5044 2267
tri 4985 2210 4998 2223 se
rect 4998 2210 5044 2233
rect 6076 2232 6131 2872
rect 7513 2969 7519 3003
rect 7553 2969 7559 3003
rect 7513 2930 7559 2969
rect 7513 2896 7519 2930
rect 7553 2896 7559 2930
rect 7513 2857 7559 2896
rect 6278 2825 6330 2833
rect 6278 2761 6330 2773
rect 6278 2363 6330 2709
rect 7158 2825 7210 2833
rect 7158 2761 7210 2773
rect 7158 2703 7210 2709
rect 7513 2823 7519 2857
rect 7553 2823 7559 2857
rect 7513 2784 7559 2823
rect 7513 2750 7519 2784
rect 7553 2750 7559 2784
rect 7513 2711 7559 2750
rect 6278 2299 6330 2311
rect 6278 2241 6330 2247
rect 7513 2677 7519 2711
rect 7553 2677 7559 2711
rect 7513 2638 7559 2677
rect 7513 2604 7519 2638
rect 7553 2604 7559 2638
rect 7513 2565 7559 2604
rect 7513 2531 7519 2565
rect 7553 2531 7559 2565
rect 7513 2492 7559 2531
rect 7513 2458 7519 2492
rect 7553 2458 7559 2492
rect 7513 2419 7559 2458
rect 7513 2385 7519 2419
rect 7553 2385 7559 2419
rect 7513 2346 7559 2385
rect 7513 2312 7519 2346
rect 7553 2312 7559 2346
rect 7513 2273 7559 2312
rect 7513 2239 7519 2273
rect 7553 2239 7559 2273
tri 5044 2210 5057 2223 sw
tri 5277 2210 5290 2223 se
tri 4975 2200 4985 2210 se
rect 4985 2200 5057 2210
tri 5057 2200 5067 2210 sw
tri 5267 2200 5277 2210 se
rect 5277 2200 5290 2210
tri 4970 2195 4975 2200 se
rect 4975 2195 5067 2200
tri 4964 2189 4970 2195 se
rect 4970 2189 5004 2195
rect 3471 2188 5004 2189
rect 3471 2136 3477 2188
rect 3529 2136 3586 2188
rect 3638 2136 3695 2188
rect 3747 2136 3803 2188
rect 3855 2136 3911 2188
rect 3963 2136 4019 2188
rect 4071 2161 5004 2188
rect 5038 2189 5067 2195
tri 5067 2189 5078 2200 sw
tri 5256 2189 5267 2200 se
rect 5267 2189 5290 2200
rect 7513 2200 7559 2239
rect 5038 2161 5305 2189
rect 4071 2136 5305 2161
rect 3471 2123 5305 2136
rect 3471 2106 5004 2123
rect 3471 2054 3477 2106
rect 3529 2054 3586 2106
rect 3638 2054 3695 2106
rect 3747 2054 3803 2106
rect 3855 2054 3911 2106
rect 3963 2054 4019 2106
rect 4071 2089 5004 2106
rect 5038 2089 5305 2123
rect 4071 2054 5305 2089
rect 3471 2051 5305 2054
rect 3471 2024 5004 2051
rect 3471 1972 3477 2024
rect 3529 1972 3586 2024
rect 3638 1972 3695 2024
rect 3747 1972 3803 2024
rect 3855 1972 3911 2024
rect 3963 1972 4019 2024
rect 4071 2017 5004 2024
rect 5038 2017 5305 2051
rect 4071 1979 5305 2017
rect 4071 1972 5004 1979
rect 3471 1945 5004 1972
rect 5038 1945 5305 1979
rect 3471 1942 5305 1945
rect 3471 1890 3477 1942
rect 3529 1890 3586 1942
rect 3638 1890 3695 1942
rect 3747 1890 3803 1942
rect 3855 1890 3911 1942
rect 3963 1890 4019 1942
rect 4071 1907 5305 1942
rect 4071 1890 5004 1907
rect 3471 1889 5004 1890
tri 4964 1873 4980 1889 ne
rect 4980 1873 5004 1889
rect 5038 1889 5305 1907
rect 7513 2166 7519 2200
rect 7553 2166 7559 2200
rect 7513 2127 7559 2166
rect 7513 2093 7519 2127
rect 7553 2093 7559 2127
rect 7513 2054 7559 2093
rect 7513 2020 7519 2054
rect 7553 2020 7559 2054
rect 7513 1981 7559 2020
rect 7513 1947 7519 1981
rect 7553 1947 7559 1981
rect 7513 1908 7559 1947
rect 5038 1874 5063 1889
tri 5063 1874 5078 1889 nw
rect 7513 1874 7519 1908
rect 7553 1874 7559 1908
rect 5038 1873 5044 1874
tri 4980 1855 4998 1873 ne
rect 4998 1835 5044 1873
tri 5044 1855 5063 1874 nw
rect 4998 1801 5004 1835
rect 5038 1801 5044 1835
rect 7513 1835 7559 1874
tri 5044 1801 5046 1803 sw
tri 7511 1801 7513 1803 se
rect 7513 1801 7519 1835
rect 7553 1801 7559 1835
rect 4998 1772 5046 1801
tri 5046 1772 5075 1801 sw
tri 7482 1772 7511 1801 se
rect 7511 1772 7559 1801
rect 4998 1769 5075 1772
tri 5075 1769 5078 1772 sw
tri 7479 1769 7482 1772 se
rect 7482 1769 7559 1772
rect 4998 1763 7559 1769
rect 4998 1729 5076 1763
rect 5110 1729 5151 1763
rect 5185 1729 5225 1763
rect 5259 1729 5299 1763
rect 5333 1729 5373 1763
rect 5407 1729 5447 1763
rect 5481 1729 5521 1763
rect 5555 1729 5595 1763
rect 5629 1729 5669 1763
rect 5703 1729 5743 1763
rect 5777 1729 5817 1763
rect 5851 1729 5891 1763
rect 5925 1729 5965 1763
rect 5999 1729 6039 1763
rect 6073 1729 6113 1763
rect 6147 1729 6187 1763
rect 6221 1729 6261 1763
rect 6295 1729 6335 1763
rect 6369 1729 6409 1763
rect 6443 1729 6483 1763
rect 6517 1729 6557 1763
rect 6591 1729 6631 1763
rect 6665 1729 6705 1763
rect 6739 1729 6779 1763
rect 6813 1729 6853 1763
rect 6887 1729 6927 1763
rect 6961 1729 7001 1763
rect 7035 1729 7075 1763
rect 7109 1729 7149 1763
rect 7183 1729 7223 1763
rect 7257 1729 7297 1763
rect 7331 1729 7371 1763
rect 7405 1729 7445 1763
rect 7479 1729 7559 1763
rect 4998 1723 7559 1729
rect 7870 2395 7876 17549
rect 9278 2395 9284 17549
rect 7870 2356 9284 2395
rect 7870 2322 7876 2356
rect 7910 2322 7948 2356
rect 7982 2322 8020 2356
rect 8054 2322 8092 2356
rect 8126 2322 8164 2356
rect 8198 2322 8236 2356
rect 8270 2322 8308 2356
rect 8342 2322 8380 2356
rect 8414 2322 8452 2356
rect 8486 2322 8524 2356
rect 8558 2322 8596 2356
rect 8630 2322 8668 2356
rect 8702 2322 8740 2356
rect 8774 2322 8812 2356
rect 8846 2322 8884 2356
rect 8918 2322 8956 2356
rect 8990 2322 9028 2356
rect 9062 2322 9100 2356
rect 9134 2322 9172 2356
rect 9206 2322 9244 2356
rect 9278 2322 9284 2356
rect 7870 2283 9284 2322
rect 7870 2249 7876 2283
rect 7910 2249 7948 2283
rect 7982 2249 8020 2283
rect 8054 2249 8092 2283
rect 8126 2249 8164 2283
rect 8198 2249 8236 2283
rect 8270 2249 8308 2283
rect 8342 2249 8380 2283
rect 8414 2249 8452 2283
rect 8486 2249 8524 2283
rect 8558 2249 8596 2283
rect 8630 2249 8668 2283
rect 8702 2249 8740 2283
rect 8774 2249 8812 2283
rect 8846 2249 8884 2283
rect 8918 2249 8956 2283
rect 8990 2249 9028 2283
rect 9062 2249 9100 2283
rect 9134 2249 9172 2283
rect 9206 2249 9244 2283
rect 9278 2249 9284 2283
rect 7870 2210 9284 2249
rect 7870 2176 7876 2210
rect 7910 2176 7948 2210
rect 7982 2176 8020 2210
rect 8054 2176 8092 2210
rect 8126 2176 8164 2210
rect 8198 2176 8236 2210
rect 8270 2176 8308 2210
rect 8342 2176 8380 2210
rect 8414 2176 8452 2210
rect 8486 2176 8524 2210
rect 8558 2176 8596 2210
rect 8630 2176 8668 2210
rect 8702 2176 8740 2210
rect 8774 2176 8812 2210
rect 8846 2176 8884 2210
rect 8918 2176 8956 2210
rect 8990 2176 9028 2210
rect 9062 2176 9100 2210
rect 9134 2176 9172 2210
rect 9206 2176 9244 2210
rect 9278 2176 9284 2210
rect 7870 2137 9284 2176
rect 7870 2103 7876 2137
rect 7910 2103 7948 2137
rect 7982 2103 8020 2137
rect 8054 2103 8092 2137
rect 8126 2103 8164 2137
rect 8198 2103 8236 2137
rect 8270 2103 8308 2137
rect 8342 2103 8380 2137
rect 8414 2103 8452 2137
rect 8486 2103 8524 2137
rect 8558 2103 8596 2137
rect 8630 2103 8668 2137
rect 8702 2103 8740 2137
rect 8774 2103 8812 2137
rect 8846 2103 8884 2137
rect 8918 2103 8956 2137
rect 8990 2103 9028 2137
rect 9062 2103 9100 2137
rect 9134 2103 9172 2137
rect 9206 2103 9244 2137
rect 9278 2103 9284 2137
rect 7870 2064 9284 2103
rect 7870 2030 7876 2064
rect 7910 2030 7948 2064
rect 7982 2030 8020 2064
rect 8054 2030 8092 2064
rect 8126 2030 8164 2064
rect 8198 2030 8236 2064
rect 8270 2030 8308 2064
rect 8342 2030 8380 2064
rect 8414 2030 8452 2064
rect 8486 2030 8524 2064
rect 8558 2030 8596 2064
rect 8630 2030 8668 2064
rect 8702 2030 8740 2064
rect 8774 2030 8812 2064
rect 8846 2030 8884 2064
rect 8918 2030 8956 2064
rect 8990 2030 9028 2064
rect 9062 2030 9100 2064
rect 9134 2030 9172 2064
rect 9206 2030 9244 2064
rect 9278 2030 9284 2064
rect 7870 1991 9284 2030
rect 7870 1957 7876 1991
rect 7910 1957 7948 1991
rect 7982 1957 8020 1991
rect 8054 1957 8092 1991
rect 8126 1957 8164 1991
rect 8198 1957 8236 1991
rect 8270 1957 8308 1991
rect 8342 1957 8380 1991
rect 8414 1957 8452 1991
rect 8486 1957 8524 1991
rect 8558 1957 8596 1991
rect 8630 1957 8668 1991
rect 8702 1957 8740 1991
rect 8774 1957 8812 1991
rect 8846 1957 8884 1991
rect 8918 1957 8956 1991
rect 8990 1957 9028 1991
rect 9062 1957 9100 1991
rect 9134 1957 9172 1991
rect 9206 1957 9244 1991
rect 9278 1957 9284 1991
rect 7870 1918 9284 1957
rect 7870 1884 7876 1918
rect 7910 1884 7948 1918
rect 7982 1884 8020 1918
rect 8054 1884 8092 1918
rect 8126 1884 8164 1918
rect 8198 1884 8236 1918
rect 8270 1884 8308 1918
rect 8342 1884 8380 1918
rect 8414 1884 8452 1918
rect 8486 1884 8524 1918
rect 8558 1884 8596 1918
rect 8630 1884 8668 1918
rect 8702 1884 8740 1918
rect 8774 1884 8812 1918
rect 8846 1884 8884 1918
rect 8918 1884 8956 1918
rect 8990 1884 9028 1918
rect 9062 1884 9100 1918
rect 9134 1884 9172 1918
rect 9206 1884 9244 1918
rect 9278 1884 9284 1918
rect 7870 1845 9284 1884
rect 7870 1811 7876 1845
rect 7910 1811 7948 1845
rect 7982 1811 8020 1845
rect 8054 1811 8092 1845
rect 8126 1811 8164 1845
rect 8198 1811 8236 1845
rect 8270 1811 8308 1845
rect 8342 1811 8380 1845
rect 8414 1811 8452 1845
rect 8486 1811 8524 1845
rect 8558 1811 8596 1845
rect 8630 1811 8668 1845
rect 8702 1811 8740 1845
rect 8774 1811 8812 1845
rect 8846 1811 8884 1845
rect 8918 1811 8956 1845
rect 8990 1811 9028 1845
rect 9062 1811 9100 1845
rect 9134 1811 9172 1845
rect 9206 1811 9244 1845
rect 9278 1811 9284 1845
rect 7870 1772 9284 1811
rect 7870 1738 7876 1772
rect 7910 1738 7948 1772
rect 7982 1738 8020 1772
rect 8054 1738 8092 1772
rect 8126 1738 8164 1772
rect 8198 1738 8236 1772
rect 8270 1738 8308 1772
rect 8342 1738 8380 1772
rect 8414 1738 8452 1772
rect 8486 1738 8524 1772
rect 8558 1738 8596 1772
rect 8630 1738 8668 1772
rect 8702 1738 8740 1772
rect 8774 1738 8812 1772
rect 8846 1738 8884 1772
rect 8918 1738 8956 1772
rect 8990 1738 9028 1772
rect 9062 1738 9100 1772
rect 9134 1738 9172 1772
rect 9206 1738 9244 1772
rect 9278 1738 9284 1772
rect 7870 1699 9284 1738
rect 7870 1665 7876 1699
rect 7910 1665 7948 1699
rect 7982 1665 8020 1699
rect 8054 1665 8092 1699
rect 8126 1665 8164 1699
rect 8198 1665 8236 1699
rect 8270 1665 8308 1699
rect 8342 1665 8380 1699
rect 8414 1665 8452 1699
rect 8486 1665 8524 1699
rect 8558 1665 8596 1699
rect 8630 1665 8668 1699
rect 8702 1665 8740 1699
rect 8774 1665 8812 1699
rect 8846 1665 8884 1699
rect 8918 1665 8956 1699
rect 8990 1665 9028 1699
rect 9062 1665 9100 1699
rect 9134 1665 9172 1699
rect 9206 1665 9244 1699
rect 9278 1665 9284 1699
rect 7870 1626 9284 1665
rect 7870 1592 7876 1626
rect 7910 1592 7948 1626
rect 7982 1592 8020 1626
rect 8054 1592 8092 1626
rect 8126 1592 8164 1626
rect 8198 1592 8236 1626
rect 8270 1592 8308 1626
rect 8342 1592 8380 1626
rect 8414 1592 8452 1626
rect 8486 1592 8524 1626
rect 8558 1592 8596 1626
rect 8630 1592 8668 1626
rect 8702 1592 8740 1626
rect 8774 1592 8812 1626
rect 8846 1592 8884 1626
rect 8918 1592 8956 1626
rect 8990 1592 9028 1626
rect 9062 1592 9100 1626
rect 9134 1592 9172 1626
rect 9206 1592 9244 1626
rect 9278 1592 9284 1626
rect 7870 1553 9284 1592
rect 7870 1519 7876 1553
rect 7910 1519 7948 1553
rect 7982 1519 8020 1553
rect 8054 1519 8092 1553
rect 8126 1519 8164 1553
rect 8198 1519 8236 1553
rect 8270 1519 8308 1553
rect 8342 1519 8380 1553
rect 8414 1519 8452 1553
rect 8486 1519 8524 1553
rect 8558 1519 8596 1553
rect 8630 1519 8668 1553
rect 8702 1519 8740 1553
rect 8774 1519 8812 1553
rect 8846 1519 8884 1553
rect 8918 1519 8956 1553
rect 8990 1519 9028 1553
rect 9062 1519 9100 1553
rect 9134 1519 9172 1553
rect 9206 1519 9244 1553
rect 9278 1519 9284 1553
rect 7870 1480 9284 1519
rect 7870 1446 7876 1480
rect 7910 1446 7948 1480
rect 7982 1446 8020 1480
rect 8054 1446 8092 1480
rect 8126 1446 8164 1480
rect 8198 1446 8236 1480
rect 8270 1446 8308 1480
rect 8342 1446 8380 1480
rect 8414 1446 8452 1480
rect 8486 1446 8524 1480
rect 8558 1446 8596 1480
rect 8630 1446 8668 1480
rect 8702 1446 8740 1480
rect 8774 1446 8812 1480
rect 8846 1446 8884 1480
rect 8918 1446 8956 1480
rect 8990 1446 9028 1480
rect 9062 1446 9100 1480
rect 9134 1446 9172 1480
rect 9206 1446 9244 1480
rect 9278 1446 9284 1480
rect 7870 1407 9284 1446
rect 7870 1373 7876 1407
rect 7910 1373 7948 1407
rect 7982 1373 8020 1407
rect 8054 1373 8092 1407
rect 8126 1373 8164 1407
rect 8198 1373 8236 1407
rect 8270 1373 8308 1407
rect 8342 1373 8380 1407
rect 8414 1373 8452 1407
rect 8486 1373 8524 1407
rect 8558 1373 8596 1407
rect 8630 1373 8668 1407
rect 8702 1373 8740 1407
rect 8774 1373 8812 1407
rect 8846 1373 8884 1407
rect 8918 1373 8956 1407
rect 8990 1373 9028 1407
rect 9062 1373 9100 1407
rect 9134 1373 9172 1407
rect 9206 1373 9244 1407
rect 9278 1373 9284 1407
rect 7870 1334 9284 1373
rect 7870 1300 7876 1334
rect 7910 1300 7948 1334
rect 7982 1300 8020 1334
rect 8054 1300 8092 1334
rect 8126 1300 8164 1334
rect 8198 1300 8236 1334
rect 8270 1300 8308 1334
rect 8342 1300 8380 1334
rect 8414 1300 8452 1334
rect 8486 1300 8524 1334
rect 8558 1300 8596 1334
rect 8630 1300 8668 1334
rect 8702 1300 8740 1334
rect 8774 1300 8812 1334
rect 8846 1300 8884 1334
rect 8918 1300 8956 1334
rect 8990 1300 9028 1334
rect 9062 1300 9100 1334
rect 9134 1300 9172 1334
rect 9206 1300 9244 1334
rect 9278 1300 9284 1334
rect 7870 1261 9284 1300
rect 7870 1227 7876 1261
rect 7910 1227 7948 1261
rect 7982 1227 8020 1261
rect 8054 1227 8092 1261
rect 8126 1227 8164 1261
rect 8198 1227 8236 1261
rect 8270 1227 8308 1261
rect 8342 1227 8380 1261
rect 8414 1227 8452 1261
rect 8486 1227 8524 1261
rect 8558 1227 8596 1261
rect 8630 1227 8668 1261
rect 8702 1227 8740 1261
rect 8774 1227 8812 1261
rect 8846 1227 8884 1261
rect 8918 1227 8956 1261
rect 8990 1227 9028 1261
rect 9062 1227 9100 1261
rect 9134 1227 9172 1261
rect 9206 1227 9244 1261
rect 9278 1227 9284 1261
rect 7870 1188 9284 1227
rect 7870 1154 7876 1188
rect 7910 1154 7948 1188
rect 7982 1154 8020 1188
rect 8054 1154 8092 1188
rect 8126 1154 8164 1188
rect 8198 1154 8236 1188
rect 8270 1154 8308 1188
rect 8342 1154 8380 1188
rect 8414 1154 8452 1188
rect 8486 1154 8524 1188
rect 8558 1154 8596 1188
rect 8630 1154 8668 1188
rect 8702 1154 8740 1188
rect 8774 1154 8812 1188
rect 8846 1154 8884 1188
rect 8918 1154 8956 1188
rect 8990 1154 9028 1188
rect 9062 1154 9100 1188
rect 9134 1154 9172 1188
rect 9206 1154 9244 1188
rect 9278 1154 9284 1188
rect 7870 1115 9284 1154
rect 7870 1081 7876 1115
rect 7910 1081 7948 1115
rect 7982 1081 8020 1115
rect 8054 1081 8092 1115
rect 8126 1081 8164 1115
rect 8198 1081 8236 1115
rect 8270 1081 8308 1115
rect 8342 1081 8380 1115
rect 8414 1081 8452 1115
rect 8486 1081 8524 1115
rect 8558 1081 8596 1115
rect 8630 1081 8668 1115
rect 8702 1081 8740 1115
rect 8774 1081 8812 1115
rect 8846 1081 8884 1115
rect 8918 1081 8956 1115
rect 8990 1081 9028 1115
rect 9062 1081 9100 1115
rect 9134 1081 9172 1115
rect 9206 1081 9244 1115
rect 9278 1081 9284 1115
rect 7870 1042 9284 1081
rect 7870 1008 7876 1042
rect 7910 1008 7948 1042
rect 7982 1008 8020 1042
rect 8054 1008 8092 1042
rect 8126 1008 8164 1042
rect 8198 1008 8236 1042
rect 8270 1008 8308 1042
rect 8342 1008 8380 1042
rect 8414 1008 8452 1042
rect 8486 1008 8524 1042
rect 8558 1008 8596 1042
rect 8630 1008 8668 1042
rect 8702 1008 8740 1042
rect 8774 1008 8812 1042
rect 8846 1008 8884 1042
rect 8918 1008 8956 1042
rect 8990 1008 9028 1042
rect 9062 1008 9100 1042
rect 9134 1008 9172 1042
rect 9206 1008 9244 1042
rect 9278 1008 9284 1042
rect 7870 969 9284 1008
rect 7870 935 7876 969
rect 7910 935 7948 969
rect 7982 935 8020 969
rect 8054 935 8092 969
rect 8126 935 8164 969
rect 8198 935 8236 969
rect 8270 935 8308 969
rect 8342 935 8380 969
rect 8414 935 8452 969
rect 8486 935 8524 969
rect 8558 935 8596 969
rect 8630 935 8668 969
rect 8702 935 8740 969
rect 8774 935 8812 969
rect 8846 935 8884 969
rect 8918 935 8956 969
rect 8990 935 9028 969
rect 9062 935 9100 969
rect 9134 935 9172 969
rect 9206 935 9244 969
rect 9278 935 9284 969
rect 7870 896 9284 935
rect 7870 862 7876 896
rect 7910 862 7948 896
rect 7982 862 8020 896
rect 8054 862 8092 896
rect 8126 862 8164 896
rect 8198 862 8236 896
rect 8270 862 8308 896
rect 8342 862 8380 896
rect 8414 862 8452 896
rect 8486 862 8524 896
rect 8558 862 8596 896
rect 8630 862 8668 896
rect 8702 862 8740 896
rect 8774 862 8812 896
rect 8846 862 8884 896
rect 8918 862 8956 896
rect 8990 862 9028 896
rect 9062 862 9100 896
rect 9134 862 9172 896
rect 9206 862 9244 896
rect 9278 862 9284 896
rect 7870 823 9284 862
rect 7870 789 7876 823
rect 7910 789 7948 823
rect 7982 789 8020 823
rect 8054 789 8092 823
rect 8126 789 8164 823
rect 8198 789 8236 823
rect 8270 789 8308 823
rect 8342 789 8380 823
rect 8414 789 8452 823
rect 8486 789 8524 823
rect 8558 789 8596 823
rect 8630 789 8668 823
rect 8702 789 8740 823
rect 8774 789 8812 823
rect 8846 789 8884 823
rect 8918 789 8956 823
rect 8990 789 9028 823
rect 9062 789 9100 823
rect 9134 789 9172 823
rect 9206 789 9244 823
rect 9278 789 9284 823
rect 7870 750 9284 789
rect 7870 716 7876 750
rect 7910 716 7948 750
rect 7982 716 8020 750
rect 8054 716 8092 750
rect 8126 716 8164 750
rect 8198 716 8236 750
rect 8270 716 8308 750
rect 8342 716 8380 750
rect 8414 716 8452 750
rect 8486 716 8524 750
rect 8558 716 8596 750
rect 8630 716 8668 750
rect 8702 716 8740 750
rect 8774 716 8812 750
rect 8846 716 8884 750
rect 8918 716 8956 750
rect 8990 716 9028 750
rect 9062 716 9100 750
rect 9134 716 9172 750
rect 9206 716 9244 750
rect 9278 716 9284 750
rect 7870 677 9284 716
rect 7870 643 7876 677
rect 7910 643 7948 677
rect 7982 643 8020 677
rect 8054 643 8092 677
rect 8126 643 8164 677
rect 8198 643 8236 677
rect 8270 643 8308 677
rect 8342 643 8380 677
rect 8414 643 8452 677
rect 8486 643 8524 677
rect 8558 643 8596 677
rect 8630 643 8668 677
rect 8702 643 8740 677
rect 8774 643 8812 677
rect 8846 643 8884 677
rect 8918 643 8956 677
rect 8990 643 9028 677
rect 9062 643 9100 677
rect 9134 643 9172 677
rect 9206 643 9244 677
rect 9278 643 9284 677
rect 7870 604 9284 643
rect 7870 570 7876 604
rect 7910 570 7948 604
rect 7982 570 8020 604
rect 8054 570 8092 604
rect 8126 570 8164 604
rect 8198 570 8236 604
rect 8270 570 8308 604
rect 8342 570 8380 604
rect 8414 570 8452 604
rect 8486 570 8524 604
rect 8558 570 8596 604
rect 8630 570 8668 604
rect 8702 570 8740 604
rect 8774 570 8812 604
rect 8846 570 8884 604
rect 8918 570 8956 604
rect 8990 570 9028 604
rect 9062 570 9100 604
rect 9134 570 9172 604
rect 9206 570 9244 604
rect 9278 570 9284 604
rect 7870 531 9284 570
rect 7870 497 7876 531
rect 7910 497 7948 531
rect 7982 497 8020 531
rect 8054 497 8092 531
rect 8126 497 8164 531
rect 8198 497 8236 531
rect 8270 497 8308 531
rect 8342 497 8380 531
rect 8414 497 8452 531
rect 8486 497 8524 531
rect 8558 497 8596 531
rect 8630 497 8668 531
rect 8702 497 8740 531
rect 8774 497 8812 531
rect 8846 497 8884 531
rect 8918 497 8956 531
rect 8990 497 9028 531
rect 9062 497 9100 531
rect 9134 497 9172 531
rect 9206 497 9244 531
rect 9278 497 9284 531
rect 7870 458 9284 497
rect 7870 424 7876 458
rect 7910 424 7948 458
rect 7982 424 8020 458
rect 8054 424 8092 458
rect 8126 424 8164 458
rect 8198 424 8236 458
rect 8270 424 8308 458
rect 8342 424 8380 458
rect 8414 424 8452 458
rect 8486 424 8524 458
rect 8558 424 8596 458
rect 8630 424 8668 458
rect 8702 424 8740 458
rect 8774 424 8812 458
rect 8846 424 8884 458
rect 8918 424 8956 458
rect 8990 424 9028 458
rect 9062 424 9100 458
rect 9134 424 9172 458
rect 9206 424 9244 458
rect 9278 424 9284 458
rect 7870 385 9284 424
rect 7870 351 7876 385
rect 7910 351 7948 385
rect 7982 351 8020 385
rect 8054 351 8092 385
rect 8126 351 8164 385
rect 8198 351 8236 385
rect 8270 351 8308 385
rect 8342 351 8380 385
rect 8414 351 8452 385
rect 8486 351 8524 385
rect 8558 351 8596 385
rect 8630 351 8668 385
rect 8702 351 8740 385
rect 8774 351 8812 385
rect 8846 351 8884 385
rect 8918 351 8956 385
rect 8990 351 9028 385
rect 9062 351 9100 385
rect 9134 351 9172 385
rect 9206 351 9244 385
rect 9278 351 9284 385
rect 7870 312 9284 351
rect 7870 278 7876 312
rect 7910 278 7948 312
rect 7982 278 8020 312
rect 8054 278 8092 312
rect 8126 278 8164 312
rect 8198 278 8236 312
rect 8270 278 8308 312
rect 8342 278 8380 312
rect 8414 278 8452 312
rect 8486 278 8524 312
rect 8558 278 8596 312
rect 8630 278 8668 312
rect 8702 278 8740 312
rect 8774 278 8812 312
rect 8846 278 8884 312
rect 8918 278 8956 312
rect 8990 278 9028 312
rect 9062 278 9100 312
rect 9134 278 9172 312
rect 9206 278 9244 312
rect 9278 278 9284 312
rect 7870 239 9284 278
rect 7870 205 7876 239
rect 7910 205 7948 239
rect 7982 205 8020 239
rect 8054 205 8092 239
rect 8126 205 8164 239
rect 8198 205 8236 239
rect 8270 205 8308 239
rect 8342 205 8380 239
rect 8414 205 8452 239
rect 8486 205 8524 239
rect 8558 205 8596 239
rect 8630 205 8668 239
rect 8702 205 8740 239
rect 8774 205 8812 239
rect 8846 205 8884 239
rect 8918 205 8956 239
rect 8990 205 9028 239
rect 9062 205 9100 239
rect 9134 205 9172 239
rect 9206 205 9244 239
rect 9278 205 9284 239
rect 7870 166 9284 205
rect 7870 132 7876 166
rect 7910 132 7948 166
rect 7982 132 8020 166
rect 8054 132 8092 166
rect 8126 132 8164 166
rect 8198 132 8236 166
rect 8270 132 8308 166
rect 8342 132 8380 166
rect 8414 132 8452 166
rect 8486 132 8524 166
rect 8558 132 8596 166
rect 8630 132 8668 166
rect 8702 132 8740 166
rect 8774 132 8812 166
rect 8846 132 8884 166
rect 8918 132 8956 166
rect 8990 132 9028 166
rect 9062 132 9100 166
rect 9134 132 9172 166
rect 9206 132 9244 166
rect 9278 132 9284 166
rect 2656 58 2708 70
rect 2656 0 2708 6
rect 6278 122 6330 128
rect 6278 58 6330 70
rect 6278 0 6330 6
rect 7158 122 7210 128
rect 7158 58 7210 70
rect 7870 93 9284 132
rect 7870 59 7876 93
rect 7910 59 7948 93
rect 7982 59 8020 93
rect 8054 59 8092 93
rect 8126 59 8164 93
rect 8198 59 8236 93
rect 8270 59 8308 93
rect 8342 59 8380 93
rect 8414 59 8452 93
rect 8486 59 8524 93
rect 8558 59 8596 93
rect 8630 59 8668 93
rect 8702 59 8740 93
rect 8774 59 8812 93
rect 8846 59 8884 93
rect 8918 59 8956 93
rect 8990 59 9028 93
rect 9062 59 9100 93
rect 9134 59 9172 93
rect 9206 59 9244 93
rect 9278 59 9284 93
rect 7870 27 9284 59
rect 7158 0 7210 6
<< via1 >>
rect 3808 29351 3860 29403
rect 3872 29351 3924 29403
rect 5226 29351 5278 29403
rect 5290 29351 5342 29403
rect 315 9189 321 9241
rect 321 9189 367 9241
rect 379 9189 431 9241
rect 315 9123 321 9175
rect 321 9123 367 9175
rect 379 9123 431 9175
rect 315 9057 321 9109
rect 321 9057 367 9109
rect 379 9057 431 9109
rect 315 8991 321 9043
rect 321 8991 367 9043
rect 379 8991 431 9043
rect 315 8925 321 8977
rect 321 8925 367 8977
rect 379 8925 431 8977
rect 315 8859 321 8911
rect 321 8859 367 8911
rect 379 8859 431 8911
rect 315 8792 321 8844
rect 321 8792 367 8844
rect 379 8792 431 8844
rect 315 8725 321 8777
rect 321 8725 367 8777
rect 379 8725 431 8777
rect 315 8658 321 8710
rect 321 8658 367 8710
rect 379 8658 431 8710
rect 315 8591 321 8643
rect 321 8591 367 8643
rect 379 8591 431 8643
rect 315 8524 321 8576
rect 321 8524 367 8576
rect 379 8524 431 8576
rect 315 8457 321 8509
rect 321 8457 367 8509
rect 379 8457 431 8509
rect 315 8390 321 8442
rect 321 8390 367 8442
rect 379 8390 431 8442
rect 315 8323 321 8375
rect 321 8323 367 8375
rect 379 8323 431 8375
rect 418 4083 470 4135
rect 525 4083 577 4135
rect 632 4083 684 4135
rect 739 4083 791 4135
rect 845 4083 897 4135
rect 951 4083 1003 4135
rect 418 3993 470 4045
rect 525 3993 577 4045
rect 632 3993 684 4045
rect 739 3993 791 4045
rect 845 3993 897 4045
rect 951 3993 1003 4045
rect 3938 29267 3990 29319
rect 4002 29267 4054 29319
rect 5325 29267 5377 29319
rect 5389 29267 5441 29319
rect 4045 29183 4097 29235
rect 4109 29183 4161 29235
rect 5431 29183 5483 29235
rect 5495 29183 5547 29235
rect 4151 29099 4203 29151
rect 4215 29099 4267 29151
rect 5538 29099 5590 29151
rect 5602 29099 5654 29151
rect 1144 7520 1196 7572
rect 1144 7456 1196 7508
rect 4250 29015 4302 29067
rect 4314 29015 4366 29067
rect 5668 29015 5720 29067
rect 5732 29015 5784 29067
rect 1312 10636 1364 10688
rect 1312 10572 1364 10624
rect 1228 6698 1280 6750
rect 1228 6634 1280 6686
rect 1312 10197 1364 10249
rect 1312 10133 1364 10185
rect 4627 22731 4679 22783
rect 4627 22641 4679 22693
rect 4627 22551 4679 22603
rect 5004 18602 5056 18654
rect 5072 18602 5124 18654
rect 5140 18602 5192 18654
rect 5004 18536 5056 18588
rect 5072 18536 5124 18588
rect 5140 18536 5192 18588
rect 1648 15684 1700 15736
rect 1648 15620 1700 15672
rect 1564 14786 1616 14838
rect 1564 14722 1616 14774
rect 1648 15245 1700 15297
rect 1648 15181 1700 15233
rect 1480 9738 1532 9790
rect 1480 9674 1532 9726
rect 1396 3906 1448 3958
rect 1396 3842 1448 3894
rect 1312 70 1364 122
rect 1312 6 1364 58
rect 1732 11746 1784 11798
rect 1732 11682 1784 11734
rect 5004 16429 5056 16481
rect 5072 16472 5124 16481
rect 5072 16438 5080 16472
rect 5080 16438 5114 16472
rect 5114 16438 5124 16472
rect 5072 16429 5124 16438
rect 5140 16472 5192 16481
rect 5140 16438 5156 16472
rect 5156 16438 5190 16472
rect 5190 16438 5192 16472
rect 5140 16429 5192 16438
rect 7044 15820 7096 15872
rect 7160 15820 7212 15872
rect 7044 15753 7096 15805
rect 7160 15753 7212 15805
rect 7044 15685 7096 15737
rect 7160 15685 7212 15737
rect 1900 12568 1952 12620
rect 1900 12504 1952 12556
rect 4422 15514 4474 15566
rect 4490 15514 4542 15566
rect 4558 15514 4610 15566
rect 2089 15457 2141 15509
rect 2173 15457 2225 15509
rect 2257 15457 2309 15509
rect 2341 15457 2393 15509
rect 2425 15457 2477 15509
rect 2089 15367 2141 15419
rect 2173 15367 2225 15419
rect 2257 15367 2309 15419
rect 2341 15367 2393 15419
rect 2425 15367 2477 15419
rect 2882 15457 2934 15509
rect 2995 15457 3047 15509
rect 3107 15457 3159 15509
rect 4422 15430 4474 15482
rect 4490 15430 4542 15482
rect 4558 15430 4610 15482
rect 2882 15367 2934 15419
rect 2995 15367 3047 15419
rect 3107 15367 3159 15419
rect 1816 5588 1868 5640
rect 1816 5524 1868 5576
rect 1900 12187 1952 12239
rect 1900 12123 1952 12175
rect 1648 70 1700 122
rect 1648 6 1700 58
rect 3877 14626 3929 14678
rect 3951 14626 4003 14678
rect 4025 14626 4077 14678
rect 3877 14558 3929 14610
rect 3951 14558 4003 14610
rect 4025 14558 4077 14610
rect 3877 14490 3929 14542
rect 3951 14490 4003 14542
rect 4025 14490 4077 14542
rect 4422 14371 4474 14423
rect 4490 14371 4542 14423
rect 4558 14371 4610 14423
rect 4422 14287 4474 14339
rect 4490 14287 4542 14339
rect 4558 14287 4610 14339
rect 7044 14101 7096 14153
rect 7160 14101 7212 14153
rect 7044 14034 7096 14086
rect 7160 14034 7212 14086
rect 7044 13966 7096 14018
rect 7160 13966 7212 14018
rect 2944 13737 2996 13789
rect 2944 13669 2996 13721
rect 2944 13601 2996 13653
rect 4422 12990 4474 13042
rect 4490 12990 4542 13042
rect 4558 12990 4610 13042
rect 4422 12906 4474 12958
rect 4490 12906 4542 12958
rect 4558 12906 4610 12958
rect 3877 12800 3929 12852
rect 3951 12800 4003 12852
rect 4025 12800 4077 12852
rect 3877 12732 3929 12784
rect 3951 12732 4003 12784
rect 4025 12732 4077 12784
rect 3877 12664 3929 12716
rect 3951 12664 4003 12716
rect 4025 12664 4077 12716
rect 2089 11923 2141 11975
rect 2173 11923 2225 11975
rect 2257 11923 2309 11975
rect 2341 11923 2393 11975
rect 2425 11923 2477 11975
rect 2089 11833 2141 11885
rect 2173 11833 2225 11885
rect 2257 11833 2309 11885
rect 2341 11833 2393 11885
rect 2425 11833 2477 11885
rect 2882 11923 2934 11975
rect 2995 11923 3047 11975
rect 3107 11923 3159 11975
rect 2882 11833 2934 11885
rect 2995 11833 3047 11885
rect 3107 11833 3159 11885
rect 4422 11857 4474 11909
rect 4490 11857 4542 11909
rect 4558 11857 4610 11909
rect 4422 11773 4474 11825
rect 4490 11773 4542 11825
rect 4558 11773 4610 11825
rect 4433 11409 4485 11461
rect 4558 11409 4610 11461
rect 4433 11325 4485 11377
rect 4558 11325 4610 11377
rect 7044 13379 7096 13431
rect 7160 13379 7212 13431
rect 7044 13312 7096 13364
rect 7160 13312 7212 13364
rect 7044 13244 7096 13296
rect 7160 13244 7212 13296
rect 7044 11580 7096 11632
rect 7160 11580 7212 11632
rect 7044 11513 7096 11565
rect 7160 11513 7212 11565
rect 7044 11445 7096 11497
rect 7160 11445 7212 11497
rect 2089 10409 2141 10461
rect 2173 10409 2225 10461
rect 2257 10409 2309 10461
rect 2341 10409 2393 10461
rect 2425 10409 2477 10461
rect 2089 10319 2141 10371
rect 2173 10319 2225 10371
rect 2257 10319 2309 10371
rect 2341 10319 2393 10371
rect 2425 10319 2477 10371
rect 2882 10409 2934 10461
rect 2995 10409 3047 10461
rect 3107 10409 3159 10461
rect 2882 10319 2934 10371
rect 2995 10319 3047 10371
rect 3107 10319 3159 10371
rect 4422 10459 4474 10511
rect 4490 10459 4542 10511
rect 4558 10459 4610 10511
rect 4422 10375 4474 10427
rect 4490 10375 4542 10427
rect 4558 10375 4610 10427
rect 3877 9578 3929 9630
rect 3951 9578 4003 9630
rect 4025 9578 4077 9630
rect 3877 9510 3929 9562
rect 3951 9510 4003 9562
rect 4025 9510 4077 9562
rect 3877 9442 3929 9494
rect 3951 9442 4003 9494
rect 4025 9442 4077 9494
rect 2085 9189 2137 9241
rect 2171 9189 2223 9241
rect 2257 9189 2309 9241
rect 2343 9189 2395 9241
rect 2429 9189 2481 9241
rect 2085 9108 2137 9160
rect 2171 9108 2223 9160
rect 2257 9108 2309 9160
rect 2343 9108 2395 9160
rect 2429 9108 2481 9160
rect 2085 9027 2137 9079
rect 2171 9027 2223 9079
rect 2257 9027 2309 9079
rect 2343 9027 2395 9079
rect 2429 9027 2481 9079
rect 2085 8945 2137 8997
rect 2171 8945 2223 8997
rect 2257 8945 2309 8997
rect 2343 8945 2395 8997
rect 2429 8945 2481 8997
rect 2085 8863 2137 8915
rect 2171 8863 2223 8915
rect 2257 8863 2309 8915
rect 2343 8863 2395 8915
rect 2429 8863 2481 8915
rect 2085 8781 2137 8833
rect 2171 8781 2223 8833
rect 2257 8781 2309 8833
rect 2343 8781 2395 8833
rect 2429 8781 2481 8833
rect 4422 9337 4474 9389
rect 4490 9337 4542 9389
rect 4558 9337 4610 9389
rect 4422 9253 4474 9305
rect 4490 9253 4542 9305
rect 4558 9253 4610 9305
rect 2944 8658 2996 8710
rect 2944 8590 2996 8642
rect 2944 8522 2996 8574
rect 7044 10892 7096 10944
rect 7160 10892 7212 10944
rect 7044 10825 7096 10877
rect 7160 10825 7212 10877
rect 7044 10757 7096 10809
rect 7160 10757 7212 10809
rect 7044 9146 7096 9198
rect 7160 9146 7212 9198
rect 7044 9079 7096 9131
rect 7160 9079 7212 9131
rect 7044 9011 7096 9063
rect 7160 9011 7212 9063
rect 4422 7950 4474 8002
rect 4490 7950 4542 8002
rect 4558 7950 4610 8002
rect 4422 7866 4474 7918
rect 4490 7866 4542 7918
rect 4558 7866 4610 7918
rect 3877 7752 3929 7804
rect 3951 7752 4003 7804
rect 4025 7752 4077 7804
rect 3877 7684 3929 7736
rect 3951 7684 4003 7736
rect 4025 7684 4077 7736
rect 3877 7616 3929 7668
rect 3951 7616 4003 7668
rect 4025 7616 4077 7668
rect 2089 6875 2141 6927
rect 2173 6875 2225 6927
rect 2257 6875 2309 6927
rect 2341 6875 2393 6927
rect 2425 6875 2477 6927
rect 2089 6785 2141 6837
rect 2173 6785 2225 6837
rect 2257 6785 2309 6837
rect 2341 6785 2393 6837
rect 2425 6785 2477 6837
rect 2089 5361 2141 5413
rect 2173 5361 2225 5413
rect 2257 5361 2309 5413
rect 2341 5361 2393 5413
rect 2425 5361 2477 5413
rect 2089 5271 2141 5323
rect 2173 5271 2225 5323
rect 2257 5271 2309 5323
rect 2341 5271 2393 5323
rect 2425 5271 2477 5323
rect 2656 7139 2708 7191
rect 2656 7075 2708 7127
rect 1900 70 1952 122
rect 1900 6 1952 58
rect 2152 5149 2204 5201
rect 2152 5085 2204 5137
rect 2152 70 2204 122
rect 2152 6 2204 58
rect 2404 4347 2456 4399
rect 2404 4283 2456 4335
rect 2404 70 2456 122
rect 2404 6 2456 58
rect 2882 6875 2934 6927
rect 2995 6875 3047 6927
rect 3107 6875 3159 6927
rect 2882 6785 2934 6837
rect 2995 6785 3047 6837
rect 3107 6785 3159 6837
rect 4422 6828 4474 6880
rect 4490 6828 4542 6880
rect 4558 6828 4610 6880
rect 4422 6744 4474 6796
rect 4490 6744 4542 6796
rect 4558 6744 4610 6796
rect 7044 8377 7096 8429
rect 7160 8377 7212 8429
rect 7044 8310 7096 8362
rect 7160 8310 7212 8362
rect 7044 8242 7096 8294
rect 7160 8242 7212 8294
rect 7044 6645 7096 6697
rect 7160 6645 7212 6697
rect 7044 6578 7096 6630
rect 7160 6578 7212 6630
rect 7044 6510 7096 6562
rect 7160 6510 7212 6562
rect 4422 5434 4474 5486
rect 4490 5434 4542 5486
rect 4558 5434 4610 5486
rect 2882 5361 2934 5413
rect 2995 5361 3047 5413
rect 3107 5361 3159 5413
rect 2882 5271 2934 5323
rect 2995 5271 3047 5323
rect 3107 5271 3159 5323
rect 4422 5350 4474 5402
rect 4490 5350 4542 5402
rect 4558 5350 4610 5402
rect 2882 4083 2934 4135
rect 2995 4083 3047 4135
rect 3107 4083 3159 4135
rect 2882 3993 2934 4045
rect 2995 3993 3047 4045
rect 3107 3993 3159 4045
rect 7044 5858 7096 5910
rect 7160 5858 7212 5910
rect 7044 5791 7096 5843
rect 7160 5791 7212 5843
rect 7044 5723 7096 5775
rect 7160 5723 7212 5775
rect 7044 4809 7096 4861
rect 7160 4809 7212 4861
rect 7044 4742 7096 4794
rect 7160 4742 7212 4794
rect 7044 4674 7096 4726
rect 7160 4674 7212 4726
rect 4422 4006 4474 4058
rect 4490 4006 4542 4058
rect 4558 4006 4610 4058
rect 4422 3922 4474 3974
rect 4490 3922 4542 3974
rect 4558 3922 4610 3974
rect 2944 3259 2996 3311
rect 2944 3191 2996 3243
rect 2944 3123 2996 3175
rect 3877 3259 3929 3311
rect 3951 3259 4003 3311
rect 4025 3259 4077 3311
rect 3877 3191 3929 3243
rect 3951 3191 4003 3243
rect 4025 3191 4077 3243
rect 3877 3123 3929 3175
rect 3951 3123 4003 3175
rect 4025 3123 4077 3175
rect 7044 3673 7096 3725
rect 7160 3673 7212 3725
rect 7044 3606 7096 3658
rect 7160 3606 7212 3658
rect 7044 3538 7096 3590
rect 7160 3538 7212 3590
rect 4416 3264 4468 3316
rect 4490 3264 4542 3316
rect 4564 3264 4616 3316
rect 4416 3136 4468 3188
rect 4490 3136 4542 3188
rect 4564 3136 4616 3188
rect 4416 3008 4468 3060
rect 4490 3008 4542 3060
rect 4564 3008 4616 3060
rect 4416 2880 4468 2932
rect 4490 2880 4542 2932
rect 4564 2880 4616 2932
rect 4736 3229 4788 3281
rect 4736 3165 4788 3217
rect 4656 2992 4708 3044
rect 4656 2928 4708 2980
rect 7044 3163 7096 3215
rect 7160 3163 7212 3215
rect 7044 3096 7096 3148
rect 7160 3096 7212 3148
rect 7044 3028 7096 3080
rect 7160 3028 7212 3080
rect 4416 2752 4468 2804
rect 4490 2752 4542 2804
rect 4564 2752 4616 2804
rect 4416 2624 4468 2676
rect 4490 2624 4542 2676
rect 4564 2624 4616 2676
rect 4416 2495 4468 2547
rect 4490 2495 4542 2547
rect 4564 2495 4616 2547
rect 4416 2366 4468 2418
rect 4490 2366 4542 2418
rect 4564 2366 4616 2418
rect 6079 2936 6131 2988
rect 6079 2872 6131 2924
rect 5989 2775 6041 2827
rect 5989 2711 6041 2763
rect 6278 2773 6330 2825
rect 6278 2709 6330 2761
rect 7158 2773 7210 2825
rect 7158 2709 7210 2761
rect 6278 2311 6330 2363
rect 6278 2247 6330 2299
rect 3477 2136 3529 2188
rect 3586 2136 3638 2188
rect 3695 2136 3747 2188
rect 3803 2136 3855 2188
rect 3911 2136 3963 2188
rect 4019 2136 4071 2188
rect 3477 2054 3529 2106
rect 3586 2054 3638 2106
rect 3695 2054 3747 2106
rect 3803 2054 3855 2106
rect 3911 2054 3963 2106
rect 4019 2054 4071 2106
rect 3477 1972 3529 2024
rect 3586 1972 3638 2024
rect 3695 1972 3747 2024
rect 3803 1972 3855 2024
rect 3911 1972 3963 2024
rect 4019 1972 4071 2024
rect 3477 1890 3529 1942
rect 3586 1890 3638 1942
rect 3695 1890 3747 1942
rect 3803 1890 3855 1942
rect 3911 1890 3963 1942
rect 4019 1890 4071 1942
rect 8534 9189 8586 9241
rect 8598 9189 8650 9241
rect 8662 9189 8714 9241
rect 8726 9189 8778 9241
rect 8790 9189 8842 9241
rect 8854 9189 8906 9241
rect 8918 9189 8970 9241
rect 8982 9189 9034 9241
rect 9046 9189 9098 9241
rect 9110 9189 9162 9241
rect 9174 9189 9226 9241
rect 8534 9123 8586 9175
rect 8598 9123 8650 9175
rect 8662 9123 8714 9175
rect 8726 9123 8778 9175
rect 8790 9123 8842 9175
rect 8854 9123 8906 9175
rect 8918 9123 8970 9175
rect 8982 9123 9034 9175
rect 9046 9123 9098 9175
rect 9110 9123 9162 9175
rect 9174 9123 9226 9175
rect 8534 9057 8586 9109
rect 8598 9057 8650 9109
rect 8662 9057 8714 9109
rect 8726 9057 8778 9109
rect 8790 9057 8842 9109
rect 8854 9057 8906 9109
rect 8918 9057 8970 9109
rect 8982 9057 9034 9109
rect 9046 9057 9098 9109
rect 9110 9057 9162 9109
rect 9174 9057 9226 9109
rect 8534 8991 8586 9043
rect 8598 8991 8650 9043
rect 8662 8991 8714 9043
rect 8726 8991 8778 9043
rect 8790 8991 8842 9043
rect 8854 8991 8906 9043
rect 8918 8991 8970 9043
rect 8982 8991 9034 9043
rect 9046 8991 9098 9043
rect 9110 8991 9162 9043
rect 9174 8991 9226 9043
rect 8534 8925 8586 8977
rect 8598 8925 8650 8977
rect 8662 8925 8714 8977
rect 8726 8925 8778 8977
rect 8790 8925 8842 8977
rect 8854 8925 8906 8977
rect 8918 8925 8970 8977
rect 8982 8925 9034 8977
rect 9046 8925 9098 8977
rect 9110 8925 9162 8977
rect 9174 8925 9226 8977
rect 8534 8859 8586 8911
rect 8598 8859 8650 8911
rect 8662 8859 8714 8911
rect 8726 8859 8778 8911
rect 8790 8859 8842 8911
rect 8854 8859 8906 8911
rect 8918 8859 8970 8911
rect 8982 8859 9034 8911
rect 9046 8859 9098 8911
rect 9110 8859 9162 8911
rect 9174 8859 9226 8911
rect 8534 8792 8586 8844
rect 8598 8792 8650 8844
rect 8662 8792 8714 8844
rect 8726 8792 8778 8844
rect 8790 8792 8842 8844
rect 8854 8792 8906 8844
rect 8918 8792 8970 8844
rect 8982 8792 9034 8844
rect 9046 8792 9098 8844
rect 9110 8792 9162 8844
rect 9174 8792 9226 8844
rect 8534 8725 8586 8777
rect 8598 8725 8650 8777
rect 8662 8725 8714 8777
rect 8726 8725 8778 8777
rect 8790 8725 8842 8777
rect 8854 8725 8906 8777
rect 8918 8725 8970 8777
rect 8982 8725 9034 8777
rect 9046 8725 9098 8777
rect 9110 8725 9162 8777
rect 9174 8725 9226 8777
rect 8534 8658 8586 8710
rect 8598 8658 8650 8710
rect 8662 8658 8714 8710
rect 8726 8658 8778 8710
rect 8790 8658 8842 8710
rect 8854 8658 8906 8710
rect 8918 8658 8970 8710
rect 8982 8658 9034 8710
rect 9046 8658 9098 8710
rect 9110 8658 9162 8710
rect 9174 8658 9226 8710
rect 8534 8591 8586 8643
rect 8598 8591 8650 8643
rect 8662 8591 8714 8643
rect 8726 8591 8778 8643
rect 8790 8591 8842 8643
rect 8854 8591 8906 8643
rect 8918 8591 8970 8643
rect 8982 8591 9034 8643
rect 9046 8591 9098 8643
rect 9110 8591 9162 8643
rect 9174 8591 9226 8643
rect 8534 8524 8586 8576
rect 8598 8524 8650 8576
rect 8662 8524 8714 8576
rect 8726 8524 8778 8576
rect 8790 8524 8842 8576
rect 8854 8524 8906 8576
rect 8918 8524 8970 8576
rect 8982 8524 9034 8576
rect 9046 8524 9098 8576
rect 9110 8524 9162 8576
rect 9174 8524 9226 8576
rect 8534 8457 8586 8509
rect 8598 8457 8650 8509
rect 8662 8457 8714 8509
rect 8726 8457 8778 8509
rect 8790 8457 8842 8509
rect 8854 8457 8906 8509
rect 8918 8457 8970 8509
rect 8982 8457 9034 8509
rect 9046 8457 9098 8509
rect 9110 8457 9162 8509
rect 9174 8457 9226 8509
rect 8534 8390 8586 8442
rect 8598 8390 8650 8442
rect 8662 8390 8714 8442
rect 8726 8390 8778 8442
rect 8790 8390 8842 8442
rect 8854 8390 8906 8442
rect 8918 8390 8970 8442
rect 8982 8390 9034 8442
rect 9046 8390 9098 8442
rect 9110 8390 9162 8442
rect 9174 8390 9226 8442
rect 8534 8323 8586 8375
rect 8598 8323 8650 8375
rect 8662 8323 8714 8375
rect 8726 8323 8778 8375
rect 8790 8323 8842 8375
rect 8854 8323 8906 8375
rect 8918 8323 8970 8375
rect 8982 8323 9034 8375
rect 9046 8323 9098 8375
rect 9110 8323 9162 8375
rect 9174 8323 9226 8375
rect 2656 70 2708 122
rect 2656 6 2708 58
rect 6278 70 6330 122
rect 6278 6 6330 58
rect 7158 70 7210 122
rect 7158 6 7210 58
<< metal2 >>
rect 1949 39865 2593 39874
rect 2005 39809 2033 39865
rect 2089 39809 2117 39865
rect 2173 39809 2201 39865
rect 2257 39809 2285 39865
rect 2341 39809 2369 39865
rect 2425 39809 2453 39865
rect 2509 39809 2537 39865
rect 1949 39785 2593 39809
rect 2005 39729 2033 39785
rect 2089 39729 2117 39785
rect 2173 39729 2201 39785
rect 2257 39729 2285 39785
rect 2341 39729 2369 39785
rect 2425 39729 2453 39785
rect 2509 39729 2537 39785
rect 1949 39705 2593 39729
rect 2005 39649 2033 39705
rect 2089 39649 2117 39705
rect 2173 39649 2201 39705
rect 2257 39649 2285 39705
rect 2341 39649 2369 39705
rect 2425 39649 2453 39705
rect 2509 39649 2537 39705
rect 1949 39625 2593 39649
rect 2005 39569 2033 39625
rect 2089 39569 2117 39625
rect 2173 39569 2201 39625
rect 2257 39569 2285 39625
rect 2341 39569 2369 39625
rect 2425 39569 2453 39625
rect 2509 39569 2537 39625
rect 1949 39545 2593 39569
rect 2005 39489 2033 39545
rect 2089 39489 2117 39545
rect 2173 39489 2201 39545
rect 2257 39489 2285 39545
rect 2341 39489 2369 39545
rect 2425 39489 2453 39545
rect 2509 39489 2537 39545
rect 1949 39465 2593 39489
rect 2005 39409 2033 39465
rect 2089 39409 2117 39465
rect 2173 39409 2201 39465
rect 2257 39409 2285 39465
rect 2341 39409 2369 39465
rect 2425 39409 2453 39465
rect 2509 39409 2537 39465
rect 1949 39385 2593 39409
rect 2005 39329 2033 39385
rect 2089 39329 2117 39385
rect 2173 39329 2201 39385
rect 2257 39329 2285 39385
rect 2341 39329 2369 39385
rect 2425 39329 2453 39385
rect 2509 39329 2537 39385
rect 1949 39305 2593 39329
rect 2005 39249 2033 39305
rect 2089 39249 2117 39305
rect 2173 39249 2201 39305
rect 2257 39249 2285 39305
rect 2341 39249 2369 39305
rect 2425 39249 2453 39305
rect 2509 39249 2537 39305
rect 1949 39225 2593 39249
rect 2005 39169 2033 39225
rect 2089 39169 2117 39225
rect 2173 39169 2201 39225
rect 2257 39169 2285 39225
rect 2341 39169 2369 39225
rect 2425 39169 2453 39225
rect 2509 39169 2537 39225
rect 1949 39145 2593 39169
rect 2005 39089 2033 39145
rect 2089 39089 2117 39145
rect 2173 39089 2201 39145
rect 2257 39089 2285 39145
rect 2341 39089 2369 39145
rect 2425 39089 2453 39145
rect 2509 39089 2537 39145
rect 1949 39065 2593 39089
rect 2005 39009 2033 39065
rect 2089 39009 2117 39065
rect 2173 39009 2201 39065
rect 2257 39009 2285 39065
rect 2341 39009 2369 39065
rect 2425 39009 2453 39065
rect 2509 39009 2537 39065
rect 1949 38985 2593 39009
rect 2005 38929 2033 38985
rect 2089 38929 2117 38985
rect 2173 38929 2201 38985
rect 2257 38929 2285 38985
rect 2341 38929 2369 38985
rect 2425 38929 2453 38985
rect 2509 38929 2537 38985
rect 1949 38905 2593 38929
rect 2005 38849 2033 38905
rect 2089 38849 2117 38905
rect 2173 38849 2201 38905
rect 2257 38849 2285 38905
rect 2341 38849 2369 38905
rect 2425 38849 2453 38905
rect 2509 38849 2537 38905
rect 1949 38825 2593 38849
rect 2005 38769 2033 38825
rect 2089 38769 2117 38825
rect 2173 38769 2201 38825
rect 2257 38769 2285 38825
rect 2341 38769 2369 38825
rect 2425 38769 2453 38825
rect 2509 38769 2537 38825
rect 1949 38745 2593 38769
rect 2005 38689 2033 38745
rect 2089 38689 2117 38745
rect 2173 38689 2201 38745
rect 2257 38689 2285 38745
rect 2341 38689 2369 38745
rect 2425 38689 2453 38745
rect 2509 38689 2537 38745
rect 1949 38665 2593 38689
rect 2005 38609 2033 38665
rect 2089 38609 2117 38665
rect 2173 38609 2201 38665
rect 2257 38609 2285 38665
rect 2341 38609 2369 38665
rect 2425 38609 2453 38665
rect 2509 38609 2537 38665
rect 1949 38585 2593 38609
rect 2005 38529 2033 38585
rect 2089 38529 2117 38585
rect 2173 38529 2201 38585
rect 2257 38529 2285 38585
rect 2341 38529 2369 38585
rect 2425 38529 2453 38585
rect 2509 38529 2537 38585
rect 1949 38505 2593 38529
rect 2005 38449 2033 38505
rect 2089 38449 2117 38505
rect 2173 38449 2201 38505
rect 2257 38449 2285 38505
rect 2341 38449 2369 38505
rect 2425 38449 2453 38505
rect 2509 38449 2537 38505
rect 1949 38425 2593 38449
rect 2005 38369 2033 38425
rect 2089 38369 2117 38425
rect 2173 38369 2201 38425
rect 2257 38369 2285 38425
rect 2341 38369 2369 38425
rect 2425 38369 2453 38425
rect 2509 38369 2537 38425
rect 1949 38345 2593 38369
rect 2005 38289 2033 38345
rect 2089 38289 2117 38345
rect 2173 38289 2201 38345
rect 2257 38289 2285 38345
rect 2341 38289 2369 38345
rect 2425 38289 2453 38345
rect 2509 38289 2537 38345
rect 1949 38265 2593 38289
rect 2005 38209 2033 38265
rect 2089 38209 2117 38265
rect 2173 38209 2201 38265
rect 2257 38209 2285 38265
rect 2341 38209 2369 38265
rect 2425 38209 2453 38265
rect 2509 38209 2537 38265
rect 1949 38185 2593 38209
rect 2005 38129 2033 38185
rect 2089 38129 2117 38185
rect 2173 38129 2201 38185
rect 2257 38129 2285 38185
rect 2341 38129 2369 38185
rect 2425 38129 2453 38185
rect 2509 38129 2537 38185
rect 1949 38105 2593 38129
rect 2005 38049 2033 38105
rect 2089 38049 2117 38105
rect 2173 38049 2201 38105
rect 2257 38049 2285 38105
rect 2341 38049 2369 38105
rect 2425 38049 2453 38105
rect 2509 38049 2537 38105
rect 1949 38025 2593 38049
rect 2005 37969 2033 38025
rect 2089 37969 2117 38025
rect 2173 37969 2201 38025
rect 2257 37969 2285 38025
rect 2341 37969 2369 38025
rect 2425 37969 2453 38025
rect 2509 37969 2537 38025
rect 1949 37945 2593 37969
rect 2005 37889 2033 37945
rect 2089 37889 2117 37945
rect 2173 37889 2201 37945
rect 2257 37889 2285 37945
rect 2341 37889 2369 37945
rect 2425 37889 2453 37945
rect 2509 37889 2537 37945
rect 1949 37865 2593 37889
rect 2005 37809 2033 37865
rect 2089 37809 2117 37865
rect 2173 37809 2201 37865
rect 2257 37809 2285 37865
rect 2341 37809 2369 37865
rect 2425 37809 2453 37865
rect 2509 37809 2537 37865
rect 1949 37785 2593 37809
rect 2005 37729 2033 37785
rect 2089 37729 2117 37785
rect 2173 37729 2201 37785
rect 2257 37729 2285 37785
rect 2341 37729 2369 37785
rect 2425 37729 2453 37785
rect 2509 37729 2537 37785
rect 1949 37705 2593 37729
rect 2005 37649 2033 37705
rect 2089 37649 2117 37705
rect 2173 37649 2201 37705
rect 2257 37649 2285 37705
rect 2341 37649 2369 37705
rect 2425 37649 2453 37705
rect 2509 37649 2537 37705
rect 1949 37625 2593 37649
rect 2005 37569 2033 37625
rect 2089 37569 2117 37625
rect 2173 37569 2201 37625
rect 2257 37569 2285 37625
rect 2341 37569 2369 37625
rect 2425 37569 2453 37625
rect 2509 37569 2537 37625
rect 1949 37545 2593 37569
rect 2005 37489 2033 37545
rect 2089 37489 2117 37545
rect 2173 37489 2201 37545
rect 2257 37489 2285 37545
rect 2341 37489 2369 37545
rect 2425 37489 2453 37545
rect 2509 37489 2537 37545
rect 1949 37465 2593 37489
rect 2005 37409 2033 37465
rect 2089 37409 2117 37465
rect 2173 37409 2201 37465
rect 2257 37409 2285 37465
rect 2341 37409 2369 37465
rect 2425 37409 2453 37465
rect 2509 37409 2537 37465
rect 1949 37385 2593 37409
rect 2005 37329 2033 37385
rect 2089 37329 2117 37385
rect 2173 37329 2201 37385
rect 2257 37329 2285 37385
rect 2341 37329 2369 37385
rect 2425 37329 2453 37385
rect 2509 37329 2537 37385
rect 1949 37305 2593 37329
rect 2005 37249 2033 37305
rect 2089 37249 2117 37305
rect 2173 37249 2201 37305
rect 2257 37249 2285 37305
rect 2341 37249 2369 37305
rect 2425 37249 2453 37305
rect 2509 37249 2537 37305
rect 1949 37225 2593 37249
rect 2005 37169 2033 37225
rect 2089 37169 2117 37225
rect 2173 37169 2201 37225
rect 2257 37169 2285 37225
rect 2341 37169 2369 37225
rect 2425 37169 2453 37225
rect 2509 37169 2537 37225
rect 1949 37145 2593 37169
rect 2005 37089 2033 37145
rect 2089 37089 2117 37145
rect 2173 37089 2201 37145
rect 2257 37089 2285 37145
rect 2341 37089 2369 37145
rect 2425 37089 2453 37145
rect 2509 37089 2537 37145
rect 6900 39870 7502 39879
rect 6900 39814 6903 39870
rect 6959 39814 6993 39870
rect 7049 39814 7083 39870
rect 7139 39814 7173 39870
rect 7229 39814 7263 39870
rect 7319 39814 7353 39870
rect 7409 39814 7443 39870
rect 7499 39814 7502 39870
rect 6900 39790 7502 39814
rect 6900 39734 6903 39790
rect 6959 39734 6993 39790
rect 7049 39734 7083 39790
rect 7139 39734 7173 39790
rect 7229 39734 7263 39790
rect 7319 39734 7353 39790
rect 7409 39734 7443 39790
rect 7499 39734 7502 39790
rect 6900 39710 7502 39734
rect 6900 39654 6903 39710
rect 6959 39654 6993 39710
rect 7049 39654 7083 39710
rect 7139 39654 7173 39710
rect 7229 39654 7263 39710
rect 7319 39654 7353 39710
rect 7409 39654 7443 39710
rect 7499 39654 7502 39710
rect 6900 39630 7502 39654
rect 6900 39574 6903 39630
rect 6959 39574 6993 39630
rect 7049 39574 7083 39630
rect 7139 39574 7173 39630
rect 7229 39574 7263 39630
rect 7319 39574 7353 39630
rect 7409 39574 7443 39630
rect 7499 39574 7502 39630
rect 6900 39550 7502 39574
rect 6900 39494 6903 39550
rect 6959 39494 6993 39550
rect 7049 39494 7083 39550
rect 7139 39494 7173 39550
rect 7229 39494 7263 39550
rect 7319 39494 7353 39550
rect 7409 39494 7443 39550
rect 7499 39494 7502 39550
rect 6900 39470 7502 39494
rect 6900 39414 6903 39470
rect 6959 39414 6993 39470
rect 7049 39414 7083 39470
rect 7139 39414 7173 39470
rect 7229 39414 7263 39470
rect 7319 39414 7353 39470
rect 7409 39414 7443 39470
rect 7499 39414 7502 39470
rect 6900 39390 7502 39414
rect 6900 39334 6903 39390
rect 6959 39334 6993 39390
rect 7049 39334 7083 39390
rect 7139 39334 7173 39390
rect 7229 39334 7263 39390
rect 7319 39334 7353 39390
rect 7409 39334 7443 39390
rect 7499 39334 7502 39390
rect 6900 39310 7502 39334
rect 6900 39254 6903 39310
rect 6959 39254 6993 39310
rect 7049 39254 7083 39310
rect 7139 39254 7173 39310
rect 7229 39254 7263 39310
rect 7319 39254 7353 39310
rect 7409 39254 7443 39310
rect 7499 39254 7502 39310
rect 6900 39230 7502 39254
rect 6900 39174 6903 39230
rect 6959 39174 6993 39230
rect 7049 39174 7083 39230
rect 7139 39174 7173 39230
rect 7229 39174 7263 39230
rect 7319 39174 7353 39230
rect 7409 39174 7443 39230
rect 7499 39174 7502 39230
rect 6900 39150 7502 39174
rect 6900 39094 6903 39150
rect 6959 39094 6993 39150
rect 7049 39094 7083 39150
rect 7139 39094 7173 39150
rect 7229 39094 7263 39150
rect 7319 39094 7353 39150
rect 7409 39094 7443 39150
rect 7499 39094 7502 39150
rect 6900 39070 7502 39094
rect 6900 39014 6903 39070
rect 6959 39014 6993 39070
rect 7049 39014 7083 39070
rect 7139 39014 7173 39070
rect 7229 39014 7263 39070
rect 7319 39014 7353 39070
rect 7409 39014 7443 39070
rect 7499 39014 7502 39070
rect 6900 38990 7502 39014
rect 6900 38934 6903 38990
rect 6959 38934 6993 38990
rect 7049 38934 7083 38990
rect 7139 38934 7173 38990
rect 7229 38934 7263 38990
rect 7319 38934 7353 38990
rect 7409 38934 7443 38990
rect 7499 38934 7502 38990
rect 6900 38910 7502 38934
rect 6900 38854 6903 38910
rect 6959 38854 6993 38910
rect 7049 38854 7083 38910
rect 7139 38854 7173 38910
rect 7229 38854 7263 38910
rect 7319 38854 7353 38910
rect 7409 38854 7443 38910
rect 7499 38854 7502 38910
rect 6900 38830 7502 38854
rect 6900 38774 6903 38830
rect 6959 38774 6993 38830
rect 7049 38774 7083 38830
rect 7139 38774 7173 38830
rect 7229 38774 7263 38830
rect 7319 38774 7353 38830
rect 7409 38774 7443 38830
rect 7499 38774 7502 38830
rect 6900 38750 7502 38774
rect 6900 38694 6903 38750
rect 6959 38694 6993 38750
rect 7049 38694 7083 38750
rect 7139 38694 7173 38750
rect 7229 38694 7263 38750
rect 7319 38694 7353 38750
rect 7409 38694 7443 38750
rect 7499 38694 7502 38750
rect 6900 38670 7502 38694
rect 6900 38614 6903 38670
rect 6959 38614 6993 38670
rect 7049 38614 7083 38670
rect 7139 38614 7173 38670
rect 7229 38614 7263 38670
rect 7319 38614 7353 38670
rect 7409 38614 7443 38670
rect 7499 38614 7502 38670
rect 6900 38590 7502 38614
rect 6900 38534 6903 38590
rect 6959 38534 6993 38590
rect 7049 38534 7083 38590
rect 7139 38534 7173 38590
rect 7229 38534 7263 38590
rect 7319 38534 7353 38590
rect 7409 38534 7443 38590
rect 7499 38534 7502 38590
rect 6900 38510 7502 38534
rect 6900 38454 6903 38510
rect 6959 38454 6993 38510
rect 7049 38454 7083 38510
rect 7139 38454 7173 38510
rect 7229 38454 7263 38510
rect 7319 38454 7353 38510
rect 7409 38454 7443 38510
rect 7499 38454 7502 38510
rect 6900 38430 7502 38454
rect 6900 38374 6903 38430
rect 6959 38374 6993 38430
rect 7049 38374 7083 38430
rect 7139 38374 7173 38430
rect 7229 38374 7263 38430
rect 7319 38374 7353 38430
rect 7409 38374 7443 38430
rect 7499 38374 7502 38430
rect 6900 38350 7502 38374
rect 6900 38294 6903 38350
rect 6959 38294 6993 38350
rect 7049 38294 7083 38350
rect 7139 38294 7173 38350
rect 7229 38294 7263 38350
rect 7319 38294 7353 38350
rect 7409 38294 7443 38350
rect 7499 38294 7502 38350
rect 6900 38270 7502 38294
rect 6900 38214 6903 38270
rect 6959 38214 6993 38270
rect 7049 38214 7083 38270
rect 7139 38214 7173 38270
rect 7229 38214 7263 38270
rect 7319 38214 7353 38270
rect 7409 38214 7443 38270
rect 7499 38214 7502 38270
rect 6900 38190 7502 38214
rect 6900 38134 6903 38190
rect 6959 38134 6993 38190
rect 7049 38134 7083 38190
rect 7139 38134 7173 38190
rect 7229 38134 7263 38190
rect 7319 38134 7353 38190
rect 7409 38134 7443 38190
rect 7499 38134 7502 38190
rect 6900 38110 7502 38134
rect 6900 38054 6903 38110
rect 6959 38054 6993 38110
rect 7049 38054 7083 38110
rect 7139 38054 7173 38110
rect 7229 38054 7263 38110
rect 7319 38054 7353 38110
rect 7409 38054 7443 38110
rect 7499 38054 7502 38110
rect 6900 38030 7502 38054
rect 6900 37974 6903 38030
rect 6959 37974 6993 38030
rect 7049 37974 7083 38030
rect 7139 37974 7173 38030
rect 7229 37974 7263 38030
rect 7319 37974 7353 38030
rect 7409 37974 7443 38030
rect 7499 37974 7502 38030
rect 6900 37950 7502 37974
rect 6900 37894 6903 37950
rect 6959 37894 6993 37950
rect 7049 37894 7083 37950
rect 7139 37894 7173 37950
rect 7229 37894 7263 37950
rect 7319 37894 7353 37950
rect 7409 37894 7443 37950
rect 7499 37894 7502 37950
rect 6900 37870 7502 37894
rect 6900 37814 6903 37870
rect 6959 37814 6993 37870
rect 7049 37814 7083 37870
rect 7139 37814 7173 37870
rect 7229 37814 7263 37870
rect 7319 37814 7353 37870
rect 7409 37814 7443 37870
rect 7499 37814 7502 37870
rect 6900 37790 7502 37814
rect 6900 37734 6903 37790
rect 6959 37734 6993 37790
rect 7049 37734 7083 37790
rect 7139 37734 7173 37790
rect 7229 37734 7263 37790
rect 7319 37734 7353 37790
rect 7409 37734 7443 37790
rect 7499 37734 7502 37790
rect 6900 37710 7502 37734
rect 6900 37654 6903 37710
rect 6959 37654 6993 37710
rect 7049 37654 7083 37710
rect 7139 37654 7173 37710
rect 7229 37654 7263 37710
rect 7319 37654 7353 37710
rect 7409 37654 7443 37710
rect 7499 37654 7502 37710
rect 6900 37630 7502 37654
rect 6900 37574 6903 37630
rect 6959 37574 6993 37630
rect 7049 37574 7083 37630
rect 7139 37574 7173 37630
rect 7229 37574 7263 37630
rect 7319 37574 7353 37630
rect 7409 37574 7443 37630
rect 7499 37574 7502 37630
rect 6900 37550 7502 37574
rect 6900 37494 6903 37550
rect 6959 37494 6993 37550
rect 7049 37494 7083 37550
rect 7139 37494 7173 37550
rect 7229 37494 7263 37550
rect 7319 37494 7353 37550
rect 7409 37494 7443 37550
rect 7499 37494 7502 37550
rect 6900 37470 7502 37494
rect 6900 37414 6903 37470
rect 6959 37414 6993 37470
rect 7049 37414 7083 37470
rect 7139 37414 7173 37470
rect 7229 37414 7263 37470
rect 7319 37414 7353 37470
rect 7409 37414 7443 37470
rect 7499 37414 7502 37470
rect 6900 37390 7502 37414
rect 6900 37334 6903 37390
rect 6959 37334 6993 37390
rect 7049 37334 7083 37390
rect 7139 37334 7173 37390
rect 7229 37334 7263 37390
rect 7319 37334 7353 37390
rect 7409 37334 7443 37390
rect 7499 37334 7502 37390
rect 6900 37310 7502 37334
rect 6900 37254 6903 37310
rect 6959 37254 6993 37310
rect 7049 37254 7083 37310
rect 7139 37254 7173 37310
rect 7229 37254 7263 37310
rect 7319 37254 7353 37310
rect 7409 37254 7443 37310
rect 7499 37254 7502 37310
rect 6900 37230 7502 37254
rect 6900 37174 6903 37230
rect 6959 37174 6993 37230
rect 7049 37174 7083 37230
rect 7139 37174 7173 37230
rect 7229 37174 7263 37230
rect 7319 37174 7353 37230
rect 7409 37174 7443 37230
rect 7499 37174 7502 37230
rect 6900 37150 7502 37174
rect 1949 37065 2593 37089
rect 2005 37009 2033 37065
rect 2089 37009 2117 37065
rect 2173 37009 2201 37065
rect 2257 37009 2285 37065
rect 2341 37009 2369 37065
rect 2425 37009 2453 37065
rect 2509 37009 2537 37065
rect 1949 36985 2593 37009
rect 2005 36929 2033 36985
rect 2089 36929 2117 36985
rect 2173 36929 2201 36985
rect 2257 36929 2285 36985
rect 2341 36929 2369 36985
rect 2425 36929 2453 36985
rect 2509 36929 2537 36985
rect 1949 36905 2593 36929
rect 2005 36849 2033 36905
rect 2089 36849 2117 36905
rect 2173 36849 2201 36905
rect 2257 36849 2285 36905
rect 2341 36849 2369 36905
rect 2425 36849 2453 36905
rect 2509 36849 2537 36905
rect 1949 36825 2593 36849
rect 2005 36769 2033 36825
rect 2089 36769 2117 36825
rect 2173 36769 2201 36825
rect 2257 36769 2285 36825
rect 2341 36769 2369 36825
rect 2425 36769 2453 36825
rect 2509 36769 2537 36825
rect 1949 36745 2593 36769
rect 2005 36689 2033 36745
rect 2089 36689 2117 36745
rect 2173 36689 2201 36745
rect 2257 36689 2285 36745
rect 2341 36689 2369 36745
rect 2425 36689 2453 36745
rect 2509 36689 2537 36745
rect 1949 36665 2593 36689
rect 2005 36609 2033 36665
rect 2089 36609 2117 36665
rect 2173 36609 2201 36665
rect 2257 36609 2285 36665
rect 2341 36609 2369 36665
rect 2425 36609 2453 36665
rect 2509 36609 2537 36665
rect 1949 36585 2593 36609
rect 2005 36529 2033 36585
rect 2089 36529 2117 36585
rect 2173 36529 2201 36585
rect 2257 36529 2285 36585
rect 2341 36529 2369 36585
rect 2425 36529 2453 36585
rect 2509 36529 2537 36585
rect 1949 36505 2593 36529
rect 2005 36449 2033 36505
rect 2089 36449 2117 36505
rect 2173 36449 2201 36505
rect 2257 36449 2285 36505
rect 2341 36449 2369 36505
rect 2425 36449 2453 36505
rect 2509 36449 2537 36505
rect 1949 36425 2593 36449
rect 2005 36369 2033 36425
rect 2089 36369 2117 36425
rect 2173 36369 2201 36425
rect 2257 36369 2285 36425
rect 2341 36369 2369 36425
rect 2425 36369 2453 36425
rect 2509 36369 2537 36425
rect 1949 36345 2593 36369
rect 2005 36289 2033 36345
rect 2089 36289 2117 36345
rect 2173 36289 2201 36345
rect 2257 36289 2285 36345
rect 2341 36289 2369 36345
rect 2425 36289 2453 36345
rect 2509 36289 2537 36345
rect 1949 36265 2593 36289
rect 2005 36209 2033 36265
rect 2089 36209 2117 36265
rect 2173 36209 2201 36265
rect 2257 36209 2285 36265
rect 2341 36209 2369 36265
rect 2425 36209 2453 36265
rect 2509 36209 2537 36265
rect 1949 36185 2593 36209
rect 2005 36129 2033 36185
rect 2089 36129 2117 36185
rect 2173 36129 2201 36185
rect 2257 36129 2285 36185
rect 2341 36129 2369 36185
rect 2425 36129 2453 36185
rect 2509 36129 2537 36185
rect 1949 36105 2593 36129
rect 2005 36049 2033 36105
rect 2089 36049 2117 36105
rect 2173 36049 2201 36105
rect 2257 36049 2285 36105
rect 2341 36049 2369 36105
rect 2425 36049 2453 36105
rect 2509 36049 2537 36105
rect 1949 36025 2593 36049
rect 2005 35969 2033 36025
rect 2089 35969 2117 36025
rect 2173 35969 2201 36025
rect 2257 35969 2285 36025
rect 2341 35969 2369 36025
rect 2425 35969 2453 36025
rect 2509 35969 2537 36025
rect 1949 35945 2593 35969
rect 2005 35889 2033 35945
rect 2089 35889 2117 35945
rect 2173 35889 2201 35945
rect 2257 35889 2285 35945
rect 2341 35889 2369 35945
rect 2425 35889 2453 35945
rect 2509 35889 2537 35945
rect 1949 35865 2593 35889
rect 2005 35809 2033 35865
rect 2089 35809 2117 35865
rect 2173 35809 2201 35865
rect 2257 35809 2285 35865
rect 2341 35809 2369 35865
rect 2425 35809 2453 35865
rect 2509 35809 2537 35865
rect 1949 35785 2593 35809
rect 2005 35729 2033 35785
rect 2089 35729 2117 35785
rect 2173 35729 2201 35785
rect 2257 35729 2285 35785
rect 2341 35729 2369 35785
rect 2425 35729 2453 35785
rect 2509 35729 2537 35785
rect 1949 35705 2593 35729
rect 2005 35649 2033 35705
rect 2089 35649 2117 35705
rect 2173 35649 2201 35705
rect 2257 35649 2285 35705
rect 2341 35649 2369 35705
rect 2425 35649 2453 35705
rect 2509 35649 2537 35705
rect 1949 35625 2593 35649
rect 2005 35569 2033 35625
rect 2089 35569 2117 35625
rect 2173 35569 2201 35625
rect 2257 35569 2285 35625
rect 2341 35569 2369 35625
rect 2425 35569 2453 35625
rect 2509 35569 2537 35625
rect 1949 35545 2593 35569
rect 2005 35489 2033 35545
rect 2089 35489 2117 35545
rect 2173 35489 2201 35545
rect 2257 35489 2285 35545
rect 2341 35489 2369 35545
rect 2425 35489 2453 35545
rect 2509 35489 2537 35545
rect 1949 35465 2593 35489
rect 2005 35409 2033 35465
rect 2089 35409 2117 35465
rect 2173 35409 2201 35465
rect 2257 35409 2285 35465
rect 2341 35409 2369 35465
rect 2425 35409 2453 35465
rect 2509 35409 2537 35465
rect 1949 35385 2593 35409
rect 2005 35329 2033 35385
rect 2089 35329 2117 35385
rect 2173 35329 2201 35385
rect 2257 35329 2285 35385
rect 2341 35329 2369 35385
rect 2425 35329 2453 35385
rect 2509 35329 2537 35385
rect 1949 35305 2593 35329
rect 2005 35249 2033 35305
rect 2089 35249 2117 35305
rect 2173 35249 2201 35305
rect 2257 35249 2285 35305
rect 2341 35249 2369 35305
rect 2425 35249 2453 35305
rect 2509 35249 2537 35305
rect 1949 35225 2593 35249
rect 2005 35169 2033 35225
rect 2089 35169 2117 35225
rect 2173 35169 2201 35225
rect 2257 35169 2285 35225
rect 2341 35169 2369 35225
rect 2425 35169 2453 35225
rect 2509 35169 2537 35225
rect 1949 35145 2593 35169
rect 2005 35089 2033 35145
rect 2089 35089 2117 35145
rect 2173 35089 2201 35145
rect 2257 35089 2285 35145
rect 2341 35089 2369 35145
rect 2425 35089 2453 35145
rect 2509 35089 2537 35145
rect 1949 35065 2593 35089
rect 2005 35009 2033 35065
rect 2089 35009 2117 35065
rect 2173 35009 2201 35065
rect 2257 35009 2285 35065
rect 2341 35009 2369 35065
rect 2425 35009 2453 35065
rect 2509 35009 2537 35065
rect 1949 34985 2593 35009
rect 2005 34929 2033 34985
rect 2089 34929 2117 34985
rect 2173 34929 2201 34985
rect 2257 34929 2285 34985
rect 2341 34929 2369 34985
rect 2425 34929 2453 34985
rect 2509 34929 2537 34985
rect 1949 34905 2593 34929
rect 2005 34849 2033 34905
rect 2089 34849 2117 34905
rect 2173 34849 2201 34905
rect 2257 34849 2285 34905
rect 2341 34849 2369 34905
rect 2425 34849 2453 34905
rect 2509 34849 2537 34905
rect 1949 34825 2593 34849
rect 2005 34769 2033 34825
rect 2089 34769 2117 34825
rect 2173 34769 2201 34825
rect 2257 34769 2285 34825
rect 2341 34769 2369 34825
rect 2425 34769 2453 34825
rect 2509 34769 2537 34825
rect 1949 34745 2593 34769
rect 2005 34689 2033 34745
rect 2089 34689 2117 34745
rect 2173 34689 2201 34745
rect 2257 34689 2285 34745
rect 2341 34689 2369 34745
rect 2425 34689 2453 34745
rect 2509 34689 2537 34745
rect 1949 34665 2593 34689
rect 2005 34609 2033 34665
rect 2089 34609 2117 34665
rect 2173 34609 2201 34665
rect 2257 34609 2285 34665
rect 2341 34609 2369 34665
rect 2425 34609 2453 34665
rect 2509 34609 2537 34665
rect 1949 34585 2593 34609
rect 2005 34529 2033 34585
rect 2089 34529 2117 34585
rect 2173 34529 2201 34585
rect 2257 34529 2285 34585
rect 2341 34529 2369 34585
rect 2425 34529 2453 34585
rect 2509 34529 2537 34585
rect 1949 34505 2593 34529
rect 2005 34449 2033 34505
rect 2089 34449 2117 34505
rect 2173 34449 2201 34505
rect 2257 34449 2285 34505
rect 2341 34449 2369 34505
rect 2425 34449 2453 34505
rect 2509 34449 2537 34505
rect 1949 34425 2593 34449
rect 2005 34369 2033 34425
rect 2089 34369 2117 34425
rect 2173 34369 2201 34425
rect 2257 34369 2285 34425
rect 2341 34369 2369 34425
rect 2425 34369 2453 34425
rect 2509 34369 2537 34425
rect 1949 34345 2593 34369
rect 2005 34289 2033 34345
rect 2089 34289 2117 34345
rect 2173 34289 2201 34345
rect 2257 34289 2285 34345
rect 2341 34289 2369 34345
rect 2425 34289 2453 34345
rect 2509 34289 2537 34345
rect 1949 34265 2593 34289
rect 2005 34209 2033 34265
rect 2089 34209 2117 34265
rect 2173 34209 2201 34265
rect 2257 34209 2285 34265
rect 2341 34209 2369 34265
rect 2425 34209 2453 34265
rect 2509 34209 2537 34265
rect 1949 34185 2593 34209
rect 2005 34129 2033 34185
rect 2089 34129 2117 34185
rect 2173 34129 2201 34185
rect 2257 34129 2285 34185
rect 2341 34129 2369 34185
rect 2425 34129 2453 34185
rect 2509 34129 2537 34185
rect 1949 34105 2593 34129
rect 2005 34049 2033 34105
rect 2089 34049 2117 34105
rect 2173 34049 2201 34105
rect 2257 34049 2285 34105
rect 2341 34049 2369 34105
rect 2425 34049 2453 34105
rect 2509 34049 2537 34105
rect 1949 34025 2593 34049
rect 2005 33969 2033 34025
rect 2089 33969 2117 34025
rect 2173 33969 2201 34025
rect 2257 33969 2285 34025
rect 2341 33969 2369 34025
rect 2425 33969 2453 34025
rect 2509 33969 2537 34025
rect 1949 33945 2593 33969
rect 2005 33889 2033 33945
rect 2089 33889 2117 33945
rect 2173 33889 2201 33945
rect 2257 33889 2285 33945
rect 2341 33889 2369 33945
rect 2425 33889 2453 33945
rect 2509 33889 2537 33945
rect 1949 33865 2593 33889
rect 2005 33809 2033 33865
rect 2089 33809 2117 33865
rect 2173 33809 2201 33865
rect 2257 33809 2285 33865
rect 2341 33809 2369 33865
rect 2425 33809 2453 33865
rect 2509 33809 2537 33865
rect 1949 33785 2593 33809
rect 2005 33729 2033 33785
rect 2089 33729 2117 33785
rect 2173 33729 2201 33785
rect 2257 33729 2285 33785
rect 2341 33729 2369 33785
rect 2425 33729 2453 33785
rect 2509 33729 2537 33785
rect 1949 33705 2593 33729
rect 2005 33649 2033 33705
rect 2089 33649 2117 33705
rect 2173 33649 2201 33705
rect 2257 33649 2285 33705
rect 2341 33649 2369 33705
rect 2425 33649 2453 33705
rect 2509 33649 2537 33705
rect 1949 33625 2593 33649
rect 2005 33569 2033 33625
rect 2089 33569 2117 33625
rect 2173 33569 2201 33625
rect 2257 33569 2285 33625
rect 2341 33569 2369 33625
rect 2425 33569 2453 33625
rect 2509 33569 2537 33625
rect 1949 33545 2593 33569
rect 2005 33489 2033 33545
rect 2089 33489 2117 33545
rect 2173 33489 2201 33545
rect 2257 33489 2285 33545
rect 2341 33489 2369 33545
rect 2425 33489 2453 33545
rect 2509 33489 2537 33545
rect 1949 33465 2593 33489
rect 2005 33409 2033 33465
rect 2089 33409 2117 33465
rect 2173 33409 2201 33465
rect 2257 33409 2285 33465
rect 2341 33409 2369 33465
rect 2425 33409 2453 33465
rect 2509 33409 2537 33465
rect 1949 33385 2593 33409
rect 2005 33329 2033 33385
rect 2089 33329 2117 33385
rect 2173 33329 2201 33385
rect 2257 33329 2285 33385
rect 2341 33329 2369 33385
rect 2425 33329 2453 33385
rect 2509 33329 2537 33385
rect 1949 33305 2593 33329
rect 2005 33249 2033 33305
rect 2089 33249 2117 33305
rect 2173 33249 2201 33305
rect 2257 33249 2285 33305
rect 2341 33249 2369 33305
rect 2425 33249 2453 33305
rect 2509 33249 2537 33305
rect 1949 33225 2593 33249
rect 2005 33169 2033 33225
rect 2089 33169 2117 33225
rect 2173 33169 2201 33225
rect 2257 33169 2285 33225
rect 2341 33169 2369 33225
rect 2425 33169 2453 33225
rect 2509 33169 2537 33225
rect 1949 33145 2593 33169
rect 2005 33089 2033 33145
rect 2089 33089 2117 33145
rect 2173 33089 2201 33145
rect 2257 33089 2285 33145
rect 2341 33089 2369 33145
rect 2425 33089 2453 33145
rect 2509 33089 2537 33145
rect 1949 33065 2593 33089
rect 2005 33009 2033 33065
rect 2089 33009 2117 33065
rect 2173 33009 2201 33065
rect 2257 33009 2285 33065
rect 2341 33009 2369 33065
rect 2425 33009 2453 33065
rect 2509 33009 2537 33065
rect 1949 32985 2593 33009
rect 2005 32929 2033 32985
rect 2089 32929 2117 32985
rect 2173 32929 2201 32985
rect 2257 32929 2285 32985
rect 2341 32929 2369 32985
rect 2425 32929 2453 32985
rect 2509 32929 2537 32985
rect 1949 32905 2593 32929
rect 2005 32849 2033 32905
rect 2089 32849 2117 32905
rect 2173 32849 2201 32905
rect 2257 32849 2285 32905
rect 2341 32849 2369 32905
rect 2425 32849 2453 32905
rect 2509 32849 2537 32905
rect 1949 32825 2593 32849
rect 2005 32769 2033 32825
rect 2089 32769 2117 32825
rect 2173 32769 2201 32825
rect 2257 32769 2285 32825
rect 2341 32769 2369 32825
rect 2425 32769 2453 32825
rect 2509 32769 2537 32825
rect 1949 32745 2593 32769
rect 2005 32689 2033 32745
rect 2089 32689 2117 32745
rect 2173 32689 2201 32745
rect 2257 32689 2285 32745
rect 2341 32689 2369 32745
rect 2425 32689 2453 32745
rect 2509 32689 2537 32745
rect 1949 32664 2593 32689
rect 2005 32608 2033 32664
rect 2089 32608 2117 32664
rect 2173 32608 2201 32664
rect 2257 32608 2285 32664
rect 2341 32608 2369 32664
rect 2425 32608 2453 32664
rect 2509 32608 2537 32664
rect 1949 32583 2593 32608
rect 2005 32527 2033 32583
rect 2089 32527 2117 32583
rect 2173 32527 2201 32583
rect 2257 32527 2285 32583
rect 2341 32527 2369 32583
rect 2425 32527 2453 32583
rect 2509 32527 2537 32583
rect 1949 32502 2593 32527
rect 2005 32446 2033 32502
rect 2089 32446 2117 32502
rect 2173 32446 2201 32502
rect 2257 32446 2285 32502
rect 2341 32446 2369 32502
rect 2425 32446 2453 32502
rect 2509 32446 2537 32502
rect 1949 32421 2593 32446
rect 2005 32365 2033 32421
rect 2089 32365 2117 32421
rect 2173 32365 2201 32421
rect 2257 32365 2285 32421
rect 2341 32365 2369 32421
rect 2425 32365 2453 32421
rect 2509 32365 2537 32421
rect 1949 32340 2593 32365
rect 2005 32284 2033 32340
rect 2089 32284 2117 32340
rect 2173 32284 2201 32340
rect 2257 32284 2285 32340
rect 2341 32284 2369 32340
rect 2425 32284 2453 32340
rect 2509 32284 2537 32340
rect 1949 32259 2593 32284
rect 2005 32203 2033 32259
rect 2089 32203 2117 32259
rect 2173 32203 2201 32259
rect 2257 32203 2285 32259
rect 2341 32203 2369 32259
rect 2425 32203 2453 32259
rect 2509 32203 2537 32259
rect 1949 32178 2593 32203
rect 2005 32122 2033 32178
rect 2089 32122 2117 32178
rect 2173 32122 2201 32178
rect 2257 32122 2285 32178
rect 2341 32122 2369 32178
rect 2425 32122 2453 32178
rect 2509 32122 2537 32178
rect 1949 32097 2593 32122
rect 2005 32041 2033 32097
rect 2089 32041 2117 32097
rect 2173 32041 2201 32097
rect 2257 32041 2285 32097
rect 2341 32041 2369 32097
rect 2425 32041 2453 32097
rect 2509 32041 2537 32097
rect 1949 32016 2593 32041
rect 2005 31960 2033 32016
rect 2089 31960 2117 32016
rect 2173 31960 2201 32016
rect 2257 31960 2285 32016
rect 2341 31960 2369 32016
rect 2425 31960 2453 32016
rect 2509 31960 2537 32016
rect 1949 31935 2593 31960
rect 2005 31879 2033 31935
rect 2089 31879 2117 31935
rect 2173 31879 2201 31935
rect 2257 31879 2285 31935
rect 2341 31879 2369 31935
rect 2425 31879 2453 31935
rect 2509 31879 2537 31935
rect 1949 31854 2593 31879
rect 2005 31798 2033 31854
rect 2089 31798 2117 31854
rect 2173 31798 2201 31854
rect 2257 31798 2285 31854
rect 2341 31798 2369 31854
rect 2425 31798 2453 31854
rect 2509 31798 2537 31854
rect 1949 31773 2593 31798
rect 2005 31717 2033 31773
rect 2089 31717 2117 31773
rect 2173 31717 2201 31773
rect 2257 31717 2285 31773
rect 2341 31717 2369 31773
rect 2425 31717 2453 31773
rect 2509 31717 2537 31773
rect 1949 31692 2593 31717
rect 2005 31636 2033 31692
rect 2089 31636 2117 31692
rect 2173 31636 2201 31692
rect 2257 31636 2285 31692
rect 2341 31636 2369 31692
rect 2425 31636 2453 31692
rect 2509 31636 2537 31692
rect 1949 31611 2593 31636
rect 2005 31555 2033 31611
rect 2089 31555 2117 31611
rect 2173 31555 2201 31611
rect 2257 31555 2285 31611
rect 2341 31555 2369 31611
rect 2425 31555 2453 31611
rect 2509 31555 2537 31611
rect 1949 31530 2593 31555
rect 2005 31474 2033 31530
rect 2089 31474 2117 31530
rect 2173 31474 2201 31530
rect 2257 31474 2285 31530
rect 2341 31474 2369 31530
rect 2425 31474 2453 31530
rect 2509 31474 2537 31530
rect 1949 31449 2593 31474
rect 2005 31393 2033 31449
rect 2089 31393 2117 31449
rect 2173 31393 2201 31449
rect 2257 31393 2285 31449
rect 2341 31393 2369 31449
rect 2425 31393 2453 31449
rect 2509 31393 2537 31449
rect 1949 31368 2593 31393
rect 2005 31312 2033 31368
rect 2089 31312 2117 31368
rect 2173 31312 2201 31368
rect 2257 31312 2285 31368
rect 2341 31312 2369 31368
rect 2425 31312 2453 31368
rect 2509 31312 2537 31368
rect 1949 31287 2593 31312
rect 2005 31231 2033 31287
rect 2089 31231 2117 31287
rect 2173 31231 2201 31287
rect 2257 31231 2285 31287
rect 2341 31231 2369 31287
rect 2425 31231 2453 31287
rect 2509 31231 2537 31287
rect 1949 31206 2593 31231
rect 2005 31150 2033 31206
rect 2089 31150 2117 31206
rect 2173 31150 2201 31206
rect 2257 31150 2285 31206
rect 2341 31150 2369 31206
rect 2425 31150 2453 31206
rect 2509 31150 2537 31206
rect 1949 31125 2593 31150
rect 2005 31069 2033 31125
rect 2089 31069 2117 31125
rect 2173 31069 2201 31125
rect 2257 31069 2285 31125
rect 2341 31069 2369 31125
rect 2425 31069 2453 31125
rect 2509 31069 2537 31125
rect 1949 31044 2593 31069
rect 2005 30988 2033 31044
rect 2089 30988 2117 31044
rect 2173 30988 2201 31044
rect 2257 30988 2285 31044
rect 2341 30988 2369 31044
rect 2425 30988 2453 31044
rect 2509 30988 2537 31044
rect 1949 30963 2593 30988
rect 2005 30907 2033 30963
rect 2089 30907 2117 30963
rect 2173 30907 2201 30963
rect 2257 30907 2285 30963
rect 2341 30907 2369 30963
rect 2425 30907 2453 30963
rect 2509 30907 2537 30963
rect 1949 30882 2593 30907
rect 2005 30826 2033 30882
rect 2089 30826 2117 30882
rect 2173 30826 2201 30882
rect 2257 30826 2285 30882
rect 2341 30826 2369 30882
rect 2425 30826 2453 30882
rect 2509 30826 2537 30882
rect 1949 30801 2593 30826
rect 2005 30745 2033 30801
rect 2089 30745 2117 30801
rect 2173 30745 2201 30801
rect 2257 30745 2285 30801
rect 2341 30745 2369 30801
rect 2425 30745 2453 30801
rect 2509 30745 2537 30801
rect 1949 30720 2593 30745
rect 2005 30664 2033 30720
rect 2089 30664 2117 30720
rect 2173 30664 2201 30720
rect 2257 30664 2285 30720
rect 2341 30664 2369 30720
rect 2425 30664 2453 30720
rect 2509 30664 2537 30720
rect 1949 30639 2593 30664
rect 2005 30583 2033 30639
rect 2089 30583 2117 30639
rect 2173 30583 2201 30639
rect 2257 30583 2285 30639
rect 2341 30583 2369 30639
rect 2425 30583 2453 30639
rect 2509 30583 2537 30639
rect 1949 30558 2593 30583
rect 2005 30502 2033 30558
rect 2089 30502 2117 30558
rect 2173 30502 2201 30558
rect 2257 30502 2285 30558
rect 2341 30502 2369 30558
rect 2425 30502 2453 30558
rect 2509 30502 2537 30558
rect 1949 30477 2593 30502
rect 2005 30421 2033 30477
rect 2089 30421 2117 30477
rect 2173 30421 2201 30477
rect 2257 30421 2285 30477
rect 2341 30421 2369 30477
rect 2425 30421 2453 30477
rect 2509 30421 2537 30477
rect 1949 30396 2593 30421
rect 2005 30340 2033 30396
rect 2089 30340 2117 30396
rect 2173 30340 2201 30396
rect 2257 30340 2285 30396
rect 2341 30340 2369 30396
rect 2425 30340 2453 30396
rect 2509 30340 2537 30396
rect 1949 30315 2593 30340
rect 2005 30259 2033 30315
rect 2089 30259 2117 30315
rect 2173 30259 2201 30315
rect 2257 30259 2285 30315
rect 2341 30259 2369 30315
rect 2425 30259 2453 30315
rect 2509 30259 2537 30315
rect 1949 30234 2593 30259
rect 2005 30178 2033 30234
rect 2089 30178 2117 30234
rect 2173 30178 2201 30234
rect 2257 30178 2285 30234
rect 2341 30178 2369 30234
rect 2425 30178 2453 30234
rect 2509 30178 2537 30234
rect 1949 30169 2593 30178
rect 2900 34795 3491 34804
rect 2900 34739 2915 34795
rect 2971 34739 3001 34795
rect 3057 34739 3087 34795
rect 3143 34739 3173 34795
rect 3229 34739 3259 34795
rect 3315 34739 3345 34795
rect 3401 34739 3431 34795
rect 3487 34739 3491 34795
rect 2900 34715 3491 34739
rect 2900 34659 2915 34715
rect 2971 34659 3001 34715
rect 3057 34659 3087 34715
rect 3143 34659 3173 34715
rect 3229 34659 3259 34715
rect 3315 34659 3345 34715
rect 3401 34659 3431 34715
rect 3487 34659 3491 34715
rect 2900 34635 3491 34659
rect 2900 34579 2915 34635
rect 2971 34579 3001 34635
rect 3057 34579 3087 34635
rect 3143 34579 3173 34635
rect 3229 34579 3259 34635
rect 3315 34579 3345 34635
rect 3401 34579 3431 34635
rect 3487 34579 3491 34635
rect 2900 34555 3491 34579
rect 2900 34499 2915 34555
rect 2971 34499 3001 34555
rect 3057 34499 3087 34555
rect 3143 34499 3173 34555
rect 3229 34499 3259 34555
rect 3315 34499 3345 34555
rect 3401 34499 3431 34555
rect 3487 34499 3491 34555
rect 2900 34475 3491 34499
rect 2900 34419 2915 34475
rect 2971 34419 3001 34475
rect 3057 34419 3087 34475
rect 3143 34419 3173 34475
rect 3229 34419 3259 34475
rect 3315 34419 3345 34475
rect 3401 34419 3431 34475
rect 3487 34419 3491 34475
rect 2900 34395 3491 34419
rect 2900 34339 2915 34395
rect 2971 34339 3001 34395
rect 3057 34339 3087 34395
rect 3143 34339 3173 34395
rect 3229 34339 3259 34395
rect 3315 34339 3345 34395
rect 3401 34339 3431 34395
rect 3487 34339 3491 34395
rect 2900 34315 3491 34339
rect 2900 34259 2915 34315
rect 2971 34259 3001 34315
rect 3057 34259 3087 34315
rect 3143 34259 3173 34315
rect 3229 34259 3259 34315
rect 3315 34259 3345 34315
rect 3401 34259 3431 34315
rect 3487 34259 3491 34315
rect 2900 34235 3491 34259
rect 2900 34179 2915 34235
rect 2971 34179 3001 34235
rect 3057 34179 3087 34235
rect 3143 34179 3173 34235
rect 3229 34179 3259 34235
rect 3315 34179 3345 34235
rect 3401 34179 3431 34235
rect 3487 34179 3491 34235
rect 2900 34155 3491 34179
rect 2900 34099 2915 34155
rect 2971 34099 3001 34155
rect 3057 34099 3087 34155
rect 3143 34099 3173 34155
rect 3229 34099 3259 34155
rect 3315 34099 3345 34155
rect 3401 34099 3431 34155
rect 3487 34099 3491 34155
rect 2900 34075 3491 34099
rect 2900 34019 2915 34075
rect 2971 34019 3001 34075
rect 3057 34019 3087 34075
rect 3143 34019 3173 34075
rect 3229 34019 3259 34075
rect 3315 34019 3345 34075
rect 3401 34019 3431 34075
rect 3487 34019 3491 34075
rect 2900 33995 3491 34019
rect 2900 33939 2915 33995
rect 2971 33939 3001 33995
rect 3057 33939 3087 33995
rect 3143 33939 3173 33995
rect 3229 33939 3259 33995
rect 3315 33939 3345 33995
rect 3401 33939 3431 33995
rect 3487 33939 3491 33995
rect 2900 33915 3491 33939
rect 2900 33859 2915 33915
rect 2971 33859 3001 33915
rect 3057 33859 3087 33915
rect 3143 33859 3173 33915
rect 3229 33859 3259 33915
rect 3315 33859 3345 33915
rect 3401 33859 3431 33915
rect 3487 33859 3491 33915
rect 2900 33835 3491 33859
rect 2900 33779 2915 33835
rect 2971 33779 3001 33835
rect 3057 33779 3087 33835
rect 3143 33779 3173 33835
rect 3229 33779 3259 33835
rect 3315 33779 3345 33835
rect 3401 33779 3431 33835
rect 3487 33779 3491 33835
rect 2900 33755 3491 33779
rect 2900 33699 2915 33755
rect 2971 33699 3001 33755
rect 3057 33699 3087 33755
rect 3143 33699 3173 33755
rect 3229 33699 3259 33755
rect 3315 33699 3345 33755
rect 3401 33699 3431 33755
rect 3487 33699 3491 33755
rect 2900 33675 3491 33699
rect 2900 33619 2915 33675
rect 2971 33619 3001 33675
rect 3057 33619 3087 33675
rect 3143 33619 3173 33675
rect 3229 33619 3259 33675
rect 3315 33619 3345 33675
rect 3401 33619 3431 33675
rect 3487 33619 3491 33675
rect 2900 33595 3491 33619
rect 2900 33539 2915 33595
rect 2971 33539 3001 33595
rect 3057 33539 3087 33595
rect 3143 33539 3173 33595
rect 3229 33539 3259 33595
rect 3315 33539 3345 33595
rect 3401 33539 3431 33595
rect 3487 33539 3491 33595
rect 2900 33515 3491 33539
rect 2900 33459 2915 33515
rect 2971 33459 3001 33515
rect 3057 33459 3087 33515
rect 3143 33459 3173 33515
rect 3229 33459 3259 33515
rect 3315 33459 3345 33515
rect 3401 33459 3431 33515
rect 3487 33459 3491 33515
rect 2900 33435 3491 33459
rect 2900 33379 2915 33435
rect 2971 33379 3001 33435
rect 3057 33379 3087 33435
rect 3143 33379 3173 33435
rect 3229 33379 3259 33435
rect 3315 33379 3345 33435
rect 3401 33379 3431 33435
rect 3487 33379 3491 33435
rect 2900 33355 3491 33379
rect 2900 33299 2915 33355
rect 2971 33299 3001 33355
rect 3057 33299 3087 33355
rect 3143 33299 3173 33355
rect 3229 33299 3259 33355
rect 3315 33299 3345 33355
rect 3401 33299 3431 33355
rect 3487 33299 3491 33355
rect 2900 33275 3491 33299
rect 2900 33219 2915 33275
rect 2971 33219 3001 33275
rect 3057 33219 3087 33275
rect 3143 33219 3173 33275
rect 3229 33219 3259 33275
rect 3315 33219 3345 33275
rect 3401 33219 3431 33275
rect 3487 33219 3491 33275
rect 2900 33195 3491 33219
rect 2900 33139 2915 33195
rect 2971 33139 3001 33195
rect 3057 33139 3087 33195
rect 3143 33139 3173 33195
rect 3229 33139 3259 33195
rect 3315 33139 3345 33195
rect 3401 33139 3431 33195
rect 3487 33139 3491 33195
rect 2900 33115 3491 33139
rect 2900 33059 2915 33115
rect 2971 33059 3001 33115
rect 3057 33059 3087 33115
rect 3143 33059 3173 33115
rect 3229 33059 3259 33115
rect 3315 33059 3345 33115
rect 3401 33059 3431 33115
rect 3487 33059 3491 33115
rect 2900 33035 3491 33059
rect 2900 32979 2915 33035
rect 2971 32979 3001 33035
rect 3057 32979 3087 33035
rect 3143 32979 3173 33035
rect 3229 32979 3259 33035
rect 3315 32979 3345 33035
rect 3401 32979 3431 33035
rect 3487 32979 3491 33035
rect 2900 32955 3491 32979
rect 2900 32899 2915 32955
rect 2971 32899 3001 32955
rect 3057 32899 3087 32955
rect 3143 32899 3173 32955
rect 3229 32899 3259 32955
rect 3315 32899 3345 32955
rect 3401 32899 3431 32955
rect 3487 32899 3491 32955
rect 2900 32875 3491 32899
rect 2900 32819 2915 32875
rect 2971 32819 3001 32875
rect 3057 32819 3087 32875
rect 3143 32819 3173 32875
rect 3229 32819 3259 32875
rect 3315 32819 3345 32875
rect 3401 32819 3431 32875
rect 3487 32819 3491 32875
rect 2900 32795 3491 32819
rect 2900 32739 2915 32795
rect 2971 32739 3001 32795
rect 3057 32739 3087 32795
rect 3143 32739 3173 32795
rect 3229 32739 3259 32795
rect 3315 32739 3345 32795
rect 3401 32739 3431 32795
rect 3487 32739 3491 32795
rect 2900 32715 3491 32739
rect 2900 32659 2915 32715
rect 2971 32659 3001 32715
rect 3057 32659 3087 32715
rect 3143 32659 3173 32715
rect 3229 32659 3259 32715
rect 3315 32659 3345 32715
rect 3401 32659 3431 32715
rect 3487 32659 3491 32715
rect 2900 32635 3491 32659
rect 2900 32579 2915 32635
rect 2971 32579 3001 32635
rect 3057 32579 3087 32635
rect 3143 32579 3173 32635
rect 3229 32579 3259 32635
rect 3315 32579 3345 32635
rect 3401 32579 3431 32635
rect 3487 32579 3491 32635
rect 2900 32555 3491 32579
rect 2900 32499 2915 32555
rect 2971 32499 3001 32555
rect 3057 32499 3087 32555
rect 3143 32499 3173 32555
rect 3229 32499 3259 32555
rect 3315 32499 3345 32555
rect 3401 32499 3431 32555
rect 3487 32499 3491 32555
rect 2900 32475 3491 32499
rect 2900 32419 2915 32475
rect 2971 32419 3001 32475
rect 3057 32419 3087 32475
rect 3143 32419 3173 32475
rect 3229 32419 3259 32475
rect 3315 32419 3345 32475
rect 3401 32419 3431 32475
rect 3487 32419 3491 32475
rect 2900 32395 3491 32419
rect 2900 32339 2915 32395
rect 2971 32339 3001 32395
rect 3057 32339 3087 32395
rect 3143 32339 3173 32395
rect 3229 32339 3259 32395
rect 3315 32339 3345 32395
rect 3401 32339 3431 32395
rect 3487 32339 3491 32395
rect 2900 32315 3491 32339
rect 2900 32259 2915 32315
rect 2971 32259 3001 32315
rect 3057 32259 3087 32315
rect 3143 32259 3173 32315
rect 3229 32259 3259 32315
rect 3315 32259 3345 32315
rect 3401 32259 3431 32315
rect 3487 32259 3491 32315
rect 2900 32235 3491 32259
rect 2900 32179 2915 32235
rect 2971 32179 3001 32235
rect 3057 32179 3087 32235
rect 3143 32179 3173 32235
rect 3229 32179 3259 32235
rect 3315 32179 3345 32235
rect 3401 32179 3431 32235
rect 3487 32179 3491 32235
rect 2900 32155 3491 32179
rect 2900 32099 2915 32155
rect 2971 32099 3001 32155
rect 3057 32099 3087 32155
rect 3143 32099 3173 32155
rect 3229 32099 3259 32155
rect 3315 32099 3345 32155
rect 3401 32099 3431 32155
rect 3487 32099 3491 32155
rect 2900 32075 3491 32099
rect 2900 32019 2915 32075
rect 2971 32019 3001 32075
rect 3057 32019 3087 32075
rect 3143 32019 3173 32075
rect 3229 32019 3259 32075
rect 3315 32019 3345 32075
rect 3401 32019 3431 32075
rect 3487 32019 3491 32075
rect 2900 31995 3491 32019
rect 2900 31939 2915 31995
rect 2971 31939 3001 31995
rect 3057 31939 3087 31995
rect 3143 31939 3173 31995
rect 3229 31939 3259 31995
rect 3315 31939 3345 31995
rect 3401 31939 3431 31995
rect 3487 31939 3491 31995
rect 2900 31915 3491 31939
rect 2900 31859 2915 31915
rect 2971 31859 3001 31915
rect 3057 31859 3087 31915
rect 3143 31859 3173 31915
rect 3229 31859 3259 31915
rect 3315 31859 3345 31915
rect 3401 31859 3431 31915
rect 3487 31859 3491 31915
rect 2900 31835 3491 31859
rect 2900 31779 2915 31835
rect 2971 31779 3001 31835
rect 3057 31779 3087 31835
rect 3143 31779 3173 31835
rect 3229 31779 3259 31835
rect 3315 31779 3345 31835
rect 3401 31779 3431 31835
rect 3487 31779 3491 31835
rect 2900 31755 3491 31779
rect 2900 31699 2915 31755
rect 2971 31699 3001 31755
rect 3057 31699 3087 31755
rect 3143 31699 3173 31755
rect 3229 31699 3259 31755
rect 3315 31699 3345 31755
rect 3401 31699 3431 31755
rect 3487 31699 3491 31755
rect 2900 31675 3491 31699
rect 2900 31619 2915 31675
rect 2971 31619 3001 31675
rect 3057 31619 3087 31675
rect 3143 31619 3173 31675
rect 3229 31619 3259 31675
rect 3315 31619 3345 31675
rect 3401 31619 3431 31675
rect 3487 31619 3491 31675
rect 2900 31595 3491 31619
rect 2900 31539 2915 31595
rect 2971 31539 3001 31595
rect 3057 31539 3087 31595
rect 3143 31539 3173 31595
rect 3229 31539 3259 31595
rect 3315 31539 3345 31595
rect 3401 31539 3431 31595
rect 3487 31539 3491 31595
rect 2900 31515 3491 31539
rect 2900 31459 2915 31515
rect 2971 31459 3001 31515
rect 3057 31459 3087 31515
rect 3143 31459 3173 31515
rect 3229 31459 3259 31515
rect 3315 31459 3345 31515
rect 3401 31459 3431 31515
rect 3487 31459 3491 31515
rect 2900 31435 3491 31459
rect 2900 31379 2915 31435
rect 2971 31379 3001 31435
rect 3057 31379 3087 31435
rect 3143 31379 3173 31435
rect 3229 31379 3259 31435
rect 3315 31379 3345 31435
rect 3401 31379 3431 31435
rect 3487 31379 3491 31435
rect 2900 31355 3491 31379
rect 2900 31299 2915 31355
rect 2971 31299 3001 31355
rect 3057 31299 3087 31355
rect 3143 31299 3173 31355
rect 3229 31299 3259 31355
rect 3315 31299 3345 31355
rect 3401 31299 3431 31355
rect 3487 31299 3491 31355
rect 2900 31275 3491 31299
rect 2900 31219 2915 31275
rect 2971 31219 3001 31275
rect 3057 31219 3087 31275
rect 3143 31219 3173 31275
rect 3229 31219 3259 31275
rect 3315 31219 3345 31275
rect 3401 31219 3431 31275
rect 3487 31219 3491 31275
rect 2900 31195 3491 31219
rect 2900 31139 2915 31195
rect 2971 31139 3001 31195
rect 3057 31139 3087 31195
rect 3143 31139 3173 31195
rect 3229 31139 3259 31195
rect 3315 31139 3345 31195
rect 3401 31139 3431 31195
rect 3487 31139 3491 31195
rect 2900 31115 3491 31139
rect 2900 31059 2915 31115
rect 2971 31059 3001 31115
rect 3057 31059 3087 31115
rect 3143 31059 3173 31115
rect 3229 31059 3259 31115
rect 3315 31059 3345 31115
rect 3401 31059 3431 31115
rect 3487 31059 3491 31115
rect 2900 31035 3491 31059
rect 2900 30979 2915 31035
rect 2971 30979 3001 31035
rect 3057 30979 3087 31035
rect 3143 30979 3173 31035
rect 3229 30979 3259 31035
rect 3315 30979 3345 31035
rect 3401 30979 3431 31035
rect 3487 30979 3491 31035
rect 2900 30955 3491 30979
rect 2900 30899 2915 30955
rect 2971 30899 3001 30955
rect 3057 30899 3087 30955
rect 3143 30899 3173 30955
rect 3229 30899 3259 30955
rect 3315 30899 3345 30955
rect 3401 30899 3431 30955
rect 3487 30899 3491 30955
rect 2900 30875 3491 30899
rect 2900 30819 2915 30875
rect 2971 30819 3001 30875
rect 3057 30819 3087 30875
rect 3143 30819 3173 30875
rect 3229 30819 3259 30875
rect 3315 30819 3345 30875
rect 3401 30819 3431 30875
rect 3487 30819 3491 30875
rect 2900 30795 3491 30819
rect 2900 30739 2915 30795
rect 2971 30739 3001 30795
rect 3057 30739 3087 30795
rect 3143 30739 3173 30795
rect 3229 30739 3259 30795
rect 3315 30739 3345 30795
rect 3401 30739 3431 30795
rect 3487 30739 3491 30795
rect 2900 30715 3491 30739
rect 2900 30659 2915 30715
rect 2971 30659 3001 30715
rect 3057 30659 3087 30715
rect 3143 30659 3173 30715
rect 3229 30659 3259 30715
rect 3315 30659 3345 30715
rect 3401 30659 3431 30715
rect 3487 30659 3491 30715
rect 2900 30635 3491 30659
rect 2900 30579 2915 30635
rect 2971 30579 3001 30635
rect 3057 30579 3087 30635
rect 3143 30579 3173 30635
rect 3229 30579 3259 30635
rect 3315 30579 3345 30635
rect 3401 30579 3431 30635
rect 3487 30579 3491 30635
rect 2900 30555 3491 30579
rect 2900 30499 2915 30555
rect 2971 30499 3001 30555
rect 3057 30499 3087 30555
rect 3143 30499 3173 30555
rect 3229 30499 3259 30555
rect 3315 30499 3345 30555
rect 3401 30499 3431 30555
rect 3487 30499 3491 30555
rect 2900 30475 3491 30499
rect 2900 30419 2915 30475
rect 2971 30419 3001 30475
rect 3057 30419 3087 30475
rect 3143 30419 3173 30475
rect 3229 30419 3259 30475
rect 3315 30419 3345 30475
rect 3401 30419 3431 30475
rect 3487 30419 3491 30475
rect 2900 30395 3491 30419
rect 2900 30339 2915 30395
rect 2971 30339 3001 30395
rect 3057 30339 3087 30395
rect 3143 30339 3173 30395
rect 3229 30339 3259 30395
rect 3315 30339 3345 30395
rect 3401 30339 3431 30395
rect 3487 30339 3491 30395
rect 2900 30315 3491 30339
rect 2900 30259 2915 30315
rect 2971 30259 3001 30315
rect 3057 30259 3087 30315
rect 3143 30259 3173 30315
rect 3229 30259 3259 30315
rect 3315 30259 3345 30315
rect 3401 30259 3431 30315
rect 3487 30259 3491 30315
rect 2900 30235 3491 30259
rect 2900 30179 2915 30235
rect 2971 30179 3001 30235
rect 3057 30179 3087 30235
rect 3143 30179 3173 30235
rect 3229 30179 3259 30235
rect 3315 30179 3345 30235
rect 3401 30179 3431 30235
rect 3487 30179 3491 30235
rect 2900 30155 3491 30179
rect 2900 30099 2915 30155
rect 2971 30099 3001 30155
rect 3057 30099 3087 30155
rect 3143 30099 3173 30155
rect 3229 30099 3259 30155
rect 3315 30099 3345 30155
rect 3401 30099 3431 30155
rect 3487 30099 3491 30155
rect 2900 30075 3491 30099
rect 2900 30019 2915 30075
rect 2971 30019 3001 30075
rect 3057 30019 3087 30075
rect 3143 30019 3173 30075
rect 3229 30019 3259 30075
rect 3315 30019 3345 30075
rect 3401 30019 3431 30075
rect 3487 30019 3491 30075
rect 2900 30010 3491 30019
tri 4501 29761 4535 29795 se
rect 4535 29761 4587 30399
rect 3878 29709 4587 29761
tri 3844 29403 3878 29437 se
rect 3878 29403 3930 29709
tri 3930 29675 3964 29709 nw
tri 4685 29675 4711 29701 se
rect 4711 29675 4763 37104
tri 4677 29667 4685 29675 se
rect 4685 29667 4763 29675
rect 1938 28963 2598 29376
rect 3802 29351 3808 29403
rect 3860 29351 3872 29403
rect 3924 29351 3930 29403
rect 4008 29615 4763 29667
rect 4008 29593 4072 29615
tri 4072 29593 4094 29615 nw
tri 4006 29351 4008 29353 se
rect 4008 29351 4060 29593
tri 4060 29581 4072 29593 nw
tri 4818 29581 4830 29593 se
rect 4830 29581 4882 37107
rect 6900 37094 6903 37150
rect 6959 37094 6993 37150
rect 7049 37094 7083 37150
rect 7139 37094 7173 37150
rect 7229 37094 7263 37150
rect 7319 37094 7353 37150
rect 7409 37094 7443 37150
rect 7499 37094 7502 37150
rect 6900 37070 7502 37094
rect 6900 37014 6903 37070
rect 6959 37014 6993 37070
rect 7049 37014 7083 37070
rect 7139 37014 7173 37070
rect 7229 37014 7263 37070
rect 7319 37014 7353 37070
rect 7409 37014 7443 37070
rect 7499 37014 7502 37070
rect 6900 36990 7502 37014
rect 6900 36934 6903 36990
rect 6959 36934 6993 36990
rect 7049 36934 7083 36990
rect 7139 36934 7173 36990
rect 7229 36934 7263 36990
rect 7319 36934 7353 36990
rect 7409 36934 7443 36990
rect 7499 36934 7502 36990
rect 6900 36910 7502 36934
rect 6900 36854 6903 36910
rect 6959 36854 6993 36910
rect 7049 36854 7083 36910
rect 7139 36854 7173 36910
rect 7229 36854 7263 36910
rect 7319 36854 7353 36910
rect 7409 36854 7443 36910
rect 7499 36854 7502 36910
rect 6900 36830 7502 36854
rect 6900 36774 6903 36830
rect 6959 36774 6993 36830
rect 7049 36774 7083 36830
rect 7139 36774 7173 36830
rect 7229 36774 7263 36830
rect 7319 36774 7353 36830
rect 7409 36774 7443 36830
rect 7499 36774 7502 36830
rect 6900 36750 7502 36774
rect 6900 36694 6903 36750
rect 6959 36694 6993 36750
rect 7049 36694 7083 36750
rect 7139 36694 7173 36750
rect 7229 36694 7263 36750
rect 7319 36694 7353 36750
rect 7409 36694 7443 36750
rect 7499 36694 7502 36750
rect 6900 36670 7502 36694
rect 6900 36614 6903 36670
rect 6959 36614 6993 36670
rect 7049 36614 7083 36670
rect 7139 36614 7173 36670
rect 7229 36614 7263 36670
rect 7319 36614 7353 36670
rect 7409 36614 7443 36670
rect 7499 36614 7502 36670
rect 6900 36590 7502 36614
rect 6900 36534 6903 36590
rect 6959 36534 6993 36590
rect 7049 36534 7083 36590
rect 7139 36534 7173 36590
rect 7229 36534 7263 36590
rect 7319 36534 7353 36590
rect 7409 36534 7443 36590
rect 7499 36534 7502 36590
rect 6900 36510 7502 36534
rect 6900 36454 6903 36510
rect 6959 36454 6993 36510
rect 7049 36454 7083 36510
rect 7139 36454 7173 36510
rect 7229 36454 7263 36510
rect 7319 36454 7353 36510
rect 7409 36454 7443 36510
rect 7499 36454 7502 36510
rect 6900 36430 7502 36454
rect 6900 36374 6903 36430
rect 6959 36374 6993 36430
rect 7049 36374 7083 36430
rect 7139 36374 7173 36430
rect 7229 36374 7263 36430
rect 7319 36374 7353 36430
rect 7409 36374 7443 36430
rect 7499 36374 7502 36430
rect 6900 36350 7502 36374
rect 6900 36294 6903 36350
rect 6959 36294 6993 36350
rect 7049 36294 7083 36350
rect 7139 36294 7173 36350
rect 7229 36294 7263 36350
rect 7319 36294 7353 36350
rect 7409 36294 7443 36350
rect 7499 36294 7502 36350
rect 6900 36270 7502 36294
rect 6900 36214 6903 36270
rect 6959 36214 6993 36270
rect 7049 36214 7083 36270
rect 7139 36214 7173 36270
rect 7229 36214 7263 36270
rect 7319 36214 7353 36270
rect 7409 36214 7443 36270
rect 7499 36214 7502 36270
rect 6900 36190 7502 36214
rect 6900 36134 6903 36190
rect 6959 36134 6993 36190
rect 7049 36134 7083 36190
rect 7139 36134 7173 36190
rect 7229 36134 7263 36190
rect 7319 36134 7353 36190
rect 7409 36134 7443 36190
rect 7499 36134 7502 36190
rect 6900 36110 7502 36134
rect 6900 36054 6903 36110
rect 6959 36054 6993 36110
rect 7049 36054 7083 36110
rect 7139 36054 7173 36110
rect 7229 36054 7263 36110
rect 7319 36054 7353 36110
rect 7409 36054 7443 36110
rect 7499 36054 7502 36110
rect 6900 36030 7502 36054
rect 6900 35974 6903 36030
rect 6959 35974 6993 36030
rect 7049 35974 7083 36030
rect 7139 35974 7173 36030
rect 7229 35974 7263 36030
rect 7319 35974 7353 36030
rect 7409 35974 7443 36030
rect 7499 35974 7502 36030
rect 6900 35950 7502 35974
rect 6900 35894 6903 35950
rect 6959 35894 6993 35950
rect 7049 35894 7083 35950
rect 7139 35894 7173 35950
rect 7229 35894 7263 35950
rect 7319 35894 7353 35950
rect 7409 35894 7443 35950
rect 7499 35894 7502 35950
rect 6900 35870 7502 35894
rect 6900 35814 6903 35870
rect 6959 35814 6993 35870
rect 7049 35814 7083 35870
rect 7139 35814 7173 35870
rect 7229 35814 7263 35870
rect 7319 35814 7353 35870
rect 7409 35814 7443 35870
rect 7499 35814 7502 35870
rect 6900 35790 7502 35814
rect 6900 35734 6903 35790
rect 6959 35734 6993 35790
rect 7049 35734 7083 35790
rect 7139 35734 7173 35790
rect 7229 35734 7263 35790
rect 7319 35734 7353 35790
rect 7409 35734 7443 35790
rect 7499 35734 7502 35790
tri 4931 35517 5005 35591 se
rect 5005 35569 5057 35722
tri 5005 35517 5057 35569 nw
rect 6900 35710 7502 35734
rect 6900 35654 6903 35710
rect 6959 35654 6993 35710
rect 7049 35654 7083 35710
rect 7139 35654 7173 35710
rect 7229 35654 7263 35710
rect 7319 35654 7353 35710
rect 7409 35654 7443 35710
rect 7499 35654 7502 35710
rect 6900 35630 7502 35654
rect 6900 35574 6903 35630
rect 6959 35574 6993 35630
rect 7049 35574 7083 35630
rect 7139 35574 7173 35630
rect 7229 35574 7263 35630
rect 7319 35574 7353 35630
rect 7409 35574 7443 35630
rect 7499 35574 7502 35630
rect 6900 35550 7502 35574
tri 4796 29559 4818 29581 se
rect 4818 29559 4882 29581
tri 3974 29319 4006 29351 se
rect 4006 29319 4060 29351
rect 3932 29267 3938 29319
rect 3990 29267 4002 29319
rect 4054 29267 4060 29319
rect 4115 29507 4882 29559
tri 4921 35507 4931 35517 se
rect 4931 35507 4995 35517
tri 4995 35507 5005 35517 nw
tri 4113 29267 4115 29269 se
rect 4115 29267 4167 29507
tri 4167 29473 4201 29507 nw
tri 4909 29473 4921 29485 se
rect 4921 29473 4973 35507
tri 4973 35485 4995 35507 nw
rect 6900 35494 6903 35550
rect 6959 35494 6993 35550
rect 7049 35494 7083 35550
rect 7139 35494 7173 35550
rect 7229 35494 7263 35550
rect 7319 35494 7353 35550
rect 7409 35494 7443 35550
rect 7499 35494 7502 35550
rect 6900 35470 7502 35494
rect 6900 35414 6903 35470
rect 6959 35414 6993 35470
rect 7049 35414 7083 35470
rect 7139 35414 7173 35470
rect 7229 35414 7263 35470
rect 7319 35414 7353 35470
rect 7409 35414 7443 35470
rect 7499 35414 7502 35470
rect 6900 35390 7502 35414
rect 6900 35334 6903 35390
rect 6959 35334 6993 35390
rect 7049 35334 7083 35390
rect 7139 35334 7173 35390
rect 7229 35334 7263 35390
rect 7319 35334 7353 35390
rect 7409 35334 7443 35390
rect 7499 35334 7502 35390
rect 6900 35310 7502 35334
rect 6900 35254 6903 35310
rect 6959 35254 6993 35310
rect 7049 35254 7083 35310
rect 7139 35254 7173 35310
rect 7229 35254 7263 35310
rect 7319 35254 7353 35310
rect 7409 35254 7443 35310
rect 7499 35254 7502 35310
rect 6900 35230 7502 35254
rect 6900 35174 6903 35230
rect 6959 35174 6993 35230
rect 7049 35174 7083 35230
rect 7139 35174 7173 35230
rect 7229 35174 7263 35230
rect 7319 35174 7353 35230
rect 7409 35174 7443 35230
rect 7499 35174 7502 35230
rect 6900 35150 7502 35174
rect 6900 35094 6903 35150
rect 6959 35094 6993 35150
rect 7049 35094 7083 35150
rect 7139 35094 7173 35150
rect 7229 35094 7263 35150
rect 7319 35094 7353 35150
rect 7409 35094 7443 35150
rect 7499 35094 7502 35150
rect 6900 35070 7502 35094
rect 6900 35014 6903 35070
rect 6959 35014 6993 35070
rect 7049 35014 7083 35070
rect 7139 35014 7173 35070
rect 7229 35014 7263 35070
rect 7319 35014 7353 35070
rect 7409 35014 7443 35070
rect 7499 35014 7502 35070
rect 6900 34990 7502 35014
rect 6900 34934 6903 34990
rect 6959 34934 6993 34990
rect 7049 34934 7083 34990
rect 7139 34934 7173 34990
rect 7229 34934 7263 34990
rect 7319 34934 7353 34990
rect 7409 34934 7443 34990
rect 7499 34934 7502 34990
rect 6900 34910 7502 34934
rect 6900 34854 6903 34910
rect 6959 34854 6993 34910
rect 7049 34854 7083 34910
rect 7139 34854 7173 34910
rect 7229 34854 7263 34910
rect 7319 34854 7353 34910
rect 7409 34854 7443 34910
rect 7499 34854 7502 34910
rect 6900 34830 7502 34854
rect 5901 34795 6481 34804
rect 5901 34739 5905 34795
rect 5961 34739 5991 34795
rect 6047 34739 6077 34795
rect 6133 34739 6163 34795
rect 6219 34739 6249 34795
rect 6305 34739 6335 34795
rect 6391 34739 6421 34795
rect 6477 34739 6481 34795
rect 5901 34715 6481 34739
rect 5901 34659 5905 34715
rect 5961 34659 5991 34715
rect 6047 34659 6077 34715
rect 6133 34659 6163 34715
rect 6219 34659 6249 34715
rect 6305 34659 6335 34715
rect 6391 34659 6421 34715
rect 6477 34659 6481 34715
rect 5901 34635 6481 34659
rect 5901 34579 5905 34635
rect 5961 34579 5991 34635
rect 6047 34579 6077 34635
rect 6133 34579 6163 34635
rect 6219 34579 6249 34635
rect 6305 34579 6335 34635
rect 6391 34579 6421 34635
rect 6477 34579 6481 34635
rect 5901 34555 6481 34579
rect 5901 34499 5905 34555
rect 5961 34499 5991 34555
rect 6047 34499 6077 34555
rect 6133 34499 6163 34555
rect 6219 34499 6249 34555
rect 6305 34499 6335 34555
rect 6391 34499 6421 34555
rect 6477 34499 6481 34555
rect 5901 34475 6481 34499
rect 5901 34419 5905 34475
rect 5961 34419 5991 34475
rect 6047 34419 6077 34475
rect 6133 34419 6163 34475
rect 6219 34419 6249 34475
rect 6305 34419 6335 34475
rect 6391 34419 6421 34475
rect 6477 34419 6481 34475
rect 5901 34395 6481 34419
rect 5901 34339 5905 34395
rect 5961 34339 5991 34395
rect 6047 34339 6077 34395
rect 6133 34339 6163 34395
rect 6219 34339 6249 34395
rect 6305 34339 6335 34395
rect 6391 34339 6421 34395
rect 6477 34339 6481 34395
rect 5901 34315 6481 34339
rect 5901 34259 5905 34315
rect 5961 34259 5991 34315
rect 6047 34259 6077 34315
rect 6133 34259 6163 34315
rect 6219 34259 6249 34315
rect 6305 34259 6335 34315
rect 6391 34259 6421 34315
rect 6477 34259 6481 34315
rect 5901 34235 6481 34259
rect 5901 34179 5905 34235
rect 5961 34179 5991 34235
rect 6047 34179 6077 34235
rect 6133 34179 6163 34235
rect 6219 34179 6249 34235
rect 6305 34179 6335 34235
rect 6391 34179 6421 34235
rect 6477 34179 6481 34235
rect 5901 34155 6481 34179
rect 5901 34099 5905 34155
rect 5961 34099 5991 34155
rect 6047 34099 6077 34155
rect 6133 34099 6163 34155
rect 6219 34099 6249 34155
rect 6305 34099 6335 34155
rect 6391 34099 6421 34155
rect 6477 34099 6481 34155
rect 5901 34075 6481 34099
rect 5901 34019 5905 34075
rect 5961 34019 5991 34075
rect 6047 34019 6077 34075
rect 6133 34019 6163 34075
rect 6219 34019 6249 34075
rect 6305 34019 6335 34075
rect 6391 34019 6421 34075
rect 6477 34019 6481 34075
rect 5901 33995 6481 34019
rect 5901 33939 5905 33995
rect 5961 33939 5991 33995
rect 6047 33939 6077 33995
rect 6133 33939 6163 33995
rect 6219 33939 6249 33995
rect 6305 33939 6335 33995
rect 6391 33939 6421 33995
rect 6477 33939 6481 33995
rect 5901 33915 6481 33939
rect 5901 33859 5905 33915
rect 5961 33859 5991 33915
rect 6047 33859 6077 33915
rect 6133 33859 6163 33915
rect 6219 33859 6249 33915
rect 6305 33859 6335 33915
rect 6391 33859 6421 33915
rect 6477 33859 6481 33915
rect 5901 33835 6481 33859
rect 5901 33779 5905 33835
rect 5961 33779 5991 33835
rect 6047 33779 6077 33835
rect 6133 33779 6163 33835
rect 6219 33779 6249 33835
rect 6305 33779 6335 33835
rect 6391 33779 6421 33835
rect 6477 33779 6481 33835
rect 5901 33755 6481 33779
rect 5901 33699 5905 33755
rect 5961 33699 5991 33755
rect 6047 33699 6077 33755
rect 6133 33699 6163 33755
rect 6219 33699 6249 33755
rect 6305 33699 6335 33755
rect 6391 33699 6421 33755
rect 6477 33699 6481 33755
rect 5901 33675 6481 33699
rect 5901 33619 5905 33675
rect 5961 33619 5991 33675
rect 6047 33619 6077 33675
rect 6133 33619 6163 33675
rect 6219 33619 6249 33675
rect 6305 33619 6335 33675
rect 6391 33619 6421 33675
rect 6477 33619 6481 33675
rect 5901 33595 6481 33619
rect 5901 33539 5905 33595
rect 5961 33539 5991 33595
rect 6047 33539 6077 33595
rect 6133 33539 6163 33595
rect 6219 33539 6249 33595
rect 6305 33539 6335 33595
rect 6391 33539 6421 33595
rect 6477 33539 6481 33595
rect 5901 33515 6481 33539
rect 5901 33459 5905 33515
rect 5961 33459 5991 33515
rect 6047 33459 6077 33515
rect 6133 33459 6163 33515
rect 6219 33459 6249 33515
rect 6305 33459 6335 33515
rect 6391 33459 6421 33515
rect 6477 33459 6481 33515
rect 5901 33435 6481 33459
rect 5901 33379 5905 33435
rect 5961 33379 5991 33435
rect 6047 33379 6077 33435
rect 6133 33379 6163 33435
rect 6219 33379 6249 33435
rect 6305 33379 6335 33435
rect 6391 33379 6421 33435
rect 6477 33379 6481 33435
rect 5901 33355 6481 33379
rect 5901 33299 5905 33355
rect 5961 33299 5991 33355
rect 6047 33299 6077 33355
rect 6133 33299 6163 33355
rect 6219 33299 6249 33355
rect 6305 33299 6335 33355
rect 6391 33299 6421 33355
rect 6477 33299 6481 33355
rect 5901 33275 6481 33299
rect 5901 33219 5905 33275
rect 5961 33219 5991 33275
rect 6047 33219 6077 33275
rect 6133 33219 6163 33275
rect 6219 33219 6249 33275
rect 6305 33219 6335 33275
rect 6391 33219 6421 33275
rect 6477 33219 6481 33275
rect 5901 33195 6481 33219
rect 5901 33139 5905 33195
rect 5961 33139 5991 33195
rect 6047 33139 6077 33195
rect 6133 33139 6163 33195
rect 6219 33139 6249 33195
rect 6305 33139 6335 33195
rect 6391 33139 6421 33195
rect 6477 33139 6481 33195
rect 5901 33115 6481 33139
rect 5901 33059 5905 33115
rect 5961 33059 5991 33115
rect 6047 33059 6077 33115
rect 6133 33059 6163 33115
rect 6219 33059 6249 33115
rect 6305 33059 6335 33115
rect 6391 33059 6421 33115
rect 6477 33059 6481 33115
rect 5901 33035 6481 33059
rect 5901 32979 5905 33035
rect 5961 32979 5991 33035
rect 6047 32979 6077 33035
rect 6133 32979 6163 33035
rect 6219 32979 6249 33035
rect 6305 32979 6335 33035
rect 6391 32979 6421 33035
rect 6477 32979 6481 33035
rect 5901 32955 6481 32979
rect 5901 32899 5905 32955
rect 5961 32899 5991 32955
rect 6047 32899 6077 32955
rect 6133 32899 6163 32955
rect 6219 32899 6249 32955
rect 6305 32899 6335 32955
rect 6391 32899 6421 32955
rect 6477 32899 6481 32955
rect 5901 32875 6481 32899
rect 5901 32819 5905 32875
rect 5961 32819 5991 32875
rect 6047 32819 6077 32875
rect 6133 32819 6163 32875
rect 6219 32819 6249 32875
rect 6305 32819 6335 32875
rect 6391 32819 6421 32875
rect 6477 32819 6481 32875
rect 5901 32795 6481 32819
rect 5901 32739 5905 32795
rect 5961 32739 5991 32795
rect 6047 32739 6077 32795
rect 6133 32739 6163 32795
rect 6219 32739 6249 32795
rect 6305 32739 6335 32795
rect 6391 32739 6421 32795
rect 6477 32739 6481 32795
rect 5901 32715 6481 32739
rect 5901 32659 5905 32715
rect 5961 32659 5991 32715
rect 6047 32659 6077 32715
rect 6133 32659 6163 32715
rect 6219 32659 6249 32715
rect 6305 32659 6335 32715
rect 6391 32659 6421 32715
rect 6477 32659 6481 32715
rect 5901 32635 6481 32659
rect 5901 32579 5905 32635
rect 5961 32579 5991 32635
rect 6047 32579 6077 32635
rect 6133 32579 6163 32635
rect 6219 32579 6249 32635
rect 6305 32579 6335 32635
rect 6391 32579 6421 32635
rect 6477 32579 6481 32635
rect 5901 32555 6481 32579
rect 5901 32499 5905 32555
rect 5961 32499 5991 32555
rect 6047 32499 6077 32555
rect 6133 32499 6163 32555
rect 6219 32499 6249 32555
rect 6305 32499 6335 32555
rect 6391 32499 6421 32555
rect 6477 32499 6481 32555
rect 5901 32475 6481 32499
rect 5901 32419 5905 32475
rect 5961 32419 5991 32475
rect 6047 32419 6077 32475
rect 6133 32419 6163 32475
rect 6219 32419 6249 32475
rect 6305 32419 6335 32475
rect 6391 32419 6421 32475
rect 6477 32419 6481 32475
rect 5901 32395 6481 32419
rect 5901 32339 5905 32395
rect 5961 32339 5991 32395
rect 6047 32339 6077 32395
rect 6133 32339 6163 32395
rect 6219 32339 6249 32395
rect 6305 32339 6335 32395
rect 6391 32339 6421 32395
rect 6477 32339 6481 32395
rect 5901 32315 6481 32339
rect 5901 32259 5905 32315
rect 5961 32259 5991 32315
rect 6047 32259 6077 32315
rect 6133 32259 6163 32315
rect 6219 32259 6249 32315
rect 6305 32259 6335 32315
rect 6391 32259 6421 32315
rect 6477 32259 6481 32315
rect 5901 32235 6481 32259
rect 5901 32179 5905 32235
rect 5961 32179 5991 32235
rect 6047 32179 6077 32235
rect 6133 32179 6163 32235
rect 6219 32179 6249 32235
rect 6305 32179 6335 32235
rect 6391 32179 6421 32235
rect 6477 32179 6481 32235
rect 5901 32155 6481 32179
rect 5901 32099 5905 32155
rect 5961 32099 5991 32155
rect 6047 32099 6077 32155
rect 6133 32099 6163 32155
rect 6219 32099 6249 32155
rect 6305 32099 6335 32155
rect 6391 32099 6421 32155
rect 6477 32099 6481 32155
rect 5901 32075 6481 32099
rect 5901 32019 5905 32075
rect 5961 32019 5991 32075
rect 6047 32019 6077 32075
rect 6133 32019 6163 32075
rect 6219 32019 6249 32075
rect 6305 32019 6335 32075
rect 6391 32019 6421 32075
rect 6477 32019 6481 32075
rect 5901 31995 6481 32019
rect 5901 31939 5905 31995
rect 5961 31939 5991 31995
rect 6047 31939 6077 31995
rect 6133 31939 6163 31995
rect 6219 31939 6249 31995
rect 6305 31939 6335 31995
rect 6391 31939 6421 31995
rect 6477 31939 6481 31995
rect 5901 31915 6481 31939
rect 5901 31859 5905 31915
rect 5961 31859 5991 31915
rect 6047 31859 6077 31915
rect 6133 31859 6163 31915
rect 6219 31859 6249 31915
rect 6305 31859 6335 31915
rect 6391 31859 6421 31915
rect 6477 31859 6481 31915
rect 5901 31835 6481 31859
rect 5901 31779 5905 31835
rect 5961 31779 5991 31835
rect 6047 31779 6077 31835
rect 6133 31779 6163 31835
rect 6219 31779 6249 31835
rect 6305 31779 6335 31835
rect 6391 31779 6421 31835
rect 6477 31779 6481 31835
rect 5901 31755 6481 31779
rect 5901 31699 5905 31755
rect 5961 31699 5991 31755
rect 6047 31699 6077 31755
rect 6133 31699 6163 31755
rect 6219 31699 6249 31755
rect 6305 31699 6335 31755
rect 6391 31699 6421 31755
rect 6477 31699 6481 31755
rect 5901 31675 6481 31699
rect 5901 31619 5905 31675
rect 5961 31619 5991 31675
rect 6047 31619 6077 31675
rect 6133 31619 6163 31675
rect 6219 31619 6249 31675
rect 6305 31619 6335 31675
rect 6391 31619 6421 31675
rect 6477 31619 6481 31675
rect 5901 31595 6481 31619
rect 5901 31539 5905 31595
rect 5961 31539 5991 31595
rect 6047 31539 6077 31595
rect 6133 31539 6163 31595
rect 6219 31539 6249 31595
rect 6305 31539 6335 31595
rect 6391 31539 6421 31595
rect 6477 31539 6481 31595
rect 5901 31515 6481 31539
rect 5901 31459 5905 31515
rect 5961 31459 5991 31515
rect 6047 31459 6077 31515
rect 6133 31459 6163 31515
rect 6219 31459 6249 31515
rect 6305 31459 6335 31515
rect 6391 31459 6421 31515
rect 6477 31459 6481 31515
rect 5901 31435 6481 31459
rect 5901 31379 5905 31435
rect 5961 31379 5991 31435
rect 6047 31379 6077 31435
rect 6133 31379 6163 31435
rect 6219 31379 6249 31435
rect 6305 31379 6335 31435
rect 6391 31379 6421 31435
rect 6477 31379 6481 31435
rect 5901 31355 6481 31379
rect 5901 31299 5905 31355
rect 5961 31299 5991 31355
rect 6047 31299 6077 31355
rect 6133 31299 6163 31355
rect 6219 31299 6249 31355
rect 6305 31299 6335 31355
rect 6391 31299 6421 31355
rect 6477 31299 6481 31355
rect 5901 31275 6481 31299
rect 5901 31219 5905 31275
rect 5961 31219 5991 31275
rect 6047 31219 6077 31275
rect 6133 31219 6163 31275
rect 6219 31219 6249 31275
rect 6305 31219 6335 31275
rect 6391 31219 6421 31275
rect 6477 31219 6481 31275
rect 5901 31195 6481 31219
rect 5901 31139 5905 31195
rect 5961 31139 5991 31195
rect 6047 31139 6077 31195
rect 6133 31139 6163 31195
rect 6219 31139 6249 31195
rect 6305 31139 6335 31195
rect 6391 31139 6421 31195
rect 6477 31139 6481 31195
rect 5901 31115 6481 31139
rect 5901 31059 5905 31115
rect 5961 31059 5991 31115
rect 6047 31059 6077 31115
rect 6133 31059 6163 31115
rect 6219 31059 6249 31115
rect 6305 31059 6335 31115
rect 6391 31059 6421 31115
rect 6477 31059 6481 31115
rect 5901 31035 6481 31059
rect 5901 30979 5905 31035
rect 5961 30979 5991 31035
rect 6047 30979 6077 31035
rect 6133 30979 6163 31035
rect 6219 30979 6249 31035
rect 6305 30979 6335 31035
rect 6391 30979 6421 31035
rect 6477 30979 6481 31035
rect 5901 30955 6481 30979
rect 5901 30899 5905 30955
rect 5961 30899 5991 30955
rect 6047 30899 6077 30955
rect 6133 30899 6163 30955
rect 6219 30899 6249 30955
rect 6305 30899 6335 30955
rect 6391 30899 6421 30955
rect 6477 30899 6481 30955
rect 5901 30875 6481 30899
rect 5901 30819 5905 30875
rect 5961 30819 5991 30875
rect 6047 30819 6077 30875
rect 6133 30819 6163 30875
rect 6219 30819 6249 30875
rect 6305 30819 6335 30875
rect 6391 30819 6421 30875
rect 6477 30819 6481 30875
rect 5901 30795 6481 30819
rect 5901 30739 5905 30795
rect 5961 30739 5991 30795
rect 6047 30739 6077 30795
rect 6133 30739 6163 30795
rect 6219 30739 6249 30795
rect 6305 30739 6335 30795
rect 6391 30739 6421 30795
rect 6477 30739 6481 30795
rect 5901 30715 6481 30739
rect 5901 30659 5905 30715
rect 5961 30659 5991 30715
rect 6047 30659 6077 30715
rect 6133 30659 6163 30715
rect 6219 30659 6249 30715
rect 6305 30659 6335 30715
rect 6391 30659 6421 30715
rect 6477 30659 6481 30715
rect 5901 30635 6481 30659
rect 5901 30579 5905 30635
rect 5961 30579 5991 30635
rect 6047 30579 6077 30635
rect 6133 30579 6163 30635
rect 6219 30579 6249 30635
rect 6305 30579 6335 30635
rect 6391 30579 6421 30635
rect 6477 30579 6481 30635
rect 5901 30555 6481 30579
rect 5901 30499 5905 30555
rect 5961 30499 5991 30555
rect 6047 30499 6077 30555
rect 6133 30499 6163 30555
rect 6219 30499 6249 30555
rect 6305 30499 6335 30555
rect 6391 30499 6421 30555
rect 6477 30499 6481 30555
rect 5901 30475 6481 30499
rect 5901 30419 5905 30475
rect 5961 30419 5991 30475
rect 6047 30419 6077 30475
rect 6133 30419 6163 30475
rect 6219 30419 6249 30475
rect 6305 30419 6335 30475
rect 6391 30419 6421 30475
rect 6477 30419 6481 30475
tri 4887 29451 4909 29473 se
rect 4909 29451 4973 29473
tri 4081 29235 4113 29267 se
rect 4113 29235 4167 29267
rect 4039 29183 4045 29235
rect 4097 29183 4109 29235
rect 4161 29183 4167 29235
rect 4221 29399 4973 29451
tri 4219 29183 4221 29185 se
rect 4221 29183 4273 29399
tri 4273 29365 4307 29399 nw
tri 4993 29365 5005 29377 se
rect 5005 29365 5057 30400
rect 5901 30395 6481 30419
rect 5901 30339 5905 30395
rect 5961 30339 5991 30395
rect 6047 30339 6077 30395
rect 6133 30339 6163 30395
rect 6219 30339 6249 30395
rect 6305 30339 6335 30395
rect 6391 30339 6421 30395
rect 6477 30339 6481 30395
rect 5901 30315 6481 30339
rect 5901 30259 5905 30315
rect 5961 30259 5991 30315
rect 6047 30259 6077 30315
rect 6133 30259 6163 30315
rect 6219 30259 6249 30315
rect 6305 30259 6335 30315
rect 6391 30259 6421 30315
rect 6477 30259 6481 30315
rect 5901 30235 6481 30259
rect 5901 30179 5905 30235
rect 5961 30179 5991 30235
rect 6047 30179 6077 30235
rect 6133 30179 6163 30235
rect 6219 30179 6249 30235
rect 6305 30179 6335 30235
rect 6391 30179 6421 30235
rect 6477 30179 6481 30235
rect 5901 30155 6481 30179
rect 5901 30099 5905 30155
rect 5961 30099 5991 30155
rect 6047 30099 6077 30155
rect 6133 30099 6163 30155
rect 6219 30099 6249 30155
rect 6305 30099 6335 30155
rect 6391 30099 6421 30155
rect 6477 30099 6481 30155
rect 5901 30075 6481 30099
rect 5901 30019 5905 30075
rect 5961 30019 5991 30075
rect 6047 30019 6077 30075
rect 6133 30019 6163 30075
rect 6219 30019 6249 30075
rect 6305 30019 6335 30075
rect 6391 30019 6421 30075
rect 6477 30019 6481 30075
rect 6900 34774 6903 34830
rect 6959 34774 6993 34830
rect 7049 34774 7083 34830
rect 7139 34774 7173 34830
rect 7229 34774 7263 34830
rect 7319 34774 7353 34830
rect 7409 34774 7443 34830
rect 7499 34774 7502 34830
rect 6900 34750 7502 34774
rect 6900 34694 6903 34750
rect 6959 34694 6993 34750
rect 7049 34694 7083 34750
rect 7139 34694 7173 34750
rect 7229 34694 7263 34750
rect 7319 34694 7353 34750
rect 7409 34694 7443 34750
rect 7499 34694 7502 34750
rect 6900 34670 7502 34694
rect 6900 34614 6903 34670
rect 6959 34614 6993 34670
rect 7049 34614 7083 34670
rect 7139 34614 7173 34670
rect 7229 34614 7263 34670
rect 7319 34614 7353 34670
rect 7409 34614 7443 34670
rect 7499 34614 7502 34670
rect 6900 34590 7502 34614
rect 6900 34534 6903 34590
rect 6959 34534 6993 34590
rect 7049 34534 7083 34590
rect 7139 34534 7173 34590
rect 7229 34534 7263 34590
rect 7319 34534 7353 34590
rect 7409 34534 7443 34590
rect 7499 34534 7502 34590
rect 6900 34510 7502 34534
rect 6900 34454 6903 34510
rect 6959 34454 6993 34510
rect 7049 34454 7083 34510
rect 7139 34454 7173 34510
rect 7229 34454 7263 34510
rect 7319 34454 7353 34510
rect 7409 34454 7443 34510
rect 7499 34454 7502 34510
rect 6900 34430 7502 34454
rect 6900 34374 6903 34430
rect 6959 34374 6993 34430
rect 7049 34374 7083 34430
rect 7139 34374 7173 34430
rect 7229 34374 7263 34430
rect 7319 34374 7353 34430
rect 7409 34374 7443 34430
rect 7499 34374 7502 34430
rect 6900 34350 7502 34374
rect 6900 34294 6903 34350
rect 6959 34294 6993 34350
rect 7049 34294 7083 34350
rect 7139 34294 7173 34350
rect 7229 34294 7263 34350
rect 7319 34294 7353 34350
rect 7409 34294 7443 34350
rect 7499 34294 7502 34350
rect 6900 34270 7502 34294
rect 6900 34214 6903 34270
rect 6959 34214 6993 34270
rect 7049 34214 7083 34270
rect 7139 34214 7173 34270
rect 7229 34214 7263 34270
rect 7319 34214 7353 34270
rect 7409 34214 7443 34270
rect 7499 34214 7502 34270
rect 6900 34190 7502 34214
rect 6900 34134 6903 34190
rect 6959 34134 6993 34190
rect 7049 34134 7083 34190
rect 7139 34134 7173 34190
rect 7229 34134 7263 34190
rect 7319 34134 7353 34190
rect 7409 34134 7443 34190
rect 7499 34134 7502 34190
rect 6900 34110 7502 34134
rect 6900 34054 6903 34110
rect 6959 34054 6993 34110
rect 7049 34054 7083 34110
rect 7139 34054 7173 34110
rect 7229 34054 7263 34110
rect 7319 34054 7353 34110
rect 7409 34054 7443 34110
rect 7499 34054 7502 34110
rect 6900 34030 7502 34054
rect 6900 33974 6903 34030
rect 6959 33974 6993 34030
rect 7049 33974 7083 34030
rect 7139 33974 7173 34030
rect 7229 33974 7263 34030
rect 7319 33974 7353 34030
rect 7409 33974 7443 34030
rect 7499 33974 7502 34030
rect 6900 33950 7502 33974
rect 6900 33894 6903 33950
rect 6959 33894 6993 33950
rect 7049 33894 7083 33950
rect 7139 33894 7173 33950
rect 7229 33894 7263 33950
rect 7319 33894 7353 33950
rect 7409 33894 7443 33950
rect 7499 33894 7502 33950
rect 6900 33870 7502 33894
rect 6900 33814 6903 33870
rect 6959 33814 6993 33870
rect 7049 33814 7083 33870
rect 7139 33814 7173 33870
rect 7229 33814 7263 33870
rect 7319 33814 7353 33870
rect 7409 33814 7443 33870
rect 7499 33814 7502 33870
rect 6900 33790 7502 33814
rect 6900 33734 6903 33790
rect 6959 33734 6993 33790
rect 7049 33734 7083 33790
rect 7139 33734 7173 33790
rect 7229 33734 7263 33790
rect 7319 33734 7353 33790
rect 7409 33734 7443 33790
rect 7499 33734 7502 33790
rect 6900 33710 7502 33734
rect 6900 33654 6903 33710
rect 6959 33654 6993 33710
rect 7049 33654 7083 33710
rect 7139 33654 7173 33710
rect 7229 33654 7263 33710
rect 7319 33654 7353 33710
rect 7409 33654 7443 33710
rect 7499 33654 7502 33710
rect 6900 33630 7502 33654
rect 6900 33574 6903 33630
rect 6959 33574 6993 33630
rect 7049 33574 7083 33630
rect 7139 33574 7173 33630
rect 7229 33574 7263 33630
rect 7319 33574 7353 33630
rect 7409 33574 7443 33630
rect 7499 33574 7502 33630
rect 6900 33550 7502 33574
rect 6900 33494 6903 33550
rect 6959 33494 6993 33550
rect 7049 33494 7083 33550
rect 7139 33494 7173 33550
rect 7229 33494 7263 33550
rect 7319 33494 7353 33550
rect 7409 33494 7443 33550
rect 7499 33494 7502 33550
rect 6900 33470 7502 33494
rect 6900 33414 6903 33470
rect 6959 33414 6993 33470
rect 7049 33414 7083 33470
rect 7139 33414 7173 33470
rect 7229 33414 7263 33470
rect 7319 33414 7353 33470
rect 7409 33414 7443 33470
rect 7499 33414 7502 33470
rect 6900 33390 7502 33414
rect 6900 33334 6903 33390
rect 6959 33334 6993 33390
rect 7049 33334 7083 33390
rect 7139 33334 7173 33390
rect 7229 33334 7263 33390
rect 7319 33334 7353 33390
rect 7409 33334 7443 33390
rect 7499 33334 7502 33390
rect 6900 33310 7502 33334
rect 6900 33254 6903 33310
rect 6959 33254 6993 33310
rect 7049 33254 7083 33310
rect 7139 33254 7173 33310
rect 7229 33254 7263 33310
rect 7319 33254 7353 33310
rect 7409 33254 7443 33310
rect 7499 33254 7502 33310
rect 6900 33230 7502 33254
rect 6900 33174 6903 33230
rect 6959 33174 6993 33230
rect 7049 33174 7083 33230
rect 7139 33174 7173 33230
rect 7229 33174 7263 33230
rect 7319 33174 7353 33230
rect 7409 33174 7443 33230
rect 7499 33174 7502 33230
rect 6900 33150 7502 33174
rect 6900 33094 6903 33150
rect 6959 33094 6993 33150
rect 7049 33094 7083 33150
rect 7139 33094 7173 33150
rect 7229 33094 7263 33150
rect 7319 33094 7353 33150
rect 7409 33094 7443 33150
rect 7499 33094 7502 33150
rect 6900 33070 7502 33094
rect 6900 33014 6903 33070
rect 6959 33014 6993 33070
rect 7049 33014 7083 33070
rect 7139 33014 7173 33070
rect 7229 33014 7263 33070
rect 7319 33014 7353 33070
rect 7409 33014 7443 33070
rect 7499 33014 7502 33070
rect 6900 32990 7502 33014
rect 6900 32934 6903 32990
rect 6959 32934 6993 32990
rect 7049 32934 7083 32990
rect 7139 32934 7173 32990
rect 7229 32934 7263 32990
rect 7319 32934 7353 32990
rect 7409 32934 7443 32990
rect 7499 32934 7502 32990
rect 6900 32910 7502 32934
rect 6900 32854 6903 32910
rect 6959 32854 6993 32910
rect 7049 32854 7083 32910
rect 7139 32854 7173 32910
rect 7229 32854 7263 32910
rect 7319 32854 7353 32910
rect 7409 32854 7443 32910
rect 7499 32854 7502 32910
rect 6900 32830 7502 32854
rect 6900 32774 6903 32830
rect 6959 32774 6993 32830
rect 7049 32774 7083 32830
rect 7139 32774 7173 32830
rect 7229 32774 7263 32830
rect 7319 32774 7353 32830
rect 7409 32774 7443 32830
rect 7499 32774 7502 32830
rect 6900 32750 7502 32774
rect 6900 32694 6903 32750
rect 6959 32694 6993 32750
rect 7049 32694 7083 32750
rect 7139 32694 7173 32750
rect 7229 32694 7263 32750
rect 7319 32694 7353 32750
rect 7409 32694 7443 32750
rect 7499 32694 7502 32750
rect 6900 32670 7502 32694
rect 6900 32614 6903 32670
rect 6959 32614 6993 32670
rect 7049 32614 7083 32670
rect 7139 32614 7173 32670
rect 7229 32614 7263 32670
rect 7319 32614 7353 32670
rect 7409 32614 7443 32670
rect 7499 32614 7502 32670
rect 6900 32590 7502 32614
rect 6900 32534 6903 32590
rect 6959 32534 6993 32590
rect 7049 32534 7083 32590
rect 7139 32534 7173 32590
rect 7229 32534 7263 32590
rect 7319 32534 7353 32590
rect 7409 32534 7443 32590
rect 7499 32534 7502 32590
rect 6900 32510 7502 32534
rect 6900 32454 6903 32510
rect 6959 32454 6993 32510
rect 7049 32454 7083 32510
rect 7139 32454 7173 32510
rect 7229 32454 7263 32510
rect 7319 32454 7353 32510
rect 7409 32454 7443 32510
rect 7499 32454 7502 32510
rect 6900 32430 7502 32454
rect 6900 32374 6903 32430
rect 6959 32374 6993 32430
rect 7049 32374 7083 32430
rect 7139 32374 7173 32430
rect 7229 32374 7263 32430
rect 7319 32374 7353 32430
rect 7409 32374 7443 32430
rect 7499 32374 7502 32430
rect 6900 32350 7502 32374
rect 6900 32294 6903 32350
rect 6959 32294 6993 32350
rect 7049 32294 7083 32350
rect 7139 32294 7173 32350
rect 7229 32294 7263 32350
rect 7319 32294 7353 32350
rect 7409 32294 7443 32350
rect 7499 32294 7502 32350
rect 6900 32270 7502 32294
rect 6900 32214 6903 32270
rect 6959 32214 6993 32270
rect 7049 32214 7083 32270
rect 7139 32214 7173 32270
rect 7229 32214 7263 32270
rect 7319 32214 7353 32270
rect 7409 32214 7443 32270
rect 7499 32214 7502 32270
rect 6900 32190 7502 32214
rect 6900 32134 6903 32190
rect 6959 32134 6993 32190
rect 7049 32134 7083 32190
rect 7139 32134 7173 32190
rect 7229 32134 7263 32190
rect 7319 32134 7353 32190
rect 7409 32134 7443 32190
rect 7499 32134 7502 32190
rect 6900 32110 7502 32134
rect 6900 32054 6903 32110
rect 6959 32054 6993 32110
rect 7049 32054 7083 32110
rect 7139 32054 7173 32110
rect 7229 32054 7263 32110
rect 7319 32054 7353 32110
rect 7409 32054 7443 32110
rect 7499 32054 7502 32110
rect 6900 32030 7502 32054
rect 6900 31974 6903 32030
rect 6959 31974 6993 32030
rect 7049 31974 7083 32030
rect 7139 31974 7173 32030
rect 7229 31974 7263 32030
rect 7319 31974 7353 32030
rect 7409 31974 7443 32030
rect 7499 31974 7502 32030
rect 6900 31950 7502 31974
rect 6900 31894 6903 31950
rect 6959 31894 6993 31950
rect 7049 31894 7083 31950
rect 7139 31894 7173 31950
rect 7229 31894 7263 31950
rect 7319 31894 7353 31950
rect 7409 31894 7443 31950
rect 7499 31894 7502 31950
rect 6900 31870 7502 31894
rect 6900 31814 6903 31870
rect 6959 31814 6993 31870
rect 7049 31814 7083 31870
rect 7139 31814 7173 31870
rect 7229 31814 7263 31870
rect 7319 31814 7353 31870
rect 7409 31814 7443 31870
rect 7499 31814 7502 31870
rect 6900 31790 7502 31814
rect 6900 31734 6903 31790
rect 6959 31734 6993 31790
rect 7049 31734 7083 31790
rect 7139 31734 7173 31790
rect 7229 31734 7263 31790
rect 7319 31734 7353 31790
rect 7409 31734 7443 31790
rect 7499 31734 7502 31790
rect 6900 31710 7502 31734
rect 6900 31654 6903 31710
rect 6959 31654 6993 31710
rect 7049 31654 7083 31710
rect 7139 31654 7173 31710
rect 7229 31654 7263 31710
rect 7319 31654 7353 31710
rect 7409 31654 7443 31710
rect 7499 31654 7502 31710
rect 6900 31630 7502 31654
rect 6900 31574 6903 31630
rect 6959 31574 6993 31630
rect 7049 31574 7083 31630
rect 7139 31574 7173 31630
rect 7229 31574 7263 31630
rect 7319 31574 7353 31630
rect 7409 31574 7443 31630
rect 7499 31574 7502 31630
rect 6900 31550 7502 31574
rect 6900 31494 6903 31550
rect 6959 31494 6993 31550
rect 7049 31494 7083 31550
rect 7139 31494 7173 31550
rect 7229 31494 7263 31550
rect 7319 31494 7353 31550
rect 7409 31494 7443 31550
rect 7499 31494 7502 31550
rect 6900 31470 7502 31494
rect 6900 31414 6903 31470
rect 6959 31414 6993 31470
rect 7049 31414 7083 31470
rect 7139 31414 7173 31470
rect 7229 31414 7263 31470
rect 7319 31414 7353 31470
rect 7409 31414 7443 31470
rect 7499 31414 7502 31470
rect 6900 31390 7502 31414
rect 6900 31334 6903 31390
rect 6959 31334 6993 31390
rect 7049 31334 7083 31390
rect 7139 31334 7173 31390
rect 7229 31334 7263 31390
rect 7319 31334 7353 31390
rect 7409 31334 7443 31390
rect 7499 31334 7502 31390
rect 6900 31310 7502 31334
rect 6900 31254 6903 31310
rect 6959 31254 6993 31310
rect 7049 31254 7083 31310
rect 7139 31254 7173 31310
rect 7229 31254 7263 31310
rect 7319 31254 7353 31310
rect 7409 31254 7443 31310
rect 7499 31254 7502 31310
rect 6900 31230 7502 31254
rect 6900 31174 6903 31230
rect 6959 31174 6993 31230
rect 7049 31174 7083 31230
rect 7139 31174 7173 31230
rect 7229 31174 7263 31230
rect 7319 31174 7353 31230
rect 7409 31174 7443 31230
rect 7499 31174 7502 31230
rect 6900 31150 7502 31174
rect 6900 31094 6903 31150
rect 6959 31094 6993 31150
rect 7049 31094 7083 31150
rect 7139 31094 7173 31150
rect 7229 31094 7263 31150
rect 7319 31094 7353 31150
rect 7409 31094 7443 31150
rect 7499 31094 7502 31150
rect 6900 31070 7502 31094
rect 6900 31014 6903 31070
rect 6959 31014 6993 31070
rect 7049 31014 7083 31070
rect 7139 31014 7173 31070
rect 7229 31014 7263 31070
rect 7319 31014 7353 31070
rect 7409 31014 7443 31070
rect 7499 31014 7502 31070
rect 6900 30990 7502 31014
rect 6900 30934 6903 30990
rect 6959 30934 6993 30990
rect 7049 30934 7083 30990
rect 7139 30934 7173 30990
rect 7229 30934 7263 30990
rect 7319 30934 7353 30990
rect 7409 30934 7443 30990
rect 7499 30934 7502 30990
rect 6900 30910 7502 30934
rect 6900 30854 6903 30910
rect 6959 30854 6993 30910
rect 7049 30854 7083 30910
rect 7139 30854 7173 30910
rect 7229 30854 7263 30910
rect 7319 30854 7353 30910
rect 7409 30854 7443 30910
rect 7499 30854 7502 30910
rect 6900 30830 7502 30854
rect 6900 30774 6903 30830
rect 6959 30774 6993 30830
rect 7049 30774 7083 30830
rect 7139 30774 7173 30830
rect 7229 30774 7263 30830
rect 7319 30774 7353 30830
rect 7409 30774 7443 30830
rect 7499 30774 7502 30830
rect 6900 30750 7502 30774
rect 6900 30694 6903 30750
rect 6959 30694 6993 30750
rect 7049 30694 7083 30750
rect 7139 30694 7173 30750
rect 7229 30694 7263 30750
rect 7319 30694 7353 30750
rect 7409 30694 7443 30750
rect 7499 30694 7502 30750
rect 6900 30670 7502 30694
rect 6900 30614 6903 30670
rect 6959 30614 6993 30670
rect 7049 30614 7083 30670
rect 7139 30614 7173 30670
rect 7229 30614 7263 30670
rect 7319 30614 7353 30670
rect 7409 30614 7443 30670
rect 7499 30614 7502 30670
rect 6900 30590 7502 30614
rect 6900 30534 6903 30590
rect 6959 30534 6993 30590
rect 7049 30534 7083 30590
rect 7139 30534 7173 30590
rect 7229 30534 7263 30590
rect 7319 30534 7353 30590
rect 7409 30534 7443 30590
rect 7499 30534 7502 30590
rect 6900 30510 7502 30534
rect 6900 30454 6903 30510
rect 6959 30454 6993 30510
rect 7049 30454 7083 30510
rect 7139 30454 7173 30510
rect 7229 30454 7263 30510
rect 7319 30454 7353 30510
rect 7409 30454 7443 30510
rect 7499 30454 7502 30510
rect 6900 30430 7502 30454
rect 6900 30374 6903 30430
rect 6959 30374 6993 30430
rect 7049 30374 7083 30430
rect 7139 30374 7173 30430
rect 7229 30374 7263 30430
rect 7319 30374 7353 30430
rect 7409 30374 7443 30430
rect 7499 30374 7502 30430
rect 6900 30350 7502 30374
rect 6900 30294 6903 30350
rect 6959 30294 6993 30350
rect 7049 30294 7083 30350
rect 7139 30294 7173 30350
rect 7229 30294 7263 30350
rect 7319 30294 7353 30350
rect 7409 30294 7443 30350
rect 7499 30294 7502 30350
rect 6900 30270 7502 30294
rect 6900 30214 6903 30270
rect 6959 30214 6993 30270
rect 7049 30214 7083 30270
rect 7139 30214 7173 30270
rect 7229 30214 7263 30270
rect 7319 30214 7353 30270
rect 7409 30214 7443 30270
rect 7499 30214 7502 30270
rect 6900 30189 7502 30214
rect 6900 30133 6903 30189
rect 6959 30133 6993 30189
rect 7049 30133 7083 30189
rect 7139 30133 7173 30189
rect 7229 30133 7263 30189
rect 7319 30133 7353 30189
rect 7409 30133 7443 30189
rect 7499 30133 7502 30189
rect 6900 30108 7502 30133
rect 6900 30052 6903 30108
rect 6959 30052 6993 30108
rect 7049 30052 7083 30108
rect 7139 30052 7173 30108
rect 7229 30052 7263 30108
rect 7319 30052 7353 30108
rect 7409 30052 7443 30108
rect 7499 30052 7502 30108
rect 6900 30043 7502 30052
rect 5901 30010 6481 30019
tri 4979 29351 4993 29365 se
rect 4993 29351 5057 29365
tri 4971 29343 4979 29351 se
rect 4979 29343 5057 29351
tri 4187 29151 4219 29183 se
rect 4219 29151 4273 29183
rect 4145 29099 4151 29151
rect 4203 29099 4215 29151
rect 4267 29099 4273 29151
rect 4320 29291 5057 29343
rect 5220 29351 5226 29403
rect 5278 29351 5290 29403
rect 5342 29351 5348 29403
rect 5220 29319 5274 29351
tri 5274 29319 5306 29351 nw
rect 4320 29267 4382 29291
tri 4382 29267 4406 29291 nw
tri 4318 29099 4320 29101 se
rect 4320 29099 4372 29267
tri 4372 29257 4382 29267 nw
tri 5210 29151 5220 29161 se
rect 5220 29151 5272 29319
tri 5272 29317 5274 29319 nw
tri 5186 29127 5210 29151 se
rect 5210 29127 5272 29151
tri 4286 29067 4318 29099 se
rect 4318 29067 4372 29099
rect 4244 29015 4250 29067
rect 4302 29015 4314 29067
rect 4366 29015 4372 29067
rect 4535 29075 5272 29127
rect 5319 29267 5325 29319
rect 5377 29267 5389 29319
rect 5441 29267 5447 29319
rect 5319 29235 5373 29267
tri 5373 29235 5405 29267 nw
rect 4535 29067 4613 29075
tri 4613 29067 4621 29075 nw
rect 4535 28018 4587 29067
tri 4587 29041 4613 29067 nw
tri 5307 29041 5319 29053 se
rect 5319 29041 5371 29235
tri 5371 29233 5373 29235 nw
tri 5285 29019 5307 29041 se
rect 5307 29019 5371 29041
rect 4627 28967 5371 29019
rect 5425 29183 5431 29235
rect 5483 29183 5495 29235
rect 5547 29183 5553 29235
rect 5425 29151 5479 29183
tri 5479 29151 5511 29183 nw
rect 2911 24037 3491 24046
rect 2911 23981 2915 24037
rect 2971 23981 3001 24037
rect 3057 23981 3087 24037
rect 3143 23981 3173 24037
rect 3229 23981 3259 24037
rect 3315 23981 3345 24037
rect 3401 23981 3431 24037
rect 3487 23981 3491 24037
rect 2911 23957 3491 23981
rect 2911 23901 2915 23957
rect 2971 23901 3001 23957
rect 3057 23901 3087 23957
rect 3143 23901 3173 23957
rect 3229 23901 3259 23957
rect 3315 23901 3345 23957
rect 3401 23901 3431 23957
rect 3487 23901 3491 23957
rect 2911 23877 3491 23901
rect 2911 23821 2915 23877
rect 2971 23821 3001 23877
rect 3057 23821 3087 23877
rect 3143 23821 3173 23877
rect 3229 23821 3259 23877
rect 3315 23821 3345 23877
rect 3401 23821 3431 23877
rect 3487 23821 3491 23877
rect 2911 23797 3491 23821
rect 2911 23741 2915 23797
rect 2971 23741 3001 23797
rect 3057 23741 3087 23797
rect 3143 23741 3173 23797
rect 3229 23741 3259 23797
rect 3315 23741 3345 23797
rect 3401 23741 3431 23797
rect 3487 23741 3491 23797
rect 2911 23717 3491 23741
rect 2911 23661 2915 23717
rect 2971 23661 3001 23717
rect 3057 23661 3087 23717
rect 3143 23661 3173 23717
rect 3229 23661 3259 23717
rect 3315 23661 3345 23717
rect 3401 23661 3431 23717
rect 3487 23661 3491 23717
rect 2911 23637 3491 23661
rect 2911 23581 2915 23637
rect 2971 23581 3001 23637
rect 3057 23581 3087 23637
rect 3143 23581 3173 23637
rect 3229 23581 3259 23637
rect 3315 23581 3345 23637
rect 3401 23581 3431 23637
rect 3487 23581 3491 23637
rect 2911 23557 3491 23581
rect 2911 23501 2915 23557
rect 2971 23501 3001 23557
rect 3057 23501 3087 23557
rect 3143 23501 3173 23557
rect 3229 23501 3259 23557
rect 3315 23501 3345 23557
rect 3401 23501 3431 23557
rect 3487 23501 3491 23557
rect 2911 23477 3491 23501
rect 2911 23421 2915 23477
rect 2971 23421 3001 23477
rect 3057 23421 3087 23477
rect 3143 23421 3173 23477
rect 3229 23421 3259 23477
rect 3315 23421 3345 23477
rect 3401 23421 3431 23477
rect 3487 23421 3491 23477
rect 2911 23397 3491 23421
rect 2911 23341 2915 23397
rect 2971 23341 3001 23397
rect 3057 23341 3087 23397
rect 3143 23341 3173 23397
rect 3229 23341 3259 23397
rect 3315 23341 3345 23397
rect 3401 23341 3431 23397
rect 3487 23341 3491 23397
rect 2911 23317 3491 23341
rect 2911 23261 2915 23317
rect 2971 23261 3001 23317
rect 3057 23261 3087 23317
rect 3143 23261 3173 23317
rect 3229 23261 3259 23317
rect 3315 23261 3345 23317
rect 3401 23261 3431 23317
rect 3487 23261 3491 23317
rect 2911 23237 3491 23261
rect 2911 23181 2915 23237
rect 2971 23181 3001 23237
rect 3057 23181 3087 23237
rect 3143 23181 3173 23237
rect 3229 23181 3259 23237
rect 3315 23181 3345 23237
rect 3401 23181 3431 23237
rect 3487 23181 3491 23237
rect 2911 23157 3491 23181
rect 2911 23101 2915 23157
rect 2971 23101 3001 23157
rect 3057 23101 3087 23157
rect 3143 23101 3173 23157
rect 3229 23101 3259 23157
rect 3315 23101 3345 23157
rect 3401 23101 3431 23157
rect 3487 23101 3491 23157
rect 2911 23077 3491 23101
rect 2911 23021 2915 23077
rect 2971 23021 3001 23077
rect 3057 23021 3087 23077
rect 3143 23021 3173 23077
rect 3229 23021 3259 23077
rect 3315 23021 3345 23077
rect 3401 23021 3431 23077
rect 3487 23021 3491 23077
rect 2911 22997 3491 23021
rect 2911 22941 2915 22997
rect 2971 22941 3001 22997
rect 3057 22941 3087 22997
rect 3143 22941 3173 22997
rect 3229 22941 3259 22997
rect 3315 22941 3345 22997
rect 3401 22941 3431 22997
rect 3487 22941 3491 22997
rect 2911 22917 3491 22941
rect 2911 22861 2915 22917
rect 2971 22861 3001 22917
rect 3057 22861 3087 22917
rect 3143 22861 3173 22917
rect 3229 22861 3259 22917
rect 3315 22861 3345 22917
rect 3401 22861 3431 22917
rect 3487 22861 3491 22917
rect 2911 22837 3491 22861
rect 2911 22781 2915 22837
rect 2971 22781 3001 22837
rect 3057 22781 3087 22837
rect 3143 22781 3173 22837
rect 3229 22781 3259 22837
rect 3315 22781 3345 22837
rect 3401 22781 3431 22837
rect 3487 22781 3491 22837
rect 2911 22757 3491 22781
rect 2911 22701 2915 22757
rect 2971 22701 3001 22757
rect 3057 22701 3087 22757
rect 3143 22701 3173 22757
rect 3229 22701 3259 22757
rect 3315 22701 3345 22757
rect 3401 22701 3431 22757
rect 3487 22701 3491 22757
rect 2911 22677 3491 22701
rect 2911 22621 2915 22677
rect 2971 22621 3001 22677
rect 3057 22621 3087 22677
rect 3143 22621 3173 22677
rect 3229 22621 3259 22677
rect 3315 22621 3345 22677
rect 3401 22621 3431 22677
rect 3487 22621 3491 22677
rect 2911 22597 3491 22621
rect 2911 22541 2915 22597
rect 2971 22541 3001 22597
rect 3057 22541 3087 22597
rect 3143 22541 3173 22597
rect 3229 22541 3259 22597
rect 3315 22541 3345 22597
rect 3401 22541 3431 22597
rect 3487 22541 3491 22597
rect 4627 22783 4679 28967
tri 4679 28933 4713 28967 nw
tri 5413 28933 5425 28945 se
rect 5425 28933 5477 29151
tri 5477 29149 5479 29151 nw
tri 5391 28911 5413 28933 se
rect 5413 28911 5477 28933
rect 4627 22693 4679 22731
rect 4627 22603 4679 22641
rect 4627 22545 4679 22551
rect 4711 28859 5477 28911
rect 5532 29099 5538 29151
rect 5590 29099 5602 29151
rect 5654 29099 5660 29151
rect 5532 29067 5586 29099
tri 5586 29067 5618 29099 nw
rect 2911 22517 3491 22541
rect 2911 22461 2915 22517
rect 2971 22461 3001 22517
rect 3057 22461 3087 22517
rect 3143 22461 3173 22517
rect 3229 22461 3259 22517
rect 3315 22461 3345 22517
rect 3401 22461 3431 22517
rect 3487 22461 3491 22517
rect 2911 22437 3491 22461
rect 2911 22381 2915 22437
rect 2971 22381 3001 22437
rect 3057 22381 3087 22437
rect 3143 22381 3173 22437
rect 3229 22381 3259 22437
rect 3315 22381 3345 22437
rect 3401 22381 3431 22437
rect 3487 22381 3491 22437
rect 2911 22357 3491 22381
rect 2911 22301 2915 22357
rect 2971 22301 3001 22357
rect 3057 22301 3087 22357
rect 3143 22301 3173 22357
rect 3229 22301 3259 22357
rect 3315 22301 3345 22357
rect 3401 22301 3431 22357
rect 3487 22301 3491 22357
rect 2911 22277 3491 22301
rect 2911 22221 2915 22277
rect 2971 22221 3001 22277
rect 3057 22221 3087 22277
rect 3143 22221 3173 22277
rect 3229 22221 3259 22277
rect 3315 22221 3345 22277
rect 3401 22221 3431 22277
rect 3487 22221 3491 22277
rect 2911 22197 3491 22221
rect 2911 22141 2915 22197
rect 2971 22141 3001 22197
rect 3057 22141 3087 22197
rect 3143 22141 3173 22197
rect 3229 22141 3259 22197
rect 3315 22141 3345 22197
rect 3401 22141 3431 22197
rect 3487 22141 3491 22197
rect 2911 22117 3491 22141
rect 2911 22061 2915 22117
rect 2971 22061 3001 22117
rect 3057 22061 3087 22117
rect 3143 22061 3173 22117
rect 3229 22061 3259 22117
rect 3315 22061 3345 22117
rect 3401 22061 3431 22117
rect 3487 22061 3491 22117
rect 2911 22037 3491 22061
rect 2911 21981 2915 22037
rect 2971 21981 3001 22037
rect 3057 21981 3087 22037
rect 3143 21981 3173 22037
rect 3229 21981 3259 22037
rect 3315 21981 3345 22037
rect 3401 21981 3431 22037
rect 3487 21981 3491 22037
rect 2911 21957 3491 21981
rect 2911 21901 2915 21957
rect 2971 21901 3001 21957
rect 3057 21901 3087 21957
rect 3143 21901 3173 21957
rect 3229 21901 3259 21957
rect 3315 21901 3345 21957
rect 3401 21901 3431 21957
rect 3487 21901 3491 21957
rect 2911 21877 3491 21901
rect 2911 21821 2915 21877
rect 2971 21821 3001 21877
rect 3057 21821 3087 21877
rect 3143 21821 3173 21877
rect 3229 21821 3259 21877
rect 3315 21821 3345 21877
rect 3401 21821 3431 21877
rect 3487 21821 3491 21877
rect 2911 21797 3491 21821
rect 2911 21741 2915 21797
rect 2971 21741 3001 21797
rect 3057 21741 3087 21797
rect 3143 21741 3173 21797
rect 3229 21741 3259 21797
rect 3315 21741 3345 21797
rect 3401 21741 3431 21797
rect 3487 21741 3491 21797
rect 2911 21717 3491 21741
rect 2911 21661 2915 21717
rect 2971 21661 3001 21717
rect 3057 21661 3087 21717
rect 3143 21661 3173 21717
rect 3229 21661 3259 21717
rect 3315 21661 3345 21717
rect 3401 21661 3431 21717
rect 3487 21661 3491 21717
rect 2911 21637 3491 21661
rect 2911 21581 2915 21637
rect 2971 21581 3001 21637
rect 3057 21581 3087 21637
rect 3143 21581 3173 21637
rect 3229 21581 3259 21637
rect 3315 21581 3345 21637
rect 3401 21581 3431 21637
rect 3487 21581 3491 21637
rect 2911 21557 3491 21581
rect 2911 21501 2915 21557
rect 2971 21501 3001 21557
rect 3057 21501 3087 21557
rect 3143 21501 3173 21557
rect 3229 21501 3259 21557
rect 3315 21501 3345 21557
rect 3401 21501 3431 21557
rect 3487 21501 3491 21557
rect 2911 21477 3491 21501
rect 2911 21421 2915 21477
rect 2971 21421 3001 21477
rect 3057 21421 3087 21477
rect 3143 21421 3173 21477
rect 3229 21421 3259 21477
rect 3315 21421 3345 21477
rect 3401 21421 3431 21477
rect 3487 21421 3491 21477
rect 2911 21397 3491 21421
rect 2911 21341 2915 21397
rect 2971 21341 3001 21397
rect 3057 21341 3087 21397
rect 3143 21341 3173 21397
rect 3229 21341 3259 21397
rect 3315 21341 3345 21397
rect 3401 21341 3431 21397
rect 3487 21341 3491 21397
rect 2911 21317 3491 21341
rect 2911 21261 2915 21317
rect 2971 21261 3001 21317
rect 3057 21261 3087 21317
rect 3143 21261 3173 21317
rect 3229 21261 3259 21317
rect 3315 21261 3345 21317
rect 3401 21261 3431 21317
rect 3487 21261 3491 21317
rect 4711 21296 4763 28859
tri 4763 28825 4797 28859 nw
tri 5520 28825 5532 28837 se
rect 5532 28825 5584 29067
tri 5584 29065 5586 29067 nw
tri 5498 28803 5520 28825 se
rect 5520 28803 5584 28825
rect 4830 28751 5584 28803
rect 5662 29015 5668 29067
rect 5720 29015 5732 29067
rect 5784 29015 5790 29067
rect 4830 21294 4882 28751
tri 4882 28717 4916 28751 nw
tri 5636 28717 5662 28743 se
rect 5662 28717 5714 29015
tri 5714 28981 5748 29015 nw
rect 6890 28963 7528 29376
tri 5628 28709 5636 28717 se
rect 5636 28709 5714 28717
rect 5005 28657 5714 28709
rect 5005 28052 5057 28657
tri 5057 28623 5091 28657 nw
rect 5899 24037 6479 24046
rect 5899 23981 5903 24037
rect 5959 23981 5989 24037
rect 6045 23981 6075 24037
rect 6131 23981 6161 24037
rect 6217 23981 6247 24037
rect 6303 23981 6333 24037
rect 6389 23981 6419 24037
rect 6475 23981 6479 24037
rect 5899 23957 6479 23981
rect 5899 23901 5903 23957
rect 5959 23901 5989 23957
rect 6045 23901 6075 23957
rect 6131 23901 6161 23957
rect 6217 23901 6247 23957
rect 6303 23901 6333 23957
rect 6389 23901 6419 23957
rect 6475 23901 6479 23957
rect 5899 23877 6479 23901
rect 5899 23821 5903 23877
rect 5959 23821 5989 23877
rect 6045 23821 6075 23877
rect 6131 23821 6161 23877
rect 6217 23821 6247 23877
rect 6303 23821 6333 23877
rect 6389 23821 6419 23877
rect 6475 23821 6479 23877
rect 5899 23797 6479 23821
rect 5899 23741 5903 23797
rect 5959 23741 5989 23797
rect 6045 23741 6075 23797
rect 6131 23741 6161 23797
rect 6217 23741 6247 23797
rect 6303 23741 6333 23797
rect 6389 23741 6419 23797
rect 6475 23741 6479 23797
rect 5899 23717 6479 23741
rect 5899 23661 5903 23717
rect 5959 23661 5989 23717
rect 6045 23661 6075 23717
rect 6131 23661 6161 23717
rect 6217 23661 6247 23717
rect 6303 23661 6333 23717
rect 6389 23661 6419 23717
rect 6475 23661 6479 23717
rect 5899 23637 6479 23661
rect 5899 23581 5903 23637
rect 5959 23581 5989 23637
rect 6045 23581 6075 23637
rect 6131 23581 6161 23637
rect 6217 23581 6247 23637
rect 6303 23581 6333 23637
rect 6389 23581 6419 23637
rect 6475 23581 6479 23637
rect 5899 23557 6479 23581
rect 5899 23501 5903 23557
rect 5959 23501 5989 23557
rect 6045 23501 6075 23557
rect 6131 23501 6161 23557
rect 6217 23501 6247 23557
rect 6303 23501 6333 23557
rect 6389 23501 6419 23557
rect 6475 23501 6479 23557
rect 5899 23477 6479 23501
rect 5899 23421 5903 23477
rect 5959 23421 5989 23477
rect 6045 23421 6075 23477
rect 6131 23421 6161 23477
rect 6217 23421 6247 23477
rect 6303 23421 6333 23477
rect 6389 23421 6419 23477
rect 6475 23421 6479 23477
rect 5899 23397 6479 23421
rect 5899 23341 5903 23397
rect 5959 23341 5989 23397
rect 6045 23341 6075 23397
rect 6131 23341 6161 23397
rect 6217 23341 6247 23397
rect 6303 23341 6333 23397
rect 6389 23341 6419 23397
rect 6475 23341 6479 23397
rect 5899 23317 6479 23341
rect 5899 23261 5903 23317
rect 5959 23261 5989 23317
rect 6045 23261 6075 23317
rect 6131 23261 6161 23317
rect 6217 23261 6247 23317
rect 6303 23261 6333 23317
rect 6389 23261 6419 23317
rect 6475 23261 6479 23317
rect 5899 23237 6479 23261
rect 5899 23181 5903 23237
rect 5959 23181 5989 23237
rect 6045 23181 6075 23237
rect 6131 23181 6161 23237
rect 6217 23181 6247 23237
rect 6303 23181 6333 23237
rect 6389 23181 6419 23237
rect 6475 23181 6479 23237
rect 5899 23157 6479 23181
rect 5899 23101 5903 23157
rect 5959 23101 5989 23157
rect 6045 23101 6075 23157
rect 6131 23101 6161 23157
rect 6217 23101 6247 23157
rect 6303 23101 6333 23157
rect 6389 23101 6419 23157
rect 6475 23101 6479 23157
rect 5899 23077 6479 23101
rect 5899 23021 5903 23077
rect 5959 23021 5989 23077
rect 6045 23021 6075 23077
rect 6131 23021 6161 23077
rect 6217 23021 6247 23077
rect 6303 23021 6333 23077
rect 6389 23021 6419 23077
rect 6475 23021 6479 23077
rect 5899 22997 6479 23021
rect 5899 22941 5903 22997
rect 5959 22941 5989 22997
rect 6045 22941 6075 22997
rect 6131 22941 6161 22997
rect 6217 22941 6247 22997
rect 6303 22941 6333 22997
rect 6389 22941 6419 22997
rect 6475 22941 6479 22997
rect 5899 22917 6479 22941
rect 5899 22861 5903 22917
rect 5959 22861 5989 22917
rect 6045 22861 6075 22917
rect 6131 22861 6161 22917
rect 6217 22861 6247 22917
rect 6303 22861 6333 22917
rect 6389 22861 6419 22917
rect 6475 22861 6479 22917
rect 5899 22837 6479 22861
rect 5899 22781 5903 22837
rect 5959 22781 5989 22837
rect 6045 22781 6075 22837
rect 6131 22781 6161 22837
rect 6217 22781 6247 22837
rect 6303 22781 6333 22837
rect 6389 22781 6419 22837
rect 6475 22781 6479 22837
rect 5899 22757 6479 22781
rect 5899 22701 5903 22757
rect 5959 22701 5989 22757
rect 6045 22701 6075 22757
rect 6131 22701 6161 22757
rect 6217 22701 6247 22757
rect 6303 22701 6333 22757
rect 6389 22701 6419 22757
rect 6475 22701 6479 22757
rect 5899 22677 6479 22701
rect 5899 22621 5903 22677
rect 5959 22621 5989 22677
rect 6045 22621 6075 22677
rect 6131 22621 6161 22677
rect 6217 22621 6247 22677
rect 6303 22621 6333 22677
rect 6389 22621 6419 22677
rect 6475 22621 6479 22677
rect 5899 22597 6479 22621
rect 5899 22541 5903 22597
rect 5959 22541 5989 22597
rect 6045 22541 6075 22597
rect 6131 22541 6161 22597
rect 6217 22541 6247 22597
rect 6303 22541 6333 22597
rect 6389 22541 6419 22597
rect 6475 22541 6479 22597
rect 5899 22517 6479 22541
rect 5899 22461 5903 22517
rect 5959 22461 5989 22517
rect 6045 22461 6075 22517
rect 6131 22461 6161 22517
rect 6217 22461 6247 22517
rect 6303 22461 6333 22517
rect 6389 22461 6419 22517
rect 6475 22461 6479 22517
rect 5899 22437 6479 22461
rect 5899 22381 5903 22437
rect 5959 22381 5989 22437
rect 6045 22381 6075 22437
rect 6131 22381 6161 22437
rect 6217 22381 6247 22437
rect 6303 22381 6333 22437
rect 6389 22381 6419 22437
rect 6475 22381 6479 22437
rect 5899 22357 6479 22381
rect 5899 22301 5903 22357
rect 5959 22301 5989 22357
rect 6045 22301 6075 22357
rect 6131 22301 6161 22357
rect 6217 22301 6247 22357
rect 6303 22301 6333 22357
rect 6389 22301 6419 22357
rect 6475 22301 6479 22357
rect 5899 22277 6479 22301
rect 5899 22221 5903 22277
rect 5959 22221 5989 22277
rect 6045 22221 6075 22277
rect 6131 22221 6161 22277
rect 6217 22221 6247 22277
rect 6303 22221 6333 22277
rect 6389 22221 6419 22277
rect 6475 22221 6479 22277
rect 5899 22197 6479 22221
rect 5899 22141 5903 22197
rect 5959 22141 5989 22197
rect 6045 22141 6075 22197
rect 6131 22141 6161 22197
rect 6217 22141 6247 22197
rect 6303 22141 6333 22197
rect 6389 22141 6419 22197
rect 6475 22141 6479 22197
rect 5899 22117 6479 22141
rect 5899 22061 5903 22117
rect 5959 22061 5989 22117
rect 6045 22061 6075 22117
rect 6131 22061 6161 22117
rect 6217 22061 6247 22117
rect 6303 22061 6333 22117
rect 6389 22061 6419 22117
rect 6475 22061 6479 22117
rect 5899 22037 6479 22061
rect 5899 21981 5903 22037
rect 5959 21981 5989 22037
rect 6045 21981 6075 22037
rect 6131 21981 6161 22037
rect 6217 21981 6247 22037
rect 6303 21981 6333 22037
rect 6389 21981 6419 22037
rect 6475 21981 6479 22037
rect 5899 21957 6479 21981
rect 5899 21901 5903 21957
rect 5959 21901 5989 21957
rect 6045 21901 6075 21957
rect 6131 21901 6161 21957
rect 6217 21901 6247 21957
rect 6303 21901 6333 21957
rect 6389 21901 6419 21957
rect 6475 21901 6479 21957
rect 5899 21877 6479 21901
rect 5899 21821 5903 21877
rect 5959 21821 5989 21877
rect 6045 21821 6075 21877
rect 6131 21821 6161 21877
rect 6217 21821 6247 21877
rect 6303 21821 6333 21877
rect 6389 21821 6419 21877
rect 6475 21821 6479 21877
rect 5899 21797 6479 21821
rect 5899 21741 5903 21797
rect 5959 21741 5989 21797
rect 6045 21741 6075 21797
rect 6131 21741 6161 21797
rect 6217 21741 6247 21797
rect 6303 21741 6333 21797
rect 6389 21741 6419 21797
rect 6475 21741 6479 21797
rect 5899 21717 6479 21741
rect 5899 21661 5903 21717
rect 5959 21661 5989 21717
rect 6045 21661 6075 21717
rect 6131 21661 6161 21717
rect 6217 21661 6247 21717
rect 6303 21661 6333 21717
rect 6389 21661 6419 21717
rect 6475 21661 6479 21717
rect 5899 21637 6479 21661
rect 5899 21581 5903 21637
rect 5959 21581 5989 21637
rect 6045 21581 6075 21637
rect 6131 21581 6161 21637
rect 6217 21581 6247 21637
rect 6303 21581 6333 21637
rect 6389 21581 6419 21637
rect 6475 21581 6479 21637
rect 5899 21557 6479 21581
rect 5899 21501 5903 21557
rect 5959 21501 5989 21557
rect 6045 21501 6075 21557
rect 6131 21501 6161 21557
rect 6217 21501 6247 21557
rect 6303 21501 6333 21557
rect 6389 21501 6419 21557
rect 6475 21501 6479 21557
rect 5899 21477 6479 21501
rect 5899 21421 5903 21477
rect 5959 21421 5989 21477
rect 6045 21421 6075 21477
rect 6131 21421 6161 21477
rect 6217 21421 6247 21477
rect 6303 21421 6333 21477
rect 6389 21421 6419 21477
rect 6475 21421 6479 21477
rect 5899 21397 6479 21421
rect 5899 21341 5903 21397
rect 5959 21341 5989 21397
rect 6045 21341 6075 21397
rect 6131 21341 6161 21397
rect 6217 21341 6247 21397
rect 6303 21341 6333 21397
rect 6389 21341 6419 21397
rect 6475 21341 6479 21397
rect 5899 21317 6479 21341
rect 2911 21237 3491 21261
rect 2911 21181 2915 21237
rect 2971 21181 3001 21237
rect 3057 21181 3087 21237
rect 3143 21181 3173 21237
rect 3229 21181 3259 21237
rect 3315 21181 3345 21237
rect 3401 21181 3431 21237
rect 3487 21181 3491 21237
rect 2911 21157 3491 21181
rect 2911 21101 2915 21157
rect 2971 21101 3001 21157
rect 3057 21101 3087 21157
rect 3143 21101 3173 21157
rect 3229 21101 3259 21157
rect 3315 21101 3345 21157
rect 3401 21101 3431 21157
rect 3487 21101 3491 21157
rect 2911 21077 3491 21101
rect 2911 21021 2915 21077
rect 2971 21021 3001 21077
rect 3057 21021 3087 21077
rect 3143 21021 3173 21077
rect 3229 21021 3259 21077
rect 3315 21021 3345 21077
rect 3401 21021 3431 21077
rect 3487 21021 3491 21077
rect 2911 20997 3491 21021
rect 2911 20941 2915 20997
rect 2971 20941 3001 20997
rect 3057 20941 3087 20997
rect 3143 20941 3173 20997
rect 3229 20941 3259 20997
rect 3315 20941 3345 20997
rect 3401 20941 3431 20997
rect 3487 20941 3491 20997
rect 2911 20917 3491 20941
rect 2911 20861 2915 20917
rect 2971 20861 3001 20917
rect 3057 20861 3087 20917
rect 3143 20861 3173 20917
rect 3229 20861 3259 20917
rect 3315 20861 3345 20917
rect 3401 20861 3431 20917
rect 3487 20861 3491 20917
rect 2911 20837 3491 20861
rect 2911 20781 2915 20837
rect 2971 20781 3001 20837
rect 3057 20781 3087 20837
rect 3143 20781 3173 20837
rect 3229 20781 3259 20837
rect 3315 20781 3345 20837
rect 3401 20781 3431 20837
rect 3487 20781 3491 20837
rect 2911 20757 3491 20781
rect 2911 20701 2915 20757
rect 2971 20701 3001 20757
rect 3057 20701 3087 20757
rect 3143 20701 3173 20757
rect 3229 20701 3259 20757
rect 3315 20701 3345 20757
rect 3401 20701 3431 20757
rect 3487 20701 3491 20757
rect 2911 20677 3491 20701
rect 2911 20621 2915 20677
rect 2971 20621 3001 20677
rect 3057 20621 3087 20677
rect 3143 20621 3173 20677
rect 3229 20621 3259 20677
rect 3315 20621 3345 20677
rect 3401 20621 3431 20677
rect 3487 20621 3491 20677
rect 2911 20597 3491 20621
rect 2911 20541 2915 20597
rect 2971 20541 3001 20597
rect 3057 20541 3087 20597
rect 3143 20541 3173 20597
rect 3229 20541 3259 20597
rect 3315 20541 3345 20597
rect 3401 20541 3431 20597
rect 3487 20541 3491 20597
rect 2911 20517 3491 20541
rect 2911 20461 2915 20517
rect 2971 20461 3001 20517
rect 3057 20461 3087 20517
rect 3143 20461 3173 20517
rect 3229 20461 3259 20517
rect 3315 20461 3345 20517
rect 3401 20461 3431 20517
rect 3487 20461 3491 20517
rect 2911 20437 3491 20461
rect 2911 20381 2915 20437
rect 2971 20381 3001 20437
rect 3057 20381 3087 20437
rect 3143 20381 3173 20437
rect 3229 20381 3259 20437
rect 3315 20381 3345 20437
rect 3401 20381 3431 20437
rect 3487 20381 3491 20437
rect 2911 20357 3491 20381
rect 2911 20301 2915 20357
rect 2971 20301 3001 20357
rect 3057 20301 3087 20357
rect 3143 20301 3173 20357
rect 3229 20301 3259 20357
rect 3315 20301 3345 20357
rect 3401 20301 3431 20357
rect 3487 20301 3491 20357
rect 2911 20277 3491 20301
rect 2911 20221 2915 20277
rect 2971 20221 3001 20277
rect 3057 20221 3087 20277
rect 3143 20221 3173 20277
rect 3229 20221 3259 20277
rect 3315 20221 3345 20277
rect 3401 20221 3431 20277
rect 3487 20221 3491 20277
rect 2911 20197 3491 20221
rect 2911 20141 2915 20197
rect 2971 20141 3001 20197
rect 3057 20141 3087 20197
rect 3143 20141 3173 20197
rect 3229 20141 3259 20197
rect 3315 20141 3345 20197
rect 3401 20141 3431 20197
rect 3487 20141 3491 20197
rect 2911 20117 3491 20141
rect 2911 20061 2915 20117
rect 2971 20061 3001 20117
rect 3057 20061 3087 20117
rect 3143 20061 3173 20117
rect 3229 20061 3259 20117
rect 3315 20061 3345 20117
rect 3401 20061 3431 20117
rect 3487 20061 3491 20117
rect 2911 20037 3491 20061
rect 2911 19981 2915 20037
rect 2971 19981 3001 20037
rect 3057 19981 3087 20037
rect 3143 19981 3173 20037
rect 3229 19981 3259 20037
rect 3315 19981 3345 20037
rect 3401 19981 3431 20037
rect 3487 19981 3491 20037
rect 2911 19957 3491 19981
rect 2911 19901 2915 19957
rect 2971 19901 3001 19957
rect 3057 19901 3087 19957
rect 3143 19901 3173 19957
rect 3229 19901 3259 19957
rect 3315 19901 3345 19957
rect 3401 19901 3431 19957
rect 3487 19901 3491 19957
rect 2911 19877 3491 19901
rect 2911 19821 2915 19877
rect 2971 19821 3001 19877
rect 3057 19821 3087 19877
rect 3143 19821 3173 19877
rect 3229 19821 3259 19877
rect 3315 19821 3345 19877
rect 3401 19821 3431 19877
rect 3487 19821 3491 19877
rect 2911 19797 3491 19821
rect 2911 19741 2915 19797
rect 2971 19741 3001 19797
rect 3057 19741 3087 19797
rect 3143 19741 3173 19797
rect 3229 19741 3259 19797
rect 3315 19741 3345 19797
rect 3401 19741 3431 19797
rect 3487 19741 3491 19797
rect 2911 19717 3491 19741
rect 2911 19661 2915 19717
rect 2971 19661 3001 19717
rect 3057 19661 3087 19717
rect 3143 19661 3173 19717
rect 3229 19661 3259 19717
rect 3315 19661 3345 19717
rect 3401 19661 3431 19717
rect 3487 19661 3491 19717
rect 2911 19637 3491 19661
rect 2911 19581 2915 19637
rect 2971 19581 3001 19637
rect 3057 19581 3087 19637
rect 3143 19581 3173 19637
rect 3229 19581 3259 19637
rect 3315 19581 3345 19637
rect 3401 19581 3431 19637
rect 3487 19581 3491 19637
rect 2911 19557 3491 19581
rect 2911 19501 2915 19557
rect 2971 19501 3001 19557
rect 3057 19501 3087 19557
rect 3143 19501 3173 19557
rect 3229 19501 3259 19557
rect 3315 19501 3345 19557
rect 3401 19501 3431 19557
rect 3487 19501 3491 19557
rect 2911 19477 3491 19501
rect 2911 19421 2915 19477
rect 2971 19421 3001 19477
rect 3057 19421 3087 19477
rect 3143 19421 3173 19477
rect 3229 19421 3259 19477
rect 3315 19421 3345 19477
rect 3401 19421 3431 19477
rect 3487 19421 3491 19477
rect 2911 19397 3491 19421
rect 2911 19341 2915 19397
rect 2971 19341 3001 19397
rect 3057 19341 3087 19397
rect 3143 19341 3173 19397
rect 3229 19341 3259 19397
rect 3315 19341 3345 19397
rect 3401 19341 3431 19397
rect 3487 19341 3491 19397
rect 2911 19317 3491 19341
rect 2911 19261 2915 19317
rect 2971 19261 3001 19317
rect 3057 19261 3087 19317
rect 3143 19261 3173 19317
rect 3229 19261 3259 19317
rect 3315 19261 3345 19317
rect 3401 19261 3431 19317
rect 3487 19261 3491 19317
rect 2911 19252 3491 19261
rect 5899 21261 5903 21317
rect 5959 21261 5989 21317
rect 6045 21261 6075 21317
rect 6131 21261 6161 21317
rect 6217 21261 6247 21317
rect 6303 21261 6333 21317
rect 6389 21261 6419 21317
rect 6475 21261 6479 21317
rect 5899 21237 6479 21261
rect 5899 21181 5903 21237
rect 5959 21181 5989 21237
rect 6045 21181 6075 21237
rect 6131 21181 6161 21237
rect 6217 21181 6247 21237
rect 6303 21181 6333 21237
rect 6389 21181 6419 21237
rect 6475 21181 6479 21237
rect 5899 21157 6479 21181
rect 5899 21101 5903 21157
rect 5959 21101 5989 21157
rect 6045 21101 6075 21157
rect 6131 21101 6161 21157
rect 6217 21101 6247 21157
rect 6303 21101 6333 21157
rect 6389 21101 6419 21157
rect 6475 21101 6479 21157
rect 5899 21077 6479 21101
rect 5899 21021 5903 21077
rect 5959 21021 5989 21077
rect 6045 21021 6075 21077
rect 6131 21021 6161 21077
rect 6217 21021 6247 21077
rect 6303 21021 6333 21077
rect 6389 21021 6419 21077
rect 6475 21021 6479 21077
rect 5899 20997 6479 21021
rect 5899 20941 5903 20997
rect 5959 20941 5989 20997
rect 6045 20941 6075 20997
rect 6131 20941 6161 20997
rect 6217 20941 6247 20997
rect 6303 20941 6333 20997
rect 6389 20941 6419 20997
rect 6475 20941 6479 20997
rect 5899 20917 6479 20941
rect 5899 20861 5903 20917
rect 5959 20861 5989 20917
rect 6045 20861 6075 20917
rect 6131 20861 6161 20917
rect 6217 20861 6247 20917
rect 6303 20861 6333 20917
rect 6389 20861 6419 20917
rect 6475 20861 6479 20917
rect 5899 20837 6479 20861
rect 5899 20781 5903 20837
rect 5959 20781 5989 20837
rect 6045 20781 6075 20837
rect 6131 20781 6161 20837
rect 6217 20781 6247 20837
rect 6303 20781 6333 20837
rect 6389 20781 6419 20837
rect 6475 20781 6479 20837
rect 5899 20757 6479 20781
rect 5899 20701 5903 20757
rect 5959 20701 5989 20757
rect 6045 20701 6075 20757
rect 6131 20701 6161 20757
rect 6217 20701 6247 20757
rect 6303 20701 6333 20757
rect 6389 20701 6419 20757
rect 6475 20701 6479 20757
rect 5899 20677 6479 20701
rect 5899 20621 5903 20677
rect 5959 20621 5989 20677
rect 6045 20621 6075 20677
rect 6131 20621 6161 20677
rect 6217 20621 6247 20677
rect 6303 20621 6333 20677
rect 6389 20621 6419 20677
rect 6475 20621 6479 20677
rect 5899 20597 6479 20621
rect 5899 20541 5903 20597
rect 5959 20541 5989 20597
rect 6045 20541 6075 20597
rect 6131 20541 6161 20597
rect 6217 20541 6247 20597
rect 6303 20541 6333 20597
rect 6389 20541 6419 20597
rect 6475 20541 6479 20597
rect 5899 20517 6479 20541
rect 5899 20461 5903 20517
rect 5959 20461 5989 20517
rect 6045 20461 6075 20517
rect 6131 20461 6161 20517
rect 6217 20461 6247 20517
rect 6303 20461 6333 20517
rect 6389 20461 6419 20517
rect 6475 20461 6479 20517
rect 5899 20437 6479 20461
rect 5899 20381 5903 20437
rect 5959 20381 5989 20437
rect 6045 20381 6075 20437
rect 6131 20381 6161 20437
rect 6217 20381 6247 20437
rect 6303 20381 6333 20437
rect 6389 20381 6419 20437
rect 6475 20381 6479 20437
rect 5899 20357 6479 20381
rect 5899 20301 5903 20357
rect 5959 20301 5989 20357
rect 6045 20301 6075 20357
rect 6131 20301 6161 20357
rect 6217 20301 6247 20357
rect 6303 20301 6333 20357
rect 6389 20301 6419 20357
rect 6475 20301 6479 20357
rect 5899 20277 6479 20301
rect 5899 20221 5903 20277
rect 5959 20221 5989 20277
rect 6045 20221 6075 20277
rect 6131 20221 6161 20277
rect 6217 20221 6247 20277
rect 6303 20221 6333 20277
rect 6389 20221 6419 20277
rect 6475 20221 6479 20277
rect 5899 20197 6479 20221
rect 5899 20141 5903 20197
rect 5959 20141 5989 20197
rect 6045 20141 6075 20197
rect 6131 20141 6161 20197
rect 6217 20141 6247 20197
rect 6303 20141 6333 20197
rect 6389 20141 6419 20197
rect 6475 20141 6479 20197
rect 5899 20117 6479 20141
rect 5899 20061 5903 20117
rect 5959 20061 5989 20117
rect 6045 20061 6075 20117
rect 6131 20061 6161 20117
rect 6217 20061 6247 20117
rect 6303 20061 6333 20117
rect 6389 20061 6419 20117
rect 6475 20061 6479 20117
rect 5899 20037 6479 20061
rect 5899 19981 5903 20037
rect 5959 19981 5989 20037
rect 6045 19981 6075 20037
rect 6131 19981 6161 20037
rect 6217 19981 6247 20037
rect 6303 19981 6333 20037
rect 6389 19981 6419 20037
rect 6475 19981 6479 20037
rect 5899 19957 6479 19981
rect 5899 19901 5903 19957
rect 5959 19901 5989 19957
rect 6045 19901 6075 19957
rect 6131 19901 6161 19957
rect 6217 19901 6247 19957
rect 6303 19901 6333 19957
rect 6389 19901 6419 19957
rect 6475 19901 6479 19957
rect 5899 19877 6479 19901
rect 5899 19821 5903 19877
rect 5959 19821 5989 19877
rect 6045 19821 6075 19877
rect 6131 19821 6161 19877
rect 6217 19821 6247 19877
rect 6303 19821 6333 19877
rect 6389 19821 6419 19877
rect 6475 19821 6479 19877
rect 5899 19797 6479 19821
rect 5899 19741 5903 19797
rect 5959 19741 5989 19797
rect 6045 19741 6075 19797
rect 6131 19741 6161 19797
rect 6217 19741 6247 19797
rect 6303 19741 6333 19797
rect 6389 19741 6419 19797
rect 6475 19741 6479 19797
rect 5899 19717 6479 19741
rect 5899 19661 5903 19717
rect 5959 19661 5989 19717
rect 6045 19661 6075 19717
rect 6131 19661 6161 19717
rect 6217 19661 6247 19717
rect 6303 19661 6333 19717
rect 6389 19661 6419 19717
rect 6475 19661 6479 19717
rect 5899 19637 6479 19661
rect 5899 19581 5903 19637
rect 5959 19581 5989 19637
rect 6045 19581 6075 19637
rect 6131 19581 6161 19637
rect 6217 19581 6247 19637
rect 6303 19581 6333 19637
rect 6389 19581 6419 19637
rect 6475 19581 6479 19637
rect 5899 19557 6479 19581
rect 5899 19501 5903 19557
rect 5959 19501 5989 19557
rect 6045 19501 6075 19557
rect 6131 19501 6161 19557
rect 6217 19501 6247 19557
rect 6303 19501 6333 19557
rect 6389 19501 6419 19557
rect 6475 19501 6479 19557
rect 5899 19477 6479 19501
rect 5899 19421 5903 19477
rect 5959 19421 5989 19477
rect 6045 19421 6075 19477
rect 6131 19421 6161 19477
rect 6217 19421 6247 19477
rect 6303 19421 6333 19477
rect 6389 19421 6419 19477
rect 6475 19421 6479 19477
rect 5899 19397 6479 19421
rect 5899 19341 5903 19397
rect 5959 19341 5989 19397
rect 6045 19341 6075 19397
rect 6131 19341 6161 19397
rect 6217 19341 6247 19397
rect 6303 19341 6333 19397
rect 6389 19341 6419 19397
rect 6475 19341 6479 19397
rect 5899 19317 6479 19341
rect 5899 19261 5903 19317
rect 5959 19261 5989 19317
rect 6045 19261 6075 19317
rect 6131 19261 6161 19317
rect 6217 19261 6247 19317
rect 6303 19261 6333 19317
rect 6389 19261 6419 19317
rect 6475 19261 6479 19317
rect 5899 19252 6479 19261
rect 4998 18602 5004 18654
rect 5056 18623 5072 18654
rect 5063 18602 5072 18623
rect 5124 18623 5140 18654
rect 5124 18602 5133 18623
rect 5192 18602 5198 18654
rect 4998 18588 5007 18602
rect 5063 18588 5133 18602
rect 5189 18588 5198 18602
rect 4998 18536 5004 18588
rect 5063 18567 5072 18588
rect 5056 18536 5072 18567
rect 5124 18567 5133 18588
rect 5124 18536 5140 18567
rect 5192 18536 5198 18588
rect 1660 17767 8434 17776
rect 1716 17711 2526 17767
rect 2582 17711 2739 17767
rect 2795 17711 3605 17767
rect 3661 17711 5728 17767
rect 5784 17711 6594 17767
rect 6650 17711 6807 17767
rect 6863 17711 7673 17767
rect 7729 17745 8434 17767
rect 7729 17711 7843 17745
rect 1660 17689 7843 17711
rect 7899 17689 7949 17745
rect 8005 17689 8054 17745
rect 8110 17689 8159 17745
rect 8215 17689 8264 17745
rect 8320 17689 8369 17745
rect 8425 17689 8434 17745
rect 1660 17680 8434 17689
rect 1716 17624 2526 17680
rect 2582 17624 2739 17680
rect 2795 17624 3605 17680
rect 3661 17624 5728 17680
rect 5784 17624 6594 17680
rect 6650 17624 6807 17680
rect 6863 17624 7673 17680
rect 7729 17645 8434 17680
rect 7729 17624 7843 17645
rect 1660 17593 7843 17624
rect 1716 17537 2526 17593
rect 2582 17537 2739 17593
rect 2795 17537 3605 17593
rect 3661 17537 5728 17593
rect 5784 17537 6594 17593
rect 6650 17537 6807 17593
rect 6863 17537 7673 17593
rect 7729 17589 7843 17593
rect 7899 17589 7949 17645
rect 8005 17589 8054 17645
rect 8110 17589 8159 17645
rect 8215 17589 8264 17645
rect 8320 17589 8369 17645
rect 8425 17589 8434 17645
rect 7729 17545 8434 17589
rect 7729 17537 7843 17545
rect 1660 17505 7843 17537
rect 1716 17449 2526 17505
rect 2582 17449 2739 17505
rect 2795 17449 3605 17505
rect 3661 17449 5728 17505
rect 5784 17449 6594 17505
rect 6650 17449 6807 17505
rect 6863 17449 7673 17505
rect 7729 17489 7843 17505
rect 7899 17489 7949 17545
rect 8005 17489 8054 17545
rect 8110 17489 8159 17545
rect 8215 17489 8264 17545
rect 8320 17489 8369 17545
rect 8425 17489 8434 17545
rect 7729 17449 8434 17489
rect 1660 17445 8434 17449
rect 1660 17417 7843 17445
rect 1716 17361 2526 17417
rect 2582 17361 2739 17417
rect 2795 17361 3605 17417
rect 3661 17361 5728 17417
rect 5784 17361 6594 17417
rect 6650 17361 6807 17417
rect 6863 17361 7673 17417
rect 7729 17389 7843 17417
rect 7899 17389 7949 17445
rect 8005 17389 8054 17445
rect 8110 17389 8159 17445
rect 8215 17389 8264 17445
rect 8320 17389 8369 17445
rect 8425 17389 8434 17445
rect 7729 17361 8434 17389
rect 1660 17345 8434 17361
rect 1660 17329 7843 17345
rect 1716 17273 2526 17329
rect 2582 17273 2739 17329
rect 2795 17273 3605 17329
rect 3661 17273 5728 17329
rect 5784 17273 6594 17329
rect 6650 17273 6807 17329
rect 6863 17273 7673 17329
rect 7729 17289 7843 17329
rect 7899 17289 7949 17345
rect 8005 17289 8054 17345
rect 8110 17289 8159 17345
rect 8215 17289 8264 17345
rect 8320 17289 8369 17345
rect 8425 17289 8434 17345
rect 7729 17273 8434 17289
rect 1660 17245 8434 17273
rect 1660 17241 7843 17245
rect 1716 17185 2526 17241
rect 2582 17185 2739 17241
rect 2795 17185 3605 17241
rect 3661 17185 5728 17241
rect 5784 17185 6594 17241
rect 6650 17185 6807 17241
rect 6863 17185 7673 17241
rect 7729 17189 7843 17241
rect 7899 17189 7949 17245
rect 8005 17189 8054 17245
rect 8110 17189 8159 17245
rect 8215 17189 8264 17245
rect 8320 17189 8369 17245
rect 8425 17189 8434 17245
rect 7729 17185 8434 17189
rect 1660 17176 8434 17185
rect 4994 16425 5003 16481
rect 5059 16429 5072 16481
rect 5124 16429 5137 16481
rect 5059 16425 5137 16429
rect 5193 16425 5202 16481
rect 7044 15872 7843 15879
rect 7096 15820 7160 15872
rect 7212 15823 7843 15872
rect 7899 15823 7949 15879
rect 8005 15823 8054 15879
rect 8110 15823 8159 15879
rect 8215 15823 8264 15879
rect 8320 15823 8369 15879
rect 8425 15823 8434 15879
rect 7212 15820 8434 15823
rect 7044 15805 8434 15820
rect 7096 15753 7160 15805
rect 7212 15753 8434 15805
rect 1648 15736 1700 15742
rect 7044 15737 8434 15753
tri 1700 15685 1715 15700 sw
rect 7096 15685 7160 15737
rect 7212 15735 8434 15737
rect 7212 15685 7843 15735
rect 1700 15684 1715 15685
rect 1648 15672 1715 15684
rect 1700 15666 1715 15672
tri 1715 15666 1734 15685 sw
rect 7044 15679 7843 15685
rect 7899 15679 7949 15735
rect 8005 15679 8054 15735
rect 8110 15679 8159 15735
rect 8215 15679 8264 15735
rect 8320 15679 8369 15735
rect 8425 15679 8434 15735
rect 1700 15620 3550 15666
rect 1648 15614 3550 15620
rect 4416 15514 4422 15566
rect 4481 15514 4490 15566
rect 4542 15514 4551 15566
rect 4610 15514 4616 15566
rect 4416 15510 4425 15514
rect 4481 15510 4551 15514
rect 4607 15510 4616 15514
rect 2083 15457 2089 15509
rect 2141 15457 2173 15509
rect 2225 15457 2257 15509
rect 2309 15457 2341 15509
rect 2393 15457 2425 15509
rect 2477 15457 2882 15509
rect 2934 15457 2995 15509
rect 3047 15457 3107 15509
rect 3159 15457 3165 15509
rect 2083 15419 3165 15457
rect 4416 15486 4616 15510
rect 4416 15482 4425 15486
rect 4481 15482 4551 15486
rect 4607 15482 4616 15486
rect 4416 15430 4422 15482
rect 4481 15430 4490 15482
rect 4542 15430 4551 15482
rect 4610 15430 4616 15482
rect 2083 15367 2089 15419
rect 2141 15367 2173 15419
rect 2225 15367 2257 15419
rect 2309 15367 2341 15419
rect 2393 15367 2425 15419
rect 2477 15367 2882 15419
rect 2934 15367 2995 15419
rect 3047 15367 3107 15419
rect 3159 15367 3165 15419
rect 1648 15297 1700 15303
rect 1648 15233 1700 15245
tri 1700 15225 1734 15259 sw
rect 1700 15181 3354 15225
rect 1648 15175 3354 15181
tri 3320 15141 3354 15175 ne
rect 1564 14838 1616 14844
rect 1564 14774 1616 14786
tri 1616 14768 1650 14802 sw
rect 1616 14722 4906 14768
rect 1564 14716 4906 14722
tri 4870 14684 4902 14716 ne
rect 4902 14684 4904 14716
rect 954 14628 963 14684
rect 1019 14628 1069 14684
rect 1125 14628 1174 14684
rect 1230 14628 1279 14684
rect 1335 14628 1384 14684
rect 1440 14628 1489 14684
rect 1545 14678 4077 14684
tri 4902 14682 4904 14684 ne
rect 1545 14628 3877 14678
rect 954 14626 3877 14628
rect 3929 14626 3951 14678
rect 4003 14626 4025 14678
rect 954 14610 4077 14626
rect 954 14558 3877 14610
rect 3929 14558 3951 14610
rect 4003 14558 4025 14610
rect 954 14542 4077 14558
rect 954 14540 3877 14542
rect 954 14484 963 14540
rect 1019 14484 1069 14540
rect 1125 14484 1174 14540
rect 1230 14484 1279 14540
rect 1335 14484 1384 14540
rect 1440 14484 1489 14540
rect 1545 14490 3877 14540
rect 3929 14490 3951 14542
rect 4003 14490 4025 14542
rect 1545 14484 4077 14490
rect 4416 14371 4422 14423
rect 4481 14371 4490 14423
rect 4542 14371 4551 14423
rect 4610 14371 4616 14423
rect 4416 14367 4425 14371
rect 4481 14367 4551 14371
rect 4607 14367 4616 14371
rect 4416 14343 4616 14367
rect 4416 14339 4425 14343
rect 4481 14339 4551 14343
rect 4607 14339 4616 14343
rect 4416 14287 4422 14339
rect 4481 14287 4490 14339
rect 4542 14287 4551 14339
rect 4610 14287 4616 14339
rect 7044 14153 7843 14160
rect 7096 14101 7160 14153
rect 7212 14104 7843 14153
rect 7899 14104 7949 14160
rect 8005 14104 8054 14160
rect 8110 14104 8159 14160
rect 8215 14104 8264 14160
rect 8320 14104 8369 14160
rect 8425 14104 8434 14160
rect 7212 14101 8434 14104
rect 7044 14086 8434 14101
rect 7096 14034 7160 14086
rect 7212 14034 8434 14086
rect 7044 14018 8434 14034
rect 7096 13966 7160 14018
rect 7212 14016 8434 14018
rect 7212 13966 7843 14016
rect 7044 13960 7843 13966
rect 7899 13960 7949 14016
rect 8005 13960 8054 14016
rect 8110 13960 8159 14016
rect 8215 13960 8264 14016
rect 8320 13960 8369 14016
rect 8425 13960 8434 14016
rect 453 13739 462 13795
rect 518 13739 571 13795
rect 627 13739 680 13795
rect 736 13739 788 13795
rect 844 13789 3023 13795
rect 844 13739 2944 13789
rect 453 13737 2944 13739
rect 2996 13737 3023 13789
rect 453 13721 3023 13737
rect 453 13669 2944 13721
rect 2996 13669 3023 13721
rect 453 13653 3023 13669
rect 453 13651 2944 13653
rect 453 13595 462 13651
rect 518 13595 571 13651
rect 627 13595 680 13651
rect 736 13595 788 13651
rect 844 13601 2944 13651
rect 2996 13601 3023 13653
rect 844 13595 3023 13601
rect 7044 13431 7843 13438
rect 7096 13379 7160 13431
rect 7212 13382 7843 13431
rect 7899 13382 7949 13438
rect 8005 13382 8054 13438
rect 8110 13382 8159 13438
rect 8215 13382 8264 13438
rect 8320 13382 8369 13438
rect 8425 13382 8434 13438
rect 7212 13379 8434 13382
rect 7044 13364 8434 13379
rect 7096 13312 7160 13364
rect 7212 13312 8434 13364
rect 7044 13296 8434 13312
rect 7096 13244 7160 13296
rect 7212 13294 8434 13296
rect 7212 13244 7843 13294
rect 7044 13238 7843 13244
rect 7899 13238 7949 13294
rect 8005 13238 8054 13294
rect 8110 13238 8159 13294
rect 8215 13238 8264 13294
rect 8320 13238 8369 13294
rect 8425 13238 8434 13294
rect 4416 12990 4422 13042
rect 4481 12990 4490 13042
rect 4542 12990 4551 13042
rect 4610 12990 4616 13042
rect 4416 12986 4425 12990
rect 4481 12986 4551 12990
rect 4607 12986 4616 12990
rect 4416 12962 4616 12986
rect 4416 12958 4425 12962
rect 4481 12958 4551 12962
rect 4607 12958 4616 12962
rect 4416 12906 4422 12958
rect 4481 12906 4490 12958
rect 4542 12906 4551 12958
rect 4610 12906 4616 12958
rect 954 12802 963 12858
rect 1019 12802 1069 12858
rect 1125 12802 1174 12858
rect 1230 12802 1279 12858
rect 1335 12802 1384 12858
rect 1440 12802 1489 12858
rect 1545 12852 4077 12858
rect 1545 12802 3877 12852
rect 954 12800 3877 12802
rect 3929 12800 3951 12852
rect 4003 12800 4025 12852
rect 954 12784 4077 12800
rect 954 12732 3877 12784
rect 3929 12732 3951 12784
rect 4003 12732 4025 12784
rect 954 12716 4077 12732
rect 954 12714 3877 12716
rect 954 12658 963 12714
rect 1019 12658 1069 12714
rect 1125 12658 1174 12714
rect 1230 12658 1279 12714
rect 1335 12658 1384 12714
rect 1440 12658 1489 12714
rect 1545 12664 3877 12714
rect 3929 12664 3951 12716
rect 4003 12664 4025 12716
rect 1545 12658 4077 12664
tri 4902 12658 4904 12660 se
tri 4870 12626 4902 12658 se
rect 4902 12626 4904 12658
rect 1900 12620 4906 12626
rect 1952 12574 4906 12620
rect 1900 12556 1952 12568
tri 1952 12540 1986 12574 nw
rect 1900 12498 1952 12504
rect 1900 12239 1952 12245
rect 1900 12175 1952 12187
tri 1952 12167 1986 12201 sw
tri 3320 12167 3354 12201 se
rect 1952 12123 3354 12167
rect 1900 12117 3354 12123
rect 2083 11923 2089 11975
rect 2141 11923 2173 11975
rect 2225 11923 2257 11975
rect 2309 11923 2341 11975
rect 2393 11923 2425 11975
rect 2477 11923 2882 11975
rect 2934 11923 2995 11975
rect 3047 11923 3107 11975
rect 3159 11923 3165 11975
rect 2083 11885 3165 11923
rect 2083 11833 2089 11885
rect 2141 11833 2173 11885
rect 2225 11833 2257 11885
rect 2309 11833 2341 11885
rect 2393 11833 2425 11885
rect 2477 11833 2882 11885
rect 2934 11833 2995 11885
rect 3047 11833 3107 11885
rect 3159 11833 3165 11885
rect 4416 11857 4422 11909
rect 4481 11857 4490 11909
rect 4542 11857 4551 11909
rect 4610 11857 4616 11909
rect 4416 11853 4425 11857
rect 4481 11853 4551 11857
rect 4607 11853 4616 11857
rect 4416 11829 4616 11853
rect 4416 11825 4425 11829
rect 4481 11825 4551 11829
rect 4607 11825 4616 11829
rect 1732 11798 1784 11804
rect 4416 11773 4422 11825
rect 4481 11773 4490 11825
rect 4542 11773 4551 11825
rect 4610 11773 4616 11825
rect 1732 11734 1784 11746
tri 1784 11728 1818 11762 sw
rect 1784 11682 3550 11728
rect 1732 11676 3550 11682
rect 7044 11632 7843 11639
rect 7096 11580 7160 11632
rect 7212 11583 7843 11632
rect 7899 11583 7949 11639
rect 8005 11583 8054 11639
rect 8110 11583 8159 11639
rect 8215 11583 8264 11639
rect 8320 11583 8369 11639
rect 8425 11583 8434 11639
rect 7212 11580 8434 11583
rect 7044 11565 8434 11580
rect 7096 11513 7160 11565
rect 7212 11513 8434 11565
rect 7044 11497 8434 11513
rect 4427 11409 4433 11461
rect 4427 11405 4436 11409
rect 4492 11405 4551 11461
rect 4610 11409 4616 11461
rect 7096 11445 7160 11497
rect 7212 11495 8434 11497
rect 7212 11445 7843 11495
rect 7044 11439 7843 11445
rect 7899 11439 7949 11495
rect 8005 11439 8054 11495
rect 8110 11439 8159 11495
rect 8215 11439 8264 11495
rect 8320 11439 8369 11495
rect 8425 11439 8434 11495
rect 4607 11405 4616 11409
rect 4427 11381 4616 11405
rect 4427 11377 4436 11381
rect 4427 11325 4433 11377
rect 4492 11325 4551 11381
rect 4607 11377 4616 11381
rect 4610 11325 4616 11377
rect 7044 10944 7843 10951
rect 7096 10892 7160 10944
rect 7212 10895 7843 10944
rect 7899 10895 7949 10951
rect 8005 10895 8054 10951
rect 8110 10895 8159 10951
rect 8215 10895 8264 10951
rect 8320 10895 8369 10951
rect 8425 10895 8434 10951
rect 7212 10892 8434 10895
rect 7044 10877 8434 10892
rect 7096 10825 7160 10877
rect 7212 10825 8434 10877
rect 7044 10809 8434 10825
rect 7096 10757 7160 10809
rect 7212 10807 8434 10809
rect 7212 10757 7843 10807
rect 7044 10751 7843 10757
rect 7899 10751 7949 10807
rect 8005 10751 8054 10807
rect 8110 10751 8159 10807
rect 8215 10751 8264 10807
rect 8320 10751 8369 10807
rect 8425 10751 8434 10807
rect 1312 10688 1364 10694
rect 1312 10624 1364 10636
tri 1364 10618 1398 10652 sw
rect 1364 10572 3574 10618
rect 1312 10566 3574 10572
rect 2083 10409 2089 10461
rect 2141 10409 2173 10461
rect 2225 10409 2257 10461
rect 2309 10409 2341 10461
rect 2393 10409 2425 10461
rect 2477 10409 2882 10461
rect 2934 10409 2995 10461
rect 3047 10409 3107 10461
rect 3159 10409 3165 10461
rect 2083 10371 3165 10409
rect 4416 10459 4422 10511
rect 4481 10459 4490 10511
rect 4542 10459 4551 10511
rect 4610 10459 4616 10511
rect 4416 10455 4425 10459
rect 4481 10455 4551 10459
rect 4607 10455 4616 10459
rect 4416 10431 4616 10455
rect 4416 10427 4425 10431
rect 4481 10427 4551 10431
rect 4607 10427 4616 10431
rect 4416 10375 4422 10427
rect 4481 10375 4490 10427
rect 4542 10375 4551 10427
rect 4610 10375 4616 10427
rect 2083 10319 2089 10371
rect 2141 10319 2173 10371
rect 2225 10319 2257 10371
rect 2309 10319 2341 10371
rect 2393 10319 2425 10371
rect 2477 10319 2882 10371
rect 2934 10319 2995 10371
rect 3047 10319 3107 10371
rect 3159 10319 3165 10371
rect 1312 10249 1364 10255
rect 1312 10185 1364 10197
tri 1364 10177 1398 10211 sw
rect 1364 10133 3354 10177
rect 1312 10127 3354 10133
tri 3320 10093 3354 10127 ne
rect 1480 9790 1532 9796
rect 1480 9726 1532 9738
tri 1532 9720 1566 9754 sw
rect 1532 9674 4906 9720
rect 1480 9668 4906 9674
tri 4870 9636 4902 9668 ne
rect 4902 9636 4904 9668
rect 954 9580 963 9636
rect 1019 9580 1069 9636
rect 1125 9580 1174 9636
rect 1230 9580 1279 9636
rect 1335 9580 1384 9636
rect 1440 9580 1489 9636
rect 1545 9630 4077 9636
tri 4902 9634 4904 9636 ne
rect 1545 9580 3877 9630
rect 954 9578 3877 9580
rect 3929 9578 3951 9630
rect 4003 9578 4025 9630
rect 954 9562 4077 9578
rect 954 9510 3877 9562
rect 3929 9510 3951 9562
rect 4003 9510 4025 9562
rect 954 9494 4077 9510
rect 954 9492 3877 9494
rect 954 9436 963 9492
rect 1019 9436 1069 9492
rect 1125 9436 1174 9492
rect 1230 9436 1279 9492
rect 1335 9436 1384 9492
rect 1440 9436 1489 9492
rect 1545 9442 3877 9492
rect 3929 9442 3951 9494
rect 4003 9442 4025 9494
rect 1545 9436 4077 9442
rect 4416 9337 4422 9389
rect 4481 9337 4490 9389
rect 4542 9337 4551 9389
rect 4610 9337 4616 9389
rect 4416 9333 4425 9337
rect 4481 9333 4551 9337
rect 4607 9333 4616 9337
rect 4416 9309 4616 9333
rect 4416 9305 4425 9309
rect 4481 9305 4551 9309
rect 4607 9305 4616 9309
rect 4416 9253 4422 9305
rect 4481 9253 4490 9305
rect 4542 9253 4551 9305
rect 4610 9253 4616 9305
rect 315 9241 431 9247
rect 367 9238 379 9241
rect 376 9189 379 9238
rect 315 9182 320 9189
rect 376 9182 431 9189
rect 315 9175 431 9182
rect 367 9153 379 9175
rect 376 9123 379 9153
rect 315 9109 320 9123
rect 376 9109 431 9123
rect 376 9097 379 9109
rect 367 9068 379 9097
rect 376 9057 379 9068
rect 315 9043 320 9057
rect 376 9043 431 9057
rect 376 9012 379 9043
rect 367 8991 379 9012
rect 315 8983 431 8991
rect 315 8977 320 8983
rect 376 8977 431 8983
rect 376 8927 379 8977
rect 367 8925 379 8927
rect 315 8911 431 8925
rect 367 8898 379 8911
rect 376 8859 379 8898
rect 315 8844 320 8859
rect 376 8844 431 8859
rect 376 8842 379 8844
rect 367 8812 379 8842
rect 376 8792 379 8812
rect 315 8777 320 8792
rect 376 8777 431 8792
rect 376 8756 379 8777
rect 367 8726 379 8756
rect 376 8725 379 8726
rect 2083 9241 2483 9247
rect 2083 9238 2085 9241
rect 2137 9238 2171 9241
rect 2223 9238 2257 9241
rect 2083 9182 2084 9238
rect 2140 9189 2171 9238
rect 2254 9189 2257 9238
rect 2309 9238 2343 9241
rect 2395 9238 2429 9241
rect 2481 9238 2483 9241
rect 2309 9189 2312 9238
rect 2395 9189 2426 9238
rect 2140 9182 2198 9189
rect 2254 9182 2312 9189
rect 2368 9182 2426 9189
rect 2482 9182 2483 9238
rect 8532 9241 9228 9247
rect 8532 9238 8534 9241
rect 8586 9238 8598 9241
rect 8650 9238 8662 9241
rect 8714 9238 8726 9241
rect 8778 9238 8790 9241
rect 8842 9238 8854 9241
rect 8906 9238 8918 9241
rect 8970 9238 8982 9241
rect 9034 9238 9046 9241
rect 9098 9238 9110 9241
rect 9162 9238 9174 9241
rect 9226 9238 9228 9241
rect 2083 9160 2483 9182
rect 2083 9108 2085 9160
rect 2137 9108 2171 9160
rect 2223 9108 2257 9160
rect 2309 9108 2343 9160
rect 2395 9108 2429 9160
rect 2481 9108 2483 9160
rect 2083 9106 2483 9108
rect 2083 9050 2084 9106
rect 2140 9079 2198 9106
rect 2254 9079 2312 9106
rect 2368 9079 2426 9106
rect 2140 9050 2171 9079
rect 2254 9050 2257 9079
rect 2083 9027 2085 9050
rect 2137 9027 2171 9050
rect 2223 9027 2257 9050
rect 2309 9050 2312 9079
rect 2395 9050 2426 9079
rect 2482 9050 2483 9106
rect 2309 9027 2343 9050
rect 2395 9027 2429 9050
rect 2481 9027 2483 9050
rect 2083 8997 2483 9027
rect 7044 9198 7843 9205
rect 7096 9146 7160 9198
rect 7212 9149 7843 9198
rect 7899 9149 7949 9205
rect 8005 9149 8054 9205
rect 8110 9149 8159 9205
rect 8215 9149 8264 9205
rect 8320 9149 8369 9205
rect 8425 9149 8434 9205
rect 7212 9146 8434 9149
rect 7044 9131 8434 9146
rect 7096 9079 7160 9131
rect 7212 9079 8434 9131
rect 7044 9063 8434 9079
rect 7096 9011 7160 9063
rect 7212 9061 8434 9063
rect 7212 9011 7843 9061
rect 7044 9005 7843 9011
rect 7899 9005 7949 9061
rect 8005 9005 8054 9061
rect 8110 9005 8159 9061
rect 8215 9005 8264 9061
rect 8320 9005 8369 9061
rect 8425 9005 8434 9061
rect 8588 9189 8598 9238
rect 8842 9189 8852 9238
rect 8908 9189 8918 9238
rect 9162 9189 9172 9238
rect 8588 9182 8612 9189
rect 8668 9182 8692 9189
rect 8748 9182 8772 9189
rect 8828 9182 8852 9189
rect 8908 9182 8932 9189
rect 8988 9182 9012 9189
rect 9068 9182 9092 9189
rect 9148 9182 9172 9189
rect 8532 9175 9228 9182
rect 8532 9153 8534 9175
rect 8586 9153 8598 9175
rect 8650 9153 8662 9175
rect 8714 9153 8726 9175
rect 8778 9153 8790 9175
rect 8842 9153 8854 9175
rect 8906 9153 8918 9175
rect 8970 9153 8982 9175
rect 9034 9153 9046 9175
rect 9098 9153 9110 9175
rect 9162 9153 9174 9175
rect 9226 9153 9228 9175
rect 8588 9123 8598 9153
rect 8842 9123 8852 9153
rect 8908 9123 8918 9153
rect 9162 9123 9172 9153
rect 8588 9109 8612 9123
rect 8668 9109 8692 9123
rect 8748 9109 8772 9123
rect 8828 9109 8852 9123
rect 8908 9109 8932 9123
rect 8988 9109 9012 9123
rect 9068 9109 9092 9123
rect 9148 9109 9172 9123
rect 8588 9097 8598 9109
rect 8842 9097 8852 9109
rect 8908 9097 8918 9109
rect 9162 9097 9172 9109
rect 8532 9068 8534 9097
rect 8586 9068 8598 9097
rect 8650 9068 8662 9097
rect 8714 9068 8726 9097
rect 8778 9068 8790 9097
rect 8842 9068 8854 9097
rect 8906 9068 8918 9097
rect 8970 9068 8982 9097
rect 9034 9068 9046 9097
rect 9098 9068 9110 9097
rect 9162 9068 9174 9097
rect 9226 9068 9228 9097
rect 8588 9057 8598 9068
rect 8842 9057 8852 9068
rect 8908 9057 8918 9068
rect 9162 9057 9172 9068
rect 8588 9043 8612 9057
rect 8668 9043 8692 9057
rect 8748 9043 8772 9057
rect 8828 9043 8852 9057
rect 8908 9043 8932 9057
rect 8988 9043 9012 9057
rect 9068 9043 9092 9057
rect 9148 9043 9172 9057
rect 8588 9012 8598 9043
rect 8842 9012 8852 9043
rect 8908 9012 8918 9043
rect 9162 9012 9172 9043
rect 2083 8973 2085 8997
rect 2137 8973 2171 8997
rect 2223 8973 2257 8997
rect 2083 8917 2084 8973
rect 2140 8945 2171 8973
rect 2254 8945 2257 8973
rect 2309 8973 2343 8997
rect 2395 8973 2429 8997
rect 2481 8973 2483 8997
rect 2309 8945 2312 8973
rect 2395 8945 2426 8973
rect 2140 8917 2198 8945
rect 2254 8917 2312 8945
rect 2368 8917 2426 8945
rect 2482 8917 2483 8973
rect 2083 8915 2483 8917
rect 2083 8863 2085 8915
rect 2137 8863 2171 8915
rect 2223 8863 2257 8915
rect 2309 8863 2343 8915
rect 2395 8863 2429 8915
rect 2481 8863 2483 8915
rect 2083 8840 2483 8863
rect 2083 8784 2084 8840
rect 2140 8833 2198 8840
rect 2254 8833 2312 8840
rect 2368 8833 2426 8840
rect 2140 8784 2171 8833
rect 2254 8784 2257 8833
rect 2083 8781 2085 8784
rect 2137 8781 2171 8784
rect 2223 8781 2257 8784
rect 2309 8784 2312 8833
rect 2395 8784 2426 8833
rect 2482 8784 2483 8840
rect 2309 8781 2343 8784
rect 2395 8781 2429 8784
rect 2481 8781 2483 8784
rect 2083 8775 2483 8781
rect 8532 8991 8534 9012
rect 8586 8991 8598 9012
rect 8650 8991 8662 9012
rect 8714 8991 8726 9012
rect 8778 8991 8790 9012
rect 8842 8991 8854 9012
rect 8906 8991 8918 9012
rect 8970 8991 8982 9012
rect 9034 8991 9046 9012
rect 9098 8991 9110 9012
rect 9162 8991 9174 9012
rect 9226 8991 9228 9012
rect 8532 8983 9228 8991
rect 8588 8977 8612 8983
rect 8668 8977 8692 8983
rect 8748 8977 8772 8983
rect 8828 8977 8852 8983
rect 8908 8977 8932 8983
rect 8988 8977 9012 8983
rect 9068 8977 9092 8983
rect 9148 8977 9172 8983
rect 8588 8927 8598 8977
rect 8842 8927 8852 8977
rect 8908 8927 8918 8977
rect 9162 8927 9172 8977
rect 8532 8925 8534 8927
rect 8586 8925 8598 8927
rect 8650 8925 8662 8927
rect 8714 8925 8726 8927
rect 8778 8925 8790 8927
rect 8842 8925 8854 8927
rect 8906 8925 8918 8927
rect 8970 8925 8982 8927
rect 9034 8925 9046 8927
rect 9098 8925 9110 8927
rect 9162 8925 9174 8927
rect 9226 8925 9228 8927
rect 8532 8911 9228 8925
rect 8532 8898 8534 8911
rect 8586 8898 8598 8911
rect 8650 8898 8662 8911
rect 8714 8898 8726 8911
rect 8778 8898 8790 8911
rect 8842 8898 8854 8911
rect 8906 8898 8918 8911
rect 8970 8898 8982 8911
rect 9034 8898 9046 8911
rect 9098 8898 9110 8911
rect 9162 8898 9174 8911
rect 9226 8898 9228 8911
rect 8588 8859 8598 8898
rect 8842 8859 8852 8898
rect 8908 8859 8918 8898
rect 9162 8859 9172 8898
rect 8588 8844 8612 8859
rect 8668 8844 8692 8859
rect 8748 8844 8772 8859
rect 8828 8844 8852 8859
rect 8908 8844 8932 8859
rect 8988 8844 9012 8859
rect 9068 8844 9092 8859
rect 9148 8844 9172 8859
rect 8588 8842 8598 8844
rect 8842 8842 8852 8844
rect 8908 8842 8918 8844
rect 9162 8842 9172 8844
rect 8532 8812 8534 8842
rect 8586 8812 8598 8842
rect 8650 8812 8662 8842
rect 8714 8812 8726 8842
rect 8778 8812 8790 8842
rect 8842 8812 8854 8842
rect 8906 8812 8918 8842
rect 8970 8812 8982 8842
rect 9034 8812 9046 8842
rect 9098 8812 9110 8842
rect 9162 8812 9174 8842
rect 9226 8812 9228 8842
rect 8588 8792 8598 8812
rect 8842 8792 8852 8812
rect 8908 8792 8918 8812
rect 9162 8792 9172 8812
rect 8588 8777 8612 8792
rect 8668 8777 8692 8792
rect 8748 8777 8772 8792
rect 8828 8777 8852 8792
rect 8908 8777 8932 8792
rect 8988 8777 9012 8792
rect 9068 8777 9092 8792
rect 9148 8777 9172 8792
rect 315 8710 320 8725
rect 376 8710 431 8725
rect 8588 8756 8598 8777
rect 8842 8756 8852 8777
rect 8908 8756 8918 8777
rect 9162 8756 9172 8777
rect 8532 8726 8534 8756
rect 8586 8726 8598 8756
rect 8650 8726 8662 8756
rect 8714 8726 8726 8756
rect 8778 8726 8790 8756
rect 8842 8726 8854 8756
rect 8906 8726 8918 8756
rect 8970 8726 8982 8756
rect 9034 8726 9046 8756
rect 9098 8726 9110 8756
rect 9162 8726 9174 8756
rect 9226 8726 9228 8756
rect 8588 8725 8598 8726
rect 8842 8725 8852 8726
rect 8908 8725 8918 8726
rect 9162 8725 9172 8726
rect 376 8670 379 8710
rect 367 8658 379 8670
rect 315 8643 431 8658
rect 367 8640 379 8643
rect 376 8591 379 8640
rect 315 8584 320 8591
rect 376 8584 431 8591
rect 315 8576 431 8584
rect 367 8554 379 8576
rect 376 8524 379 8554
rect 315 8509 320 8524
rect 376 8509 431 8524
rect 467 8660 476 8716
rect 532 8660 580 8716
rect 636 8660 684 8716
rect 740 8660 788 8716
rect 844 8710 3023 8716
rect 844 8660 2944 8710
rect 467 8658 2944 8660
rect 2996 8658 3023 8710
rect 467 8642 3023 8658
rect 467 8590 2944 8642
rect 2996 8590 3023 8642
rect 467 8574 3023 8590
rect 467 8572 2944 8574
rect 467 8516 476 8572
rect 532 8516 580 8572
rect 636 8516 684 8572
rect 740 8516 788 8572
rect 844 8522 2944 8572
rect 2996 8522 3023 8574
rect 844 8516 3023 8522
rect 8588 8710 8612 8725
rect 8668 8710 8692 8725
rect 8748 8710 8772 8725
rect 8828 8710 8852 8725
rect 8908 8710 8932 8725
rect 8988 8710 9012 8725
rect 9068 8710 9092 8725
rect 9148 8710 9172 8725
rect 8588 8670 8598 8710
rect 8842 8670 8852 8710
rect 8908 8670 8918 8710
rect 9162 8670 9172 8710
rect 8532 8658 8534 8670
rect 8586 8658 8598 8670
rect 8650 8658 8662 8670
rect 8714 8658 8726 8670
rect 8778 8658 8790 8670
rect 8842 8658 8854 8670
rect 8906 8658 8918 8670
rect 8970 8658 8982 8670
rect 9034 8658 9046 8670
rect 9098 8658 9110 8670
rect 9162 8658 9174 8670
rect 9226 8658 9228 8670
rect 8532 8643 9228 8658
rect 8532 8640 8534 8643
rect 8586 8640 8598 8643
rect 8650 8640 8662 8643
rect 8714 8640 8726 8643
rect 8778 8640 8790 8643
rect 8842 8640 8854 8643
rect 8906 8640 8918 8643
rect 8970 8640 8982 8643
rect 9034 8640 9046 8643
rect 9098 8640 9110 8643
rect 9162 8640 9174 8643
rect 9226 8640 9228 8643
rect 8588 8591 8598 8640
rect 8842 8591 8852 8640
rect 8908 8591 8918 8640
rect 9162 8591 9172 8640
rect 8588 8584 8612 8591
rect 8668 8584 8692 8591
rect 8748 8584 8772 8591
rect 8828 8584 8852 8591
rect 8908 8584 8932 8591
rect 8988 8584 9012 8591
rect 9068 8584 9092 8591
rect 9148 8584 9172 8591
rect 8532 8576 9228 8584
rect 8532 8554 8534 8576
rect 8586 8554 8598 8576
rect 8650 8554 8662 8576
rect 8714 8554 8726 8576
rect 8778 8554 8790 8576
rect 8842 8554 8854 8576
rect 8906 8554 8918 8576
rect 8970 8554 8982 8576
rect 9034 8554 9046 8576
rect 9098 8554 9110 8576
rect 9162 8554 9174 8576
rect 9226 8554 9228 8576
rect 8588 8524 8598 8554
rect 8842 8524 8852 8554
rect 8908 8524 8918 8554
rect 9162 8524 9172 8554
rect 376 8498 379 8509
rect 367 8468 379 8498
rect 376 8457 379 8468
rect 315 8442 320 8457
rect 376 8442 431 8457
rect 376 8412 379 8442
rect 367 8390 379 8412
rect 8588 8509 8612 8524
rect 8668 8509 8692 8524
rect 8748 8509 8772 8524
rect 8828 8509 8852 8524
rect 8908 8509 8932 8524
rect 8988 8509 9012 8524
rect 9068 8509 9092 8524
rect 9148 8509 9172 8524
rect 8588 8498 8598 8509
rect 8842 8498 8852 8509
rect 8908 8498 8918 8509
rect 9162 8498 9172 8509
rect 8532 8468 8534 8498
rect 8586 8468 8598 8498
rect 8650 8468 8662 8498
rect 8714 8468 8726 8498
rect 8778 8468 8790 8498
rect 8842 8468 8854 8498
rect 8906 8468 8918 8498
rect 8970 8468 8982 8498
rect 9034 8468 9046 8498
rect 9098 8468 9110 8498
rect 9162 8468 9174 8498
rect 9226 8468 9228 8498
rect 8588 8457 8598 8468
rect 8842 8457 8852 8468
rect 8908 8457 8918 8468
rect 9162 8457 9172 8468
rect 8588 8442 8612 8457
rect 8668 8442 8692 8457
rect 8748 8442 8772 8457
rect 8828 8442 8852 8457
rect 8908 8442 8932 8457
rect 8988 8442 9012 8457
rect 9068 8442 9092 8457
rect 9148 8442 9172 8457
rect 315 8382 431 8390
rect 315 8375 320 8382
rect 376 8375 431 8382
rect 376 8326 379 8375
rect 367 8323 379 8326
rect 315 8317 431 8323
rect 7044 8429 7843 8436
rect 7096 8377 7160 8429
rect 7212 8380 7843 8429
rect 7899 8380 7949 8436
rect 8005 8380 8054 8436
rect 8110 8380 8159 8436
rect 8215 8380 8264 8436
rect 8320 8380 8369 8436
rect 8425 8380 8434 8436
rect 7212 8377 8434 8380
rect 7044 8362 8434 8377
rect 7096 8310 7160 8362
rect 7212 8310 8434 8362
rect 8588 8412 8598 8442
rect 8842 8412 8852 8442
rect 8908 8412 8918 8442
rect 9162 8412 9172 8442
rect 8532 8390 8534 8412
rect 8586 8390 8598 8412
rect 8650 8390 8662 8412
rect 8714 8390 8726 8412
rect 8778 8390 8790 8412
rect 8842 8390 8854 8412
rect 8906 8390 8918 8412
rect 8970 8390 8982 8412
rect 9034 8390 9046 8412
rect 9098 8390 9110 8412
rect 9162 8390 9174 8412
rect 9226 8390 9228 8412
rect 8532 8382 9228 8390
rect 8588 8375 8612 8382
rect 8668 8375 8692 8382
rect 8748 8375 8772 8382
rect 8828 8375 8852 8382
rect 8908 8375 8932 8382
rect 8988 8375 9012 8382
rect 9068 8375 9092 8382
rect 9148 8375 9172 8382
rect 8588 8326 8598 8375
rect 8842 8326 8852 8375
rect 8908 8326 8918 8375
rect 9162 8326 9172 8375
rect 8532 8323 8534 8326
rect 8586 8323 8598 8326
rect 8650 8323 8662 8326
rect 8714 8323 8726 8326
rect 8778 8323 8790 8326
rect 8842 8323 8854 8326
rect 8906 8323 8918 8326
rect 8970 8323 8982 8326
rect 9034 8323 9046 8326
rect 9098 8323 9110 8326
rect 9162 8323 9174 8326
rect 9226 8323 9228 8326
rect 8532 8317 9228 8323
rect 7044 8294 8434 8310
rect 7096 8242 7160 8294
rect 7212 8292 8434 8294
rect 7212 8242 7843 8292
rect 7044 8236 7843 8242
rect 7899 8236 7949 8292
rect 8005 8236 8054 8292
rect 8110 8236 8159 8292
rect 8215 8236 8264 8292
rect 8320 8236 8369 8292
rect 8425 8236 8434 8292
rect 4416 7950 4422 8002
rect 4481 7950 4490 8002
rect 4542 7950 4551 8002
rect 4610 7950 4616 8002
rect 4416 7946 4425 7950
rect 4481 7946 4551 7950
rect 4607 7946 4616 7950
rect 4416 7922 4616 7946
rect 4416 7918 4425 7922
rect 4481 7918 4551 7922
rect 4607 7918 4616 7922
rect 4416 7866 4422 7918
rect 4481 7866 4490 7918
rect 4542 7866 4551 7918
rect 4610 7866 4616 7918
rect 954 7754 963 7810
rect 1019 7754 1069 7810
rect 1125 7754 1174 7810
rect 1230 7754 1279 7810
rect 1335 7754 1384 7810
rect 1440 7754 1489 7810
rect 1545 7804 4077 7810
rect 1545 7754 3877 7804
rect 954 7752 3877 7754
rect 3929 7752 3951 7804
rect 4003 7752 4025 7804
rect 954 7736 4077 7752
rect 954 7684 3877 7736
rect 3929 7684 3951 7736
rect 4003 7684 4025 7736
rect 954 7668 4077 7684
rect 954 7666 3877 7668
rect 954 7610 963 7666
rect 1019 7610 1069 7666
rect 1125 7610 1174 7666
rect 1230 7610 1279 7666
rect 1335 7610 1384 7666
rect 1440 7610 1489 7666
rect 1545 7616 3877 7666
rect 3929 7616 3951 7668
rect 4003 7616 4025 7668
rect 1545 7610 4077 7616
tri 4902 7610 4904 7612 se
tri 4870 7578 4902 7610 se
rect 4902 7578 4904 7610
rect 1144 7572 4910 7578
rect 1196 7526 4910 7572
rect 1144 7508 1196 7520
tri 1196 7492 1230 7526 nw
rect 1144 7450 1196 7456
rect 2656 7191 2708 7197
rect 2656 7127 2708 7139
tri 2708 7119 2742 7153 sw
tri 3320 7119 3354 7153 se
rect 2708 7075 3354 7119
rect 2656 7069 3354 7075
rect 2083 6875 2089 6927
rect 2141 6875 2173 6927
rect 2225 6875 2257 6927
rect 2309 6875 2341 6927
rect 2393 6875 2425 6927
rect 2477 6875 2882 6927
rect 2934 6875 2995 6927
rect 3047 6875 3107 6927
rect 3159 6875 3165 6927
rect 2083 6837 3165 6875
rect 2083 6785 2089 6837
rect 2141 6785 2173 6837
rect 2225 6785 2257 6837
rect 2309 6785 2341 6837
rect 2393 6785 2425 6837
rect 2477 6785 2882 6837
rect 2934 6785 2995 6837
rect 3047 6785 3107 6837
rect 3159 6785 3165 6837
rect 4416 6828 4422 6880
rect 4481 6828 4490 6880
rect 4542 6828 4551 6880
rect 4610 6828 4616 6880
rect 4416 6824 4425 6828
rect 4481 6824 4551 6828
rect 4607 6824 4616 6828
rect 4416 6800 4616 6824
rect 4416 6796 4425 6800
rect 4481 6796 4551 6800
rect 4607 6796 4616 6800
rect 1228 6750 1280 6756
rect 4416 6744 4422 6796
rect 4481 6744 4490 6796
rect 4542 6744 4551 6796
rect 4610 6744 4616 6796
rect 1228 6697 1280 6698
tri 1280 6697 1297 6714 sw
rect 7044 6697 7843 6704
rect 1228 6686 1297 6697
rect 1280 6680 1297 6686
tri 1297 6680 1314 6697 sw
rect 1280 6634 3558 6680
rect 1228 6628 3558 6634
rect 7096 6645 7160 6697
rect 7212 6648 7843 6697
rect 7899 6648 7949 6704
rect 8005 6648 8054 6704
rect 8110 6648 8159 6704
rect 8215 6648 8264 6704
rect 8320 6648 8369 6704
rect 8425 6648 8434 6704
rect 7212 6645 8434 6648
rect 7044 6630 8434 6645
rect 7096 6578 7160 6630
rect 7212 6578 8434 6630
rect 7044 6562 8434 6578
rect 7096 6510 7160 6562
rect 7212 6560 8434 6562
rect 7212 6510 7843 6560
rect 7044 6504 7843 6510
rect 7899 6504 7949 6560
rect 8005 6504 8054 6560
rect 8110 6504 8159 6560
rect 8215 6504 8264 6560
rect 8320 6504 8369 6560
rect 8425 6504 8434 6560
rect 7044 5910 7843 5917
rect 7096 5858 7160 5910
rect 7212 5861 7843 5910
rect 7899 5861 7949 5917
rect 8005 5861 8054 5917
rect 8110 5861 8159 5917
rect 8215 5861 8264 5917
rect 8320 5861 8369 5917
rect 8425 5861 8434 5917
rect 7212 5858 8434 5861
rect 7044 5843 8434 5858
rect 7096 5791 7160 5843
rect 7212 5791 8434 5843
rect 7044 5775 8434 5791
rect 7096 5723 7160 5775
rect 7212 5773 8434 5775
rect 7212 5723 7843 5773
rect 7044 5717 7843 5723
rect 7899 5717 7949 5773
rect 8005 5717 8054 5773
rect 8110 5717 8159 5773
rect 8215 5717 8264 5773
rect 8320 5717 8369 5773
rect 8425 5717 8434 5773
rect 1816 5640 1868 5646
rect 1816 5576 1868 5588
tri 1868 5570 1902 5604 sw
rect 1868 5524 3550 5570
rect 1816 5518 3550 5524
rect 4416 5434 4422 5486
rect 4481 5434 4490 5486
rect 4542 5434 4551 5486
rect 4610 5434 4616 5486
rect 4416 5430 4425 5434
rect 4481 5430 4551 5434
rect 4607 5430 4616 5434
rect 2083 5361 2089 5413
rect 2141 5361 2173 5413
rect 2225 5361 2257 5413
rect 2309 5361 2341 5413
rect 2393 5361 2425 5413
rect 2477 5361 2882 5413
rect 2934 5361 2995 5413
rect 3047 5361 3107 5413
rect 3159 5361 3165 5413
rect 2083 5323 3165 5361
rect 4416 5406 4616 5430
rect 4416 5402 4425 5406
rect 4481 5402 4551 5406
rect 4607 5402 4616 5406
rect 4416 5350 4422 5402
rect 4481 5350 4490 5402
rect 4542 5350 4551 5402
rect 4610 5350 4616 5402
rect 2083 5271 2089 5323
rect 2141 5271 2173 5323
rect 2225 5271 2257 5323
rect 2309 5271 2341 5323
rect 2393 5271 2425 5323
rect 2477 5271 2882 5323
rect 2934 5271 2995 5323
rect 3047 5271 3107 5323
rect 3159 5271 3165 5323
rect 2152 5201 2204 5207
rect 2152 5137 2204 5149
tri 2204 5129 2238 5163 sw
rect 2204 5085 3354 5129
rect 2152 5079 3354 5085
tri 3320 5045 3354 5079 ne
rect 7044 4861 7843 4868
rect 7096 4809 7160 4861
rect 7212 4812 7843 4861
rect 7899 4812 7949 4868
rect 8005 4812 8054 4868
rect 8110 4812 8159 4868
rect 8215 4812 8264 4868
rect 8320 4812 8369 4868
rect 8425 4812 8434 4868
rect 7212 4809 8434 4812
rect 7044 4794 8434 4809
rect 7096 4742 7160 4794
rect 7212 4742 8434 4794
rect 7044 4726 8434 4742
rect 7096 4674 7160 4726
rect 7212 4724 8434 4726
rect 7212 4674 7843 4724
rect 7044 4668 7843 4674
rect 7899 4668 7949 4724
rect 8005 4668 8054 4724
rect 8110 4668 8159 4724
rect 8215 4668 8264 4724
rect 8320 4668 8369 4724
rect 8425 4668 8434 4724
rect 2404 4399 2456 4405
rect 2404 4335 2456 4347
tri 2456 4327 2490 4361 sw
tri 3320 4327 3354 4361 se
rect 2456 4283 3354 4327
rect 2404 4277 3354 4283
rect 412 4083 418 4135
rect 470 4083 525 4135
rect 577 4083 632 4135
rect 684 4083 739 4135
rect 791 4083 845 4135
rect 897 4083 951 4135
rect 1003 4083 2882 4135
rect 2934 4083 2995 4135
rect 3047 4083 3107 4135
rect 3159 4083 3165 4135
rect 412 4045 3165 4083
rect 412 3993 418 4045
rect 470 3993 525 4045
rect 577 3993 632 4045
rect 684 3993 739 4045
rect 791 3993 845 4045
rect 897 3993 951 4045
rect 1003 3993 2882 4045
rect 2934 3993 2995 4045
rect 3047 3993 3107 4045
rect 3159 3993 3165 4045
rect 4416 4006 4422 4058
rect 4481 4006 4490 4058
rect 4542 4006 4551 4058
rect 4610 4006 4616 4058
rect 4416 4002 4425 4006
rect 4481 4002 4551 4006
rect 4607 4002 4616 4006
rect 4416 3978 4616 4002
rect 4416 3974 4425 3978
rect 4481 3974 4551 3978
rect 4607 3974 4616 3978
rect 1396 3958 1448 3964
rect 4416 3922 4422 3974
rect 4481 3922 4490 3974
rect 4542 3922 4551 3974
rect 4610 3922 4616 3974
rect 1396 3894 1448 3906
tri 1448 3888 1482 3922 sw
rect 1448 3842 3553 3888
rect 1396 3836 3553 3842
rect 7044 3725 7843 3732
rect 7096 3673 7160 3725
rect 7212 3676 7843 3725
rect 7899 3676 7949 3732
rect 8005 3676 8054 3732
rect 8110 3676 8159 3732
rect 8215 3676 8264 3732
rect 8320 3676 8369 3732
rect 8425 3676 8434 3732
rect 7212 3673 8434 3676
rect 7044 3658 8434 3673
rect 7096 3606 7160 3658
rect 7212 3606 8434 3658
rect 7044 3590 8434 3606
rect 7096 3538 7160 3590
rect 7212 3588 8434 3590
rect 7212 3538 7843 3588
rect 7044 3532 7843 3538
rect 7899 3532 7949 3588
rect 8005 3532 8054 3588
rect 8110 3532 8159 3588
rect 8215 3532 8264 3588
rect 8320 3532 8369 3588
rect 8425 3532 8434 3588
rect 954 3261 963 3317
rect 1019 3261 1069 3317
rect 1125 3261 1174 3317
rect 1230 3261 1279 3317
rect 1335 3261 1384 3317
rect 1440 3261 1489 3317
rect 1545 3311 4077 3317
rect 1545 3261 2944 3311
rect 954 3259 2944 3261
rect 2996 3259 3877 3311
rect 3929 3259 3951 3311
rect 4003 3259 4025 3311
rect 954 3243 4077 3259
rect 954 3191 2944 3243
rect 2996 3191 3877 3243
rect 3929 3191 3951 3243
rect 4003 3191 4025 3243
rect 954 3175 4077 3191
rect 954 3173 2944 3175
rect 954 3117 963 3173
rect 1019 3117 1069 3173
rect 1125 3117 1174 3173
rect 1230 3117 1279 3173
rect 1335 3117 1384 3173
rect 1440 3117 1489 3173
rect 1545 3123 2944 3173
rect 2996 3123 3877 3175
rect 3929 3123 3951 3175
rect 4003 3123 4025 3175
rect 1545 3117 4077 3123
rect 4416 3316 4616 3322
rect 4468 3312 4490 3316
rect 4542 3312 4564 3316
rect 4416 3256 4452 3264
rect 4508 3256 4532 3264
rect 4588 3256 4616 3264
rect 4416 3231 4616 3256
rect 4416 3188 4452 3231
rect 4508 3188 4532 3231
rect 4588 3188 4616 3231
rect 4468 3150 4490 3175
rect 4542 3150 4564 3175
rect 4736 3281 4788 3287
rect 4736 3217 4788 3229
tri 4788 3215 4818 3245 sw
rect 7044 3215 7843 3222
rect 4788 3211 4818 3215
tri 4818 3211 4822 3215 sw
rect 4788 3208 6054 3211
tri 6054 3208 6057 3211 sw
rect 4788 3165 6057 3208
rect 4736 3163 6057 3165
tri 6057 3163 6102 3208 sw
rect 7096 3163 7160 3215
rect 7212 3166 7843 3215
rect 7899 3166 7949 3222
rect 8005 3166 8054 3222
rect 8110 3166 8159 3222
rect 8215 3166 8264 3222
rect 8320 3166 8369 3222
rect 8425 3166 8434 3222
rect 7212 3163 8434 3166
rect 4736 3159 6102 3163
tri 6102 3159 6106 3163 sw
tri 6032 3148 6043 3159 ne
rect 6043 3148 6106 3159
tri 6106 3148 6117 3159 sw
rect 7044 3148 8434 3163
rect 4416 3094 4452 3136
rect 4508 3094 4532 3136
rect 4588 3094 4616 3136
tri 6043 3134 6057 3148 ne
rect 6057 3134 6117 3148
tri 6117 3134 6131 3148 sw
tri 6057 3112 6079 3134 ne
rect 4416 3069 4616 3094
rect 4416 3060 4452 3069
rect 4508 3060 4532 3069
rect 4588 3060 4616 3069
rect 4468 3008 4490 3013
rect 4542 3008 4564 3013
rect 4416 2988 4616 3008
rect 4416 2932 4452 2988
rect 4508 2932 4532 2988
rect 4588 2932 4616 2988
rect 4468 2907 4490 2932
rect 4542 2907 4564 2932
rect 4656 3047 5964 3050
tri 5964 3047 5967 3050 sw
rect 4656 3044 5967 3047
rect 4708 3028 5967 3044
tri 5967 3028 5986 3047 sw
rect 4708 2998 5986 3028
rect 4708 2992 4732 2998
rect 4656 2988 4732 2992
tri 4732 2988 4742 2998 nw
tri 5942 2988 5952 2998 ne
rect 5952 2988 5986 2998
tri 5986 2988 6026 3028 sw
rect 6079 2988 6131 3134
rect 7096 3096 7160 3148
rect 7212 3096 8434 3148
rect 7044 3080 8434 3096
rect 7096 3028 7160 3080
rect 7212 3078 8434 3080
rect 7212 3028 7843 3078
rect 7044 3022 7843 3028
rect 7899 3022 7949 3078
rect 8005 3022 8054 3078
rect 8110 3022 8159 3078
rect 8215 3022 8264 3078
rect 8320 3022 8369 3078
rect 8425 3022 8434 3078
rect 4656 2980 4717 2988
rect 4708 2973 4717 2980
tri 4717 2973 4732 2988 nw
tri 5952 2973 5967 2988 ne
rect 5967 2973 6026 2988
tri 6026 2973 6041 2988 sw
tri 4708 2964 4717 2973 nw
tri 5967 2964 5976 2973 ne
rect 5976 2964 6041 2973
tri 5976 2951 5989 2964 ne
rect 4656 2922 4708 2928
rect 4416 2851 4452 2880
rect 4508 2851 4532 2880
rect 4588 2851 4616 2880
rect 4416 2826 4616 2851
rect 4416 2804 4452 2826
rect 4508 2804 4532 2826
rect 4588 2804 4616 2826
rect 4468 2752 4490 2770
rect 4542 2752 4564 2770
rect 4416 2744 4616 2752
rect 4416 2688 4452 2744
rect 4508 2688 4532 2744
rect 4588 2688 4616 2744
rect 5989 2827 6041 2964
rect 6079 2924 6131 2936
rect 6079 2866 6131 2872
rect 5989 2763 6041 2775
rect 5989 2705 6041 2711
rect 6278 2825 6330 2831
rect 6278 2761 6330 2773
rect 6278 2703 6330 2709
rect 7158 2825 7210 2831
rect 7158 2761 7210 2773
rect 4416 2676 4616 2688
rect 4468 2662 4490 2676
rect 4542 2662 4564 2676
rect 4416 2606 4452 2624
rect 4508 2606 4532 2624
rect 4588 2606 4616 2624
rect 4416 2580 4616 2606
rect 4416 2547 4452 2580
rect 4508 2547 4532 2580
rect 4588 2547 4616 2580
rect 4468 2498 4490 2524
rect 4542 2498 4564 2524
rect 4416 2442 4452 2495
rect 4508 2442 4532 2495
rect 4588 2442 4616 2495
rect 4416 2418 4616 2442
rect 4468 2416 4490 2418
rect 4542 2416 4564 2418
rect 4416 2360 4452 2366
rect 4508 2360 4532 2366
rect 4588 2360 4616 2366
rect 4416 2334 4616 2360
rect 4416 2278 4452 2334
rect 4508 2278 4532 2334
rect 4588 2278 4616 2334
rect 4416 2252 4616 2278
rect 4416 2196 4452 2252
rect 4508 2196 4532 2252
rect 4588 2196 4616 2252
rect 954 2133 963 2189
rect 1019 2133 1069 2189
rect 1125 2133 1174 2189
rect 1230 2133 1279 2189
rect 1335 2133 1384 2189
rect 1440 2133 1489 2189
rect 1545 2188 4077 2189
rect 1545 2136 3477 2188
rect 3529 2136 3586 2188
rect 3638 2136 3695 2188
rect 3747 2136 3803 2188
rect 3855 2136 3911 2188
rect 3963 2136 4019 2188
rect 4071 2136 4077 2188
rect 1545 2133 4077 2136
rect 954 2106 4077 2133
rect 954 2067 3477 2106
rect 954 2011 963 2067
rect 1019 2011 1069 2067
rect 1125 2011 1174 2067
rect 1230 2011 1279 2067
rect 1335 2011 1384 2067
rect 1440 2011 1489 2067
rect 1545 2054 3477 2067
rect 3529 2054 3586 2106
rect 3638 2054 3695 2106
rect 3747 2054 3803 2106
rect 3855 2054 3911 2106
rect 3963 2054 4019 2106
rect 4071 2054 4077 2106
rect 1545 2024 4077 2054
rect 1545 2011 3477 2024
rect 954 1972 3477 2011
rect 3529 1972 3586 2024
rect 3638 1972 3695 2024
rect 3747 1972 3803 2024
rect 3855 1972 3911 2024
rect 3963 1972 4019 2024
rect 4071 1972 4077 2024
rect 954 1945 4077 1972
rect 954 1889 963 1945
rect 1019 1889 1069 1945
rect 1125 1889 1174 1945
rect 1230 1889 1279 1945
rect 1335 1889 1384 1945
rect 1440 1889 1489 1945
rect 1545 1942 4077 1945
rect 1545 1890 3477 1942
rect 3529 1890 3586 1942
rect 3638 1890 3695 1942
rect 3747 1890 3803 1942
rect 3855 1890 3911 1942
rect 3963 1890 4019 1942
rect 4071 1890 4077 1942
rect 1545 1889 4077 1890
rect 4416 2170 4616 2196
rect 4416 2114 4452 2170
rect 4508 2114 4532 2170
rect 4588 2114 4616 2170
rect 4416 2088 4616 2114
rect 4416 2032 4452 2088
rect 4508 2032 4532 2088
rect 4588 2032 4616 2088
rect 4416 2006 4616 2032
rect 4416 1950 4452 2006
rect 4508 1950 4532 2006
rect 4588 1950 4616 2006
rect 4416 1924 4616 1950
rect 4416 1868 4452 1924
rect 4508 1868 4532 1924
rect 4588 1868 4616 1924
rect 4416 1842 4616 1868
rect 4416 1786 4452 1842
rect 4508 1786 4532 1842
rect 4588 1786 4616 1842
rect 4416 1777 4616 1786
rect 6278 2363 6330 2369
rect 6278 2299 6330 2311
rect 1312 122 1364 128
rect 1312 58 1364 70
rect 1312 0 1364 6
rect 1648 122 1700 128
rect 1648 58 1700 70
rect 1648 0 1700 6
rect 1900 122 1952 128
rect 1900 58 1952 70
rect 1900 0 1952 6
rect 2152 122 2204 128
rect 2152 58 2204 70
rect 2152 0 2204 6
rect 2404 122 2456 128
rect 2404 58 2456 70
rect 2404 0 2456 6
rect 2656 122 2708 128
rect 2656 58 2708 70
rect 2656 0 2708 6
rect 6278 122 6330 2247
rect 6278 58 6330 70
rect 6278 0 6330 6
rect 7158 122 7210 2709
rect 7158 58 7210 70
rect 7158 0 7210 6
<< via2 >>
rect 1949 39809 2005 39865
rect 2033 39809 2089 39865
rect 2117 39809 2173 39865
rect 2201 39809 2257 39865
rect 2285 39809 2341 39865
rect 2369 39809 2425 39865
rect 2453 39809 2509 39865
rect 2537 39809 2593 39865
rect 1949 39729 2005 39785
rect 2033 39729 2089 39785
rect 2117 39729 2173 39785
rect 2201 39729 2257 39785
rect 2285 39729 2341 39785
rect 2369 39729 2425 39785
rect 2453 39729 2509 39785
rect 2537 39729 2593 39785
rect 1949 39649 2005 39705
rect 2033 39649 2089 39705
rect 2117 39649 2173 39705
rect 2201 39649 2257 39705
rect 2285 39649 2341 39705
rect 2369 39649 2425 39705
rect 2453 39649 2509 39705
rect 2537 39649 2593 39705
rect 1949 39569 2005 39625
rect 2033 39569 2089 39625
rect 2117 39569 2173 39625
rect 2201 39569 2257 39625
rect 2285 39569 2341 39625
rect 2369 39569 2425 39625
rect 2453 39569 2509 39625
rect 2537 39569 2593 39625
rect 1949 39489 2005 39545
rect 2033 39489 2089 39545
rect 2117 39489 2173 39545
rect 2201 39489 2257 39545
rect 2285 39489 2341 39545
rect 2369 39489 2425 39545
rect 2453 39489 2509 39545
rect 2537 39489 2593 39545
rect 1949 39409 2005 39465
rect 2033 39409 2089 39465
rect 2117 39409 2173 39465
rect 2201 39409 2257 39465
rect 2285 39409 2341 39465
rect 2369 39409 2425 39465
rect 2453 39409 2509 39465
rect 2537 39409 2593 39465
rect 1949 39329 2005 39385
rect 2033 39329 2089 39385
rect 2117 39329 2173 39385
rect 2201 39329 2257 39385
rect 2285 39329 2341 39385
rect 2369 39329 2425 39385
rect 2453 39329 2509 39385
rect 2537 39329 2593 39385
rect 1949 39249 2005 39305
rect 2033 39249 2089 39305
rect 2117 39249 2173 39305
rect 2201 39249 2257 39305
rect 2285 39249 2341 39305
rect 2369 39249 2425 39305
rect 2453 39249 2509 39305
rect 2537 39249 2593 39305
rect 1949 39169 2005 39225
rect 2033 39169 2089 39225
rect 2117 39169 2173 39225
rect 2201 39169 2257 39225
rect 2285 39169 2341 39225
rect 2369 39169 2425 39225
rect 2453 39169 2509 39225
rect 2537 39169 2593 39225
rect 1949 39089 2005 39145
rect 2033 39089 2089 39145
rect 2117 39089 2173 39145
rect 2201 39089 2257 39145
rect 2285 39089 2341 39145
rect 2369 39089 2425 39145
rect 2453 39089 2509 39145
rect 2537 39089 2593 39145
rect 1949 39009 2005 39065
rect 2033 39009 2089 39065
rect 2117 39009 2173 39065
rect 2201 39009 2257 39065
rect 2285 39009 2341 39065
rect 2369 39009 2425 39065
rect 2453 39009 2509 39065
rect 2537 39009 2593 39065
rect 1949 38929 2005 38985
rect 2033 38929 2089 38985
rect 2117 38929 2173 38985
rect 2201 38929 2257 38985
rect 2285 38929 2341 38985
rect 2369 38929 2425 38985
rect 2453 38929 2509 38985
rect 2537 38929 2593 38985
rect 1949 38849 2005 38905
rect 2033 38849 2089 38905
rect 2117 38849 2173 38905
rect 2201 38849 2257 38905
rect 2285 38849 2341 38905
rect 2369 38849 2425 38905
rect 2453 38849 2509 38905
rect 2537 38849 2593 38905
rect 1949 38769 2005 38825
rect 2033 38769 2089 38825
rect 2117 38769 2173 38825
rect 2201 38769 2257 38825
rect 2285 38769 2341 38825
rect 2369 38769 2425 38825
rect 2453 38769 2509 38825
rect 2537 38769 2593 38825
rect 1949 38689 2005 38745
rect 2033 38689 2089 38745
rect 2117 38689 2173 38745
rect 2201 38689 2257 38745
rect 2285 38689 2341 38745
rect 2369 38689 2425 38745
rect 2453 38689 2509 38745
rect 2537 38689 2593 38745
rect 1949 38609 2005 38665
rect 2033 38609 2089 38665
rect 2117 38609 2173 38665
rect 2201 38609 2257 38665
rect 2285 38609 2341 38665
rect 2369 38609 2425 38665
rect 2453 38609 2509 38665
rect 2537 38609 2593 38665
rect 1949 38529 2005 38585
rect 2033 38529 2089 38585
rect 2117 38529 2173 38585
rect 2201 38529 2257 38585
rect 2285 38529 2341 38585
rect 2369 38529 2425 38585
rect 2453 38529 2509 38585
rect 2537 38529 2593 38585
rect 1949 38449 2005 38505
rect 2033 38449 2089 38505
rect 2117 38449 2173 38505
rect 2201 38449 2257 38505
rect 2285 38449 2341 38505
rect 2369 38449 2425 38505
rect 2453 38449 2509 38505
rect 2537 38449 2593 38505
rect 1949 38369 2005 38425
rect 2033 38369 2089 38425
rect 2117 38369 2173 38425
rect 2201 38369 2257 38425
rect 2285 38369 2341 38425
rect 2369 38369 2425 38425
rect 2453 38369 2509 38425
rect 2537 38369 2593 38425
rect 1949 38289 2005 38345
rect 2033 38289 2089 38345
rect 2117 38289 2173 38345
rect 2201 38289 2257 38345
rect 2285 38289 2341 38345
rect 2369 38289 2425 38345
rect 2453 38289 2509 38345
rect 2537 38289 2593 38345
rect 1949 38209 2005 38265
rect 2033 38209 2089 38265
rect 2117 38209 2173 38265
rect 2201 38209 2257 38265
rect 2285 38209 2341 38265
rect 2369 38209 2425 38265
rect 2453 38209 2509 38265
rect 2537 38209 2593 38265
rect 1949 38129 2005 38185
rect 2033 38129 2089 38185
rect 2117 38129 2173 38185
rect 2201 38129 2257 38185
rect 2285 38129 2341 38185
rect 2369 38129 2425 38185
rect 2453 38129 2509 38185
rect 2537 38129 2593 38185
rect 1949 38049 2005 38105
rect 2033 38049 2089 38105
rect 2117 38049 2173 38105
rect 2201 38049 2257 38105
rect 2285 38049 2341 38105
rect 2369 38049 2425 38105
rect 2453 38049 2509 38105
rect 2537 38049 2593 38105
rect 1949 37969 2005 38025
rect 2033 37969 2089 38025
rect 2117 37969 2173 38025
rect 2201 37969 2257 38025
rect 2285 37969 2341 38025
rect 2369 37969 2425 38025
rect 2453 37969 2509 38025
rect 2537 37969 2593 38025
rect 1949 37889 2005 37945
rect 2033 37889 2089 37945
rect 2117 37889 2173 37945
rect 2201 37889 2257 37945
rect 2285 37889 2341 37945
rect 2369 37889 2425 37945
rect 2453 37889 2509 37945
rect 2537 37889 2593 37945
rect 1949 37809 2005 37865
rect 2033 37809 2089 37865
rect 2117 37809 2173 37865
rect 2201 37809 2257 37865
rect 2285 37809 2341 37865
rect 2369 37809 2425 37865
rect 2453 37809 2509 37865
rect 2537 37809 2593 37865
rect 1949 37729 2005 37785
rect 2033 37729 2089 37785
rect 2117 37729 2173 37785
rect 2201 37729 2257 37785
rect 2285 37729 2341 37785
rect 2369 37729 2425 37785
rect 2453 37729 2509 37785
rect 2537 37729 2593 37785
rect 1949 37649 2005 37705
rect 2033 37649 2089 37705
rect 2117 37649 2173 37705
rect 2201 37649 2257 37705
rect 2285 37649 2341 37705
rect 2369 37649 2425 37705
rect 2453 37649 2509 37705
rect 2537 37649 2593 37705
rect 1949 37569 2005 37625
rect 2033 37569 2089 37625
rect 2117 37569 2173 37625
rect 2201 37569 2257 37625
rect 2285 37569 2341 37625
rect 2369 37569 2425 37625
rect 2453 37569 2509 37625
rect 2537 37569 2593 37625
rect 1949 37489 2005 37545
rect 2033 37489 2089 37545
rect 2117 37489 2173 37545
rect 2201 37489 2257 37545
rect 2285 37489 2341 37545
rect 2369 37489 2425 37545
rect 2453 37489 2509 37545
rect 2537 37489 2593 37545
rect 1949 37409 2005 37465
rect 2033 37409 2089 37465
rect 2117 37409 2173 37465
rect 2201 37409 2257 37465
rect 2285 37409 2341 37465
rect 2369 37409 2425 37465
rect 2453 37409 2509 37465
rect 2537 37409 2593 37465
rect 1949 37329 2005 37385
rect 2033 37329 2089 37385
rect 2117 37329 2173 37385
rect 2201 37329 2257 37385
rect 2285 37329 2341 37385
rect 2369 37329 2425 37385
rect 2453 37329 2509 37385
rect 2537 37329 2593 37385
rect 1949 37249 2005 37305
rect 2033 37249 2089 37305
rect 2117 37249 2173 37305
rect 2201 37249 2257 37305
rect 2285 37249 2341 37305
rect 2369 37249 2425 37305
rect 2453 37249 2509 37305
rect 2537 37249 2593 37305
rect 1949 37169 2005 37225
rect 2033 37169 2089 37225
rect 2117 37169 2173 37225
rect 2201 37169 2257 37225
rect 2285 37169 2341 37225
rect 2369 37169 2425 37225
rect 2453 37169 2509 37225
rect 2537 37169 2593 37225
rect 1949 37089 2005 37145
rect 2033 37089 2089 37145
rect 2117 37089 2173 37145
rect 2201 37089 2257 37145
rect 2285 37089 2341 37145
rect 2369 37089 2425 37145
rect 2453 37089 2509 37145
rect 2537 37089 2593 37145
rect 6903 39814 6959 39870
rect 6993 39814 7049 39870
rect 7083 39814 7139 39870
rect 7173 39814 7229 39870
rect 7263 39814 7319 39870
rect 7353 39814 7409 39870
rect 7443 39814 7499 39870
rect 6903 39734 6959 39790
rect 6993 39734 7049 39790
rect 7083 39734 7139 39790
rect 7173 39734 7229 39790
rect 7263 39734 7319 39790
rect 7353 39734 7409 39790
rect 7443 39734 7499 39790
rect 6903 39654 6959 39710
rect 6993 39654 7049 39710
rect 7083 39654 7139 39710
rect 7173 39654 7229 39710
rect 7263 39654 7319 39710
rect 7353 39654 7409 39710
rect 7443 39654 7499 39710
rect 6903 39574 6959 39630
rect 6993 39574 7049 39630
rect 7083 39574 7139 39630
rect 7173 39574 7229 39630
rect 7263 39574 7319 39630
rect 7353 39574 7409 39630
rect 7443 39574 7499 39630
rect 6903 39494 6959 39550
rect 6993 39494 7049 39550
rect 7083 39494 7139 39550
rect 7173 39494 7229 39550
rect 7263 39494 7319 39550
rect 7353 39494 7409 39550
rect 7443 39494 7499 39550
rect 6903 39414 6959 39470
rect 6993 39414 7049 39470
rect 7083 39414 7139 39470
rect 7173 39414 7229 39470
rect 7263 39414 7319 39470
rect 7353 39414 7409 39470
rect 7443 39414 7499 39470
rect 6903 39334 6959 39390
rect 6993 39334 7049 39390
rect 7083 39334 7139 39390
rect 7173 39334 7229 39390
rect 7263 39334 7319 39390
rect 7353 39334 7409 39390
rect 7443 39334 7499 39390
rect 6903 39254 6959 39310
rect 6993 39254 7049 39310
rect 7083 39254 7139 39310
rect 7173 39254 7229 39310
rect 7263 39254 7319 39310
rect 7353 39254 7409 39310
rect 7443 39254 7499 39310
rect 6903 39174 6959 39230
rect 6993 39174 7049 39230
rect 7083 39174 7139 39230
rect 7173 39174 7229 39230
rect 7263 39174 7319 39230
rect 7353 39174 7409 39230
rect 7443 39174 7499 39230
rect 6903 39094 6959 39150
rect 6993 39094 7049 39150
rect 7083 39094 7139 39150
rect 7173 39094 7229 39150
rect 7263 39094 7319 39150
rect 7353 39094 7409 39150
rect 7443 39094 7499 39150
rect 6903 39014 6959 39070
rect 6993 39014 7049 39070
rect 7083 39014 7139 39070
rect 7173 39014 7229 39070
rect 7263 39014 7319 39070
rect 7353 39014 7409 39070
rect 7443 39014 7499 39070
rect 6903 38934 6959 38990
rect 6993 38934 7049 38990
rect 7083 38934 7139 38990
rect 7173 38934 7229 38990
rect 7263 38934 7319 38990
rect 7353 38934 7409 38990
rect 7443 38934 7499 38990
rect 6903 38854 6959 38910
rect 6993 38854 7049 38910
rect 7083 38854 7139 38910
rect 7173 38854 7229 38910
rect 7263 38854 7319 38910
rect 7353 38854 7409 38910
rect 7443 38854 7499 38910
rect 6903 38774 6959 38830
rect 6993 38774 7049 38830
rect 7083 38774 7139 38830
rect 7173 38774 7229 38830
rect 7263 38774 7319 38830
rect 7353 38774 7409 38830
rect 7443 38774 7499 38830
rect 6903 38694 6959 38750
rect 6993 38694 7049 38750
rect 7083 38694 7139 38750
rect 7173 38694 7229 38750
rect 7263 38694 7319 38750
rect 7353 38694 7409 38750
rect 7443 38694 7499 38750
rect 6903 38614 6959 38670
rect 6993 38614 7049 38670
rect 7083 38614 7139 38670
rect 7173 38614 7229 38670
rect 7263 38614 7319 38670
rect 7353 38614 7409 38670
rect 7443 38614 7499 38670
rect 6903 38534 6959 38590
rect 6993 38534 7049 38590
rect 7083 38534 7139 38590
rect 7173 38534 7229 38590
rect 7263 38534 7319 38590
rect 7353 38534 7409 38590
rect 7443 38534 7499 38590
rect 6903 38454 6959 38510
rect 6993 38454 7049 38510
rect 7083 38454 7139 38510
rect 7173 38454 7229 38510
rect 7263 38454 7319 38510
rect 7353 38454 7409 38510
rect 7443 38454 7499 38510
rect 6903 38374 6959 38430
rect 6993 38374 7049 38430
rect 7083 38374 7139 38430
rect 7173 38374 7229 38430
rect 7263 38374 7319 38430
rect 7353 38374 7409 38430
rect 7443 38374 7499 38430
rect 6903 38294 6959 38350
rect 6993 38294 7049 38350
rect 7083 38294 7139 38350
rect 7173 38294 7229 38350
rect 7263 38294 7319 38350
rect 7353 38294 7409 38350
rect 7443 38294 7499 38350
rect 6903 38214 6959 38270
rect 6993 38214 7049 38270
rect 7083 38214 7139 38270
rect 7173 38214 7229 38270
rect 7263 38214 7319 38270
rect 7353 38214 7409 38270
rect 7443 38214 7499 38270
rect 6903 38134 6959 38190
rect 6993 38134 7049 38190
rect 7083 38134 7139 38190
rect 7173 38134 7229 38190
rect 7263 38134 7319 38190
rect 7353 38134 7409 38190
rect 7443 38134 7499 38190
rect 6903 38054 6959 38110
rect 6993 38054 7049 38110
rect 7083 38054 7139 38110
rect 7173 38054 7229 38110
rect 7263 38054 7319 38110
rect 7353 38054 7409 38110
rect 7443 38054 7499 38110
rect 6903 37974 6959 38030
rect 6993 37974 7049 38030
rect 7083 37974 7139 38030
rect 7173 37974 7229 38030
rect 7263 37974 7319 38030
rect 7353 37974 7409 38030
rect 7443 37974 7499 38030
rect 6903 37894 6959 37950
rect 6993 37894 7049 37950
rect 7083 37894 7139 37950
rect 7173 37894 7229 37950
rect 7263 37894 7319 37950
rect 7353 37894 7409 37950
rect 7443 37894 7499 37950
rect 6903 37814 6959 37870
rect 6993 37814 7049 37870
rect 7083 37814 7139 37870
rect 7173 37814 7229 37870
rect 7263 37814 7319 37870
rect 7353 37814 7409 37870
rect 7443 37814 7499 37870
rect 6903 37734 6959 37790
rect 6993 37734 7049 37790
rect 7083 37734 7139 37790
rect 7173 37734 7229 37790
rect 7263 37734 7319 37790
rect 7353 37734 7409 37790
rect 7443 37734 7499 37790
rect 6903 37654 6959 37710
rect 6993 37654 7049 37710
rect 7083 37654 7139 37710
rect 7173 37654 7229 37710
rect 7263 37654 7319 37710
rect 7353 37654 7409 37710
rect 7443 37654 7499 37710
rect 6903 37574 6959 37630
rect 6993 37574 7049 37630
rect 7083 37574 7139 37630
rect 7173 37574 7229 37630
rect 7263 37574 7319 37630
rect 7353 37574 7409 37630
rect 7443 37574 7499 37630
rect 6903 37494 6959 37550
rect 6993 37494 7049 37550
rect 7083 37494 7139 37550
rect 7173 37494 7229 37550
rect 7263 37494 7319 37550
rect 7353 37494 7409 37550
rect 7443 37494 7499 37550
rect 6903 37414 6959 37470
rect 6993 37414 7049 37470
rect 7083 37414 7139 37470
rect 7173 37414 7229 37470
rect 7263 37414 7319 37470
rect 7353 37414 7409 37470
rect 7443 37414 7499 37470
rect 6903 37334 6959 37390
rect 6993 37334 7049 37390
rect 7083 37334 7139 37390
rect 7173 37334 7229 37390
rect 7263 37334 7319 37390
rect 7353 37334 7409 37390
rect 7443 37334 7499 37390
rect 6903 37254 6959 37310
rect 6993 37254 7049 37310
rect 7083 37254 7139 37310
rect 7173 37254 7229 37310
rect 7263 37254 7319 37310
rect 7353 37254 7409 37310
rect 7443 37254 7499 37310
rect 6903 37174 6959 37230
rect 6993 37174 7049 37230
rect 7083 37174 7139 37230
rect 7173 37174 7229 37230
rect 7263 37174 7319 37230
rect 7353 37174 7409 37230
rect 7443 37174 7499 37230
rect 1949 37009 2005 37065
rect 2033 37009 2089 37065
rect 2117 37009 2173 37065
rect 2201 37009 2257 37065
rect 2285 37009 2341 37065
rect 2369 37009 2425 37065
rect 2453 37009 2509 37065
rect 2537 37009 2593 37065
rect 1949 36929 2005 36985
rect 2033 36929 2089 36985
rect 2117 36929 2173 36985
rect 2201 36929 2257 36985
rect 2285 36929 2341 36985
rect 2369 36929 2425 36985
rect 2453 36929 2509 36985
rect 2537 36929 2593 36985
rect 1949 36849 2005 36905
rect 2033 36849 2089 36905
rect 2117 36849 2173 36905
rect 2201 36849 2257 36905
rect 2285 36849 2341 36905
rect 2369 36849 2425 36905
rect 2453 36849 2509 36905
rect 2537 36849 2593 36905
rect 1949 36769 2005 36825
rect 2033 36769 2089 36825
rect 2117 36769 2173 36825
rect 2201 36769 2257 36825
rect 2285 36769 2341 36825
rect 2369 36769 2425 36825
rect 2453 36769 2509 36825
rect 2537 36769 2593 36825
rect 1949 36689 2005 36745
rect 2033 36689 2089 36745
rect 2117 36689 2173 36745
rect 2201 36689 2257 36745
rect 2285 36689 2341 36745
rect 2369 36689 2425 36745
rect 2453 36689 2509 36745
rect 2537 36689 2593 36745
rect 1949 36609 2005 36665
rect 2033 36609 2089 36665
rect 2117 36609 2173 36665
rect 2201 36609 2257 36665
rect 2285 36609 2341 36665
rect 2369 36609 2425 36665
rect 2453 36609 2509 36665
rect 2537 36609 2593 36665
rect 1949 36529 2005 36585
rect 2033 36529 2089 36585
rect 2117 36529 2173 36585
rect 2201 36529 2257 36585
rect 2285 36529 2341 36585
rect 2369 36529 2425 36585
rect 2453 36529 2509 36585
rect 2537 36529 2593 36585
rect 1949 36449 2005 36505
rect 2033 36449 2089 36505
rect 2117 36449 2173 36505
rect 2201 36449 2257 36505
rect 2285 36449 2341 36505
rect 2369 36449 2425 36505
rect 2453 36449 2509 36505
rect 2537 36449 2593 36505
rect 1949 36369 2005 36425
rect 2033 36369 2089 36425
rect 2117 36369 2173 36425
rect 2201 36369 2257 36425
rect 2285 36369 2341 36425
rect 2369 36369 2425 36425
rect 2453 36369 2509 36425
rect 2537 36369 2593 36425
rect 1949 36289 2005 36345
rect 2033 36289 2089 36345
rect 2117 36289 2173 36345
rect 2201 36289 2257 36345
rect 2285 36289 2341 36345
rect 2369 36289 2425 36345
rect 2453 36289 2509 36345
rect 2537 36289 2593 36345
rect 1949 36209 2005 36265
rect 2033 36209 2089 36265
rect 2117 36209 2173 36265
rect 2201 36209 2257 36265
rect 2285 36209 2341 36265
rect 2369 36209 2425 36265
rect 2453 36209 2509 36265
rect 2537 36209 2593 36265
rect 1949 36129 2005 36185
rect 2033 36129 2089 36185
rect 2117 36129 2173 36185
rect 2201 36129 2257 36185
rect 2285 36129 2341 36185
rect 2369 36129 2425 36185
rect 2453 36129 2509 36185
rect 2537 36129 2593 36185
rect 1949 36049 2005 36105
rect 2033 36049 2089 36105
rect 2117 36049 2173 36105
rect 2201 36049 2257 36105
rect 2285 36049 2341 36105
rect 2369 36049 2425 36105
rect 2453 36049 2509 36105
rect 2537 36049 2593 36105
rect 1949 35969 2005 36025
rect 2033 35969 2089 36025
rect 2117 35969 2173 36025
rect 2201 35969 2257 36025
rect 2285 35969 2341 36025
rect 2369 35969 2425 36025
rect 2453 35969 2509 36025
rect 2537 35969 2593 36025
rect 1949 35889 2005 35945
rect 2033 35889 2089 35945
rect 2117 35889 2173 35945
rect 2201 35889 2257 35945
rect 2285 35889 2341 35945
rect 2369 35889 2425 35945
rect 2453 35889 2509 35945
rect 2537 35889 2593 35945
rect 1949 35809 2005 35865
rect 2033 35809 2089 35865
rect 2117 35809 2173 35865
rect 2201 35809 2257 35865
rect 2285 35809 2341 35865
rect 2369 35809 2425 35865
rect 2453 35809 2509 35865
rect 2537 35809 2593 35865
rect 1949 35729 2005 35785
rect 2033 35729 2089 35785
rect 2117 35729 2173 35785
rect 2201 35729 2257 35785
rect 2285 35729 2341 35785
rect 2369 35729 2425 35785
rect 2453 35729 2509 35785
rect 2537 35729 2593 35785
rect 1949 35649 2005 35705
rect 2033 35649 2089 35705
rect 2117 35649 2173 35705
rect 2201 35649 2257 35705
rect 2285 35649 2341 35705
rect 2369 35649 2425 35705
rect 2453 35649 2509 35705
rect 2537 35649 2593 35705
rect 1949 35569 2005 35625
rect 2033 35569 2089 35625
rect 2117 35569 2173 35625
rect 2201 35569 2257 35625
rect 2285 35569 2341 35625
rect 2369 35569 2425 35625
rect 2453 35569 2509 35625
rect 2537 35569 2593 35625
rect 1949 35489 2005 35545
rect 2033 35489 2089 35545
rect 2117 35489 2173 35545
rect 2201 35489 2257 35545
rect 2285 35489 2341 35545
rect 2369 35489 2425 35545
rect 2453 35489 2509 35545
rect 2537 35489 2593 35545
rect 1949 35409 2005 35465
rect 2033 35409 2089 35465
rect 2117 35409 2173 35465
rect 2201 35409 2257 35465
rect 2285 35409 2341 35465
rect 2369 35409 2425 35465
rect 2453 35409 2509 35465
rect 2537 35409 2593 35465
rect 1949 35329 2005 35385
rect 2033 35329 2089 35385
rect 2117 35329 2173 35385
rect 2201 35329 2257 35385
rect 2285 35329 2341 35385
rect 2369 35329 2425 35385
rect 2453 35329 2509 35385
rect 2537 35329 2593 35385
rect 1949 35249 2005 35305
rect 2033 35249 2089 35305
rect 2117 35249 2173 35305
rect 2201 35249 2257 35305
rect 2285 35249 2341 35305
rect 2369 35249 2425 35305
rect 2453 35249 2509 35305
rect 2537 35249 2593 35305
rect 1949 35169 2005 35225
rect 2033 35169 2089 35225
rect 2117 35169 2173 35225
rect 2201 35169 2257 35225
rect 2285 35169 2341 35225
rect 2369 35169 2425 35225
rect 2453 35169 2509 35225
rect 2537 35169 2593 35225
rect 1949 35089 2005 35145
rect 2033 35089 2089 35145
rect 2117 35089 2173 35145
rect 2201 35089 2257 35145
rect 2285 35089 2341 35145
rect 2369 35089 2425 35145
rect 2453 35089 2509 35145
rect 2537 35089 2593 35145
rect 1949 35009 2005 35065
rect 2033 35009 2089 35065
rect 2117 35009 2173 35065
rect 2201 35009 2257 35065
rect 2285 35009 2341 35065
rect 2369 35009 2425 35065
rect 2453 35009 2509 35065
rect 2537 35009 2593 35065
rect 1949 34929 2005 34985
rect 2033 34929 2089 34985
rect 2117 34929 2173 34985
rect 2201 34929 2257 34985
rect 2285 34929 2341 34985
rect 2369 34929 2425 34985
rect 2453 34929 2509 34985
rect 2537 34929 2593 34985
rect 1949 34849 2005 34905
rect 2033 34849 2089 34905
rect 2117 34849 2173 34905
rect 2201 34849 2257 34905
rect 2285 34849 2341 34905
rect 2369 34849 2425 34905
rect 2453 34849 2509 34905
rect 2537 34849 2593 34905
rect 1949 34769 2005 34825
rect 2033 34769 2089 34825
rect 2117 34769 2173 34825
rect 2201 34769 2257 34825
rect 2285 34769 2341 34825
rect 2369 34769 2425 34825
rect 2453 34769 2509 34825
rect 2537 34769 2593 34825
rect 1949 34689 2005 34745
rect 2033 34689 2089 34745
rect 2117 34689 2173 34745
rect 2201 34689 2257 34745
rect 2285 34689 2341 34745
rect 2369 34689 2425 34745
rect 2453 34689 2509 34745
rect 2537 34689 2593 34745
rect 1949 34609 2005 34665
rect 2033 34609 2089 34665
rect 2117 34609 2173 34665
rect 2201 34609 2257 34665
rect 2285 34609 2341 34665
rect 2369 34609 2425 34665
rect 2453 34609 2509 34665
rect 2537 34609 2593 34665
rect 1949 34529 2005 34585
rect 2033 34529 2089 34585
rect 2117 34529 2173 34585
rect 2201 34529 2257 34585
rect 2285 34529 2341 34585
rect 2369 34529 2425 34585
rect 2453 34529 2509 34585
rect 2537 34529 2593 34585
rect 1949 34449 2005 34505
rect 2033 34449 2089 34505
rect 2117 34449 2173 34505
rect 2201 34449 2257 34505
rect 2285 34449 2341 34505
rect 2369 34449 2425 34505
rect 2453 34449 2509 34505
rect 2537 34449 2593 34505
rect 1949 34369 2005 34425
rect 2033 34369 2089 34425
rect 2117 34369 2173 34425
rect 2201 34369 2257 34425
rect 2285 34369 2341 34425
rect 2369 34369 2425 34425
rect 2453 34369 2509 34425
rect 2537 34369 2593 34425
rect 1949 34289 2005 34345
rect 2033 34289 2089 34345
rect 2117 34289 2173 34345
rect 2201 34289 2257 34345
rect 2285 34289 2341 34345
rect 2369 34289 2425 34345
rect 2453 34289 2509 34345
rect 2537 34289 2593 34345
rect 1949 34209 2005 34265
rect 2033 34209 2089 34265
rect 2117 34209 2173 34265
rect 2201 34209 2257 34265
rect 2285 34209 2341 34265
rect 2369 34209 2425 34265
rect 2453 34209 2509 34265
rect 2537 34209 2593 34265
rect 1949 34129 2005 34185
rect 2033 34129 2089 34185
rect 2117 34129 2173 34185
rect 2201 34129 2257 34185
rect 2285 34129 2341 34185
rect 2369 34129 2425 34185
rect 2453 34129 2509 34185
rect 2537 34129 2593 34185
rect 1949 34049 2005 34105
rect 2033 34049 2089 34105
rect 2117 34049 2173 34105
rect 2201 34049 2257 34105
rect 2285 34049 2341 34105
rect 2369 34049 2425 34105
rect 2453 34049 2509 34105
rect 2537 34049 2593 34105
rect 1949 33969 2005 34025
rect 2033 33969 2089 34025
rect 2117 33969 2173 34025
rect 2201 33969 2257 34025
rect 2285 33969 2341 34025
rect 2369 33969 2425 34025
rect 2453 33969 2509 34025
rect 2537 33969 2593 34025
rect 1949 33889 2005 33945
rect 2033 33889 2089 33945
rect 2117 33889 2173 33945
rect 2201 33889 2257 33945
rect 2285 33889 2341 33945
rect 2369 33889 2425 33945
rect 2453 33889 2509 33945
rect 2537 33889 2593 33945
rect 1949 33809 2005 33865
rect 2033 33809 2089 33865
rect 2117 33809 2173 33865
rect 2201 33809 2257 33865
rect 2285 33809 2341 33865
rect 2369 33809 2425 33865
rect 2453 33809 2509 33865
rect 2537 33809 2593 33865
rect 1949 33729 2005 33785
rect 2033 33729 2089 33785
rect 2117 33729 2173 33785
rect 2201 33729 2257 33785
rect 2285 33729 2341 33785
rect 2369 33729 2425 33785
rect 2453 33729 2509 33785
rect 2537 33729 2593 33785
rect 1949 33649 2005 33705
rect 2033 33649 2089 33705
rect 2117 33649 2173 33705
rect 2201 33649 2257 33705
rect 2285 33649 2341 33705
rect 2369 33649 2425 33705
rect 2453 33649 2509 33705
rect 2537 33649 2593 33705
rect 1949 33569 2005 33625
rect 2033 33569 2089 33625
rect 2117 33569 2173 33625
rect 2201 33569 2257 33625
rect 2285 33569 2341 33625
rect 2369 33569 2425 33625
rect 2453 33569 2509 33625
rect 2537 33569 2593 33625
rect 1949 33489 2005 33545
rect 2033 33489 2089 33545
rect 2117 33489 2173 33545
rect 2201 33489 2257 33545
rect 2285 33489 2341 33545
rect 2369 33489 2425 33545
rect 2453 33489 2509 33545
rect 2537 33489 2593 33545
rect 1949 33409 2005 33465
rect 2033 33409 2089 33465
rect 2117 33409 2173 33465
rect 2201 33409 2257 33465
rect 2285 33409 2341 33465
rect 2369 33409 2425 33465
rect 2453 33409 2509 33465
rect 2537 33409 2593 33465
rect 1949 33329 2005 33385
rect 2033 33329 2089 33385
rect 2117 33329 2173 33385
rect 2201 33329 2257 33385
rect 2285 33329 2341 33385
rect 2369 33329 2425 33385
rect 2453 33329 2509 33385
rect 2537 33329 2593 33385
rect 1949 33249 2005 33305
rect 2033 33249 2089 33305
rect 2117 33249 2173 33305
rect 2201 33249 2257 33305
rect 2285 33249 2341 33305
rect 2369 33249 2425 33305
rect 2453 33249 2509 33305
rect 2537 33249 2593 33305
rect 1949 33169 2005 33225
rect 2033 33169 2089 33225
rect 2117 33169 2173 33225
rect 2201 33169 2257 33225
rect 2285 33169 2341 33225
rect 2369 33169 2425 33225
rect 2453 33169 2509 33225
rect 2537 33169 2593 33225
rect 1949 33089 2005 33145
rect 2033 33089 2089 33145
rect 2117 33089 2173 33145
rect 2201 33089 2257 33145
rect 2285 33089 2341 33145
rect 2369 33089 2425 33145
rect 2453 33089 2509 33145
rect 2537 33089 2593 33145
rect 1949 33009 2005 33065
rect 2033 33009 2089 33065
rect 2117 33009 2173 33065
rect 2201 33009 2257 33065
rect 2285 33009 2341 33065
rect 2369 33009 2425 33065
rect 2453 33009 2509 33065
rect 2537 33009 2593 33065
rect 1949 32929 2005 32985
rect 2033 32929 2089 32985
rect 2117 32929 2173 32985
rect 2201 32929 2257 32985
rect 2285 32929 2341 32985
rect 2369 32929 2425 32985
rect 2453 32929 2509 32985
rect 2537 32929 2593 32985
rect 1949 32849 2005 32905
rect 2033 32849 2089 32905
rect 2117 32849 2173 32905
rect 2201 32849 2257 32905
rect 2285 32849 2341 32905
rect 2369 32849 2425 32905
rect 2453 32849 2509 32905
rect 2537 32849 2593 32905
rect 1949 32769 2005 32825
rect 2033 32769 2089 32825
rect 2117 32769 2173 32825
rect 2201 32769 2257 32825
rect 2285 32769 2341 32825
rect 2369 32769 2425 32825
rect 2453 32769 2509 32825
rect 2537 32769 2593 32825
rect 1949 32689 2005 32745
rect 2033 32689 2089 32745
rect 2117 32689 2173 32745
rect 2201 32689 2257 32745
rect 2285 32689 2341 32745
rect 2369 32689 2425 32745
rect 2453 32689 2509 32745
rect 2537 32689 2593 32745
rect 1949 32608 2005 32664
rect 2033 32608 2089 32664
rect 2117 32608 2173 32664
rect 2201 32608 2257 32664
rect 2285 32608 2341 32664
rect 2369 32608 2425 32664
rect 2453 32608 2509 32664
rect 2537 32608 2593 32664
rect 1949 32527 2005 32583
rect 2033 32527 2089 32583
rect 2117 32527 2173 32583
rect 2201 32527 2257 32583
rect 2285 32527 2341 32583
rect 2369 32527 2425 32583
rect 2453 32527 2509 32583
rect 2537 32527 2593 32583
rect 1949 32446 2005 32502
rect 2033 32446 2089 32502
rect 2117 32446 2173 32502
rect 2201 32446 2257 32502
rect 2285 32446 2341 32502
rect 2369 32446 2425 32502
rect 2453 32446 2509 32502
rect 2537 32446 2593 32502
rect 1949 32365 2005 32421
rect 2033 32365 2089 32421
rect 2117 32365 2173 32421
rect 2201 32365 2257 32421
rect 2285 32365 2341 32421
rect 2369 32365 2425 32421
rect 2453 32365 2509 32421
rect 2537 32365 2593 32421
rect 1949 32284 2005 32340
rect 2033 32284 2089 32340
rect 2117 32284 2173 32340
rect 2201 32284 2257 32340
rect 2285 32284 2341 32340
rect 2369 32284 2425 32340
rect 2453 32284 2509 32340
rect 2537 32284 2593 32340
rect 1949 32203 2005 32259
rect 2033 32203 2089 32259
rect 2117 32203 2173 32259
rect 2201 32203 2257 32259
rect 2285 32203 2341 32259
rect 2369 32203 2425 32259
rect 2453 32203 2509 32259
rect 2537 32203 2593 32259
rect 1949 32122 2005 32178
rect 2033 32122 2089 32178
rect 2117 32122 2173 32178
rect 2201 32122 2257 32178
rect 2285 32122 2341 32178
rect 2369 32122 2425 32178
rect 2453 32122 2509 32178
rect 2537 32122 2593 32178
rect 1949 32041 2005 32097
rect 2033 32041 2089 32097
rect 2117 32041 2173 32097
rect 2201 32041 2257 32097
rect 2285 32041 2341 32097
rect 2369 32041 2425 32097
rect 2453 32041 2509 32097
rect 2537 32041 2593 32097
rect 1949 31960 2005 32016
rect 2033 31960 2089 32016
rect 2117 31960 2173 32016
rect 2201 31960 2257 32016
rect 2285 31960 2341 32016
rect 2369 31960 2425 32016
rect 2453 31960 2509 32016
rect 2537 31960 2593 32016
rect 1949 31879 2005 31935
rect 2033 31879 2089 31935
rect 2117 31879 2173 31935
rect 2201 31879 2257 31935
rect 2285 31879 2341 31935
rect 2369 31879 2425 31935
rect 2453 31879 2509 31935
rect 2537 31879 2593 31935
rect 1949 31798 2005 31854
rect 2033 31798 2089 31854
rect 2117 31798 2173 31854
rect 2201 31798 2257 31854
rect 2285 31798 2341 31854
rect 2369 31798 2425 31854
rect 2453 31798 2509 31854
rect 2537 31798 2593 31854
rect 1949 31717 2005 31773
rect 2033 31717 2089 31773
rect 2117 31717 2173 31773
rect 2201 31717 2257 31773
rect 2285 31717 2341 31773
rect 2369 31717 2425 31773
rect 2453 31717 2509 31773
rect 2537 31717 2593 31773
rect 1949 31636 2005 31692
rect 2033 31636 2089 31692
rect 2117 31636 2173 31692
rect 2201 31636 2257 31692
rect 2285 31636 2341 31692
rect 2369 31636 2425 31692
rect 2453 31636 2509 31692
rect 2537 31636 2593 31692
rect 1949 31555 2005 31611
rect 2033 31555 2089 31611
rect 2117 31555 2173 31611
rect 2201 31555 2257 31611
rect 2285 31555 2341 31611
rect 2369 31555 2425 31611
rect 2453 31555 2509 31611
rect 2537 31555 2593 31611
rect 1949 31474 2005 31530
rect 2033 31474 2089 31530
rect 2117 31474 2173 31530
rect 2201 31474 2257 31530
rect 2285 31474 2341 31530
rect 2369 31474 2425 31530
rect 2453 31474 2509 31530
rect 2537 31474 2593 31530
rect 1949 31393 2005 31449
rect 2033 31393 2089 31449
rect 2117 31393 2173 31449
rect 2201 31393 2257 31449
rect 2285 31393 2341 31449
rect 2369 31393 2425 31449
rect 2453 31393 2509 31449
rect 2537 31393 2593 31449
rect 1949 31312 2005 31368
rect 2033 31312 2089 31368
rect 2117 31312 2173 31368
rect 2201 31312 2257 31368
rect 2285 31312 2341 31368
rect 2369 31312 2425 31368
rect 2453 31312 2509 31368
rect 2537 31312 2593 31368
rect 1949 31231 2005 31287
rect 2033 31231 2089 31287
rect 2117 31231 2173 31287
rect 2201 31231 2257 31287
rect 2285 31231 2341 31287
rect 2369 31231 2425 31287
rect 2453 31231 2509 31287
rect 2537 31231 2593 31287
rect 1949 31150 2005 31206
rect 2033 31150 2089 31206
rect 2117 31150 2173 31206
rect 2201 31150 2257 31206
rect 2285 31150 2341 31206
rect 2369 31150 2425 31206
rect 2453 31150 2509 31206
rect 2537 31150 2593 31206
rect 1949 31069 2005 31125
rect 2033 31069 2089 31125
rect 2117 31069 2173 31125
rect 2201 31069 2257 31125
rect 2285 31069 2341 31125
rect 2369 31069 2425 31125
rect 2453 31069 2509 31125
rect 2537 31069 2593 31125
rect 1949 30988 2005 31044
rect 2033 30988 2089 31044
rect 2117 30988 2173 31044
rect 2201 30988 2257 31044
rect 2285 30988 2341 31044
rect 2369 30988 2425 31044
rect 2453 30988 2509 31044
rect 2537 30988 2593 31044
rect 1949 30907 2005 30963
rect 2033 30907 2089 30963
rect 2117 30907 2173 30963
rect 2201 30907 2257 30963
rect 2285 30907 2341 30963
rect 2369 30907 2425 30963
rect 2453 30907 2509 30963
rect 2537 30907 2593 30963
rect 1949 30826 2005 30882
rect 2033 30826 2089 30882
rect 2117 30826 2173 30882
rect 2201 30826 2257 30882
rect 2285 30826 2341 30882
rect 2369 30826 2425 30882
rect 2453 30826 2509 30882
rect 2537 30826 2593 30882
rect 1949 30745 2005 30801
rect 2033 30745 2089 30801
rect 2117 30745 2173 30801
rect 2201 30745 2257 30801
rect 2285 30745 2341 30801
rect 2369 30745 2425 30801
rect 2453 30745 2509 30801
rect 2537 30745 2593 30801
rect 1949 30664 2005 30720
rect 2033 30664 2089 30720
rect 2117 30664 2173 30720
rect 2201 30664 2257 30720
rect 2285 30664 2341 30720
rect 2369 30664 2425 30720
rect 2453 30664 2509 30720
rect 2537 30664 2593 30720
rect 1949 30583 2005 30639
rect 2033 30583 2089 30639
rect 2117 30583 2173 30639
rect 2201 30583 2257 30639
rect 2285 30583 2341 30639
rect 2369 30583 2425 30639
rect 2453 30583 2509 30639
rect 2537 30583 2593 30639
rect 1949 30502 2005 30558
rect 2033 30502 2089 30558
rect 2117 30502 2173 30558
rect 2201 30502 2257 30558
rect 2285 30502 2341 30558
rect 2369 30502 2425 30558
rect 2453 30502 2509 30558
rect 2537 30502 2593 30558
rect 1949 30421 2005 30477
rect 2033 30421 2089 30477
rect 2117 30421 2173 30477
rect 2201 30421 2257 30477
rect 2285 30421 2341 30477
rect 2369 30421 2425 30477
rect 2453 30421 2509 30477
rect 2537 30421 2593 30477
rect 1949 30340 2005 30396
rect 2033 30340 2089 30396
rect 2117 30340 2173 30396
rect 2201 30340 2257 30396
rect 2285 30340 2341 30396
rect 2369 30340 2425 30396
rect 2453 30340 2509 30396
rect 2537 30340 2593 30396
rect 1949 30259 2005 30315
rect 2033 30259 2089 30315
rect 2117 30259 2173 30315
rect 2201 30259 2257 30315
rect 2285 30259 2341 30315
rect 2369 30259 2425 30315
rect 2453 30259 2509 30315
rect 2537 30259 2593 30315
rect 1949 30178 2005 30234
rect 2033 30178 2089 30234
rect 2117 30178 2173 30234
rect 2201 30178 2257 30234
rect 2285 30178 2341 30234
rect 2369 30178 2425 30234
rect 2453 30178 2509 30234
rect 2537 30178 2593 30234
rect 2915 34739 2971 34795
rect 3001 34739 3057 34795
rect 3087 34739 3143 34795
rect 3173 34739 3229 34795
rect 3259 34739 3315 34795
rect 3345 34739 3401 34795
rect 3431 34739 3487 34795
rect 2915 34659 2971 34715
rect 3001 34659 3057 34715
rect 3087 34659 3143 34715
rect 3173 34659 3229 34715
rect 3259 34659 3315 34715
rect 3345 34659 3401 34715
rect 3431 34659 3487 34715
rect 2915 34579 2971 34635
rect 3001 34579 3057 34635
rect 3087 34579 3143 34635
rect 3173 34579 3229 34635
rect 3259 34579 3315 34635
rect 3345 34579 3401 34635
rect 3431 34579 3487 34635
rect 2915 34499 2971 34555
rect 3001 34499 3057 34555
rect 3087 34499 3143 34555
rect 3173 34499 3229 34555
rect 3259 34499 3315 34555
rect 3345 34499 3401 34555
rect 3431 34499 3487 34555
rect 2915 34419 2971 34475
rect 3001 34419 3057 34475
rect 3087 34419 3143 34475
rect 3173 34419 3229 34475
rect 3259 34419 3315 34475
rect 3345 34419 3401 34475
rect 3431 34419 3487 34475
rect 2915 34339 2971 34395
rect 3001 34339 3057 34395
rect 3087 34339 3143 34395
rect 3173 34339 3229 34395
rect 3259 34339 3315 34395
rect 3345 34339 3401 34395
rect 3431 34339 3487 34395
rect 2915 34259 2971 34315
rect 3001 34259 3057 34315
rect 3087 34259 3143 34315
rect 3173 34259 3229 34315
rect 3259 34259 3315 34315
rect 3345 34259 3401 34315
rect 3431 34259 3487 34315
rect 2915 34179 2971 34235
rect 3001 34179 3057 34235
rect 3087 34179 3143 34235
rect 3173 34179 3229 34235
rect 3259 34179 3315 34235
rect 3345 34179 3401 34235
rect 3431 34179 3487 34235
rect 2915 34099 2971 34155
rect 3001 34099 3057 34155
rect 3087 34099 3143 34155
rect 3173 34099 3229 34155
rect 3259 34099 3315 34155
rect 3345 34099 3401 34155
rect 3431 34099 3487 34155
rect 2915 34019 2971 34075
rect 3001 34019 3057 34075
rect 3087 34019 3143 34075
rect 3173 34019 3229 34075
rect 3259 34019 3315 34075
rect 3345 34019 3401 34075
rect 3431 34019 3487 34075
rect 2915 33939 2971 33995
rect 3001 33939 3057 33995
rect 3087 33939 3143 33995
rect 3173 33939 3229 33995
rect 3259 33939 3315 33995
rect 3345 33939 3401 33995
rect 3431 33939 3487 33995
rect 2915 33859 2971 33915
rect 3001 33859 3057 33915
rect 3087 33859 3143 33915
rect 3173 33859 3229 33915
rect 3259 33859 3315 33915
rect 3345 33859 3401 33915
rect 3431 33859 3487 33915
rect 2915 33779 2971 33835
rect 3001 33779 3057 33835
rect 3087 33779 3143 33835
rect 3173 33779 3229 33835
rect 3259 33779 3315 33835
rect 3345 33779 3401 33835
rect 3431 33779 3487 33835
rect 2915 33699 2971 33755
rect 3001 33699 3057 33755
rect 3087 33699 3143 33755
rect 3173 33699 3229 33755
rect 3259 33699 3315 33755
rect 3345 33699 3401 33755
rect 3431 33699 3487 33755
rect 2915 33619 2971 33675
rect 3001 33619 3057 33675
rect 3087 33619 3143 33675
rect 3173 33619 3229 33675
rect 3259 33619 3315 33675
rect 3345 33619 3401 33675
rect 3431 33619 3487 33675
rect 2915 33539 2971 33595
rect 3001 33539 3057 33595
rect 3087 33539 3143 33595
rect 3173 33539 3229 33595
rect 3259 33539 3315 33595
rect 3345 33539 3401 33595
rect 3431 33539 3487 33595
rect 2915 33459 2971 33515
rect 3001 33459 3057 33515
rect 3087 33459 3143 33515
rect 3173 33459 3229 33515
rect 3259 33459 3315 33515
rect 3345 33459 3401 33515
rect 3431 33459 3487 33515
rect 2915 33379 2971 33435
rect 3001 33379 3057 33435
rect 3087 33379 3143 33435
rect 3173 33379 3229 33435
rect 3259 33379 3315 33435
rect 3345 33379 3401 33435
rect 3431 33379 3487 33435
rect 2915 33299 2971 33355
rect 3001 33299 3057 33355
rect 3087 33299 3143 33355
rect 3173 33299 3229 33355
rect 3259 33299 3315 33355
rect 3345 33299 3401 33355
rect 3431 33299 3487 33355
rect 2915 33219 2971 33275
rect 3001 33219 3057 33275
rect 3087 33219 3143 33275
rect 3173 33219 3229 33275
rect 3259 33219 3315 33275
rect 3345 33219 3401 33275
rect 3431 33219 3487 33275
rect 2915 33139 2971 33195
rect 3001 33139 3057 33195
rect 3087 33139 3143 33195
rect 3173 33139 3229 33195
rect 3259 33139 3315 33195
rect 3345 33139 3401 33195
rect 3431 33139 3487 33195
rect 2915 33059 2971 33115
rect 3001 33059 3057 33115
rect 3087 33059 3143 33115
rect 3173 33059 3229 33115
rect 3259 33059 3315 33115
rect 3345 33059 3401 33115
rect 3431 33059 3487 33115
rect 2915 32979 2971 33035
rect 3001 32979 3057 33035
rect 3087 32979 3143 33035
rect 3173 32979 3229 33035
rect 3259 32979 3315 33035
rect 3345 32979 3401 33035
rect 3431 32979 3487 33035
rect 2915 32899 2971 32955
rect 3001 32899 3057 32955
rect 3087 32899 3143 32955
rect 3173 32899 3229 32955
rect 3259 32899 3315 32955
rect 3345 32899 3401 32955
rect 3431 32899 3487 32955
rect 2915 32819 2971 32875
rect 3001 32819 3057 32875
rect 3087 32819 3143 32875
rect 3173 32819 3229 32875
rect 3259 32819 3315 32875
rect 3345 32819 3401 32875
rect 3431 32819 3487 32875
rect 2915 32739 2971 32795
rect 3001 32739 3057 32795
rect 3087 32739 3143 32795
rect 3173 32739 3229 32795
rect 3259 32739 3315 32795
rect 3345 32739 3401 32795
rect 3431 32739 3487 32795
rect 2915 32659 2971 32715
rect 3001 32659 3057 32715
rect 3087 32659 3143 32715
rect 3173 32659 3229 32715
rect 3259 32659 3315 32715
rect 3345 32659 3401 32715
rect 3431 32659 3487 32715
rect 2915 32579 2971 32635
rect 3001 32579 3057 32635
rect 3087 32579 3143 32635
rect 3173 32579 3229 32635
rect 3259 32579 3315 32635
rect 3345 32579 3401 32635
rect 3431 32579 3487 32635
rect 2915 32499 2971 32555
rect 3001 32499 3057 32555
rect 3087 32499 3143 32555
rect 3173 32499 3229 32555
rect 3259 32499 3315 32555
rect 3345 32499 3401 32555
rect 3431 32499 3487 32555
rect 2915 32419 2971 32475
rect 3001 32419 3057 32475
rect 3087 32419 3143 32475
rect 3173 32419 3229 32475
rect 3259 32419 3315 32475
rect 3345 32419 3401 32475
rect 3431 32419 3487 32475
rect 2915 32339 2971 32395
rect 3001 32339 3057 32395
rect 3087 32339 3143 32395
rect 3173 32339 3229 32395
rect 3259 32339 3315 32395
rect 3345 32339 3401 32395
rect 3431 32339 3487 32395
rect 2915 32259 2971 32315
rect 3001 32259 3057 32315
rect 3087 32259 3143 32315
rect 3173 32259 3229 32315
rect 3259 32259 3315 32315
rect 3345 32259 3401 32315
rect 3431 32259 3487 32315
rect 2915 32179 2971 32235
rect 3001 32179 3057 32235
rect 3087 32179 3143 32235
rect 3173 32179 3229 32235
rect 3259 32179 3315 32235
rect 3345 32179 3401 32235
rect 3431 32179 3487 32235
rect 2915 32099 2971 32155
rect 3001 32099 3057 32155
rect 3087 32099 3143 32155
rect 3173 32099 3229 32155
rect 3259 32099 3315 32155
rect 3345 32099 3401 32155
rect 3431 32099 3487 32155
rect 2915 32019 2971 32075
rect 3001 32019 3057 32075
rect 3087 32019 3143 32075
rect 3173 32019 3229 32075
rect 3259 32019 3315 32075
rect 3345 32019 3401 32075
rect 3431 32019 3487 32075
rect 2915 31939 2971 31995
rect 3001 31939 3057 31995
rect 3087 31939 3143 31995
rect 3173 31939 3229 31995
rect 3259 31939 3315 31995
rect 3345 31939 3401 31995
rect 3431 31939 3487 31995
rect 2915 31859 2971 31915
rect 3001 31859 3057 31915
rect 3087 31859 3143 31915
rect 3173 31859 3229 31915
rect 3259 31859 3315 31915
rect 3345 31859 3401 31915
rect 3431 31859 3487 31915
rect 2915 31779 2971 31835
rect 3001 31779 3057 31835
rect 3087 31779 3143 31835
rect 3173 31779 3229 31835
rect 3259 31779 3315 31835
rect 3345 31779 3401 31835
rect 3431 31779 3487 31835
rect 2915 31699 2971 31755
rect 3001 31699 3057 31755
rect 3087 31699 3143 31755
rect 3173 31699 3229 31755
rect 3259 31699 3315 31755
rect 3345 31699 3401 31755
rect 3431 31699 3487 31755
rect 2915 31619 2971 31675
rect 3001 31619 3057 31675
rect 3087 31619 3143 31675
rect 3173 31619 3229 31675
rect 3259 31619 3315 31675
rect 3345 31619 3401 31675
rect 3431 31619 3487 31675
rect 2915 31539 2971 31595
rect 3001 31539 3057 31595
rect 3087 31539 3143 31595
rect 3173 31539 3229 31595
rect 3259 31539 3315 31595
rect 3345 31539 3401 31595
rect 3431 31539 3487 31595
rect 2915 31459 2971 31515
rect 3001 31459 3057 31515
rect 3087 31459 3143 31515
rect 3173 31459 3229 31515
rect 3259 31459 3315 31515
rect 3345 31459 3401 31515
rect 3431 31459 3487 31515
rect 2915 31379 2971 31435
rect 3001 31379 3057 31435
rect 3087 31379 3143 31435
rect 3173 31379 3229 31435
rect 3259 31379 3315 31435
rect 3345 31379 3401 31435
rect 3431 31379 3487 31435
rect 2915 31299 2971 31355
rect 3001 31299 3057 31355
rect 3087 31299 3143 31355
rect 3173 31299 3229 31355
rect 3259 31299 3315 31355
rect 3345 31299 3401 31355
rect 3431 31299 3487 31355
rect 2915 31219 2971 31275
rect 3001 31219 3057 31275
rect 3087 31219 3143 31275
rect 3173 31219 3229 31275
rect 3259 31219 3315 31275
rect 3345 31219 3401 31275
rect 3431 31219 3487 31275
rect 2915 31139 2971 31195
rect 3001 31139 3057 31195
rect 3087 31139 3143 31195
rect 3173 31139 3229 31195
rect 3259 31139 3315 31195
rect 3345 31139 3401 31195
rect 3431 31139 3487 31195
rect 2915 31059 2971 31115
rect 3001 31059 3057 31115
rect 3087 31059 3143 31115
rect 3173 31059 3229 31115
rect 3259 31059 3315 31115
rect 3345 31059 3401 31115
rect 3431 31059 3487 31115
rect 2915 30979 2971 31035
rect 3001 30979 3057 31035
rect 3087 30979 3143 31035
rect 3173 30979 3229 31035
rect 3259 30979 3315 31035
rect 3345 30979 3401 31035
rect 3431 30979 3487 31035
rect 2915 30899 2971 30955
rect 3001 30899 3057 30955
rect 3087 30899 3143 30955
rect 3173 30899 3229 30955
rect 3259 30899 3315 30955
rect 3345 30899 3401 30955
rect 3431 30899 3487 30955
rect 2915 30819 2971 30875
rect 3001 30819 3057 30875
rect 3087 30819 3143 30875
rect 3173 30819 3229 30875
rect 3259 30819 3315 30875
rect 3345 30819 3401 30875
rect 3431 30819 3487 30875
rect 2915 30739 2971 30795
rect 3001 30739 3057 30795
rect 3087 30739 3143 30795
rect 3173 30739 3229 30795
rect 3259 30739 3315 30795
rect 3345 30739 3401 30795
rect 3431 30739 3487 30795
rect 2915 30659 2971 30715
rect 3001 30659 3057 30715
rect 3087 30659 3143 30715
rect 3173 30659 3229 30715
rect 3259 30659 3315 30715
rect 3345 30659 3401 30715
rect 3431 30659 3487 30715
rect 2915 30579 2971 30635
rect 3001 30579 3057 30635
rect 3087 30579 3143 30635
rect 3173 30579 3229 30635
rect 3259 30579 3315 30635
rect 3345 30579 3401 30635
rect 3431 30579 3487 30635
rect 2915 30499 2971 30555
rect 3001 30499 3057 30555
rect 3087 30499 3143 30555
rect 3173 30499 3229 30555
rect 3259 30499 3315 30555
rect 3345 30499 3401 30555
rect 3431 30499 3487 30555
rect 2915 30419 2971 30475
rect 3001 30419 3057 30475
rect 3087 30419 3143 30475
rect 3173 30419 3229 30475
rect 3259 30419 3315 30475
rect 3345 30419 3401 30475
rect 3431 30419 3487 30475
rect 2915 30339 2971 30395
rect 3001 30339 3057 30395
rect 3087 30339 3143 30395
rect 3173 30339 3229 30395
rect 3259 30339 3315 30395
rect 3345 30339 3401 30395
rect 3431 30339 3487 30395
rect 2915 30259 2971 30315
rect 3001 30259 3057 30315
rect 3087 30259 3143 30315
rect 3173 30259 3229 30315
rect 3259 30259 3315 30315
rect 3345 30259 3401 30315
rect 3431 30259 3487 30315
rect 2915 30179 2971 30235
rect 3001 30179 3057 30235
rect 3087 30179 3143 30235
rect 3173 30179 3229 30235
rect 3259 30179 3315 30235
rect 3345 30179 3401 30235
rect 3431 30179 3487 30235
rect 2915 30099 2971 30155
rect 3001 30099 3057 30155
rect 3087 30099 3143 30155
rect 3173 30099 3229 30155
rect 3259 30099 3315 30155
rect 3345 30099 3401 30155
rect 3431 30099 3487 30155
rect 2915 30019 2971 30075
rect 3001 30019 3057 30075
rect 3087 30019 3143 30075
rect 3173 30019 3229 30075
rect 3259 30019 3315 30075
rect 3345 30019 3401 30075
rect 3431 30019 3487 30075
rect 6903 37094 6959 37150
rect 6993 37094 7049 37150
rect 7083 37094 7139 37150
rect 7173 37094 7229 37150
rect 7263 37094 7319 37150
rect 7353 37094 7409 37150
rect 7443 37094 7499 37150
rect 6903 37014 6959 37070
rect 6993 37014 7049 37070
rect 7083 37014 7139 37070
rect 7173 37014 7229 37070
rect 7263 37014 7319 37070
rect 7353 37014 7409 37070
rect 7443 37014 7499 37070
rect 6903 36934 6959 36990
rect 6993 36934 7049 36990
rect 7083 36934 7139 36990
rect 7173 36934 7229 36990
rect 7263 36934 7319 36990
rect 7353 36934 7409 36990
rect 7443 36934 7499 36990
rect 6903 36854 6959 36910
rect 6993 36854 7049 36910
rect 7083 36854 7139 36910
rect 7173 36854 7229 36910
rect 7263 36854 7319 36910
rect 7353 36854 7409 36910
rect 7443 36854 7499 36910
rect 6903 36774 6959 36830
rect 6993 36774 7049 36830
rect 7083 36774 7139 36830
rect 7173 36774 7229 36830
rect 7263 36774 7319 36830
rect 7353 36774 7409 36830
rect 7443 36774 7499 36830
rect 6903 36694 6959 36750
rect 6993 36694 7049 36750
rect 7083 36694 7139 36750
rect 7173 36694 7229 36750
rect 7263 36694 7319 36750
rect 7353 36694 7409 36750
rect 7443 36694 7499 36750
rect 6903 36614 6959 36670
rect 6993 36614 7049 36670
rect 7083 36614 7139 36670
rect 7173 36614 7229 36670
rect 7263 36614 7319 36670
rect 7353 36614 7409 36670
rect 7443 36614 7499 36670
rect 6903 36534 6959 36590
rect 6993 36534 7049 36590
rect 7083 36534 7139 36590
rect 7173 36534 7229 36590
rect 7263 36534 7319 36590
rect 7353 36534 7409 36590
rect 7443 36534 7499 36590
rect 6903 36454 6959 36510
rect 6993 36454 7049 36510
rect 7083 36454 7139 36510
rect 7173 36454 7229 36510
rect 7263 36454 7319 36510
rect 7353 36454 7409 36510
rect 7443 36454 7499 36510
rect 6903 36374 6959 36430
rect 6993 36374 7049 36430
rect 7083 36374 7139 36430
rect 7173 36374 7229 36430
rect 7263 36374 7319 36430
rect 7353 36374 7409 36430
rect 7443 36374 7499 36430
rect 6903 36294 6959 36350
rect 6993 36294 7049 36350
rect 7083 36294 7139 36350
rect 7173 36294 7229 36350
rect 7263 36294 7319 36350
rect 7353 36294 7409 36350
rect 7443 36294 7499 36350
rect 6903 36214 6959 36270
rect 6993 36214 7049 36270
rect 7083 36214 7139 36270
rect 7173 36214 7229 36270
rect 7263 36214 7319 36270
rect 7353 36214 7409 36270
rect 7443 36214 7499 36270
rect 6903 36134 6959 36190
rect 6993 36134 7049 36190
rect 7083 36134 7139 36190
rect 7173 36134 7229 36190
rect 7263 36134 7319 36190
rect 7353 36134 7409 36190
rect 7443 36134 7499 36190
rect 6903 36054 6959 36110
rect 6993 36054 7049 36110
rect 7083 36054 7139 36110
rect 7173 36054 7229 36110
rect 7263 36054 7319 36110
rect 7353 36054 7409 36110
rect 7443 36054 7499 36110
rect 6903 35974 6959 36030
rect 6993 35974 7049 36030
rect 7083 35974 7139 36030
rect 7173 35974 7229 36030
rect 7263 35974 7319 36030
rect 7353 35974 7409 36030
rect 7443 35974 7499 36030
rect 6903 35894 6959 35950
rect 6993 35894 7049 35950
rect 7083 35894 7139 35950
rect 7173 35894 7229 35950
rect 7263 35894 7319 35950
rect 7353 35894 7409 35950
rect 7443 35894 7499 35950
rect 6903 35814 6959 35870
rect 6993 35814 7049 35870
rect 7083 35814 7139 35870
rect 7173 35814 7229 35870
rect 7263 35814 7319 35870
rect 7353 35814 7409 35870
rect 7443 35814 7499 35870
rect 6903 35734 6959 35790
rect 6993 35734 7049 35790
rect 7083 35734 7139 35790
rect 7173 35734 7229 35790
rect 7263 35734 7319 35790
rect 7353 35734 7409 35790
rect 7443 35734 7499 35790
rect 6903 35654 6959 35710
rect 6993 35654 7049 35710
rect 7083 35654 7139 35710
rect 7173 35654 7229 35710
rect 7263 35654 7319 35710
rect 7353 35654 7409 35710
rect 7443 35654 7499 35710
rect 6903 35574 6959 35630
rect 6993 35574 7049 35630
rect 7083 35574 7139 35630
rect 7173 35574 7229 35630
rect 7263 35574 7319 35630
rect 7353 35574 7409 35630
rect 7443 35574 7499 35630
rect 6903 35494 6959 35550
rect 6993 35494 7049 35550
rect 7083 35494 7139 35550
rect 7173 35494 7229 35550
rect 7263 35494 7319 35550
rect 7353 35494 7409 35550
rect 7443 35494 7499 35550
rect 6903 35414 6959 35470
rect 6993 35414 7049 35470
rect 7083 35414 7139 35470
rect 7173 35414 7229 35470
rect 7263 35414 7319 35470
rect 7353 35414 7409 35470
rect 7443 35414 7499 35470
rect 6903 35334 6959 35390
rect 6993 35334 7049 35390
rect 7083 35334 7139 35390
rect 7173 35334 7229 35390
rect 7263 35334 7319 35390
rect 7353 35334 7409 35390
rect 7443 35334 7499 35390
rect 6903 35254 6959 35310
rect 6993 35254 7049 35310
rect 7083 35254 7139 35310
rect 7173 35254 7229 35310
rect 7263 35254 7319 35310
rect 7353 35254 7409 35310
rect 7443 35254 7499 35310
rect 6903 35174 6959 35230
rect 6993 35174 7049 35230
rect 7083 35174 7139 35230
rect 7173 35174 7229 35230
rect 7263 35174 7319 35230
rect 7353 35174 7409 35230
rect 7443 35174 7499 35230
rect 6903 35094 6959 35150
rect 6993 35094 7049 35150
rect 7083 35094 7139 35150
rect 7173 35094 7229 35150
rect 7263 35094 7319 35150
rect 7353 35094 7409 35150
rect 7443 35094 7499 35150
rect 6903 35014 6959 35070
rect 6993 35014 7049 35070
rect 7083 35014 7139 35070
rect 7173 35014 7229 35070
rect 7263 35014 7319 35070
rect 7353 35014 7409 35070
rect 7443 35014 7499 35070
rect 6903 34934 6959 34990
rect 6993 34934 7049 34990
rect 7083 34934 7139 34990
rect 7173 34934 7229 34990
rect 7263 34934 7319 34990
rect 7353 34934 7409 34990
rect 7443 34934 7499 34990
rect 6903 34854 6959 34910
rect 6993 34854 7049 34910
rect 7083 34854 7139 34910
rect 7173 34854 7229 34910
rect 7263 34854 7319 34910
rect 7353 34854 7409 34910
rect 7443 34854 7499 34910
rect 5905 34739 5961 34795
rect 5991 34739 6047 34795
rect 6077 34739 6133 34795
rect 6163 34739 6219 34795
rect 6249 34739 6305 34795
rect 6335 34739 6391 34795
rect 6421 34739 6477 34795
rect 5905 34659 5961 34715
rect 5991 34659 6047 34715
rect 6077 34659 6133 34715
rect 6163 34659 6219 34715
rect 6249 34659 6305 34715
rect 6335 34659 6391 34715
rect 6421 34659 6477 34715
rect 5905 34579 5961 34635
rect 5991 34579 6047 34635
rect 6077 34579 6133 34635
rect 6163 34579 6219 34635
rect 6249 34579 6305 34635
rect 6335 34579 6391 34635
rect 6421 34579 6477 34635
rect 5905 34499 5961 34555
rect 5991 34499 6047 34555
rect 6077 34499 6133 34555
rect 6163 34499 6219 34555
rect 6249 34499 6305 34555
rect 6335 34499 6391 34555
rect 6421 34499 6477 34555
rect 5905 34419 5961 34475
rect 5991 34419 6047 34475
rect 6077 34419 6133 34475
rect 6163 34419 6219 34475
rect 6249 34419 6305 34475
rect 6335 34419 6391 34475
rect 6421 34419 6477 34475
rect 5905 34339 5961 34395
rect 5991 34339 6047 34395
rect 6077 34339 6133 34395
rect 6163 34339 6219 34395
rect 6249 34339 6305 34395
rect 6335 34339 6391 34395
rect 6421 34339 6477 34395
rect 5905 34259 5961 34315
rect 5991 34259 6047 34315
rect 6077 34259 6133 34315
rect 6163 34259 6219 34315
rect 6249 34259 6305 34315
rect 6335 34259 6391 34315
rect 6421 34259 6477 34315
rect 5905 34179 5961 34235
rect 5991 34179 6047 34235
rect 6077 34179 6133 34235
rect 6163 34179 6219 34235
rect 6249 34179 6305 34235
rect 6335 34179 6391 34235
rect 6421 34179 6477 34235
rect 5905 34099 5961 34155
rect 5991 34099 6047 34155
rect 6077 34099 6133 34155
rect 6163 34099 6219 34155
rect 6249 34099 6305 34155
rect 6335 34099 6391 34155
rect 6421 34099 6477 34155
rect 5905 34019 5961 34075
rect 5991 34019 6047 34075
rect 6077 34019 6133 34075
rect 6163 34019 6219 34075
rect 6249 34019 6305 34075
rect 6335 34019 6391 34075
rect 6421 34019 6477 34075
rect 5905 33939 5961 33995
rect 5991 33939 6047 33995
rect 6077 33939 6133 33995
rect 6163 33939 6219 33995
rect 6249 33939 6305 33995
rect 6335 33939 6391 33995
rect 6421 33939 6477 33995
rect 5905 33859 5961 33915
rect 5991 33859 6047 33915
rect 6077 33859 6133 33915
rect 6163 33859 6219 33915
rect 6249 33859 6305 33915
rect 6335 33859 6391 33915
rect 6421 33859 6477 33915
rect 5905 33779 5961 33835
rect 5991 33779 6047 33835
rect 6077 33779 6133 33835
rect 6163 33779 6219 33835
rect 6249 33779 6305 33835
rect 6335 33779 6391 33835
rect 6421 33779 6477 33835
rect 5905 33699 5961 33755
rect 5991 33699 6047 33755
rect 6077 33699 6133 33755
rect 6163 33699 6219 33755
rect 6249 33699 6305 33755
rect 6335 33699 6391 33755
rect 6421 33699 6477 33755
rect 5905 33619 5961 33675
rect 5991 33619 6047 33675
rect 6077 33619 6133 33675
rect 6163 33619 6219 33675
rect 6249 33619 6305 33675
rect 6335 33619 6391 33675
rect 6421 33619 6477 33675
rect 5905 33539 5961 33595
rect 5991 33539 6047 33595
rect 6077 33539 6133 33595
rect 6163 33539 6219 33595
rect 6249 33539 6305 33595
rect 6335 33539 6391 33595
rect 6421 33539 6477 33595
rect 5905 33459 5961 33515
rect 5991 33459 6047 33515
rect 6077 33459 6133 33515
rect 6163 33459 6219 33515
rect 6249 33459 6305 33515
rect 6335 33459 6391 33515
rect 6421 33459 6477 33515
rect 5905 33379 5961 33435
rect 5991 33379 6047 33435
rect 6077 33379 6133 33435
rect 6163 33379 6219 33435
rect 6249 33379 6305 33435
rect 6335 33379 6391 33435
rect 6421 33379 6477 33435
rect 5905 33299 5961 33355
rect 5991 33299 6047 33355
rect 6077 33299 6133 33355
rect 6163 33299 6219 33355
rect 6249 33299 6305 33355
rect 6335 33299 6391 33355
rect 6421 33299 6477 33355
rect 5905 33219 5961 33275
rect 5991 33219 6047 33275
rect 6077 33219 6133 33275
rect 6163 33219 6219 33275
rect 6249 33219 6305 33275
rect 6335 33219 6391 33275
rect 6421 33219 6477 33275
rect 5905 33139 5961 33195
rect 5991 33139 6047 33195
rect 6077 33139 6133 33195
rect 6163 33139 6219 33195
rect 6249 33139 6305 33195
rect 6335 33139 6391 33195
rect 6421 33139 6477 33195
rect 5905 33059 5961 33115
rect 5991 33059 6047 33115
rect 6077 33059 6133 33115
rect 6163 33059 6219 33115
rect 6249 33059 6305 33115
rect 6335 33059 6391 33115
rect 6421 33059 6477 33115
rect 5905 32979 5961 33035
rect 5991 32979 6047 33035
rect 6077 32979 6133 33035
rect 6163 32979 6219 33035
rect 6249 32979 6305 33035
rect 6335 32979 6391 33035
rect 6421 32979 6477 33035
rect 5905 32899 5961 32955
rect 5991 32899 6047 32955
rect 6077 32899 6133 32955
rect 6163 32899 6219 32955
rect 6249 32899 6305 32955
rect 6335 32899 6391 32955
rect 6421 32899 6477 32955
rect 5905 32819 5961 32875
rect 5991 32819 6047 32875
rect 6077 32819 6133 32875
rect 6163 32819 6219 32875
rect 6249 32819 6305 32875
rect 6335 32819 6391 32875
rect 6421 32819 6477 32875
rect 5905 32739 5961 32795
rect 5991 32739 6047 32795
rect 6077 32739 6133 32795
rect 6163 32739 6219 32795
rect 6249 32739 6305 32795
rect 6335 32739 6391 32795
rect 6421 32739 6477 32795
rect 5905 32659 5961 32715
rect 5991 32659 6047 32715
rect 6077 32659 6133 32715
rect 6163 32659 6219 32715
rect 6249 32659 6305 32715
rect 6335 32659 6391 32715
rect 6421 32659 6477 32715
rect 5905 32579 5961 32635
rect 5991 32579 6047 32635
rect 6077 32579 6133 32635
rect 6163 32579 6219 32635
rect 6249 32579 6305 32635
rect 6335 32579 6391 32635
rect 6421 32579 6477 32635
rect 5905 32499 5961 32555
rect 5991 32499 6047 32555
rect 6077 32499 6133 32555
rect 6163 32499 6219 32555
rect 6249 32499 6305 32555
rect 6335 32499 6391 32555
rect 6421 32499 6477 32555
rect 5905 32419 5961 32475
rect 5991 32419 6047 32475
rect 6077 32419 6133 32475
rect 6163 32419 6219 32475
rect 6249 32419 6305 32475
rect 6335 32419 6391 32475
rect 6421 32419 6477 32475
rect 5905 32339 5961 32395
rect 5991 32339 6047 32395
rect 6077 32339 6133 32395
rect 6163 32339 6219 32395
rect 6249 32339 6305 32395
rect 6335 32339 6391 32395
rect 6421 32339 6477 32395
rect 5905 32259 5961 32315
rect 5991 32259 6047 32315
rect 6077 32259 6133 32315
rect 6163 32259 6219 32315
rect 6249 32259 6305 32315
rect 6335 32259 6391 32315
rect 6421 32259 6477 32315
rect 5905 32179 5961 32235
rect 5991 32179 6047 32235
rect 6077 32179 6133 32235
rect 6163 32179 6219 32235
rect 6249 32179 6305 32235
rect 6335 32179 6391 32235
rect 6421 32179 6477 32235
rect 5905 32099 5961 32155
rect 5991 32099 6047 32155
rect 6077 32099 6133 32155
rect 6163 32099 6219 32155
rect 6249 32099 6305 32155
rect 6335 32099 6391 32155
rect 6421 32099 6477 32155
rect 5905 32019 5961 32075
rect 5991 32019 6047 32075
rect 6077 32019 6133 32075
rect 6163 32019 6219 32075
rect 6249 32019 6305 32075
rect 6335 32019 6391 32075
rect 6421 32019 6477 32075
rect 5905 31939 5961 31995
rect 5991 31939 6047 31995
rect 6077 31939 6133 31995
rect 6163 31939 6219 31995
rect 6249 31939 6305 31995
rect 6335 31939 6391 31995
rect 6421 31939 6477 31995
rect 5905 31859 5961 31915
rect 5991 31859 6047 31915
rect 6077 31859 6133 31915
rect 6163 31859 6219 31915
rect 6249 31859 6305 31915
rect 6335 31859 6391 31915
rect 6421 31859 6477 31915
rect 5905 31779 5961 31835
rect 5991 31779 6047 31835
rect 6077 31779 6133 31835
rect 6163 31779 6219 31835
rect 6249 31779 6305 31835
rect 6335 31779 6391 31835
rect 6421 31779 6477 31835
rect 5905 31699 5961 31755
rect 5991 31699 6047 31755
rect 6077 31699 6133 31755
rect 6163 31699 6219 31755
rect 6249 31699 6305 31755
rect 6335 31699 6391 31755
rect 6421 31699 6477 31755
rect 5905 31619 5961 31675
rect 5991 31619 6047 31675
rect 6077 31619 6133 31675
rect 6163 31619 6219 31675
rect 6249 31619 6305 31675
rect 6335 31619 6391 31675
rect 6421 31619 6477 31675
rect 5905 31539 5961 31595
rect 5991 31539 6047 31595
rect 6077 31539 6133 31595
rect 6163 31539 6219 31595
rect 6249 31539 6305 31595
rect 6335 31539 6391 31595
rect 6421 31539 6477 31595
rect 5905 31459 5961 31515
rect 5991 31459 6047 31515
rect 6077 31459 6133 31515
rect 6163 31459 6219 31515
rect 6249 31459 6305 31515
rect 6335 31459 6391 31515
rect 6421 31459 6477 31515
rect 5905 31379 5961 31435
rect 5991 31379 6047 31435
rect 6077 31379 6133 31435
rect 6163 31379 6219 31435
rect 6249 31379 6305 31435
rect 6335 31379 6391 31435
rect 6421 31379 6477 31435
rect 5905 31299 5961 31355
rect 5991 31299 6047 31355
rect 6077 31299 6133 31355
rect 6163 31299 6219 31355
rect 6249 31299 6305 31355
rect 6335 31299 6391 31355
rect 6421 31299 6477 31355
rect 5905 31219 5961 31275
rect 5991 31219 6047 31275
rect 6077 31219 6133 31275
rect 6163 31219 6219 31275
rect 6249 31219 6305 31275
rect 6335 31219 6391 31275
rect 6421 31219 6477 31275
rect 5905 31139 5961 31195
rect 5991 31139 6047 31195
rect 6077 31139 6133 31195
rect 6163 31139 6219 31195
rect 6249 31139 6305 31195
rect 6335 31139 6391 31195
rect 6421 31139 6477 31195
rect 5905 31059 5961 31115
rect 5991 31059 6047 31115
rect 6077 31059 6133 31115
rect 6163 31059 6219 31115
rect 6249 31059 6305 31115
rect 6335 31059 6391 31115
rect 6421 31059 6477 31115
rect 5905 30979 5961 31035
rect 5991 30979 6047 31035
rect 6077 30979 6133 31035
rect 6163 30979 6219 31035
rect 6249 30979 6305 31035
rect 6335 30979 6391 31035
rect 6421 30979 6477 31035
rect 5905 30899 5961 30955
rect 5991 30899 6047 30955
rect 6077 30899 6133 30955
rect 6163 30899 6219 30955
rect 6249 30899 6305 30955
rect 6335 30899 6391 30955
rect 6421 30899 6477 30955
rect 5905 30819 5961 30875
rect 5991 30819 6047 30875
rect 6077 30819 6133 30875
rect 6163 30819 6219 30875
rect 6249 30819 6305 30875
rect 6335 30819 6391 30875
rect 6421 30819 6477 30875
rect 5905 30739 5961 30795
rect 5991 30739 6047 30795
rect 6077 30739 6133 30795
rect 6163 30739 6219 30795
rect 6249 30739 6305 30795
rect 6335 30739 6391 30795
rect 6421 30739 6477 30795
rect 5905 30659 5961 30715
rect 5991 30659 6047 30715
rect 6077 30659 6133 30715
rect 6163 30659 6219 30715
rect 6249 30659 6305 30715
rect 6335 30659 6391 30715
rect 6421 30659 6477 30715
rect 5905 30579 5961 30635
rect 5991 30579 6047 30635
rect 6077 30579 6133 30635
rect 6163 30579 6219 30635
rect 6249 30579 6305 30635
rect 6335 30579 6391 30635
rect 6421 30579 6477 30635
rect 5905 30499 5961 30555
rect 5991 30499 6047 30555
rect 6077 30499 6133 30555
rect 6163 30499 6219 30555
rect 6249 30499 6305 30555
rect 6335 30499 6391 30555
rect 6421 30499 6477 30555
rect 5905 30419 5961 30475
rect 5991 30419 6047 30475
rect 6077 30419 6133 30475
rect 6163 30419 6219 30475
rect 6249 30419 6305 30475
rect 6335 30419 6391 30475
rect 6421 30419 6477 30475
rect 5905 30339 5961 30395
rect 5991 30339 6047 30395
rect 6077 30339 6133 30395
rect 6163 30339 6219 30395
rect 6249 30339 6305 30395
rect 6335 30339 6391 30395
rect 6421 30339 6477 30395
rect 5905 30259 5961 30315
rect 5991 30259 6047 30315
rect 6077 30259 6133 30315
rect 6163 30259 6219 30315
rect 6249 30259 6305 30315
rect 6335 30259 6391 30315
rect 6421 30259 6477 30315
rect 5905 30179 5961 30235
rect 5991 30179 6047 30235
rect 6077 30179 6133 30235
rect 6163 30179 6219 30235
rect 6249 30179 6305 30235
rect 6335 30179 6391 30235
rect 6421 30179 6477 30235
rect 5905 30099 5961 30155
rect 5991 30099 6047 30155
rect 6077 30099 6133 30155
rect 6163 30099 6219 30155
rect 6249 30099 6305 30155
rect 6335 30099 6391 30155
rect 6421 30099 6477 30155
rect 5905 30019 5961 30075
rect 5991 30019 6047 30075
rect 6077 30019 6133 30075
rect 6163 30019 6219 30075
rect 6249 30019 6305 30075
rect 6335 30019 6391 30075
rect 6421 30019 6477 30075
rect 6903 34774 6959 34830
rect 6993 34774 7049 34830
rect 7083 34774 7139 34830
rect 7173 34774 7229 34830
rect 7263 34774 7319 34830
rect 7353 34774 7409 34830
rect 7443 34774 7499 34830
rect 6903 34694 6959 34750
rect 6993 34694 7049 34750
rect 7083 34694 7139 34750
rect 7173 34694 7229 34750
rect 7263 34694 7319 34750
rect 7353 34694 7409 34750
rect 7443 34694 7499 34750
rect 6903 34614 6959 34670
rect 6993 34614 7049 34670
rect 7083 34614 7139 34670
rect 7173 34614 7229 34670
rect 7263 34614 7319 34670
rect 7353 34614 7409 34670
rect 7443 34614 7499 34670
rect 6903 34534 6959 34590
rect 6993 34534 7049 34590
rect 7083 34534 7139 34590
rect 7173 34534 7229 34590
rect 7263 34534 7319 34590
rect 7353 34534 7409 34590
rect 7443 34534 7499 34590
rect 6903 34454 6959 34510
rect 6993 34454 7049 34510
rect 7083 34454 7139 34510
rect 7173 34454 7229 34510
rect 7263 34454 7319 34510
rect 7353 34454 7409 34510
rect 7443 34454 7499 34510
rect 6903 34374 6959 34430
rect 6993 34374 7049 34430
rect 7083 34374 7139 34430
rect 7173 34374 7229 34430
rect 7263 34374 7319 34430
rect 7353 34374 7409 34430
rect 7443 34374 7499 34430
rect 6903 34294 6959 34350
rect 6993 34294 7049 34350
rect 7083 34294 7139 34350
rect 7173 34294 7229 34350
rect 7263 34294 7319 34350
rect 7353 34294 7409 34350
rect 7443 34294 7499 34350
rect 6903 34214 6959 34270
rect 6993 34214 7049 34270
rect 7083 34214 7139 34270
rect 7173 34214 7229 34270
rect 7263 34214 7319 34270
rect 7353 34214 7409 34270
rect 7443 34214 7499 34270
rect 6903 34134 6959 34190
rect 6993 34134 7049 34190
rect 7083 34134 7139 34190
rect 7173 34134 7229 34190
rect 7263 34134 7319 34190
rect 7353 34134 7409 34190
rect 7443 34134 7499 34190
rect 6903 34054 6959 34110
rect 6993 34054 7049 34110
rect 7083 34054 7139 34110
rect 7173 34054 7229 34110
rect 7263 34054 7319 34110
rect 7353 34054 7409 34110
rect 7443 34054 7499 34110
rect 6903 33974 6959 34030
rect 6993 33974 7049 34030
rect 7083 33974 7139 34030
rect 7173 33974 7229 34030
rect 7263 33974 7319 34030
rect 7353 33974 7409 34030
rect 7443 33974 7499 34030
rect 6903 33894 6959 33950
rect 6993 33894 7049 33950
rect 7083 33894 7139 33950
rect 7173 33894 7229 33950
rect 7263 33894 7319 33950
rect 7353 33894 7409 33950
rect 7443 33894 7499 33950
rect 6903 33814 6959 33870
rect 6993 33814 7049 33870
rect 7083 33814 7139 33870
rect 7173 33814 7229 33870
rect 7263 33814 7319 33870
rect 7353 33814 7409 33870
rect 7443 33814 7499 33870
rect 6903 33734 6959 33790
rect 6993 33734 7049 33790
rect 7083 33734 7139 33790
rect 7173 33734 7229 33790
rect 7263 33734 7319 33790
rect 7353 33734 7409 33790
rect 7443 33734 7499 33790
rect 6903 33654 6959 33710
rect 6993 33654 7049 33710
rect 7083 33654 7139 33710
rect 7173 33654 7229 33710
rect 7263 33654 7319 33710
rect 7353 33654 7409 33710
rect 7443 33654 7499 33710
rect 6903 33574 6959 33630
rect 6993 33574 7049 33630
rect 7083 33574 7139 33630
rect 7173 33574 7229 33630
rect 7263 33574 7319 33630
rect 7353 33574 7409 33630
rect 7443 33574 7499 33630
rect 6903 33494 6959 33550
rect 6993 33494 7049 33550
rect 7083 33494 7139 33550
rect 7173 33494 7229 33550
rect 7263 33494 7319 33550
rect 7353 33494 7409 33550
rect 7443 33494 7499 33550
rect 6903 33414 6959 33470
rect 6993 33414 7049 33470
rect 7083 33414 7139 33470
rect 7173 33414 7229 33470
rect 7263 33414 7319 33470
rect 7353 33414 7409 33470
rect 7443 33414 7499 33470
rect 6903 33334 6959 33390
rect 6993 33334 7049 33390
rect 7083 33334 7139 33390
rect 7173 33334 7229 33390
rect 7263 33334 7319 33390
rect 7353 33334 7409 33390
rect 7443 33334 7499 33390
rect 6903 33254 6959 33310
rect 6993 33254 7049 33310
rect 7083 33254 7139 33310
rect 7173 33254 7229 33310
rect 7263 33254 7319 33310
rect 7353 33254 7409 33310
rect 7443 33254 7499 33310
rect 6903 33174 6959 33230
rect 6993 33174 7049 33230
rect 7083 33174 7139 33230
rect 7173 33174 7229 33230
rect 7263 33174 7319 33230
rect 7353 33174 7409 33230
rect 7443 33174 7499 33230
rect 6903 33094 6959 33150
rect 6993 33094 7049 33150
rect 7083 33094 7139 33150
rect 7173 33094 7229 33150
rect 7263 33094 7319 33150
rect 7353 33094 7409 33150
rect 7443 33094 7499 33150
rect 6903 33014 6959 33070
rect 6993 33014 7049 33070
rect 7083 33014 7139 33070
rect 7173 33014 7229 33070
rect 7263 33014 7319 33070
rect 7353 33014 7409 33070
rect 7443 33014 7499 33070
rect 6903 32934 6959 32990
rect 6993 32934 7049 32990
rect 7083 32934 7139 32990
rect 7173 32934 7229 32990
rect 7263 32934 7319 32990
rect 7353 32934 7409 32990
rect 7443 32934 7499 32990
rect 6903 32854 6959 32910
rect 6993 32854 7049 32910
rect 7083 32854 7139 32910
rect 7173 32854 7229 32910
rect 7263 32854 7319 32910
rect 7353 32854 7409 32910
rect 7443 32854 7499 32910
rect 6903 32774 6959 32830
rect 6993 32774 7049 32830
rect 7083 32774 7139 32830
rect 7173 32774 7229 32830
rect 7263 32774 7319 32830
rect 7353 32774 7409 32830
rect 7443 32774 7499 32830
rect 6903 32694 6959 32750
rect 6993 32694 7049 32750
rect 7083 32694 7139 32750
rect 7173 32694 7229 32750
rect 7263 32694 7319 32750
rect 7353 32694 7409 32750
rect 7443 32694 7499 32750
rect 6903 32614 6959 32670
rect 6993 32614 7049 32670
rect 7083 32614 7139 32670
rect 7173 32614 7229 32670
rect 7263 32614 7319 32670
rect 7353 32614 7409 32670
rect 7443 32614 7499 32670
rect 6903 32534 6959 32590
rect 6993 32534 7049 32590
rect 7083 32534 7139 32590
rect 7173 32534 7229 32590
rect 7263 32534 7319 32590
rect 7353 32534 7409 32590
rect 7443 32534 7499 32590
rect 6903 32454 6959 32510
rect 6993 32454 7049 32510
rect 7083 32454 7139 32510
rect 7173 32454 7229 32510
rect 7263 32454 7319 32510
rect 7353 32454 7409 32510
rect 7443 32454 7499 32510
rect 6903 32374 6959 32430
rect 6993 32374 7049 32430
rect 7083 32374 7139 32430
rect 7173 32374 7229 32430
rect 7263 32374 7319 32430
rect 7353 32374 7409 32430
rect 7443 32374 7499 32430
rect 6903 32294 6959 32350
rect 6993 32294 7049 32350
rect 7083 32294 7139 32350
rect 7173 32294 7229 32350
rect 7263 32294 7319 32350
rect 7353 32294 7409 32350
rect 7443 32294 7499 32350
rect 6903 32214 6959 32270
rect 6993 32214 7049 32270
rect 7083 32214 7139 32270
rect 7173 32214 7229 32270
rect 7263 32214 7319 32270
rect 7353 32214 7409 32270
rect 7443 32214 7499 32270
rect 6903 32134 6959 32190
rect 6993 32134 7049 32190
rect 7083 32134 7139 32190
rect 7173 32134 7229 32190
rect 7263 32134 7319 32190
rect 7353 32134 7409 32190
rect 7443 32134 7499 32190
rect 6903 32054 6959 32110
rect 6993 32054 7049 32110
rect 7083 32054 7139 32110
rect 7173 32054 7229 32110
rect 7263 32054 7319 32110
rect 7353 32054 7409 32110
rect 7443 32054 7499 32110
rect 6903 31974 6959 32030
rect 6993 31974 7049 32030
rect 7083 31974 7139 32030
rect 7173 31974 7229 32030
rect 7263 31974 7319 32030
rect 7353 31974 7409 32030
rect 7443 31974 7499 32030
rect 6903 31894 6959 31950
rect 6993 31894 7049 31950
rect 7083 31894 7139 31950
rect 7173 31894 7229 31950
rect 7263 31894 7319 31950
rect 7353 31894 7409 31950
rect 7443 31894 7499 31950
rect 6903 31814 6959 31870
rect 6993 31814 7049 31870
rect 7083 31814 7139 31870
rect 7173 31814 7229 31870
rect 7263 31814 7319 31870
rect 7353 31814 7409 31870
rect 7443 31814 7499 31870
rect 6903 31734 6959 31790
rect 6993 31734 7049 31790
rect 7083 31734 7139 31790
rect 7173 31734 7229 31790
rect 7263 31734 7319 31790
rect 7353 31734 7409 31790
rect 7443 31734 7499 31790
rect 6903 31654 6959 31710
rect 6993 31654 7049 31710
rect 7083 31654 7139 31710
rect 7173 31654 7229 31710
rect 7263 31654 7319 31710
rect 7353 31654 7409 31710
rect 7443 31654 7499 31710
rect 6903 31574 6959 31630
rect 6993 31574 7049 31630
rect 7083 31574 7139 31630
rect 7173 31574 7229 31630
rect 7263 31574 7319 31630
rect 7353 31574 7409 31630
rect 7443 31574 7499 31630
rect 6903 31494 6959 31550
rect 6993 31494 7049 31550
rect 7083 31494 7139 31550
rect 7173 31494 7229 31550
rect 7263 31494 7319 31550
rect 7353 31494 7409 31550
rect 7443 31494 7499 31550
rect 6903 31414 6959 31470
rect 6993 31414 7049 31470
rect 7083 31414 7139 31470
rect 7173 31414 7229 31470
rect 7263 31414 7319 31470
rect 7353 31414 7409 31470
rect 7443 31414 7499 31470
rect 6903 31334 6959 31390
rect 6993 31334 7049 31390
rect 7083 31334 7139 31390
rect 7173 31334 7229 31390
rect 7263 31334 7319 31390
rect 7353 31334 7409 31390
rect 7443 31334 7499 31390
rect 6903 31254 6959 31310
rect 6993 31254 7049 31310
rect 7083 31254 7139 31310
rect 7173 31254 7229 31310
rect 7263 31254 7319 31310
rect 7353 31254 7409 31310
rect 7443 31254 7499 31310
rect 6903 31174 6959 31230
rect 6993 31174 7049 31230
rect 7083 31174 7139 31230
rect 7173 31174 7229 31230
rect 7263 31174 7319 31230
rect 7353 31174 7409 31230
rect 7443 31174 7499 31230
rect 6903 31094 6959 31150
rect 6993 31094 7049 31150
rect 7083 31094 7139 31150
rect 7173 31094 7229 31150
rect 7263 31094 7319 31150
rect 7353 31094 7409 31150
rect 7443 31094 7499 31150
rect 6903 31014 6959 31070
rect 6993 31014 7049 31070
rect 7083 31014 7139 31070
rect 7173 31014 7229 31070
rect 7263 31014 7319 31070
rect 7353 31014 7409 31070
rect 7443 31014 7499 31070
rect 6903 30934 6959 30990
rect 6993 30934 7049 30990
rect 7083 30934 7139 30990
rect 7173 30934 7229 30990
rect 7263 30934 7319 30990
rect 7353 30934 7409 30990
rect 7443 30934 7499 30990
rect 6903 30854 6959 30910
rect 6993 30854 7049 30910
rect 7083 30854 7139 30910
rect 7173 30854 7229 30910
rect 7263 30854 7319 30910
rect 7353 30854 7409 30910
rect 7443 30854 7499 30910
rect 6903 30774 6959 30830
rect 6993 30774 7049 30830
rect 7083 30774 7139 30830
rect 7173 30774 7229 30830
rect 7263 30774 7319 30830
rect 7353 30774 7409 30830
rect 7443 30774 7499 30830
rect 6903 30694 6959 30750
rect 6993 30694 7049 30750
rect 7083 30694 7139 30750
rect 7173 30694 7229 30750
rect 7263 30694 7319 30750
rect 7353 30694 7409 30750
rect 7443 30694 7499 30750
rect 6903 30614 6959 30670
rect 6993 30614 7049 30670
rect 7083 30614 7139 30670
rect 7173 30614 7229 30670
rect 7263 30614 7319 30670
rect 7353 30614 7409 30670
rect 7443 30614 7499 30670
rect 6903 30534 6959 30590
rect 6993 30534 7049 30590
rect 7083 30534 7139 30590
rect 7173 30534 7229 30590
rect 7263 30534 7319 30590
rect 7353 30534 7409 30590
rect 7443 30534 7499 30590
rect 6903 30454 6959 30510
rect 6993 30454 7049 30510
rect 7083 30454 7139 30510
rect 7173 30454 7229 30510
rect 7263 30454 7319 30510
rect 7353 30454 7409 30510
rect 7443 30454 7499 30510
rect 6903 30374 6959 30430
rect 6993 30374 7049 30430
rect 7083 30374 7139 30430
rect 7173 30374 7229 30430
rect 7263 30374 7319 30430
rect 7353 30374 7409 30430
rect 7443 30374 7499 30430
rect 6903 30294 6959 30350
rect 6993 30294 7049 30350
rect 7083 30294 7139 30350
rect 7173 30294 7229 30350
rect 7263 30294 7319 30350
rect 7353 30294 7409 30350
rect 7443 30294 7499 30350
rect 6903 30214 6959 30270
rect 6993 30214 7049 30270
rect 7083 30214 7139 30270
rect 7173 30214 7229 30270
rect 7263 30214 7319 30270
rect 7353 30214 7409 30270
rect 7443 30214 7499 30270
rect 6903 30133 6959 30189
rect 6993 30133 7049 30189
rect 7083 30133 7139 30189
rect 7173 30133 7229 30189
rect 7263 30133 7319 30189
rect 7353 30133 7409 30189
rect 7443 30133 7499 30189
rect 6903 30052 6959 30108
rect 6993 30052 7049 30108
rect 7083 30052 7139 30108
rect 7173 30052 7229 30108
rect 7263 30052 7319 30108
rect 7353 30052 7409 30108
rect 7443 30052 7499 30108
rect 2915 23981 2971 24037
rect 3001 23981 3057 24037
rect 3087 23981 3143 24037
rect 3173 23981 3229 24037
rect 3259 23981 3315 24037
rect 3345 23981 3401 24037
rect 3431 23981 3487 24037
rect 2915 23901 2971 23957
rect 3001 23901 3057 23957
rect 3087 23901 3143 23957
rect 3173 23901 3229 23957
rect 3259 23901 3315 23957
rect 3345 23901 3401 23957
rect 3431 23901 3487 23957
rect 2915 23821 2971 23877
rect 3001 23821 3057 23877
rect 3087 23821 3143 23877
rect 3173 23821 3229 23877
rect 3259 23821 3315 23877
rect 3345 23821 3401 23877
rect 3431 23821 3487 23877
rect 2915 23741 2971 23797
rect 3001 23741 3057 23797
rect 3087 23741 3143 23797
rect 3173 23741 3229 23797
rect 3259 23741 3315 23797
rect 3345 23741 3401 23797
rect 3431 23741 3487 23797
rect 2915 23661 2971 23717
rect 3001 23661 3057 23717
rect 3087 23661 3143 23717
rect 3173 23661 3229 23717
rect 3259 23661 3315 23717
rect 3345 23661 3401 23717
rect 3431 23661 3487 23717
rect 2915 23581 2971 23637
rect 3001 23581 3057 23637
rect 3087 23581 3143 23637
rect 3173 23581 3229 23637
rect 3259 23581 3315 23637
rect 3345 23581 3401 23637
rect 3431 23581 3487 23637
rect 2915 23501 2971 23557
rect 3001 23501 3057 23557
rect 3087 23501 3143 23557
rect 3173 23501 3229 23557
rect 3259 23501 3315 23557
rect 3345 23501 3401 23557
rect 3431 23501 3487 23557
rect 2915 23421 2971 23477
rect 3001 23421 3057 23477
rect 3087 23421 3143 23477
rect 3173 23421 3229 23477
rect 3259 23421 3315 23477
rect 3345 23421 3401 23477
rect 3431 23421 3487 23477
rect 2915 23341 2971 23397
rect 3001 23341 3057 23397
rect 3087 23341 3143 23397
rect 3173 23341 3229 23397
rect 3259 23341 3315 23397
rect 3345 23341 3401 23397
rect 3431 23341 3487 23397
rect 2915 23261 2971 23317
rect 3001 23261 3057 23317
rect 3087 23261 3143 23317
rect 3173 23261 3229 23317
rect 3259 23261 3315 23317
rect 3345 23261 3401 23317
rect 3431 23261 3487 23317
rect 2915 23181 2971 23237
rect 3001 23181 3057 23237
rect 3087 23181 3143 23237
rect 3173 23181 3229 23237
rect 3259 23181 3315 23237
rect 3345 23181 3401 23237
rect 3431 23181 3487 23237
rect 2915 23101 2971 23157
rect 3001 23101 3057 23157
rect 3087 23101 3143 23157
rect 3173 23101 3229 23157
rect 3259 23101 3315 23157
rect 3345 23101 3401 23157
rect 3431 23101 3487 23157
rect 2915 23021 2971 23077
rect 3001 23021 3057 23077
rect 3087 23021 3143 23077
rect 3173 23021 3229 23077
rect 3259 23021 3315 23077
rect 3345 23021 3401 23077
rect 3431 23021 3487 23077
rect 2915 22941 2971 22997
rect 3001 22941 3057 22997
rect 3087 22941 3143 22997
rect 3173 22941 3229 22997
rect 3259 22941 3315 22997
rect 3345 22941 3401 22997
rect 3431 22941 3487 22997
rect 2915 22861 2971 22917
rect 3001 22861 3057 22917
rect 3087 22861 3143 22917
rect 3173 22861 3229 22917
rect 3259 22861 3315 22917
rect 3345 22861 3401 22917
rect 3431 22861 3487 22917
rect 2915 22781 2971 22837
rect 3001 22781 3057 22837
rect 3087 22781 3143 22837
rect 3173 22781 3229 22837
rect 3259 22781 3315 22837
rect 3345 22781 3401 22837
rect 3431 22781 3487 22837
rect 2915 22701 2971 22757
rect 3001 22701 3057 22757
rect 3087 22701 3143 22757
rect 3173 22701 3229 22757
rect 3259 22701 3315 22757
rect 3345 22701 3401 22757
rect 3431 22701 3487 22757
rect 2915 22621 2971 22677
rect 3001 22621 3057 22677
rect 3087 22621 3143 22677
rect 3173 22621 3229 22677
rect 3259 22621 3315 22677
rect 3345 22621 3401 22677
rect 3431 22621 3487 22677
rect 2915 22541 2971 22597
rect 3001 22541 3057 22597
rect 3087 22541 3143 22597
rect 3173 22541 3229 22597
rect 3259 22541 3315 22597
rect 3345 22541 3401 22597
rect 3431 22541 3487 22597
rect 2915 22461 2971 22517
rect 3001 22461 3057 22517
rect 3087 22461 3143 22517
rect 3173 22461 3229 22517
rect 3259 22461 3315 22517
rect 3345 22461 3401 22517
rect 3431 22461 3487 22517
rect 2915 22381 2971 22437
rect 3001 22381 3057 22437
rect 3087 22381 3143 22437
rect 3173 22381 3229 22437
rect 3259 22381 3315 22437
rect 3345 22381 3401 22437
rect 3431 22381 3487 22437
rect 2915 22301 2971 22357
rect 3001 22301 3057 22357
rect 3087 22301 3143 22357
rect 3173 22301 3229 22357
rect 3259 22301 3315 22357
rect 3345 22301 3401 22357
rect 3431 22301 3487 22357
rect 2915 22221 2971 22277
rect 3001 22221 3057 22277
rect 3087 22221 3143 22277
rect 3173 22221 3229 22277
rect 3259 22221 3315 22277
rect 3345 22221 3401 22277
rect 3431 22221 3487 22277
rect 2915 22141 2971 22197
rect 3001 22141 3057 22197
rect 3087 22141 3143 22197
rect 3173 22141 3229 22197
rect 3259 22141 3315 22197
rect 3345 22141 3401 22197
rect 3431 22141 3487 22197
rect 2915 22061 2971 22117
rect 3001 22061 3057 22117
rect 3087 22061 3143 22117
rect 3173 22061 3229 22117
rect 3259 22061 3315 22117
rect 3345 22061 3401 22117
rect 3431 22061 3487 22117
rect 2915 21981 2971 22037
rect 3001 21981 3057 22037
rect 3087 21981 3143 22037
rect 3173 21981 3229 22037
rect 3259 21981 3315 22037
rect 3345 21981 3401 22037
rect 3431 21981 3487 22037
rect 2915 21901 2971 21957
rect 3001 21901 3057 21957
rect 3087 21901 3143 21957
rect 3173 21901 3229 21957
rect 3259 21901 3315 21957
rect 3345 21901 3401 21957
rect 3431 21901 3487 21957
rect 2915 21821 2971 21877
rect 3001 21821 3057 21877
rect 3087 21821 3143 21877
rect 3173 21821 3229 21877
rect 3259 21821 3315 21877
rect 3345 21821 3401 21877
rect 3431 21821 3487 21877
rect 2915 21741 2971 21797
rect 3001 21741 3057 21797
rect 3087 21741 3143 21797
rect 3173 21741 3229 21797
rect 3259 21741 3315 21797
rect 3345 21741 3401 21797
rect 3431 21741 3487 21797
rect 2915 21661 2971 21717
rect 3001 21661 3057 21717
rect 3087 21661 3143 21717
rect 3173 21661 3229 21717
rect 3259 21661 3315 21717
rect 3345 21661 3401 21717
rect 3431 21661 3487 21717
rect 2915 21581 2971 21637
rect 3001 21581 3057 21637
rect 3087 21581 3143 21637
rect 3173 21581 3229 21637
rect 3259 21581 3315 21637
rect 3345 21581 3401 21637
rect 3431 21581 3487 21637
rect 2915 21501 2971 21557
rect 3001 21501 3057 21557
rect 3087 21501 3143 21557
rect 3173 21501 3229 21557
rect 3259 21501 3315 21557
rect 3345 21501 3401 21557
rect 3431 21501 3487 21557
rect 2915 21421 2971 21477
rect 3001 21421 3057 21477
rect 3087 21421 3143 21477
rect 3173 21421 3229 21477
rect 3259 21421 3315 21477
rect 3345 21421 3401 21477
rect 3431 21421 3487 21477
rect 2915 21341 2971 21397
rect 3001 21341 3057 21397
rect 3087 21341 3143 21397
rect 3173 21341 3229 21397
rect 3259 21341 3315 21397
rect 3345 21341 3401 21397
rect 3431 21341 3487 21397
rect 2915 21261 2971 21317
rect 3001 21261 3057 21317
rect 3087 21261 3143 21317
rect 3173 21261 3229 21317
rect 3259 21261 3315 21317
rect 3345 21261 3401 21317
rect 3431 21261 3487 21317
rect 5903 23981 5959 24037
rect 5989 23981 6045 24037
rect 6075 23981 6131 24037
rect 6161 23981 6217 24037
rect 6247 23981 6303 24037
rect 6333 23981 6389 24037
rect 6419 23981 6475 24037
rect 5903 23901 5959 23957
rect 5989 23901 6045 23957
rect 6075 23901 6131 23957
rect 6161 23901 6217 23957
rect 6247 23901 6303 23957
rect 6333 23901 6389 23957
rect 6419 23901 6475 23957
rect 5903 23821 5959 23877
rect 5989 23821 6045 23877
rect 6075 23821 6131 23877
rect 6161 23821 6217 23877
rect 6247 23821 6303 23877
rect 6333 23821 6389 23877
rect 6419 23821 6475 23877
rect 5903 23741 5959 23797
rect 5989 23741 6045 23797
rect 6075 23741 6131 23797
rect 6161 23741 6217 23797
rect 6247 23741 6303 23797
rect 6333 23741 6389 23797
rect 6419 23741 6475 23797
rect 5903 23661 5959 23717
rect 5989 23661 6045 23717
rect 6075 23661 6131 23717
rect 6161 23661 6217 23717
rect 6247 23661 6303 23717
rect 6333 23661 6389 23717
rect 6419 23661 6475 23717
rect 5903 23581 5959 23637
rect 5989 23581 6045 23637
rect 6075 23581 6131 23637
rect 6161 23581 6217 23637
rect 6247 23581 6303 23637
rect 6333 23581 6389 23637
rect 6419 23581 6475 23637
rect 5903 23501 5959 23557
rect 5989 23501 6045 23557
rect 6075 23501 6131 23557
rect 6161 23501 6217 23557
rect 6247 23501 6303 23557
rect 6333 23501 6389 23557
rect 6419 23501 6475 23557
rect 5903 23421 5959 23477
rect 5989 23421 6045 23477
rect 6075 23421 6131 23477
rect 6161 23421 6217 23477
rect 6247 23421 6303 23477
rect 6333 23421 6389 23477
rect 6419 23421 6475 23477
rect 5903 23341 5959 23397
rect 5989 23341 6045 23397
rect 6075 23341 6131 23397
rect 6161 23341 6217 23397
rect 6247 23341 6303 23397
rect 6333 23341 6389 23397
rect 6419 23341 6475 23397
rect 5903 23261 5959 23317
rect 5989 23261 6045 23317
rect 6075 23261 6131 23317
rect 6161 23261 6217 23317
rect 6247 23261 6303 23317
rect 6333 23261 6389 23317
rect 6419 23261 6475 23317
rect 5903 23181 5959 23237
rect 5989 23181 6045 23237
rect 6075 23181 6131 23237
rect 6161 23181 6217 23237
rect 6247 23181 6303 23237
rect 6333 23181 6389 23237
rect 6419 23181 6475 23237
rect 5903 23101 5959 23157
rect 5989 23101 6045 23157
rect 6075 23101 6131 23157
rect 6161 23101 6217 23157
rect 6247 23101 6303 23157
rect 6333 23101 6389 23157
rect 6419 23101 6475 23157
rect 5903 23021 5959 23077
rect 5989 23021 6045 23077
rect 6075 23021 6131 23077
rect 6161 23021 6217 23077
rect 6247 23021 6303 23077
rect 6333 23021 6389 23077
rect 6419 23021 6475 23077
rect 5903 22941 5959 22997
rect 5989 22941 6045 22997
rect 6075 22941 6131 22997
rect 6161 22941 6217 22997
rect 6247 22941 6303 22997
rect 6333 22941 6389 22997
rect 6419 22941 6475 22997
rect 5903 22861 5959 22917
rect 5989 22861 6045 22917
rect 6075 22861 6131 22917
rect 6161 22861 6217 22917
rect 6247 22861 6303 22917
rect 6333 22861 6389 22917
rect 6419 22861 6475 22917
rect 5903 22781 5959 22837
rect 5989 22781 6045 22837
rect 6075 22781 6131 22837
rect 6161 22781 6217 22837
rect 6247 22781 6303 22837
rect 6333 22781 6389 22837
rect 6419 22781 6475 22837
rect 5903 22701 5959 22757
rect 5989 22701 6045 22757
rect 6075 22701 6131 22757
rect 6161 22701 6217 22757
rect 6247 22701 6303 22757
rect 6333 22701 6389 22757
rect 6419 22701 6475 22757
rect 5903 22621 5959 22677
rect 5989 22621 6045 22677
rect 6075 22621 6131 22677
rect 6161 22621 6217 22677
rect 6247 22621 6303 22677
rect 6333 22621 6389 22677
rect 6419 22621 6475 22677
rect 5903 22541 5959 22597
rect 5989 22541 6045 22597
rect 6075 22541 6131 22597
rect 6161 22541 6217 22597
rect 6247 22541 6303 22597
rect 6333 22541 6389 22597
rect 6419 22541 6475 22597
rect 5903 22461 5959 22517
rect 5989 22461 6045 22517
rect 6075 22461 6131 22517
rect 6161 22461 6217 22517
rect 6247 22461 6303 22517
rect 6333 22461 6389 22517
rect 6419 22461 6475 22517
rect 5903 22381 5959 22437
rect 5989 22381 6045 22437
rect 6075 22381 6131 22437
rect 6161 22381 6217 22437
rect 6247 22381 6303 22437
rect 6333 22381 6389 22437
rect 6419 22381 6475 22437
rect 5903 22301 5959 22357
rect 5989 22301 6045 22357
rect 6075 22301 6131 22357
rect 6161 22301 6217 22357
rect 6247 22301 6303 22357
rect 6333 22301 6389 22357
rect 6419 22301 6475 22357
rect 5903 22221 5959 22277
rect 5989 22221 6045 22277
rect 6075 22221 6131 22277
rect 6161 22221 6217 22277
rect 6247 22221 6303 22277
rect 6333 22221 6389 22277
rect 6419 22221 6475 22277
rect 5903 22141 5959 22197
rect 5989 22141 6045 22197
rect 6075 22141 6131 22197
rect 6161 22141 6217 22197
rect 6247 22141 6303 22197
rect 6333 22141 6389 22197
rect 6419 22141 6475 22197
rect 5903 22061 5959 22117
rect 5989 22061 6045 22117
rect 6075 22061 6131 22117
rect 6161 22061 6217 22117
rect 6247 22061 6303 22117
rect 6333 22061 6389 22117
rect 6419 22061 6475 22117
rect 5903 21981 5959 22037
rect 5989 21981 6045 22037
rect 6075 21981 6131 22037
rect 6161 21981 6217 22037
rect 6247 21981 6303 22037
rect 6333 21981 6389 22037
rect 6419 21981 6475 22037
rect 5903 21901 5959 21957
rect 5989 21901 6045 21957
rect 6075 21901 6131 21957
rect 6161 21901 6217 21957
rect 6247 21901 6303 21957
rect 6333 21901 6389 21957
rect 6419 21901 6475 21957
rect 5903 21821 5959 21877
rect 5989 21821 6045 21877
rect 6075 21821 6131 21877
rect 6161 21821 6217 21877
rect 6247 21821 6303 21877
rect 6333 21821 6389 21877
rect 6419 21821 6475 21877
rect 5903 21741 5959 21797
rect 5989 21741 6045 21797
rect 6075 21741 6131 21797
rect 6161 21741 6217 21797
rect 6247 21741 6303 21797
rect 6333 21741 6389 21797
rect 6419 21741 6475 21797
rect 5903 21661 5959 21717
rect 5989 21661 6045 21717
rect 6075 21661 6131 21717
rect 6161 21661 6217 21717
rect 6247 21661 6303 21717
rect 6333 21661 6389 21717
rect 6419 21661 6475 21717
rect 5903 21581 5959 21637
rect 5989 21581 6045 21637
rect 6075 21581 6131 21637
rect 6161 21581 6217 21637
rect 6247 21581 6303 21637
rect 6333 21581 6389 21637
rect 6419 21581 6475 21637
rect 5903 21501 5959 21557
rect 5989 21501 6045 21557
rect 6075 21501 6131 21557
rect 6161 21501 6217 21557
rect 6247 21501 6303 21557
rect 6333 21501 6389 21557
rect 6419 21501 6475 21557
rect 5903 21421 5959 21477
rect 5989 21421 6045 21477
rect 6075 21421 6131 21477
rect 6161 21421 6217 21477
rect 6247 21421 6303 21477
rect 6333 21421 6389 21477
rect 6419 21421 6475 21477
rect 5903 21341 5959 21397
rect 5989 21341 6045 21397
rect 6075 21341 6131 21397
rect 6161 21341 6217 21397
rect 6247 21341 6303 21397
rect 6333 21341 6389 21397
rect 6419 21341 6475 21397
rect 2915 21181 2971 21237
rect 3001 21181 3057 21237
rect 3087 21181 3143 21237
rect 3173 21181 3229 21237
rect 3259 21181 3315 21237
rect 3345 21181 3401 21237
rect 3431 21181 3487 21237
rect 2915 21101 2971 21157
rect 3001 21101 3057 21157
rect 3087 21101 3143 21157
rect 3173 21101 3229 21157
rect 3259 21101 3315 21157
rect 3345 21101 3401 21157
rect 3431 21101 3487 21157
rect 2915 21021 2971 21077
rect 3001 21021 3057 21077
rect 3087 21021 3143 21077
rect 3173 21021 3229 21077
rect 3259 21021 3315 21077
rect 3345 21021 3401 21077
rect 3431 21021 3487 21077
rect 2915 20941 2971 20997
rect 3001 20941 3057 20997
rect 3087 20941 3143 20997
rect 3173 20941 3229 20997
rect 3259 20941 3315 20997
rect 3345 20941 3401 20997
rect 3431 20941 3487 20997
rect 2915 20861 2971 20917
rect 3001 20861 3057 20917
rect 3087 20861 3143 20917
rect 3173 20861 3229 20917
rect 3259 20861 3315 20917
rect 3345 20861 3401 20917
rect 3431 20861 3487 20917
rect 2915 20781 2971 20837
rect 3001 20781 3057 20837
rect 3087 20781 3143 20837
rect 3173 20781 3229 20837
rect 3259 20781 3315 20837
rect 3345 20781 3401 20837
rect 3431 20781 3487 20837
rect 2915 20701 2971 20757
rect 3001 20701 3057 20757
rect 3087 20701 3143 20757
rect 3173 20701 3229 20757
rect 3259 20701 3315 20757
rect 3345 20701 3401 20757
rect 3431 20701 3487 20757
rect 2915 20621 2971 20677
rect 3001 20621 3057 20677
rect 3087 20621 3143 20677
rect 3173 20621 3229 20677
rect 3259 20621 3315 20677
rect 3345 20621 3401 20677
rect 3431 20621 3487 20677
rect 2915 20541 2971 20597
rect 3001 20541 3057 20597
rect 3087 20541 3143 20597
rect 3173 20541 3229 20597
rect 3259 20541 3315 20597
rect 3345 20541 3401 20597
rect 3431 20541 3487 20597
rect 2915 20461 2971 20517
rect 3001 20461 3057 20517
rect 3087 20461 3143 20517
rect 3173 20461 3229 20517
rect 3259 20461 3315 20517
rect 3345 20461 3401 20517
rect 3431 20461 3487 20517
rect 2915 20381 2971 20437
rect 3001 20381 3057 20437
rect 3087 20381 3143 20437
rect 3173 20381 3229 20437
rect 3259 20381 3315 20437
rect 3345 20381 3401 20437
rect 3431 20381 3487 20437
rect 2915 20301 2971 20357
rect 3001 20301 3057 20357
rect 3087 20301 3143 20357
rect 3173 20301 3229 20357
rect 3259 20301 3315 20357
rect 3345 20301 3401 20357
rect 3431 20301 3487 20357
rect 2915 20221 2971 20277
rect 3001 20221 3057 20277
rect 3087 20221 3143 20277
rect 3173 20221 3229 20277
rect 3259 20221 3315 20277
rect 3345 20221 3401 20277
rect 3431 20221 3487 20277
rect 2915 20141 2971 20197
rect 3001 20141 3057 20197
rect 3087 20141 3143 20197
rect 3173 20141 3229 20197
rect 3259 20141 3315 20197
rect 3345 20141 3401 20197
rect 3431 20141 3487 20197
rect 2915 20061 2971 20117
rect 3001 20061 3057 20117
rect 3087 20061 3143 20117
rect 3173 20061 3229 20117
rect 3259 20061 3315 20117
rect 3345 20061 3401 20117
rect 3431 20061 3487 20117
rect 2915 19981 2971 20037
rect 3001 19981 3057 20037
rect 3087 19981 3143 20037
rect 3173 19981 3229 20037
rect 3259 19981 3315 20037
rect 3345 19981 3401 20037
rect 3431 19981 3487 20037
rect 2915 19901 2971 19957
rect 3001 19901 3057 19957
rect 3087 19901 3143 19957
rect 3173 19901 3229 19957
rect 3259 19901 3315 19957
rect 3345 19901 3401 19957
rect 3431 19901 3487 19957
rect 2915 19821 2971 19877
rect 3001 19821 3057 19877
rect 3087 19821 3143 19877
rect 3173 19821 3229 19877
rect 3259 19821 3315 19877
rect 3345 19821 3401 19877
rect 3431 19821 3487 19877
rect 2915 19741 2971 19797
rect 3001 19741 3057 19797
rect 3087 19741 3143 19797
rect 3173 19741 3229 19797
rect 3259 19741 3315 19797
rect 3345 19741 3401 19797
rect 3431 19741 3487 19797
rect 2915 19661 2971 19717
rect 3001 19661 3057 19717
rect 3087 19661 3143 19717
rect 3173 19661 3229 19717
rect 3259 19661 3315 19717
rect 3345 19661 3401 19717
rect 3431 19661 3487 19717
rect 2915 19581 2971 19637
rect 3001 19581 3057 19637
rect 3087 19581 3143 19637
rect 3173 19581 3229 19637
rect 3259 19581 3315 19637
rect 3345 19581 3401 19637
rect 3431 19581 3487 19637
rect 2915 19501 2971 19557
rect 3001 19501 3057 19557
rect 3087 19501 3143 19557
rect 3173 19501 3229 19557
rect 3259 19501 3315 19557
rect 3345 19501 3401 19557
rect 3431 19501 3487 19557
rect 2915 19421 2971 19477
rect 3001 19421 3057 19477
rect 3087 19421 3143 19477
rect 3173 19421 3229 19477
rect 3259 19421 3315 19477
rect 3345 19421 3401 19477
rect 3431 19421 3487 19477
rect 2915 19341 2971 19397
rect 3001 19341 3057 19397
rect 3087 19341 3143 19397
rect 3173 19341 3229 19397
rect 3259 19341 3315 19397
rect 3345 19341 3401 19397
rect 3431 19341 3487 19397
rect 2915 19261 2971 19317
rect 3001 19261 3057 19317
rect 3087 19261 3143 19317
rect 3173 19261 3229 19317
rect 3259 19261 3315 19317
rect 3345 19261 3401 19317
rect 3431 19261 3487 19317
rect 5903 21261 5959 21317
rect 5989 21261 6045 21317
rect 6075 21261 6131 21317
rect 6161 21261 6217 21317
rect 6247 21261 6303 21317
rect 6333 21261 6389 21317
rect 6419 21261 6475 21317
rect 5903 21181 5959 21237
rect 5989 21181 6045 21237
rect 6075 21181 6131 21237
rect 6161 21181 6217 21237
rect 6247 21181 6303 21237
rect 6333 21181 6389 21237
rect 6419 21181 6475 21237
rect 5903 21101 5959 21157
rect 5989 21101 6045 21157
rect 6075 21101 6131 21157
rect 6161 21101 6217 21157
rect 6247 21101 6303 21157
rect 6333 21101 6389 21157
rect 6419 21101 6475 21157
rect 5903 21021 5959 21077
rect 5989 21021 6045 21077
rect 6075 21021 6131 21077
rect 6161 21021 6217 21077
rect 6247 21021 6303 21077
rect 6333 21021 6389 21077
rect 6419 21021 6475 21077
rect 5903 20941 5959 20997
rect 5989 20941 6045 20997
rect 6075 20941 6131 20997
rect 6161 20941 6217 20997
rect 6247 20941 6303 20997
rect 6333 20941 6389 20997
rect 6419 20941 6475 20997
rect 5903 20861 5959 20917
rect 5989 20861 6045 20917
rect 6075 20861 6131 20917
rect 6161 20861 6217 20917
rect 6247 20861 6303 20917
rect 6333 20861 6389 20917
rect 6419 20861 6475 20917
rect 5903 20781 5959 20837
rect 5989 20781 6045 20837
rect 6075 20781 6131 20837
rect 6161 20781 6217 20837
rect 6247 20781 6303 20837
rect 6333 20781 6389 20837
rect 6419 20781 6475 20837
rect 5903 20701 5959 20757
rect 5989 20701 6045 20757
rect 6075 20701 6131 20757
rect 6161 20701 6217 20757
rect 6247 20701 6303 20757
rect 6333 20701 6389 20757
rect 6419 20701 6475 20757
rect 5903 20621 5959 20677
rect 5989 20621 6045 20677
rect 6075 20621 6131 20677
rect 6161 20621 6217 20677
rect 6247 20621 6303 20677
rect 6333 20621 6389 20677
rect 6419 20621 6475 20677
rect 5903 20541 5959 20597
rect 5989 20541 6045 20597
rect 6075 20541 6131 20597
rect 6161 20541 6217 20597
rect 6247 20541 6303 20597
rect 6333 20541 6389 20597
rect 6419 20541 6475 20597
rect 5903 20461 5959 20517
rect 5989 20461 6045 20517
rect 6075 20461 6131 20517
rect 6161 20461 6217 20517
rect 6247 20461 6303 20517
rect 6333 20461 6389 20517
rect 6419 20461 6475 20517
rect 5903 20381 5959 20437
rect 5989 20381 6045 20437
rect 6075 20381 6131 20437
rect 6161 20381 6217 20437
rect 6247 20381 6303 20437
rect 6333 20381 6389 20437
rect 6419 20381 6475 20437
rect 5903 20301 5959 20357
rect 5989 20301 6045 20357
rect 6075 20301 6131 20357
rect 6161 20301 6217 20357
rect 6247 20301 6303 20357
rect 6333 20301 6389 20357
rect 6419 20301 6475 20357
rect 5903 20221 5959 20277
rect 5989 20221 6045 20277
rect 6075 20221 6131 20277
rect 6161 20221 6217 20277
rect 6247 20221 6303 20277
rect 6333 20221 6389 20277
rect 6419 20221 6475 20277
rect 5903 20141 5959 20197
rect 5989 20141 6045 20197
rect 6075 20141 6131 20197
rect 6161 20141 6217 20197
rect 6247 20141 6303 20197
rect 6333 20141 6389 20197
rect 6419 20141 6475 20197
rect 5903 20061 5959 20117
rect 5989 20061 6045 20117
rect 6075 20061 6131 20117
rect 6161 20061 6217 20117
rect 6247 20061 6303 20117
rect 6333 20061 6389 20117
rect 6419 20061 6475 20117
rect 5903 19981 5959 20037
rect 5989 19981 6045 20037
rect 6075 19981 6131 20037
rect 6161 19981 6217 20037
rect 6247 19981 6303 20037
rect 6333 19981 6389 20037
rect 6419 19981 6475 20037
rect 5903 19901 5959 19957
rect 5989 19901 6045 19957
rect 6075 19901 6131 19957
rect 6161 19901 6217 19957
rect 6247 19901 6303 19957
rect 6333 19901 6389 19957
rect 6419 19901 6475 19957
rect 5903 19821 5959 19877
rect 5989 19821 6045 19877
rect 6075 19821 6131 19877
rect 6161 19821 6217 19877
rect 6247 19821 6303 19877
rect 6333 19821 6389 19877
rect 6419 19821 6475 19877
rect 5903 19741 5959 19797
rect 5989 19741 6045 19797
rect 6075 19741 6131 19797
rect 6161 19741 6217 19797
rect 6247 19741 6303 19797
rect 6333 19741 6389 19797
rect 6419 19741 6475 19797
rect 5903 19661 5959 19717
rect 5989 19661 6045 19717
rect 6075 19661 6131 19717
rect 6161 19661 6217 19717
rect 6247 19661 6303 19717
rect 6333 19661 6389 19717
rect 6419 19661 6475 19717
rect 5903 19581 5959 19637
rect 5989 19581 6045 19637
rect 6075 19581 6131 19637
rect 6161 19581 6217 19637
rect 6247 19581 6303 19637
rect 6333 19581 6389 19637
rect 6419 19581 6475 19637
rect 5903 19501 5959 19557
rect 5989 19501 6045 19557
rect 6075 19501 6131 19557
rect 6161 19501 6217 19557
rect 6247 19501 6303 19557
rect 6333 19501 6389 19557
rect 6419 19501 6475 19557
rect 5903 19421 5959 19477
rect 5989 19421 6045 19477
rect 6075 19421 6131 19477
rect 6161 19421 6217 19477
rect 6247 19421 6303 19477
rect 6333 19421 6389 19477
rect 6419 19421 6475 19477
rect 5903 19341 5959 19397
rect 5989 19341 6045 19397
rect 6075 19341 6131 19397
rect 6161 19341 6217 19397
rect 6247 19341 6303 19397
rect 6333 19341 6389 19397
rect 6419 19341 6475 19397
rect 5903 19261 5959 19317
rect 5989 19261 6045 19317
rect 6075 19261 6131 19317
rect 6161 19261 6217 19317
rect 6247 19261 6303 19317
rect 6333 19261 6389 19317
rect 6419 19261 6475 19317
rect 5007 18602 5056 18623
rect 5056 18602 5063 18623
rect 5133 18602 5140 18623
rect 5140 18602 5189 18623
rect 5007 18588 5063 18602
rect 5133 18588 5189 18602
rect 5007 18567 5056 18588
rect 5056 18567 5063 18588
rect 5133 18567 5140 18588
rect 5140 18567 5189 18588
rect 1660 17711 1716 17767
rect 2526 17711 2582 17767
rect 2739 17711 2795 17767
rect 3605 17711 3661 17767
rect 5728 17711 5784 17767
rect 6594 17711 6650 17767
rect 6807 17711 6863 17767
rect 7673 17711 7729 17767
rect 7843 17689 7899 17745
rect 7949 17689 8005 17745
rect 8054 17689 8110 17745
rect 8159 17689 8215 17745
rect 8264 17689 8320 17745
rect 8369 17689 8425 17745
rect 1660 17624 1716 17680
rect 2526 17624 2582 17680
rect 2739 17624 2795 17680
rect 3605 17624 3661 17680
rect 5728 17624 5784 17680
rect 6594 17624 6650 17680
rect 6807 17624 6863 17680
rect 7673 17624 7729 17680
rect 1660 17537 1716 17593
rect 2526 17537 2582 17593
rect 2739 17537 2795 17593
rect 3605 17537 3661 17593
rect 5728 17537 5784 17593
rect 6594 17537 6650 17593
rect 6807 17537 6863 17593
rect 7673 17537 7729 17593
rect 7843 17589 7899 17645
rect 7949 17589 8005 17645
rect 8054 17589 8110 17645
rect 8159 17589 8215 17645
rect 8264 17589 8320 17645
rect 8369 17589 8425 17645
rect 1660 17449 1716 17505
rect 2526 17449 2582 17505
rect 2739 17449 2795 17505
rect 3605 17449 3661 17505
rect 5728 17449 5784 17505
rect 6594 17449 6650 17505
rect 6807 17449 6863 17505
rect 7673 17449 7729 17505
rect 7843 17489 7899 17545
rect 7949 17489 8005 17545
rect 8054 17489 8110 17545
rect 8159 17489 8215 17545
rect 8264 17489 8320 17545
rect 8369 17489 8425 17545
rect 1660 17361 1716 17417
rect 2526 17361 2582 17417
rect 2739 17361 2795 17417
rect 3605 17361 3661 17417
rect 5728 17361 5784 17417
rect 6594 17361 6650 17417
rect 6807 17361 6863 17417
rect 7673 17361 7729 17417
rect 7843 17389 7899 17445
rect 7949 17389 8005 17445
rect 8054 17389 8110 17445
rect 8159 17389 8215 17445
rect 8264 17389 8320 17445
rect 8369 17389 8425 17445
rect 1660 17273 1716 17329
rect 2526 17273 2582 17329
rect 2739 17273 2795 17329
rect 3605 17273 3661 17329
rect 5728 17273 5784 17329
rect 6594 17273 6650 17329
rect 6807 17273 6863 17329
rect 7673 17273 7729 17329
rect 7843 17289 7899 17345
rect 7949 17289 8005 17345
rect 8054 17289 8110 17345
rect 8159 17289 8215 17345
rect 8264 17289 8320 17345
rect 8369 17289 8425 17345
rect 1660 17185 1716 17241
rect 2526 17185 2582 17241
rect 2739 17185 2795 17241
rect 3605 17185 3661 17241
rect 5728 17185 5784 17241
rect 6594 17185 6650 17241
rect 6807 17185 6863 17241
rect 7673 17185 7729 17241
rect 7843 17189 7899 17245
rect 7949 17189 8005 17245
rect 8054 17189 8110 17245
rect 8159 17189 8215 17245
rect 8264 17189 8320 17245
rect 8369 17189 8425 17245
rect 5003 16429 5004 16481
rect 5004 16429 5056 16481
rect 5056 16429 5059 16481
rect 5137 16429 5140 16481
rect 5140 16429 5192 16481
rect 5192 16429 5193 16481
rect 5003 16425 5059 16429
rect 5137 16425 5193 16429
rect 7843 15823 7899 15879
rect 7949 15823 8005 15879
rect 8054 15823 8110 15879
rect 8159 15823 8215 15879
rect 8264 15823 8320 15879
rect 8369 15823 8425 15879
rect 7843 15679 7899 15735
rect 7949 15679 8005 15735
rect 8054 15679 8110 15735
rect 8159 15679 8215 15735
rect 8264 15679 8320 15735
rect 8369 15679 8425 15735
rect 4425 15514 4474 15566
rect 4474 15514 4481 15566
rect 4551 15514 4558 15566
rect 4558 15514 4607 15566
rect 4425 15510 4481 15514
rect 4551 15510 4607 15514
rect 4425 15482 4481 15486
rect 4551 15482 4607 15486
rect 4425 15430 4474 15482
rect 4474 15430 4481 15482
rect 4551 15430 4558 15482
rect 4558 15430 4607 15482
rect 963 14628 1019 14684
rect 1069 14628 1125 14684
rect 1174 14628 1230 14684
rect 1279 14628 1335 14684
rect 1384 14628 1440 14684
rect 1489 14628 1545 14684
rect 963 14484 1019 14540
rect 1069 14484 1125 14540
rect 1174 14484 1230 14540
rect 1279 14484 1335 14540
rect 1384 14484 1440 14540
rect 1489 14484 1545 14540
rect 4425 14371 4474 14423
rect 4474 14371 4481 14423
rect 4551 14371 4558 14423
rect 4558 14371 4607 14423
rect 4425 14367 4481 14371
rect 4551 14367 4607 14371
rect 4425 14339 4481 14343
rect 4551 14339 4607 14343
rect 4425 14287 4474 14339
rect 4474 14287 4481 14339
rect 4551 14287 4558 14339
rect 4558 14287 4607 14339
rect 7843 14104 7899 14160
rect 7949 14104 8005 14160
rect 8054 14104 8110 14160
rect 8159 14104 8215 14160
rect 8264 14104 8320 14160
rect 8369 14104 8425 14160
rect 7843 13960 7899 14016
rect 7949 13960 8005 14016
rect 8054 13960 8110 14016
rect 8159 13960 8215 14016
rect 8264 13960 8320 14016
rect 8369 13960 8425 14016
rect 462 13739 518 13795
rect 571 13739 627 13795
rect 680 13739 736 13795
rect 788 13739 844 13795
rect 462 13595 518 13651
rect 571 13595 627 13651
rect 680 13595 736 13651
rect 788 13595 844 13651
rect 7843 13382 7899 13438
rect 7949 13382 8005 13438
rect 8054 13382 8110 13438
rect 8159 13382 8215 13438
rect 8264 13382 8320 13438
rect 8369 13382 8425 13438
rect 7843 13238 7899 13294
rect 7949 13238 8005 13294
rect 8054 13238 8110 13294
rect 8159 13238 8215 13294
rect 8264 13238 8320 13294
rect 8369 13238 8425 13294
rect 4425 12990 4474 13042
rect 4474 12990 4481 13042
rect 4551 12990 4558 13042
rect 4558 12990 4607 13042
rect 4425 12986 4481 12990
rect 4551 12986 4607 12990
rect 4425 12958 4481 12962
rect 4551 12958 4607 12962
rect 4425 12906 4474 12958
rect 4474 12906 4481 12958
rect 4551 12906 4558 12958
rect 4558 12906 4607 12958
rect 963 12802 1019 12858
rect 1069 12802 1125 12858
rect 1174 12802 1230 12858
rect 1279 12802 1335 12858
rect 1384 12802 1440 12858
rect 1489 12802 1545 12858
rect 963 12658 1019 12714
rect 1069 12658 1125 12714
rect 1174 12658 1230 12714
rect 1279 12658 1335 12714
rect 1384 12658 1440 12714
rect 1489 12658 1545 12714
rect 4425 11857 4474 11909
rect 4474 11857 4481 11909
rect 4551 11857 4558 11909
rect 4558 11857 4607 11909
rect 4425 11853 4481 11857
rect 4551 11853 4607 11857
rect 4425 11825 4481 11829
rect 4551 11825 4607 11829
rect 4425 11773 4474 11825
rect 4474 11773 4481 11825
rect 4551 11773 4558 11825
rect 4558 11773 4607 11825
rect 7843 11583 7899 11639
rect 7949 11583 8005 11639
rect 8054 11583 8110 11639
rect 8159 11583 8215 11639
rect 8264 11583 8320 11639
rect 8369 11583 8425 11639
rect 4436 11409 4485 11461
rect 4485 11409 4492 11461
rect 4436 11405 4492 11409
rect 4551 11409 4558 11461
rect 4558 11409 4607 11461
rect 7843 11439 7899 11495
rect 7949 11439 8005 11495
rect 8054 11439 8110 11495
rect 8159 11439 8215 11495
rect 8264 11439 8320 11495
rect 8369 11439 8425 11495
rect 4551 11405 4607 11409
rect 4436 11377 4492 11381
rect 4436 11325 4485 11377
rect 4485 11325 4492 11377
rect 4551 11377 4607 11381
rect 4551 11325 4558 11377
rect 4558 11325 4607 11377
rect 7843 10895 7899 10951
rect 7949 10895 8005 10951
rect 8054 10895 8110 10951
rect 8159 10895 8215 10951
rect 8264 10895 8320 10951
rect 8369 10895 8425 10951
rect 7843 10751 7899 10807
rect 7949 10751 8005 10807
rect 8054 10751 8110 10807
rect 8159 10751 8215 10807
rect 8264 10751 8320 10807
rect 8369 10751 8425 10807
rect 4425 10459 4474 10511
rect 4474 10459 4481 10511
rect 4551 10459 4558 10511
rect 4558 10459 4607 10511
rect 4425 10455 4481 10459
rect 4551 10455 4607 10459
rect 4425 10427 4481 10431
rect 4551 10427 4607 10431
rect 4425 10375 4474 10427
rect 4474 10375 4481 10427
rect 4551 10375 4558 10427
rect 4558 10375 4607 10427
rect 963 9580 1019 9636
rect 1069 9580 1125 9636
rect 1174 9580 1230 9636
rect 1279 9580 1335 9636
rect 1384 9580 1440 9636
rect 1489 9580 1545 9636
rect 963 9436 1019 9492
rect 1069 9436 1125 9492
rect 1174 9436 1230 9492
rect 1279 9436 1335 9492
rect 1384 9436 1440 9492
rect 1489 9436 1545 9492
rect 4425 9337 4474 9389
rect 4474 9337 4481 9389
rect 4551 9337 4558 9389
rect 4558 9337 4607 9389
rect 4425 9333 4481 9337
rect 4551 9333 4607 9337
rect 4425 9305 4481 9309
rect 4551 9305 4607 9309
rect 4425 9253 4474 9305
rect 4474 9253 4481 9305
rect 4551 9253 4558 9305
rect 4558 9253 4607 9305
rect 320 9189 367 9238
rect 367 9189 376 9238
rect 320 9182 376 9189
rect 320 9123 367 9153
rect 367 9123 376 9153
rect 320 9109 376 9123
rect 320 9097 367 9109
rect 367 9097 376 9109
rect 320 9057 367 9068
rect 367 9057 376 9068
rect 320 9043 376 9057
rect 320 9012 367 9043
rect 367 9012 376 9043
rect 320 8977 376 8983
rect 320 8927 367 8977
rect 367 8927 376 8977
rect 320 8859 367 8898
rect 367 8859 376 8898
rect 320 8844 376 8859
rect 320 8842 367 8844
rect 367 8842 376 8844
rect 320 8792 367 8812
rect 367 8792 376 8812
rect 320 8777 376 8792
rect 320 8756 367 8777
rect 367 8756 376 8777
rect 320 8725 367 8726
rect 367 8725 376 8726
rect 2084 9189 2085 9238
rect 2085 9189 2137 9238
rect 2137 9189 2140 9238
rect 2198 9189 2223 9238
rect 2223 9189 2254 9238
rect 2312 9189 2343 9238
rect 2343 9189 2368 9238
rect 2426 9189 2429 9238
rect 2429 9189 2481 9238
rect 2481 9189 2482 9238
rect 2084 9182 2140 9189
rect 2198 9182 2254 9189
rect 2312 9182 2368 9189
rect 2426 9182 2482 9189
rect 2084 9079 2140 9106
rect 2198 9079 2254 9106
rect 2312 9079 2368 9106
rect 2426 9079 2482 9106
rect 2084 9050 2085 9079
rect 2085 9050 2137 9079
rect 2137 9050 2140 9079
rect 2198 9050 2223 9079
rect 2223 9050 2254 9079
rect 2312 9050 2343 9079
rect 2343 9050 2368 9079
rect 2426 9050 2429 9079
rect 2429 9050 2481 9079
rect 2481 9050 2482 9079
rect 7843 9149 7899 9205
rect 7949 9149 8005 9205
rect 8054 9149 8110 9205
rect 8159 9149 8215 9205
rect 8264 9149 8320 9205
rect 8369 9149 8425 9205
rect 7843 9005 7899 9061
rect 7949 9005 8005 9061
rect 8054 9005 8110 9061
rect 8159 9005 8215 9061
rect 8264 9005 8320 9061
rect 8369 9005 8425 9061
rect 8532 9189 8534 9238
rect 8534 9189 8586 9238
rect 8586 9189 8588 9238
rect 8612 9189 8650 9238
rect 8650 9189 8662 9238
rect 8662 9189 8668 9238
rect 8692 9189 8714 9238
rect 8714 9189 8726 9238
rect 8726 9189 8748 9238
rect 8772 9189 8778 9238
rect 8778 9189 8790 9238
rect 8790 9189 8828 9238
rect 8852 9189 8854 9238
rect 8854 9189 8906 9238
rect 8906 9189 8908 9238
rect 8932 9189 8970 9238
rect 8970 9189 8982 9238
rect 8982 9189 8988 9238
rect 9012 9189 9034 9238
rect 9034 9189 9046 9238
rect 9046 9189 9068 9238
rect 9092 9189 9098 9238
rect 9098 9189 9110 9238
rect 9110 9189 9148 9238
rect 9172 9189 9174 9238
rect 9174 9189 9226 9238
rect 9226 9189 9228 9238
rect 8532 9182 8588 9189
rect 8612 9182 8668 9189
rect 8692 9182 8748 9189
rect 8772 9182 8828 9189
rect 8852 9182 8908 9189
rect 8932 9182 8988 9189
rect 9012 9182 9068 9189
rect 9092 9182 9148 9189
rect 9172 9182 9228 9189
rect 8532 9123 8534 9153
rect 8534 9123 8586 9153
rect 8586 9123 8588 9153
rect 8612 9123 8650 9153
rect 8650 9123 8662 9153
rect 8662 9123 8668 9153
rect 8692 9123 8714 9153
rect 8714 9123 8726 9153
rect 8726 9123 8748 9153
rect 8772 9123 8778 9153
rect 8778 9123 8790 9153
rect 8790 9123 8828 9153
rect 8852 9123 8854 9153
rect 8854 9123 8906 9153
rect 8906 9123 8908 9153
rect 8932 9123 8970 9153
rect 8970 9123 8982 9153
rect 8982 9123 8988 9153
rect 9012 9123 9034 9153
rect 9034 9123 9046 9153
rect 9046 9123 9068 9153
rect 9092 9123 9098 9153
rect 9098 9123 9110 9153
rect 9110 9123 9148 9153
rect 9172 9123 9174 9153
rect 9174 9123 9226 9153
rect 9226 9123 9228 9153
rect 8532 9109 8588 9123
rect 8612 9109 8668 9123
rect 8692 9109 8748 9123
rect 8772 9109 8828 9123
rect 8852 9109 8908 9123
rect 8932 9109 8988 9123
rect 9012 9109 9068 9123
rect 9092 9109 9148 9123
rect 9172 9109 9228 9123
rect 8532 9097 8534 9109
rect 8534 9097 8586 9109
rect 8586 9097 8588 9109
rect 8612 9097 8650 9109
rect 8650 9097 8662 9109
rect 8662 9097 8668 9109
rect 8692 9097 8714 9109
rect 8714 9097 8726 9109
rect 8726 9097 8748 9109
rect 8772 9097 8778 9109
rect 8778 9097 8790 9109
rect 8790 9097 8828 9109
rect 8852 9097 8854 9109
rect 8854 9097 8906 9109
rect 8906 9097 8908 9109
rect 8932 9097 8970 9109
rect 8970 9097 8982 9109
rect 8982 9097 8988 9109
rect 9012 9097 9034 9109
rect 9034 9097 9046 9109
rect 9046 9097 9068 9109
rect 9092 9097 9098 9109
rect 9098 9097 9110 9109
rect 9110 9097 9148 9109
rect 9172 9097 9174 9109
rect 9174 9097 9226 9109
rect 9226 9097 9228 9109
rect 8532 9057 8534 9068
rect 8534 9057 8586 9068
rect 8586 9057 8588 9068
rect 8612 9057 8650 9068
rect 8650 9057 8662 9068
rect 8662 9057 8668 9068
rect 8692 9057 8714 9068
rect 8714 9057 8726 9068
rect 8726 9057 8748 9068
rect 8772 9057 8778 9068
rect 8778 9057 8790 9068
rect 8790 9057 8828 9068
rect 8852 9057 8854 9068
rect 8854 9057 8906 9068
rect 8906 9057 8908 9068
rect 8932 9057 8970 9068
rect 8970 9057 8982 9068
rect 8982 9057 8988 9068
rect 9012 9057 9034 9068
rect 9034 9057 9046 9068
rect 9046 9057 9068 9068
rect 9092 9057 9098 9068
rect 9098 9057 9110 9068
rect 9110 9057 9148 9068
rect 9172 9057 9174 9068
rect 9174 9057 9226 9068
rect 9226 9057 9228 9068
rect 8532 9043 8588 9057
rect 8612 9043 8668 9057
rect 8692 9043 8748 9057
rect 8772 9043 8828 9057
rect 8852 9043 8908 9057
rect 8932 9043 8988 9057
rect 9012 9043 9068 9057
rect 9092 9043 9148 9057
rect 9172 9043 9228 9057
rect 8532 9012 8534 9043
rect 8534 9012 8586 9043
rect 8586 9012 8588 9043
rect 8612 9012 8650 9043
rect 8650 9012 8662 9043
rect 8662 9012 8668 9043
rect 8692 9012 8714 9043
rect 8714 9012 8726 9043
rect 8726 9012 8748 9043
rect 8772 9012 8778 9043
rect 8778 9012 8790 9043
rect 8790 9012 8828 9043
rect 8852 9012 8854 9043
rect 8854 9012 8906 9043
rect 8906 9012 8908 9043
rect 8932 9012 8970 9043
rect 8970 9012 8982 9043
rect 8982 9012 8988 9043
rect 9012 9012 9034 9043
rect 9034 9012 9046 9043
rect 9046 9012 9068 9043
rect 9092 9012 9098 9043
rect 9098 9012 9110 9043
rect 9110 9012 9148 9043
rect 9172 9012 9174 9043
rect 9174 9012 9226 9043
rect 9226 9012 9228 9043
rect 2084 8945 2085 8973
rect 2085 8945 2137 8973
rect 2137 8945 2140 8973
rect 2198 8945 2223 8973
rect 2223 8945 2254 8973
rect 2312 8945 2343 8973
rect 2343 8945 2368 8973
rect 2426 8945 2429 8973
rect 2429 8945 2481 8973
rect 2481 8945 2482 8973
rect 2084 8917 2140 8945
rect 2198 8917 2254 8945
rect 2312 8917 2368 8945
rect 2426 8917 2482 8945
rect 2084 8833 2140 8840
rect 2198 8833 2254 8840
rect 2312 8833 2368 8840
rect 2426 8833 2482 8840
rect 2084 8784 2085 8833
rect 2085 8784 2137 8833
rect 2137 8784 2140 8833
rect 2198 8784 2223 8833
rect 2223 8784 2254 8833
rect 2312 8784 2343 8833
rect 2343 8784 2368 8833
rect 2426 8784 2429 8833
rect 2429 8784 2481 8833
rect 2481 8784 2482 8833
rect 8532 8977 8588 8983
rect 8612 8977 8668 8983
rect 8692 8977 8748 8983
rect 8772 8977 8828 8983
rect 8852 8977 8908 8983
rect 8932 8977 8988 8983
rect 9012 8977 9068 8983
rect 9092 8977 9148 8983
rect 9172 8977 9228 8983
rect 8532 8927 8534 8977
rect 8534 8927 8586 8977
rect 8586 8927 8588 8977
rect 8612 8927 8650 8977
rect 8650 8927 8662 8977
rect 8662 8927 8668 8977
rect 8692 8927 8714 8977
rect 8714 8927 8726 8977
rect 8726 8927 8748 8977
rect 8772 8927 8778 8977
rect 8778 8927 8790 8977
rect 8790 8927 8828 8977
rect 8852 8927 8854 8977
rect 8854 8927 8906 8977
rect 8906 8927 8908 8977
rect 8932 8927 8970 8977
rect 8970 8927 8982 8977
rect 8982 8927 8988 8977
rect 9012 8927 9034 8977
rect 9034 8927 9046 8977
rect 9046 8927 9068 8977
rect 9092 8927 9098 8977
rect 9098 8927 9110 8977
rect 9110 8927 9148 8977
rect 9172 8927 9174 8977
rect 9174 8927 9226 8977
rect 9226 8927 9228 8977
rect 8532 8859 8534 8898
rect 8534 8859 8586 8898
rect 8586 8859 8588 8898
rect 8612 8859 8650 8898
rect 8650 8859 8662 8898
rect 8662 8859 8668 8898
rect 8692 8859 8714 8898
rect 8714 8859 8726 8898
rect 8726 8859 8748 8898
rect 8772 8859 8778 8898
rect 8778 8859 8790 8898
rect 8790 8859 8828 8898
rect 8852 8859 8854 8898
rect 8854 8859 8906 8898
rect 8906 8859 8908 8898
rect 8932 8859 8970 8898
rect 8970 8859 8982 8898
rect 8982 8859 8988 8898
rect 9012 8859 9034 8898
rect 9034 8859 9046 8898
rect 9046 8859 9068 8898
rect 9092 8859 9098 8898
rect 9098 8859 9110 8898
rect 9110 8859 9148 8898
rect 9172 8859 9174 8898
rect 9174 8859 9226 8898
rect 9226 8859 9228 8898
rect 8532 8844 8588 8859
rect 8612 8844 8668 8859
rect 8692 8844 8748 8859
rect 8772 8844 8828 8859
rect 8852 8844 8908 8859
rect 8932 8844 8988 8859
rect 9012 8844 9068 8859
rect 9092 8844 9148 8859
rect 9172 8844 9228 8859
rect 8532 8842 8534 8844
rect 8534 8842 8586 8844
rect 8586 8842 8588 8844
rect 8612 8842 8650 8844
rect 8650 8842 8662 8844
rect 8662 8842 8668 8844
rect 8692 8842 8714 8844
rect 8714 8842 8726 8844
rect 8726 8842 8748 8844
rect 8772 8842 8778 8844
rect 8778 8842 8790 8844
rect 8790 8842 8828 8844
rect 8852 8842 8854 8844
rect 8854 8842 8906 8844
rect 8906 8842 8908 8844
rect 8932 8842 8970 8844
rect 8970 8842 8982 8844
rect 8982 8842 8988 8844
rect 9012 8842 9034 8844
rect 9034 8842 9046 8844
rect 9046 8842 9068 8844
rect 9092 8842 9098 8844
rect 9098 8842 9110 8844
rect 9110 8842 9148 8844
rect 9172 8842 9174 8844
rect 9174 8842 9226 8844
rect 9226 8842 9228 8844
rect 8532 8792 8534 8812
rect 8534 8792 8586 8812
rect 8586 8792 8588 8812
rect 8612 8792 8650 8812
rect 8650 8792 8662 8812
rect 8662 8792 8668 8812
rect 8692 8792 8714 8812
rect 8714 8792 8726 8812
rect 8726 8792 8748 8812
rect 8772 8792 8778 8812
rect 8778 8792 8790 8812
rect 8790 8792 8828 8812
rect 8852 8792 8854 8812
rect 8854 8792 8906 8812
rect 8906 8792 8908 8812
rect 8932 8792 8970 8812
rect 8970 8792 8982 8812
rect 8982 8792 8988 8812
rect 9012 8792 9034 8812
rect 9034 8792 9046 8812
rect 9046 8792 9068 8812
rect 9092 8792 9098 8812
rect 9098 8792 9110 8812
rect 9110 8792 9148 8812
rect 9172 8792 9174 8812
rect 9174 8792 9226 8812
rect 9226 8792 9228 8812
rect 8532 8777 8588 8792
rect 8612 8777 8668 8792
rect 8692 8777 8748 8792
rect 8772 8777 8828 8792
rect 8852 8777 8908 8792
rect 8932 8777 8988 8792
rect 9012 8777 9068 8792
rect 9092 8777 9148 8792
rect 9172 8777 9228 8792
rect 320 8710 376 8725
rect 8532 8756 8534 8777
rect 8534 8756 8586 8777
rect 8586 8756 8588 8777
rect 8612 8756 8650 8777
rect 8650 8756 8662 8777
rect 8662 8756 8668 8777
rect 8692 8756 8714 8777
rect 8714 8756 8726 8777
rect 8726 8756 8748 8777
rect 8772 8756 8778 8777
rect 8778 8756 8790 8777
rect 8790 8756 8828 8777
rect 8852 8756 8854 8777
rect 8854 8756 8906 8777
rect 8906 8756 8908 8777
rect 8932 8756 8970 8777
rect 8970 8756 8982 8777
rect 8982 8756 8988 8777
rect 9012 8756 9034 8777
rect 9034 8756 9046 8777
rect 9046 8756 9068 8777
rect 9092 8756 9098 8777
rect 9098 8756 9110 8777
rect 9110 8756 9148 8777
rect 9172 8756 9174 8777
rect 9174 8756 9226 8777
rect 9226 8756 9228 8777
rect 8532 8725 8534 8726
rect 8534 8725 8586 8726
rect 8586 8725 8588 8726
rect 8612 8725 8650 8726
rect 8650 8725 8662 8726
rect 8662 8725 8668 8726
rect 8692 8725 8714 8726
rect 8714 8725 8726 8726
rect 8726 8725 8748 8726
rect 8772 8725 8778 8726
rect 8778 8725 8790 8726
rect 8790 8725 8828 8726
rect 8852 8725 8854 8726
rect 8854 8725 8906 8726
rect 8906 8725 8908 8726
rect 8932 8725 8970 8726
rect 8970 8725 8982 8726
rect 8982 8725 8988 8726
rect 9012 8725 9034 8726
rect 9034 8725 9046 8726
rect 9046 8725 9068 8726
rect 9092 8725 9098 8726
rect 9098 8725 9110 8726
rect 9110 8725 9148 8726
rect 9172 8725 9174 8726
rect 9174 8725 9226 8726
rect 9226 8725 9228 8726
rect 320 8670 367 8710
rect 367 8670 376 8710
rect 320 8591 367 8640
rect 367 8591 376 8640
rect 320 8584 376 8591
rect 320 8524 367 8554
rect 367 8524 376 8554
rect 320 8509 376 8524
rect 476 8660 532 8716
rect 580 8660 636 8716
rect 684 8660 740 8716
rect 788 8660 844 8716
rect 476 8516 532 8572
rect 580 8516 636 8572
rect 684 8516 740 8572
rect 788 8516 844 8572
rect 8532 8710 8588 8725
rect 8612 8710 8668 8725
rect 8692 8710 8748 8725
rect 8772 8710 8828 8725
rect 8852 8710 8908 8725
rect 8932 8710 8988 8725
rect 9012 8710 9068 8725
rect 9092 8710 9148 8725
rect 9172 8710 9228 8725
rect 8532 8670 8534 8710
rect 8534 8670 8586 8710
rect 8586 8670 8588 8710
rect 8612 8670 8650 8710
rect 8650 8670 8662 8710
rect 8662 8670 8668 8710
rect 8692 8670 8714 8710
rect 8714 8670 8726 8710
rect 8726 8670 8748 8710
rect 8772 8670 8778 8710
rect 8778 8670 8790 8710
rect 8790 8670 8828 8710
rect 8852 8670 8854 8710
rect 8854 8670 8906 8710
rect 8906 8670 8908 8710
rect 8932 8670 8970 8710
rect 8970 8670 8982 8710
rect 8982 8670 8988 8710
rect 9012 8670 9034 8710
rect 9034 8670 9046 8710
rect 9046 8670 9068 8710
rect 9092 8670 9098 8710
rect 9098 8670 9110 8710
rect 9110 8670 9148 8710
rect 9172 8670 9174 8710
rect 9174 8670 9226 8710
rect 9226 8670 9228 8710
rect 8532 8591 8534 8640
rect 8534 8591 8586 8640
rect 8586 8591 8588 8640
rect 8612 8591 8650 8640
rect 8650 8591 8662 8640
rect 8662 8591 8668 8640
rect 8692 8591 8714 8640
rect 8714 8591 8726 8640
rect 8726 8591 8748 8640
rect 8772 8591 8778 8640
rect 8778 8591 8790 8640
rect 8790 8591 8828 8640
rect 8852 8591 8854 8640
rect 8854 8591 8906 8640
rect 8906 8591 8908 8640
rect 8932 8591 8970 8640
rect 8970 8591 8982 8640
rect 8982 8591 8988 8640
rect 9012 8591 9034 8640
rect 9034 8591 9046 8640
rect 9046 8591 9068 8640
rect 9092 8591 9098 8640
rect 9098 8591 9110 8640
rect 9110 8591 9148 8640
rect 9172 8591 9174 8640
rect 9174 8591 9226 8640
rect 9226 8591 9228 8640
rect 8532 8584 8588 8591
rect 8612 8584 8668 8591
rect 8692 8584 8748 8591
rect 8772 8584 8828 8591
rect 8852 8584 8908 8591
rect 8932 8584 8988 8591
rect 9012 8584 9068 8591
rect 9092 8584 9148 8591
rect 9172 8584 9228 8591
rect 8532 8524 8534 8554
rect 8534 8524 8586 8554
rect 8586 8524 8588 8554
rect 8612 8524 8650 8554
rect 8650 8524 8662 8554
rect 8662 8524 8668 8554
rect 8692 8524 8714 8554
rect 8714 8524 8726 8554
rect 8726 8524 8748 8554
rect 8772 8524 8778 8554
rect 8778 8524 8790 8554
rect 8790 8524 8828 8554
rect 8852 8524 8854 8554
rect 8854 8524 8906 8554
rect 8906 8524 8908 8554
rect 8932 8524 8970 8554
rect 8970 8524 8982 8554
rect 8982 8524 8988 8554
rect 9012 8524 9034 8554
rect 9034 8524 9046 8554
rect 9046 8524 9068 8554
rect 9092 8524 9098 8554
rect 9098 8524 9110 8554
rect 9110 8524 9148 8554
rect 9172 8524 9174 8554
rect 9174 8524 9226 8554
rect 9226 8524 9228 8554
rect 320 8498 367 8509
rect 367 8498 376 8509
rect 320 8457 367 8468
rect 367 8457 376 8468
rect 320 8442 376 8457
rect 320 8412 367 8442
rect 367 8412 376 8442
rect 8532 8509 8588 8524
rect 8612 8509 8668 8524
rect 8692 8509 8748 8524
rect 8772 8509 8828 8524
rect 8852 8509 8908 8524
rect 8932 8509 8988 8524
rect 9012 8509 9068 8524
rect 9092 8509 9148 8524
rect 9172 8509 9228 8524
rect 8532 8498 8534 8509
rect 8534 8498 8586 8509
rect 8586 8498 8588 8509
rect 8612 8498 8650 8509
rect 8650 8498 8662 8509
rect 8662 8498 8668 8509
rect 8692 8498 8714 8509
rect 8714 8498 8726 8509
rect 8726 8498 8748 8509
rect 8772 8498 8778 8509
rect 8778 8498 8790 8509
rect 8790 8498 8828 8509
rect 8852 8498 8854 8509
rect 8854 8498 8906 8509
rect 8906 8498 8908 8509
rect 8932 8498 8970 8509
rect 8970 8498 8982 8509
rect 8982 8498 8988 8509
rect 9012 8498 9034 8509
rect 9034 8498 9046 8509
rect 9046 8498 9068 8509
rect 9092 8498 9098 8509
rect 9098 8498 9110 8509
rect 9110 8498 9148 8509
rect 9172 8498 9174 8509
rect 9174 8498 9226 8509
rect 9226 8498 9228 8509
rect 8532 8457 8534 8468
rect 8534 8457 8586 8468
rect 8586 8457 8588 8468
rect 8612 8457 8650 8468
rect 8650 8457 8662 8468
rect 8662 8457 8668 8468
rect 8692 8457 8714 8468
rect 8714 8457 8726 8468
rect 8726 8457 8748 8468
rect 8772 8457 8778 8468
rect 8778 8457 8790 8468
rect 8790 8457 8828 8468
rect 8852 8457 8854 8468
rect 8854 8457 8906 8468
rect 8906 8457 8908 8468
rect 8932 8457 8970 8468
rect 8970 8457 8982 8468
rect 8982 8457 8988 8468
rect 9012 8457 9034 8468
rect 9034 8457 9046 8468
rect 9046 8457 9068 8468
rect 9092 8457 9098 8468
rect 9098 8457 9110 8468
rect 9110 8457 9148 8468
rect 9172 8457 9174 8468
rect 9174 8457 9226 8468
rect 9226 8457 9228 8468
rect 8532 8442 8588 8457
rect 8612 8442 8668 8457
rect 8692 8442 8748 8457
rect 8772 8442 8828 8457
rect 8852 8442 8908 8457
rect 8932 8442 8988 8457
rect 9012 8442 9068 8457
rect 9092 8442 9148 8457
rect 9172 8442 9228 8457
rect 320 8375 376 8382
rect 320 8326 367 8375
rect 367 8326 376 8375
rect 7843 8380 7899 8436
rect 7949 8380 8005 8436
rect 8054 8380 8110 8436
rect 8159 8380 8215 8436
rect 8264 8380 8320 8436
rect 8369 8380 8425 8436
rect 8532 8412 8534 8442
rect 8534 8412 8586 8442
rect 8586 8412 8588 8442
rect 8612 8412 8650 8442
rect 8650 8412 8662 8442
rect 8662 8412 8668 8442
rect 8692 8412 8714 8442
rect 8714 8412 8726 8442
rect 8726 8412 8748 8442
rect 8772 8412 8778 8442
rect 8778 8412 8790 8442
rect 8790 8412 8828 8442
rect 8852 8412 8854 8442
rect 8854 8412 8906 8442
rect 8906 8412 8908 8442
rect 8932 8412 8970 8442
rect 8970 8412 8982 8442
rect 8982 8412 8988 8442
rect 9012 8412 9034 8442
rect 9034 8412 9046 8442
rect 9046 8412 9068 8442
rect 9092 8412 9098 8442
rect 9098 8412 9110 8442
rect 9110 8412 9148 8442
rect 9172 8412 9174 8442
rect 9174 8412 9226 8442
rect 9226 8412 9228 8442
rect 8532 8375 8588 8382
rect 8612 8375 8668 8382
rect 8692 8375 8748 8382
rect 8772 8375 8828 8382
rect 8852 8375 8908 8382
rect 8932 8375 8988 8382
rect 9012 8375 9068 8382
rect 9092 8375 9148 8382
rect 9172 8375 9228 8382
rect 8532 8326 8534 8375
rect 8534 8326 8586 8375
rect 8586 8326 8588 8375
rect 8612 8326 8650 8375
rect 8650 8326 8662 8375
rect 8662 8326 8668 8375
rect 8692 8326 8714 8375
rect 8714 8326 8726 8375
rect 8726 8326 8748 8375
rect 8772 8326 8778 8375
rect 8778 8326 8790 8375
rect 8790 8326 8828 8375
rect 8852 8326 8854 8375
rect 8854 8326 8906 8375
rect 8906 8326 8908 8375
rect 8932 8326 8970 8375
rect 8970 8326 8982 8375
rect 8982 8326 8988 8375
rect 9012 8326 9034 8375
rect 9034 8326 9046 8375
rect 9046 8326 9068 8375
rect 9092 8326 9098 8375
rect 9098 8326 9110 8375
rect 9110 8326 9148 8375
rect 9172 8326 9174 8375
rect 9174 8326 9226 8375
rect 9226 8326 9228 8375
rect 7843 8236 7899 8292
rect 7949 8236 8005 8292
rect 8054 8236 8110 8292
rect 8159 8236 8215 8292
rect 8264 8236 8320 8292
rect 8369 8236 8425 8292
rect 4425 7950 4474 8002
rect 4474 7950 4481 8002
rect 4551 7950 4558 8002
rect 4558 7950 4607 8002
rect 4425 7946 4481 7950
rect 4551 7946 4607 7950
rect 4425 7918 4481 7922
rect 4551 7918 4607 7922
rect 4425 7866 4474 7918
rect 4474 7866 4481 7918
rect 4551 7866 4558 7918
rect 4558 7866 4607 7918
rect 963 7754 1019 7810
rect 1069 7754 1125 7810
rect 1174 7754 1230 7810
rect 1279 7754 1335 7810
rect 1384 7754 1440 7810
rect 1489 7754 1545 7810
rect 963 7610 1019 7666
rect 1069 7610 1125 7666
rect 1174 7610 1230 7666
rect 1279 7610 1335 7666
rect 1384 7610 1440 7666
rect 1489 7610 1545 7666
rect 4425 6828 4474 6880
rect 4474 6828 4481 6880
rect 4551 6828 4558 6880
rect 4558 6828 4607 6880
rect 4425 6824 4481 6828
rect 4551 6824 4607 6828
rect 4425 6796 4481 6800
rect 4551 6796 4607 6800
rect 4425 6744 4474 6796
rect 4474 6744 4481 6796
rect 4551 6744 4558 6796
rect 4558 6744 4607 6796
rect 7843 6648 7899 6704
rect 7949 6648 8005 6704
rect 8054 6648 8110 6704
rect 8159 6648 8215 6704
rect 8264 6648 8320 6704
rect 8369 6648 8425 6704
rect 7843 6504 7899 6560
rect 7949 6504 8005 6560
rect 8054 6504 8110 6560
rect 8159 6504 8215 6560
rect 8264 6504 8320 6560
rect 8369 6504 8425 6560
rect 7843 5861 7899 5917
rect 7949 5861 8005 5917
rect 8054 5861 8110 5917
rect 8159 5861 8215 5917
rect 8264 5861 8320 5917
rect 8369 5861 8425 5917
rect 7843 5717 7899 5773
rect 7949 5717 8005 5773
rect 8054 5717 8110 5773
rect 8159 5717 8215 5773
rect 8264 5717 8320 5773
rect 8369 5717 8425 5773
rect 4425 5434 4474 5486
rect 4474 5434 4481 5486
rect 4551 5434 4558 5486
rect 4558 5434 4607 5486
rect 4425 5430 4481 5434
rect 4551 5430 4607 5434
rect 4425 5402 4481 5406
rect 4551 5402 4607 5406
rect 4425 5350 4474 5402
rect 4474 5350 4481 5402
rect 4551 5350 4558 5402
rect 4558 5350 4607 5402
rect 7843 4812 7899 4868
rect 7949 4812 8005 4868
rect 8054 4812 8110 4868
rect 8159 4812 8215 4868
rect 8264 4812 8320 4868
rect 8369 4812 8425 4868
rect 7843 4668 7899 4724
rect 7949 4668 8005 4724
rect 8054 4668 8110 4724
rect 8159 4668 8215 4724
rect 8264 4668 8320 4724
rect 8369 4668 8425 4724
rect 4425 4006 4474 4058
rect 4474 4006 4481 4058
rect 4551 4006 4558 4058
rect 4558 4006 4607 4058
rect 4425 4002 4481 4006
rect 4551 4002 4607 4006
rect 4425 3974 4481 3978
rect 4551 3974 4607 3978
rect 4425 3922 4474 3974
rect 4474 3922 4481 3974
rect 4551 3922 4558 3974
rect 4558 3922 4607 3974
rect 7843 3676 7899 3732
rect 7949 3676 8005 3732
rect 8054 3676 8110 3732
rect 8159 3676 8215 3732
rect 8264 3676 8320 3732
rect 8369 3676 8425 3732
rect 7843 3532 7899 3588
rect 7949 3532 8005 3588
rect 8054 3532 8110 3588
rect 8159 3532 8215 3588
rect 8264 3532 8320 3588
rect 8369 3532 8425 3588
rect 963 3261 1019 3317
rect 1069 3261 1125 3317
rect 1174 3261 1230 3317
rect 1279 3261 1335 3317
rect 1384 3261 1440 3317
rect 1489 3261 1545 3317
rect 963 3117 1019 3173
rect 1069 3117 1125 3173
rect 1174 3117 1230 3173
rect 1279 3117 1335 3173
rect 1384 3117 1440 3173
rect 1489 3117 1545 3173
rect 4452 3264 4468 3312
rect 4468 3264 4490 3312
rect 4490 3264 4508 3312
rect 4532 3264 4542 3312
rect 4542 3264 4564 3312
rect 4564 3264 4588 3312
rect 4452 3256 4508 3264
rect 4532 3256 4588 3264
rect 4452 3188 4508 3231
rect 4532 3188 4588 3231
rect 4452 3175 4468 3188
rect 4468 3175 4490 3188
rect 4490 3175 4508 3188
rect 4532 3175 4542 3188
rect 4542 3175 4564 3188
rect 4564 3175 4588 3188
rect 7843 3166 7899 3222
rect 7949 3166 8005 3222
rect 8054 3166 8110 3222
rect 8159 3166 8215 3222
rect 8264 3166 8320 3222
rect 8369 3166 8425 3222
rect 4452 3136 4468 3150
rect 4468 3136 4490 3150
rect 4490 3136 4508 3150
rect 4532 3136 4542 3150
rect 4542 3136 4564 3150
rect 4564 3136 4588 3150
rect 4452 3094 4508 3136
rect 4532 3094 4588 3136
rect 4452 3060 4508 3069
rect 4532 3060 4588 3069
rect 4452 3013 4468 3060
rect 4468 3013 4490 3060
rect 4490 3013 4508 3060
rect 4532 3013 4542 3060
rect 4542 3013 4564 3060
rect 4564 3013 4588 3060
rect 4452 2932 4508 2988
rect 4532 2932 4588 2988
rect 7843 3022 7899 3078
rect 7949 3022 8005 3078
rect 8054 3022 8110 3078
rect 8159 3022 8215 3078
rect 8264 3022 8320 3078
rect 8369 3022 8425 3078
rect 4452 2880 4468 2907
rect 4468 2880 4490 2907
rect 4490 2880 4508 2907
rect 4532 2880 4542 2907
rect 4542 2880 4564 2907
rect 4564 2880 4588 2907
rect 4452 2851 4508 2880
rect 4532 2851 4588 2880
rect 4452 2804 4508 2826
rect 4532 2804 4588 2826
rect 4452 2770 4468 2804
rect 4468 2770 4490 2804
rect 4490 2770 4508 2804
rect 4532 2770 4542 2804
rect 4542 2770 4564 2804
rect 4564 2770 4588 2804
rect 4452 2688 4508 2744
rect 4532 2688 4588 2744
rect 4452 2624 4468 2662
rect 4468 2624 4490 2662
rect 4490 2624 4508 2662
rect 4532 2624 4542 2662
rect 4542 2624 4564 2662
rect 4564 2624 4588 2662
rect 4452 2606 4508 2624
rect 4532 2606 4588 2624
rect 4452 2547 4508 2580
rect 4532 2547 4588 2580
rect 4452 2524 4468 2547
rect 4468 2524 4490 2547
rect 4490 2524 4508 2547
rect 4532 2524 4542 2547
rect 4542 2524 4564 2547
rect 4564 2524 4588 2547
rect 4452 2495 4468 2498
rect 4468 2495 4490 2498
rect 4490 2495 4508 2498
rect 4532 2495 4542 2498
rect 4542 2495 4564 2498
rect 4564 2495 4588 2498
rect 4452 2442 4508 2495
rect 4532 2442 4588 2495
rect 4452 2366 4468 2416
rect 4468 2366 4490 2416
rect 4490 2366 4508 2416
rect 4532 2366 4542 2416
rect 4542 2366 4564 2416
rect 4564 2366 4588 2416
rect 4452 2360 4508 2366
rect 4532 2360 4588 2366
rect 4452 2278 4508 2334
rect 4532 2278 4588 2334
rect 4452 2196 4508 2252
rect 4532 2196 4588 2252
rect 963 2133 1019 2189
rect 1069 2133 1125 2189
rect 1174 2133 1230 2189
rect 1279 2133 1335 2189
rect 1384 2133 1440 2189
rect 1489 2133 1545 2189
rect 963 2011 1019 2067
rect 1069 2011 1125 2067
rect 1174 2011 1230 2067
rect 1279 2011 1335 2067
rect 1384 2011 1440 2067
rect 1489 2011 1545 2067
rect 963 1889 1019 1945
rect 1069 1889 1125 1945
rect 1174 1889 1230 1945
rect 1279 1889 1335 1945
rect 1384 1889 1440 1945
rect 1489 1889 1545 1945
rect 4452 2114 4508 2170
rect 4532 2114 4588 2170
rect 4452 2032 4508 2088
rect 4532 2032 4588 2088
rect 4452 1950 4508 2006
rect 4532 1950 4588 2006
rect 4452 1868 4508 1924
rect 4532 1868 4588 1924
rect 4452 1786 4508 1842
rect 4532 1786 4588 1842
<< metal3 >>
rect 1938 39865 2598 39874
rect 1938 39809 1949 39865
rect 2005 39809 2033 39865
rect 2089 39809 2117 39865
rect 2173 39809 2201 39865
rect 2257 39809 2285 39865
rect 2341 39809 2369 39865
rect 2425 39809 2453 39865
rect 2509 39809 2537 39865
rect 2593 39809 2598 39865
rect 1938 39785 2598 39809
rect 1938 39729 1949 39785
rect 2005 39729 2033 39785
rect 2089 39729 2117 39785
rect 2173 39729 2201 39785
rect 2257 39729 2285 39785
rect 2341 39729 2369 39785
rect 2425 39729 2453 39785
rect 2509 39729 2537 39785
rect 2593 39729 2598 39785
rect 1938 39705 2598 39729
rect 1938 39649 1949 39705
rect 2005 39649 2033 39705
rect 2089 39649 2117 39705
rect 2173 39649 2201 39705
rect 2257 39649 2285 39705
rect 2341 39649 2369 39705
rect 2425 39649 2453 39705
rect 2509 39649 2537 39705
rect 2593 39649 2598 39705
rect 1938 39625 2598 39649
rect 1938 39569 1949 39625
rect 2005 39569 2033 39625
rect 2089 39569 2117 39625
rect 2173 39569 2201 39625
rect 2257 39569 2285 39625
rect 2341 39569 2369 39625
rect 2425 39569 2453 39625
rect 2509 39569 2537 39625
rect 2593 39569 2598 39625
rect 1938 39545 2598 39569
rect 1938 39489 1949 39545
rect 2005 39489 2033 39545
rect 2089 39489 2117 39545
rect 2173 39489 2201 39545
rect 2257 39489 2285 39545
rect 2341 39489 2369 39545
rect 2425 39489 2453 39545
rect 2509 39489 2537 39545
rect 2593 39489 2598 39545
rect 1938 39465 2598 39489
rect 1938 39409 1949 39465
rect 2005 39409 2033 39465
rect 2089 39409 2117 39465
rect 2173 39409 2201 39465
rect 2257 39409 2285 39465
rect 2341 39409 2369 39465
rect 2425 39409 2453 39465
rect 2509 39409 2537 39465
rect 2593 39409 2598 39465
rect 1938 39385 2598 39409
rect 1938 39329 1949 39385
rect 2005 39329 2033 39385
rect 2089 39329 2117 39385
rect 2173 39329 2201 39385
rect 2257 39329 2285 39385
rect 2341 39329 2369 39385
rect 2425 39329 2453 39385
rect 2509 39329 2537 39385
rect 2593 39329 2598 39385
rect 1938 39305 2598 39329
rect 1938 39249 1949 39305
rect 2005 39249 2033 39305
rect 2089 39249 2117 39305
rect 2173 39249 2201 39305
rect 2257 39249 2285 39305
rect 2341 39249 2369 39305
rect 2425 39249 2453 39305
rect 2509 39249 2537 39305
rect 2593 39249 2598 39305
rect 1938 39225 2598 39249
rect 1938 39169 1949 39225
rect 2005 39169 2033 39225
rect 2089 39169 2117 39225
rect 2173 39169 2201 39225
rect 2257 39169 2285 39225
rect 2341 39169 2369 39225
rect 2425 39169 2453 39225
rect 2509 39169 2537 39225
rect 2593 39169 2598 39225
rect 1938 39145 2598 39169
rect 1938 39089 1949 39145
rect 2005 39089 2033 39145
rect 2089 39089 2117 39145
rect 2173 39089 2201 39145
rect 2257 39089 2285 39145
rect 2341 39089 2369 39145
rect 2425 39089 2453 39145
rect 2509 39089 2537 39145
rect 2593 39089 2598 39145
rect 1938 39065 2598 39089
rect 1938 39009 1949 39065
rect 2005 39009 2033 39065
rect 2089 39009 2117 39065
rect 2173 39009 2201 39065
rect 2257 39009 2285 39065
rect 2341 39009 2369 39065
rect 2425 39009 2453 39065
rect 2509 39009 2537 39065
rect 2593 39009 2598 39065
rect 1938 38985 2598 39009
rect 1938 38929 1949 38985
rect 2005 38929 2033 38985
rect 2089 38929 2117 38985
rect 2173 38929 2201 38985
rect 2257 38929 2285 38985
rect 2341 38929 2369 38985
rect 2425 38929 2453 38985
rect 2509 38929 2537 38985
rect 2593 38929 2598 38985
rect 1938 38905 2598 38929
rect 1938 38849 1949 38905
rect 2005 38849 2033 38905
rect 2089 38849 2117 38905
rect 2173 38849 2201 38905
rect 2257 38849 2285 38905
rect 2341 38849 2369 38905
rect 2425 38849 2453 38905
rect 2509 38849 2537 38905
rect 2593 38849 2598 38905
rect 1938 38825 2598 38849
rect 1938 38769 1949 38825
rect 2005 38769 2033 38825
rect 2089 38769 2117 38825
rect 2173 38769 2201 38825
rect 2257 38769 2285 38825
rect 2341 38769 2369 38825
rect 2425 38769 2453 38825
rect 2509 38769 2537 38825
rect 2593 38769 2598 38825
rect 1938 38745 2598 38769
rect 1938 38689 1949 38745
rect 2005 38689 2033 38745
rect 2089 38689 2117 38745
rect 2173 38689 2201 38745
rect 2257 38689 2285 38745
rect 2341 38689 2369 38745
rect 2425 38689 2453 38745
rect 2509 38689 2537 38745
rect 2593 38689 2598 38745
rect 1938 38665 2598 38689
rect 1938 38609 1949 38665
rect 2005 38609 2033 38665
rect 2089 38609 2117 38665
rect 2173 38609 2201 38665
rect 2257 38609 2285 38665
rect 2341 38609 2369 38665
rect 2425 38609 2453 38665
rect 2509 38609 2537 38665
rect 2593 38609 2598 38665
rect 1938 38585 2598 38609
rect 1938 38529 1949 38585
rect 2005 38529 2033 38585
rect 2089 38529 2117 38585
rect 2173 38529 2201 38585
rect 2257 38529 2285 38585
rect 2341 38529 2369 38585
rect 2425 38529 2453 38585
rect 2509 38529 2537 38585
rect 2593 38529 2598 38585
rect 1938 38505 2598 38529
rect 1938 38449 1949 38505
rect 2005 38449 2033 38505
rect 2089 38449 2117 38505
rect 2173 38449 2201 38505
rect 2257 38449 2285 38505
rect 2341 38449 2369 38505
rect 2425 38449 2453 38505
rect 2509 38449 2537 38505
rect 2593 38449 2598 38505
rect 1938 38425 2598 38449
rect 1938 38369 1949 38425
rect 2005 38369 2033 38425
rect 2089 38369 2117 38425
rect 2173 38369 2201 38425
rect 2257 38369 2285 38425
rect 2341 38369 2369 38425
rect 2425 38369 2453 38425
rect 2509 38369 2537 38425
rect 2593 38369 2598 38425
rect 1938 38345 2598 38369
rect 1938 38289 1949 38345
rect 2005 38289 2033 38345
rect 2089 38289 2117 38345
rect 2173 38289 2201 38345
rect 2257 38289 2285 38345
rect 2341 38289 2369 38345
rect 2425 38289 2453 38345
rect 2509 38289 2537 38345
rect 2593 38289 2598 38345
rect 1938 38265 2598 38289
rect 1938 38209 1949 38265
rect 2005 38209 2033 38265
rect 2089 38209 2117 38265
rect 2173 38209 2201 38265
rect 2257 38209 2285 38265
rect 2341 38209 2369 38265
rect 2425 38209 2453 38265
rect 2509 38209 2537 38265
rect 2593 38209 2598 38265
rect 1938 38185 2598 38209
rect 1938 38129 1949 38185
rect 2005 38129 2033 38185
rect 2089 38129 2117 38185
rect 2173 38129 2201 38185
rect 2257 38129 2285 38185
rect 2341 38129 2369 38185
rect 2425 38129 2453 38185
rect 2509 38129 2537 38185
rect 2593 38129 2598 38185
rect 1938 38105 2598 38129
rect 1938 38049 1949 38105
rect 2005 38049 2033 38105
rect 2089 38049 2117 38105
rect 2173 38049 2201 38105
rect 2257 38049 2285 38105
rect 2341 38049 2369 38105
rect 2425 38049 2453 38105
rect 2509 38049 2537 38105
rect 2593 38049 2598 38105
rect 1938 38025 2598 38049
rect 1938 37969 1949 38025
rect 2005 37969 2033 38025
rect 2089 37969 2117 38025
rect 2173 37969 2201 38025
rect 2257 37969 2285 38025
rect 2341 37969 2369 38025
rect 2425 37969 2453 38025
rect 2509 37969 2537 38025
rect 2593 37969 2598 38025
rect 1938 37945 2598 37969
rect 1938 37889 1949 37945
rect 2005 37889 2033 37945
rect 2089 37889 2117 37945
rect 2173 37889 2201 37945
rect 2257 37889 2285 37945
rect 2341 37889 2369 37945
rect 2425 37889 2453 37945
rect 2509 37889 2537 37945
rect 2593 37889 2598 37945
rect 1938 37865 2598 37889
rect 1938 37809 1949 37865
rect 2005 37809 2033 37865
rect 2089 37809 2117 37865
rect 2173 37809 2201 37865
rect 2257 37809 2285 37865
rect 2341 37809 2369 37865
rect 2425 37809 2453 37865
rect 2509 37809 2537 37865
rect 2593 37809 2598 37865
rect 1938 37785 2598 37809
rect 1938 37729 1949 37785
rect 2005 37729 2033 37785
rect 2089 37729 2117 37785
rect 2173 37729 2201 37785
rect 2257 37729 2285 37785
rect 2341 37729 2369 37785
rect 2425 37729 2453 37785
rect 2509 37729 2537 37785
rect 2593 37729 2598 37785
rect 1938 37705 2598 37729
rect 1938 37649 1949 37705
rect 2005 37649 2033 37705
rect 2089 37649 2117 37705
rect 2173 37649 2201 37705
rect 2257 37649 2285 37705
rect 2341 37649 2369 37705
rect 2425 37649 2453 37705
rect 2509 37649 2537 37705
rect 2593 37649 2598 37705
rect 1938 37625 2598 37649
rect 1938 37569 1949 37625
rect 2005 37569 2033 37625
rect 2089 37569 2117 37625
rect 2173 37569 2201 37625
rect 2257 37569 2285 37625
rect 2341 37569 2369 37625
rect 2425 37569 2453 37625
rect 2509 37569 2537 37625
rect 2593 37569 2598 37625
rect 1938 37545 2598 37569
rect 1938 37489 1949 37545
rect 2005 37489 2033 37545
rect 2089 37489 2117 37545
rect 2173 37489 2201 37545
rect 2257 37489 2285 37545
rect 2341 37489 2369 37545
rect 2425 37489 2453 37545
rect 2509 37489 2537 37545
rect 2593 37489 2598 37545
rect 1938 37465 2598 37489
rect 1938 37409 1949 37465
rect 2005 37409 2033 37465
rect 2089 37409 2117 37465
rect 2173 37409 2201 37465
rect 2257 37409 2285 37465
rect 2341 37409 2369 37465
rect 2425 37409 2453 37465
rect 2509 37409 2537 37465
rect 2593 37409 2598 37465
rect 1938 37385 2598 37409
rect 1938 37329 1949 37385
rect 2005 37329 2033 37385
rect 2089 37329 2117 37385
rect 2173 37329 2201 37385
rect 2257 37329 2285 37385
rect 2341 37329 2369 37385
rect 2425 37329 2453 37385
rect 2509 37329 2537 37385
rect 2593 37329 2598 37385
rect 1938 37305 2598 37329
rect 1938 37249 1949 37305
rect 2005 37249 2033 37305
rect 2089 37249 2117 37305
rect 2173 37249 2201 37305
rect 2257 37249 2285 37305
rect 2341 37249 2369 37305
rect 2425 37249 2453 37305
rect 2509 37249 2537 37305
rect 2593 37249 2598 37305
rect 1938 37225 2598 37249
rect 1938 37169 1949 37225
rect 2005 37169 2033 37225
rect 2089 37169 2117 37225
rect 2173 37169 2201 37225
rect 2257 37169 2285 37225
rect 2341 37169 2369 37225
rect 2425 37169 2453 37225
rect 2509 37169 2537 37225
rect 2593 37169 2598 37225
rect 1938 37145 2598 37169
rect 1938 37089 1949 37145
rect 2005 37089 2033 37145
rect 2089 37089 2117 37145
rect 2173 37089 2201 37145
rect 2257 37089 2285 37145
rect 2341 37089 2369 37145
rect 2425 37089 2453 37145
rect 2509 37089 2537 37145
rect 2593 37089 2598 37145
rect 1938 37065 2598 37089
rect 1938 37009 1949 37065
rect 2005 37009 2033 37065
rect 2089 37009 2117 37065
rect 2173 37009 2201 37065
rect 2257 37009 2285 37065
rect 2341 37009 2369 37065
rect 2425 37009 2453 37065
rect 2509 37009 2537 37065
rect 2593 37009 2598 37065
rect 1938 36985 2598 37009
rect 1938 36929 1949 36985
rect 2005 36929 2033 36985
rect 2089 36929 2117 36985
rect 2173 36929 2201 36985
rect 2257 36929 2285 36985
rect 2341 36929 2369 36985
rect 2425 36929 2453 36985
rect 2509 36929 2537 36985
rect 2593 36929 2598 36985
rect 1938 36905 2598 36929
rect 1938 36849 1949 36905
rect 2005 36849 2033 36905
rect 2089 36849 2117 36905
rect 2173 36849 2201 36905
rect 2257 36849 2285 36905
rect 2341 36849 2369 36905
rect 2425 36849 2453 36905
rect 2509 36849 2537 36905
rect 2593 36849 2598 36905
rect 1938 36825 2598 36849
rect 1938 36769 1949 36825
rect 2005 36769 2033 36825
rect 2089 36769 2117 36825
rect 2173 36769 2201 36825
rect 2257 36769 2285 36825
rect 2341 36769 2369 36825
rect 2425 36769 2453 36825
rect 2509 36769 2537 36825
rect 2593 36769 2598 36825
rect 1938 36745 2598 36769
rect 1938 36689 1949 36745
rect 2005 36689 2033 36745
rect 2089 36689 2117 36745
rect 2173 36689 2201 36745
rect 2257 36689 2285 36745
rect 2341 36689 2369 36745
rect 2425 36689 2453 36745
rect 2509 36689 2537 36745
rect 2593 36689 2598 36745
rect 1938 36665 2598 36689
rect 1938 36609 1949 36665
rect 2005 36609 2033 36665
rect 2089 36609 2117 36665
rect 2173 36609 2201 36665
rect 2257 36609 2285 36665
rect 2341 36609 2369 36665
rect 2425 36609 2453 36665
rect 2509 36609 2537 36665
rect 2593 36609 2598 36665
rect 1938 36585 2598 36609
rect 1938 36529 1949 36585
rect 2005 36529 2033 36585
rect 2089 36529 2117 36585
rect 2173 36529 2201 36585
rect 2257 36529 2285 36585
rect 2341 36529 2369 36585
rect 2425 36529 2453 36585
rect 2509 36529 2537 36585
rect 2593 36529 2598 36585
rect 1938 36505 2598 36529
rect 1938 36449 1949 36505
rect 2005 36449 2033 36505
rect 2089 36449 2117 36505
rect 2173 36449 2201 36505
rect 2257 36449 2285 36505
rect 2341 36449 2369 36505
rect 2425 36449 2453 36505
rect 2509 36449 2537 36505
rect 2593 36449 2598 36505
rect 1938 36425 2598 36449
rect 1938 36369 1949 36425
rect 2005 36369 2033 36425
rect 2089 36369 2117 36425
rect 2173 36369 2201 36425
rect 2257 36369 2285 36425
rect 2341 36369 2369 36425
rect 2425 36369 2453 36425
rect 2509 36369 2537 36425
rect 2593 36369 2598 36425
rect 1938 36345 2598 36369
rect 1938 36289 1949 36345
rect 2005 36289 2033 36345
rect 2089 36289 2117 36345
rect 2173 36289 2201 36345
rect 2257 36289 2285 36345
rect 2341 36289 2369 36345
rect 2425 36289 2453 36345
rect 2509 36289 2537 36345
rect 2593 36289 2598 36345
rect 1938 36265 2598 36289
rect 1938 36209 1949 36265
rect 2005 36209 2033 36265
rect 2089 36209 2117 36265
rect 2173 36209 2201 36265
rect 2257 36209 2285 36265
rect 2341 36209 2369 36265
rect 2425 36209 2453 36265
rect 2509 36209 2537 36265
rect 2593 36209 2598 36265
rect 1938 36185 2598 36209
rect 1938 36129 1949 36185
rect 2005 36129 2033 36185
rect 2089 36129 2117 36185
rect 2173 36129 2201 36185
rect 2257 36129 2285 36185
rect 2341 36129 2369 36185
rect 2425 36129 2453 36185
rect 2509 36129 2537 36185
rect 2593 36129 2598 36185
rect 1938 36105 2598 36129
rect 1938 36049 1949 36105
rect 2005 36049 2033 36105
rect 2089 36049 2117 36105
rect 2173 36049 2201 36105
rect 2257 36049 2285 36105
rect 2341 36049 2369 36105
rect 2425 36049 2453 36105
rect 2509 36049 2537 36105
rect 2593 36049 2598 36105
rect 1938 36025 2598 36049
rect 1938 35969 1949 36025
rect 2005 35969 2033 36025
rect 2089 35969 2117 36025
rect 2173 35969 2201 36025
rect 2257 35969 2285 36025
rect 2341 35969 2369 36025
rect 2425 35969 2453 36025
rect 2509 35969 2537 36025
rect 2593 35969 2598 36025
rect 1938 35945 2598 35969
rect 1938 35889 1949 35945
rect 2005 35889 2033 35945
rect 2089 35889 2117 35945
rect 2173 35889 2201 35945
rect 2257 35889 2285 35945
rect 2341 35889 2369 35945
rect 2425 35889 2453 35945
rect 2509 35889 2537 35945
rect 2593 35889 2598 35945
rect 1938 35865 2598 35889
rect 1938 35809 1949 35865
rect 2005 35809 2033 35865
rect 2089 35809 2117 35865
rect 2173 35809 2201 35865
rect 2257 35809 2285 35865
rect 2341 35809 2369 35865
rect 2425 35809 2453 35865
rect 2509 35809 2537 35865
rect 2593 35809 2598 35865
rect 1938 35785 2598 35809
rect 1938 35729 1949 35785
rect 2005 35729 2033 35785
rect 2089 35729 2117 35785
rect 2173 35729 2201 35785
rect 2257 35729 2285 35785
rect 2341 35729 2369 35785
rect 2425 35729 2453 35785
rect 2509 35729 2537 35785
rect 2593 35729 2598 35785
rect 1938 35705 2598 35729
rect 1938 35649 1949 35705
rect 2005 35649 2033 35705
rect 2089 35649 2117 35705
rect 2173 35649 2201 35705
rect 2257 35649 2285 35705
rect 2341 35649 2369 35705
rect 2425 35649 2453 35705
rect 2509 35649 2537 35705
rect 2593 35649 2598 35705
rect 1938 35625 2598 35649
rect 1938 35569 1949 35625
rect 2005 35569 2033 35625
rect 2089 35569 2117 35625
rect 2173 35569 2201 35625
rect 2257 35569 2285 35625
rect 2341 35569 2369 35625
rect 2425 35569 2453 35625
rect 2509 35569 2537 35625
rect 2593 35569 2598 35625
rect 1938 35545 2598 35569
rect 1938 35489 1949 35545
rect 2005 35489 2033 35545
rect 2089 35489 2117 35545
rect 2173 35489 2201 35545
rect 2257 35489 2285 35545
rect 2341 35489 2369 35545
rect 2425 35489 2453 35545
rect 2509 35489 2537 35545
rect 2593 35489 2598 35545
rect 1938 35465 2598 35489
rect 1938 35409 1949 35465
rect 2005 35409 2033 35465
rect 2089 35409 2117 35465
rect 2173 35409 2201 35465
rect 2257 35409 2285 35465
rect 2341 35409 2369 35465
rect 2425 35409 2453 35465
rect 2509 35409 2537 35465
rect 2593 35409 2598 35465
rect 1938 35385 2598 35409
rect 1938 35329 1949 35385
rect 2005 35329 2033 35385
rect 2089 35329 2117 35385
rect 2173 35329 2201 35385
rect 2257 35329 2285 35385
rect 2341 35329 2369 35385
rect 2425 35329 2453 35385
rect 2509 35329 2537 35385
rect 2593 35329 2598 35385
rect 1938 35305 2598 35329
rect 1938 35249 1949 35305
rect 2005 35249 2033 35305
rect 2089 35249 2117 35305
rect 2173 35249 2201 35305
rect 2257 35249 2285 35305
rect 2341 35249 2369 35305
rect 2425 35249 2453 35305
rect 2509 35249 2537 35305
rect 2593 35249 2598 35305
rect 1938 35225 2598 35249
rect 1938 35169 1949 35225
rect 2005 35169 2033 35225
rect 2089 35169 2117 35225
rect 2173 35169 2201 35225
rect 2257 35169 2285 35225
rect 2341 35169 2369 35225
rect 2425 35169 2453 35225
rect 2509 35169 2537 35225
rect 2593 35169 2598 35225
rect 1938 35145 2598 35169
rect 1938 35089 1949 35145
rect 2005 35089 2033 35145
rect 2089 35089 2117 35145
rect 2173 35089 2201 35145
rect 2257 35089 2285 35145
rect 2341 35089 2369 35145
rect 2425 35089 2453 35145
rect 2509 35089 2537 35145
rect 2593 35089 2598 35145
rect 6890 39870 7528 39882
rect 6890 39814 6903 39870
rect 6959 39814 6993 39870
rect 7049 39814 7083 39870
rect 7139 39814 7173 39870
rect 7229 39814 7263 39870
rect 7319 39814 7353 39870
rect 7409 39814 7443 39870
rect 7499 39814 7528 39870
rect 6890 39790 7528 39814
rect 6890 39734 6903 39790
rect 6959 39734 6993 39790
rect 7049 39734 7083 39790
rect 7139 39734 7173 39790
rect 7229 39734 7263 39790
rect 7319 39734 7353 39790
rect 7409 39734 7443 39790
rect 7499 39734 7528 39790
rect 6890 39710 7528 39734
rect 6890 39654 6903 39710
rect 6959 39654 6993 39710
rect 7049 39654 7083 39710
rect 7139 39654 7173 39710
rect 7229 39654 7263 39710
rect 7319 39654 7353 39710
rect 7409 39654 7443 39710
rect 7499 39654 7528 39710
rect 6890 39630 7528 39654
rect 6890 39574 6903 39630
rect 6959 39574 6993 39630
rect 7049 39574 7083 39630
rect 7139 39574 7173 39630
rect 7229 39574 7263 39630
rect 7319 39574 7353 39630
rect 7409 39574 7443 39630
rect 7499 39574 7528 39630
rect 6890 39550 7528 39574
rect 6890 39494 6903 39550
rect 6959 39494 6993 39550
rect 7049 39494 7083 39550
rect 7139 39494 7173 39550
rect 7229 39494 7263 39550
rect 7319 39494 7353 39550
rect 7409 39494 7443 39550
rect 7499 39494 7528 39550
rect 6890 39470 7528 39494
rect 6890 39414 6903 39470
rect 6959 39414 6993 39470
rect 7049 39414 7083 39470
rect 7139 39414 7173 39470
rect 7229 39414 7263 39470
rect 7319 39414 7353 39470
rect 7409 39414 7443 39470
rect 7499 39414 7528 39470
rect 6890 39390 7528 39414
rect 6890 39334 6903 39390
rect 6959 39334 6993 39390
rect 7049 39334 7083 39390
rect 7139 39334 7173 39390
rect 7229 39334 7263 39390
rect 7319 39334 7353 39390
rect 7409 39334 7443 39390
rect 7499 39334 7528 39390
rect 6890 39310 7528 39334
rect 6890 39254 6903 39310
rect 6959 39254 6993 39310
rect 7049 39254 7083 39310
rect 7139 39254 7173 39310
rect 7229 39254 7263 39310
rect 7319 39254 7353 39310
rect 7409 39254 7443 39310
rect 7499 39254 7528 39310
rect 6890 39230 7528 39254
rect 6890 39174 6903 39230
rect 6959 39174 6993 39230
rect 7049 39174 7083 39230
rect 7139 39174 7173 39230
rect 7229 39174 7263 39230
rect 7319 39174 7353 39230
rect 7409 39174 7443 39230
rect 7499 39174 7528 39230
rect 6890 39150 7528 39174
rect 6890 39094 6903 39150
rect 6959 39094 6993 39150
rect 7049 39094 7083 39150
rect 7139 39094 7173 39150
rect 7229 39094 7263 39150
rect 7319 39094 7353 39150
rect 7409 39094 7443 39150
rect 7499 39094 7528 39150
rect 6890 39070 7528 39094
rect 6890 39014 6903 39070
rect 6959 39014 6993 39070
rect 7049 39014 7083 39070
rect 7139 39014 7173 39070
rect 7229 39014 7263 39070
rect 7319 39014 7353 39070
rect 7409 39014 7443 39070
rect 7499 39014 7528 39070
rect 6890 38990 7528 39014
rect 6890 38934 6903 38990
rect 6959 38934 6993 38990
rect 7049 38934 7083 38990
rect 7139 38934 7173 38990
rect 7229 38934 7263 38990
rect 7319 38934 7353 38990
rect 7409 38934 7443 38990
rect 7499 38934 7528 38990
rect 6890 38910 7528 38934
rect 6890 38854 6903 38910
rect 6959 38854 6993 38910
rect 7049 38854 7083 38910
rect 7139 38854 7173 38910
rect 7229 38854 7263 38910
rect 7319 38854 7353 38910
rect 7409 38854 7443 38910
rect 7499 38854 7528 38910
rect 6890 38830 7528 38854
rect 6890 38774 6903 38830
rect 6959 38774 6993 38830
rect 7049 38774 7083 38830
rect 7139 38774 7173 38830
rect 7229 38774 7263 38830
rect 7319 38774 7353 38830
rect 7409 38774 7443 38830
rect 7499 38774 7528 38830
rect 6890 38750 7528 38774
rect 6890 38694 6903 38750
rect 6959 38694 6993 38750
rect 7049 38694 7083 38750
rect 7139 38694 7173 38750
rect 7229 38694 7263 38750
rect 7319 38694 7353 38750
rect 7409 38694 7443 38750
rect 7499 38694 7528 38750
rect 6890 38670 7528 38694
rect 6890 38614 6903 38670
rect 6959 38614 6993 38670
rect 7049 38614 7083 38670
rect 7139 38614 7173 38670
rect 7229 38614 7263 38670
rect 7319 38614 7353 38670
rect 7409 38614 7443 38670
rect 7499 38614 7528 38670
rect 6890 38590 7528 38614
rect 6890 38534 6903 38590
rect 6959 38534 6993 38590
rect 7049 38534 7083 38590
rect 7139 38534 7173 38590
rect 7229 38534 7263 38590
rect 7319 38534 7353 38590
rect 7409 38534 7443 38590
rect 7499 38534 7528 38590
rect 6890 38510 7528 38534
rect 6890 38454 6903 38510
rect 6959 38454 6993 38510
rect 7049 38454 7083 38510
rect 7139 38454 7173 38510
rect 7229 38454 7263 38510
rect 7319 38454 7353 38510
rect 7409 38454 7443 38510
rect 7499 38454 7528 38510
rect 6890 38430 7528 38454
rect 6890 38374 6903 38430
rect 6959 38374 6993 38430
rect 7049 38374 7083 38430
rect 7139 38374 7173 38430
rect 7229 38374 7263 38430
rect 7319 38374 7353 38430
rect 7409 38374 7443 38430
rect 7499 38374 7528 38430
rect 6890 38350 7528 38374
rect 6890 38294 6903 38350
rect 6959 38294 6993 38350
rect 7049 38294 7083 38350
rect 7139 38294 7173 38350
rect 7229 38294 7263 38350
rect 7319 38294 7353 38350
rect 7409 38294 7443 38350
rect 7499 38294 7528 38350
rect 6890 38270 7528 38294
rect 6890 38214 6903 38270
rect 6959 38214 6993 38270
rect 7049 38214 7083 38270
rect 7139 38214 7173 38270
rect 7229 38214 7263 38270
rect 7319 38214 7353 38270
rect 7409 38214 7443 38270
rect 7499 38214 7528 38270
rect 6890 38190 7528 38214
rect 6890 38134 6903 38190
rect 6959 38134 6993 38190
rect 7049 38134 7083 38190
rect 7139 38134 7173 38190
rect 7229 38134 7263 38190
rect 7319 38134 7353 38190
rect 7409 38134 7443 38190
rect 7499 38134 7528 38190
rect 6890 38110 7528 38134
rect 6890 38054 6903 38110
rect 6959 38054 6993 38110
rect 7049 38054 7083 38110
rect 7139 38054 7173 38110
rect 7229 38054 7263 38110
rect 7319 38054 7353 38110
rect 7409 38054 7443 38110
rect 7499 38054 7528 38110
rect 6890 38030 7528 38054
rect 6890 37974 6903 38030
rect 6959 37974 6993 38030
rect 7049 37974 7083 38030
rect 7139 37974 7173 38030
rect 7229 37974 7263 38030
rect 7319 37974 7353 38030
rect 7409 37974 7443 38030
rect 7499 37974 7528 38030
rect 6890 37950 7528 37974
rect 6890 37894 6903 37950
rect 6959 37894 6993 37950
rect 7049 37894 7083 37950
rect 7139 37894 7173 37950
rect 7229 37894 7263 37950
rect 7319 37894 7353 37950
rect 7409 37894 7443 37950
rect 7499 37894 7528 37950
rect 6890 37870 7528 37894
rect 6890 37814 6903 37870
rect 6959 37814 6993 37870
rect 7049 37814 7083 37870
rect 7139 37814 7173 37870
rect 7229 37814 7263 37870
rect 7319 37814 7353 37870
rect 7409 37814 7443 37870
rect 7499 37814 7528 37870
rect 6890 37790 7528 37814
rect 6890 37734 6903 37790
rect 6959 37734 6993 37790
rect 7049 37734 7083 37790
rect 7139 37734 7173 37790
rect 7229 37734 7263 37790
rect 7319 37734 7353 37790
rect 7409 37734 7443 37790
rect 7499 37734 7528 37790
rect 6890 37710 7528 37734
rect 6890 37654 6903 37710
rect 6959 37654 6993 37710
rect 7049 37654 7083 37710
rect 7139 37654 7173 37710
rect 7229 37654 7263 37710
rect 7319 37654 7353 37710
rect 7409 37654 7443 37710
rect 7499 37654 7528 37710
rect 6890 37630 7528 37654
rect 6890 37574 6903 37630
rect 6959 37574 6993 37630
rect 7049 37574 7083 37630
rect 7139 37574 7173 37630
rect 7229 37574 7263 37630
rect 7319 37574 7353 37630
rect 7409 37574 7443 37630
rect 7499 37574 7528 37630
rect 6890 37550 7528 37574
rect 6890 37494 6903 37550
rect 6959 37494 6993 37550
rect 7049 37494 7083 37550
rect 7139 37494 7173 37550
rect 7229 37494 7263 37550
rect 7319 37494 7353 37550
rect 7409 37494 7443 37550
rect 7499 37494 7528 37550
rect 6890 37470 7528 37494
rect 6890 37414 6903 37470
rect 6959 37414 6993 37470
rect 7049 37414 7083 37470
rect 7139 37414 7173 37470
rect 7229 37414 7263 37470
rect 7319 37414 7353 37470
rect 7409 37414 7443 37470
rect 7499 37414 7528 37470
rect 6890 37390 7528 37414
rect 6890 37334 6903 37390
rect 6959 37334 6993 37390
rect 7049 37334 7083 37390
rect 7139 37334 7173 37390
rect 7229 37334 7263 37390
rect 7319 37334 7353 37390
rect 7409 37334 7443 37390
rect 7499 37334 7528 37390
rect 6890 37310 7528 37334
rect 6890 37254 6903 37310
rect 6959 37254 6993 37310
rect 7049 37254 7083 37310
rect 7139 37254 7173 37310
rect 7229 37254 7263 37310
rect 7319 37254 7353 37310
rect 7409 37254 7443 37310
rect 7499 37254 7528 37310
rect 6890 37230 7528 37254
rect 6890 37174 6903 37230
rect 6959 37174 6993 37230
rect 7049 37174 7083 37230
rect 7139 37174 7173 37230
rect 7229 37174 7263 37230
rect 7319 37174 7353 37230
rect 7409 37174 7443 37230
rect 7499 37174 7528 37230
rect 6890 37150 7528 37174
rect 6890 37094 6903 37150
rect 6959 37094 6993 37150
rect 7049 37094 7083 37150
rect 7139 37094 7173 37150
rect 7229 37094 7263 37150
rect 7319 37094 7353 37150
rect 7409 37094 7443 37150
rect 7499 37094 7528 37150
rect 6890 37070 7528 37094
rect 6890 37014 6903 37070
rect 6959 37014 6993 37070
rect 7049 37014 7083 37070
rect 7139 37014 7173 37070
rect 7229 37014 7263 37070
rect 7319 37014 7353 37070
rect 7409 37014 7443 37070
rect 7499 37014 7528 37070
rect 6890 36990 7528 37014
rect 6890 36934 6903 36990
rect 6959 36934 6993 36990
rect 7049 36934 7083 36990
rect 7139 36934 7173 36990
rect 7229 36934 7263 36990
rect 7319 36934 7353 36990
rect 7409 36934 7443 36990
rect 7499 36934 7528 36990
rect 6890 36910 7528 36934
rect 6890 36854 6903 36910
rect 6959 36854 6993 36910
rect 7049 36854 7083 36910
rect 7139 36854 7173 36910
rect 7229 36854 7263 36910
rect 7319 36854 7353 36910
rect 7409 36854 7443 36910
rect 7499 36854 7528 36910
rect 6890 36830 7528 36854
rect 6890 36774 6903 36830
rect 6959 36774 6993 36830
rect 7049 36774 7083 36830
rect 7139 36774 7173 36830
rect 7229 36774 7263 36830
rect 7319 36774 7353 36830
rect 7409 36774 7443 36830
rect 7499 36774 7528 36830
rect 6890 36750 7528 36774
rect 6890 36694 6903 36750
rect 6959 36694 6993 36750
rect 7049 36694 7083 36750
rect 7139 36694 7173 36750
rect 7229 36694 7263 36750
rect 7319 36694 7353 36750
rect 7409 36694 7443 36750
rect 7499 36694 7528 36750
rect 6890 36670 7528 36694
rect 6890 36614 6903 36670
rect 6959 36614 6993 36670
rect 7049 36614 7083 36670
rect 7139 36614 7173 36670
rect 7229 36614 7263 36670
rect 7319 36614 7353 36670
rect 7409 36614 7443 36670
rect 7499 36614 7528 36670
rect 6890 36590 7528 36614
rect 6890 36534 6903 36590
rect 6959 36534 6993 36590
rect 7049 36534 7083 36590
rect 7139 36534 7173 36590
rect 7229 36534 7263 36590
rect 7319 36534 7353 36590
rect 7409 36534 7443 36590
rect 7499 36534 7528 36590
rect 6890 36510 7528 36534
rect 6890 36454 6903 36510
rect 6959 36454 6993 36510
rect 7049 36454 7083 36510
rect 7139 36454 7173 36510
rect 7229 36454 7263 36510
rect 7319 36454 7353 36510
rect 7409 36454 7443 36510
rect 7499 36454 7528 36510
rect 6890 36430 7528 36454
rect 6890 36374 6903 36430
rect 6959 36374 6993 36430
rect 7049 36374 7083 36430
rect 7139 36374 7173 36430
rect 7229 36374 7263 36430
rect 7319 36374 7353 36430
rect 7409 36374 7443 36430
rect 7499 36374 7528 36430
rect 6890 36350 7528 36374
rect 6890 36294 6903 36350
rect 6959 36294 6993 36350
rect 7049 36294 7083 36350
rect 7139 36294 7173 36350
rect 7229 36294 7263 36350
rect 7319 36294 7353 36350
rect 7409 36294 7443 36350
rect 7499 36294 7528 36350
rect 6890 36270 7528 36294
rect 6890 36214 6903 36270
rect 6959 36214 6993 36270
rect 7049 36214 7083 36270
rect 7139 36214 7173 36270
rect 7229 36214 7263 36270
rect 7319 36214 7353 36270
rect 7409 36214 7443 36270
rect 7499 36214 7528 36270
rect 6890 36190 7528 36214
rect 6890 36134 6903 36190
rect 6959 36134 6993 36190
rect 7049 36134 7083 36190
rect 7139 36134 7173 36190
rect 7229 36134 7263 36190
rect 7319 36134 7353 36190
rect 7409 36134 7443 36190
rect 7499 36134 7528 36190
rect 6890 36110 7528 36134
rect 6890 36054 6903 36110
rect 6959 36054 6993 36110
rect 7049 36054 7083 36110
rect 7139 36054 7173 36110
rect 7229 36054 7263 36110
rect 7319 36054 7353 36110
rect 7409 36054 7443 36110
rect 7499 36054 7528 36110
rect 6890 36030 7528 36054
rect 6890 35974 6903 36030
rect 6959 35974 6993 36030
rect 7049 35974 7083 36030
rect 7139 35974 7173 36030
rect 7229 35974 7263 36030
rect 7319 35974 7353 36030
rect 7409 35974 7443 36030
rect 7499 35974 7528 36030
rect 6890 35950 7528 35974
rect 6890 35894 6903 35950
rect 6959 35894 6993 35950
rect 7049 35894 7083 35950
rect 7139 35894 7173 35950
rect 7229 35894 7263 35950
rect 7319 35894 7353 35950
rect 7409 35894 7443 35950
rect 7499 35894 7528 35950
rect 6890 35870 7528 35894
rect 6890 35814 6903 35870
rect 6959 35814 6993 35870
rect 7049 35814 7083 35870
rect 7139 35814 7173 35870
rect 7229 35814 7263 35870
rect 7319 35814 7353 35870
rect 7409 35814 7443 35870
rect 7499 35814 7528 35870
rect 6890 35790 7528 35814
rect 6890 35734 6903 35790
rect 6959 35734 6993 35790
rect 7049 35734 7083 35790
rect 7139 35734 7173 35790
rect 7229 35734 7263 35790
rect 7319 35734 7353 35790
rect 7409 35734 7443 35790
rect 7499 35734 7528 35790
rect 6890 35710 7528 35734
rect 6890 35654 6903 35710
rect 6959 35654 6993 35710
rect 7049 35654 7083 35710
rect 7139 35654 7173 35710
rect 7229 35654 7263 35710
rect 7319 35654 7353 35710
rect 7409 35654 7443 35710
rect 7499 35654 7528 35710
rect 6890 35630 7528 35654
rect 6890 35574 6903 35630
rect 6959 35574 6993 35630
rect 7049 35574 7083 35630
rect 7139 35574 7173 35630
rect 7229 35574 7263 35630
rect 7319 35574 7353 35630
rect 7409 35574 7443 35630
rect 7499 35574 7528 35630
rect 6890 35550 7528 35574
rect 6890 35494 6903 35550
rect 6959 35494 6993 35550
rect 7049 35494 7083 35550
rect 7139 35494 7173 35550
rect 7229 35494 7263 35550
rect 7319 35494 7353 35550
rect 7409 35494 7443 35550
rect 7499 35494 7528 35550
rect 6890 35470 7528 35494
rect 6890 35414 6903 35470
rect 6959 35414 6993 35470
rect 7049 35414 7083 35470
rect 7139 35414 7173 35470
rect 7229 35414 7263 35470
rect 7319 35414 7353 35470
rect 7409 35414 7443 35470
rect 7499 35414 7528 35470
rect 6890 35390 7528 35414
rect 6890 35334 6903 35390
rect 6959 35334 6993 35390
rect 7049 35334 7083 35390
rect 7139 35334 7173 35390
rect 7229 35334 7263 35390
rect 7319 35334 7353 35390
rect 7409 35334 7443 35390
rect 7499 35334 7528 35390
rect 6890 35310 7528 35334
rect 6890 35254 6903 35310
rect 6959 35254 6993 35310
rect 7049 35254 7083 35310
rect 7139 35254 7173 35310
rect 7229 35254 7263 35310
rect 7319 35254 7353 35310
rect 7409 35254 7443 35310
rect 7499 35254 7528 35310
rect 6890 35230 7528 35254
rect 6890 35174 6903 35230
rect 6959 35174 6993 35230
rect 7049 35174 7083 35230
rect 7139 35174 7173 35230
rect 7229 35174 7263 35230
rect 7319 35174 7353 35230
rect 7409 35174 7443 35230
rect 7499 35174 7528 35230
rect 6890 35150 7528 35174
rect 1938 35065 2598 35089
rect 1938 35009 1949 35065
rect 2005 35009 2033 35065
rect 2089 35009 2117 35065
rect 2173 35009 2201 35065
rect 2257 35009 2285 35065
rect 2341 35009 2369 35065
rect 2425 35009 2453 35065
rect 2509 35009 2537 35065
rect 2593 35009 2598 35065
rect 1938 34985 2598 35009
rect 1938 34929 1949 34985
rect 2005 34929 2033 34985
rect 2089 34929 2117 34985
rect 2173 34929 2201 34985
rect 2257 34929 2285 34985
rect 2341 34929 2369 34985
rect 2425 34929 2453 34985
rect 2509 34929 2537 34985
rect 2593 34929 2598 34985
rect 1938 34905 2598 34929
rect 1938 34849 1949 34905
rect 2005 34849 2033 34905
rect 2089 34849 2117 34905
rect 2173 34849 2201 34905
rect 2257 34849 2285 34905
rect 2341 34849 2369 34905
rect 2425 34849 2453 34905
rect 2509 34849 2537 34905
rect 2593 34849 2598 34905
rect 1938 34825 2598 34849
rect 1938 34769 1949 34825
rect 2005 34769 2033 34825
rect 2089 34769 2117 34825
rect 2173 34769 2201 34825
rect 2257 34769 2285 34825
rect 2341 34769 2369 34825
rect 2425 34769 2453 34825
rect 2509 34769 2537 34825
rect 2593 34769 2598 34825
rect 1938 34745 2598 34769
rect 1938 34689 1949 34745
rect 2005 34689 2033 34745
rect 2089 34689 2117 34745
rect 2173 34689 2201 34745
rect 2257 34689 2285 34745
rect 2341 34689 2369 34745
rect 2425 34689 2453 34745
rect 2509 34689 2537 34745
rect 2593 34689 2598 34745
rect 1938 34665 2598 34689
rect 1938 34609 1949 34665
rect 2005 34609 2033 34665
rect 2089 34609 2117 34665
rect 2173 34609 2201 34665
rect 2257 34609 2285 34665
rect 2341 34609 2369 34665
rect 2425 34609 2453 34665
rect 2509 34609 2537 34665
rect 2593 34609 2598 34665
rect 1938 34585 2598 34609
rect 1938 34529 1949 34585
rect 2005 34529 2033 34585
rect 2089 34529 2117 34585
rect 2173 34529 2201 34585
rect 2257 34529 2285 34585
rect 2341 34529 2369 34585
rect 2425 34529 2453 34585
rect 2509 34529 2537 34585
rect 2593 34529 2598 34585
rect 1938 34505 2598 34529
rect 1938 34449 1949 34505
rect 2005 34449 2033 34505
rect 2089 34449 2117 34505
rect 2173 34449 2201 34505
rect 2257 34449 2285 34505
rect 2341 34449 2369 34505
rect 2425 34449 2453 34505
rect 2509 34449 2537 34505
rect 2593 34449 2598 34505
rect 1938 34425 2598 34449
rect 1938 34369 1949 34425
rect 2005 34369 2033 34425
rect 2089 34369 2117 34425
rect 2173 34369 2201 34425
rect 2257 34369 2285 34425
rect 2341 34369 2369 34425
rect 2425 34369 2453 34425
rect 2509 34369 2537 34425
rect 2593 34369 2598 34425
rect 1938 34345 2598 34369
rect 1938 34289 1949 34345
rect 2005 34289 2033 34345
rect 2089 34289 2117 34345
rect 2173 34289 2201 34345
rect 2257 34289 2285 34345
rect 2341 34289 2369 34345
rect 2425 34289 2453 34345
rect 2509 34289 2537 34345
rect 2593 34289 2598 34345
rect 1938 34265 2598 34289
rect 1938 34209 1949 34265
rect 2005 34209 2033 34265
rect 2089 34209 2117 34265
rect 2173 34209 2201 34265
rect 2257 34209 2285 34265
rect 2341 34209 2369 34265
rect 2425 34209 2453 34265
rect 2509 34209 2537 34265
rect 2593 34209 2598 34265
rect 1938 34185 2598 34209
rect 1938 34129 1949 34185
rect 2005 34129 2033 34185
rect 2089 34129 2117 34185
rect 2173 34129 2201 34185
rect 2257 34129 2285 34185
rect 2341 34129 2369 34185
rect 2425 34129 2453 34185
rect 2509 34129 2537 34185
rect 2593 34129 2598 34185
rect 1938 34105 2598 34129
rect 1938 34049 1949 34105
rect 2005 34049 2033 34105
rect 2089 34049 2117 34105
rect 2173 34049 2201 34105
rect 2257 34049 2285 34105
rect 2341 34049 2369 34105
rect 2425 34049 2453 34105
rect 2509 34049 2537 34105
rect 2593 34049 2598 34105
rect 1938 34025 2598 34049
rect 1938 33969 1949 34025
rect 2005 33969 2033 34025
rect 2089 33969 2117 34025
rect 2173 33969 2201 34025
rect 2257 33969 2285 34025
rect 2341 33969 2369 34025
rect 2425 33969 2453 34025
rect 2509 33969 2537 34025
rect 2593 33969 2598 34025
rect 1938 33945 2598 33969
rect 1938 33889 1949 33945
rect 2005 33889 2033 33945
rect 2089 33889 2117 33945
rect 2173 33889 2201 33945
rect 2257 33889 2285 33945
rect 2341 33889 2369 33945
rect 2425 33889 2453 33945
rect 2509 33889 2537 33945
rect 2593 33889 2598 33945
rect 1938 33865 2598 33889
rect 1938 33809 1949 33865
rect 2005 33809 2033 33865
rect 2089 33809 2117 33865
rect 2173 33809 2201 33865
rect 2257 33809 2285 33865
rect 2341 33809 2369 33865
rect 2425 33809 2453 33865
rect 2509 33809 2537 33865
rect 2593 33809 2598 33865
rect 1938 33785 2598 33809
rect 1938 33729 1949 33785
rect 2005 33729 2033 33785
rect 2089 33729 2117 33785
rect 2173 33729 2201 33785
rect 2257 33729 2285 33785
rect 2341 33729 2369 33785
rect 2425 33729 2453 33785
rect 2509 33729 2537 33785
rect 2593 33729 2598 33785
rect 1938 33705 2598 33729
rect 1938 33649 1949 33705
rect 2005 33649 2033 33705
rect 2089 33649 2117 33705
rect 2173 33649 2201 33705
rect 2257 33649 2285 33705
rect 2341 33649 2369 33705
rect 2425 33649 2453 33705
rect 2509 33649 2537 33705
rect 2593 33649 2598 33705
rect 1938 33625 2598 33649
rect 1938 33569 1949 33625
rect 2005 33569 2033 33625
rect 2089 33569 2117 33625
rect 2173 33569 2201 33625
rect 2257 33569 2285 33625
rect 2341 33569 2369 33625
rect 2425 33569 2453 33625
rect 2509 33569 2537 33625
rect 2593 33569 2598 33625
rect 1938 33545 2598 33569
rect 1938 33489 1949 33545
rect 2005 33489 2033 33545
rect 2089 33489 2117 33545
rect 2173 33489 2201 33545
rect 2257 33489 2285 33545
rect 2341 33489 2369 33545
rect 2425 33489 2453 33545
rect 2509 33489 2537 33545
rect 2593 33489 2598 33545
rect 1938 33465 2598 33489
rect 1938 33409 1949 33465
rect 2005 33409 2033 33465
rect 2089 33409 2117 33465
rect 2173 33409 2201 33465
rect 2257 33409 2285 33465
rect 2341 33409 2369 33465
rect 2425 33409 2453 33465
rect 2509 33409 2537 33465
rect 2593 33409 2598 33465
rect 1938 33385 2598 33409
rect 1938 33329 1949 33385
rect 2005 33329 2033 33385
rect 2089 33329 2117 33385
rect 2173 33329 2201 33385
rect 2257 33329 2285 33385
rect 2341 33329 2369 33385
rect 2425 33329 2453 33385
rect 2509 33329 2537 33385
rect 2593 33329 2598 33385
rect 1938 33305 2598 33329
rect 1938 33249 1949 33305
rect 2005 33249 2033 33305
rect 2089 33249 2117 33305
rect 2173 33249 2201 33305
rect 2257 33249 2285 33305
rect 2341 33249 2369 33305
rect 2425 33249 2453 33305
rect 2509 33249 2537 33305
rect 2593 33249 2598 33305
rect 1938 33225 2598 33249
rect 1938 33169 1949 33225
rect 2005 33169 2033 33225
rect 2089 33169 2117 33225
rect 2173 33169 2201 33225
rect 2257 33169 2285 33225
rect 2341 33169 2369 33225
rect 2425 33169 2453 33225
rect 2509 33169 2537 33225
rect 2593 33169 2598 33225
rect 1938 33145 2598 33169
rect 1938 33089 1949 33145
rect 2005 33089 2033 33145
rect 2089 33089 2117 33145
rect 2173 33089 2201 33145
rect 2257 33089 2285 33145
rect 2341 33089 2369 33145
rect 2425 33089 2453 33145
rect 2509 33089 2537 33145
rect 2593 33089 2598 33145
rect 1938 33065 2598 33089
rect 1938 33009 1949 33065
rect 2005 33009 2033 33065
rect 2089 33009 2117 33065
rect 2173 33009 2201 33065
rect 2257 33009 2285 33065
rect 2341 33009 2369 33065
rect 2425 33009 2453 33065
rect 2509 33009 2537 33065
rect 2593 33009 2598 33065
rect 1938 32985 2598 33009
rect 1938 32929 1949 32985
rect 2005 32929 2033 32985
rect 2089 32929 2117 32985
rect 2173 32929 2201 32985
rect 2257 32929 2285 32985
rect 2341 32929 2369 32985
rect 2425 32929 2453 32985
rect 2509 32929 2537 32985
rect 2593 32929 2598 32985
rect 1938 32905 2598 32929
rect 1938 32849 1949 32905
rect 2005 32849 2033 32905
rect 2089 32849 2117 32905
rect 2173 32849 2201 32905
rect 2257 32849 2285 32905
rect 2341 32849 2369 32905
rect 2425 32849 2453 32905
rect 2509 32849 2537 32905
rect 2593 32849 2598 32905
rect 1938 32825 2598 32849
rect 1938 32769 1949 32825
rect 2005 32769 2033 32825
rect 2089 32769 2117 32825
rect 2173 32769 2201 32825
rect 2257 32769 2285 32825
rect 2341 32769 2369 32825
rect 2425 32769 2453 32825
rect 2509 32769 2537 32825
rect 2593 32769 2598 32825
rect 1938 32745 2598 32769
rect 1938 32689 1949 32745
rect 2005 32689 2033 32745
rect 2089 32689 2117 32745
rect 2173 32689 2201 32745
rect 2257 32689 2285 32745
rect 2341 32689 2369 32745
rect 2425 32689 2453 32745
rect 2509 32689 2537 32745
rect 2593 32689 2598 32745
rect 1938 32664 2598 32689
rect 1938 32608 1949 32664
rect 2005 32608 2033 32664
rect 2089 32608 2117 32664
rect 2173 32608 2201 32664
rect 2257 32608 2285 32664
rect 2341 32608 2369 32664
rect 2425 32608 2453 32664
rect 2509 32608 2537 32664
rect 2593 32608 2598 32664
rect 1938 32583 2598 32608
rect 1938 32527 1949 32583
rect 2005 32527 2033 32583
rect 2089 32527 2117 32583
rect 2173 32527 2201 32583
rect 2257 32527 2285 32583
rect 2341 32527 2369 32583
rect 2425 32527 2453 32583
rect 2509 32527 2537 32583
rect 2593 32527 2598 32583
rect 1938 32502 2598 32527
rect 1938 32446 1949 32502
rect 2005 32446 2033 32502
rect 2089 32446 2117 32502
rect 2173 32446 2201 32502
rect 2257 32446 2285 32502
rect 2341 32446 2369 32502
rect 2425 32446 2453 32502
rect 2509 32446 2537 32502
rect 2593 32446 2598 32502
rect 1938 32421 2598 32446
rect 1938 32365 1949 32421
rect 2005 32365 2033 32421
rect 2089 32365 2117 32421
rect 2173 32365 2201 32421
rect 2257 32365 2285 32421
rect 2341 32365 2369 32421
rect 2425 32365 2453 32421
rect 2509 32365 2537 32421
rect 2593 32365 2598 32421
rect 1938 32340 2598 32365
rect 1938 32284 1949 32340
rect 2005 32284 2033 32340
rect 2089 32284 2117 32340
rect 2173 32284 2201 32340
rect 2257 32284 2285 32340
rect 2341 32284 2369 32340
rect 2425 32284 2453 32340
rect 2509 32284 2537 32340
rect 2593 32284 2598 32340
rect 1938 32259 2598 32284
rect 1938 32203 1949 32259
rect 2005 32203 2033 32259
rect 2089 32203 2117 32259
rect 2173 32203 2201 32259
rect 2257 32203 2285 32259
rect 2341 32203 2369 32259
rect 2425 32203 2453 32259
rect 2509 32203 2537 32259
rect 2593 32203 2598 32259
rect 1938 32178 2598 32203
rect 1938 32122 1949 32178
rect 2005 32122 2033 32178
rect 2089 32122 2117 32178
rect 2173 32122 2201 32178
rect 2257 32122 2285 32178
rect 2341 32122 2369 32178
rect 2425 32122 2453 32178
rect 2509 32122 2537 32178
rect 2593 32122 2598 32178
rect 1938 32097 2598 32122
rect 1938 32041 1949 32097
rect 2005 32041 2033 32097
rect 2089 32041 2117 32097
rect 2173 32041 2201 32097
rect 2257 32041 2285 32097
rect 2341 32041 2369 32097
rect 2425 32041 2453 32097
rect 2509 32041 2537 32097
rect 2593 32041 2598 32097
rect 1938 32016 2598 32041
rect 1938 31960 1949 32016
rect 2005 31960 2033 32016
rect 2089 31960 2117 32016
rect 2173 31960 2201 32016
rect 2257 31960 2285 32016
rect 2341 31960 2369 32016
rect 2425 31960 2453 32016
rect 2509 31960 2537 32016
rect 2593 31960 2598 32016
rect 1938 31935 2598 31960
rect 1938 31879 1949 31935
rect 2005 31879 2033 31935
rect 2089 31879 2117 31935
rect 2173 31879 2201 31935
rect 2257 31879 2285 31935
rect 2341 31879 2369 31935
rect 2425 31879 2453 31935
rect 2509 31879 2537 31935
rect 2593 31879 2598 31935
rect 1938 31854 2598 31879
rect 1938 31798 1949 31854
rect 2005 31798 2033 31854
rect 2089 31798 2117 31854
rect 2173 31798 2201 31854
rect 2257 31798 2285 31854
rect 2341 31798 2369 31854
rect 2425 31798 2453 31854
rect 2509 31798 2537 31854
rect 2593 31798 2598 31854
rect 1938 31773 2598 31798
rect 1938 31717 1949 31773
rect 2005 31717 2033 31773
rect 2089 31717 2117 31773
rect 2173 31717 2201 31773
rect 2257 31717 2285 31773
rect 2341 31717 2369 31773
rect 2425 31717 2453 31773
rect 2509 31717 2537 31773
rect 2593 31717 2598 31773
rect 1938 31692 2598 31717
rect 1938 31636 1949 31692
rect 2005 31636 2033 31692
rect 2089 31636 2117 31692
rect 2173 31636 2201 31692
rect 2257 31636 2285 31692
rect 2341 31636 2369 31692
rect 2425 31636 2453 31692
rect 2509 31636 2537 31692
rect 2593 31636 2598 31692
rect 1938 31611 2598 31636
rect 1938 31555 1949 31611
rect 2005 31555 2033 31611
rect 2089 31555 2117 31611
rect 2173 31555 2201 31611
rect 2257 31555 2285 31611
rect 2341 31555 2369 31611
rect 2425 31555 2453 31611
rect 2509 31555 2537 31611
rect 2593 31555 2598 31611
rect 1938 31530 2598 31555
rect 1938 31474 1949 31530
rect 2005 31474 2033 31530
rect 2089 31474 2117 31530
rect 2173 31474 2201 31530
rect 2257 31474 2285 31530
rect 2341 31474 2369 31530
rect 2425 31474 2453 31530
rect 2509 31474 2537 31530
rect 2593 31474 2598 31530
rect 1938 31449 2598 31474
rect 1938 31393 1949 31449
rect 2005 31393 2033 31449
rect 2089 31393 2117 31449
rect 2173 31393 2201 31449
rect 2257 31393 2285 31449
rect 2341 31393 2369 31449
rect 2425 31393 2453 31449
rect 2509 31393 2537 31449
rect 2593 31393 2598 31449
rect 1938 31368 2598 31393
rect 1938 31312 1949 31368
rect 2005 31312 2033 31368
rect 2089 31312 2117 31368
rect 2173 31312 2201 31368
rect 2257 31312 2285 31368
rect 2341 31312 2369 31368
rect 2425 31312 2453 31368
rect 2509 31312 2537 31368
rect 2593 31312 2598 31368
rect 1938 31287 2598 31312
rect 1938 31231 1949 31287
rect 2005 31231 2033 31287
rect 2089 31231 2117 31287
rect 2173 31231 2201 31287
rect 2257 31231 2285 31287
rect 2341 31231 2369 31287
rect 2425 31231 2453 31287
rect 2509 31231 2537 31287
rect 2593 31231 2598 31287
rect 1938 31206 2598 31231
rect 1938 31150 1949 31206
rect 2005 31150 2033 31206
rect 2089 31150 2117 31206
rect 2173 31150 2201 31206
rect 2257 31150 2285 31206
rect 2341 31150 2369 31206
rect 2425 31150 2453 31206
rect 2509 31150 2537 31206
rect 2593 31150 2598 31206
rect 1938 31125 2598 31150
rect 1938 31069 1949 31125
rect 2005 31069 2033 31125
rect 2089 31069 2117 31125
rect 2173 31069 2201 31125
rect 2257 31069 2285 31125
rect 2341 31069 2369 31125
rect 2425 31069 2453 31125
rect 2509 31069 2537 31125
rect 2593 31069 2598 31125
rect 1938 31044 2598 31069
rect 1938 30988 1949 31044
rect 2005 30988 2033 31044
rect 2089 30988 2117 31044
rect 2173 30988 2201 31044
rect 2257 30988 2285 31044
rect 2341 30988 2369 31044
rect 2425 30988 2453 31044
rect 2509 30988 2537 31044
rect 2593 30988 2598 31044
rect 1938 30963 2598 30988
rect 1938 30907 1949 30963
rect 2005 30907 2033 30963
rect 2089 30907 2117 30963
rect 2173 30907 2201 30963
rect 2257 30907 2285 30963
rect 2341 30907 2369 30963
rect 2425 30907 2453 30963
rect 2509 30907 2537 30963
rect 2593 30907 2598 30963
rect 1938 30882 2598 30907
rect 1938 30826 1949 30882
rect 2005 30826 2033 30882
rect 2089 30826 2117 30882
rect 2173 30826 2201 30882
rect 2257 30826 2285 30882
rect 2341 30826 2369 30882
rect 2425 30826 2453 30882
rect 2509 30826 2537 30882
rect 2593 30826 2598 30882
rect 1938 30801 2598 30826
rect 1938 30745 1949 30801
rect 2005 30745 2033 30801
rect 2089 30745 2117 30801
rect 2173 30745 2201 30801
rect 2257 30745 2285 30801
rect 2341 30745 2369 30801
rect 2425 30745 2453 30801
rect 2509 30745 2537 30801
rect 2593 30745 2598 30801
rect 1938 30720 2598 30745
rect 1938 30664 1949 30720
rect 2005 30664 2033 30720
rect 2089 30664 2117 30720
rect 2173 30664 2201 30720
rect 2257 30664 2285 30720
rect 2341 30664 2369 30720
rect 2425 30664 2453 30720
rect 2509 30664 2537 30720
rect 2593 30664 2598 30720
rect 1938 30639 2598 30664
rect 1938 30583 1949 30639
rect 2005 30583 2033 30639
rect 2089 30583 2117 30639
rect 2173 30583 2201 30639
rect 2257 30583 2285 30639
rect 2341 30583 2369 30639
rect 2425 30583 2453 30639
rect 2509 30583 2537 30639
rect 2593 30583 2598 30639
rect 1938 30558 2598 30583
rect 1938 30502 1949 30558
rect 2005 30502 2033 30558
rect 2089 30502 2117 30558
rect 2173 30502 2201 30558
rect 2257 30502 2285 30558
rect 2341 30502 2369 30558
rect 2425 30502 2453 30558
rect 2509 30502 2537 30558
rect 2593 30502 2598 30558
rect 1938 30477 2598 30502
rect 1938 30421 1949 30477
rect 2005 30421 2033 30477
rect 2089 30421 2117 30477
rect 2173 30421 2201 30477
rect 2257 30421 2285 30477
rect 2341 30421 2369 30477
rect 2425 30421 2453 30477
rect 2509 30421 2537 30477
rect 2593 30421 2598 30477
rect 1938 30396 2598 30421
rect 1938 30340 1949 30396
rect 2005 30340 2033 30396
rect 2089 30340 2117 30396
rect 2173 30340 2201 30396
rect 2257 30340 2285 30396
rect 2341 30340 2369 30396
rect 2425 30340 2453 30396
rect 2509 30340 2537 30396
rect 2593 30340 2598 30396
rect 1938 30315 2598 30340
rect 1938 30259 1949 30315
rect 2005 30259 2033 30315
rect 2089 30259 2117 30315
rect 2173 30259 2201 30315
rect 2257 30259 2285 30315
rect 2341 30259 2369 30315
rect 2425 30259 2453 30315
rect 2509 30259 2537 30315
rect 2593 30259 2598 30315
rect 1938 30234 2598 30259
tri 1929 30178 1938 30187 se
rect 1938 30178 1949 30234
rect 2005 30178 2033 30234
rect 2089 30178 2117 30234
rect 2173 30178 2201 30234
rect 2257 30178 2285 30234
rect 2341 30178 2369 30234
rect 2425 30178 2453 30234
rect 2509 30178 2537 30234
rect 2593 30178 2598 30234
tri 1906 30155 1929 30178 se
rect 1929 30155 2598 30178
tri 1850 30099 1906 30155 se
rect 1906 30099 2598 30155
tri 1826 30075 1850 30099 se
rect 1850 30075 2598 30099
tri 1804 30053 1826 30075 se
rect 1826 30053 2598 30075
tri 1770 30019 1804 30053 se
rect 1804 30019 2598 30053
tri 1731 29980 1770 30019 se
rect 1770 29997 2598 30019
rect 1770 29980 2581 29997
tri 2581 29980 2598 29997 nw
rect 2734 35032 3666 35132
rect 2734 35014 2853 35032
tri 2853 35014 2871 35032 nw
tri 3529 35014 3547 35032 ne
rect 3547 35014 3666 35032
rect 2734 34990 2829 35014
tri 2829 34990 2853 35014 nw
tri 3547 34990 3571 35014 ne
rect 3571 34990 3666 35014
tri 1660 29909 1731 29980 se
rect 1731 29909 2510 29980
tri 2510 29909 2581 29980 nw
tri 2663 29909 2734 29980 se
rect 2734 29952 2800 34990
tri 2800 34961 2829 34990 nw
tri 3571 34961 3600 34990 ne
rect 2734 29909 2757 29952
tri 2757 29909 2800 29952 nw
rect 2900 34795 3500 34804
rect 2900 34739 2915 34795
rect 2971 34739 3001 34795
rect 3057 34739 3087 34795
rect 3143 34739 3173 34795
rect 3229 34739 3259 34795
rect 3315 34739 3345 34795
rect 3401 34739 3431 34795
rect 3487 34739 3500 34795
rect 2900 34715 3500 34739
rect 2900 34659 2915 34715
rect 2971 34659 3001 34715
rect 3057 34659 3087 34715
rect 3143 34659 3173 34715
rect 3229 34659 3259 34715
rect 3315 34659 3345 34715
rect 3401 34659 3431 34715
rect 3487 34659 3500 34715
rect 2900 34635 3500 34659
rect 2900 34579 2915 34635
rect 2971 34579 3001 34635
rect 3057 34579 3087 34635
rect 3143 34579 3173 34635
rect 3229 34579 3259 34635
rect 3315 34579 3345 34635
rect 3401 34579 3431 34635
rect 3487 34579 3500 34635
rect 2900 34555 3500 34579
rect 2900 34499 2915 34555
rect 2971 34499 3001 34555
rect 3057 34499 3087 34555
rect 3143 34499 3173 34555
rect 3229 34499 3259 34555
rect 3315 34499 3345 34555
rect 3401 34499 3431 34555
rect 3487 34499 3500 34555
rect 2900 34475 3500 34499
rect 2900 34419 2915 34475
rect 2971 34419 3001 34475
rect 3057 34419 3087 34475
rect 3143 34419 3173 34475
rect 3229 34419 3259 34475
rect 3315 34419 3345 34475
rect 3401 34419 3431 34475
rect 3487 34419 3500 34475
rect 2900 34395 3500 34419
rect 2900 34339 2915 34395
rect 2971 34339 3001 34395
rect 3057 34339 3087 34395
rect 3143 34339 3173 34395
rect 3229 34339 3259 34395
rect 3315 34339 3345 34395
rect 3401 34339 3431 34395
rect 3487 34339 3500 34395
rect 2900 34315 3500 34339
rect 2900 34259 2915 34315
rect 2971 34259 3001 34315
rect 3057 34259 3087 34315
rect 3143 34259 3173 34315
rect 3229 34259 3259 34315
rect 3315 34259 3345 34315
rect 3401 34259 3431 34315
rect 3487 34259 3500 34315
rect 2900 34235 3500 34259
rect 2900 34179 2915 34235
rect 2971 34179 3001 34235
rect 3057 34179 3087 34235
rect 3143 34179 3173 34235
rect 3229 34179 3259 34235
rect 3315 34179 3345 34235
rect 3401 34179 3431 34235
rect 3487 34179 3500 34235
rect 2900 34155 3500 34179
rect 2900 34099 2915 34155
rect 2971 34099 3001 34155
rect 3057 34099 3087 34155
rect 3143 34099 3173 34155
rect 3229 34099 3259 34155
rect 3315 34099 3345 34155
rect 3401 34099 3431 34155
rect 3487 34099 3500 34155
rect 2900 34075 3500 34099
rect 2900 34019 2915 34075
rect 2971 34019 3001 34075
rect 3057 34019 3087 34075
rect 3143 34019 3173 34075
rect 3229 34019 3259 34075
rect 3315 34019 3345 34075
rect 3401 34019 3431 34075
rect 3487 34019 3500 34075
rect 2900 33995 3500 34019
rect 2900 33939 2915 33995
rect 2971 33939 3001 33995
rect 3057 33939 3087 33995
rect 3143 33939 3173 33995
rect 3229 33939 3259 33995
rect 3315 33939 3345 33995
rect 3401 33939 3431 33995
rect 3487 33939 3500 33995
rect 2900 33915 3500 33939
rect 2900 33859 2915 33915
rect 2971 33859 3001 33915
rect 3057 33859 3087 33915
rect 3143 33859 3173 33915
rect 3229 33859 3259 33915
rect 3315 33859 3345 33915
rect 3401 33859 3431 33915
rect 3487 33859 3500 33915
rect 2900 33835 3500 33859
rect 2900 33779 2915 33835
rect 2971 33779 3001 33835
rect 3057 33779 3087 33835
rect 3143 33779 3173 33835
rect 3229 33779 3259 33835
rect 3315 33779 3345 33835
rect 3401 33779 3431 33835
rect 3487 33779 3500 33835
rect 2900 33755 3500 33779
rect 2900 33699 2915 33755
rect 2971 33699 3001 33755
rect 3057 33699 3087 33755
rect 3143 33699 3173 33755
rect 3229 33699 3259 33755
rect 3315 33699 3345 33755
rect 3401 33699 3431 33755
rect 3487 33699 3500 33755
rect 2900 33675 3500 33699
rect 2900 33619 2915 33675
rect 2971 33619 3001 33675
rect 3057 33619 3087 33675
rect 3143 33619 3173 33675
rect 3229 33619 3259 33675
rect 3315 33619 3345 33675
rect 3401 33619 3431 33675
rect 3487 33619 3500 33675
rect 2900 33595 3500 33619
rect 2900 33539 2915 33595
rect 2971 33539 3001 33595
rect 3057 33539 3087 33595
rect 3143 33539 3173 33595
rect 3229 33539 3259 33595
rect 3315 33539 3345 33595
rect 3401 33539 3431 33595
rect 3487 33539 3500 33595
rect 2900 33515 3500 33539
rect 2900 33459 2915 33515
rect 2971 33459 3001 33515
rect 3057 33459 3087 33515
rect 3143 33459 3173 33515
rect 3229 33459 3259 33515
rect 3315 33459 3345 33515
rect 3401 33459 3431 33515
rect 3487 33459 3500 33515
rect 2900 33435 3500 33459
rect 2900 33379 2915 33435
rect 2971 33379 3001 33435
rect 3057 33379 3087 33435
rect 3143 33379 3173 33435
rect 3229 33379 3259 33435
rect 3315 33379 3345 33435
rect 3401 33379 3431 33435
rect 3487 33379 3500 33435
rect 2900 33355 3500 33379
rect 2900 33299 2915 33355
rect 2971 33299 3001 33355
rect 3057 33299 3087 33355
rect 3143 33299 3173 33355
rect 3229 33299 3259 33355
rect 3315 33299 3345 33355
rect 3401 33299 3431 33355
rect 3487 33299 3500 33355
rect 2900 33275 3500 33299
rect 2900 33219 2915 33275
rect 2971 33219 3001 33275
rect 3057 33219 3087 33275
rect 3143 33219 3173 33275
rect 3229 33219 3259 33275
rect 3315 33219 3345 33275
rect 3401 33219 3431 33275
rect 3487 33219 3500 33275
rect 2900 33195 3500 33219
rect 2900 33139 2915 33195
rect 2971 33139 3001 33195
rect 3057 33139 3087 33195
rect 3143 33139 3173 33195
rect 3229 33139 3259 33195
rect 3315 33139 3345 33195
rect 3401 33139 3431 33195
rect 3487 33139 3500 33195
rect 2900 33115 3500 33139
rect 2900 33059 2915 33115
rect 2971 33059 3001 33115
rect 3057 33059 3087 33115
rect 3143 33059 3173 33115
rect 3229 33059 3259 33115
rect 3315 33059 3345 33115
rect 3401 33059 3431 33115
rect 3487 33059 3500 33115
rect 2900 33035 3500 33059
rect 2900 32979 2915 33035
rect 2971 32979 3001 33035
rect 3057 32979 3087 33035
rect 3143 32979 3173 33035
rect 3229 32979 3259 33035
rect 3315 32979 3345 33035
rect 3401 32979 3431 33035
rect 3487 32979 3500 33035
rect 2900 32955 3500 32979
rect 2900 32899 2915 32955
rect 2971 32899 3001 32955
rect 3057 32899 3087 32955
rect 3143 32899 3173 32955
rect 3229 32899 3259 32955
rect 3315 32899 3345 32955
rect 3401 32899 3431 32955
rect 3487 32899 3500 32955
rect 2900 32875 3500 32899
rect 2900 32819 2915 32875
rect 2971 32819 3001 32875
rect 3057 32819 3087 32875
rect 3143 32819 3173 32875
rect 3229 32819 3259 32875
rect 3315 32819 3345 32875
rect 3401 32819 3431 32875
rect 3487 32819 3500 32875
rect 2900 32795 3500 32819
rect 2900 32739 2915 32795
rect 2971 32739 3001 32795
rect 3057 32739 3087 32795
rect 3143 32739 3173 32795
rect 3229 32739 3259 32795
rect 3315 32739 3345 32795
rect 3401 32739 3431 32795
rect 3487 32739 3500 32795
rect 2900 32715 3500 32739
rect 2900 32659 2915 32715
rect 2971 32659 3001 32715
rect 3057 32659 3087 32715
rect 3143 32659 3173 32715
rect 3229 32659 3259 32715
rect 3315 32659 3345 32715
rect 3401 32659 3431 32715
rect 3487 32659 3500 32715
rect 2900 32635 3500 32659
rect 2900 32579 2915 32635
rect 2971 32579 3001 32635
rect 3057 32579 3087 32635
rect 3143 32579 3173 32635
rect 3229 32579 3259 32635
rect 3315 32579 3345 32635
rect 3401 32579 3431 32635
rect 3487 32579 3500 32635
rect 2900 32555 3500 32579
rect 2900 32499 2915 32555
rect 2971 32499 3001 32555
rect 3057 32499 3087 32555
rect 3143 32499 3173 32555
rect 3229 32499 3259 32555
rect 3315 32499 3345 32555
rect 3401 32499 3431 32555
rect 3487 32499 3500 32555
rect 2900 32475 3500 32499
rect 2900 32419 2915 32475
rect 2971 32419 3001 32475
rect 3057 32419 3087 32475
rect 3143 32419 3173 32475
rect 3229 32419 3259 32475
rect 3315 32419 3345 32475
rect 3401 32419 3431 32475
rect 3487 32419 3500 32475
rect 2900 32395 3500 32419
rect 2900 32339 2915 32395
rect 2971 32339 3001 32395
rect 3057 32339 3087 32395
rect 3143 32339 3173 32395
rect 3229 32339 3259 32395
rect 3315 32339 3345 32395
rect 3401 32339 3431 32395
rect 3487 32339 3500 32395
rect 2900 32315 3500 32339
rect 2900 32259 2915 32315
rect 2971 32259 3001 32315
rect 3057 32259 3087 32315
rect 3143 32259 3173 32315
rect 3229 32259 3259 32315
rect 3315 32259 3345 32315
rect 3401 32259 3431 32315
rect 3487 32259 3500 32315
rect 2900 32235 3500 32259
rect 2900 32179 2915 32235
rect 2971 32179 3001 32235
rect 3057 32179 3087 32235
rect 3143 32179 3173 32235
rect 3229 32179 3259 32235
rect 3315 32179 3345 32235
rect 3401 32179 3431 32235
rect 3487 32179 3500 32235
rect 2900 32155 3500 32179
rect 2900 32099 2915 32155
rect 2971 32099 3001 32155
rect 3057 32099 3087 32155
rect 3143 32099 3173 32155
rect 3229 32099 3259 32155
rect 3315 32099 3345 32155
rect 3401 32099 3431 32155
rect 3487 32099 3500 32155
rect 2900 32075 3500 32099
rect 2900 32019 2915 32075
rect 2971 32019 3001 32075
rect 3057 32019 3087 32075
rect 3143 32019 3173 32075
rect 3229 32019 3259 32075
rect 3315 32019 3345 32075
rect 3401 32019 3431 32075
rect 3487 32019 3500 32075
rect 2900 31995 3500 32019
rect 2900 31939 2915 31995
rect 2971 31939 3001 31995
rect 3057 31939 3087 31995
rect 3143 31939 3173 31995
rect 3229 31939 3259 31995
rect 3315 31939 3345 31995
rect 3401 31939 3431 31995
rect 3487 31939 3500 31995
rect 2900 31915 3500 31939
rect 2900 31859 2915 31915
rect 2971 31859 3001 31915
rect 3057 31859 3087 31915
rect 3143 31859 3173 31915
rect 3229 31859 3259 31915
rect 3315 31859 3345 31915
rect 3401 31859 3431 31915
rect 3487 31859 3500 31915
rect 2900 31835 3500 31859
rect 2900 31779 2915 31835
rect 2971 31779 3001 31835
rect 3057 31779 3087 31835
rect 3143 31779 3173 31835
rect 3229 31779 3259 31835
rect 3315 31779 3345 31835
rect 3401 31779 3431 31835
rect 3487 31779 3500 31835
rect 2900 31755 3500 31779
rect 2900 31699 2915 31755
rect 2971 31699 3001 31755
rect 3057 31699 3087 31755
rect 3143 31699 3173 31755
rect 3229 31699 3259 31755
rect 3315 31699 3345 31755
rect 3401 31699 3431 31755
rect 3487 31699 3500 31755
rect 2900 31675 3500 31699
rect 2900 31619 2915 31675
rect 2971 31619 3001 31675
rect 3057 31619 3087 31675
rect 3143 31619 3173 31675
rect 3229 31619 3259 31675
rect 3315 31619 3345 31675
rect 3401 31619 3431 31675
rect 3487 31619 3500 31675
rect 2900 31595 3500 31619
rect 2900 31539 2915 31595
rect 2971 31539 3001 31595
rect 3057 31539 3087 31595
rect 3143 31539 3173 31595
rect 3229 31539 3259 31595
rect 3315 31539 3345 31595
rect 3401 31539 3431 31595
rect 3487 31539 3500 31595
rect 2900 31515 3500 31539
rect 2900 31459 2915 31515
rect 2971 31459 3001 31515
rect 3057 31459 3087 31515
rect 3143 31459 3173 31515
rect 3229 31459 3259 31515
rect 3315 31459 3345 31515
rect 3401 31459 3431 31515
rect 3487 31459 3500 31515
rect 2900 31435 3500 31459
rect 2900 31379 2915 31435
rect 2971 31379 3001 31435
rect 3057 31379 3087 31435
rect 3143 31379 3173 31435
rect 3229 31379 3259 31435
rect 3315 31379 3345 31435
rect 3401 31379 3431 31435
rect 3487 31379 3500 31435
rect 2900 31355 3500 31379
rect 2900 31299 2915 31355
rect 2971 31299 3001 31355
rect 3057 31299 3087 31355
rect 3143 31299 3173 31355
rect 3229 31299 3259 31355
rect 3315 31299 3345 31355
rect 3401 31299 3431 31355
rect 3487 31299 3500 31355
rect 2900 31275 3500 31299
rect 2900 31219 2915 31275
rect 2971 31219 3001 31275
rect 3057 31219 3087 31275
rect 3143 31219 3173 31275
rect 3229 31219 3259 31275
rect 3315 31219 3345 31275
rect 3401 31219 3431 31275
rect 3487 31219 3500 31275
rect 2900 31195 3500 31219
rect 2900 31139 2915 31195
rect 2971 31139 3001 31195
rect 3057 31139 3087 31195
rect 3143 31139 3173 31195
rect 3229 31139 3259 31195
rect 3315 31139 3345 31195
rect 3401 31139 3431 31195
rect 3487 31139 3500 31195
rect 2900 31115 3500 31139
rect 2900 31059 2915 31115
rect 2971 31059 3001 31115
rect 3057 31059 3087 31115
rect 3143 31059 3173 31115
rect 3229 31059 3259 31115
rect 3315 31059 3345 31115
rect 3401 31059 3431 31115
rect 3487 31059 3500 31115
rect 2900 31035 3500 31059
rect 2900 30979 2915 31035
rect 2971 30979 3001 31035
rect 3057 30979 3087 31035
rect 3143 30979 3173 31035
rect 3229 30979 3259 31035
rect 3315 30979 3345 31035
rect 3401 30979 3431 31035
rect 3487 30979 3500 31035
rect 2900 30955 3500 30979
rect 2900 30899 2915 30955
rect 2971 30899 3001 30955
rect 3057 30899 3087 30955
rect 3143 30899 3173 30955
rect 3229 30899 3259 30955
rect 3315 30899 3345 30955
rect 3401 30899 3431 30955
rect 3487 30899 3500 30955
rect 2900 30875 3500 30899
rect 2900 30819 2915 30875
rect 2971 30819 3001 30875
rect 3057 30819 3087 30875
rect 3143 30819 3173 30875
rect 3229 30819 3259 30875
rect 3315 30819 3345 30875
rect 3401 30819 3431 30875
rect 3487 30819 3500 30875
rect 2900 30795 3500 30819
rect 2900 30739 2915 30795
rect 2971 30739 3001 30795
rect 3057 30739 3087 30795
rect 3143 30739 3173 30795
rect 3229 30739 3259 30795
rect 3315 30739 3345 30795
rect 3401 30739 3431 30795
rect 3487 30739 3500 30795
rect 2900 30715 3500 30739
rect 2900 30659 2915 30715
rect 2971 30659 3001 30715
rect 3057 30659 3087 30715
rect 3143 30659 3173 30715
rect 3229 30659 3259 30715
rect 3315 30659 3345 30715
rect 3401 30659 3431 30715
rect 3487 30659 3500 30715
rect 2900 30635 3500 30659
rect 2900 30579 2915 30635
rect 2971 30579 3001 30635
rect 3057 30579 3087 30635
rect 3143 30579 3173 30635
rect 3229 30579 3259 30635
rect 3315 30579 3345 30635
rect 3401 30579 3431 30635
rect 3487 30579 3500 30635
rect 2900 30555 3500 30579
rect 2900 30499 2915 30555
rect 2971 30499 3001 30555
rect 3057 30499 3087 30555
rect 3143 30499 3173 30555
rect 3229 30499 3259 30555
rect 3315 30499 3345 30555
rect 3401 30499 3431 30555
rect 3487 30499 3500 30555
rect 2900 30475 3500 30499
rect 2900 30419 2915 30475
rect 2971 30419 3001 30475
rect 3057 30419 3087 30475
rect 3143 30419 3173 30475
rect 3229 30419 3259 30475
rect 3315 30419 3345 30475
rect 3401 30419 3431 30475
rect 3487 30419 3500 30475
rect 2900 30395 3500 30419
rect 2900 30339 2915 30395
rect 2971 30339 3001 30395
rect 3057 30339 3087 30395
rect 3143 30339 3173 30395
rect 3229 30339 3259 30395
rect 3315 30339 3345 30395
rect 3401 30339 3431 30395
rect 3487 30339 3500 30395
rect 2900 30315 3500 30339
rect 2900 30259 2915 30315
rect 2971 30259 3001 30315
rect 3057 30259 3087 30315
rect 3143 30259 3173 30315
rect 3229 30259 3259 30315
rect 3315 30259 3345 30315
rect 3401 30259 3431 30315
rect 3487 30259 3500 30315
rect 2900 30235 3500 30259
rect 2900 30179 2915 30235
rect 2971 30179 3001 30235
rect 3057 30179 3087 30235
rect 3143 30179 3173 30235
rect 3229 30179 3259 30235
rect 3315 30179 3345 30235
rect 3401 30179 3431 30235
rect 3487 30179 3500 30235
rect 2900 30155 3500 30179
rect 2900 30099 2915 30155
rect 2971 30099 3001 30155
rect 3057 30099 3087 30155
rect 3143 30099 3173 30155
rect 3229 30099 3259 30155
rect 3315 30099 3345 30155
rect 3401 30099 3431 30155
rect 3487 30099 3500 30155
rect 2900 30075 3500 30099
rect 2900 30019 2915 30075
rect 2971 30019 3001 30075
rect 3057 30019 3087 30075
rect 3143 30019 3173 30075
rect 3229 30019 3259 30075
rect 3315 30019 3345 30075
rect 3401 30019 3431 30075
rect 3487 30019 3500 30075
tri 1637 29886 1660 29909 se
rect 1660 29886 2487 29909
tri 2487 29886 2510 29909 nw
tri 2640 29886 2663 29909 se
rect 2663 29886 2734 29909
tri 2734 29886 2757 29909 nw
tri 2877 29886 2900 29909 se
rect 2900 29886 3500 30019
tri 1543 29792 1637 29886 se
rect 1637 29844 2445 29886
tri 2445 29844 2487 29886 nw
tri 2598 29844 2640 29886 se
rect 2640 29844 2671 29886
rect 1637 29792 2393 29844
tri 2393 29792 2445 29844 nw
tri 2546 29792 2598 29844 se
rect 2598 29823 2671 29844
tri 2671 29823 2734 29886 nw
tri 2814 29823 2877 29886 se
rect 2877 29823 3500 29886
rect 2598 29792 2640 29823
tri 2640 29792 2671 29823 nw
tri 2783 29792 2814 29823 se
rect 2814 29792 3500 29823
tri 1449 29698 1543 29792 se
rect 1543 29698 2299 29792
tri 2299 29698 2393 29792 nw
tri 2452 29698 2546 29792 se
rect 2546 29750 2598 29792
tri 2598 29750 2640 29792 nw
tri 2741 29750 2783 29792 se
rect 2783 29750 3500 29792
tri 2546 29698 2598 29750 nw
tri 2689 29698 2741 29750 se
rect 2741 29698 3500 29750
tri 1431 29680 1449 29698 se
rect 1449 29680 2281 29698
tri 2281 29680 2299 29698 nw
tri 2434 29680 2452 29698 se
rect 2452 29680 2528 29698
tri 2528 29680 2546 29698 nw
tri 2671 29680 2689 29698 se
rect 2689 29680 3500 29698
tri 1355 29604 1431 29680 se
rect 1431 29604 2205 29680
tri 2205 29604 2281 29680 nw
tri 2358 29604 2434 29680 se
rect 2434 29604 2452 29680
tri 2452 29604 2528 29680 nw
tri 2603 29612 2671 29680 se
rect 2671 29659 3500 29680
rect 2671 29612 3453 29659
tri 3453 29612 3500 29659 nw
tri 2598 29607 2603 29612 se
rect 2603 29607 3445 29612
tri 2595 29604 2598 29607 se
rect 2598 29604 3445 29607
tri 3445 29604 3453 29612 nw
tri 3592 29604 3600 29612 se
rect 3600 29604 3666 34990
tri 1261 29510 1355 29604 se
rect 1355 29510 2111 29604
tri 2111 29510 2205 29604 nw
tri 2264 29510 2358 29604 se
tri 2358 29510 2452 29604 nw
tri 2509 29518 2595 29604 se
rect 2595 29518 3359 29604
tri 3359 29518 3445 29604 nw
tri 3506 29518 3592 29604 se
rect 3592 29584 3666 29604
rect 3592 29518 3600 29584
tri 3600 29518 3666 29584 nw
rect 5723 35032 6655 35132
rect 5723 35014 5842 35032
tri 5842 35014 5860 35032 nw
tri 6518 35014 6536 35032 ne
rect 6536 35014 6655 35032
rect 5723 34990 5818 35014
tri 5818 34990 5842 35014 nw
tri 6536 34990 6560 35014 ne
rect 6560 34990 6655 35014
rect 5723 29584 5789 34990
tri 5789 34961 5818 34990 nw
tri 6560 34961 6589 34990 ne
rect 5889 34795 6489 34804
rect 5889 34739 5905 34795
rect 5961 34739 5991 34795
rect 6047 34739 6077 34795
rect 6133 34739 6163 34795
rect 6219 34739 6249 34795
rect 6305 34739 6335 34795
rect 6391 34739 6421 34795
rect 6477 34739 6489 34795
rect 5889 34715 6489 34739
rect 5889 34659 5905 34715
rect 5961 34659 5991 34715
rect 6047 34659 6077 34715
rect 6133 34659 6163 34715
rect 6219 34659 6249 34715
rect 6305 34659 6335 34715
rect 6391 34659 6421 34715
rect 6477 34659 6489 34715
rect 5889 34635 6489 34659
rect 5889 34579 5905 34635
rect 5961 34579 5991 34635
rect 6047 34579 6077 34635
rect 6133 34579 6163 34635
rect 6219 34579 6249 34635
rect 6305 34579 6335 34635
rect 6391 34579 6421 34635
rect 6477 34579 6489 34635
rect 5889 34555 6489 34579
rect 5889 34499 5905 34555
rect 5961 34499 5991 34555
rect 6047 34499 6077 34555
rect 6133 34499 6163 34555
rect 6219 34499 6249 34555
rect 6305 34499 6335 34555
rect 6391 34499 6421 34555
rect 6477 34499 6489 34555
rect 5889 34475 6489 34499
rect 5889 34419 5905 34475
rect 5961 34419 5991 34475
rect 6047 34419 6077 34475
rect 6133 34419 6163 34475
rect 6219 34419 6249 34475
rect 6305 34419 6335 34475
rect 6391 34419 6421 34475
rect 6477 34419 6489 34475
rect 5889 34395 6489 34419
rect 5889 34339 5905 34395
rect 5961 34339 5991 34395
rect 6047 34339 6077 34395
rect 6133 34339 6163 34395
rect 6219 34339 6249 34395
rect 6305 34339 6335 34395
rect 6391 34339 6421 34395
rect 6477 34339 6489 34395
rect 5889 34315 6489 34339
rect 5889 34259 5905 34315
rect 5961 34259 5991 34315
rect 6047 34259 6077 34315
rect 6133 34259 6163 34315
rect 6219 34259 6249 34315
rect 6305 34259 6335 34315
rect 6391 34259 6421 34315
rect 6477 34259 6489 34315
rect 5889 34235 6489 34259
rect 5889 34179 5905 34235
rect 5961 34179 5991 34235
rect 6047 34179 6077 34235
rect 6133 34179 6163 34235
rect 6219 34179 6249 34235
rect 6305 34179 6335 34235
rect 6391 34179 6421 34235
rect 6477 34179 6489 34235
rect 5889 34155 6489 34179
rect 5889 34099 5905 34155
rect 5961 34099 5991 34155
rect 6047 34099 6077 34155
rect 6133 34099 6163 34155
rect 6219 34099 6249 34155
rect 6305 34099 6335 34155
rect 6391 34099 6421 34155
rect 6477 34099 6489 34155
rect 5889 34075 6489 34099
rect 5889 34019 5905 34075
rect 5961 34019 5991 34075
rect 6047 34019 6077 34075
rect 6133 34019 6163 34075
rect 6219 34019 6249 34075
rect 6305 34019 6335 34075
rect 6391 34019 6421 34075
rect 6477 34019 6489 34075
rect 5889 33995 6489 34019
rect 5889 33939 5905 33995
rect 5961 33939 5991 33995
rect 6047 33939 6077 33995
rect 6133 33939 6163 33995
rect 6219 33939 6249 33995
rect 6305 33939 6335 33995
rect 6391 33939 6421 33995
rect 6477 33939 6489 33995
rect 5889 33915 6489 33939
rect 5889 33859 5905 33915
rect 5961 33859 5991 33915
rect 6047 33859 6077 33915
rect 6133 33859 6163 33915
rect 6219 33859 6249 33915
rect 6305 33859 6335 33915
rect 6391 33859 6421 33915
rect 6477 33859 6489 33915
rect 5889 33835 6489 33859
rect 5889 33779 5905 33835
rect 5961 33779 5991 33835
rect 6047 33779 6077 33835
rect 6133 33779 6163 33835
rect 6219 33779 6249 33835
rect 6305 33779 6335 33835
rect 6391 33779 6421 33835
rect 6477 33779 6489 33835
rect 5889 33755 6489 33779
rect 5889 33699 5905 33755
rect 5961 33699 5991 33755
rect 6047 33699 6077 33755
rect 6133 33699 6163 33755
rect 6219 33699 6249 33755
rect 6305 33699 6335 33755
rect 6391 33699 6421 33755
rect 6477 33699 6489 33755
rect 5889 33675 6489 33699
rect 5889 33619 5905 33675
rect 5961 33619 5991 33675
rect 6047 33619 6077 33675
rect 6133 33619 6163 33675
rect 6219 33619 6249 33675
rect 6305 33619 6335 33675
rect 6391 33619 6421 33675
rect 6477 33619 6489 33675
rect 5889 33595 6489 33619
rect 5889 33539 5905 33595
rect 5961 33539 5991 33595
rect 6047 33539 6077 33595
rect 6133 33539 6163 33595
rect 6219 33539 6249 33595
rect 6305 33539 6335 33595
rect 6391 33539 6421 33595
rect 6477 33539 6489 33595
rect 5889 33515 6489 33539
rect 5889 33459 5905 33515
rect 5961 33459 5991 33515
rect 6047 33459 6077 33515
rect 6133 33459 6163 33515
rect 6219 33459 6249 33515
rect 6305 33459 6335 33515
rect 6391 33459 6421 33515
rect 6477 33459 6489 33515
rect 5889 33435 6489 33459
rect 5889 33379 5905 33435
rect 5961 33379 5991 33435
rect 6047 33379 6077 33435
rect 6133 33379 6163 33435
rect 6219 33379 6249 33435
rect 6305 33379 6335 33435
rect 6391 33379 6421 33435
rect 6477 33379 6489 33435
rect 5889 33355 6489 33379
rect 5889 33299 5905 33355
rect 5961 33299 5991 33355
rect 6047 33299 6077 33355
rect 6133 33299 6163 33355
rect 6219 33299 6249 33355
rect 6305 33299 6335 33355
rect 6391 33299 6421 33355
rect 6477 33299 6489 33355
rect 5889 33275 6489 33299
rect 5889 33219 5905 33275
rect 5961 33219 5991 33275
rect 6047 33219 6077 33275
rect 6133 33219 6163 33275
rect 6219 33219 6249 33275
rect 6305 33219 6335 33275
rect 6391 33219 6421 33275
rect 6477 33219 6489 33275
rect 5889 33195 6489 33219
rect 5889 33139 5905 33195
rect 5961 33139 5991 33195
rect 6047 33139 6077 33195
rect 6133 33139 6163 33195
rect 6219 33139 6249 33195
rect 6305 33139 6335 33195
rect 6391 33139 6421 33195
rect 6477 33139 6489 33195
rect 5889 33115 6489 33139
rect 5889 33059 5905 33115
rect 5961 33059 5991 33115
rect 6047 33059 6077 33115
rect 6133 33059 6163 33115
rect 6219 33059 6249 33115
rect 6305 33059 6335 33115
rect 6391 33059 6421 33115
rect 6477 33059 6489 33115
rect 5889 33035 6489 33059
rect 5889 32979 5905 33035
rect 5961 32979 5991 33035
rect 6047 32979 6077 33035
rect 6133 32979 6163 33035
rect 6219 32979 6249 33035
rect 6305 32979 6335 33035
rect 6391 32979 6421 33035
rect 6477 32979 6489 33035
rect 5889 32955 6489 32979
rect 5889 32899 5905 32955
rect 5961 32899 5991 32955
rect 6047 32899 6077 32955
rect 6133 32899 6163 32955
rect 6219 32899 6249 32955
rect 6305 32899 6335 32955
rect 6391 32899 6421 32955
rect 6477 32899 6489 32955
rect 5889 32875 6489 32899
rect 5889 32819 5905 32875
rect 5961 32819 5991 32875
rect 6047 32819 6077 32875
rect 6133 32819 6163 32875
rect 6219 32819 6249 32875
rect 6305 32819 6335 32875
rect 6391 32819 6421 32875
rect 6477 32819 6489 32875
rect 5889 32795 6489 32819
rect 5889 32739 5905 32795
rect 5961 32739 5991 32795
rect 6047 32739 6077 32795
rect 6133 32739 6163 32795
rect 6219 32739 6249 32795
rect 6305 32739 6335 32795
rect 6391 32739 6421 32795
rect 6477 32739 6489 32795
rect 5889 32715 6489 32739
rect 5889 32659 5905 32715
rect 5961 32659 5991 32715
rect 6047 32659 6077 32715
rect 6133 32659 6163 32715
rect 6219 32659 6249 32715
rect 6305 32659 6335 32715
rect 6391 32659 6421 32715
rect 6477 32659 6489 32715
rect 5889 32635 6489 32659
rect 5889 32579 5905 32635
rect 5961 32579 5991 32635
rect 6047 32579 6077 32635
rect 6133 32579 6163 32635
rect 6219 32579 6249 32635
rect 6305 32579 6335 32635
rect 6391 32579 6421 32635
rect 6477 32579 6489 32635
rect 5889 32555 6489 32579
rect 5889 32499 5905 32555
rect 5961 32499 5991 32555
rect 6047 32499 6077 32555
rect 6133 32499 6163 32555
rect 6219 32499 6249 32555
rect 6305 32499 6335 32555
rect 6391 32499 6421 32555
rect 6477 32499 6489 32555
rect 5889 32475 6489 32499
rect 5889 32419 5905 32475
rect 5961 32419 5991 32475
rect 6047 32419 6077 32475
rect 6133 32419 6163 32475
rect 6219 32419 6249 32475
rect 6305 32419 6335 32475
rect 6391 32419 6421 32475
rect 6477 32419 6489 32475
rect 5889 32395 6489 32419
rect 5889 32339 5905 32395
rect 5961 32339 5991 32395
rect 6047 32339 6077 32395
rect 6133 32339 6163 32395
rect 6219 32339 6249 32395
rect 6305 32339 6335 32395
rect 6391 32339 6421 32395
rect 6477 32339 6489 32395
rect 5889 32315 6489 32339
rect 5889 32259 5905 32315
rect 5961 32259 5991 32315
rect 6047 32259 6077 32315
rect 6133 32259 6163 32315
rect 6219 32259 6249 32315
rect 6305 32259 6335 32315
rect 6391 32259 6421 32315
rect 6477 32259 6489 32315
rect 5889 32235 6489 32259
rect 5889 32179 5905 32235
rect 5961 32179 5991 32235
rect 6047 32179 6077 32235
rect 6133 32179 6163 32235
rect 6219 32179 6249 32235
rect 6305 32179 6335 32235
rect 6391 32179 6421 32235
rect 6477 32179 6489 32235
rect 5889 32155 6489 32179
rect 5889 32099 5905 32155
rect 5961 32099 5991 32155
rect 6047 32099 6077 32155
rect 6133 32099 6163 32155
rect 6219 32099 6249 32155
rect 6305 32099 6335 32155
rect 6391 32099 6421 32155
rect 6477 32099 6489 32155
rect 5889 32075 6489 32099
rect 5889 32019 5905 32075
rect 5961 32019 5991 32075
rect 6047 32019 6077 32075
rect 6133 32019 6163 32075
rect 6219 32019 6249 32075
rect 6305 32019 6335 32075
rect 6391 32019 6421 32075
rect 6477 32019 6489 32075
rect 5889 31995 6489 32019
rect 5889 31939 5905 31995
rect 5961 31939 5991 31995
rect 6047 31939 6077 31995
rect 6133 31939 6163 31995
rect 6219 31939 6249 31995
rect 6305 31939 6335 31995
rect 6391 31939 6421 31995
rect 6477 31939 6489 31995
rect 5889 31915 6489 31939
rect 5889 31859 5905 31915
rect 5961 31859 5991 31915
rect 6047 31859 6077 31915
rect 6133 31859 6163 31915
rect 6219 31859 6249 31915
rect 6305 31859 6335 31915
rect 6391 31859 6421 31915
rect 6477 31859 6489 31915
rect 5889 31835 6489 31859
rect 5889 31779 5905 31835
rect 5961 31779 5991 31835
rect 6047 31779 6077 31835
rect 6133 31779 6163 31835
rect 6219 31779 6249 31835
rect 6305 31779 6335 31835
rect 6391 31779 6421 31835
rect 6477 31779 6489 31835
rect 5889 31755 6489 31779
rect 5889 31699 5905 31755
rect 5961 31699 5991 31755
rect 6047 31699 6077 31755
rect 6133 31699 6163 31755
rect 6219 31699 6249 31755
rect 6305 31699 6335 31755
rect 6391 31699 6421 31755
rect 6477 31699 6489 31755
rect 5889 31675 6489 31699
rect 5889 31619 5905 31675
rect 5961 31619 5991 31675
rect 6047 31619 6077 31675
rect 6133 31619 6163 31675
rect 6219 31619 6249 31675
rect 6305 31619 6335 31675
rect 6391 31619 6421 31675
rect 6477 31619 6489 31675
rect 5889 31595 6489 31619
rect 5889 31539 5905 31595
rect 5961 31539 5991 31595
rect 6047 31539 6077 31595
rect 6133 31539 6163 31595
rect 6219 31539 6249 31595
rect 6305 31539 6335 31595
rect 6391 31539 6421 31595
rect 6477 31539 6489 31595
rect 5889 31515 6489 31539
rect 5889 31459 5905 31515
rect 5961 31459 5991 31515
rect 6047 31459 6077 31515
rect 6133 31459 6163 31515
rect 6219 31459 6249 31515
rect 6305 31459 6335 31515
rect 6391 31459 6421 31515
rect 6477 31459 6489 31515
rect 5889 31435 6489 31459
rect 5889 31379 5905 31435
rect 5961 31379 5991 31435
rect 6047 31379 6077 31435
rect 6133 31379 6163 31435
rect 6219 31379 6249 31435
rect 6305 31379 6335 31435
rect 6391 31379 6421 31435
rect 6477 31379 6489 31435
rect 5889 31355 6489 31379
rect 5889 31299 5905 31355
rect 5961 31299 5991 31355
rect 6047 31299 6077 31355
rect 6133 31299 6163 31355
rect 6219 31299 6249 31355
rect 6305 31299 6335 31355
rect 6391 31299 6421 31355
rect 6477 31299 6489 31355
rect 5889 31275 6489 31299
rect 5889 31219 5905 31275
rect 5961 31219 5991 31275
rect 6047 31219 6077 31275
rect 6133 31219 6163 31275
rect 6219 31219 6249 31275
rect 6305 31219 6335 31275
rect 6391 31219 6421 31275
rect 6477 31219 6489 31275
rect 5889 31195 6489 31219
rect 5889 31139 5905 31195
rect 5961 31139 5991 31195
rect 6047 31139 6077 31195
rect 6133 31139 6163 31195
rect 6219 31139 6249 31195
rect 6305 31139 6335 31195
rect 6391 31139 6421 31195
rect 6477 31139 6489 31195
rect 5889 31115 6489 31139
rect 5889 31059 5905 31115
rect 5961 31059 5991 31115
rect 6047 31059 6077 31115
rect 6133 31059 6163 31115
rect 6219 31059 6249 31115
rect 6305 31059 6335 31115
rect 6391 31059 6421 31115
rect 6477 31059 6489 31115
rect 5889 31035 6489 31059
rect 5889 30979 5905 31035
rect 5961 30979 5991 31035
rect 6047 30979 6077 31035
rect 6133 30979 6163 31035
rect 6219 30979 6249 31035
rect 6305 30979 6335 31035
rect 6391 30979 6421 31035
rect 6477 30979 6489 31035
rect 5889 30955 6489 30979
rect 5889 30899 5905 30955
rect 5961 30899 5991 30955
rect 6047 30899 6077 30955
rect 6133 30899 6163 30955
rect 6219 30899 6249 30955
rect 6305 30899 6335 30955
rect 6391 30899 6421 30955
rect 6477 30899 6489 30955
rect 5889 30875 6489 30899
rect 5889 30819 5905 30875
rect 5961 30819 5991 30875
rect 6047 30819 6077 30875
rect 6133 30819 6163 30875
rect 6219 30819 6249 30875
rect 6305 30819 6335 30875
rect 6391 30819 6421 30875
rect 6477 30819 6489 30875
rect 5889 30795 6489 30819
rect 5889 30739 5905 30795
rect 5961 30739 5991 30795
rect 6047 30739 6077 30795
rect 6133 30739 6163 30795
rect 6219 30739 6249 30795
rect 6305 30739 6335 30795
rect 6391 30739 6421 30795
rect 6477 30739 6489 30795
rect 5889 30715 6489 30739
rect 5889 30659 5905 30715
rect 5961 30659 5991 30715
rect 6047 30659 6077 30715
rect 6133 30659 6163 30715
rect 6219 30659 6249 30715
rect 6305 30659 6335 30715
rect 6391 30659 6421 30715
rect 6477 30659 6489 30715
rect 5889 30635 6489 30659
rect 5889 30579 5905 30635
rect 5961 30579 5991 30635
rect 6047 30579 6077 30635
rect 6133 30579 6163 30635
rect 6219 30579 6249 30635
rect 6305 30579 6335 30635
rect 6391 30579 6421 30635
rect 6477 30579 6489 30635
rect 5889 30555 6489 30579
rect 5889 30499 5905 30555
rect 5961 30499 5991 30555
rect 6047 30499 6077 30555
rect 6133 30499 6163 30555
rect 6219 30499 6249 30555
rect 6305 30499 6335 30555
rect 6391 30499 6421 30555
rect 6477 30499 6489 30555
rect 5889 30475 6489 30499
rect 5889 30419 5905 30475
rect 5961 30419 5991 30475
rect 6047 30419 6077 30475
rect 6133 30419 6163 30475
rect 6219 30419 6249 30475
rect 6305 30419 6335 30475
rect 6391 30419 6421 30475
rect 6477 30419 6489 30475
rect 5889 30395 6489 30419
rect 5889 30339 5905 30395
rect 5961 30339 5991 30395
rect 6047 30339 6077 30395
rect 6133 30339 6163 30395
rect 6219 30339 6249 30395
rect 6305 30339 6335 30395
rect 6391 30339 6421 30395
rect 6477 30339 6489 30395
rect 5889 30315 6489 30339
rect 5889 30259 5905 30315
rect 5961 30259 5991 30315
rect 6047 30259 6077 30315
rect 6133 30259 6163 30315
rect 6219 30259 6249 30315
rect 6305 30259 6335 30315
rect 6391 30259 6421 30315
rect 6477 30259 6489 30315
rect 5889 30235 6489 30259
rect 5889 30179 5905 30235
rect 5961 30179 5991 30235
rect 6047 30179 6077 30235
rect 6133 30179 6163 30235
rect 6219 30179 6249 30235
rect 6305 30179 6335 30235
rect 6391 30179 6421 30235
rect 6477 30179 6489 30235
rect 5889 30155 6489 30179
rect 5889 30099 5905 30155
rect 5961 30099 5991 30155
rect 6047 30099 6077 30155
rect 6133 30099 6163 30155
rect 6219 30099 6249 30155
rect 6305 30099 6335 30155
rect 6391 30099 6421 30155
rect 6477 30099 6489 30155
rect 5889 30075 6489 30099
rect 5889 30019 5905 30075
rect 5961 30019 5991 30075
rect 6047 30019 6077 30075
rect 6133 30019 6163 30075
rect 6219 30019 6249 30075
rect 6305 30019 6335 30075
rect 6391 30019 6421 30075
rect 6477 30019 6489 30075
rect 5889 29890 6489 30019
rect 6589 29956 6655 34990
rect 6890 35094 6903 35150
rect 6959 35094 6993 35150
rect 7049 35094 7083 35150
rect 7139 35094 7173 35150
rect 7229 35094 7263 35150
rect 7319 35094 7353 35150
rect 7409 35094 7443 35150
rect 7499 35094 7528 35150
rect 6890 35070 7528 35094
rect 6890 35014 6903 35070
rect 6959 35014 6993 35070
rect 7049 35014 7083 35070
rect 7139 35014 7173 35070
rect 7229 35014 7263 35070
rect 7319 35014 7353 35070
rect 7409 35014 7443 35070
rect 7499 35014 7528 35070
rect 6890 34990 7528 35014
rect 6890 34934 6903 34990
rect 6959 34934 6993 34990
rect 7049 34934 7083 34990
rect 7139 34934 7173 34990
rect 7229 34934 7263 34990
rect 7319 34934 7353 34990
rect 7409 34934 7443 34990
rect 7499 34934 7528 34990
rect 6890 34910 7528 34934
rect 6890 34854 6903 34910
rect 6959 34854 6993 34910
rect 7049 34854 7083 34910
rect 7139 34854 7173 34910
rect 7229 34854 7263 34910
rect 7319 34854 7353 34910
rect 7409 34854 7443 34910
rect 7499 34854 7528 34910
rect 6890 34830 7528 34854
rect 6890 34774 6903 34830
rect 6959 34774 6993 34830
rect 7049 34774 7083 34830
rect 7139 34774 7173 34830
rect 7229 34774 7263 34830
rect 7319 34774 7353 34830
rect 7409 34774 7443 34830
rect 7499 34774 7528 34830
rect 6890 34750 7528 34774
rect 6890 34694 6903 34750
rect 6959 34694 6993 34750
rect 7049 34694 7083 34750
rect 7139 34694 7173 34750
rect 7229 34694 7263 34750
rect 7319 34694 7353 34750
rect 7409 34694 7443 34750
rect 7499 34694 7528 34750
rect 6890 34670 7528 34694
rect 6890 34614 6903 34670
rect 6959 34614 6993 34670
rect 7049 34614 7083 34670
rect 7139 34614 7173 34670
rect 7229 34614 7263 34670
rect 7319 34614 7353 34670
rect 7409 34614 7443 34670
rect 7499 34614 7528 34670
rect 6890 34590 7528 34614
rect 6890 34534 6903 34590
rect 6959 34534 6993 34590
rect 7049 34534 7083 34590
rect 7139 34534 7173 34590
rect 7229 34534 7263 34590
rect 7319 34534 7353 34590
rect 7409 34534 7443 34590
rect 7499 34534 7528 34590
rect 6890 34510 7528 34534
rect 6890 34454 6903 34510
rect 6959 34454 6993 34510
rect 7049 34454 7083 34510
rect 7139 34454 7173 34510
rect 7229 34454 7263 34510
rect 7319 34454 7353 34510
rect 7409 34454 7443 34510
rect 7499 34454 7528 34510
rect 6890 34430 7528 34454
rect 6890 34374 6903 34430
rect 6959 34374 6993 34430
rect 7049 34374 7083 34430
rect 7139 34374 7173 34430
rect 7229 34374 7263 34430
rect 7319 34374 7353 34430
rect 7409 34374 7443 34430
rect 7499 34374 7528 34430
rect 6890 34350 7528 34374
rect 6890 34294 6903 34350
rect 6959 34294 6993 34350
rect 7049 34294 7083 34350
rect 7139 34294 7173 34350
rect 7229 34294 7263 34350
rect 7319 34294 7353 34350
rect 7409 34294 7443 34350
rect 7499 34294 7528 34350
rect 6890 34270 7528 34294
rect 6890 34214 6903 34270
rect 6959 34214 6993 34270
rect 7049 34214 7083 34270
rect 7139 34214 7173 34270
rect 7229 34214 7263 34270
rect 7319 34214 7353 34270
rect 7409 34214 7443 34270
rect 7499 34214 7528 34270
rect 6890 34190 7528 34214
rect 6890 34134 6903 34190
rect 6959 34134 6993 34190
rect 7049 34134 7083 34190
rect 7139 34134 7173 34190
rect 7229 34134 7263 34190
rect 7319 34134 7353 34190
rect 7409 34134 7443 34190
rect 7499 34134 7528 34190
rect 6890 34110 7528 34134
rect 6890 34054 6903 34110
rect 6959 34054 6993 34110
rect 7049 34054 7083 34110
rect 7139 34054 7173 34110
rect 7229 34054 7263 34110
rect 7319 34054 7353 34110
rect 7409 34054 7443 34110
rect 7499 34054 7528 34110
rect 6890 34030 7528 34054
rect 6890 33974 6903 34030
rect 6959 33974 6993 34030
rect 7049 33974 7083 34030
rect 7139 33974 7173 34030
rect 7229 33974 7263 34030
rect 7319 33974 7353 34030
rect 7409 33974 7443 34030
rect 7499 33974 7528 34030
rect 6890 33950 7528 33974
rect 6890 33894 6903 33950
rect 6959 33894 6993 33950
rect 7049 33894 7083 33950
rect 7139 33894 7173 33950
rect 7229 33894 7263 33950
rect 7319 33894 7353 33950
rect 7409 33894 7443 33950
rect 7499 33894 7528 33950
rect 6890 33870 7528 33894
rect 6890 33814 6903 33870
rect 6959 33814 6993 33870
rect 7049 33814 7083 33870
rect 7139 33814 7173 33870
rect 7229 33814 7263 33870
rect 7319 33814 7353 33870
rect 7409 33814 7443 33870
rect 7499 33814 7528 33870
rect 6890 33790 7528 33814
rect 6890 33734 6903 33790
rect 6959 33734 6993 33790
rect 7049 33734 7083 33790
rect 7139 33734 7173 33790
rect 7229 33734 7263 33790
rect 7319 33734 7353 33790
rect 7409 33734 7443 33790
rect 7499 33734 7528 33790
rect 6890 33710 7528 33734
rect 6890 33654 6903 33710
rect 6959 33654 6993 33710
rect 7049 33654 7083 33710
rect 7139 33654 7173 33710
rect 7229 33654 7263 33710
rect 7319 33654 7353 33710
rect 7409 33654 7443 33710
rect 7499 33654 7528 33710
rect 6890 33630 7528 33654
rect 6890 33574 6903 33630
rect 6959 33574 6993 33630
rect 7049 33574 7083 33630
rect 7139 33574 7173 33630
rect 7229 33574 7263 33630
rect 7319 33574 7353 33630
rect 7409 33574 7443 33630
rect 7499 33574 7528 33630
rect 6890 33550 7528 33574
rect 6890 33494 6903 33550
rect 6959 33494 6993 33550
rect 7049 33494 7083 33550
rect 7139 33494 7173 33550
rect 7229 33494 7263 33550
rect 7319 33494 7353 33550
rect 7409 33494 7443 33550
rect 7499 33494 7528 33550
rect 6890 33470 7528 33494
rect 6890 33414 6903 33470
rect 6959 33414 6993 33470
rect 7049 33414 7083 33470
rect 7139 33414 7173 33470
rect 7229 33414 7263 33470
rect 7319 33414 7353 33470
rect 7409 33414 7443 33470
rect 7499 33414 7528 33470
rect 6890 33390 7528 33414
rect 6890 33334 6903 33390
rect 6959 33334 6993 33390
rect 7049 33334 7083 33390
rect 7139 33334 7173 33390
rect 7229 33334 7263 33390
rect 7319 33334 7353 33390
rect 7409 33334 7443 33390
rect 7499 33334 7528 33390
rect 6890 33310 7528 33334
rect 6890 33254 6903 33310
rect 6959 33254 6993 33310
rect 7049 33254 7083 33310
rect 7139 33254 7173 33310
rect 7229 33254 7263 33310
rect 7319 33254 7353 33310
rect 7409 33254 7443 33310
rect 7499 33254 7528 33310
rect 6890 33230 7528 33254
rect 6890 33174 6903 33230
rect 6959 33174 6993 33230
rect 7049 33174 7083 33230
rect 7139 33174 7173 33230
rect 7229 33174 7263 33230
rect 7319 33174 7353 33230
rect 7409 33174 7443 33230
rect 7499 33174 7528 33230
rect 6890 33150 7528 33174
rect 6890 33094 6903 33150
rect 6959 33094 6993 33150
rect 7049 33094 7083 33150
rect 7139 33094 7173 33150
rect 7229 33094 7263 33150
rect 7319 33094 7353 33150
rect 7409 33094 7443 33150
rect 7499 33094 7528 33150
rect 6890 33070 7528 33094
rect 6890 33014 6903 33070
rect 6959 33014 6993 33070
rect 7049 33014 7083 33070
rect 7139 33014 7173 33070
rect 7229 33014 7263 33070
rect 7319 33014 7353 33070
rect 7409 33014 7443 33070
rect 7499 33014 7528 33070
rect 6890 32990 7528 33014
rect 6890 32934 6903 32990
rect 6959 32934 6993 32990
rect 7049 32934 7083 32990
rect 7139 32934 7173 32990
rect 7229 32934 7263 32990
rect 7319 32934 7353 32990
rect 7409 32934 7443 32990
rect 7499 32934 7528 32990
rect 6890 32910 7528 32934
rect 6890 32854 6903 32910
rect 6959 32854 6993 32910
rect 7049 32854 7083 32910
rect 7139 32854 7173 32910
rect 7229 32854 7263 32910
rect 7319 32854 7353 32910
rect 7409 32854 7443 32910
rect 7499 32854 7528 32910
rect 6890 32830 7528 32854
rect 6890 32774 6903 32830
rect 6959 32774 6993 32830
rect 7049 32774 7083 32830
rect 7139 32774 7173 32830
rect 7229 32774 7263 32830
rect 7319 32774 7353 32830
rect 7409 32774 7443 32830
rect 7499 32774 7528 32830
rect 6890 32750 7528 32774
rect 6890 32694 6903 32750
rect 6959 32694 6993 32750
rect 7049 32694 7083 32750
rect 7139 32694 7173 32750
rect 7229 32694 7263 32750
rect 7319 32694 7353 32750
rect 7409 32694 7443 32750
rect 7499 32694 7528 32750
rect 6890 32670 7528 32694
rect 6890 32614 6903 32670
rect 6959 32614 6993 32670
rect 7049 32614 7083 32670
rect 7139 32614 7173 32670
rect 7229 32614 7263 32670
rect 7319 32614 7353 32670
rect 7409 32614 7443 32670
rect 7499 32614 7528 32670
rect 6890 32590 7528 32614
rect 6890 32534 6903 32590
rect 6959 32534 6993 32590
rect 7049 32534 7083 32590
rect 7139 32534 7173 32590
rect 7229 32534 7263 32590
rect 7319 32534 7353 32590
rect 7409 32534 7443 32590
rect 7499 32534 7528 32590
rect 6890 32510 7528 32534
rect 6890 32454 6903 32510
rect 6959 32454 6993 32510
rect 7049 32454 7083 32510
rect 7139 32454 7173 32510
rect 7229 32454 7263 32510
rect 7319 32454 7353 32510
rect 7409 32454 7443 32510
rect 7499 32454 7528 32510
rect 6890 32430 7528 32454
rect 6890 32374 6903 32430
rect 6959 32374 6993 32430
rect 7049 32374 7083 32430
rect 7139 32374 7173 32430
rect 7229 32374 7263 32430
rect 7319 32374 7353 32430
rect 7409 32374 7443 32430
rect 7499 32374 7528 32430
rect 6890 32350 7528 32374
rect 6890 32294 6903 32350
rect 6959 32294 6993 32350
rect 7049 32294 7083 32350
rect 7139 32294 7173 32350
rect 7229 32294 7263 32350
rect 7319 32294 7353 32350
rect 7409 32294 7443 32350
rect 7499 32294 7528 32350
rect 6890 32270 7528 32294
rect 6890 32214 6903 32270
rect 6959 32214 6993 32270
rect 7049 32214 7083 32270
rect 7139 32214 7173 32270
rect 7229 32214 7263 32270
rect 7319 32214 7353 32270
rect 7409 32214 7443 32270
rect 7499 32214 7528 32270
rect 6890 32190 7528 32214
rect 6890 32134 6903 32190
rect 6959 32134 6993 32190
rect 7049 32134 7083 32190
rect 7139 32134 7173 32190
rect 7229 32134 7263 32190
rect 7319 32134 7353 32190
rect 7409 32134 7443 32190
rect 7499 32134 7528 32190
rect 6890 32110 7528 32134
rect 6890 32054 6903 32110
rect 6959 32054 6993 32110
rect 7049 32054 7083 32110
rect 7139 32054 7173 32110
rect 7229 32054 7263 32110
rect 7319 32054 7353 32110
rect 7409 32054 7443 32110
rect 7499 32054 7528 32110
rect 6890 32030 7528 32054
rect 6890 31974 6903 32030
rect 6959 31974 6993 32030
rect 7049 31974 7083 32030
rect 7139 31974 7173 32030
rect 7229 31974 7263 32030
rect 7319 31974 7353 32030
rect 7409 31974 7443 32030
rect 7499 31974 7528 32030
rect 6890 31950 7528 31974
rect 6890 31894 6903 31950
rect 6959 31894 6993 31950
rect 7049 31894 7083 31950
rect 7139 31894 7173 31950
rect 7229 31894 7263 31950
rect 7319 31894 7353 31950
rect 7409 31894 7443 31950
rect 7499 31894 7528 31950
rect 6890 31870 7528 31894
rect 6890 31814 6903 31870
rect 6959 31814 6993 31870
rect 7049 31814 7083 31870
rect 7139 31814 7173 31870
rect 7229 31814 7263 31870
rect 7319 31814 7353 31870
rect 7409 31814 7443 31870
rect 7499 31814 7528 31870
rect 6890 31790 7528 31814
rect 6890 31734 6903 31790
rect 6959 31734 6993 31790
rect 7049 31734 7083 31790
rect 7139 31734 7173 31790
rect 7229 31734 7263 31790
rect 7319 31734 7353 31790
rect 7409 31734 7443 31790
rect 7499 31734 7528 31790
rect 6890 31710 7528 31734
rect 6890 31654 6903 31710
rect 6959 31654 6993 31710
rect 7049 31654 7083 31710
rect 7139 31654 7173 31710
rect 7229 31654 7263 31710
rect 7319 31654 7353 31710
rect 7409 31654 7443 31710
rect 7499 31654 7528 31710
rect 6890 31630 7528 31654
rect 6890 31574 6903 31630
rect 6959 31574 6993 31630
rect 7049 31574 7083 31630
rect 7139 31574 7173 31630
rect 7229 31574 7263 31630
rect 7319 31574 7353 31630
rect 7409 31574 7443 31630
rect 7499 31574 7528 31630
rect 6890 31550 7528 31574
rect 6890 31494 6903 31550
rect 6959 31494 6993 31550
rect 7049 31494 7083 31550
rect 7139 31494 7173 31550
rect 7229 31494 7263 31550
rect 7319 31494 7353 31550
rect 7409 31494 7443 31550
rect 7499 31494 7528 31550
rect 6890 31470 7528 31494
rect 6890 31414 6903 31470
rect 6959 31414 6993 31470
rect 7049 31414 7083 31470
rect 7139 31414 7173 31470
rect 7229 31414 7263 31470
rect 7319 31414 7353 31470
rect 7409 31414 7443 31470
rect 7499 31414 7528 31470
rect 6890 31390 7528 31414
rect 6890 31334 6903 31390
rect 6959 31334 6993 31390
rect 7049 31334 7083 31390
rect 7139 31334 7173 31390
rect 7229 31334 7263 31390
rect 7319 31334 7353 31390
rect 7409 31334 7443 31390
rect 7499 31334 7528 31390
rect 6890 31310 7528 31334
rect 6890 31254 6903 31310
rect 6959 31254 6993 31310
rect 7049 31254 7083 31310
rect 7139 31254 7173 31310
rect 7229 31254 7263 31310
rect 7319 31254 7353 31310
rect 7409 31254 7443 31310
rect 7499 31254 7528 31310
rect 6890 31230 7528 31254
rect 6890 31174 6903 31230
rect 6959 31174 6993 31230
rect 7049 31174 7083 31230
rect 7139 31174 7173 31230
rect 7229 31174 7263 31230
rect 7319 31174 7353 31230
rect 7409 31174 7443 31230
rect 7499 31174 7528 31230
rect 6890 31150 7528 31174
rect 6890 31094 6903 31150
rect 6959 31094 6993 31150
rect 7049 31094 7083 31150
rect 7139 31094 7173 31150
rect 7229 31094 7263 31150
rect 7319 31094 7353 31150
rect 7409 31094 7443 31150
rect 7499 31094 7528 31150
rect 6890 31070 7528 31094
rect 6890 31014 6903 31070
rect 6959 31014 6993 31070
rect 7049 31014 7083 31070
rect 7139 31014 7173 31070
rect 7229 31014 7263 31070
rect 7319 31014 7353 31070
rect 7409 31014 7443 31070
rect 7499 31014 7528 31070
rect 6890 30990 7528 31014
rect 6890 30934 6903 30990
rect 6959 30934 6993 30990
rect 7049 30934 7083 30990
rect 7139 30934 7173 30990
rect 7229 30934 7263 30990
rect 7319 30934 7353 30990
rect 7409 30934 7443 30990
rect 7499 30934 7528 30990
rect 6890 30910 7528 30934
rect 6890 30854 6903 30910
rect 6959 30854 6993 30910
rect 7049 30854 7083 30910
rect 7139 30854 7173 30910
rect 7229 30854 7263 30910
rect 7319 30854 7353 30910
rect 7409 30854 7443 30910
rect 7499 30854 7528 30910
rect 6890 30830 7528 30854
rect 6890 30774 6903 30830
rect 6959 30774 6993 30830
rect 7049 30774 7083 30830
rect 7139 30774 7173 30830
rect 7229 30774 7263 30830
rect 7319 30774 7353 30830
rect 7409 30774 7443 30830
rect 7499 30774 7528 30830
rect 6890 30750 7528 30774
rect 6890 30694 6903 30750
rect 6959 30694 6993 30750
rect 7049 30694 7083 30750
rect 7139 30694 7173 30750
rect 7229 30694 7263 30750
rect 7319 30694 7353 30750
rect 7409 30694 7443 30750
rect 7499 30694 7528 30750
rect 6890 30670 7528 30694
rect 6890 30614 6903 30670
rect 6959 30614 6993 30670
rect 7049 30614 7083 30670
rect 7139 30614 7173 30670
rect 7229 30614 7263 30670
rect 7319 30614 7353 30670
rect 7409 30614 7443 30670
rect 7499 30614 7528 30670
rect 6890 30590 7528 30614
rect 6890 30534 6903 30590
rect 6959 30534 6993 30590
rect 7049 30534 7083 30590
rect 7139 30534 7173 30590
rect 7229 30534 7263 30590
rect 7319 30534 7353 30590
rect 7409 30534 7443 30590
rect 7499 30534 7528 30590
rect 6890 30510 7528 30534
rect 6890 30454 6903 30510
rect 6959 30454 6993 30510
rect 7049 30454 7083 30510
rect 7139 30454 7173 30510
rect 7229 30454 7263 30510
rect 7319 30454 7353 30510
rect 7409 30454 7443 30510
rect 7499 30454 7528 30510
rect 6890 30430 7528 30454
rect 6890 30374 6903 30430
rect 6959 30374 6993 30430
rect 7049 30374 7083 30430
rect 7139 30374 7173 30430
rect 7229 30374 7263 30430
rect 7319 30374 7353 30430
rect 7409 30374 7443 30430
rect 7499 30374 7528 30430
rect 6890 30350 7528 30374
rect 6890 30294 6903 30350
rect 6959 30294 6993 30350
rect 7049 30294 7083 30350
rect 7139 30294 7173 30350
rect 7229 30294 7263 30350
rect 7319 30294 7353 30350
rect 7409 30294 7443 30350
rect 7499 30294 7528 30350
rect 6890 30270 7528 30294
rect 6890 30214 6903 30270
rect 6959 30214 6993 30270
rect 7049 30214 7083 30270
rect 7139 30214 7173 30270
rect 7229 30214 7263 30270
rect 7319 30214 7353 30270
rect 7409 30214 7443 30270
rect 7499 30214 7528 30270
rect 6890 30189 7528 30214
rect 6890 30133 6903 30189
rect 6959 30133 6993 30189
rect 7049 30133 7083 30189
rect 7139 30133 7173 30189
rect 7229 30133 7263 30189
rect 7319 30133 7353 30189
rect 7409 30133 7443 30189
rect 7499 30133 7528 30189
rect 6890 30108 7528 30133
rect 6890 30052 6903 30108
rect 6959 30052 6993 30108
rect 7049 30052 7083 30108
rect 7139 30052 7173 30108
rect 7229 30052 7263 30108
rect 7319 30052 7353 30108
rect 7409 30052 7443 30108
rect 7499 30053 7528 30108
tri 7528 30053 7584 30109 sw
rect 7499 30052 7584 30053
rect 6890 30043 7584 30052
tri 7584 30043 7594 30053 sw
rect 6890 29984 7594 30043
tri 7594 29984 7653 30043 sw
tri 6589 29939 6606 29956 ne
rect 6606 29939 6655 29956
tri 6655 29939 6700 29984 sw
rect 6890 29939 7653 29984
tri 7653 29939 7698 29984 sw
tri 6606 29909 6636 29939 ne
rect 6636 29909 6700 29939
tri 6700 29909 6730 29939 sw
rect 6890 29909 7698 29939
tri 7698 29909 7728 29939 sw
tri 6489 29890 6508 29909 sw
tri 6636 29890 6655 29909 ne
rect 6655 29890 6730 29909
rect 5889 29845 6508 29890
tri 6508 29845 6553 29890 sw
tri 6655 29845 6700 29890 ne
rect 6700 29845 6730 29890
tri 6730 29845 6794 29909 sw
rect 6890 29897 7728 29909
tri 6890 29845 6942 29897 ne
rect 6942 29845 7728 29897
tri 7728 29845 7792 29909 sw
rect 5889 29827 6553 29845
tri 6553 29827 6571 29845 sw
tri 6700 29827 6718 29845 ne
rect 6718 29827 6794 29845
rect 5889 29751 6571 29827
tri 6571 29751 6647 29827 sw
tri 6718 29751 6794 29827 ne
tri 6794 29751 6888 29845 sw
tri 6942 29751 7036 29845 ne
rect 7036 29751 7792 29845
tri 7792 29751 7886 29845 sw
rect 5889 29680 6647 29751
tri 6647 29680 6718 29751 sw
tri 6794 29680 6865 29751 ne
rect 6865 29749 6888 29751
tri 6888 29749 6890 29751 sw
tri 7036 29749 7038 29751 ne
rect 7038 29749 7886 29751
rect 6865 29680 6890 29749
tri 6890 29680 6959 29749 sw
tri 7038 29680 7107 29749 ne
rect 7107 29680 7886 29749
tri 7886 29680 7957 29751 sw
rect 5889 29659 6718 29680
tri 5889 29612 5936 29659 ne
rect 5936 29657 6718 29659
tri 6718 29657 6741 29680 sw
tri 6865 29657 6888 29680 ne
rect 6888 29657 6959 29680
tri 6959 29657 6982 29680 sw
tri 7107 29657 7130 29680 ne
rect 7130 29657 7957 29680
tri 7957 29657 7980 29680 sw
rect 5936 29612 6741 29657
tri 6741 29612 6786 29657 sw
tri 6888 29655 6890 29657 ne
rect 6890 29655 6982 29657
tri 6890 29612 6933 29655 ne
rect 6933 29612 6982 29655
tri 5723 29567 5740 29584 ne
rect 5740 29567 5789 29584
tri 5789 29567 5834 29612 sw
tri 5936 29567 5981 29612 ne
rect 5981 29567 6786 29612
tri 6786 29567 6831 29612 sw
tri 6933 29567 6978 29612 ne
rect 6978 29567 6982 29612
tri 5740 29518 5789 29567 ne
rect 5789 29563 5834 29567
tri 5834 29563 5838 29567 sw
tri 5981 29563 5985 29567 ne
rect 5985 29563 6831 29567
tri 6831 29563 6835 29567 sw
tri 6978 29563 6982 29567 ne
tri 6982 29563 7076 29657 sw
tri 7130 29563 7224 29657 ne
rect 7224 29563 7980 29657
tri 7980 29563 8074 29657 sw
rect 5789 29518 5838 29563
tri 5838 29518 5883 29563 sw
tri 5985 29518 6030 29563 ne
rect 6030 29518 6835 29563
tri 6835 29518 6880 29563 sw
tri 6982 29518 7027 29563 ne
rect 7027 29518 7076 29563
tri 7076 29518 7121 29563 sw
tri 7224 29518 7269 29563 ne
rect 7269 29518 8074 29563
tri 8074 29518 8119 29563 sw
tri 2501 29510 2509 29518 se
rect 2509 29512 3353 29518
tri 3353 29512 3359 29518 nw
tri 3500 29512 3506 29518 se
rect 2509 29510 3351 29512
tri 3351 29510 3353 29512 nw
tri 3498 29510 3500 29512 se
rect 3500 29510 3506 29512
tri 1167 29416 1261 29510 se
rect 1261 29416 2017 29510
tri 2017 29416 2111 29510 nw
tri 2170 29416 2264 29510 se
tri 2264 29416 2358 29510 nw
tri 2415 29424 2501 29510 se
rect 2501 29424 3265 29510
tri 3265 29424 3351 29510 nw
tri 3412 29424 3498 29510 se
rect 3498 29424 3506 29510
tri 3506 29424 3600 29518 nw
tri 5789 29473 5834 29518 ne
rect 5834 29512 5883 29518
tri 5883 29512 5889 29518 sw
tri 6030 29512 6036 29518 ne
rect 6036 29512 6880 29518
rect 5834 29473 5889 29512
tri 5889 29473 5928 29512 sw
tri 6036 29473 6075 29512 ne
rect 6075 29508 6880 29512
tri 6880 29508 6890 29518 sw
tri 7027 29508 7037 29518 ne
rect 7037 29508 7121 29518
rect 6075 29473 6890 29508
tri 6890 29473 6925 29508 sw
tri 7037 29473 7072 29508 ne
rect 7072 29473 7121 29508
tri 5834 29424 5883 29473 ne
rect 5883 29469 5928 29473
tri 5928 29469 5932 29473 sw
tri 6075 29469 6079 29473 ne
rect 6079 29469 6925 29473
tri 6925 29469 6929 29473 sw
tri 7072 29469 7076 29473 ne
rect 7076 29469 7121 29473
tri 7121 29469 7170 29518 sw
tri 7269 29469 7318 29518 ne
rect 7318 29469 8119 29518
tri 8119 29469 8168 29518 sw
rect 5883 29424 5932 29469
tri 5932 29424 5977 29469 sw
tri 6079 29424 6124 29469 ne
rect 6124 29424 6929 29469
tri 6929 29424 6974 29469 sw
tri 7076 29424 7121 29469 ne
rect 7121 29424 7170 29469
tri 7170 29424 7215 29469 sw
tri 7318 29424 7363 29469 ne
rect 7363 29424 8168 29469
tri 8168 29424 8213 29469 sw
tri 2407 29416 2415 29424 se
rect 2415 29416 3257 29424
tri 3257 29416 3265 29424 nw
tri 3404 29416 3412 29424 se
rect 3412 29418 3500 29424
tri 3500 29418 3506 29424 nw
tri 5883 29418 5889 29424 ne
rect 5889 29418 5977 29424
tri 1073 29322 1167 29416 se
rect 1167 29322 1923 29416
tri 1923 29322 2017 29416 nw
tri 2076 29322 2170 29416 se
tri 2170 29322 2264 29416 nw
tri 2321 29330 2407 29416 se
rect 2407 29330 3171 29416
tri 3171 29330 3257 29416 nw
tri 3318 29330 3404 29416 se
rect 3404 29330 3412 29416
tri 3412 29330 3500 29418 nw
tri 5889 29379 5928 29418 ne
rect 5928 29379 5977 29418
tri 5977 29379 6022 29424 sw
tri 6124 29379 6169 29424 ne
rect 6169 29379 6974 29424
tri 6974 29379 7019 29424 sw
tri 7121 29379 7166 29424 ne
rect 7166 29379 7215 29424
tri 5928 29330 5977 29379 ne
rect 5977 29375 6022 29379
tri 6022 29375 6026 29379 sw
tri 6169 29375 6173 29379 ne
rect 6173 29375 7019 29379
tri 7019 29375 7023 29379 sw
tri 7166 29375 7170 29379 ne
rect 7170 29375 7215 29379
tri 7215 29375 7264 29424 sw
tri 7363 29375 7412 29424 ne
rect 7412 29375 8213 29424
tri 8213 29375 8262 29424 sw
rect 5977 29330 6026 29375
tri 6026 29330 6071 29375 sw
tri 6173 29330 6218 29375 ne
rect 6218 29330 7023 29375
tri 7023 29330 7068 29375 sw
tri 7170 29330 7215 29375 ne
rect 7215 29330 7264 29375
tri 7264 29330 7309 29375 sw
tri 7412 29330 7457 29375 ne
rect 7457 29330 8262 29375
tri 8262 29330 8307 29375 sw
tri 2313 29322 2321 29330 se
rect 2321 29322 3163 29330
tri 3163 29322 3171 29330 nw
tri 3310 29322 3318 29330 se
tri 979 29228 1073 29322 se
rect 1073 29228 1829 29322
tri 1829 29228 1923 29322 nw
tri 1982 29228 2076 29322 se
tri 2076 29228 2170 29322 nw
tri 2227 29236 2313 29322 se
rect 2313 29236 3077 29322
tri 3077 29236 3163 29322 nw
tri 3224 29236 3310 29322 se
rect 3310 29236 3318 29322
tri 3318 29236 3412 29330 nw
tri 5977 29285 6022 29330 ne
rect 6022 29285 6071 29330
tri 6071 29285 6116 29330 sw
tri 6218 29285 6263 29330 ne
rect 6263 29285 7068 29330
tri 7068 29285 7113 29330 sw
tri 7215 29285 7260 29330 ne
rect 7260 29285 7309 29330
tri 6022 29236 6071 29285 ne
rect 6071 29281 6116 29285
tri 6116 29281 6120 29285 sw
tri 6263 29281 6267 29285 ne
rect 6267 29281 7113 29285
tri 7113 29281 7117 29285 sw
tri 7260 29281 7264 29285 ne
rect 7264 29281 7309 29285
tri 7309 29281 7358 29330 sw
tri 7457 29281 7506 29330 ne
rect 7506 29281 8307 29330
tri 8307 29281 8356 29330 sw
rect 6071 29236 6120 29281
tri 6120 29236 6165 29281 sw
tri 6267 29236 6312 29281 ne
rect 6312 29236 7117 29281
tri 7117 29236 7162 29281 sw
tri 7264 29236 7309 29281 ne
rect 7309 29236 7358 29281
tri 7358 29236 7403 29281 sw
tri 7506 29236 7551 29281 ne
rect 7551 29236 8356 29281
tri 8356 29236 8401 29281 sw
tri 2219 29228 2227 29236 se
rect 2227 29228 3069 29236
tri 3069 29228 3077 29236 nw
tri 3216 29228 3224 29236 se
tri 954 29203 979 29228 se
rect 979 29203 1804 29228
tri 1804 29203 1829 29228 nw
tri 1957 29203 1982 29228 se
rect 1982 29203 2051 29228
tri 2051 29203 2076 29228 nw
tri 2194 29203 2219 29228 se
rect 2219 29203 2983 29228
rect 954 29134 1735 29203
tri 1735 29134 1804 29203 nw
tri 1888 29134 1957 29203 se
rect 1957 29134 1982 29203
tri 1982 29134 2051 29203 nw
tri 2133 29142 2194 29203 se
rect 2194 29142 2983 29203
tri 2983 29142 3069 29228 nw
tri 3130 29142 3216 29228 se
rect 3216 29142 3224 29228
tri 3224 29142 3318 29236 nw
tri 6071 29191 6116 29236 ne
rect 6116 29191 6165 29236
tri 6165 29191 6210 29236 sw
tri 6312 29191 6357 29236 ne
rect 6357 29203 7162 29236
tri 7162 29203 7195 29236 sw
tri 7309 29203 7342 29236 ne
rect 7342 29203 7403 29236
tri 7403 29203 7436 29236 sw
tri 7551 29203 7584 29236 ne
rect 7584 29203 8401 29236
tri 8401 29203 8434 29236 sw
rect 6357 29191 7195 29203
tri 7195 29191 7207 29203 sw
tri 7342 29191 7354 29203 ne
rect 7354 29191 7436 29203
tri 6116 29142 6165 29191 ne
rect 6165 29187 6210 29191
tri 6210 29187 6214 29191 sw
tri 6357 29187 6361 29191 ne
rect 6361 29187 7207 29191
tri 7207 29187 7211 29191 sw
tri 7354 29187 7358 29191 ne
rect 7358 29187 7436 29191
tri 7436 29187 7452 29203 sw
tri 7584 29187 7600 29203 ne
rect 7600 29187 8434 29203
rect 6165 29142 6214 29187
tri 6214 29142 6259 29187 sw
tri 6361 29142 6406 29187 ne
rect 6406 29142 7211 29187
tri 7211 29142 7256 29187 sw
tri 7358 29142 7403 29187 ne
rect 7403 29142 7452 29187
tri 7452 29142 7497 29187 sw
tri 7600 29142 7645 29187 ne
rect 7645 29142 8434 29187
tri 2125 29134 2133 29142 se
rect 2133 29134 2975 29142
tri 2975 29134 2983 29142 nw
tri 3122 29134 3130 29142 se
rect 954 29067 1668 29134
tri 1668 29067 1735 29134 nw
tri 1821 29067 1888 29134 se
rect 954 29050 1651 29067
tri 1651 29050 1668 29067 nw
tri 1804 29050 1821 29067 se
rect 1821 29050 1888 29067
rect 954 29040 1641 29050
tri 1641 29040 1651 29050 nw
tri 1794 29040 1804 29050 se
rect 1804 29040 1888 29050
tri 1888 29040 1982 29134 nw
tri 2039 29048 2125 29134 se
rect 2125 29048 2889 29134
tri 2889 29048 2975 29134 nw
tri 3036 29048 3122 29134 se
rect 3122 29048 3130 29134
tri 3130 29048 3224 29142 nw
tri 6165 29097 6210 29142 ne
rect 6210 29097 6259 29142
tri 6259 29097 6304 29142 sw
tri 6406 29097 6451 29142 ne
rect 6451 29097 7256 29142
tri 7256 29097 7301 29142 sw
tri 7403 29097 7448 29142 ne
rect 7448 29097 7497 29142
tri 6210 29048 6259 29097 ne
rect 6259 29093 6304 29097
tri 6304 29093 6308 29097 sw
tri 6451 29093 6455 29097 ne
rect 6455 29093 7301 29097
tri 7301 29093 7305 29097 sw
tri 7448 29093 7452 29097 ne
rect 7452 29093 7497 29097
tri 7497 29093 7546 29142 sw
tri 7645 29093 7694 29142 ne
rect 7694 29093 8434 29142
rect 6259 29048 6308 29093
tri 6308 29048 6353 29093 sw
tri 6455 29048 6500 29093 ne
rect 6500 29048 7305 29093
tri 7305 29048 7350 29093 sw
tri 7452 29048 7497 29093 ne
rect 7497 29071 7546 29093
tri 7546 29071 7568 29093 sw
tri 7694 29071 7716 29093 ne
rect 7716 29071 8434 29093
rect 7497 29055 7568 29071
tri 7568 29055 7584 29071 sw
tri 7716 29055 7732 29071 ne
rect 7732 29055 8434 29071
rect 7497 29048 7584 29055
tri 7584 29048 7591 29055 sw
tri 7732 29048 7739 29055 ne
rect 7739 29048 8434 29055
tri 2031 29040 2039 29048 se
rect 2039 29040 2881 29048
tri 2881 29040 2889 29048 nw
tri 3028 29040 3036 29048 se
rect 954 14684 1554 29040
tri 1554 28953 1641 29040 nw
tri 1707 28953 1794 29040 se
rect 1794 28973 1821 29040
tri 1821 28973 1888 29040 nw
tri 1964 28973 2031 29040 se
rect 2031 28973 2795 29040
rect 1794 28956 1804 28973
tri 1804 28956 1821 28973 nw
tri 1947 28956 1964 28973 se
rect 1964 28956 2795 28973
rect 1794 28953 1801 28956
tri 1801 28953 1804 28956 nw
tri 1945 28954 1947 28956 se
rect 1947 28954 2795 28956
tri 2795 28954 2881 29040 nw
tri 2942 28954 3028 29040 se
rect 3028 28954 3036 29040
tri 3036 28954 3130 29048 nw
tri 6259 29003 6304 29048 ne
rect 6304 29003 6353 29048
tri 6353 29003 6398 29048 sw
tri 6500 29003 6545 29048 ne
rect 6545 29003 7350 29048
tri 7350 29003 7395 29048 sw
tri 7497 29003 7542 29048 ne
rect 7542 29003 7591 29048
tri 6304 28954 6353 29003 ne
rect 6353 28999 6398 29003
tri 6398 28999 6402 29003 sw
tri 6545 28999 6549 29003 ne
rect 6549 28999 7395 29003
tri 7395 28999 7399 29003 sw
tri 7542 28999 7546 29003 ne
rect 7546 28999 7591 29003
tri 7591 28999 7640 29048 sw
tri 7739 28999 7788 29048 ne
rect 7788 28999 8434 29048
rect 6353 28954 6402 28999
tri 6402 28954 6447 28999 sw
tri 6549 28954 6594 28999 ne
rect 6594 28977 7399 28999
tri 7399 28977 7421 28999 sw
tri 7546 28977 7568 28999 ne
rect 7568 28977 7640 28999
rect 6594 28954 7421 28977
tri 7421 28954 7444 28977 sw
tri 7568 28961 7584 28977 ne
rect 7584 28961 7640 28977
tri 7584 28954 7591 28961 ne
rect 7591 28954 7640 28961
tri 7640 28954 7685 28999 sw
tri 7788 28954 7833 28999 ne
rect 7833 28954 8434 28999
tri 1944 28953 1945 28954 se
rect 1945 28953 2787 28954
tri 1700 28946 1707 28953 se
rect 1707 28946 1794 28953
tri 1794 28946 1801 28953 nw
tri 1937 28946 1944 28953 se
rect 1944 28946 2787 28953
tri 2787 28946 2795 28954 nw
tri 2934 28946 2942 28954 se
rect 954 14628 963 14684
rect 1019 14628 1069 14684
rect 1125 14628 1174 14684
rect 1230 14628 1279 14684
rect 1335 14628 1384 14684
rect 1440 14628 1489 14684
rect 1545 14628 1554 14684
rect 954 14540 1554 14628
rect 954 14484 963 14540
rect 1019 14484 1069 14540
rect 1125 14484 1174 14540
rect 1230 14484 1279 14540
rect 1335 14484 1384 14540
rect 1440 14484 1489 14540
rect 1545 14484 1554 14540
rect 453 13795 853 13800
rect 453 13739 462 13795
rect 518 13739 571 13795
rect 627 13739 680 13795
rect 736 13739 788 13795
rect 844 13739 853 13795
rect 453 13651 853 13739
rect 453 13595 462 13651
rect 518 13595 571 13651
rect 627 13595 680 13651
rect 736 13595 788 13651
rect 844 13595 853 13651
rect 315 9241 381 9247
rect 315 9177 316 9241
rect 380 9177 381 9241
rect 315 9156 381 9177
rect 315 9092 316 9156
rect 380 9092 381 9156
rect 315 9071 381 9092
rect 315 9007 316 9071
rect 380 9007 381 9071
rect 315 8986 381 9007
rect 315 8922 316 8986
rect 380 8922 381 8986
rect 315 8901 381 8922
rect 315 8837 316 8901
rect 380 8837 381 8901
rect 315 8816 381 8837
rect 315 8752 316 8816
rect 380 8752 381 8816
rect 315 8731 381 8752
rect 315 8667 316 8731
rect 380 8667 381 8731
rect 315 8645 381 8667
rect 315 8581 316 8645
rect 380 8581 381 8645
rect 315 8559 381 8581
rect 315 8495 316 8559
rect 380 8495 381 8559
rect 315 8473 381 8495
rect 315 8409 316 8473
rect 380 8409 381 8473
rect 315 8387 381 8409
rect 315 8323 316 8387
rect 380 8323 381 8387
rect 315 8317 381 8323
rect 453 8716 853 13595
rect 453 8660 476 8716
rect 532 8660 580 8716
rect 636 8660 684 8716
rect 740 8660 788 8716
rect 844 8660 853 8716
rect 453 8572 853 8660
rect 453 8516 476 8572
rect 532 8516 580 8572
rect 636 8516 684 8572
rect 740 8516 788 8572
rect 844 8516 853 8572
rect 453 7041 853 8516
rect 453 6977 490 7041
rect 554 6977 580 7041
rect 644 6977 670 7041
rect 734 6977 760 7041
rect 824 6977 853 7041
rect 453 6960 853 6977
rect 453 6896 490 6960
rect 554 6896 580 6960
rect 644 6896 670 6960
rect 734 6896 760 6960
rect 824 6896 853 6960
rect 453 6878 853 6896
rect 453 6814 490 6878
rect 554 6814 580 6878
rect 644 6814 670 6878
rect 734 6814 760 6878
rect 824 6814 853 6878
rect 453 6796 853 6814
rect 453 6732 490 6796
rect 554 6732 580 6796
rect 644 6732 670 6796
rect 734 6732 760 6796
rect 824 6732 853 6796
rect 453 6714 853 6732
rect 453 6650 490 6714
rect 554 6650 580 6714
rect 644 6650 670 6714
rect 734 6650 760 6714
rect 824 6650 853 6714
rect 453 6632 853 6650
rect 453 6568 490 6632
rect 554 6568 580 6632
rect 644 6568 670 6632
rect 734 6568 760 6632
rect 824 6568 853 6632
rect 453 6550 853 6568
rect 453 6486 490 6550
rect 554 6486 580 6550
rect 644 6486 670 6550
rect 734 6486 760 6550
rect 824 6486 853 6550
rect 453 6468 853 6486
rect 453 6404 490 6468
rect 554 6404 580 6468
rect 644 6404 670 6468
rect 734 6404 760 6468
rect 824 6404 853 6468
rect 453 6377 853 6404
rect 954 12858 1554 14484
rect 954 12802 963 12858
rect 1019 12802 1069 12858
rect 1125 12802 1174 12858
rect 1230 12802 1279 12858
rect 1335 12802 1384 12858
rect 1440 12802 1489 12858
rect 1545 12802 1554 12858
rect 954 12714 1554 12802
rect 954 12658 963 12714
rect 1019 12658 1069 12714
rect 1125 12658 1174 12714
rect 1230 12658 1279 12714
rect 1335 12658 1384 12714
rect 1440 12658 1489 12714
rect 1545 12658 1554 12714
rect 954 9636 1554 12658
rect 954 9580 963 9636
rect 1019 9580 1069 9636
rect 1125 9580 1174 9636
rect 1230 9580 1279 9636
rect 1335 9580 1384 9636
rect 1440 9580 1489 9636
rect 1545 9580 1554 9636
rect 954 9492 1554 9580
tri 1655 28901 1700 28946 se
rect 1700 28901 1749 28946
tri 1749 28901 1794 28946 nw
tri 1892 28901 1937 28946 se
rect 1937 28901 2742 28946
tri 2742 28901 2787 28946 nw
tri 2889 28901 2934 28946 se
rect 2934 28901 2942 28946
rect 1655 17767 1721 28901
tri 1721 28873 1749 28901 nw
tri 1864 28873 1892 28901 se
rect 1892 28873 2714 28901
tri 2714 28873 2742 28901 nw
tri 2861 28873 2889 28901 se
rect 2889 28873 2942 28901
tri 1851 28860 1864 28873 se
rect 1864 28860 2701 28873
tri 2701 28860 2714 28873 nw
tri 2848 28860 2861 28873 se
rect 2861 28860 2942 28873
tri 2942 28860 3036 28954 nw
tri 6353 28909 6398 28954 ne
rect 6398 28909 6447 28954
tri 6447 28909 6492 28954 sw
tri 6594 28909 6639 28954 ne
rect 6639 28909 7444 28954
tri 7444 28909 7489 28954 sw
tri 7591 28953 7592 28954 ne
rect 7592 28953 7685 28954
tri 7685 28953 7686 28954 sw
tri 7833 28953 7834 28954 ne
tri 7592 28909 7636 28953 ne
rect 7636 28909 7686 28953
tri 6398 28860 6447 28909 ne
rect 6447 28905 6492 28909
tri 6492 28905 6496 28909 sw
tri 6639 28905 6643 28909 ne
rect 6643 28905 7489 28909
tri 7489 28905 7493 28909 sw
tri 7636 28905 7640 28909 ne
rect 7640 28905 7686 28909
tri 7686 28905 7734 28953 sw
rect 6447 28877 6496 28905
tri 6496 28877 6524 28905 sw
tri 6643 28877 6671 28905 ne
rect 6671 28877 7493 28905
tri 7493 28877 7521 28905 sw
tri 7640 28877 7668 28905 ne
rect 6447 28860 6524 28877
tri 6524 28860 6541 28877 sw
tri 6671 28860 6688 28877 ne
rect 6688 28860 7521 28877
tri 7521 28860 7538 28877 sw
rect 1655 17711 1660 17767
rect 1716 17711 1721 17767
rect 1655 17680 1721 17711
rect 1655 17624 1660 17680
rect 1716 17624 1721 17680
rect 1655 17593 1721 17624
rect 1655 17537 1660 17593
rect 1716 17537 1721 17593
rect 1655 17505 1721 17537
rect 1655 17449 1660 17505
rect 1716 17449 1721 17505
rect 1655 17417 1721 17449
rect 1655 17361 1660 17417
rect 1716 17361 1721 17417
rect 1655 17329 1721 17361
rect 1655 17273 1660 17329
rect 1716 17273 1721 17329
rect 1655 17241 1721 17273
rect 1655 17185 1660 17241
rect 1716 17185 1721 17241
rect 1655 9547 1721 17185
tri 1821 28830 1851 28860 se
rect 1851 28830 2671 28860
tri 2671 28830 2701 28860 nw
tri 2818 28830 2848 28860 se
rect 2848 28830 2912 28860
tri 2912 28830 2942 28860 nw
tri 6447 28830 6477 28860 ne
rect 6477 28830 6541 28860
tri 6541 28830 6571 28860 sw
tri 6688 28830 6718 28860 ne
rect 6718 28830 7538 28860
tri 7538 28830 7568 28860 sw
rect 1821 28766 2607 28830
tri 2607 28766 2671 28830 nw
tri 2754 28766 2818 28830 se
rect 2818 28766 2848 28830
tri 2848 28766 2912 28830 nw
tri 6477 28815 6492 28830 ne
rect 6492 28815 6571 28830
tri 6571 28815 6586 28830 sw
tri 6718 28815 6733 28830 ne
rect 6733 28815 7568 28830
tri 6492 28766 6541 28815 ne
rect 6541 28766 6586 28815
tri 6586 28766 6635 28815 sw
tri 6733 28766 6782 28815 ne
rect 6782 28766 7568 28815
rect 1821 28683 2524 28766
tri 2524 28683 2607 28766 nw
tri 2671 28683 2754 28766 se
rect 1821 28672 2513 28683
tri 2513 28672 2524 28683 nw
tri 2660 28672 2671 28683 se
rect 2671 28672 2754 28683
tri 2754 28672 2848 28766 nw
tri 6541 28721 6586 28766 ne
rect 6586 28721 6635 28766
tri 6635 28721 6680 28766 sw
tri 6782 28721 6827 28766 ne
rect 6827 28721 7568 28766
tri 6586 28672 6635 28721 ne
rect 6635 28683 6680 28721
tri 6680 28683 6718 28721 sw
tri 6827 28683 6865 28721 ne
rect 6865 28683 7568 28721
rect 6635 28672 6718 28683
tri 6718 28672 6729 28683 sw
tri 6865 28672 6876 28683 ne
rect 6876 28672 7568 28683
rect 1821 11192 2421 28672
tri 2421 28580 2513 28672 nw
tri 2568 28580 2660 28672 se
rect 2660 28589 2671 28672
tri 2671 28589 2754 28672 nw
tri 6635 28627 6680 28672 ne
rect 6680 28627 6729 28672
tri 6729 28627 6774 28672 sw
tri 6876 28627 6921 28672 ne
rect 6921 28627 7568 28672
tri 6680 28589 6718 28627 ne
rect 6718 28589 6774 28627
rect 2660 28580 2662 28589
tri 2662 28580 2671 28589 nw
tri 6718 28580 6727 28589 ne
rect 6727 28580 6774 28589
tri 6774 28580 6821 28627 sw
tri 6921 28580 6968 28627 ne
tri 2566 28578 2568 28580 se
rect 2568 28578 2660 28580
tri 2660 28578 2662 28580 nw
tri 6727 28578 6729 28580 ne
rect 6729 28578 6821 28580
tri 6821 28578 6823 28580 sw
rect 1821 11128 1856 11192
rect 1920 11128 1936 11192
rect 2000 11128 2016 11192
rect 2080 11128 2096 11192
rect 2160 11128 2176 11192
rect 2240 11128 2256 11192
rect 2320 11128 2336 11192
rect 2400 11128 2421 11192
rect 1821 11097 2421 11128
rect 1821 11033 1856 11097
rect 1920 11033 1936 11097
rect 2000 11033 2016 11097
rect 2080 11033 2096 11097
rect 2160 11033 2176 11097
rect 2240 11033 2256 11097
rect 2320 11033 2336 11097
rect 2400 11033 2421 11097
rect 1821 11001 2421 11033
rect 1821 10937 1856 11001
rect 1920 10937 1936 11001
rect 2000 10937 2016 11001
rect 2080 10937 2096 11001
rect 2160 10937 2176 11001
rect 2240 10937 2256 11001
rect 2320 10937 2336 11001
rect 2400 10937 2421 11001
rect 1821 10905 2421 10937
rect 1821 10841 1856 10905
rect 1920 10841 1936 10905
rect 2000 10841 2016 10905
rect 2080 10841 2096 10905
rect 2160 10841 2176 10905
rect 2240 10841 2256 10905
rect 2320 10841 2336 10905
rect 2400 10841 2421 10905
rect 1821 10809 2421 10841
rect 1821 10745 1856 10809
rect 1920 10745 1936 10809
rect 2000 10745 2016 10809
rect 2080 10745 2096 10809
rect 2160 10745 2176 10809
rect 2240 10745 2256 10809
rect 2320 10745 2336 10809
rect 2400 10745 2421 10809
rect 1821 10713 2421 10745
rect 1821 10649 1856 10713
rect 1920 10649 1936 10713
rect 2000 10649 2016 10713
rect 2080 10649 2096 10713
rect 2160 10649 2176 10713
rect 2240 10649 2256 10713
rect 2320 10649 2336 10713
rect 2400 10649 2421 10713
rect 1821 9547 2421 10649
tri 2521 28533 2566 28578 se
rect 2566 28533 2615 28578
tri 2615 28533 2660 28578 nw
tri 6729 28533 6774 28578 ne
rect 6774 28533 6823 28578
tri 6823 28533 6868 28578 sw
rect 2521 17767 2587 28533
tri 2587 28505 2615 28533 nw
tri 6774 28505 6802 28533 ne
rect 2521 17711 2526 17767
rect 2582 17711 2587 17767
rect 2521 17680 2587 17711
rect 2521 17624 2526 17680
rect 2582 17624 2587 17680
rect 2521 17593 2587 17624
rect 2521 17537 2526 17593
rect 2582 17537 2587 17593
rect 2521 17505 2587 17537
rect 2521 17449 2526 17505
rect 2582 17449 2587 17505
rect 2521 17417 2587 17449
rect 2521 17361 2526 17417
rect 2582 17361 2587 17417
rect 2521 17329 2587 17361
rect 2521 17273 2526 17329
rect 2582 17273 2587 17329
rect 2521 17241 2587 17273
rect 2521 17185 2526 17241
rect 2582 17185 2587 17241
rect 2521 9547 2587 17185
rect 2734 24279 3666 24379
rect 2734 17767 2800 24279
tri 2800 24208 2871 24279 nw
tri 3529 24208 3600 24279 ne
rect 2734 17711 2739 17767
rect 2795 17711 2800 17767
rect 2734 17680 2800 17711
rect 2734 17624 2739 17680
rect 2795 17624 2800 17680
rect 2734 17593 2800 17624
rect 2734 17537 2739 17593
rect 2795 17537 2800 17593
rect 2734 17505 2800 17537
rect 2734 17449 2739 17505
rect 2795 17449 2800 17505
rect 2734 17417 2800 17449
rect 2734 17361 2739 17417
rect 2795 17361 2800 17417
rect 2734 17329 2800 17361
rect 2734 17273 2739 17329
rect 2795 17273 2800 17329
rect 2734 17241 2800 17273
rect 2734 17185 2739 17241
rect 2795 17185 2800 17241
rect 2734 9547 2800 17185
rect 2900 24037 3500 24052
rect 2900 23981 2915 24037
rect 2971 23981 3001 24037
rect 3057 23981 3087 24037
rect 3143 23981 3173 24037
rect 3229 23981 3259 24037
rect 3315 23981 3345 24037
rect 3401 23981 3431 24037
rect 3487 23981 3500 24037
rect 2900 23957 3500 23981
rect 2900 23901 2915 23957
rect 2971 23901 3001 23957
rect 3057 23901 3087 23957
rect 3143 23901 3173 23957
rect 3229 23901 3259 23957
rect 3315 23901 3345 23957
rect 3401 23901 3431 23957
rect 3487 23901 3500 23957
rect 2900 23877 3500 23901
rect 2900 23821 2915 23877
rect 2971 23821 3001 23877
rect 3057 23821 3087 23877
rect 3143 23821 3173 23877
rect 3229 23821 3259 23877
rect 3315 23821 3345 23877
rect 3401 23821 3431 23877
rect 3487 23821 3500 23877
rect 2900 23797 3500 23821
rect 2900 23741 2915 23797
rect 2971 23741 3001 23797
rect 3057 23741 3087 23797
rect 3143 23741 3173 23797
rect 3229 23741 3259 23797
rect 3315 23741 3345 23797
rect 3401 23741 3431 23797
rect 3487 23741 3500 23797
rect 2900 23717 3500 23741
rect 2900 23661 2915 23717
rect 2971 23661 3001 23717
rect 3057 23661 3087 23717
rect 3143 23661 3173 23717
rect 3229 23661 3259 23717
rect 3315 23661 3345 23717
rect 3401 23661 3431 23717
rect 3487 23661 3500 23717
rect 2900 23637 3500 23661
rect 2900 23581 2915 23637
rect 2971 23581 3001 23637
rect 3057 23581 3087 23637
rect 3143 23581 3173 23637
rect 3229 23581 3259 23637
rect 3315 23581 3345 23637
rect 3401 23581 3431 23637
rect 3487 23581 3500 23637
rect 2900 23557 3500 23581
rect 2900 23501 2915 23557
rect 2971 23501 3001 23557
rect 3057 23501 3087 23557
rect 3143 23501 3173 23557
rect 3229 23501 3259 23557
rect 3315 23501 3345 23557
rect 3401 23501 3431 23557
rect 3487 23501 3500 23557
rect 2900 23477 3500 23501
rect 2900 23421 2915 23477
rect 2971 23421 3001 23477
rect 3057 23421 3087 23477
rect 3143 23421 3173 23477
rect 3229 23421 3259 23477
rect 3315 23421 3345 23477
rect 3401 23421 3431 23477
rect 3487 23421 3500 23477
rect 2900 23397 3500 23421
rect 2900 23341 2915 23397
rect 2971 23341 3001 23397
rect 3057 23341 3087 23397
rect 3143 23341 3173 23397
rect 3229 23341 3259 23397
rect 3315 23341 3345 23397
rect 3401 23341 3431 23397
rect 3487 23341 3500 23397
rect 2900 23317 3500 23341
rect 2900 23261 2915 23317
rect 2971 23261 3001 23317
rect 3057 23261 3087 23317
rect 3143 23261 3173 23317
rect 3229 23261 3259 23317
rect 3315 23261 3345 23317
rect 3401 23261 3431 23317
rect 3487 23261 3500 23317
rect 2900 23237 3500 23261
rect 2900 23181 2915 23237
rect 2971 23181 3001 23237
rect 3057 23181 3087 23237
rect 3143 23181 3173 23237
rect 3229 23181 3259 23237
rect 3315 23181 3345 23237
rect 3401 23181 3431 23237
rect 3487 23181 3500 23237
rect 2900 23157 3500 23181
rect 2900 23101 2915 23157
rect 2971 23101 3001 23157
rect 3057 23101 3087 23157
rect 3143 23101 3173 23157
rect 3229 23101 3259 23157
rect 3315 23101 3345 23157
rect 3401 23101 3431 23157
rect 3487 23101 3500 23157
rect 2900 23077 3500 23101
rect 2900 23021 2915 23077
rect 2971 23021 3001 23077
rect 3057 23021 3087 23077
rect 3143 23021 3173 23077
rect 3229 23021 3259 23077
rect 3315 23021 3345 23077
rect 3401 23021 3431 23077
rect 3487 23021 3500 23077
rect 2900 22997 3500 23021
rect 2900 22941 2915 22997
rect 2971 22941 3001 22997
rect 3057 22941 3087 22997
rect 3143 22941 3173 22997
rect 3229 22941 3259 22997
rect 3315 22941 3345 22997
rect 3401 22941 3431 22997
rect 3487 22941 3500 22997
rect 2900 22917 3500 22941
rect 2900 22861 2915 22917
rect 2971 22861 3001 22917
rect 3057 22861 3087 22917
rect 3143 22861 3173 22917
rect 3229 22861 3259 22917
rect 3315 22861 3345 22917
rect 3401 22861 3431 22917
rect 3487 22861 3500 22917
rect 2900 22837 3500 22861
rect 2900 22781 2915 22837
rect 2971 22781 3001 22837
rect 3057 22781 3087 22837
rect 3143 22781 3173 22837
rect 3229 22781 3259 22837
rect 3315 22781 3345 22837
rect 3401 22781 3431 22837
rect 3487 22781 3500 22837
rect 2900 22757 3500 22781
rect 2900 22701 2915 22757
rect 2971 22701 3001 22757
rect 3057 22701 3087 22757
rect 3143 22701 3173 22757
rect 3229 22701 3259 22757
rect 3315 22701 3345 22757
rect 3401 22701 3431 22757
rect 3487 22701 3500 22757
rect 2900 22677 3500 22701
rect 2900 22621 2915 22677
rect 2971 22621 3001 22677
rect 3057 22621 3087 22677
rect 3143 22621 3173 22677
rect 3229 22621 3259 22677
rect 3315 22621 3345 22677
rect 3401 22621 3431 22677
rect 3487 22621 3500 22677
rect 2900 22597 3500 22621
rect 2900 22541 2915 22597
rect 2971 22541 3001 22597
rect 3057 22541 3087 22597
rect 3143 22541 3173 22597
rect 3229 22541 3259 22597
rect 3315 22541 3345 22597
rect 3401 22541 3431 22597
rect 3487 22541 3500 22597
rect 2900 22517 3500 22541
rect 2900 22461 2915 22517
rect 2971 22461 3001 22517
rect 3057 22461 3087 22517
rect 3143 22461 3173 22517
rect 3229 22461 3259 22517
rect 3315 22461 3345 22517
rect 3401 22461 3431 22517
rect 3487 22461 3500 22517
rect 2900 22437 3500 22461
rect 2900 22381 2915 22437
rect 2971 22381 3001 22437
rect 3057 22381 3087 22437
rect 3143 22381 3173 22437
rect 3229 22381 3259 22437
rect 3315 22381 3345 22437
rect 3401 22381 3431 22437
rect 3487 22381 3500 22437
rect 2900 22357 3500 22381
rect 2900 22301 2915 22357
rect 2971 22301 3001 22357
rect 3057 22301 3087 22357
rect 3143 22301 3173 22357
rect 3229 22301 3259 22357
rect 3315 22301 3345 22357
rect 3401 22301 3431 22357
rect 3487 22301 3500 22357
rect 2900 22277 3500 22301
rect 2900 22221 2915 22277
rect 2971 22221 3001 22277
rect 3057 22221 3087 22277
rect 3143 22221 3173 22277
rect 3229 22221 3259 22277
rect 3315 22221 3345 22277
rect 3401 22221 3431 22277
rect 3487 22221 3500 22277
rect 2900 22197 3500 22221
rect 2900 22141 2915 22197
rect 2971 22141 3001 22197
rect 3057 22141 3087 22197
rect 3143 22141 3173 22197
rect 3229 22141 3259 22197
rect 3315 22141 3345 22197
rect 3401 22141 3431 22197
rect 3487 22141 3500 22197
rect 2900 22117 3500 22141
rect 2900 22061 2915 22117
rect 2971 22061 3001 22117
rect 3057 22061 3087 22117
rect 3143 22061 3173 22117
rect 3229 22061 3259 22117
rect 3315 22061 3345 22117
rect 3401 22061 3431 22117
rect 3487 22061 3500 22117
rect 2900 22037 3500 22061
rect 2900 21981 2915 22037
rect 2971 21981 3001 22037
rect 3057 21981 3087 22037
rect 3143 21981 3173 22037
rect 3229 21981 3259 22037
rect 3315 21981 3345 22037
rect 3401 21981 3431 22037
rect 3487 21981 3500 22037
rect 2900 21957 3500 21981
rect 2900 21901 2915 21957
rect 2971 21901 3001 21957
rect 3057 21901 3087 21957
rect 3143 21901 3173 21957
rect 3229 21901 3259 21957
rect 3315 21901 3345 21957
rect 3401 21901 3431 21957
rect 3487 21901 3500 21957
rect 2900 21877 3500 21901
rect 2900 21821 2915 21877
rect 2971 21821 3001 21877
rect 3057 21821 3087 21877
rect 3143 21821 3173 21877
rect 3229 21821 3259 21877
rect 3315 21821 3345 21877
rect 3401 21821 3431 21877
rect 3487 21821 3500 21877
rect 2900 21797 3500 21821
rect 2900 21741 2915 21797
rect 2971 21741 3001 21797
rect 3057 21741 3087 21797
rect 3143 21741 3173 21797
rect 3229 21741 3259 21797
rect 3315 21741 3345 21797
rect 3401 21741 3431 21797
rect 3487 21741 3500 21797
rect 2900 21717 3500 21741
rect 2900 21661 2915 21717
rect 2971 21661 3001 21717
rect 3057 21661 3087 21717
rect 3143 21661 3173 21717
rect 3229 21661 3259 21717
rect 3315 21661 3345 21717
rect 3401 21661 3431 21717
rect 3487 21661 3500 21717
rect 2900 21637 3500 21661
rect 2900 21581 2915 21637
rect 2971 21581 3001 21637
rect 3057 21581 3087 21637
rect 3143 21581 3173 21637
rect 3229 21581 3259 21637
rect 3315 21581 3345 21637
rect 3401 21581 3431 21637
rect 3487 21581 3500 21637
rect 2900 21557 3500 21581
rect 2900 21501 2915 21557
rect 2971 21501 3001 21557
rect 3057 21501 3087 21557
rect 3143 21501 3173 21557
rect 3229 21501 3259 21557
rect 3315 21501 3345 21557
rect 3401 21501 3431 21557
rect 3487 21501 3500 21557
rect 2900 21477 3500 21501
rect 2900 21421 2915 21477
rect 2971 21421 3001 21477
rect 3057 21421 3087 21477
rect 3143 21421 3173 21477
rect 3229 21421 3259 21477
rect 3315 21421 3345 21477
rect 3401 21421 3431 21477
rect 3487 21421 3500 21477
rect 2900 21397 3500 21421
rect 2900 21341 2915 21397
rect 2971 21341 3001 21397
rect 3057 21341 3087 21397
rect 3143 21341 3173 21397
rect 3229 21341 3259 21397
rect 3315 21341 3345 21397
rect 3401 21341 3431 21397
rect 3487 21341 3500 21397
rect 2900 21317 3500 21341
rect 2900 21261 2915 21317
rect 2971 21261 3001 21317
rect 3057 21261 3087 21317
rect 3143 21261 3173 21317
rect 3229 21261 3259 21317
rect 3315 21261 3345 21317
rect 3401 21261 3431 21317
rect 3487 21261 3500 21317
rect 2900 21237 3500 21261
rect 2900 21181 2915 21237
rect 2971 21181 3001 21237
rect 3057 21181 3087 21237
rect 3143 21181 3173 21237
rect 3229 21181 3259 21237
rect 3315 21181 3345 21237
rect 3401 21181 3431 21237
rect 3487 21181 3500 21237
rect 2900 21157 3500 21181
rect 2900 21101 2915 21157
rect 2971 21101 3001 21157
rect 3057 21101 3087 21157
rect 3143 21101 3173 21157
rect 3229 21101 3259 21157
rect 3315 21101 3345 21157
rect 3401 21101 3431 21157
rect 3487 21101 3500 21157
rect 2900 21077 3500 21101
rect 2900 21021 2915 21077
rect 2971 21021 3001 21077
rect 3057 21021 3087 21077
rect 3143 21021 3173 21077
rect 3229 21021 3259 21077
rect 3315 21021 3345 21077
rect 3401 21021 3431 21077
rect 3487 21021 3500 21077
rect 2900 20997 3500 21021
rect 2900 20941 2915 20997
rect 2971 20941 3001 20997
rect 3057 20941 3087 20997
rect 3143 20941 3173 20997
rect 3229 20941 3259 20997
rect 3315 20941 3345 20997
rect 3401 20941 3431 20997
rect 3487 20941 3500 20997
rect 2900 20917 3500 20941
rect 2900 20861 2915 20917
rect 2971 20861 3001 20917
rect 3057 20861 3087 20917
rect 3143 20861 3173 20917
rect 3229 20861 3259 20917
rect 3315 20861 3345 20917
rect 3401 20861 3431 20917
rect 3487 20861 3500 20917
rect 2900 20837 3500 20861
rect 2900 20781 2915 20837
rect 2971 20781 3001 20837
rect 3057 20781 3087 20837
rect 3143 20781 3173 20837
rect 3229 20781 3259 20837
rect 3315 20781 3345 20837
rect 3401 20781 3431 20837
rect 3487 20781 3500 20837
rect 2900 20757 3500 20781
rect 2900 20701 2915 20757
rect 2971 20701 3001 20757
rect 3057 20701 3087 20757
rect 3143 20701 3173 20757
rect 3229 20701 3259 20757
rect 3315 20701 3345 20757
rect 3401 20701 3431 20757
rect 3487 20701 3500 20757
rect 2900 20677 3500 20701
rect 2900 20621 2915 20677
rect 2971 20621 3001 20677
rect 3057 20621 3087 20677
rect 3143 20621 3173 20677
rect 3229 20621 3259 20677
rect 3315 20621 3345 20677
rect 3401 20621 3431 20677
rect 3487 20621 3500 20677
rect 2900 20597 3500 20621
rect 2900 20541 2915 20597
rect 2971 20541 3001 20597
rect 3057 20541 3087 20597
rect 3143 20541 3173 20597
rect 3229 20541 3259 20597
rect 3315 20541 3345 20597
rect 3401 20541 3431 20597
rect 3487 20541 3500 20597
rect 2900 20517 3500 20541
rect 2900 20461 2915 20517
rect 2971 20461 3001 20517
rect 3057 20461 3087 20517
rect 3143 20461 3173 20517
rect 3229 20461 3259 20517
rect 3315 20461 3345 20517
rect 3401 20461 3431 20517
rect 3487 20461 3500 20517
rect 2900 20437 3500 20461
rect 2900 20381 2915 20437
rect 2971 20381 3001 20437
rect 3057 20381 3087 20437
rect 3143 20381 3173 20437
rect 3229 20381 3259 20437
rect 3315 20381 3345 20437
rect 3401 20381 3431 20437
rect 3487 20381 3500 20437
rect 2900 20357 3500 20381
rect 2900 20301 2915 20357
rect 2971 20301 3001 20357
rect 3057 20301 3087 20357
rect 3143 20301 3173 20357
rect 3229 20301 3259 20357
rect 3315 20301 3345 20357
rect 3401 20301 3431 20357
rect 3487 20301 3500 20357
rect 2900 20277 3500 20301
rect 2900 20221 2915 20277
rect 2971 20221 3001 20277
rect 3057 20221 3087 20277
rect 3143 20221 3173 20277
rect 3229 20221 3259 20277
rect 3315 20221 3345 20277
rect 3401 20221 3431 20277
rect 3487 20221 3500 20277
rect 2900 20197 3500 20221
rect 2900 20141 2915 20197
rect 2971 20141 3001 20197
rect 3057 20141 3087 20197
rect 3143 20141 3173 20197
rect 3229 20141 3259 20197
rect 3315 20141 3345 20197
rect 3401 20141 3431 20197
rect 3487 20141 3500 20197
rect 2900 20117 3500 20141
rect 2900 20061 2915 20117
rect 2971 20061 3001 20117
rect 3057 20061 3087 20117
rect 3143 20061 3173 20117
rect 3229 20061 3259 20117
rect 3315 20061 3345 20117
rect 3401 20061 3431 20117
rect 3487 20061 3500 20117
rect 2900 20037 3500 20061
rect 2900 19981 2915 20037
rect 2971 19981 3001 20037
rect 3057 19981 3087 20037
rect 3143 19981 3173 20037
rect 3229 19981 3259 20037
rect 3315 19981 3345 20037
rect 3401 19981 3431 20037
rect 3487 19981 3500 20037
rect 2900 19957 3500 19981
rect 2900 19901 2915 19957
rect 2971 19901 3001 19957
rect 3057 19901 3087 19957
rect 3143 19901 3173 19957
rect 3229 19901 3259 19957
rect 3315 19901 3345 19957
rect 3401 19901 3431 19957
rect 3487 19901 3500 19957
rect 2900 19877 3500 19901
rect 2900 19821 2915 19877
rect 2971 19821 3001 19877
rect 3057 19821 3087 19877
rect 3143 19821 3173 19877
rect 3229 19821 3259 19877
rect 3315 19821 3345 19877
rect 3401 19821 3431 19877
rect 3487 19821 3500 19877
rect 2900 19797 3500 19821
rect 2900 19741 2915 19797
rect 2971 19741 3001 19797
rect 3057 19741 3087 19797
rect 3143 19741 3173 19797
rect 3229 19741 3259 19797
rect 3315 19741 3345 19797
rect 3401 19741 3431 19797
rect 3487 19741 3500 19797
rect 2900 19717 3500 19741
rect 2900 19661 2915 19717
rect 2971 19661 3001 19717
rect 3057 19661 3087 19717
rect 3143 19661 3173 19717
rect 3229 19661 3259 19717
rect 3315 19661 3345 19717
rect 3401 19661 3431 19717
rect 3487 19661 3500 19717
rect 2900 19637 3500 19661
rect 2900 19581 2915 19637
rect 2971 19581 3001 19637
rect 3057 19581 3087 19637
rect 3143 19581 3173 19637
rect 3229 19581 3259 19637
rect 3315 19581 3345 19637
rect 3401 19581 3431 19637
rect 3487 19581 3500 19637
rect 2900 19557 3500 19581
rect 2900 19501 2915 19557
rect 2971 19501 3001 19557
rect 3057 19501 3087 19557
rect 3143 19501 3173 19557
rect 3229 19501 3259 19557
rect 3315 19501 3345 19557
rect 3401 19501 3431 19557
rect 3487 19501 3500 19557
rect 2900 19477 3500 19501
rect 2900 19421 2915 19477
rect 2971 19421 3001 19477
rect 3057 19421 3087 19477
rect 3143 19421 3173 19477
rect 3229 19421 3259 19477
rect 3315 19421 3345 19477
rect 3401 19421 3431 19477
rect 3487 19421 3500 19477
rect 2900 19397 3500 19421
rect 2900 19341 2915 19397
rect 2971 19341 3001 19397
rect 3057 19341 3087 19397
rect 3143 19341 3173 19397
rect 3229 19341 3259 19397
rect 3315 19341 3345 19397
rect 3401 19341 3431 19397
rect 3487 19341 3500 19397
rect 2900 19317 3500 19341
rect 2900 19261 2915 19317
rect 2971 19261 3001 19317
rect 3057 19261 3087 19317
rect 3143 19261 3173 19317
rect 3229 19261 3259 19317
rect 3315 19261 3345 19317
rect 3401 19261 3431 19317
rect 3487 19261 3500 19317
rect 2900 10244 3500 19261
rect 2900 10180 2921 10244
rect 2985 10180 3001 10244
rect 3065 10180 3081 10244
rect 3145 10180 3161 10244
rect 3225 10180 3241 10244
rect 3305 10180 3321 10244
rect 3385 10180 3401 10244
rect 3465 10180 3500 10244
rect 2900 10149 3500 10180
rect 2900 10085 2921 10149
rect 2985 10085 3001 10149
rect 3065 10085 3081 10149
rect 3145 10085 3161 10149
rect 3225 10085 3241 10149
rect 3305 10085 3321 10149
rect 3385 10085 3401 10149
rect 3465 10085 3500 10149
rect 2900 10053 3500 10085
rect 2900 9989 2921 10053
rect 2985 9989 3001 10053
rect 3065 9989 3081 10053
rect 3145 9989 3161 10053
rect 3225 9989 3241 10053
rect 3305 9989 3321 10053
rect 3385 9989 3401 10053
rect 3465 9989 3500 10053
rect 2900 9957 3500 9989
rect 2900 9893 2921 9957
rect 2985 9893 3001 9957
rect 3065 9893 3081 9957
rect 3145 9893 3161 9957
rect 3225 9893 3241 9957
rect 3305 9893 3321 9957
rect 3385 9893 3401 9957
rect 3465 9893 3500 9957
rect 2900 9861 3500 9893
rect 2900 9797 2921 9861
rect 2985 9797 3001 9861
rect 3065 9797 3081 9861
rect 3145 9797 3161 9861
rect 3225 9797 3241 9861
rect 3305 9797 3321 9861
rect 3385 9797 3401 9861
rect 3465 9797 3500 9861
rect 2900 9765 3500 9797
rect 2900 9701 2921 9765
rect 2985 9701 3001 9765
rect 3065 9701 3081 9765
rect 3145 9701 3161 9765
rect 3225 9701 3241 9765
rect 3305 9701 3321 9765
rect 3385 9701 3401 9765
rect 3465 9701 3500 9765
rect 2900 9547 3500 9701
rect 3600 17767 3666 24279
rect 5723 24279 6655 24379
rect 3600 17711 3605 17767
rect 3661 17711 3666 17767
rect 3600 17680 3666 17711
rect 3600 17624 3605 17680
rect 3661 17624 3666 17680
rect 3600 17593 3666 17624
rect 3600 17537 3605 17593
rect 3661 17537 3666 17593
rect 3600 17505 3666 17537
rect 3600 17449 3605 17505
rect 3661 17449 3666 17505
rect 3600 17417 3666 17449
rect 3600 17361 3605 17417
rect 3661 17361 3666 17417
rect 3600 17329 3666 17361
rect 3600 17273 3605 17329
rect 3661 17273 3666 17329
rect 3600 17241 3666 17273
rect 3600 17185 3605 17241
rect 3661 17185 3666 17241
rect 3600 9547 3666 17185
rect 4998 18623 5198 18659
rect 4998 18567 5007 18623
rect 5063 18567 5133 18623
rect 5189 18567 5198 18623
rect 4998 16481 5198 18567
rect 4998 16425 5003 16481
rect 5059 16425 5137 16481
rect 5193 16425 5198 16481
rect 4998 16420 5198 16425
rect 5723 17767 5789 24279
tri 5789 24208 5860 24279 nw
tri 6518 24208 6589 24279 ne
rect 5723 17711 5728 17767
rect 5784 17711 5789 17767
rect 5723 17680 5789 17711
rect 5723 17624 5728 17680
rect 5784 17624 5789 17680
rect 5723 17593 5789 17624
rect 5723 17537 5728 17593
rect 5784 17537 5789 17593
rect 5723 17505 5789 17537
rect 5723 17449 5728 17505
rect 5784 17449 5789 17505
rect 5723 17417 5789 17449
rect 5723 17361 5728 17417
rect 5784 17361 5789 17417
rect 5723 17329 5789 17361
rect 5723 17273 5728 17329
rect 5784 17273 5789 17329
rect 5723 17241 5789 17273
rect 5723 17185 5728 17241
rect 5784 17185 5789 17241
rect 4416 15566 4616 16094
rect 4416 15510 4425 15566
rect 4481 15510 4551 15566
rect 4607 15510 4616 15566
rect 4416 15486 4616 15510
rect 4416 15430 4425 15486
rect 4481 15430 4551 15486
rect 4607 15430 4616 15486
rect 4416 14423 4616 15430
rect 4416 14367 4425 14423
rect 4481 14367 4551 14423
rect 4607 14367 4616 14423
rect 4416 14343 4616 14367
rect 4416 14287 4425 14343
rect 4481 14287 4551 14343
rect 4607 14287 4616 14343
rect 4416 13042 4616 14287
rect 4416 12986 4425 13042
rect 4481 12986 4551 13042
rect 4607 12986 4616 13042
rect 4416 12962 4616 12986
rect 4416 12906 4425 12962
rect 4481 12906 4551 12962
rect 4607 12906 4616 12962
rect 4416 11909 4616 12906
rect 4416 11853 4425 11909
rect 4481 11853 4551 11909
rect 4607 11853 4616 11909
rect 4416 11829 4616 11853
rect 4416 11773 4425 11829
rect 4481 11773 4551 11829
rect 4607 11773 4616 11829
rect 4416 11461 4616 11773
rect 4416 11405 4436 11461
rect 4492 11405 4551 11461
rect 4607 11405 4616 11461
rect 4416 11381 4616 11405
rect 4416 11325 4436 11381
rect 4492 11325 4551 11381
rect 4607 11325 4616 11381
rect 4416 10511 4616 11325
rect 4416 10455 4425 10511
rect 4481 10455 4551 10511
rect 4607 10455 4616 10511
rect 4416 10431 4616 10455
rect 4416 10375 4425 10431
rect 4481 10375 4551 10431
rect 4607 10375 4616 10431
rect 954 9436 963 9492
rect 1019 9436 1069 9492
rect 1125 9436 1174 9492
rect 1230 9436 1279 9492
rect 1335 9436 1384 9492
rect 1440 9436 1489 9492
rect 1545 9436 1554 9492
rect 954 7810 1554 9436
rect 4416 9389 4616 10375
rect 5723 9547 5789 17185
rect 5889 24037 6489 24052
rect 5889 23981 5903 24037
rect 5959 23981 5989 24037
rect 6045 23981 6075 24037
rect 6131 23981 6161 24037
rect 6217 23981 6247 24037
rect 6303 23981 6333 24037
rect 6389 23981 6419 24037
rect 6475 23981 6489 24037
rect 5889 23957 6489 23981
rect 5889 23901 5903 23957
rect 5959 23901 5989 23957
rect 6045 23901 6075 23957
rect 6131 23901 6161 23957
rect 6217 23901 6247 23957
rect 6303 23901 6333 23957
rect 6389 23901 6419 23957
rect 6475 23901 6489 23957
rect 5889 23877 6489 23901
rect 5889 23821 5903 23877
rect 5959 23821 5989 23877
rect 6045 23821 6075 23877
rect 6131 23821 6161 23877
rect 6217 23821 6247 23877
rect 6303 23821 6333 23877
rect 6389 23821 6419 23877
rect 6475 23821 6489 23877
rect 5889 23797 6489 23821
rect 5889 23741 5903 23797
rect 5959 23741 5989 23797
rect 6045 23741 6075 23797
rect 6131 23741 6161 23797
rect 6217 23741 6247 23797
rect 6303 23741 6333 23797
rect 6389 23741 6419 23797
rect 6475 23741 6489 23797
rect 5889 23717 6489 23741
rect 5889 23661 5903 23717
rect 5959 23661 5989 23717
rect 6045 23661 6075 23717
rect 6131 23661 6161 23717
rect 6217 23661 6247 23717
rect 6303 23661 6333 23717
rect 6389 23661 6419 23717
rect 6475 23661 6489 23717
rect 5889 23637 6489 23661
rect 5889 23581 5903 23637
rect 5959 23581 5989 23637
rect 6045 23581 6075 23637
rect 6131 23581 6161 23637
rect 6217 23581 6247 23637
rect 6303 23581 6333 23637
rect 6389 23581 6419 23637
rect 6475 23581 6489 23637
rect 5889 23557 6489 23581
rect 5889 23501 5903 23557
rect 5959 23501 5989 23557
rect 6045 23501 6075 23557
rect 6131 23501 6161 23557
rect 6217 23501 6247 23557
rect 6303 23501 6333 23557
rect 6389 23501 6419 23557
rect 6475 23501 6489 23557
rect 5889 23477 6489 23501
rect 5889 23421 5903 23477
rect 5959 23421 5989 23477
rect 6045 23421 6075 23477
rect 6131 23421 6161 23477
rect 6217 23421 6247 23477
rect 6303 23421 6333 23477
rect 6389 23421 6419 23477
rect 6475 23421 6489 23477
rect 5889 23397 6489 23421
rect 5889 23341 5903 23397
rect 5959 23341 5989 23397
rect 6045 23341 6075 23397
rect 6131 23341 6161 23397
rect 6217 23341 6247 23397
rect 6303 23341 6333 23397
rect 6389 23341 6419 23397
rect 6475 23341 6489 23397
rect 5889 23317 6489 23341
rect 5889 23261 5903 23317
rect 5959 23261 5989 23317
rect 6045 23261 6075 23317
rect 6131 23261 6161 23317
rect 6217 23261 6247 23317
rect 6303 23261 6333 23317
rect 6389 23261 6419 23317
rect 6475 23261 6489 23317
rect 5889 23237 6489 23261
rect 5889 23181 5903 23237
rect 5959 23181 5989 23237
rect 6045 23181 6075 23237
rect 6131 23181 6161 23237
rect 6217 23181 6247 23237
rect 6303 23181 6333 23237
rect 6389 23181 6419 23237
rect 6475 23181 6489 23237
rect 5889 23157 6489 23181
rect 5889 23101 5903 23157
rect 5959 23101 5989 23157
rect 6045 23101 6075 23157
rect 6131 23101 6161 23157
rect 6217 23101 6247 23157
rect 6303 23101 6333 23157
rect 6389 23101 6419 23157
rect 6475 23101 6489 23157
rect 5889 23077 6489 23101
rect 5889 23021 5903 23077
rect 5959 23021 5989 23077
rect 6045 23021 6075 23077
rect 6131 23021 6161 23077
rect 6217 23021 6247 23077
rect 6303 23021 6333 23077
rect 6389 23021 6419 23077
rect 6475 23021 6489 23077
rect 5889 22997 6489 23021
rect 5889 22941 5903 22997
rect 5959 22941 5989 22997
rect 6045 22941 6075 22997
rect 6131 22941 6161 22997
rect 6217 22941 6247 22997
rect 6303 22941 6333 22997
rect 6389 22941 6419 22997
rect 6475 22941 6489 22997
rect 5889 22917 6489 22941
rect 5889 22861 5903 22917
rect 5959 22861 5989 22917
rect 6045 22861 6075 22917
rect 6131 22861 6161 22917
rect 6217 22861 6247 22917
rect 6303 22861 6333 22917
rect 6389 22861 6419 22917
rect 6475 22861 6489 22917
rect 5889 22837 6489 22861
rect 5889 22781 5903 22837
rect 5959 22781 5989 22837
rect 6045 22781 6075 22837
rect 6131 22781 6161 22837
rect 6217 22781 6247 22837
rect 6303 22781 6333 22837
rect 6389 22781 6419 22837
rect 6475 22781 6489 22837
rect 5889 22757 6489 22781
rect 5889 22701 5903 22757
rect 5959 22701 5989 22757
rect 6045 22701 6075 22757
rect 6131 22701 6161 22757
rect 6217 22701 6247 22757
rect 6303 22701 6333 22757
rect 6389 22701 6419 22757
rect 6475 22701 6489 22757
rect 5889 22677 6489 22701
rect 5889 22621 5903 22677
rect 5959 22621 5989 22677
rect 6045 22621 6075 22677
rect 6131 22621 6161 22677
rect 6217 22621 6247 22677
rect 6303 22621 6333 22677
rect 6389 22621 6419 22677
rect 6475 22621 6489 22677
rect 5889 22597 6489 22621
rect 5889 22541 5903 22597
rect 5959 22541 5989 22597
rect 6045 22541 6075 22597
rect 6131 22541 6161 22597
rect 6217 22541 6247 22597
rect 6303 22541 6333 22597
rect 6389 22541 6419 22597
rect 6475 22541 6489 22597
rect 5889 22517 6489 22541
rect 5889 22461 5903 22517
rect 5959 22461 5989 22517
rect 6045 22461 6075 22517
rect 6131 22461 6161 22517
rect 6217 22461 6247 22517
rect 6303 22461 6333 22517
rect 6389 22461 6419 22517
rect 6475 22461 6489 22517
rect 5889 22437 6489 22461
rect 5889 22381 5903 22437
rect 5959 22381 5989 22437
rect 6045 22381 6075 22437
rect 6131 22381 6161 22437
rect 6217 22381 6247 22437
rect 6303 22381 6333 22437
rect 6389 22381 6419 22437
rect 6475 22381 6489 22437
rect 5889 22357 6489 22381
rect 5889 22301 5903 22357
rect 5959 22301 5989 22357
rect 6045 22301 6075 22357
rect 6131 22301 6161 22357
rect 6217 22301 6247 22357
rect 6303 22301 6333 22357
rect 6389 22301 6419 22357
rect 6475 22301 6489 22357
rect 5889 22277 6489 22301
rect 5889 22221 5903 22277
rect 5959 22221 5989 22277
rect 6045 22221 6075 22277
rect 6131 22221 6161 22277
rect 6217 22221 6247 22277
rect 6303 22221 6333 22277
rect 6389 22221 6419 22277
rect 6475 22221 6489 22277
rect 5889 22197 6489 22221
rect 5889 22141 5903 22197
rect 5959 22141 5989 22197
rect 6045 22141 6075 22197
rect 6131 22141 6161 22197
rect 6217 22141 6247 22197
rect 6303 22141 6333 22197
rect 6389 22141 6419 22197
rect 6475 22141 6489 22197
rect 5889 22117 6489 22141
rect 5889 22061 5903 22117
rect 5959 22061 5989 22117
rect 6045 22061 6075 22117
rect 6131 22061 6161 22117
rect 6217 22061 6247 22117
rect 6303 22061 6333 22117
rect 6389 22061 6419 22117
rect 6475 22061 6489 22117
rect 5889 22037 6489 22061
rect 5889 21981 5903 22037
rect 5959 21981 5989 22037
rect 6045 21981 6075 22037
rect 6131 21981 6161 22037
rect 6217 21981 6247 22037
rect 6303 21981 6333 22037
rect 6389 21981 6419 22037
rect 6475 21981 6489 22037
rect 5889 21957 6489 21981
rect 5889 21901 5903 21957
rect 5959 21901 5989 21957
rect 6045 21901 6075 21957
rect 6131 21901 6161 21957
rect 6217 21901 6247 21957
rect 6303 21901 6333 21957
rect 6389 21901 6419 21957
rect 6475 21901 6489 21957
rect 5889 21877 6489 21901
rect 5889 21821 5903 21877
rect 5959 21821 5989 21877
rect 6045 21821 6075 21877
rect 6131 21821 6161 21877
rect 6217 21821 6247 21877
rect 6303 21821 6333 21877
rect 6389 21821 6419 21877
rect 6475 21821 6489 21877
rect 5889 21797 6489 21821
rect 5889 21741 5903 21797
rect 5959 21741 5989 21797
rect 6045 21741 6075 21797
rect 6131 21741 6161 21797
rect 6217 21741 6247 21797
rect 6303 21741 6333 21797
rect 6389 21741 6419 21797
rect 6475 21741 6489 21797
rect 5889 21717 6489 21741
rect 5889 21661 5903 21717
rect 5959 21661 5989 21717
rect 6045 21661 6075 21717
rect 6131 21661 6161 21717
rect 6217 21661 6247 21717
rect 6303 21661 6333 21717
rect 6389 21661 6419 21717
rect 6475 21661 6489 21717
rect 5889 21637 6489 21661
rect 5889 21581 5903 21637
rect 5959 21581 5989 21637
rect 6045 21581 6075 21637
rect 6131 21581 6161 21637
rect 6217 21581 6247 21637
rect 6303 21581 6333 21637
rect 6389 21581 6419 21637
rect 6475 21581 6489 21637
rect 5889 21557 6489 21581
rect 5889 21501 5903 21557
rect 5959 21501 5989 21557
rect 6045 21501 6075 21557
rect 6131 21501 6161 21557
rect 6217 21501 6247 21557
rect 6303 21501 6333 21557
rect 6389 21501 6419 21557
rect 6475 21501 6489 21557
rect 5889 21477 6489 21501
rect 5889 21421 5903 21477
rect 5959 21421 5989 21477
rect 6045 21421 6075 21477
rect 6131 21421 6161 21477
rect 6217 21421 6247 21477
rect 6303 21421 6333 21477
rect 6389 21421 6419 21477
rect 6475 21421 6489 21477
rect 5889 21397 6489 21421
rect 5889 21341 5903 21397
rect 5959 21341 5989 21397
rect 6045 21341 6075 21397
rect 6131 21341 6161 21397
rect 6217 21341 6247 21397
rect 6303 21341 6333 21397
rect 6389 21341 6419 21397
rect 6475 21341 6489 21397
rect 5889 21317 6489 21341
rect 5889 21261 5903 21317
rect 5959 21261 5989 21317
rect 6045 21261 6075 21317
rect 6131 21261 6161 21317
rect 6217 21261 6247 21317
rect 6303 21261 6333 21317
rect 6389 21261 6419 21317
rect 6475 21261 6489 21317
rect 5889 21237 6489 21261
rect 5889 21181 5903 21237
rect 5959 21181 5989 21237
rect 6045 21181 6075 21237
rect 6131 21181 6161 21237
rect 6217 21181 6247 21237
rect 6303 21181 6333 21237
rect 6389 21181 6419 21237
rect 6475 21181 6489 21237
rect 5889 21157 6489 21181
rect 5889 21101 5903 21157
rect 5959 21101 5989 21157
rect 6045 21101 6075 21157
rect 6131 21101 6161 21157
rect 6217 21101 6247 21157
rect 6303 21101 6333 21157
rect 6389 21101 6419 21157
rect 6475 21101 6489 21157
rect 5889 21077 6489 21101
rect 5889 21021 5903 21077
rect 5959 21021 5989 21077
rect 6045 21021 6075 21077
rect 6131 21021 6161 21077
rect 6217 21021 6247 21077
rect 6303 21021 6333 21077
rect 6389 21021 6419 21077
rect 6475 21021 6489 21077
rect 5889 20997 6489 21021
rect 5889 20941 5903 20997
rect 5959 20941 5989 20997
rect 6045 20941 6075 20997
rect 6131 20941 6161 20997
rect 6217 20941 6247 20997
rect 6303 20941 6333 20997
rect 6389 20941 6419 20997
rect 6475 20941 6489 20997
rect 5889 20917 6489 20941
rect 5889 20861 5903 20917
rect 5959 20861 5989 20917
rect 6045 20861 6075 20917
rect 6131 20861 6161 20917
rect 6217 20861 6247 20917
rect 6303 20861 6333 20917
rect 6389 20861 6419 20917
rect 6475 20861 6489 20917
rect 5889 20837 6489 20861
rect 5889 20781 5903 20837
rect 5959 20781 5989 20837
rect 6045 20781 6075 20837
rect 6131 20781 6161 20837
rect 6217 20781 6247 20837
rect 6303 20781 6333 20837
rect 6389 20781 6419 20837
rect 6475 20781 6489 20837
rect 5889 20757 6489 20781
rect 5889 20701 5903 20757
rect 5959 20701 5989 20757
rect 6045 20701 6075 20757
rect 6131 20701 6161 20757
rect 6217 20701 6247 20757
rect 6303 20701 6333 20757
rect 6389 20701 6419 20757
rect 6475 20701 6489 20757
rect 5889 20677 6489 20701
rect 5889 20621 5903 20677
rect 5959 20621 5989 20677
rect 6045 20621 6075 20677
rect 6131 20621 6161 20677
rect 6217 20621 6247 20677
rect 6303 20621 6333 20677
rect 6389 20621 6419 20677
rect 6475 20621 6489 20677
rect 5889 20597 6489 20621
rect 5889 20541 5903 20597
rect 5959 20541 5989 20597
rect 6045 20541 6075 20597
rect 6131 20541 6161 20597
rect 6217 20541 6247 20597
rect 6303 20541 6333 20597
rect 6389 20541 6419 20597
rect 6475 20541 6489 20597
rect 5889 20517 6489 20541
rect 5889 20461 5903 20517
rect 5959 20461 5989 20517
rect 6045 20461 6075 20517
rect 6131 20461 6161 20517
rect 6217 20461 6247 20517
rect 6303 20461 6333 20517
rect 6389 20461 6419 20517
rect 6475 20461 6489 20517
rect 5889 20437 6489 20461
rect 5889 20381 5903 20437
rect 5959 20381 5989 20437
rect 6045 20381 6075 20437
rect 6131 20381 6161 20437
rect 6217 20381 6247 20437
rect 6303 20381 6333 20437
rect 6389 20381 6419 20437
rect 6475 20381 6489 20437
rect 5889 20357 6489 20381
rect 5889 20301 5903 20357
rect 5959 20301 5989 20357
rect 6045 20301 6075 20357
rect 6131 20301 6161 20357
rect 6217 20301 6247 20357
rect 6303 20301 6333 20357
rect 6389 20301 6419 20357
rect 6475 20301 6489 20357
rect 5889 20277 6489 20301
rect 5889 20221 5903 20277
rect 5959 20221 5989 20277
rect 6045 20221 6075 20277
rect 6131 20221 6161 20277
rect 6217 20221 6247 20277
rect 6303 20221 6333 20277
rect 6389 20221 6419 20277
rect 6475 20221 6489 20277
rect 5889 20197 6489 20221
rect 5889 20141 5903 20197
rect 5959 20141 5989 20197
rect 6045 20141 6075 20197
rect 6131 20141 6161 20197
rect 6217 20141 6247 20197
rect 6303 20141 6333 20197
rect 6389 20141 6419 20197
rect 6475 20141 6489 20197
rect 5889 20117 6489 20141
rect 5889 20061 5903 20117
rect 5959 20061 5989 20117
rect 6045 20061 6075 20117
rect 6131 20061 6161 20117
rect 6217 20061 6247 20117
rect 6303 20061 6333 20117
rect 6389 20061 6419 20117
rect 6475 20061 6489 20117
rect 5889 20037 6489 20061
rect 5889 19981 5903 20037
rect 5959 19981 5989 20037
rect 6045 19981 6075 20037
rect 6131 19981 6161 20037
rect 6217 19981 6247 20037
rect 6303 19981 6333 20037
rect 6389 19981 6419 20037
rect 6475 19981 6489 20037
rect 5889 19957 6489 19981
rect 5889 19901 5903 19957
rect 5959 19901 5989 19957
rect 6045 19901 6075 19957
rect 6131 19901 6161 19957
rect 6217 19901 6247 19957
rect 6303 19901 6333 19957
rect 6389 19901 6419 19957
rect 6475 19901 6489 19957
rect 5889 19877 6489 19901
rect 5889 19821 5903 19877
rect 5959 19821 5989 19877
rect 6045 19821 6075 19877
rect 6131 19821 6161 19877
rect 6217 19821 6247 19877
rect 6303 19821 6333 19877
rect 6389 19821 6419 19877
rect 6475 19821 6489 19877
rect 5889 19797 6489 19821
rect 5889 19741 5903 19797
rect 5959 19741 5989 19797
rect 6045 19741 6075 19797
rect 6131 19741 6161 19797
rect 6217 19741 6247 19797
rect 6303 19741 6333 19797
rect 6389 19741 6419 19797
rect 6475 19741 6489 19797
rect 5889 19717 6489 19741
rect 5889 19661 5903 19717
rect 5959 19661 5989 19717
rect 6045 19661 6075 19717
rect 6131 19661 6161 19717
rect 6217 19661 6247 19717
rect 6303 19661 6333 19717
rect 6389 19661 6419 19717
rect 6475 19661 6489 19717
rect 5889 19637 6489 19661
rect 5889 19581 5903 19637
rect 5959 19581 5989 19637
rect 6045 19581 6075 19637
rect 6131 19581 6161 19637
rect 6217 19581 6247 19637
rect 6303 19581 6333 19637
rect 6389 19581 6419 19637
rect 6475 19581 6489 19637
rect 5889 19557 6489 19581
rect 5889 19501 5903 19557
rect 5959 19501 5989 19557
rect 6045 19501 6075 19557
rect 6131 19501 6161 19557
rect 6217 19501 6247 19557
rect 6303 19501 6333 19557
rect 6389 19501 6419 19557
rect 6475 19501 6489 19557
rect 5889 19477 6489 19501
rect 5889 19421 5903 19477
rect 5959 19421 5989 19477
rect 6045 19421 6075 19477
rect 6131 19421 6161 19477
rect 6217 19421 6247 19477
rect 6303 19421 6333 19477
rect 6389 19421 6419 19477
rect 6475 19421 6489 19477
rect 5889 19397 6489 19421
rect 5889 19341 5903 19397
rect 5959 19341 5989 19397
rect 6045 19341 6075 19397
rect 6131 19341 6161 19397
rect 6217 19341 6247 19397
rect 6303 19341 6333 19397
rect 6389 19341 6419 19397
rect 6475 19341 6489 19397
rect 5889 19317 6489 19341
rect 5889 19261 5903 19317
rect 5959 19261 5989 19317
rect 6045 19261 6075 19317
rect 6131 19261 6161 19317
rect 6217 19261 6247 19317
rect 6303 19261 6333 19317
rect 6389 19261 6419 19317
rect 6475 19261 6489 19317
rect 5889 10236 6489 19261
rect 5889 10172 5918 10236
rect 5982 10172 5998 10236
rect 6062 10172 6078 10236
rect 6142 10172 6158 10236
rect 6222 10172 6238 10236
rect 6302 10172 6318 10236
rect 6382 10172 6398 10236
rect 6462 10172 6489 10236
rect 5889 10141 6489 10172
rect 5889 10077 5918 10141
rect 5982 10077 5998 10141
rect 6062 10077 6078 10141
rect 6142 10077 6158 10141
rect 6222 10077 6238 10141
rect 6302 10077 6318 10141
rect 6382 10077 6398 10141
rect 6462 10077 6489 10141
rect 5889 10045 6489 10077
rect 5889 9981 5918 10045
rect 5982 9981 5998 10045
rect 6062 9981 6078 10045
rect 6142 9981 6158 10045
rect 6222 9981 6238 10045
rect 6302 9981 6318 10045
rect 6382 9981 6398 10045
rect 6462 9981 6489 10045
rect 5889 9949 6489 9981
rect 5889 9885 5918 9949
rect 5982 9885 5998 9949
rect 6062 9885 6078 9949
rect 6142 9885 6158 9949
rect 6222 9885 6238 9949
rect 6302 9885 6318 9949
rect 6382 9885 6398 9949
rect 6462 9885 6489 9949
rect 5889 9853 6489 9885
rect 5889 9789 5918 9853
rect 5982 9789 5998 9853
rect 6062 9789 6078 9853
rect 6142 9789 6158 9853
rect 6222 9789 6238 9853
rect 6302 9789 6318 9853
rect 6382 9789 6398 9853
rect 6462 9789 6489 9853
rect 5889 9757 6489 9789
rect 5889 9693 5918 9757
rect 5982 9693 5998 9757
rect 6062 9693 6078 9757
rect 6142 9693 6158 9757
rect 6222 9693 6238 9757
rect 6302 9693 6318 9757
rect 6382 9693 6398 9757
rect 6462 9693 6489 9757
rect 5889 9547 6489 9693
rect 6589 17767 6655 24279
rect 6589 17711 6594 17767
rect 6650 17711 6655 17767
rect 6589 17680 6655 17711
rect 6589 17624 6594 17680
rect 6650 17624 6655 17680
rect 6589 17593 6655 17624
rect 6589 17537 6594 17593
rect 6650 17537 6655 17593
rect 6589 17505 6655 17537
rect 6589 17449 6594 17505
rect 6650 17449 6655 17505
rect 6589 17417 6655 17449
rect 6589 17361 6594 17417
rect 6650 17361 6655 17417
rect 6589 17329 6655 17361
rect 6589 17273 6594 17329
rect 6650 17273 6655 17329
rect 6589 17241 6655 17273
rect 6589 17185 6594 17241
rect 6650 17185 6655 17241
rect 6589 9547 6655 17185
rect 6802 17767 6868 28533
rect 6802 17711 6807 17767
rect 6863 17711 6868 17767
rect 6802 17680 6868 17711
rect 6802 17624 6807 17680
rect 6863 17624 6868 17680
rect 6802 17593 6868 17624
rect 6802 17537 6807 17593
rect 6863 17537 6868 17593
rect 6802 17505 6868 17537
rect 6802 17449 6807 17505
rect 6863 17449 6868 17505
rect 6802 17417 6868 17449
rect 6802 17361 6807 17417
rect 6863 17361 6868 17417
rect 6802 17329 6868 17361
rect 6802 17273 6807 17329
rect 6863 17273 6868 17329
rect 6802 17241 6868 17273
rect 6802 17185 6807 17241
rect 6863 17185 6868 17241
rect 6802 9547 6868 17185
rect 6968 11200 7568 28627
rect 6968 11136 6993 11200
rect 7057 11136 7073 11200
rect 7137 11136 7153 11200
rect 7217 11136 7233 11200
rect 7297 11136 7313 11200
rect 7377 11136 7393 11200
rect 7457 11136 7473 11200
rect 7537 11136 7568 11200
rect 6968 11105 7568 11136
rect 6968 11041 6993 11105
rect 7057 11041 7073 11105
rect 7137 11041 7153 11105
rect 7217 11041 7233 11105
rect 7297 11041 7313 11105
rect 7377 11041 7393 11105
rect 7457 11041 7473 11105
rect 7537 11041 7568 11105
rect 6968 11009 7568 11041
rect 6968 10945 6993 11009
rect 7057 10945 7073 11009
rect 7137 10945 7153 11009
rect 7217 10945 7233 11009
rect 7297 10945 7313 11009
rect 7377 10945 7393 11009
rect 7457 10945 7473 11009
rect 7537 10945 7568 11009
rect 6968 10913 7568 10945
rect 6968 10849 6993 10913
rect 7057 10849 7073 10913
rect 7137 10849 7153 10913
rect 7217 10849 7233 10913
rect 7297 10849 7313 10913
rect 7377 10849 7393 10913
rect 7457 10849 7473 10913
rect 7537 10849 7568 10913
rect 6968 10817 7568 10849
rect 6968 10753 6993 10817
rect 7057 10753 7073 10817
rect 7137 10753 7153 10817
rect 7217 10753 7233 10817
rect 7297 10753 7313 10817
rect 7377 10753 7393 10817
rect 7457 10753 7473 10817
rect 7537 10753 7568 10817
rect 6968 10721 7568 10753
rect 6968 10657 6993 10721
rect 7057 10657 7073 10721
rect 7137 10657 7153 10721
rect 7217 10657 7233 10721
rect 7297 10657 7313 10721
rect 7377 10657 7393 10721
rect 7457 10657 7473 10721
rect 7537 10657 7568 10721
rect 6968 9547 7568 10657
rect 7668 17767 7734 28905
rect 7668 17711 7673 17767
rect 7729 17711 7734 17767
rect 7668 17680 7734 17711
rect 7668 17624 7673 17680
rect 7729 17624 7734 17680
rect 7668 17593 7734 17624
rect 7668 17537 7673 17593
rect 7729 17537 7734 17593
rect 7668 17505 7734 17537
rect 7668 17449 7673 17505
rect 7729 17449 7734 17505
rect 7668 17417 7734 17449
rect 7668 17361 7673 17417
rect 7729 17361 7734 17417
rect 7668 17329 7734 17361
rect 7668 17273 7673 17329
rect 7729 17273 7734 17329
rect 7668 17241 7734 17273
rect 7668 17185 7673 17241
rect 7729 17185 7734 17241
rect 7668 9547 7734 17185
rect 7834 17745 8434 28954
rect 7834 17689 7843 17745
rect 7899 17689 7949 17745
rect 8005 17689 8054 17745
rect 8110 17689 8159 17745
rect 8215 17689 8264 17745
rect 8320 17689 8369 17745
rect 8425 17689 8434 17745
rect 7834 17645 8434 17689
rect 7834 17589 7843 17645
rect 7899 17589 7949 17645
rect 8005 17589 8054 17645
rect 8110 17589 8159 17645
rect 8215 17589 8264 17645
rect 8320 17589 8369 17645
rect 8425 17589 8434 17645
rect 7834 17545 8434 17589
rect 7834 17489 7843 17545
rect 7899 17489 7949 17545
rect 8005 17489 8054 17545
rect 8110 17489 8159 17545
rect 8215 17489 8264 17545
rect 8320 17489 8369 17545
rect 8425 17489 8434 17545
rect 7834 17445 8434 17489
rect 7834 17389 7843 17445
rect 7899 17389 7949 17445
rect 8005 17389 8054 17445
rect 8110 17389 8159 17445
rect 8215 17389 8264 17445
rect 8320 17389 8369 17445
rect 8425 17389 8434 17445
rect 7834 17345 8434 17389
rect 7834 17289 7843 17345
rect 7899 17289 7949 17345
rect 8005 17289 8054 17345
rect 8110 17289 8159 17345
rect 8215 17289 8264 17345
rect 8320 17289 8369 17345
rect 8425 17289 8434 17345
rect 7834 17245 8434 17289
rect 7834 17189 7843 17245
rect 7899 17189 7949 17245
rect 8005 17189 8054 17245
rect 8110 17189 8159 17245
rect 8215 17189 8264 17245
rect 8320 17189 8369 17245
rect 8425 17189 8434 17245
rect 7834 15879 8434 17189
rect 7834 15823 7843 15879
rect 7899 15823 7949 15879
rect 8005 15823 8054 15879
rect 8110 15823 8159 15879
rect 8215 15823 8264 15879
rect 8320 15823 8369 15879
rect 8425 15823 8434 15879
rect 7834 15735 8434 15823
rect 7834 15679 7843 15735
rect 7899 15679 7949 15735
rect 8005 15679 8054 15735
rect 8110 15679 8159 15735
rect 8215 15679 8264 15735
rect 8320 15679 8369 15735
rect 8425 15679 8434 15735
rect 7834 14160 8434 15679
rect 7834 14104 7843 14160
rect 7899 14104 7949 14160
rect 8005 14104 8054 14160
rect 8110 14104 8159 14160
rect 8215 14104 8264 14160
rect 8320 14104 8369 14160
rect 8425 14104 8434 14160
rect 7834 14016 8434 14104
rect 7834 13960 7843 14016
rect 7899 13960 7949 14016
rect 8005 13960 8054 14016
rect 8110 13960 8159 14016
rect 8215 13960 8264 14016
rect 8320 13960 8369 14016
rect 8425 13960 8434 14016
rect 7834 13438 8434 13960
rect 7834 13382 7843 13438
rect 7899 13382 7949 13438
rect 8005 13382 8054 13438
rect 8110 13382 8159 13438
rect 8215 13382 8264 13438
rect 8320 13382 8369 13438
rect 8425 13382 8434 13438
rect 7834 13294 8434 13382
rect 7834 13238 7843 13294
rect 7899 13238 7949 13294
rect 8005 13238 8054 13294
rect 8110 13238 8159 13294
rect 8215 13238 8264 13294
rect 8320 13238 8369 13294
rect 8425 13238 8434 13294
rect 7834 11639 8434 13238
rect 7834 11583 7843 11639
rect 7899 11583 7949 11639
rect 8005 11583 8054 11639
rect 8110 11583 8159 11639
rect 8215 11583 8264 11639
rect 8320 11583 8369 11639
rect 8425 11583 8434 11639
rect 7834 11495 8434 11583
rect 7834 11439 7843 11495
rect 7899 11439 7949 11495
rect 8005 11439 8054 11495
rect 8110 11439 8159 11495
rect 8215 11439 8264 11495
rect 8320 11439 8369 11495
rect 8425 11439 8434 11495
rect 7834 10951 8434 11439
rect 7834 10895 7843 10951
rect 7899 10895 7949 10951
rect 8005 10895 8054 10951
rect 8110 10895 8159 10951
rect 8215 10895 8264 10951
rect 8320 10895 8369 10951
rect 8425 10895 8434 10951
rect 7834 10807 8434 10895
rect 7834 10751 7843 10807
rect 7899 10751 7949 10807
rect 8005 10751 8054 10807
rect 8110 10751 8159 10807
rect 8215 10751 8264 10807
rect 8320 10751 8369 10807
rect 8425 10751 8434 10807
rect 4416 9333 4425 9389
rect 4481 9333 4551 9389
rect 4607 9333 4616 9389
rect 4416 9309 4616 9333
rect 4416 9253 4425 9309
rect 4481 9253 4551 9309
rect 4607 9253 4616 9309
rect 2078 9241 2488 9247
rect 2078 9177 2083 9241
rect 2147 9177 2195 9241
rect 2259 9177 2307 9241
rect 2371 9177 2419 9241
rect 2483 9177 2488 9241
rect 2078 9109 2488 9177
rect 2078 9045 2083 9109
rect 2147 9045 2195 9109
rect 2259 9045 2307 9109
rect 2371 9045 2419 9109
rect 2483 9045 2488 9109
rect 2078 8977 2488 9045
rect 2078 8913 2083 8977
rect 2147 8913 2195 8977
rect 2259 8913 2307 8977
rect 2371 8913 2419 8977
rect 2483 8913 2488 8977
rect 2078 8845 2488 8913
rect 2078 8781 2083 8845
rect 2147 8781 2195 8845
rect 2259 8781 2307 8845
rect 2371 8781 2419 8845
rect 2483 8781 2488 8845
rect 2078 8775 2488 8781
rect 954 7754 963 7810
rect 1019 7754 1069 7810
rect 1125 7754 1174 7810
rect 1230 7754 1279 7810
rect 1335 7754 1384 7810
rect 1440 7754 1489 7810
rect 1545 7754 1554 7810
rect 954 7666 1554 7754
rect 954 7610 963 7666
rect 1019 7610 1069 7666
rect 1125 7610 1174 7666
rect 1230 7610 1279 7666
rect 1335 7610 1384 7666
rect 1440 7610 1489 7666
rect 1545 7610 1554 7666
rect 954 3666 1554 7610
rect 954 3602 975 3666
rect 1039 3602 1057 3666
rect 1121 3602 1139 3666
rect 1203 3602 1221 3666
rect 1285 3602 1303 3666
rect 1367 3602 1385 3666
rect 1449 3602 1467 3666
rect 1531 3602 1554 3666
rect 954 3581 1554 3602
rect 954 3517 975 3581
rect 1039 3517 1057 3581
rect 1121 3517 1139 3581
rect 1203 3517 1221 3581
rect 1285 3517 1303 3581
rect 1367 3517 1385 3581
rect 1449 3517 1467 3581
rect 1531 3517 1554 3581
rect 954 3495 1554 3517
rect 954 3431 975 3495
rect 1039 3431 1057 3495
rect 1121 3431 1139 3495
rect 1203 3431 1221 3495
rect 1285 3431 1303 3495
rect 1367 3431 1385 3495
rect 1449 3431 1467 3495
rect 1531 3431 1554 3495
rect 954 3409 1554 3431
rect 954 3345 975 3409
rect 1039 3345 1057 3409
rect 1121 3345 1139 3409
rect 1203 3345 1221 3409
rect 1285 3345 1303 3409
rect 1367 3345 1385 3409
rect 1449 3345 1467 3409
rect 1531 3345 1554 3409
rect 954 3323 1554 3345
rect 954 3317 975 3323
rect 954 3261 963 3317
rect 954 3259 975 3261
rect 1039 3259 1057 3323
rect 1121 3317 1139 3323
rect 1203 3317 1221 3323
rect 1285 3317 1303 3323
rect 1367 3317 1385 3323
rect 1125 3261 1139 3317
rect 1367 3261 1384 3317
rect 1121 3259 1139 3261
rect 1203 3259 1221 3261
rect 1285 3259 1303 3261
rect 1367 3259 1385 3261
rect 1449 3259 1467 3323
rect 1531 3317 1554 3323
rect 1545 3261 1554 3317
rect 1531 3259 1554 3261
rect 954 3237 1554 3259
rect 954 3173 975 3237
rect 1039 3173 1057 3237
rect 1121 3173 1139 3237
rect 1203 3173 1221 3237
rect 1285 3173 1303 3237
rect 1367 3173 1385 3237
rect 1449 3173 1467 3237
rect 1531 3173 1554 3237
rect 954 3117 963 3173
rect 1019 3151 1069 3173
rect 1125 3151 1174 3173
rect 1230 3151 1279 3173
rect 1335 3151 1384 3173
rect 1440 3151 1489 3173
rect 954 3087 975 3117
rect 1039 3087 1057 3151
rect 1125 3117 1139 3151
rect 1367 3117 1384 3151
rect 1121 3087 1139 3117
rect 1203 3087 1221 3117
rect 1285 3087 1303 3117
rect 1367 3087 1385 3117
rect 1449 3087 1467 3151
rect 1545 3117 1554 3173
rect 1531 3087 1554 3117
rect 954 3065 1554 3087
rect 954 3001 975 3065
rect 1039 3001 1057 3065
rect 1121 3001 1139 3065
rect 1203 3001 1221 3065
rect 1285 3001 1303 3065
rect 1367 3001 1385 3065
rect 1449 3001 1467 3065
rect 1531 3001 1554 3065
rect 954 2189 1554 3001
rect 954 2133 963 2189
rect 1019 2133 1069 2189
rect 1125 2133 1174 2189
rect 1230 2133 1279 2189
rect 1335 2133 1384 2189
rect 1440 2133 1489 2189
rect 1545 2133 1554 2189
rect 954 2067 1554 2133
rect 954 2011 963 2067
rect 1019 2011 1069 2067
rect 1125 2011 1174 2067
rect 1230 2011 1279 2067
rect 1335 2011 1384 2067
rect 1440 2011 1489 2067
rect 1545 2011 1554 2067
rect 954 1945 1554 2011
rect 954 1889 963 1945
rect 1019 1889 1069 1945
rect 1125 1889 1174 1945
rect 1230 1889 1279 1945
rect 1335 1889 1384 1945
rect 1440 1889 1489 1945
rect 1545 1889 1554 1945
rect 954 1568 1554 1889
rect 4416 8002 4616 9253
rect 4416 7946 4425 8002
rect 4481 7946 4551 8002
rect 4607 7946 4616 8002
rect 4416 7922 4616 7946
rect 4416 7866 4425 7922
rect 4481 7866 4551 7922
rect 4607 7866 4616 7922
rect 4416 6880 4616 7866
rect 4416 6824 4425 6880
rect 4481 6824 4551 6880
rect 4607 6824 4616 6880
rect 4416 6800 4616 6824
rect 4416 6744 4425 6800
rect 4481 6744 4551 6800
rect 4607 6744 4616 6800
rect 4416 5486 4616 6744
rect 4416 5430 4425 5486
rect 4481 5430 4551 5486
rect 4607 5430 4616 5486
rect 4416 5406 4616 5430
rect 4416 5350 4425 5406
rect 4481 5350 4551 5406
rect 4607 5350 4616 5406
rect 4416 4058 4616 5350
rect 4416 4002 4425 4058
rect 4481 4002 4551 4058
rect 4607 4002 4616 4058
rect 4416 3978 4616 4002
rect 4416 3922 4425 3978
rect 4481 3922 4551 3978
rect 4607 3922 4616 3978
rect 4416 3312 4616 3922
rect 4416 3256 4452 3312
rect 4508 3256 4532 3312
rect 4588 3256 4616 3312
rect 4416 3231 4616 3256
rect 4416 3175 4452 3231
rect 4508 3175 4532 3231
rect 4588 3175 4616 3231
rect 4416 3150 4616 3175
rect 4416 3094 4452 3150
rect 4508 3094 4532 3150
rect 4588 3094 4616 3150
rect 4416 3069 4616 3094
rect 4416 3013 4452 3069
rect 4508 3013 4532 3069
rect 4588 3013 4616 3069
rect 4416 2988 4616 3013
rect 4416 2932 4452 2988
rect 4508 2932 4532 2988
rect 4588 2932 4616 2988
rect 4416 2907 4616 2932
rect 4416 2851 4452 2907
rect 4508 2851 4532 2907
rect 4588 2851 4616 2907
rect 4416 2826 4616 2851
rect 4416 2770 4452 2826
rect 4508 2770 4532 2826
rect 4588 2770 4616 2826
rect 4416 2744 4616 2770
rect 4416 2701 4452 2744
rect 4416 2637 4428 2701
rect 4508 2688 4532 2744
rect 4588 2701 4616 2744
rect 4492 2662 4538 2688
rect 4416 2616 4452 2637
rect 4416 2552 4428 2616
rect 4508 2606 4532 2662
rect 4602 2637 4616 2701
rect 4588 2616 4616 2637
rect 4492 2580 4538 2606
rect 4416 2531 4452 2552
rect 4416 2467 4428 2531
rect 4508 2524 4532 2580
rect 4602 2552 4616 2616
rect 4588 2531 4616 2552
rect 4492 2498 4538 2524
rect 4416 2446 4452 2467
rect 4416 2382 4428 2446
rect 4508 2442 4532 2498
rect 4602 2467 4616 2531
rect 4588 2446 4616 2467
rect 4492 2416 4538 2442
rect 4416 2361 4452 2382
rect 4416 2297 4428 2361
rect 4508 2360 4532 2416
rect 4602 2382 4616 2446
rect 4588 2361 4616 2382
rect 4492 2334 4538 2360
rect 4416 2278 4452 2297
rect 4508 2278 4532 2334
rect 4602 2297 4616 2361
rect 4588 2278 4616 2297
rect 4416 2276 4616 2278
rect 4416 2212 4428 2276
rect 4492 2252 4538 2276
rect 4416 2196 4452 2212
rect 4508 2196 4532 2252
rect 4602 2212 4616 2276
rect 4588 2196 4616 2212
rect 4416 2191 4616 2196
rect 4416 2127 4428 2191
rect 4492 2170 4538 2191
rect 4416 2114 4452 2127
rect 4508 2114 4532 2170
rect 4602 2127 4616 2191
rect 4588 2114 4616 2127
rect 4416 2105 4616 2114
rect 4416 2041 4428 2105
rect 4492 2088 4538 2105
rect 4416 2032 4452 2041
rect 4508 2032 4532 2088
rect 4602 2041 4616 2105
rect 4588 2032 4616 2041
rect 4416 2019 4616 2032
rect 4416 1955 4428 2019
rect 4492 2006 4538 2019
rect 4416 1950 4452 1955
rect 4508 1950 4532 2006
rect 4602 1955 4616 2019
rect 4588 1950 4616 1955
rect 4416 1933 4616 1950
rect 4416 1869 4428 1933
rect 4492 1924 4538 1933
rect 4416 1868 4452 1869
rect 4508 1868 4532 1924
rect 4602 1869 4616 1933
rect 4588 1868 4616 1869
rect 4416 1847 4616 1868
rect 4416 1783 4428 1847
rect 4492 1842 4538 1847
rect 4508 1786 4532 1842
rect 4492 1783 4538 1786
rect 4602 1783 4616 1847
rect 4416 1777 4616 1783
rect 7834 9205 8434 10751
rect 7834 9149 7843 9205
rect 7899 9149 7949 9205
rect 8005 9149 8054 9205
rect 8110 9149 8159 9205
rect 8215 9149 8264 9205
rect 8320 9149 8369 9205
rect 8425 9149 8434 9205
rect 7834 9061 8434 9149
rect 7834 9005 7843 9061
rect 7899 9005 7949 9061
rect 8005 9005 8054 9061
rect 8110 9005 8159 9061
rect 8215 9005 8264 9061
rect 8320 9005 8369 9061
rect 8425 9005 8434 9061
rect 7834 8436 8434 9005
rect 7834 8380 7843 8436
rect 7899 8380 7949 8436
rect 8005 8380 8054 8436
rect 8110 8380 8159 8436
rect 8215 8380 8264 8436
rect 8320 8380 8369 8436
rect 8425 8380 8434 8436
rect 7834 8292 8434 8380
rect 8527 9238 9233 9247
rect 8527 9182 8532 9238
rect 8588 9236 8612 9238
rect 8668 9236 8692 9238
rect 8748 9236 8772 9238
rect 8828 9236 8852 9238
rect 8908 9236 8932 9238
rect 8988 9236 9012 9238
rect 9068 9236 9092 9238
rect 9148 9236 9172 9238
rect 9228 9182 9233 9238
rect 8527 9172 8568 9182
rect 8632 9172 8648 9182
rect 8712 9172 8728 9182
rect 8792 9172 8808 9182
rect 8872 9172 8888 9182
rect 8952 9172 8968 9182
rect 9032 9172 9048 9182
rect 9112 9172 9128 9182
rect 9192 9172 9233 9182
rect 8527 9153 9233 9172
rect 8527 9097 8532 9153
rect 9228 9097 9233 9153
rect 8527 9089 8568 9097
rect 8632 9089 8648 9097
rect 8712 9089 8728 9097
rect 8792 9089 8808 9097
rect 8872 9089 8888 9097
rect 8952 9089 8968 9097
rect 9032 9089 9048 9097
rect 9112 9089 9128 9097
rect 9192 9089 9233 9097
rect 8527 9070 9233 9089
rect 8527 9068 8568 9070
rect 8632 9068 8648 9070
rect 8712 9068 8728 9070
rect 8792 9068 8808 9070
rect 8872 9068 8888 9070
rect 8952 9068 8968 9070
rect 9032 9068 9048 9070
rect 9112 9068 9128 9070
rect 9192 9068 9233 9070
rect 8527 9012 8532 9068
rect 9228 9012 9233 9068
rect 8527 9006 8568 9012
rect 8632 9006 8648 9012
rect 8712 9006 8728 9012
rect 8792 9006 8808 9012
rect 8872 9006 8888 9012
rect 8952 9006 8968 9012
rect 9032 9006 9048 9012
rect 9112 9006 9128 9012
rect 9192 9006 9233 9012
rect 8527 8986 9233 9006
rect 8527 8983 8568 8986
rect 8632 8983 8648 8986
rect 8712 8983 8728 8986
rect 8792 8983 8808 8986
rect 8872 8983 8888 8986
rect 8952 8983 8968 8986
rect 9032 8983 9048 8986
rect 9112 8983 9128 8986
rect 9192 8983 9233 8986
rect 8527 8927 8532 8983
rect 9228 8927 9233 8983
rect 8527 8922 8568 8927
rect 8632 8922 8648 8927
rect 8712 8922 8728 8927
rect 8792 8922 8808 8927
rect 8872 8922 8888 8927
rect 8952 8922 8968 8927
rect 9032 8922 9048 8927
rect 9112 8922 9128 8927
rect 9192 8922 9233 8927
rect 8527 8902 9233 8922
rect 8527 8898 8568 8902
rect 8632 8898 8648 8902
rect 8712 8898 8728 8902
rect 8792 8898 8808 8902
rect 8872 8898 8888 8902
rect 8952 8898 8968 8902
rect 9032 8898 9048 8902
rect 9112 8898 9128 8902
rect 9192 8898 9233 8902
rect 8527 8842 8532 8898
rect 9228 8842 9233 8898
rect 8527 8838 8568 8842
rect 8632 8838 8648 8842
rect 8712 8838 8728 8842
rect 8792 8838 8808 8842
rect 8872 8838 8888 8842
rect 8952 8838 8968 8842
rect 9032 8838 9048 8842
rect 9112 8838 9128 8842
rect 9192 8838 9233 8842
rect 8527 8818 9233 8838
rect 8527 8812 8568 8818
rect 8632 8812 8648 8818
rect 8712 8812 8728 8818
rect 8792 8812 8808 8818
rect 8872 8812 8888 8818
rect 8952 8812 8968 8818
rect 9032 8812 9048 8818
rect 9112 8812 9128 8818
rect 9192 8812 9233 8818
rect 8527 8756 8532 8812
rect 9228 8756 9233 8812
rect 8527 8754 8568 8756
rect 8632 8754 8648 8756
rect 8712 8754 8728 8756
rect 8792 8754 8808 8756
rect 8872 8754 8888 8756
rect 8952 8754 8968 8756
rect 9032 8754 9048 8756
rect 9112 8754 9128 8756
rect 9192 8754 9233 8756
rect 8527 8734 9233 8754
rect 8527 8726 8568 8734
rect 8632 8726 8648 8734
rect 8712 8726 8728 8734
rect 8792 8726 8808 8734
rect 8872 8726 8888 8734
rect 8952 8726 8968 8734
rect 9032 8726 9048 8734
rect 9112 8726 9128 8734
rect 9192 8726 9233 8734
rect 8527 8670 8532 8726
rect 9228 8670 9233 8726
rect 8527 8650 9233 8670
rect 8527 8640 8568 8650
rect 8632 8640 8648 8650
rect 8712 8640 8728 8650
rect 8792 8640 8808 8650
rect 8872 8640 8888 8650
rect 8952 8640 8968 8650
rect 9032 8640 9048 8650
rect 9112 8640 9128 8650
rect 9192 8640 9233 8650
rect 8527 8584 8532 8640
rect 8588 8584 8612 8586
rect 8668 8584 8692 8586
rect 8748 8584 8772 8586
rect 8828 8584 8852 8586
rect 8908 8584 8932 8586
rect 8988 8584 9012 8586
rect 9068 8584 9092 8586
rect 9148 8584 9172 8586
rect 9228 8584 9233 8640
rect 8527 8566 9233 8584
rect 8527 8554 8568 8566
rect 8632 8554 8648 8566
rect 8712 8554 8728 8566
rect 8792 8554 8808 8566
rect 8872 8554 8888 8566
rect 8952 8554 8968 8566
rect 9032 8554 9048 8566
rect 9112 8554 9128 8566
rect 9192 8554 9233 8566
rect 8527 8498 8532 8554
rect 8588 8498 8612 8502
rect 8668 8498 8692 8502
rect 8748 8498 8772 8502
rect 8828 8498 8852 8502
rect 8908 8498 8932 8502
rect 8988 8498 9012 8502
rect 9068 8498 9092 8502
rect 9148 8498 9172 8502
rect 9228 8498 9233 8554
rect 8527 8482 9233 8498
rect 8527 8468 8568 8482
rect 8632 8468 8648 8482
rect 8712 8468 8728 8482
rect 8792 8468 8808 8482
rect 8872 8468 8888 8482
rect 8952 8468 8968 8482
rect 9032 8468 9048 8482
rect 9112 8468 9128 8482
rect 9192 8468 9233 8482
rect 8527 8412 8532 8468
rect 8588 8412 8612 8418
rect 8668 8412 8692 8418
rect 8748 8412 8772 8418
rect 8828 8412 8852 8418
rect 8908 8412 8932 8418
rect 8988 8412 9012 8418
rect 9068 8412 9092 8418
rect 9148 8412 9172 8418
rect 9228 8412 9233 8468
rect 8527 8398 9233 8412
rect 8527 8382 8568 8398
rect 8632 8382 8648 8398
rect 8712 8382 8728 8398
rect 8792 8382 8808 8398
rect 8872 8382 8888 8398
rect 8952 8382 8968 8398
rect 9032 8382 9048 8398
rect 9112 8382 9128 8398
rect 9192 8382 9233 8398
rect 8527 8326 8532 8382
rect 8588 8326 8612 8334
rect 8668 8326 8692 8334
rect 8748 8326 8772 8334
rect 8828 8326 8852 8334
rect 8908 8326 8932 8334
rect 8988 8326 9012 8334
rect 9068 8326 9092 8334
rect 9148 8326 9172 8334
rect 9228 8326 9233 8382
rect 8527 8317 9233 8326
rect 7834 8236 7843 8292
rect 7899 8236 7949 8292
rect 8005 8236 8054 8292
rect 8110 8236 8159 8292
rect 8215 8236 8264 8292
rect 8320 8236 8369 8292
rect 8425 8236 8434 8292
rect 7834 8031 8434 8236
rect 7834 7967 7865 8031
rect 7929 7967 7945 8031
rect 8009 7967 8025 8031
rect 8089 7967 8105 8031
rect 8169 7967 8185 8031
rect 8249 7967 8265 8031
rect 8329 7967 8345 8031
rect 8409 7967 8434 8031
rect 7834 7944 8434 7967
rect 7834 7880 7865 7944
rect 7929 7880 7945 7944
rect 8009 7880 8025 7944
rect 8089 7880 8105 7944
rect 8169 7880 8185 7944
rect 8249 7880 8265 7944
rect 8329 7880 8345 7944
rect 8409 7880 8434 7944
rect 7834 7857 8434 7880
rect 7834 7793 7865 7857
rect 7929 7793 7945 7857
rect 8009 7793 8025 7857
rect 8089 7793 8105 7857
rect 8169 7793 8185 7857
rect 8249 7793 8265 7857
rect 8329 7793 8345 7857
rect 8409 7793 8434 7857
rect 7834 7769 8434 7793
rect 7834 7705 7865 7769
rect 7929 7705 7945 7769
rect 8009 7705 8025 7769
rect 8089 7705 8105 7769
rect 8169 7705 8185 7769
rect 8249 7705 8265 7769
rect 8329 7705 8345 7769
rect 8409 7705 8434 7769
rect 7834 7681 8434 7705
rect 7834 7617 7865 7681
rect 7929 7617 7945 7681
rect 8009 7617 8025 7681
rect 8089 7617 8105 7681
rect 8169 7617 8185 7681
rect 8249 7617 8265 7681
rect 8329 7617 8345 7681
rect 8409 7617 8434 7681
rect 7834 7593 8434 7617
rect 7834 7529 7865 7593
rect 7929 7529 7945 7593
rect 8009 7529 8025 7593
rect 8089 7529 8105 7593
rect 8169 7529 8185 7593
rect 8249 7529 8265 7593
rect 8329 7529 8345 7593
rect 8409 7529 8434 7593
rect 7834 7505 8434 7529
rect 7834 7441 7865 7505
rect 7929 7441 7945 7505
rect 8009 7441 8025 7505
rect 8089 7441 8105 7505
rect 8169 7441 8185 7505
rect 8249 7441 8265 7505
rect 8329 7441 8345 7505
rect 8409 7441 8434 7505
rect 7834 7417 8434 7441
rect 7834 7353 7865 7417
rect 7929 7353 7945 7417
rect 8009 7353 8025 7417
rect 8089 7353 8105 7417
rect 8169 7353 8185 7417
rect 8249 7353 8265 7417
rect 8329 7353 8345 7417
rect 8409 7353 8434 7417
rect 7834 6704 8434 7353
rect 7834 6648 7843 6704
rect 7899 6648 7949 6704
rect 8005 6648 8054 6704
rect 8110 6648 8159 6704
rect 8215 6648 8264 6704
rect 8320 6648 8369 6704
rect 8425 6648 8434 6704
rect 7834 6560 8434 6648
rect 7834 6504 7843 6560
rect 7899 6504 7949 6560
rect 8005 6504 8054 6560
rect 8110 6504 8159 6560
rect 8215 6504 8264 6560
rect 8320 6504 8369 6560
rect 8425 6504 8434 6560
rect 7834 5917 8434 6504
rect 7834 5861 7843 5917
rect 7899 5861 7949 5917
rect 8005 5861 8054 5917
rect 8110 5861 8159 5917
rect 8215 5861 8264 5917
rect 8320 5861 8369 5917
rect 8425 5861 8434 5917
rect 7834 5773 8434 5861
rect 7834 5717 7843 5773
rect 7899 5717 7949 5773
rect 8005 5717 8054 5773
rect 8110 5717 8159 5773
rect 8215 5717 8264 5773
rect 8320 5717 8369 5773
rect 8425 5717 8434 5773
rect 7834 4868 8434 5717
rect 7834 4812 7843 4868
rect 7899 4812 7949 4868
rect 8005 4812 8054 4868
rect 8110 4812 8159 4868
rect 8215 4812 8264 4868
rect 8320 4812 8369 4868
rect 8425 4812 8434 4868
rect 7834 4724 8434 4812
rect 7834 4668 7843 4724
rect 7899 4668 7949 4724
rect 8005 4668 8054 4724
rect 8110 4668 8159 4724
rect 8215 4668 8264 4724
rect 8320 4668 8369 4724
rect 8425 4668 8434 4724
rect 7834 3732 8434 4668
rect 7834 3676 7843 3732
rect 7899 3676 7949 3732
rect 8005 3676 8054 3732
rect 8110 3676 8159 3732
rect 8215 3676 8264 3732
rect 8320 3676 8369 3732
rect 8425 3676 8434 3732
rect 7834 3588 8434 3676
rect 7834 3532 7843 3588
rect 7899 3532 7949 3588
rect 8005 3532 8054 3588
rect 8110 3532 8159 3588
rect 8215 3532 8264 3588
rect 8320 3532 8369 3588
rect 8425 3532 8434 3588
rect 7834 3222 8434 3532
rect 7834 3166 7843 3222
rect 7899 3166 7949 3222
rect 8005 3166 8054 3222
rect 8110 3166 8159 3222
rect 8215 3166 8264 3222
rect 8320 3166 8369 3222
rect 8425 3166 8434 3222
rect 7834 3078 8434 3166
rect 7834 3022 7843 3078
rect 7899 3022 7949 3078
rect 8005 3022 8054 3078
rect 8110 3022 8159 3078
rect 8215 3022 8264 3078
rect 8320 3022 8369 3078
rect 8425 3022 8434 3078
rect 7834 1597 8434 3022
<< via3 >>
rect 316 9238 380 9241
rect 316 9182 320 9238
rect 320 9182 376 9238
rect 376 9182 380 9238
rect 316 9177 380 9182
rect 316 9153 380 9156
rect 316 9097 320 9153
rect 320 9097 376 9153
rect 376 9097 380 9153
rect 316 9092 380 9097
rect 316 9068 380 9071
rect 316 9012 320 9068
rect 320 9012 376 9068
rect 376 9012 380 9068
rect 316 9007 380 9012
rect 316 8983 380 8986
rect 316 8927 320 8983
rect 320 8927 376 8983
rect 376 8927 380 8983
rect 316 8922 380 8927
rect 316 8898 380 8901
rect 316 8842 320 8898
rect 320 8842 376 8898
rect 376 8842 380 8898
rect 316 8837 380 8842
rect 316 8812 380 8816
rect 316 8756 320 8812
rect 320 8756 376 8812
rect 376 8756 380 8812
rect 316 8752 380 8756
rect 316 8726 380 8731
rect 316 8670 320 8726
rect 320 8670 376 8726
rect 376 8670 380 8726
rect 316 8667 380 8670
rect 316 8640 380 8645
rect 316 8584 320 8640
rect 320 8584 376 8640
rect 376 8584 380 8640
rect 316 8581 380 8584
rect 316 8554 380 8559
rect 316 8498 320 8554
rect 320 8498 376 8554
rect 376 8498 380 8554
rect 316 8495 380 8498
rect 316 8468 380 8473
rect 316 8412 320 8468
rect 320 8412 376 8468
rect 376 8412 380 8468
rect 316 8409 380 8412
rect 316 8382 380 8387
rect 316 8326 320 8382
rect 320 8326 376 8382
rect 376 8326 380 8382
rect 316 8323 380 8326
rect 490 6977 554 7041
rect 580 6977 644 7041
rect 670 6977 734 7041
rect 760 6977 824 7041
rect 490 6896 554 6960
rect 580 6896 644 6960
rect 670 6896 734 6960
rect 760 6896 824 6960
rect 490 6814 554 6878
rect 580 6814 644 6878
rect 670 6814 734 6878
rect 760 6814 824 6878
rect 490 6732 554 6796
rect 580 6732 644 6796
rect 670 6732 734 6796
rect 760 6732 824 6796
rect 490 6650 554 6714
rect 580 6650 644 6714
rect 670 6650 734 6714
rect 760 6650 824 6714
rect 490 6568 554 6632
rect 580 6568 644 6632
rect 670 6568 734 6632
rect 760 6568 824 6632
rect 490 6486 554 6550
rect 580 6486 644 6550
rect 670 6486 734 6550
rect 760 6486 824 6550
rect 490 6404 554 6468
rect 580 6404 644 6468
rect 670 6404 734 6468
rect 760 6404 824 6468
rect 1856 11128 1920 11192
rect 1936 11128 2000 11192
rect 2016 11128 2080 11192
rect 2096 11128 2160 11192
rect 2176 11128 2240 11192
rect 2256 11128 2320 11192
rect 2336 11128 2400 11192
rect 1856 11033 1920 11097
rect 1936 11033 2000 11097
rect 2016 11033 2080 11097
rect 2096 11033 2160 11097
rect 2176 11033 2240 11097
rect 2256 11033 2320 11097
rect 2336 11033 2400 11097
rect 1856 10937 1920 11001
rect 1936 10937 2000 11001
rect 2016 10937 2080 11001
rect 2096 10937 2160 11001
rect 2176 10937 2240 11001
rect 2256 10937 2320 11001
rect 2336 10937 2400 11001
rect 1856 10841 1920 10905
rect 1936 10841 2000 10905
rect 2016 10841 2080 10905
rect 2096 10841 2160 10905
rect 2176 10841 2240 10905
rect 2256 10841 2320 10905
rect 2336 10841 2400 10905
rect 1856 10745 1920 10809
rect 1936 10745 2000 10809
rect 2016 10745 2080 10809
rect 2096 10745 2160 10809
rect 2176 10745 2240 10809
rect 2256 10745 2320 10809
rect 2336 10745 2400 10809
rect 1856 10649 1920 10713
rect 1936 10649 2000 10713
rect 2016 10649 2080 10713
rect 2096 10649 2160 10713
rect 2176 10649 2240 10713
rect 2256 10649 2320 10713
rect 2336 10649 2400 10713
rect 2921 10180 2985 10244
rect 3001 10180 3065 10244
rect 3081 10180 3145 10244
rect 3161 10180 3225 10244
rect 3241 10180 3305 10244
rect 3321 10180 3385 10244
rect 3401 10180 3465 10244
rect 2921 10085 2985 10149
rect 3001 10085 3065 10149
rect 3081 10085 3145 10149
rect 3161 10085 3225 10149
rect 3241 10085 3305 10149
rect 3321 10085 3385 10149
rect 3401 10085 3465 10149
rect 2921 9989 2985 10053
rect 3001 9989 3065 10053
rect 3081 9989 3145 10053
rect 3161 9989 3225 10053
rect 3241 9989 3305 10053
rect 3321 9989 3385 10053
rect 3401 9989 3465 10053
rect 2921 9893 2985 9957
rect 3001 9893 3065 9957
rect 3081 9893 3145 9957
rect 3161 9893 3225 9957
rect 3241 9893 3305 9957
rect 3321 9893 3385 9957
rect 3401 9893 3465 9957
rect 2921 9797 2985 9861
rect 3001 9797 3065 9861
rect 3081 9797 3145 9861
rect 3161 9797 3225 9861
rect 3241 9797 3305 9861
rect 3321 9797 3385 9861
rect 3401 9797 3465 9861
rect 2921 9701 2985 9765
rect 3001 9701 3065 9765
rect 3081 9701 3145 9765
rect 3161 9701 3225 9765
rect 3241 9701 3305 9765
rect 3321 9701 3385 9765
rect 3401 9701 3465 9765
rect 5918 10172 5982 10236
rect 5998 10172 6062 10236
rect 6078 10172 6142 10236
rect 6158 10172 6222 10236
rect 6238 10172 6302 10236
rect 6318 10172 6382 10236
rect 6398 10172 6462 10236
rect 5918 10077 5982 10141
rect 5998 10077 6062 10141
rect 6078 10077 6142 10141
rect 6158 10077 6222 10141
rect 6238 10077 6302 10141
rect 6318 10077 6382 10141
rect 6398 10077 6462 10141
rect 5918 9981 5982 10045
rect 5998 9981 6062 10045
rect 6078 9981 6142 10045
rect 6158 9981 6222 10045
rect 6238 9981 6302 10045
rect 6318 9981 6382 10045
rect 6398 9981 6462 10045
rect 5918 9885 5982 9949
rect 5998 9885 6062 9949
rect 6078 9885 6142 9949
rect 6158 9885 6222 9949
rect 6238 9885 6302 9949
rect 6318 9885 6382 9949
rect 6398 9885 6462 9949
rect 5918 9789 5982 9853
rect 5998 9789 6062 9853
rect 6078 9789 6142 9853
rect 6158 9789 6222 9853
rect 6238 9789 6302 9853
rect 6318 9789 6382 9853
rect 6398 9789 6462 9853
rect 5918 9693 5982 9757
rect 5998 9693 6062 9757
rect 6078 9693 6142 9757
rect 6158 9693 6222 9757
rect 6238 9693 6302 9757
rect 6318 9693 6382 9757
rect 6398 9693 6462 9757
rect 6993 11136 7057 11200
rect 7073 11136 7137 11200
rect 7153 11136 7217 11200
rect 7233 11136 7297 11200
rect 7313 11136 7377 11200
rect 7393 11136 7457 11200
rect 7473 11136 7537 11200
rect 6993 11041 7057 11105
rect 7073 11041 7137 11105
rect 7153 11041 7217 11105
rect 7233 11041 7297 11105
rect 7313 11041 7377 11105
rect 7393 11041 7457 11105
rect 7473 11041 7537 11105
rect 6993 10945 7057 11009
rect 7073 10945 7137 11009
rect 7153 10945 7217 11009
rect 7233 10945 7297 11009
rect 7313 10945 7377 11009
rect 7393 10945 7457 11009
rect 7473 10945 7537 11009
rect 6993 10849 7057 10913
rect 7073 10849 7137 10913
rect 7153 10849 7217 10913
rect 7233 10849 7297 10913
rect 7313 10849 7377 10913
rect 7393 10849 7457 10913
rect 7473 10849 7537 10913
rect 6993 10753 7057 10817
rect 7073 10753 7137 10817
rect 7153 10753 7217 10817
rect 7233 10753 7297 10817
rect 7313 10753 7377 10817
rect 7393 10753 7457 10817
rect 7473 10753 7537 10817
rect 6993 10657 7057 10721
rect 7073 10657 7137 10721
rect 7153 10657 7217 10721
rect 7233 10657 7297 10721
rect 7313 10657 7377 10721
rect 7393 10657 7457 10721
rect 7473 10657 7537 10721
rect 2083 9238 2147 9241
rect 2083 9182 2084 9238
rect 2084 9182 2140 9238
rect 2140 9182 2147 9238
rect 2083 9177 2147 9182
rect 2195 9238 2259 9241
rect 2195 9182 2198 9238
rect 2198 9182 2254 9238
rect 2254 9182 2259 9238
rect 2195 9177 2259 9182
rect 2307 9238 2371 9241
rect 2307 9182 2312 9238
rect 2312 9182 2368 9238
rect 2368 9182 2371 9238
rect 2307 9177 2371 9182
rect 2419 9238 2483 9241
rect 2419 9182 2426 9238
rect 2426 9182 2482 9238
rect 2482 9182 2483 9238
rect 2419 9177 2483 9182
rect 2083 9106 2147 9109
rect 2083 9050 2084 9106
rect 2084 9050 2140 9106
rect 2140 9050 2147 9106
rect 2083 9045 2147 9050
rect 2195 9106 2259 9109
rect 2195 9050 2198 9106
rect 2198 9050 2254 9106
rect 2254 9050 2259 9106
rect 2195 9045 2259 9050
rect 2307 9106 2371 9109
rect 2307 9050 2312 9106
rect 2312 9050 2368 9106
rect 2368 9050 2371 9106
rect 2307 9045 2371 9050
rect 2419 9106 2483 9109
rect 2419 9050 2426 9106
rect 2426 9050 2482 9106
rect 2482 9050 2483 9106
rect 2419 9045 2483 9050
rect 2083 8973 2147 8977
rect 2083 8917 2084 8973
rect 2084 8917 2140 8973
rect 2140 8917 2147 8973
rect 2083 8913 2147 8917
rect 2195 8973 2259 8977
rect 2195 8917 2198 8973
rect 2198 8917 2254 8973
rect 2254 8917 2259 8973
rect 2195 8913 2259 8917
rect 2307 8973 2371 8977
rect 2307 8917 2312 8973
rect 2312 8917 2368 8973
rect 2368 8917 2371 8973
rect 2307 8913 2371 8917
rect 2419 8973 2483 8977
rect 2419 8917 2426 8973
rect 2426 8917 2482 8973
rect 2482 8917 2483 8973
rect 2419 8913 2483 8917
rect 2083 8840 2147 8845
rect 2083 8784 2084 8840
rect 2084 8784 2140 8840
rect 2140 8784 2147 8840
rect 2083 8781 2147 8784
rect 2195 8840 2259 8845
rect 2195 8784 2198 8840
rect 2198 8784 2254 8840
rect 2254 8784 2259 8840
rect 2195 8781 2259 8784
rect 2307 8840 2371 8845
rect 2307 8784 2312 8840
rect 2312 8784 2368 8840
rect 2368 8784 2371 8840
rect 2307 8781 2371 8784
rect 2419 8840 2483 8845
rect 2419 8784 2426 8840
rect 2426 8784 2482 8840
rect 2482 8784 2483 8840
rect 2419 8781 2483 8784
rect 975 3602 1039 3666
rect 1057 3602 1121 3666
rect 1139 3602 1203 3666
rect 1221 3602 1285 3666
rect 1303 3602 1367 3666
rect 1385 3602 1449 3666
rect 1467 3602 1531 3666
rect 975 3517 1039 3581
rect 1057 3517 1121 3581
rect 1139 3517 1203 3581
rect 1221 3517 1285 3581
rect 1303 3517 1367 3581
rect 1385 3517 1449 3581
rect 1467 3517 1531 3581
rect 975 3431 1039 3495
rect 1057 3431 1121 3495
rect 1139 3431 1203 3495
rect 1221 3431 1285 3495
rect 1303 3431 1367 3495
rect 1385 3431 1449 3495
rect 1467 3431 1531 3495
rect 975 3345 1039 3409
rect 1057 3345 1121 3409
rect 1139 3345 1203 3409
rect 1221 3345 1285 3409
rect 1303 3345 1367 3409
rect 1385 3345 1449 3409
rect 1467 3345 1531 3409
rect 975 3317 1039 3323
rect 975 3261 1019 3317
rect 1019 3261 1039 3317
rect 975 3259 1039 3261
rect 1057 3317 1121 3323
rect 1139 3317 1203 3323
rect 1221 3317 1285 3323
rect 1303 3317 1367 3323
rect 1385 3317 1449 3323
rect 1057 3261 1069 3317
rect 1069 3261 1121 3317
rect 1139 3261 1174 3317
rect 1174 3261 1203 3317
rect 1221 3261 1230 3317
rect 1230 3261 1279 3317
rect 1279 3261 1285 3317
rect 1303 3261 1335 3317
rect 1335 3261 1367 3317
rect 1385 3261 1440 3317
rect 1440 3261 1449 3317
rect 1057 3259 1121 3261
rect 1139 3259 1203 3261
rect 1221 3259 1285 3261
rect 1303 3259 1367 3261
rect 1385 3259 1449 3261
rect 1467 3317 1531 3323
rect 1467 3261 1489 3317
rect 1489 3261 1531 3317
rect 1467 3259 1531 3261
rect 975 3173 1039 3237
rect 1057 3173 1121 3237
rect 1139 3173 1203 3237
rect 1221 3173 1285 3237
rect 1303 3173 1367 3237
rect 1385 3173 1449 3237
rect 1467 3173 1531 3237
rect 975 3117 1019 3151
rect 1019 3117 1039 3151
rect 975 3087 1039 3117
rect 1057 3117 1069 3151
rect 1069 3117 1121 3151
rect 1139 3117 1174 3151
rect 1174 3117 1203 3151
rect 1221 3117 1230 3151
rect 1230 3117 1279 3151
rect 1279 3117 1285 3151
rect 1303 3117 1335 3151
rect 1335 3117 1367 3151
rect 1385 3117 1440 3151
rect 1440 3117 1449 3151
rect 1057 3087 1121 3117
rect 1139 3087 1203 3117
rect 1221 3087 1285 3117
rect 1303 3087 1367 3117
rect 1385 3087 1449 3117
rect 1467 3117 1489 3151
rect 1489 3117 1531 3151
rect 1467 3087 1531 3117
rect 975 3001 1039 3065
rect 1057 3001 1121 3065
rect 1139 3001 1203 3065
rect 1221 3001 1285 3065
rect 1303 3001 1367 3065
rect 1385 3001 1449 3065
rect 1467 3001 1531 3065
rect 4428 2688 4452 2701
rect 4452 2688 4492 2701
rect 4538 2688 4588 2701
rect 4588 2688 4602 2701
rect 4428 2662 4492 2688
rect 4538 2662 4602 2688
rect 4428 2637 4452 2662
rect 4452 2637 4492 2662
rect 4428 2606 4452 2616
rect 4452 2606 4492 2616
rect 4538 2637 4588 2662
rect 4588 2637 4602 2662
rect 4538 2606 4588 2616
rect 4588 2606 4602 2616
rect 4428 2580 4492 2606
rect 4538 2580 4602 2606
rect 4428 2552 4452 2580
rect 4452 2552 4492 2580
rect 4428 2524 4452 2531
rect 4452 2524 4492 2531
rect 4538 2552 4588 2580
rect 4588 2552 4602 2580
rect 4538 2524 4588 2531
rect 4588 2524 4602 2531
rect 4428 2498 4492 2524
rect 4538 2498 4602 2524
rect 4428 2467 4452 2498
rect 4452 2467 4492 2498
rect 4428 2442 4452 2446
rect 4452 2442 4492 2446
rect 4538 2467 4588 2498
rect 4588 2467 4602 2498
rect 4538 2442 4588 2446
rect 4588 2442 4602 2446
rect 4428 2416 4492 2442
rect 4538 2416 4602 2442
rect 4428 2382 4452 2416
rect 4452 2382 4492 2416
rect 4428 2360 4452 2361
rect 4452 2360 4492 2361
rect 4538 2382 4588 2416
rect 4588 2382 4602 2416
rect 4538 2360 4588 2361
rect 4588 2360 4602 2361
rect 4428 2334 4492 2360
rect 4538 2334 4602 2360
rect 4428 2297 4452 2334
rect 4452 2297 4492 2334
rect 4538 2297 4588 2334
rect 4588 2297 4602 2334
rect 4428 2252 4492 2276
rect 4538 2252 4602 2276
rect 4428 2212 4452 2252
rect 4452 2212 4492 2252
rect 4538 2212 4588 2252
rect 4588 2212 4602 2252
rect 4428 2170 4492 2191
rect 4538 2170 4602 2191
rect 4428 2127 4452 2170
rect 4452 2127 4492 2170
rect 4538 2127 4588 2170
rect 4588 2127 4602 2170
rect 4428 2088 4492 2105
rect 4538 2088 4602 2105
rect 4428 2041 4452 2088
rect 4452 2041 4492 2088
rect 4538 2041 4588 2088
rect 4588 2041 4602 2088
rect 4428 2006 4492 2019
rect 4538 2006 4602 2019
rect 4428 1955 4452 2006
rect 4452 1955 4492 2006
rect 4538 1955 4588 2006
rect 4588 1955 4602 2006
rect 4428 1924 4492 1933
rect 4538 1924 4602 1933
rect 4428 1869 4452 1924
rect 4452 1869 4492 1924
rect 4538 1869 4588 1924
rect 4588 1869 4602 1924
rect 4428 1842 4492 1847
rect 4538 1842 4602 1847
rect 4428 1786 4452 1842
rect 4452 1786 4492 1842
rect 4538 1786 4588 1842
rect 4588 1786 4602 1842
rect 4428 1783 4492 1786
rect 4538 1783 4602 1786
rect 8568 9182 8588 9236
rect 8588 9182 8612 9236
rect 8612 9182 8632 9236
rect 8648 9182 8668 9236
rect 8668 9182 8692 9236
rect 8692 9182 8712 9236
rect 8728 9182 8748 9236
rect 8748 9182 8772 9236
rect 8772 9182 8792 9236
rect 8808 9182 8828 9236
rect 8828 9182 8852 9236
rect 8852 9182 8872 9236
rect 8888 9182 8908 9236
rect 8908 9182 8932 9236
rect 8932 9182 8952 9236
rect 8968 9182 8988 9236
rect 8988 9182 9012 9236
rect 9012 9182 9032 9236
rect 9048 9182 9068 9236
rect 9068 9182 9092 9236
rect 9092 9182 9112 9236
rect 9128 9182 9148 9236
rect 9148 9182 9172 9236
rect 9172 9182 9192 9236
rect 8568 9172 8632 9182
rect 8648 9172 8712 9182
rect 8728 9172 8792 9182
rect 8808 9172 8872 9182
rect 8888 9172 8952 9182
rect 8968 9172 9032 9182
rect 9048 9172 9112 9182
rect 9128 9172 9192 9182
rect 8568 9097 8588 9153
rect 8588 9097 8612 9153
rect 8612 9097 8632 9153
rect 8648 9097 8668 9153
rect 8668 9097 8692 9153
rect 8692 9097 8712 9153
rect 8728 9097 8748 9153
rect 8748 9097 8772 9153
rect 8772 9097 8792 9153
rect 8808 9097 8828 9153
rect 8828 9097 8852 9153
rect 8852 9097 8872 9153
rect 8888 9097 8908 9153
rect 8908 9097 8932 9153
rect 8932 9097 8952 9153
rect 8968 9097 8988 9153
rect 8988 9097 9012 9153
rect 9012 9097 9032 9153
rect 9048 9097 9068 9153
rect 9068 9097 9092 9153
rect 9092 9097 9112 9153
rect 9128 9097 9148 9153
rect 9148 9097 9172 9153
rect 9172 9097 9192 9153
rect 8568 9089 8632 9097
rect 8648 9089 8712 9097
rect 8728 9089 8792 9097
rect 8808 9089 8872 9097
rect 8888 9089 8952 9097
rect 8968 9089 9032 9097
rect 9048 9089 9112 9097
rect 9128 9089 9192 9097
rect 8568 9068 8632 9070
rect 8648 9068 8712 9070
rect 8728 9068 8792 9070
rect 8808 9068 8872 9070
rect 8888 9068 8952 9070
rect 8968 9068 9032 9070
rect 9048 9068 9112 9070
rect 9128 9068 9192 9070
rect 8568 9012 8588 9068
rect 8588 9012 8612 9068
rect 8612 9012 8632 9068
rect 8648 9012 8668 9068
rect 8668 9012 8692 9068
rect 8692 9012 8712 9068
rect 8728 9012 8748 9068
rect 8748 9012 8772 9068
rect 8772 9012 8792 9068
rect 8808 9012 8828 9068
rect 8828 9012 8852 9068
rect 8852 9012 8872 9068
rect 8888 9012 8908 9068
rect 8908 9012 8932 9068
rect 8932 9012 8952 9068
rect 8968 9012 8988 9068
rect 8988 9012 9012 9068
rect 9012 9012 9032 9068
rect 9048 9012 9068 9068
rect 9068 9012 9092 9068
rect 9092 9012 9112 9068
rect 9128 9012 9148 9068
rect 9148 9012 9172 9068
rect 9172 9012 9192 9068
rect 8568 9006 8632 9012
rect 8648 9006 8712 9012
rect 8728 9006 8792 9012
rect 8808 9006 8872 9012
rect 8888 9006 8952 9012
rect 8968 9006 9032 9012
rect 9048 9006 9112 9012
rect 9128 9006 9192 9012
rect 8568 8983 8632 8986
rect 8648 8983 8712 8986
rect 8728 8983 8792 8986
rect 8808 8983 8872 8986
rect 8888 8983 8952 8986
rect 8968 8983 9032 8986
rect 9048 8983 9112 8986
rect 9128 8983 9192 8986
rect 8568 8927 8588 8983
rect 8588 8927 8612 8983
rect 8612 8927 8632 8983
rect 8648 8927 8668 8983
rect 8668 8927 8692 8983
rect 8692 8927 8712 8983
rect 8728 8927 8748 8983
rect 8748 8927 8772 8983
rect 8772 8927 8792 8983
rect 8808 8927 8828 8983
rect 8828 8927 8852 8983
rect 8852 8927 8872 8983
rect 8888 8927 8908 8983
rect 8908 8927 8932 8983
rect 8932 8927 8952 8983
rect 8968 8927 8988 8983
rect 8988 8927 9012 8983
rect 9012 8927 9032 8983
rect 9048 8927 9068 8983
rect 9068 8927 9092 8983
rect 9092 8927 9112 8983
rect 9128 8927 9148 8983
rect 9148 8927 9172 8983
rect 9172 8927 9192 8983
rect 8568 8922 8632 8927
rect 8648 8922 8712 8927
rect 8728 8922 8792 8927
rect 8808 8922 8872 8927
rect 8888 8922 8952 8927
rect 8968 8922 9032 8927
rect 9048 8922 9112 8927
rect 9128 8922 9192 8927
rect 8568 8898 8632 8902
rect 8648 8898 8712 8902
rect 8728 8898 8792 8902
rect 8808 8898 8872 8902
rect 8888 8898 8952 8902
rect 8968 8898 9032 8902
rect 9048 8898 9112 8902
rect 9128 8898 9192 8902
rect 8568 8842 8588 8898
rect 8588 8842 8612 8898
rect 8612 8842 8632 8898
rect 8648 8842 8668 8898
rect 8668 8842 8692 8898
rect 8692 8842 8712 8898
rect 8728 8842 8748 8898
rect 8748 8842 8772 8898
rect 8772 8842 8792 8898
rect 8808 8842 8828 8898
rect 8828 8842 8852 8898
rect 8852 8842 8872 8898
rect 8888 8842 8908 8898
rect 8908 8842 8932 8898
rect 8932 8842 8952 8898
rect 8968 8842 8988 8898
rect 8988 8842 9012 8898
rect 9012 8842 9032 8898
rect 9048 8842 9068 8898
rect 9068 8842 9092 8898
rect 9092 8842 9112 8898
rect 9128 8842 9148 8898
rect 9148 8842 9172 8898
rect 9172 8842 9192 8898
rect 8568 8838 8632 8842
rect 8648 8838 8712 8842
rect 8728 8838 8792 8842
rect 8808 8838 8872 8842
rect 8888 8838 8952 8842
rect 8968 8838 9032 8842
rect 9048 8838 9112 8842
rect 9128 8838 9192 8842
rect 8568 8812 8632 8818
rect 8648 8812 8712 8818
rect 8728 8812 8792 8818
rect 8808 8812 8872 8818
rect 8888 8812 8952 8818
rect 8968 8812 9032 8818
rect 9048 8812 9112 8818
rect 9128 8812 9192 8818
rect 8568 8756 8588 8812
rect 8588 8756 8612 8812
rect 8612 8756 8632 8812
rect 8648 8756 8668 8812
rect 8668 8756 8692 8812
rect 8692 8756 8712 8812
rect 8728 8756 8748 8812
rect 8748 8756 8772 8812
rect 8772 8756 8792 8812
rect 8808 8756 8828 8812
rect 8828 8756 8852 8812
rect 8852 8756 8872 8812
rect 8888 8756 8908 8812
rect 8908 8756 8932 8812
rect 8932 8756 8952 8812
rect 8968 8756 8988 8812
rect 8988 8756 9012 8812
rect 9012 8756 9032 8812
rect 9048 8756 9068 8812
rect 9068 8756 9092 8812
rect 9092 8756 9112 8812
rect 9128 8756 9148 8812
rect 9148 8756 9172 8812
rect 9172 8756 9192 8812
rect 8568 8754 8632 8756
rect 8648 8754 8712 8756
rect 8728 8754 8792 8756
rect 8808 8754 8872 8756
rect 8888 8754 8952 8756
rect 8968 8754 9032 8756
rect 9048 8754 9112 8756
rect 9128 8754 9192 8756
rect 8568 8726 8632 8734
rect 8648 8726 8712 8734
rect 8728 8726 8792 8734
rect 8808 8726 8872 8734
rect 8888 8726 8952 8734
rect 8968 8726 9032 8734
rect 9048 8726 9112 8734
rect 9128 8726 9192 8734
rect 8568 8670 8588 8726
rect 8588 8670 8612 8726
rect 8612 8670 8632 8726
rect 8648 8670 8668 8726
rect 8668 8670 8692 8726
rect 8692 8670 8712 8726
rect 8728 8670 8748 8726
rect 8748 8670 8772 8726
rect 8772 8670 8792 8726
rect 8808 8670 8828 8726
rect 8828 8670 8852 8726
rect 8852 8670 8872 8726
rect 8888 8670 8908 8726
rect 8908 8670 8932 8726
rect 8932 8670 8952 8726
rect 8968 8670 8988 8726
rect 8988 8670 9012 8726
rect 9012 8670 9032 8726
rect 9048 8670 9068 8726
rect 9068 8670 9092 8726
rect 9092 8670 9112 8726
rect 9128 8670 9148 8726
rect 9148 8670 9172 8726
rect 9172 8670 9192 8726
rect 8568 8640 8632 8650
rect 8648 8640 8712 8650
rect 8728 8640 8792 8650
rect 8808 8640 8872 8650
rect 8888 8640 8952 8650
rect 8968 8640 9032 8650
rect 9048 8640 9112 8650
rect 9128 8640 9192 8650
rect 8568 8586 8588 8640
rect 8588 8586 8612 8640
rect 8612 8586 8632 8640
rect 8648 8586 8668 8640
rect 8668 8586 8692 8640
rect 8692 8586 8712 8640
rect 8728 8586 8748 8640
rect 8748 8586 8772 8640
rect 8772 8586 8792 8640
rect 8808 8586 8828 8640
rect 8828 8586 8852 8640
rect 8852 8586 8872 8640
rect 8888 8586 8908 8640
rect 8908 8586 8932 8640
rect 8932 8586 8952 8640
rect 8968 8586 8988 8640
rect 8988 8586 9012 8640
rect 9012 8586 9032 8640
rect 9048 8586 9068 8640
rect 9068 8586 9092 8640
rect 9092 8586 9112 8640
rect 9128 8586 9148 8640
rect 9148 8586 9172 8640
rect 9172 8586 9192 8640
rect 8568 8554 8632 8566
rect 8648 8554 8712 8566
rect 8728 8554 8792 8566
rect 8808 8554 8872 8566
rect 8888 8554 8952 8566
rect 8968 8554 9032 8566
rect 9048 8554 9112 8566
rect 9128 8554 9192 8566
rect 8568 8502 8588 8554
rect 8588 8502 8612 8554
rect 8612 8502 8632 8554
rect 8648 8502 8668 8554
rect 8668 8502 8692 8554
rect 8692 8502 8712 8554
rect 8728 8502 8748 8554
rect 8748 8502 8772 8554
rect 8772 8502 8792 8554
rect 8808 8502 8828 8554
rect 8828 8502 8852 8554
rect 8852 8502 8872 8554
rect 8888 8502 8908 8554
rect 8908 8502 8932 8554
rect 8932 8502 8952 8554
rect 8968 8502 8988 8554
rect 8988 8502 9012 8554
rect 9012 8502 9032 8554
rect 9048 8502 9068 8554
rect 9068 8502 9092 8554
rect 9092 8502 9112 8554
rect 9128 8502 9148 8554
rect 9148 8502 9172 8554
rect 9172 8502 9192 8554
rect 8568 8468 8632 8482
rect 8648 8468 8712 8482
rect 8728 8468 8792 8482
rect 8808 8468 8872 8482
rect 8888 8468 8952 8482
rect 8968 8468 9032 8482
rect 9048 8468 9112 8482
rect 9128 8468 9192 8482
rect 8568 8418 8588 8468
rect 8588 8418 8612 8468
rect 8612 8418 8632 8468
rect 8648 8418 8668 8468
rect 8668 8418 8692 8468
rect 8692 8418 8712 8468
rect 8728 8418 8748 8468
rect 8748 8418 8772 8468
rect 8772 8418 8792 8468
rect 8808 8418 8828 8468
rect 8828 8418 8852 8468
rect 8852 8418 8872 8468
rect 8888 8418 8908 8468
rect 8908 8418 8932 8468
rect 8932 8418 8952 8468
rect 8968 8418 8988 8468
rect 8988 8418 9012 8468
rect 9012 8418 9032 8468
rect 9048 8418 9068 8468
rect 9068 8418 9092 8468
rect 9092 8418 9112 8468
rect 9128 8418 9148 8468
rect 9148 8418 9172 8468
rect 9172 8418 9192 8468
rect 8568 8382 8632 8398
rect 8648 8382 8712 8398
rect 8728 8382 8792 8398
rect 8808 8382 8872 8398
rect 8888 8382 8952 8398
rect 8968 8382 9032 8398
rect 9048 8382 9112 8398
rect 9128 8382 9192 8398
rect 8568 8334 8588 8382
rect 8588 8334 8612 8382
rect 8612 8334 8632 8382
rect 8648 8334 8668 8382
rect 8668 8334 8692 8382
rect 8692 8334 8712 8382
rect 8728 8334 8748 8382
rect 8748 8334 8772 8382
rect 8772 8334 8792 8382
rect 8808 8334 8828 8382
rect 8828 8334 8852 8382
rect 8852 8334 8872 8382
rect 8888 8334 8908 8382
rect 8908 8334 8932 8382
rect 8932 8334 8952 8382
rect 8968 8334 8988 8382
rect 8988 8334 9012 8382
rect 9012 8334 9032 8382
rect 9048 8334 9068 8382
rect 9068 8334 9092 8382
rect 9092 8334 9112 8382
rect 9128 8334 9148 8382
rect 9148 8334 9172 8382
rect 9172 8334 9192 8382
rect 7865 7967 7929 8031
rect 7945 7967 8009 8031
rect 8025 7967 8089 8031
rect 8105 7967 8169 8031
rect 8185 7967 8249 8031
rect 8265 7967 8329 8031
rect 8345 7967 8409 8031
rect 7865 7880 7929 7944
rect 7945 7880 8009 7944
rect 8025 7880 8089 7944
rect 8105 7880 8169 7944
rect 8185 7880 8249 7944
rect 8265 7880 8329 7944
rect 8345 7880 8409 7944
rect 7865 7793 7929 7857
rect 7945 7793 8009 7857
rect 8025 7793 8089 7857
rect 8105 7793 8169 7857
rect 8185 7793 8249 7857
rect 8265 7793 8329 7857
rect 8345 7793 8409 7857
rect 7865 7705 7929 7769
rect 7945 7705 8009 7769
rect 8025 7705 8089 7769
rect 8105 7705 8169 7769
rect 8185 7705 8249 7769
rect 8265 7705 8329 7769
rect 8345 7705 8409 7769
rect 7865 7617 7929 7681
rect 7945 7617 8009 7681
rect 8025 7617 8089 7681
rect 8105 7617 8169 7681
rect 8185 7617 8249 7681
rect 8265 7617 8329 7681
rect 8345 7617 8409 7681
rect 7865 7529 7929 7593
rect 7945 7529 8009 7593
rect 8025 7529 8089 7593
rect 8105 7529 8169 7593
rect 8185 7529 8249 7593
rect 8265 7529 8329 7593
rect 8345 7529 8409 7593
rect 7865 7441 7929 7505
rect 7945 7441 8009 7505
rect 8025 7441 8089 7505
rect 8105 7441 8169 7505
rect 8185 7441 8249 7505
rect 8265 7441 8329 7505
rect 8345 7441 8409 7505
rect 7865 7353 7929 7417
rect 7945 7353 8009 7417
rect 8025 7353 8089 7417
rect 8105 7353 8169 7417
rect 8185 7353 8249 7417
rect 8265 7353 8329 7417
rect 8345 7353 8409 7417
<< metal4 >>
rect 9346 11281 9600 11347
rect 0 10625 321 11221
rect 6993 11200 7537 11206
rect 1856 11192 2401 11198
rect 1920 11128 1936 11192
rect 2000 11128 2016 11192
rect 2080 11128 2096 11192
rect 2160 11128 2176 11192
rect 2240 11128 2256 11192
rect 2320 11128 2336 11192
rect 2400 11128 2401 11192
rect 1856 11097 2401 11128
rect 1920 11033 1936 11097
rect 2000 11033 2016 11097
rect 2080 11033 2096 11097
rect 2160 11033 2176 11097
rect 2240 11033 2256 11097
rect 2320 11033 2336 11097
rect 2400 11033 2401 11097
rect 1856 11001 2401 11033
rect 1920 10937 1936 11001
rect 2000 10937 2016 11001
rect 2080 10937 2096 11001
rect 2160 10937 2176 11001
rect 2240 10937 2256 11001
rect 2320 10937 2336 11001
rect 2400 10937 2401 11001
rect 1856 10905 2401 10937
rect 1920 10841 1936 10905
rect 2000 10841 2016 10905
rect 2080 10841 2096 10905
rect 2160 10841 2176 10905
rect 2240 10841 2256 10905
rect 2320 10841 2336 10905
rect 2400 10841 2401 10905
rect 1856 10809 2401 10841
rect 1920 10745 1936 10809
rect 2000 10745 2016 10809
rect 2080 10745 2096 10809
rect 2160 10745 2176 10809
rect 2240 10745 2256 10809
rect 2320 10745 2336 10809
rect 2400 10745 2401 10809
rect 1856 10713 2401 10745
rect 1920 10649 1936 10713
rect 2000 10649 2016 10713
rect 2080 10649 2096 10713
rect 2160 10649 2176 10713
rect 2240 10649 2256 10713
rect 2320 10649 2336 10713
rect 2400 10649 2401 10713
rect 7057 11136 7073 11200
rect 7137 11136 7153 11200
rect 7217 11136 7233 11200
rect 7297 11136 7313 11200
rect 7377 11136 7393 11200
rect 7457 11136 7473 11200
rect 6993 11105 7537 11136
rect 7057 11041 7073 11105
rect 7137 11041 7153 11105
rect 7217 11041 7233 11105
rect 7297 11041 7313 11105
rect 7377 11041 7393 11105
rect 7457 11041 7473 11105
rect 6993 11009 7537 11041
rect 7057 10945 7073 11009
rect 7137 10945 7153 11009
rect 7217 10945 7233 11009
rect 7297 10945 7313 11009
rect 7377 10945 7393 11009
rect 7457 10945 7473 11009
rect 6993 10913 7537 10945
rect 7057 10849 7073 10913
rect 7137 10849 7153 10913
rect 7217 10849 7233 10913
rect 7297 10849 7313 10913
rect 7377 10849 7393 10913
rect 7457 10849 7473 10913
rect 6993 10817 7537 10849
rect 7057 10753 7073 10817
rect 7137 10753 7153 10817
rect 7217 10753 7233 10817
rect 7297 10753 7313 10817
rect 7377 10753 7393 10817
rect 7457 10753 7473 10817
rect 6993 10721 7537 10753
rect 7057 10657 7073 10721
rect 7137 10657 7153 10721
rect 7217 10657 7233 10721
rect 7297 10657 7313 10721
rect 7377 10657 7393 10721
rect 7457 10657 7473 10721
rect 6993 10651 7537 10657
rect 1856 10643 2401 10649
rect 9346 10625 9600 11221
rect 0 9673 334 10269
rect 2921 10244 3465 10250
rect 2985 10180 3001 10244
rect 3065 10180 3081 10244
rect 3145 10180 3161 10244
rect 3225 10180 3241 10244
rect 3305 10180 3321 10244
rect 3385 10180 3401 10244
rect 2921 10149 3465 10180
rect 2985 10085 3001 10149
rect 3065 10085 3081 10149
rect 3145 10085 3161 10149
rect 3225 10085 3241 10149
rect 3305 10085 3321 10149
rect 3385 10085 3401 10149
rect 2921 10053 3465 10085
rect 2985 9989 3001 10053
rect 3065 9989 3081 10053
rect 3145 9989 3161 10053
rect 3225 9989 3241 10053
rect 3305 9989 3321 10053
rect 3385 9989 3401 10053
rect 2921 9957 3465 9989
rect 2985 9893 3001 9957
rect 3065 9893 3081 9957
rect 3145 9893 3161 9957
rect 3225 9893 3241 9957
rect 3305 9893 3321 9957
rect 3385 9893 3401 9957
rect 2921 9861 3465 9893
rect 2985 9797 3001 9861
rect 3065 9797 3081 9861
rect 3145 9797 3161 9861
rect 3225 9797 3241 9861
rect 3305 9797 3321 9861
rect 3385 9797 3401 9861
rect 2921 9765 3465 9797
rect 2985 9701 3001 9765
rect 3065 9701 3081 9765
rect 3145 9701 3161 9765
rect 3225 9701 3241 9765
rect 3305 9701 3321 9765
rect 3385 9701 3401 9765
rect 2921 9695 3465 9701
rect 5918 10236 6462 10242
rect 5982 10172 5998 10236
rect 6062 10172 6078 10236
rect 6142 10172 6158 10236
rect 6222 10172 6238 10236
rect 6302 10172 6318 10236
rect 6382 10172 6398 10236
rect 5918 10141 6462 10172
rect 5982 10077 5998 10141
rect 6062 10077 6078 10141
rect 6142 10077 6158 10141
rect 6222 10077 6238 10141
rect 6302 10077 6318 10141
rect 6382 10077 6398 10141
rect 5918 10045 6462 10077
rect 5982 9981 5998 10045
rect 6062 9981 6078 10045
rect 6142 9981 6158 10045
rect 6222 9981 6238 10045
rect 6302 9981 6318 10045
rect 6382 9981 6398 10045
rect 5918 9949 6462 9981
rect 5982 9885 5998 9949
rect 6062 9885 6078 9949
rect 6142 9885 6158 9949
rect 6222 9885 6238 9949
rect 6302 9885 6318 9949
rect 6382 9885 6398 9949
rect 5918 9853 6462 9885
rect 5982 9789 5998 9853
rect 6062 9789 6078 9853
rect 6142 9789 6158 9853
rect 6222 9789 6238 9853
rect 6302 9789 6318 9853
rect 6382 9789 6398 9853
rect 5918 9757 6462 9789
rect 5982 9693 5998 9757
rect 6062 9693 6078 9757
rect 6142 9693 6158 9757
rect 6222 9693 6238 9757
rect 6302 9693 6318 9757
rect 6382 9693 6398 9757
rect 5918 9687 6462 9693
rect 9308 9673 9600 10269
rect 9346 9547 9600 9613
rect 315 9241 381 9242
rect 315 9177 316 9241
rect 380 9177 381 9241
rect 315 9156 381 9177
rect 315 9092 316 9156
rect 380 9092 381 9156
rect 315 9071 381 9092
rect 315 9007 316 9071
rect 380 9007 381 9071
rect 315 8986 381 9007
rect 315 8922 316 8986
rect 380 8922 381 8986
rect 315 8901 381 8922
rect 315 8837 316 8901
rect 380 8837 381 8901
rect 315 8816 381 8837
rect 315 8752 316 8816
rect 380 8752 381 8816
rect 2083 9241 2483 9247
rect 2147 9177 2195 9241
rect 2259 9177 2307 9241
rect 2371 9177 2419 9241
rect 2083 9109 2483 9177
rect 2147 9045 2195 9109
rect 2259 9045 2307 9109
rect 2371 9045 2419 9109
rect 2083 8977 2483 9045
rect 2147 8913 2195 8977
rect 2259 8913 2307 8977
rect 2371 8913 2419 8977
rect 2083 8845 2483 8913
rect 2147 8781 2195 8845
rect 2259 8781 2307 8845
rect 2371 8781 2419 8845
rect 2083 8775 2483 8781
rect 8568 9236 9192 9242
rect 8632 9172 8648 9236
rect 8712 9172 8728 9236
rect 8792 9172 8808 9236
rect 8872 9172 8888 9236
rect 8952 9172 8968 9236
rect 9032 9172 9048 9236
rect 9112 9172 9128 9236
rect 8568 9153 9192 9172
rect 8632 9089 8648 9153
rect 8712 9089 8728 9153
rect 8792 9089 8808 9153
rect 8872 9089 8888 9153
rect 8952 9089 8968 9153
rect 9032 9089 9048 9153
rect 9112 9089 9128 9153
rect 8568 9070 9192 9089
rect 8632 9006 8648 9070
rect 8712 9006 8728 9070
rect 8792 9006 8808 9070
rect 8872 9006 8888 9070
rect 8952 9006 8968 9070
rect 9032 9006 9048 9070
rect 9112 9006 9128 9070
rect 8568 8986 9192 9006
rect 8632 8922 8648 8986
rect 8712 8922 8728 8986
rect 8792 8922 8808 8986
rect 8872 8922 8888 8986
rect 8952 8922 8968 8986
rect 9032 8922 9048 8986
rect 9112 8922 9128 8986
rect 8568 8902 9192 8922
rect 8632 8838 8648 8902
rect 8712 8838 8728 8902
rect 8792 8838 8808 8902
rect 8872 8838 8888 8902
rect 8952 8838 8968 8902
rect 9032 8838 9048 8902
rect 9112 8838 9128 8902
rect 8568 8818 9192 8838
rect 315 8731 381 8752
rect 315 8667 316 8731
rect 380 8667 381 8731
rect 315 8645 381 8667
rect 315 8581 316 8645
rect 380 8581 381 8645
rect 315 8559 381 8581
rect 315 8495 316 8559
rect 380 8495 381 8559
rect 315 8473 381 8495
rect 315 8409 316 8473
rect 380 8409 381 8473
rect 315 8387 381 8409
rect 315 8323 316 8387
rect 380 8323 381 8387
rect 8632 8754 8648 8818
rect 8712 8754 8728 8818
rect 8792 8754 8808 8818
rect 8872 8754 8888 8818
rect 8952 8754 8968 8818
rect 9032 8754 9048 8818
rect 9112 8754 9128 8818
rect 8568 8734 9192 8754
rect 8632 8670 8648 8734
rect 8712 8670 8728 8734
rect 8792 8670 8808 8734
rect 8872 8670 8888 8734
rect 8952 8670 8968 8734
rect 9032 8670 9048 8734
rect 9112 8670 9128 8734
rect 8568 8650 9192 8670
rect 8632 8586 8648 8650
rect 8712 8586 8728 8650
rect 8792 8586 8808 8650
rect 8872 8586 8888 8650
rect 8952 8586 8968 8650
rect 9032 8586 9048 8650
rect 9112 8586 9128 8650
rect 8568 8566 9192 8586
rect 8632 8502 8648 8566
rect 8712 8502 8728 8566
rect 8792 8502 8808 8566
rect 8872 8502 8888 8566
rect 8952 8502 8968 8566
rect 9032 8502 9048 8566
rect 9112 8502 9128 8566
rect 8568 8482 9192 8502
rect 8632 8418 8648 8482
rect 8712 8418 8728 8482
rect 8792 8418 8808 8482
rect 8872 8418 8888 8482
rect 8952 8418 8968 8482
rect 9032 8418 9048 8482
rect 9112 8418 9128 8482
rect 8568 8398 9192 8418
rect 8632 8334 8648 8398
rect 8712 8334 8728 8398
rect 8792 8334 8808 8398
rect 8872 8334 8888 8398
rect 8952 8334 8968 8398
rect 9032 8334 9048 8398
rect 9112 8334 9128 8398
rect 8568 8328 9192 8334
rect 315 8322 381 8323
rect 7848 8031 8409 8037
rect 7848 7967 7865 8031
rect 7929 7967 7945 8031
rect 8009 7967 8025 8031
rect 8089 7967 8105 8031
rect 8169 7967 8185 8031
rect 8249 7967 8265 8031
rect 8329 7967 8345 8031
rect 7848 7944 8409 7967
rect 7848 7880 7865 7944
rect 7929 7880 7945 7944
rect 8009 7880 8025 7944
rect 8089 7880 8105 7944
rect 8169 7880 8185 7944
rect 8249 7880 8265 7944
rect 8329 7880 8345 7944
rect 7848 7857 8409 7880
rect 7848 7793 7865 7857
rect 7929 7793 7945 7857
rect 8009 7793 8025 7857
rect 8089 7793 8105 7857
rect 8169 7793 8185 7857
rect 8249 7793 8265 7857
rect 8329 7793 8345 7857
rect 7848 7769 8409 7793
rect 7848 7705 7865 7769
rect 7929 7705 7945 7769
rect 8009 7705 8025 7769
rect 8089 7705 8105 7769
rect 8169 7705 8185 7769
rect 8249 7705 8265 7769
rect 8329 7705 8345 7769
rect 7848 7681 8409 7705
rect 7848 7617 7865 7681
rect 7929 7617 7945 7681
rect 8009 7617 8025 7681
rect 8089 7617 8105 7681
rect 8169 7617 8185 7681
rect 8249 7617 8265 7681
rect 8329 7617 8345 7681
rect 7848 7593 8409 7617
rect 7848 7529 7865 7593
rect 7929 7529 7945 7593
rect 8009 7529 8025 7593
rect 8089 7529 8105 7593
rect 8169 7529 8185 7593
rect 8249 7529 8265 7593
rect 8329 7529 8345 7593
rect 7848 7505 8409 7529
rect 7848 7441 7865 7505
rect 7929 7441 7945 7505
rect 8009 7441 8025 7505
rect 8089 7441 8105 7505
rect 8169 7441 8185 7505
rect 8249 7441 8265 7505
rect 8329 7441 8345 7505
rect 7848 7417 8409 7441
rect 7848 7353 7865 7417
rect 7929 7353 7945 7417
rect 8009 7353 8025 7417
rect 8089 7353 8105 7417
rect 8169 7353 8185 7417
rect 8249 7353 8265 7417
rect 8329 7353 8345 7417
rect 7848 7347 8409 7353
rect 490 7041 824 7047
rect 554 6977 580 7041
rect 644 6977 670 7041
rect 734 6977 760 7041
rect 490 6960 824 6977
rect 554 6896 580 6960
rect 644 6896 670 6960
rect 734 6896 760 6960
rect 490 6878 824 6896
rect 554 6814 580 6878
rect 644 6814 670 6878
rect 734 6814 760 6878
rect 490 6796 824 6814
rect 554 6732 580 6796
rect 644 6732 670 6796
rect 734 6732 760 6796
rect 490 6714 824 6732
rect 554 6650 580 6714
rect 644 6650 670 6714
rect 734 6650 760 6714
rect 490 6632 824 6650
rect 554 6568 580 6632
rect 644 6568 670 6632
rect 734 6568 760 6632
rect 490 6550 824 6568
rect 554 6486 580 6550
rect 644 6486 670 6550
rect 734 6486 760 6550
rect 490 6468 824 6486
rect 554 6404 580 6468
rect 644 6404 670 6468
rect 734 6404 760 6468
rect 490 6398 824 6404
rect 965 3666 1535 3672
rect 965 3602 975 3666
rect 1039 3602 1057 3666
rect 1121 3602 1139 3666
rect 1203 3602 1221 3666
rect 1285 3602 1303 3666
rect 1367 3602 1385 3666
rect 1449 3602 1467 3666
rect 1531 3602 1535 3666
rect 965 3581 1535 3602
rect 965 3517 975 3581
rect 1039 3517 1057 3581
rect 1121 3517 1139 3581
rect 1203 3517 1221 3581
rect 1285 3517 1303 3581
rect 1367 3517 1385 3581
rect 1449 3517 1467 3581
rect 1531 3517 1535 3581
rect 965 3495 1535 3517
rect 965 3431 975 3495
rect 1039 3431 1057 3495
rect 1121 3431 1139 3495
rect 1203 3431 1221 3495
rect 1285 3431 1303 3495
rect 1367 3431 1385 3495
rect 1449 3431 1467 3495
rect 1531 3431 1535 3495
rect 965 3409 1535 3431
rect 965 3345 975 3409
rect 1039 3345 1057 3409
rect 1121 3345 1139 3409
rect 1203 3345 1221 3409
rect 1285 3345 1303 3409
rect 1367 3345 1385 3409
rect 1449 3345 1467 3409
rect 1531 3345 1535 3409
rect 965 3323 1535 3345
rect 965 3259 975 3323
rect 1039 3259 1057 3323
rect 1121 3259 1139 3323
rect 1203 3259 1221 3323
rect 1285 3259 1303 3323
rect 1367 3259 1385 3323
rect 1449 3259 1467 3323
rect 1531 3259 1535 3323
rect 965 3237 1535 3259
rect 965 3173 975 3237
rect 1039 3173 1057 3237
rect 1121 3173 1139 3237
rect 1203 3173 1221 3237
rect 1285 3173 1303 3237
rect 1367 3173 1385 3237
rect 1449 3173 1467 3237
rect 1531 3173 1535 3237
rect 965 3151 1535 3173
rect 965 3087 975 3151
rect 1039 3087 1057 3151
rect 1121 3087 1139 3151
rect 1203 3087 1221 3151
rect 1285 3087 1303 3151
rect 1367 3087 1385 3151
rect 1449 3087 1467 3151
rect 1531 3087 1535 3151
rect 965 3065 1535 3087
rect 965 3001 975 3065
rect 1039 3001 1057 3065
rect 1121 3001 1139 3065
rect 1203 3001 1221 3065
rect 1285 3001 1303 3065
rect 1367 3001 1385 3065
rect 1449 3001 1467 3065
rect 1531 3001 1535 3065
rect 965 2995 1535 3001
rect 4427 2701 4602 2707
rect 4427 2637 4428 2701
rect 4492 2637 4538 2701
rect 4427 2616 4602 2637
rect 4427 2552 4428 2616
rect 4492 2552 4538 2616
rect 4427 2531 4602 2552
rect 4427 2467 4428 2531
rect 4492 2467 4538 2531
rect 4427 2446 4602 2467
rect 4427 2382 4428 2446
rect 4492 2382 4538 2446
rect 4427 2361 4602 2382
rect 4427 2297 4428 2361
rect 4492 2297 4538 2361
rect 4427 2276 4602 2297
rect 4427 2212 4428 2276
rect 4492 2212 4538 2276
rect 4427 2191 4602 2212
rect 4427 2127 4428 2191
rect 4492 2127 4538 2191
rect 4427 2105 4602 2127
rect 4427 2041 4428 2105
rect 4492 2041 4538 2105
rect 4427 2019 4602 2041
rect 4427 1955 4428 2019
rect 4492 1955 4538 2019
rect 4427 1933 4602 1955
rect 4427 1869 4428 1933
rect 4492 1869 4538 1933
rect 4427 1847 4602 1869
rect 4427 1783 4428 1847
rect 4492 1783 4538 1847
rect 4427 1777 4602 1783
<< metal5 >>
rect 0 35157 254 40000
rect 9346 35157 9600 40000
rect 0 14007 254 18997
rect 9346 14007 9600 18997
rect 0 12837 254 13687
rect 9346 12837 9600 13687
rect 0 11667 254 12517
rect 9346 11667 9600 12517
rect 0 9547 254 11347
rect 9346 9547 9600 11347
rect 0 8337 254 9227
rect 9346 8337 9600 9227
rect 0 7368 254 8017
rect 9346 7368 9600 8017
rect 0 6397 254 7047
rect 9346 6397 9600 7047
rect 0 5187 254 6077
rect 9346 5187 9600 6077
rect 0 3977 254 4867
rect 9346 3977 9600 4867
rect 0 3007 193 3657
rect 9407 3007 9600 3657
rect 0 1797 254 2687
rect 9346 1797 9600 2687
rect 0 427 254 1477
rect 9346 427 9600 1477
use sky130_fd_io__amuxsplitv2_busses  sky130_fd_io__amuxsplitv2_busses_0
timestamp 1707688321
transform 1 0 0 0 1 407
box 0 0 9600 39593
use sky130_fd_io__amuxsplitv2_delay  sky130_fd_io__amuxsplitv2_delay_0
timestamp 1707688321
transform -1 0 7359 0 -1 3222
box 0 0 2135 1333
use sky130_fd_io__amuxsplitv2_switch  sky130_fd_io__amuxsplitv2_switch_0
timestamp 1707688321
transform 0 -1 7760 1 0 18566
box -148 -12 10507 5940
use sky130_fd_io__amuxsplitv2_switch  sky130_fd_io__amuxsplitv2_switch_1
timestamp 1707688321
transform 0 -1 7760 -1 0 39852
box -148 -12 10507 5940
use sky130_fd_io__amuxsplitv2_switch_s0  sky130_fd_io__amuxsplitv2_switch_s0_0
timestamp 1707688321
transform 0 -1 7246 -1 0 6134
box -8 14 1474 4390
use sky130_fd_io__amuxsplitv2_switch_s0  sky130_fd_io__amuxsplitv2_switch_s0_1
timestamp 1707688321
transform 0 -1 7246 1 0 3272
box -8 14 1474 4390
use sky130_fd_io__amuxsplitv2_switch_sl  sky130_fd_io__amuxsplitv2_switch_sl_0
timestamp 1707688321
transform 0 -1 7246 -1 0 11182
box -8 14 2602 4390
use sky130_fd_io__amuxsplitv2_switch_sl  sky130_fd_io__amuxsplitv2_switch_sl_1
timestamp 1707688321
transform 0 -1 7246 -1 0 16230
box -8 14 2602 4390
use sky130_fd_io__amuxsplitv2_switch_sl  sky130_fd_io__amuxsplitv2_switch_sl_2
timestamp 1707688321
transform 0 -1 7246 1 0 6064
box -8 14 2602 4390
use sky130_fd_io__amuxsplitv2_switch_sl  sky130_fd_io__amuxsplitv2_switch_sl_3
timestamp 1707688321
transform 0 -1 7246 1 0 11112
box -8 14 2602 4390
<< labels >>
flabel metal4 s 9346 10625 9600 11221 3 FreeSans 520 90 0 0 amuxbus_a_r
port 2 nsew signal bidirectional
flabel metal4 s 0 10625 321 11221 3 FreeSans 520 90 0 0 amuxbus_a_l
port 3 nsew signal bidirectional
flabel metal4 s 9346 11281 9600 11347 3 FreeSans 520 180 0 0 vssa
port 4 nsew ground bidirectional
flabel metal4 s 9346 9547 9600 9613 3 FreeSans 520 180 0 0 vssa
port 4 nsew ground bidirectional
flabel metal4 s 9308 9673 9600 10269 3 FreeSans 520 90 0 0 amuxbus_b_r
port 5 nsew signal bidirectional
flabel metal4 s 0 9673 334 10269 3 FreeSans 520 90 0 0 amuxbus_b_l
port 6 nsew signal bidirectional
flabel metal2 s 6278 0 6330 128 3 FreeSans 520 90 0 0 enable_vdda_h
port 8 nsew signal input
flabel metal2 s 7158 0 7210 128 3 FreeSans 520 90 0 0 hld_vdda_h_n
port 9 nsew signal input
flabel metal2 s 2404 0 2456 128 3 FreeSans 520 90 0 0 switch_aa_s0
port 10 nsew signal input
flabel metal2 s 2656 0 2708 128 3 FreeSans 520 90 0 0 switch_aa_sl
port 11 nsew signal input
flabel metal2 s 1312 0 1364 128 3 FreeSans 520 90 0 0 switch_aa_sr
port 12 nsew signal input
flabel metal2 s 2152 0 2204 128 3 FreeSans 520 90 0 0 switch_bb_s0
port 13 nsew signal input
flabel metal2 s 1900 0 1952 128 3 FreeSans 520 90 0 0 switch_bb_sl
port 14 nsew signal input
flabel metal2 s 1648 0 1700 128 3 FreeSans 520 90 0 0 switch_bb_sr
port 15 nsew signal input
flabel metal5 s 9346 9547 9600 11347 3 FreeSans 520 180 0 0 vssa
port 4 nsew ground bidirectional
flabel metal5 s 9407 3007 9600 3657 3 FreeSans 520 180 0 0 vdda
port 16 nsew power bidirectional
flabel metal5 s 9346 8337 9600 9227 3 FreeSans 520 180 0 0 vssd
port 17 nsew ground bidirectional
flabel metal5 s 9346 11667 9600 12517 3 FreeSans 520 180 0 0 vssio_q
port 18 nsew ground bidirectional
flabel metal5 s 9346 5187 9600 6077 3 FreeSans 520 180 0 0 vssio
port 19 nsew ground bidirectional
flabel metal5 s 9346 6397 9600 7047 3 FreeSans 520 180 0 0 vswitch
port 20 nsew power bidirectional
flabel metal5 s 9346 7368 9600 8017 3 FreeSans 520 180 0 0 vssa
port 4 nsew ground bidirectional
flabel metal5 s 9346 1797 9600 2687 3 FreeSans 520 180 0 0 vccd
port 21 nsew power bidirectional
flabel metal5 s 9346 35157 9600 40000 3 FreeSans 520 180 0 0 vssio
port 19 nsew ground bidirectional
flabel metal5 s 9346 12837 9600 13687 3 FreeSans 520 180 0 0 vddio_q
port 22 nsew power bidirectional
flabel metal5 s 9346 14007 9600 18997 3 FreeSans 520 180 0 0 vddio
port 23 nsew power bidirectional
flabel metal5 s 0 3977 254 4867 3 FreeSans 520 0 0 0 vddio
port 23 nsew power bidirectional
flabel metal5 s 0 427 254 1477 3 FreeSans 520 0 0 0 vcchib
port 24 nsew power bidirectional
flabel metal5 s 0 14007 254 18997 3 FreeSans 520 0 0 0 vddio
port 23 nsew power bidirectional
flabel metal5 s 0 12837 254 13687 3 FreeSans 520 0 0 0 vddio_q
port 22 nsew power bidirectional
flabel metal5 s 0 1797 254 2687 3 FreeSans 520 0 0 0 vccd
port 21 nsew power bidirectional
flabel metal5 s 0 7368 254 8017 3 FreeSans 520 0 0 0 vssa
port 4 nsew ground bidirectional
flabel metal5 s 0 6397 254 7047 3 FreeSans 520 0 0 0 vswitch
port 20 nsew power bidirectional
flabel metal5 s 0 5187 254 6077 3 FreeSans 520 0 0 0 vssio
port 19 nsew ground bidirectional
flabel metal5 s 0 11667 254 12517 3 FreeSans 520 0 0 0 vssio_q
port 18 nsew ground bidirectional
flabel metal5 s 0 8337 254 9227 3 FreeSans 520 0 0 0 vssd
port 17 nsew ground bidirectional
flabel metal5 s 0 3007 193 3657 3 FreeSans 520 0 0 0 vdda
port 16 nsew power bidirectional
flabel metal5 s 0 9547 254 11347 3 FreeSans 520 0 0 0 vssa
port 4 nsew ground bidirectional
flabel metal5 s 0 35157 254 40000 3 FreeSans 520 180 0 0 vssio
port 19 nsew ground bidirectional
flabel metal5 s 9346 3977 9600 4867 3 FreeSans 520 180 0 0 vddio
port 23 nsew power bidirectional
flabel metal5 s 9346 427 9600 1477 3 FreeSans 520 180 0 0 vcchib
port 24 nsew power bidirectional
flabel metal1 s 2152 0 2204 128 3 FreeSans 520 90 0 0 switch_bb_s0
port 13 nsew signal input
flabel metal1 s 1900 0 1952 128 3 FreeSans 520 90 0 0 switch_bb_sl
port 14 nsew signal input
flabel metal1 s 1648 0 1700 128 3 FreeSans 520 90 0 0 switch_bb_sr
port 15 nsew signal input
flabel metal1 s 2404 0 2456 154 3 FreeSans 520 90 0 0 switch_aa_s0
port 10 nsew signal input
flabel metal1 s 2656 0 2708 154 3 FreeSans 520 90 0 0 switch_aa_sl
port 11 nsew signal input
flabel metal1 s 1312 0 1364 154 3 FreeSans 520 90 0 0 switch_aa_sr
port 12 nsew signal input
flabel metal1 s 6278 0 6330 128 3 FreeSans 520 90 0 0 enable_vdda_h
port 8 nsew signal input
flabel metal1 s 7158 0 7210 128 3 FreeSans 520 90 0 0 hld_vdda_h_n
port 9 nsew signal input
flabel comment s 4862 26904 4862 26904 0 FreeSans 200 90 0 0 pgate_sl_h_n
flabel comment s 5025 26904 5025 26904 0 FreeSans 200 90 0 0 ngate_sr_h
flabel comment s 8075 18518 8075 18518 0 FreeSans 200 90 0 0 pgate_sl_h_n
flabel comment s 4555 31273 4555 31273 0 FreeSans 200 90 0 0 ngate_sl_h
flabel comment s 4729 31273 4729 31273 0 FreeSans 200 90 0 0 pgate_sl_h_n
flabel comment s 4853 31273 4853 31273 0 FreeSans 200 90 0 0 pgate_sr_h_n
flabel comment s 4941 31273 4941 31273 0 FreeSans 200 90 0 0 nmid_h
flabel comment s 5028 31273 5028 31273 0 FreeSans 200 90 0 0 ngate_sr_h
flabel comment s 1496 28719 1496 28719 0 FreeSans 200 90 0 0 ngate_sr_h
flabel comment s 1413 28719 1413 28719 0 FreeSans 200 90 0 0 nmid_h
flabel comment s 1332 28719 1332 28719 0 FreeSans 200 90 0 0 pgate_sr_h_n
flabel comment s 1249 28719 1249 28719 0 FreeSans 200 90 0 0 pgate_sl_h_n
flabel comment s 1162 28719 1162 28719 0 FreeSans 200 90 0 0 ngate_sl_h
flabel comment s 1496 17899 1496 17899 0 FreeSans 200 90 0 0 ngate_sr_h
flabel comment s 1162 17899 1162 17899 0 FreeSans 200 90 0 0 ngate_sl_h
flabel comment s 1249 17899 1249 17899 0 FreeSans 200 90 0 0 pgate_sl_h_n
flabel comment s 1332 17899 1332 17899 0 FreeSans 200 90 0 0 pgate_sr_h_n
flabel comment s 1413 17899 1413 17899 0 FreeSans 200 90 0 0 nmid_h
flabel comment s 4771 26904 4771 26904 0 FreeSans 200 90 0 0 nmid_h
flabel comment s 4939 26904 4939 26904 0 FreeSans 200 90 0 0 pgate_sr_h_n
flabel comment s 8249 18518 8249 18518 0 FreeSans 200 90 0 0 ngate_sl_h
flabel comment s 8166 18518 8166 18518 0 FreeSans 200 90 0 0 nmid_h
flabel comment s 4552 26904 4552 26904 0 FreeSans 200 90 0 0 ngate_sl_h
flabel comment s 8249 26904 8249 26904 0 FreeSans 200 90 0 0 ngate_sl_h
flabel comment s 8166 26904 8166 26904 0 FreeSans 200 90 0 0 nmid_h
flabel comment s 8075 26904 8075 26904 0 FreeSans 200 90 0 0 pgate_sl_h_n
flabel comment s 7998 26904 7998 26904 0 FreeSans 200 90 0 0 pgate_sr_h_n
flabel comment s 7912 26904 7912 26904 0 FreeSans 200 90 0 0 ngate_sr_h
flabel comment s 1846 17414 1846 17414 0 FreeSans 200 90 0 0 nmid_h
flabel comment s 1755 17414 1755 17414 0 FreeSans 200 90 0 0 pgate_sl_h_n
flabel comment s 1678 17414 1678 17414 0 FreeSans 200 90 0 0 pgate_sr_h_n
flabel comment s 1592 17414 1592 17414 0 FreeSans 200 90 0 0 ngate_sr_h
flabel comment s 1929 17414 1929 17414 0 FreeSans 200 90 0 0 ngate_sl_h
flabel comment s 7912 18518 7912 18518 0 FreeSans 200 90 0 0 ngate_sr_h
flabel comment s 7998 18518 7998 18518 0 FreeSans 200 90 0 0 pgate_sr_h_n
flabel comment s 7309 5759 7309 5759 0 FreeSans 600 90 0 0 condiode
flabel comment s 1918 1668 1918 1668 0 FreeSans 200 90 0 0 switch_bb_sl
flabel comment s 2178 1668 2178 1668 0 FreeSans 200 90 0 0 switch_bb_s0
flabel comment s 1333 1668 1333 1668 0 FreeSans 200 90 0 0 switch_aa_sr
flabel comment s 2678 1668 2678 1668 0 FreeSans 200 90 0 0 switch_aa_sl
flabel comment s 2428 1668 2428 1668 0 FreeSans 200 90 0 0 switch_aa_s0
flabel comment s 1670 1668 1670 1668 0 FreeSans 200 90 0 0 switch_bb_sr
flabel comment s 1846 14890 1846 14890 0 FreeSans 200 90 0 0 nmid_h
flabel comment s 1755 14890 1755 14890 0 FreeSans 200 90 0 0 pgate_sl_h_n
flabel comment s 1678 15884 1678 15884 0 FreeSans 200 90 0 0 pgate_sr_h_n
flabel comment s 1592 14890 1592 14890 0 FreeSans 200 90 0 0 ngate_sr_h
flabel comment s 1929 14890 1929 14890 0 FreeSans 200 90 0 0 ngate_sl_h
flabel comment s 1496 10686 1496 10686 0 FreeSans 200 90 0 0 ngate_sr_h
flabel comment s 1162 10686 1162 10686 0 FreeSans 200 90 0 0 ngate_sl_h
flabel comment s 1249 10686 1249 10686 0 FreeSans 200 90 0 0 pgate_sl_h_n
flabel comment s 1332 10686 1332 10686 0 FreeSans 200 90 0 0 pgate_sr_h_n
flabel comment s 1413 10686 1413 10686 0 FreeSans 200 90 0 0 nmid_h
rlabel metal1 s 1648 0 1700 15303 1 switch_bb_sr
port 15 nsew signal input
rlabel metal1 s 1900 0 1952 12245 1 switch_bb_sl
port 14 nsew signal input
rlabel metal1 s 2152 0 2204 5207 1 switch_bb_s0
port 13 nsew signal input
rlabel metal1 s 1312 0 1364 10255 1 switch_aa_sr
port 12 nsew signal input
rlabel metal1 s 2656 0 2708 7197 1 switch_aa_sl
port 11 nsew signal input
rlabel metal1 s 2404 0 2456 4405 1 switch_aa_s0
port 10 nsew signal input
rlabel metal1 s 7158 0 7210 128 1 hld_vdda_h_n
port 9 nsew signal input
rlabel metal1 s 6278 0 6330 128 1 enable_vdda_h
port 8 nsew signal input
rlabel metal5 s 0 427 254 1477 1 vcchib
port 24 nsew power bidirectional
rlabel metal5 s 0 3977 254 4867 1 vddio
port 23 nsew power bidirectional
rlabel metal5 s 0 14007 254 18997 1 vddio
port 23 nsew power bidirectional
rlabel metal5 s 9346 14007 9600 18997 1 vddio
port 23 nsew power bidirectional
rlabel metal5 s 9346 12837 9600 13687 1 vddio_q
port 22 nsew power bidirectional
rlabel metal5 s 9346 1797 9600 2687 1 vccd
port 21 nsew power bidirectional
rlabel metal5 s 9346 6397 9600 7047 1 vswitch
port 20 nsew power bidirectional
rlabel metal5 s 9346 5187 9600 6077 1 vssio
port 19 nsew ground bidirectional
rlabel metal5 s 0 35157 254 40000 1 vssio
port 19 nsew ground bidirectional
rlabel metal5 s 9346 35157 9600 40000 1 vssio
port 19 nsew ground bidirectional
rlabel metal5 s 9346 11667 9600 12517 1 vssio_q
port 18 nsew ground bidirectional
rlabel metal5 s 9346 8337 9600 9227 1 vssd
port 17 nsew ground bidirectional
rlabel metal5 s 9407 3007 9600 3657 1 vdda
port 16 nsew power bidirectional
rlabel metal5 s 9346 7368 9600 8017 1 vssa
port 4 nsew ground bidirectional
rlabel metal5 s 0 9547 254 11347 1 vssa
port 4 nsew ground bidirectional
rlabel metal5 s 9346 9547 9600 11347 1 vssa
port 4 nsew ground bidirectional
rlabel metal4 s 9346 9547 9600 9613 1 vssa
port 4 nsew ground bidirectional
rlabel metal4 s 9346 11281 9600 11347 1 vssa
port 4 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 9600 40000
string GDS_END 2728554
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 829610
string LEFclass PAD
string LEFsymmetry X Y R90
<< end >>
