magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -82 -26 650 176
<< mvnmos >>
rect 0 0 100 150
rect 156 0 256 150
rect 312 0 412 150
rect 468 0 568 150
<< mvndiff >>
rect -56 114 0 150
rect -56 80 -45 114
rect -11 80 0 114
rect -56 46 0 80
rect -56 12 -45 46
rect -11 12 0 46
rect -56 0 0 12
rect 100 114 156 150
rect 100 80 111 114
rect 145 80 156 114
rect 100 46 156 80
rect 100 12 111 46
rect 145 12 156 46
rect 100 0 156 12
rect 256 114 312 150
rect 256 80 267 114
rect 301 80 312 114
rect 256 46 312 80
rect 256 12 267 46
rect 301 12 312 46
rect 256 0 312 12
rect 412 114 468 150
rect 412 80 423 114
rect 457 80 468 114
rect 412 46 468 80
rect 412 12 423 46
rect 457 12 468 46
rect 412 0 468 12
rect 568 114 624 150
rect 568 80 579 114
rect 613 80 624 114
rect 568 46 624 80
rect 568 12 579 46
rect 613 12 624 46
rect 568 0 624 12
<< mvndiffc >>
rect -45 80 -11 114
rect -45 12 -11 46
rect 111 80 145 114
rect 111 12 145 46
rect 267 80 301 114
rect 267 12 301 46
rect 423 80 457 114
rect 423 12 457 46
rect 579 80 613 114
rect 579 12 613 46
<< poly >>
rect 0 150 100 182
rect 156 150 256 182
rect 312 150 412 182
rect 468 150 568 182
rect 0 -32 100 0
rect 156 -32 256 0
rect 312 -32 412 0
rect 468 -32 568 0
<< locali >>
rect -45 114 -11 130
rect -45 46 -11 68
rect 111 114 145 130
rect 111 46 145 68
rect 267 114 301 130
rect 267 46 301 68
rect 423 114 457 130
rect 423 46 457 68
rect 579 114 613 130
rect 579 46 613 68
<< viali >>
rect -45 80 -11 102
rect -45 68 -11 80
rect -45 12 -11 30
rect -45 -4 -11 12
rect 111 80 145 102
rect 111 68 145 80
rect 111 12 145 30
rect 111 -4 145 12
rect 267 80 301 102
rect 267 68 301 80
rect 267 12 301 30
rect 267 -4 301 12
rect 423 80 457 102
rect 423 68 457 80
rect 423 12 457 30
rect 423 -4 457 12
rect 579 80 613 102
rect 579 68 613 80
rect 579 12 613 30
rect 579 -4 613 12
<< metal1 >>
rect -51 102 -5 114
rect -51 68 -45 102
rect -11 68 -5 102
rect -51 30 -5 68
rect -51 -4 -45 30
rect -11 -4 -5 30
rect -51 -16 -5 -4
rect 105 102 151 114
rect 105 68 111 102
rect 145 68 151 102
rect 105 30 151 68
rect 105 -4 111 30
rect 145 -4 151 30
rect 105 -16 151 -4
rect 261 102 307 114
rect 261 68 267 102
rect 301 68 307 102
rect 261 30 307 68
rect 261 -4 267 30
rect 301 -4 307 30
rect 261 -16 307 -4
rect 417 102 463 114
rect 417 68 423 102
rect 457 68 463 102
rect 417 30 463 68
rect 417 -4 423 30
rect 457 -4 463 30
rect 417 -16 463 -4
rect 573 102 619 114
rect 573 68 579 102
rect 613 68 619 102
rect 573 30 619 68
rect 573 -4 579 30
rect 613 -4 619 30
rect 573 -16 619 -4
use hvDFM1sd2_CDNS_52468879185875  hvDFM1sd2_CDNS_52468879185875_0
timestamp 1707688321
transform -1 0 0 0 1 0
box 0 0 1 1
use hvDFM1sd2_CDNS_52468879185875  hvDFM1sd2_CDNS_52468879185875_1
timestamp 1707688321
transform 1 0 568 0 1 0
box 0 0 1 1
use hvDFM1sd2_CDNS_52468879185875  hvDFM1sd2_CDNS_52468879185875_2
timestamp 1707688321
transform 1 0 412 0 1 0
box 0 0 1 1
use hvDFM1sd2_CDNS_52468879185875  hvDFM1sd2_CDNS_52468879185875_3
timestamp 1707688321
transform 1 0 256 0 1 0
box 0 0 1 1
use hvDFM1sd2_CDNS_52468879185875  hvDFM1sd2_CDNS_52468879185875_4
timestamp 1707688321
transform 1 0 100 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 49 -28 49 0 FreeSans 300 0 0 0 S
flabel comment s 128 49 128 49 0 FreeSans 300 0 0 0 D
flabel comment s 284 49 284 49 0 FreeSans 300 0 0 0 S
flabel comment s 440 49 440 49 0 FreeSans 300 0 0 0 D
flabel comment s 596 49 596 49 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 7611768
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7609374
<< end >>
