magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< poly >>
rect 770 54 930 83
rect 770 20 799 54
rect 833 20 867 54
rect 901 20 930 54
rect 770 4 930 20
<< polycont >>
rect 799 20 833 54
rect 867 20 901 54
<< locali >>
rect 834 4062 1941 4096
rect 800 4024 1941 4062
rect 834 3990 1941 4024
rect 834 3916 1173 3950
rect 800 3878 1173 3916
rect 834 3844 1173 3878
rect 60 3748 98 3782
rect 317 3748 355 3782
rect 525 3286 659 3782
rect 525 3252 539 3286
rect 573 3252 611 3286
rect 645 3252 659 3286
rect 783 3286 917 3782
rect 1039 3748 1173 3844
rect 1807 3726 1941 3990
rect 783 3252 795 3286
rect 829 3252 867 3286
rect 901 3252 917 3286
rect 525 2992 539 3026
rect 573 2992 611 3026
rect 645 2992 659 3026
rect 525 2514 659 2992
rect 783 2992 797 3026
rect 831 2992 869 3026
rect 903 2992 917 3026
rect 783 1786 917 2992
rect 783 1752 797 1786
rect 831 1752 869 1786
rect 903 1752 917 1786
rect 831 1418 869 1452
rect 831 1310 869 1344
rect 831 976 869 1010
rect 831 868 869 902
rect 831 534 869 568
rect 831 426 869 460
rect 831 92 869 126
rect 783 44 799 54
rect 783 20 797 44
rect 833 20 867 54
rect 901 44 917 54
rect 903 20 917 44
rect 831 10 869 20
<< viali >>
rect 800 4062 834 4096
rect 800 3990 834 4024
rect 800 3916 834 3950
rect 800 3844 834 3878
rect 26 3748 60 3782
rect 98 3748 132 3782
rect 283 3748 317 3782
rect 355 3748 389 3782
rect 539 3252 573 3286
rect 611 3252 645 3286
rect 795 3252 829 3286
rect 867 3252 901 3286
rect 539 2992 573 3026
rect 611 2992 645 3026
rect 797 2992 831 3026
rect 869 2992 903 3026
rect 797 1752 831 1786
rect 869 1752 903 1786
rect 797 1418 831 1452
rect 869 1418 903 1452
rect 797 1310 831 1344
rect 869 1310 903 1344
rect 797 976 831 1010
rect 869 976 903 1010
rect 797 868 831 902
rect 869 868 903 902
rect 797 534 831 568
rect 869 534 903 568
rect 797 426 831 460
rect 869 426 903 460
rect 797 92 831 126
rect 869 92 903 126
rect 797 20 799 44
rect 799 20 831 44
rect 869 20 901 44
rect 901 20 903 44
rect 797 10 831 20
rect 869 10 903 20
<< metal1 >>
rect 318 4106 846 4112
rect 370 4096 846 4106
rect 370 4062 800 4096
rect 834 4062 846 4096
rect 370 4054 846 4062
rect 318 4042 846 4054
rect 370 4024 846 4042
rect 370 3990 800 4024
rect 834 3990 846 4024
rect 318 3984 846 3990
tri 352 3950 358 3956 se
rect 358 3950 846 3956
tri 318 3916 352 3950 se
rect 352 3916 800 3950
rect 834 3916 846 3950
tri 280 3878 318 3916 se
rect 318 3878 846 3916
tri 271 3869 280 3878 se
rect 280 3869 800 3878
rect 271 3844 800 3869
rect 834 3844 846 3878
rect 271 3838 846 3844
rect 14 3782 144 3788
rect 14 3748 26 3782
rect 60 3748 98 3782
rect 132 3748 144 3782
rect 14 3129 144 3748
rect 271 3782 401 3838
tri 401 3824 415 3838 nw
rect 271 3748 283 3782
rect 317 3748 355 3782
rect 389 3748 401 3782
rect 271 3742 401 3748
rect 525 3286 915 3292
rect 525 3252 539 3286
rect 573 3252 611 3286
rect 645 3252 795 3286
rect 829 3252 867 3286
rect 901 3252 915 3286
rect 525 3246 915 3252
rect 525 3167 657 3246
tri 657 3221 682 3246 nw
tri 758 3221 783 3246 ne
rect 526 3165 656 3166
rect 783 3169 915 3246
rect 784 3167 914 3168
tri 144 3129 170 3155 sw
rect 783 3131 915 3167
rect 784 3130 914 3131
rect 14 3103 170 3129
tri 170 3103 196 3129 sw
rect 526 3128 656 3129
rect 14 3102 196 3103
tri 14 3080 36 3102 ne
rect 36 3080 196 3102
tri 196 3080 219 3103 sw
tri 502 3080 525 3103 se
rect 525 3080 657 3127
tri 36 3075 41 3080 ne
rect 41 3075 657 3080
tri 41 3032 84 3075 ne
rect 84 3032 657 3075
tri 84 3026 90 3032 ne
rect 90 3026 657 3032
tri 90 2992 124 3026 ne
rect 124 2992 539 3026
rect 573 2992 611 3026
rect 645 2992 657 3026
tri 124 2986 130 2992 ne
rect 130 2986 657 2992
rect 783 3026 915 3129
rect 783 2992 797 3026
rect 831 2992 869 3026
rect 903 2992 915 3026
rect 783 2986 915 2992
rect 785 1786 917 1792
rect 785 1752 797 1786
rect 831 1752 869 1786
rect 903 1752 917 1786
rect 785 1625 917 1752
rect 786 1623 916 1624
rect 785 1587 917 1623
rect 786 1586 916 1587
rect 785 1452 917 1585
rect 785 1418 797 1452
rect 831 1418 869 1452
rect 903 1418 917 1452
rect 785 1344 917 1418
rect 785 1310 797 1344
rect 831 1310 869 1344
rect 903 1310 917 1344
rect 785 1162 917 1310
rect 786 1160 916 1161
rect 785 1124 917 1160
rect 786 1123 916 1124
rect 785 1010 917 1122
rect 785 976 797 1010
rect 831 976 869 1010
rect 903 976 917 1010
rect 785 902 917 976
rect 785 868 797 902
rect 831 868 869 902
rect 903 868 917 902
rect 785 737 917 868
rect 786 735 916 736
rect 785 699 917 735
rect 786 698 916 699
rect 785 568 917 697
rect 785 534 797 568
rect 831 534 869 568
rect 903 534 917 568
rect 785 460 917 534
rect 785 426 797 460
rect 831 426 869 460
rect 903 426 917 460
rect 785 293 917 426
rect 786 291 916 292
rect 785 255 917 291
rect 786 254 916 255
rect 785 201 917 253
rect 785 126 917 132
rect 785 92 797 126
rect 831 92 869 126
rect 903 92 917 126
rect 785 44 917 92
rect 785 10 797 44
rect 831 10 869 44
rect 903 10 917 44
rect 785 4 917 10
<< rmetal1 >>
rect 525 3166 657 3167
rect 525 3165 526 3166
rect 656 3165 657 3166
rect 783 3168 915 3169
rect 783 3167 784 3168
rect 914 3167 915 3168
rect 783 3130 784 3131
rect 914 3130 915 3131
rect 783 3129 915 3130
rect 525 3128 526 3129
rect 656 3128 657 3129
rect 525 3127 657 3128
rect 785 1624 917 1625
rect 785 1623 786 1624
rect 916 1623 917 1624
rect 785 1586 786 1587
rect 916 1586 917 1587
rect 785 1585 917 1586
rect 785 1161 917 1162
rect 785 1160 786 1161
rect 916 1160 917 1161
rect 785 1123 786 1124
rect 916 1123 917 1124
rect 785 1122 917 1123
rect 785 736 917 737
rect 785 735 786 736
rect 916 735 917 736
rect 785 698 786 699
rect 916 698 917 699
rect 785 697 917 698
rect 785 292 917 293
rect 785 291 786 292
rect 916 291 917 292
rect 785 254 786 255
rect 916 254 917 255
rect 785 253 917 254
<< via1 >>
rect 318 4054 370 4106
rect 318 3990 370 4042
<< metal2 >>
rect 318 4106 370 4112
rect 318 4042 370 4054
rect 318 3984 370 3990
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1707688321
transform 1 0 800 0 1 3990
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_1
timestamp 1707688321
transform 1 0 800 0 1 3844
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1707688321
transform -1 0 645 0 1 2992
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1707688321
transform -1 0 645 0 1 3252
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1707688321
transform -1 0 903 0 -1 3026
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1707688321
transform 1 0 283 0 -1 3782
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1707688321
transform 1 0 26 0 -1 3782
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1707688321
transform 1 0 795 0 -1 3286
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1707688321
transform 1 0 797 0 -1 1452
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1707688321
transform 1 0 797 0 -1 1786
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1707688321
transform 1 0 797 0 1 10
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_9
timestamp 1707688321
transform 1 0 797 0 1 976
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_10
timestamp 1707688321
transform 1 0 797 0 1 1310
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_11
timestamp 1707688321
transform 1 0 797 0 1 534
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_12
timestamp 1707688321
transform 1 0 797 0 1 868
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_13
timestamp 1707688321
transform 1 0 797 0 1 92
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_14
timestamp 1707688321
transform 1 0 797 0 1 426
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1707688321
transform 0 -1 370 -1 0 4112
box 0 0 1 1
use PYbentRes_CDNS_5246887918563  PYbentRes_CDNS_5246887918563_0
timestamp 1707688321
transform 0 1 512 -1 0 3748
box -50 0 1250 160
use PYbentRes_CDNS_5246887918563  PYbentRes_CDNS_5246887918563_1
timestamp 1707688321
transform 0 1 770 -1 0 3748
box -50 0 1250 160
use PYbentRes_CDNS_524688791851509  PYbentRes_CDNS_524688791851509_0
timestamp 1707688321
transform 0 -1 1186 -1 0 3748
box -50 -768 2523 160
use PYbentRes_CDNS_524688791851510  PYbentRes_CDNS_524688791851510_0
timestamp 1707688321
transform 0 -1 160 -1 0 3748
box -50 -256 1232 160
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1707688321
transform 0 1 783 1 0 4
box 0 0 1 1
use PYres_CDNS_5246887918567  PYres_CDNS_5246887918567_0
timestamp 1707688321
transform 0 1 770 -1 0 1752
box -50 0 350 160
use PYres_CDNS_5246887918567  PYres_CDNS_5246887918567_1
timestamp 1707688321
transform 0 1 770 -1 0 1310
box -50 0 350 160
use PYres_CDNS_5246887918567  PYres_CDNS_5246887918567_2
timestamp 1707688321
transform 0 1 770 -1 0 868
box -50 0 350 160
use PYres_CDNS_5246887918567  PYres_CDNS_5246887918567_3
timestamp 1707688321
transform 0 1 770 -1 0 426
box -50 0 350 160
use sky130_fd_io__tk_em1o_CDNS_524688791851507  sky130_fd_io__tk_em1o_CDNS_524688791851507_0
timestamp 1707688321
transform 0 1 525 1 0 3075
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851508  sky130_fd_io__tk_em1s_CDNS_524688791851508_0
timestamp 1707688321
transform 0 -1 915 -1 0 3221
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851508  sky130_fd_io__tk_em1s_CDNS_524688791851508_1
timestamp 1707688321
transform 0 1 785 -1 0 1677
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851508  sky130_fd_io__tk_em1s_CDNS_524688791851508_2
timestamp 1707688321
transform 0 1 785 -1 0 1214
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851508  sky130_fd_io__tk_em1s_CDNS_524688791851508_3
timestamp 1707688321
transform 0 1 785 -1 0 789
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851508  sky130_fd_io__tk_em1s_CDNS_524688791851508_4
timestamp 1707688321
transform 0 1 785 -1 0 345
box 0 0 1 1
<< labels >>
flabel comment s 848 1773 848 1773 0 FreeSans 100 0 0 0 n<0>
<< properties >>
string GDS_END 90834894
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 90831108
<< end >>
