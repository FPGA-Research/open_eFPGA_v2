magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -36 18142 1876 18781
rect -36 15902 1876 17066
rect -36 13662 1876 14826
rect -36 11422 1876 12586
rect -36 9182 1876 10346
rect 2576 7127 3494 7805
rect 2576 6335 4258 7127
rect 2576 4185 4306 4977
rect 2576 3507 3394 4185
rect 2576 1471 3762 2149
rect 1168 1467 1976 1471
rect -8 679 1976 1467
rect 2576 679 4306 1471
rect -8 676 1176 679
<< pwell >>
rect 34 17753 136 17763
rect 402 17753 504 17763
rect 770 17753 872 17763
rect 1138 17753 1240 17763
rect 1506 17753 1608 17763
rect 34 17455 1812 17753
rect 34 17445 136 17455
rect 402 17445 504 17455
rect 770 17445 872 17455
rect 1138 17445 1240 17455
rect 1506 17445 1608 17455
rect 34 15513 136 15523
rect 402 15513 504 15523
rect 770 15513 872 15523
rect 1138 15513 1240 15523
rect 1506 15513 1608 15523
rect 34 15215 1812 15513
rect 34 15205 136 15215
rect 402 15205 504 15215
rect 770 15205 872 15215
rect 1138 15205 1240 15215
rect 1506 15205 1608 15215
rect 34 13273 136 13283
rect 402 13273 504 13283
rect 770 13273 872 13283
rect 1138 13273 1240 13283
rect 1506 13273 1608 13283
rect 34 12975 1812 13273
rect 34 12965 136 12975
rect 402 12965 504 12975
rect 770 12965 872 12975
rect 1138 12965 1240 12975
rect 1506 12965 1608 12975
rect 34 11033 136 11043
rect 402 11033 504 11043
rect 770 11033 872 11043
rect 1138 11033 1240 11043
rect 1506 11033 1608 11043
rect 34 10735 1812 11033
rect 34 10725 136 10735
rect 402 10725 504 10735
rect 770 10725 872 10735
rect 1138 10725 1240 10735
rect 1506 10725 1608 10735
rect 34 8793 136 8803
rect 402 8793 504 8803
rect 770 8793 872 8803
rect 1138 8793 1240 8803
rect 1506 8793 1608 8803
rect 34 8669 1812 8793
rect 2640 8325 3424 8459
rect 2640 8259 3320 8325
rect 3118 8007 3320 8259
rect 3992 5985 4194 6133
rect 3734 5881 4194 5985
rect 2640 5832 2942 5881
rect 2640 5805 3046 5832
rect 3476 5815 4194 5881
rect 3312 5805 4194 5815
rect 2640 5631 4194 5805
rect 2640 5507 4242 5631
rect 2844 5480 4242 5507
rect 3008 5431 4242 5480
rect 3524 5243 4242 5431
rect 3524 5179 3726 5243
rect 4040 5179 4242 5243
rect 3018 3053 3220 3241
rect 2640 2987 3220 3053
rect 2640 2803 3324 2987
rect 2640 2679 3692 2803
rect 2844 2669 3692 2679
rect 3008 2603 3588 2669
rect 3386 2415 3588 2603
rect 3782 413 4242 477
rect 2 225 1166 328
rect 1600 225 1802 413
rect 3524 329 4242 413
rect 2 159 1802 225
rect 2 25 1906 159
rect 2844 149 2946 159
rect 3266 149 4242 329
rect 2640 25 4242 149
rect 2 -43 1088 25
<< scnmos >>
rect 224 17655 254 17727
rect 592 17655 622 17727
rect 960 17655 990 17727
rect 1328 17655 1358 17727
rect 1696 17655 1726 17727
rect 224 17481 254 17553
rect 592 17481 622 17553
rect 960 17481 990 17553
rect 1328 17481 1358 17553
rect 1696 17481 1726 17553
rect 224 15415 254 15487
rect 592 15415 622 15487
rect 960 15415 990 15487
rect 1328 15415 1358 15487
rect 1696 15415 1726 15487
rect 224 15241 254 15313
rect 592 15241 622 15313
rect 960 15241 990 15313
rect 1328 15241 1358 15313
rect 1696 15241 1726 15313
rect 224 13175 254 13247
rect 592 13175 622 13247
rect 960 13175 990 13247
rect 1328 13175 1358 13247
rect 1696 13175 1726 13247
rect 224 13001 254 13073
rect 592 13001 622 13073
rect 960 13001 990 13073
rect 1328 13001 1358 13073
rect 1696 13001 1726 13073
rect 224 10935 254 11007
rect 592 10935 622 11007
rect 960 10935 990 11007
rect 1328 10935 1358 11007
rect 1696 10935 1726 11007
rect 224 10761 254 10833
rect 592 10761 622 10833
rect 960 10761 990 10833
rect 1328 10761 1358 10833
rect 1696 10761 1726 10833
rect 224 8695 254 8767
rect 592 8695 622 8767
rect 960 8695 990 8767
rect 1328 8695 1358 8767
rect 1696 8695 1726 8767
rect 2726 8285 2756 8433
rect 2826 8285 2856 8433
rect 2926 8285 2956 8433
rect 3204 8033 3234 8433
rect 2726 5707 2756 5855
rect 2826 5707 2856 5855
rect 3194 5707 3224 5779
rect 3562 5707 3592 5855
rect 3820 5707 3850 5959
rect 4078 5707 4108 6107
rect 2726 5533 2756 5605
rect 3094 5457 3124 5529
rect 3352 5457 3382 5605
rect 3610 5205 3640 5605
rect 3868 5269 3898 5605
rect 4126 5205 4156 5605
rect 2726 2879 2756 3027
rect 2826 2879 2856 3027
rect 3104 2879 3134 3215
rect 2726 2705 2756 2777
rect 3094 2629 3124 2777
rect 3194 2629 3224 2777
rect 3472 2441 3502 2777
rect 81 102 111 302
rect 167 102 197 302
rect 239 102 269 302
rect 359 102 389 302
rect 431 102 461 302
rect 517 102 547 302
rect 589 102 619 302
rect 709 102 739 302
rect 781 102 811 302
rect 867 102 897 302
rect 1057 102 1087 302
rect 1318 51 1348 199
rect 1686 51 1716 387
rect 2726 51 2756 123
rect 3094 51 3124 123
rect 3352 51 3382 303
rect 3610 51 3640 387
rect 3868 51 3898 451
rect 4126 51 4156 451
<< scpmos >>
rect 224 18449 254 18673
rect 592 18449 622 18673
rect 960 18449 990 18673
rect 1328 18449 1358 18673
rect 1696 18449 1726 18673
rect 224 16535 254 16759
rect 592 16535 622 16759
rect 960 16535 990 16759
rect 1328 16535 1358 16759
rect 1696 16535 1726 16759
rect 224 16209 254 16433
rect 592 16209 622 16433
rect 960 16209 990 16433
rect 1328 16209 1358 16433
rect 1696 16209 1726 16433
rect 224 14295 254 14519
rect 592 14295 622 14519
rect 960 14295 990 14519
rect 1328 14295 1358 14519
rect 1696 14295 1726 14519
rect 224 13969 254 14193
rect 592 13969 622 14193
rect 960 13969 990 14193
rect 1328 13969 1358 14193
rect 1696 13969 1726 14193
rect 224 12055 254 12279
rect 592 12055 622 12279
rect 960 12055 990 12279
rect 1328 12055 1358 12279
rect 1696 12055 1726 12279
rect 224 11729 254 11953
rect 592 11729 622 11953
rect 960 11729 990 11953
rect 1328 11729 1358 11953
rect 1696 11729 1726 11953
rect 224 9815 254 10039
rect 592 9815 622 10039
rect 960 9815 990 10039
rect 1328 9815 1358 10039
rect 1696 9815 1726 10039
rect 224 9489 254 9713
rect 592 9489 622 9713
rect 960 9489 990 9713
rect 1328 9489 1358 9713
rect 1696 9489 1726 9713
rect 2726 7121 2756 7345
rect 2826 7121 2856 7345
rect 2926 7121 2956 7345
rect 3204 7121 3234 7521
rect 2726 6795 2756 7019
rect 2826 6795 2856 7019
rect 3194 6795 3224 7019
rect 3562 6795 3592 7019
rect 3820 6619 3850 7019
rect 4078 6619 4108 7019
rect 2726 4293 2756 4517
rect 3094 4293 3124 4517
rect 3352 4293 3382 4517
rect 3610 4293 3640 4693
rect 3868 4293 3898 4693
rect 4126 4293 4156 4693
rect 2726 3967 2756 4191
rect 2826 3967 2856 4191
rect 3104 3791 3134 4191
rect 2726 1465 2756 1689
rect 3094 1465 3124 1689
rect 3194 1465 3224 1689
rect 3472 1465 3502 1865
rect 81 712 111 1312
rect 167 712 197 1312
rect 239 712 269 1312
rect 359 712 389 1312
rect 431 712 461 1312
rect 517 712 547 1312
rect 589 712 619 1312
rect 709 712 739 1312
rect 781 712 811 1312
rect 867 712 897 1312
rect 1057 712 1087 1312
rect 1318 1139 1348 1363
rect 1686 1033 1716 1363
rect 2726 1139 2756 1363
rect 3094 1139 3124 1363
rect 3352 1033 3382 1363
rect 3610 963 3640 1363
rect 3868 963 3898 1363
rect 4126 963 4156 1363
<< ndiff >>
rect 164 17708 224 17727
rect 164 17674 172 17708
rect 206 17674 224 17708
rect 164 17655 224 17674
rect 254 17708 314 17727
rect 254 17674 272 17708
rect 306 17674 314 17708
rect 254 17655 314 17674
rect 532 17708 592 17727
rect 532 17674 540 17708
rect 574 17674 592 17708
rect 532 17655 592 17674
rect 622 17708 682 17727
rect 622 17674 640 17708
rect 674 17674 682 17708
rect 622 17655 682 17674
rect 900 17708 960 17727
rect 900 17674 908 17708
rect 942 17674 960 17708
rect 900 17655 960 17674
rect 990 17708 1050 17727
rect 990 17674 1008 17708
rect 1042 17674 1050 17708
rect 990 17655 1050 17674
rect 1268 17708 1328 17727
rect 1268 17674 1276 17708
rect 1310 17674 1328 17708
rect 1268 17655 1328 17674
rect 1358 17708 1418 17727
rect 1358 17674 1376 17708
rect 1410 17674 1418 17708
rect 1358 17655 1418 17674
rect 1636 17708 1696 17727
rect 1636 17674 1644 17708
rect 1678 17674 1696 17708
rect 1636 17655 1696 17674
rect 1726 17708 1786 17727
rect 1726 17674 1744 17708
rect 1778 17674 1786 17708
rect 1726 17655 1786 17674
rect 164 17534 224 17553
rect 164 17500 172 17534
rect 206 17500 224 17534
rect 164 17481 224 17500
rect 254 17534 314 17553
rect 254 17500 272 17534
rect 306 17500 314 17534
rect 254 17481 314 17500
rect 532 17534 592 17553
rect 532 17500 540 17534
rect 574 17500 592 17534
rect 532 17481 592 17500
rect 622 17534 682 17553
rect 622 17500 640 17534
rect 674 17500 682 17534
rect 622 17481 682 17500
rect 900 17534 960 17553
rect 900 17500 908 17534
rect 942 17500 960 17534
rect 900 17481 960 17500
rect 990 17534 1050 17553
rect 990 17500 1008 17534
rect 1042 17500 1050 17534
rect 990 17481 1050 17500
rect 1268 17534 1328 17553
rect 1268 17500 1276 17534
rect 1310 17500 1328 17534
rect 1268 17481 1328 17500
rect 1358 17534 1418 17553
rect 1358 17500 1376 17534
rect 1410 17500 1418 17534
rect 1358 17481 1418 17500
rect 1636 17534 1696 17553
rect 1636 17500 1644 17534
rect 1678 17500 1696 17534
rect 1636 17481 1696 17500
rect 1726 17534 1786 17553
rect 1726 17500 1744 17534
rect 1778 17500 1786 17534
rect 1726 17481 1786 17500
rect 164 15468 224 15487
rect 164 15434 172 15468
rect 206 15434 224 15468
rect 164 15415 224 15434
rect 254 15468 314 15487
rect 254 15434 272 15468
rect 306 15434 314 15468
rect 254 15415 314 15434
rect 532 15468 592 15487
rect 532 15434 540 15468
rect 574 15434 592 15468
rect 532 15415 592 15434
rect 622 15468 682 15487
rect 622 15434 640 15468
rect 674 15434 682 15468
rect 622 15415 682 15434
rect 900 15468 960 15487
rect 900 15434 908 15468
rect 942 15434 960 15468
rect 900 15415 960 15434
rect 990 15468 1050 15487
rect 990 15434 1008 15468
rect 1042 15434 1050 15468
rect 990 15415 1050 15434
rect 1268 15468 1328 15487
rect 1268 15434 1276 15468
rect 1310 15434 1328 15468
rect 1268 15415 1328 15434
rect 1358 15468 1418 15487
rect 1358 15434 1376 15468
rect 1410 15434 1418 15468
rect 1358 15415 1418 15434
rect 1636 15468 1696 15487
rect 1636 15434 1644 15468
rect 1678 15434 1696 15468
rect 1636 15415 1696 15434
rect 1726 15468 1786 15487
rect 1726 15434 1744 15468
rect 1778 15434 1786 15468
rect 1726 15415 1786 15434
rect 164 15294 224 15313
rect 164 15260 172 15294
rect 206 15260 224 15294
rect 164 15241 224 15260
rect 254 15294 314 15313
rect 254 15260 272 15294
rect 306 15260 314 15294
rect 254 15241 314 15260
rect 532 15294 592 15313
rect 532 15260 540 15294
rect 574 15260 592 15294
rect 532 15241 592 15260
rect 622 15294 682 15313
rect 622 15260 640 15294
rect 674 15260 682 15294
rect 622 15241 682 15260
rect 900 15294 960 15313
rect 900 15260 908 15294
rect 942 15260 960 15294
rect 900 15241 960 15260
rect 990 15294 1050 15313
rect 990 15260 1008 15294
rect 1042 15260 1050 15294
rect 990 15241 1050 15260
rect 1268 15294 1328 15313
rect 1268 15260 1276 15294
rect 1310 15260 1328 15294
rect 1268 15241 1328 15260
rect 1358 15294 1418 15313
rect 1358 15260 1376 15294
rect 1410 15260 1418 15294
rect 1358 15241 1418 15260
rect 1636 15294 1696 15313
rect 1636 15260 1644 15294
rect 1678 15260 1696 15294
rect 1636 15241 1696 15260
rect 1726 15294 1786 15313
rect 1726 15260 1744 15294
rect 1778 15260 1786 15294
rect 1726 15241 1786 15260
rect 164 13228 224 13247
rect 164 13194 172 13228
rect 206 13194 224 13228
rect 164 13175 224 13194
rect 254 13228 314 13247
rect 254 13194 272 13228
rect 306 13194 314 13228
rect 254 13175 314 13194
rect 532 13228 592 13247
rect 532 13194 540 13228
rect 574 13194 592 13228
rect 532 13175 592 13194
rect 622 13228 682 13247
rect 622 13194 640 13228
rect 674 13194 682 13228
rect 622 13175 682 13194
rect 900 13228 960 13247
rect 900 13194 908 13228
rect 942 13194 960 13228
rect 900 13175 960 13194
rect 990 13228 1050 13247
rect 990 13194 1008 13228
rect 1042 13194 1050 13228
rect 990 13175 1050 13194
rect 1268 13228 1328 13247
rect 1268 13194 1276 13228
rect 1310 13194 1328 13228
rect 1268 13175 1328 13194
rect 1358 13228 1418 13247
rect 1358 13194 1376 13228
rect 1410 13194 1418 13228
rect 1358 13175 1418 13194
rect 1636 13228 1696 13247
rect 1636 13194 1644 13228
rect 1678 13194 1696 13228
rect 1636 13175 1696 13194
rect 1726 13228 1786 13247
rect 1726 13194 1744 13228
rect 1778 13194 1786 13228
rect 1726 13175 1786 13194
rect 164 13054 224 13073
rect 164 13020 172 13054
rect 206 13020 224 13054
rect 164 13001 224 13020
rect 254 13054 314 13073
rect 254 13020 272 13054
rect 306 13020 314 13054
rect 254 13001 314 13020
rect 532 13054 592 13073
rect 532 13020 540 13054
rect 574 13020 592 13054
rect 532 13001 592 13020
rect 622 13054 682 13073
rect 622 13020 640 13054
rect 674 13020 682 13054
rect 622 13001 682 13020
rect 900 13054 960 13073
rect 900 13020 908 13054
rect 942 13020 960 13054
rect 900 13001 960 13020
rect 990 13054 1050 13073
rect 990 13020 1008 13054
rect 1042 13020 1050 13054
rect 990 13001 1050 13020
rect 1268 13054 1328 13073
rect 1268 13020 1276 13054
rect 1310 13020 1328 13054
rect 1268 13001 1328 13020
rect 1358 13054 1418 13073
rect 1358 13020 1376 13054
rect 1410 13020 1418 13054
rect 1358 13001 1418 13020
rect 1636 13054 1696 13073
rect 1636 13020 1644 13054
rect 1678 13020 1696 13054
rect 1636 13001 1696 13020
rect 1726 13054 1786 13073
rect 1726 13020 1744 13054
rect 1778 13020 1786 13054
rect 1726 13001 1786 13020
rect 164 10988 224 11007
rect 164 10954 172 10988
rect 206 10954 224 10988
rect 164 10935 224 10954
rect 254 10988 314 11007
rect 254 10954 272 10988
rect 306 10954 314 10988
rect 254 10935 314 10954
rect 532 10988 592 11007
rect 532 10954 540 10988
rect 574 10954 592 10988
rect 532 10935 592 10954
rect 622 10988 682 11007
rect 622 10954 640 10988
rect 674 10954 682 10988
rect 622 10935 682 10954
rect 900 10988 960 11007
rect 900 10954 908 10988
rect 942 10954 960 10988
rect 900 10935 960 10954
rect 990 10988 1050 11007
rect 990 10954 1008 10988
rect 1042 10954 1050 10988
rect 990 10935 1050 10954
rect 1268 10988 1328 11007
rect 1268 10954 1276 10988
rect 1310 10954 1328 10988
rect 1268 10935 1328 10954
rect 1358 10988 1418 11007
rect 1358 10954 1376 10988
rect 1410 10954 1418 10988
rect 1358 10935 1418 10954
rect 1636 10988 1696 11007
rect 1636 10954 1644 10988
rect 1678 10954 1696 10988
rect 1636 10935 1696 10954
rect 1726 10988 1786 11007
rect 1726 10954 1744 10988
rect 1778 10954 1786 10988
rect 1726 10935 1786 10954
rect 164 10814 224 10833
rect 164 10780 172 10814
rect 206 10780 224 10814
rect 164 10761 224 10780
rect 254 10814 314 10833
rect 254 10780 272 10814
rect 306 10780 314 10814
rect 254 10761 314 10780
rect 532 10814 592 10833
rect 532 10780 540 10814
rect 574 10780 592 10814
rect 532 10761 592 10780
rect 622 10814 682 10833
rect 622 10780 640 10814
rect 674 10780 682 10814
rect 622 10761 682 10780
rect 900 10814 960 10833
rect 900 10780 908 10814
rect 942 10780 960 10814
rect 900 10761 960 10780
rect 990 10814 1050 10833
rect 990 10780 1008 10814
rect 1042 10780 1050 10814
rect 990 10761 1050 10780
rect 1268 10814 1328 10833
rect 1268 10780 1276 10814
rect 1310 10780 1328 10814
rect 1268 10761 1328 10780
rect 1358 10814 1418 10833
rect 1358 10780 1376 10814
rect 1410 10780 1418 10814
rect 1358 10761 1418 10780
rect 1636 10814 1696 10833
rect 1636 10780 1644 10814
rect 1678 10780 1696 10814
rect 1636 10761 1696 10780
rect 1726 10814 1786 10833
rect 1726 10780 1744 10814
rect 1778 10780 1786 10814
rect 1726 10761 1786 10780
rect 164 8748 224 8767
rect 164 8714 172 8748
rect 206 8714 224 8748
rect 164 8695 224 8714
rect 254 8748 314 8767
rect 254 8714 272 8748
rect 306 8714 314 8748
rect 254 8695 314 8714
rect 532 8748 592 8767
rect 532 8714 540 8748
rect 574 8714 592 8748
rect 532 8695 592 8714
rect 622 8748 682 8767
rect 622 8714 640 8748
rect 674 8714 682 8748
rect 622 8695 682 8714
rect 900 8748 960 8767
rect 900 8714 908 8748
rect 942 8714 960 8748
rect 900 8695 960 8714
rect 990 8748 1050 8767
rect 990 8714 1008 8748
rect 1042 8714 1050 8748
rect 990 8695 1050 8714
rect 1268 8748 1328 8767
rect 1268 8714 1276 8748
rect 1310 8714 1328 8748
rect 1268 8695 1328 8714
rect 1358 8748 1418 8767
rect 1358 8714 1376 8748
rect 1410 8714 1418 8748
rect 1358 8695 1418 8714
rect 1636 8748 1696 8767
rect 1636 8714 1644 8748
rect 1678 8714 1696 8748
rect 1636 8695 1696 8714
rect 1726 8748 1786 8767
rect 1726 8714 1744 8748
rect 1778 8714 1786 8748
rect 1726 8695 1786 8714
rect 2666 8376 2726 8433
rect 2666 8342 2674 8376
rect 2708 8342 2726 8376
rect 2666 8285 2726 8342
rect 2756 8285 2826 8433
rect 2856 8285 2926 8433
rect 2956 8376 3016 8433
rect 2956 8342 2974 8376
rect 3008 8342 3016 8376
rect 2956 8285 3016 8342
rect 3144 8250 3204 8433
rect 3144 8216 3152 8250
rect 3186 8216 3204 8250
rect 3144 8033 3204 8216
rect 3234 8250 3294 8433
rect 3234 8216 3252 8250
rect 3286 8216 3294 8250
rect 3234 8033 3294 8216
rect 2666 5798 2726 5855
rect 2666 5764 2674 5798
rect 2708 5764 2726 5798
rect 2666 5707 2726 5764
rect 2756 5707 2826 5855
rect 2856 5798 2916 5855
rect 2856 5764 2874 5798
rect 2908 5764 2916 5798
rect 2856 5707 2916 5764
rect 3502 5798 3562 5855
rect 3134 5760 3194 5779
rect 3134 5726 3142 5760
rect 3176 5726 3194 5760
rect 3134 5707 3194 5726
rect 3224 5760 3284 5779
rect 3224 5726 3242 5760
rect 3276 5726 3284 5760
rect 3224 5707 3284 5726
rect 3502 5764 3510 5798
rect 3544 5764 3562 5798
rect 3502 5707 3562 5764
rect 3592 5798 3652 5855
rect 3592 5764 3610 5798
rect 3644 5764 3652 5798
rect 3592 5707 3652 5764
rect 3760 5850 3820 5959
rect 3760 5816 3768 5850
rect 3802 5816 3820 5850
rect 3760 5707 3820 5816
rect 3850 5850 3910 5959
rect 3850 5816 3868 5850
rect 3902 5816 3910 5850
rect 3850 5707 3910 5816
rect 4018 5924 4078 6107
rect 4018 5890 4026 5924
rect 4060 5890 4078 5924
rect 4018 5707 4078 5890
rect 4108 5924 4168 6107
rect 4108 5890 4126 5924
rect 4160 5890 4168 5924
rect 4108 5707 4168 5890
rect 2666 5586 2726 5605
rect 2666 5552 2674 5586
rect 2708 5552 2726 5586
rect 2666 5533 2726 5552
rect 2756 5586 2816 5605
rect 2756 5552 2774 5586
rect 2808 5552 2816 5586
rect 2756 5533 2816 5552
rect 3292 5548 3352 5605
rect 3034 5510 3094 5529
rect 3034 5476 3042 5510
rect 3076 5476 3094 5510
rect 3034 5457 3094 5476
rect 3124 5510 3184 5529
rect 3124 5476 3142 5510
rect 3176 5476 3184 5510
rect 3124 5457 3184 5476
rect 3292 5514 3300 5548
rect 3334 5514 3352 5548
rect 3292 5457 3352 5514
rect 3382 5548 3442 5605
rect 3382 5514 3400 5548
rect 3434 5514 3442 5548
rect 3382 5457 3442 5514
rect 3550 5422 3610 5605
rect 3550 5388 3558 5422
rect 3592 5388 3610 5422
rect 3550 5205 3610 5388
rect 3640 5422 3700 5605
rect 3640 5388 3658 5422
rect 3692 5388 3700 5422
rect 3640 5205 3700 5388
rect 3808 5454 3868 5605
rect 3808 5420 3816 5454
rect 3850 5420 3868 5454
rect 3808 5269 3868 5420
rect 3898 5454 3958 5605
rect 3898 5420 3916 5454
rect 3950 5420 3958 5454
rect 3898 5269 3958 5420
rect 4066 5422 4126 5605
rect 4066 5388 4074 5422
rect 4108 5388 4126 5422
rect 4066 5205 4126 5388
rect 4156 5422 4216 5605
rect 4156 5388 4174 5422
rect 4208 5388 4216 5422
rect 4156 5205 4216 5388
rect 3044 3064 3104 3215
rect 3044 3030 3052 3064
rect 3086 3030 3104 3064
rect 2666 2970 2726 3027
rect 2666 2936 2674 2970
rect 2708 2936 2726 2970
rect 2666 2879 2726 2936
rect 2756 2879 2826 3027
rect 2856 2970 2916 3027
rect 2856 2936 2874 2970
rect 2908 2936 2916 2970
rect 2856 2879 2916 2936
rect 3044 2879 3104 3030
rect 3134 3064 3194 3215
rect 3134 3030 3152 3064
rect 3186 3030 3194 3064
rect 3134 2879 3194 3030
rect 2666 2758 2726 2777
rect 2666 2724 2674 2758
rect 2708 2724 2726 2758
rect 2666 2705 2726 2724
rect 2756 2758 2816 2777
rect 2756 2724 2774 2758
rect 2808 2724 2816 2758
rect 2756 2705 2816 2724
rect 3034 2720 3094 2777
rect 3034 2686 3042 2720
rect 3076 2686 3094 2720
rect 3034 2629 3094 2686
rect 3124 2629 3194 2777
rect 3224 2720 3284 2777
rect 3224 2686 3242 2720
rect 3276 2686 3284 2720
rect 3224 2629 3284 2686
rect 3412 2626 3472 2777
rect 3412 2592 3420 2626
rect 3454 2592 3472 2626
rect 3412 2441 3472 2592
rect 3502 2626 3562 2777
rect 3502 2592 3520 2626
rect 3554 2592 3562 2626
rect 3502 2441 3562 2592
rect 28 237 81 302
rect 28 203 36 237
rect 70 203 81 237
rect 28 169 81 203
rect 28 135 36 169
rect 70 135 81 169
rect 28 102 81 135
rect 111 237 167 302
rect 111 203 122 237
rect 156 203 167 237
rect 111 169 167 203
rect 111 135 122 169
rect 156 135 167 169
rect 111 102 167 135
rect 197 102 239 302
rect 269 237 359 302
rect 269 203 297 237
rect 331 203 359 237
rect 269 169 359 203
rect 269 135 297 169
rect 331 135 359 169
rect 269 102 359 135
rect 389 102 431 302
rect 461 237 517 302
rect 461 203 472 237
rect 506 203 517 237
rect 461 169 517 203
rect 461 135 472 169
rect 506 135 517 169
rect 461 102 517 135
rect 547 102 589 302
rect 619 237 709 302
rect 619 203 647 237
rect 681 203 709 237
rect 619 169 709 203
rect 619 135 647 169
rect 681 135 709 169
rect 619 102 709 135
rect 739 102 781 302
rect 811 237 867 302
rect 811 203 822 237
rect 856 203 867 237
rect 811 169 867 203
rect 811 135 822 169
rect 856 135 867 169
rect 811 102 867 135
rect 897 237 950 302
rect 897 203 908 237
rect 942 203 950 237
rect 897 169 950 203
rect 897 135 908 169
rect 942 135 950 169
rect 897 102 950 135
rect 1004 237 1057 302
rect 1004 203 1012 237
rect 1046 203 1057 237
rect 1004 169 1057 203
rect 1004 135 1012 169
rect 1046 135 1057 169
rect 1004 102 1057 135
rect 1087 237 1140 302
rect 1087 203 1098 237
rect 1132 203 1140 237
rect 1087 169 1140 203
rect 1626 236 1686 387
rect 1626 202 1634 236
rect 1668 202 1686 236
rect 1087 135 1098 169
rect 1132 135 1140 169
rect 1087 102 1140 135
rect 1258 142 1318 199
rect 1258 108 1266 142
rect 1300 108 1318 142
rect 1258 51 1318 108
rect 1348 142 1408 199
rect 1348 108 1366 142
rect 1400 108 1408 142
rect 1348 51 1408 108
rect 1626 51 1686 202
rect 1716 236 1776 387
rect 1716 202 1734 236
rect 1768 202 1776 236
rect 1716 51 1776 202
rect 2666 104 2726 123
rect 2666 70 2674 104
rect 2708 70 2726 104
rect 2666 51 2726 70
rect 2756 104 2816 123
rect 2756 70 2774 104
rect 2808 70 2816 104
rect 2756 51 2816 70
rect 3292 194 3352 303
rect 3292 160 3300 194
rect 3334 160 3352 194
rect 3034 104 3094 123
rect 3034 70 3042 104
rect 3076 70 3094 104
rect 3034 51 3094 70
rect 3124 104 3184 123
rect 3124 70 3142 104
rect 3176 70 3184 104
rect 3124 51 3184 70
rect 3292 51 3352 160
rect 3382 194 3442 303
rect 3382 160 3400 194
rect 3434 160 3442 194
rect 3382 51 3442 160
rect 3550 236 3610 387
rect 3550 202 3558 236
rect 3592 202 3610 236
rect 3550 51 3610 202
rect 3640 236 3700 387
rect 3640 202 3658 236
rect 3692 202 3700 236
rect 3640 51 3700 202
rect 3808 268 3868 451
rect 3808 234 3816 268
rect 3850 234 3868 268
rect 3808 51 3868 234
rect 3898 268 3958 451
rect 3898 234 3916 268
rect 3950 234 3958 268
rect 3898 51 3958 234
rect 4066 268 4126 451
rect 4066 234 4074 268
rect 4108 234 4126 268
rect 4066 51 4126 234
rect 4156 268 4216 451
rect 4156 234 4174 268
rect 4208 234 4216 268
rect 4156 51 4216 234
<< pdiff >>
rect 164 18578 224 18673
rect 164 18544 172 18578
rect 206 18544 224 18578
rect 164 18449 224 18544
rect 254 18578 314 18673
rect 254 18544 272 18578
rect 306 18544 314 18578
rect 254 18449 314 18544
rect 532 18578 592 18673
rect 532 18544 540 18578
rect 574 18544 592 18578
rect 532 18449 592 18544
rect 622 18578 682 18673
rect 622 18544 640 18578
rect 674 18544 682 18578
rect 622 18449 682 18544
rect 900 18578 960 18673
rect 900 18544 908 18578
rect 942 18544 960 18578
rect 900 18449 960 18544
rect 990 18578 1050 18673
rect 990 18544 1008 18578
rect 1042 18544 1050 18578
rect 990 18449 1050 18544
rect 1268 18578 1328 18673
rect 1268 18544 1276 18578
rect 1310 18544 1328 18578
rect 1268 18449 1328 18544
rect 1358 18578 1418 18673
rect 1358 18544 1376 18578
rect 1410 18544 1418 18578
rect 1358 18449 1418 18544
rect 1636 18578 1696 18673
rect 1636 18544 1644 18578
rect 1678 18544 1696 18578
rect 1636 18449 1696 18544
rect 1726 18578 1786 18673
rect 1726 18544 1744 18578
rect 1778 18544 1786 18578
rect 1726 18449 1786 18544
rect 164 16664 224 16759
rect 164 16630 172 16664
rect 206 16630 224 16664
rect 164 16535 224 16630
rect 254 16664 314 16759
rect 254 16630 272 16664
rect 306 16630 314 16664
rect 254 16535 314 16630
rect 532 16664 592 16759
rect 532 16630 540 16664
rect 574 16630 592 16664
rect 532 16535 592 16630
rect 622 16664 682 16759
rect 622 16630 640 16664
rect 674 16630 682 16664
rect 622 16535 682 16630
rect 900 16664 960 16759
rect 900 16630 908 16664
rect 942 16630 960 16664
rect 900 16535 960 16630
rect 990 16664 1050 16759
rect 990 16630 1008 16664
rect 1042 16630 1050 16664
rect 990 16535 1050 16630
rect 1268 16664 1328 16759
rect 1268 16630 1276 16664
rect 1310 16630 1328 16664
rect 1268 16535 1328 16630
rect 1358 16664 1418 16759
rect 1358 16630 1376 16664
rect 1410 16630 1418 16664
rect 1358 16535 1418 16630
rect 1636 16664 1696 16759
rect 1636 16630 1644 16664
rect 1678 16630 1696 16664
rect 1636 16535 1696 16630
rect 1726 16664 1786 16759
rect 1726 16630 1744 16664
rect 1778 16630 1786 16664
rect 1726 16535 1786 16630
rect 164 16338 224 16433
rect 164 16304 172 16338
rect 206 16304 224 16338
rect 164 16209 224 16304
rect 254 16338 314 16433
rect 254 16304 272 16338
rect 306 16304 314 16338
rect 254 16209 314 16304
rect 532 16338 592 16433
rect 532 16304 540 16338
rect 574 16304 592 16338
rect 532 16209 592 16304
rect 622 16338 682 16433
rect 622 16304 640 16338
rect 674 16304 682 16338
rect 622 16209 682 16304
rect 900 16338 960 16433
rect 900 16304 908 16338
rect 942 16304 960 16338
rect 900 16209 960 16304
rect 990 16338 1050 16433
rect 990 16304 1008 16338
rect 1042 16304 1050 16338
rect 990 16209 1050 16304
rect 1268 16338 1328 16433
rect 1268 16304 1276 16338
rect 1310 16304 1328 16338
rect 1268 16209 1328 16304
rect 1358 16338 1418 16433
rect 1358 16304 1376 16338
rect 1410 16304 1418 16338
rect 1358 16209 1418 16304
rect 1636 16338 1696 16433
rect 1636 16304 1644 16338
rect 1678 16304 1696 16338
rect 1636 16209 1696 16304
rect 1726 16338 1786 16433
rect 1726 16304 1744 16338
rect 1778 16304 1786 16338
rect 1726 16209 1786 16304
rect 164 14424 224 14519
rect 164 14390 172 14424
rect 206 14390 224 14424
rect 164 14295 224 14390
rect 254 14424 314 14519
rect 254 14390 272 14424
rect 306 14390 314 14424
rect 254 14295 314 14390
rect 532 14424 592 14519
rect 532 14390 540 14424
rect 574 14390 592 14424
rect 532 14295 592 14390
rect 622 14424 682 14519
rect 622 14390 640 14424
rect 674 14390 682 14424
rect 622 14295 682 14390
rect 900 14424 960 14519
rect 900 14390 908 14424
rect 942 14390 960 14424
rect 900 14295 960 14390
rect 990 14424 1050 14519
rect 990 14390 1008 14424
rect 1042 14390 1050 14424
rect 990 14295 1050 14390
rect 1268 14424 1328 14519
rect 1268 14390 1276 14424
rect 1310 14390 1328 14424
rect 1268 14295 1328 14390
rect 1358 14424 1418 14519
rect 1358 14390 1376 14424
rect 1410 14390 1418 14424
rect 1358 14295 1418 14390
rect 1636 14424 1696 14519
rect 1636 14390 1644 14424
rect 1678 14390 1696 14424
rect 1636 14295 1696 14390
rect 1726 14424 1786 14519
rect 1726 14390 1744 14424
rect 1778 14390 1786 14424
rect 1726 14295 1786 14390
rect 164 14098 224 14193
rect 164 14064 172 14098
rect 206 14064 224 14098
rect 164 13969 224 14064
rect 254 14098 314 14193
rect 254 14064 272 14098
rect 306 14064 314 14098
rect 254 13969 314 14064
rect 532 14098 592 14193
rect 532 14064 540 14098
rect 574 14064 592 14098
rect 532 13969 592 14064
rect 622 14098 682 14193
rect 622 14064 640 14098
rect 674 14064 682 14098
rect 622 13969 682 14064
rect 900 14098 960 14193
rect 900 14064 908 14098
rect 942 14064 960 14098
rect 900 13969 960 14064
rect 990 14098 1050 14193
rect 990 14064 1008 14098
rect 1042 14064 1050 14098
rect 990 13969 1050 14064
rect 1268 14098 1328 14193
rect 1268 14064 1276 14098
rect 1310 14064 1328 14098
rect 1268 13969 1328 14064
rect 1358 14098 1418 14193
rect 1358 14064 1376 14098
rect 1410 14064 1418 14098
rect 1358 13969 1418 14064
rect 1636 14098 1696 14193
rect 1636 14064 1644 14098
rect 1678 14064 1696 14098
rect 1636 13969 1696 14064
rect 1726 14098 1786 14193
rect 1726 14064 1744 14098
rect 1778 14064 1786 14098
rect 1726 13969 1786 14064
rect 164 12184 224 12279
rect 164 12150 172 12184
rect 206 12150 224 12184
rect 164 12055 224 12150
rect 254 12184 314 12279
rect 254 12150 272 12184
rect 306 12150 314 12184
rect 254 12055 314 12150
rect 532 12184 592 12279
rect 532 12150 540 12184
rect 574 12150 592 12184
rect 532 12055 592 12150
rect 622 12184 682 12279
rect 622 12150 640 12184
rect 674 12150 682 12184
rect 622 12055 682 12150
rect 900 12184 960 12279
rect 900 12150 908 12184
rect 942 12150 960 12184
rect 900 12055 960 12150
rect 990 12184 1050 12279
rect 990 12150 1008 12184
rect 1042 12150 1050 12184
rect 990 12055 1050 12150
rect 1268 12184 1328 12279
rect 1268 12150 1276 12184
rect 1310 12150 1328 12184
rect 1268 12055 1328 12150
rect 1358 12184 1418 12279
rect 1358 12150 1376 12184
rect 1410 12150 1418 12184
rect 1358 12055 1418 12150
rect 1636 12184 1696 12279
rect 1636 12150 1644 12184
rect 1678 12150 1696 12184
rect 1636 12055 1696 12150
rect 1726 12184 1786 12279
rect 1726 12150 1744 12184
rect 1778 12150 1786 12184
rect 1726 12055 1786 12150
rect 164 11858 224 11953
rect 164 11824 172 11858
rect 206 11824 224 11858
rect 164 11729 224 11824
rect 254 11858 314 11953
rect 254 11824 272 11858
rect 306 11824 314 11858
rect 254 11729 314 11824
rect 532 11858 592 11953
rect 532 11824 540 11858
rect 574 11824 592 11858
rect 532 11729 592 11824
rect 622 11858 682 11953
rect 622 11824 640 11858
rect 674 11824 682 11858
rect 622 11729 682 11824
rect 900 11858 960 11953
rect 900 11824 908 11858
rect 942 11824 960 11858
rect 900 11729 960 11824
rect 990 11858 1050 11953
rect 990 11824 1008 11858
rect 1042 11824 1050 11858
rect 990 11729 1050 11824
rect 1268 11858 1328 11953
rect 1268 11824 1276 11858
rect 1310 11824 1328 11858
rect 1268 11729 1328 11824
rect 1358 11858 1418 11953
rect 1358 11824 1376 11858
rect 1410 11824 1418 11858
rect 1358 11729 1418 11824
rect 1636 11858 1696 11953
rect 1636 11824 1644 11858
rect 1678 11824 1696 11858
rect 1636 11729 1696 11824
rect 1726 11858 1786 11953
rect 1726 11824 1744 11858
rect 1778 11824 1786 11858
rect 1726 11729 1786 11824
rect 164 9944 224 10039
rect 164 9910 172 9944
rect 206 9910 224 9944
rect 164 9815 224 9910
rect 254 9944 314 10039
rect 254 9910 272 9944
rect 306 9910 314 9944
rect 254 9815 314 9910
rect 532 9944 592 10039
rect 532 9910 540 9944
rect 574 9910 592 9944
rect 532 9815 592 9910
rect 622 9944 682 10039
rect 622 9910 640 9944
rect 674 9910 682 9944
rect 622 9815 682 9910
rect 900 9944 960 10039
rect 900 9910 908 9944
rect 942 9910 960 9944
rect 900 9815 960 9910
rect 990 9944 1050 10039
rect 990 9910 1008 9944
rect 1042 9910 1050 9944
rect 990 9815 1050 9910
rect 1268 9944 1328 10039
rect 1268 9910 1276 9944
rect 1310 9910 1328 9944
rect 1268 9815 1328 9910
rect 1358 9944 1418 10039
rect 1358 9910 1376 9944
rect 1410 9910 1418 9944
rect 1358 9815 1418 9910
rect 1636 9944 1696 10039
rect 1636 9910 1644 9944
rect 1678 9910 1696 9944
rect 1636 9815 1696 9910
rect 1726 9944 1786 10039
rect 1726 9910 1744 9944
rect 1778 9910 1786 9944
rect 1726 9815 1786 9910
rect 164 9618 224 9713
rect 164 9584 172 9618
rect 206 9584 224 9618
rect 164 9489 224 9584
rect 254 9618 314 9713
rect 254 9584 272 9618
rect 306 9584 314 9618
rect 254 9489 314 9584
rect 532 9618 592 9713
rect 532 9584 540 9618
rect 574 9584 592 9618
rect 532 9489 592 9584
rect 622 9618 682 9713
rect 622 9584 640 9618
rect 674 9584 682 9618
rect 622 9489 682 9584
rect 900 9618 960 9713
rect 900 9584 908 9618
rect 942 9584 960 9618
rect 900 9489 960 9584
rect 990 9618 1050 9713
rect 990 9584 1008 9618
rect 1042 9584 1050 9618
rect 990 9489 1050 9584
rect 1268 9618 1328 9713
rect 1268 9584 1276 9618
rect 1310 9584 1328 9618
rect 1268 9489 1328 9584
rect 1358 9618 1418 9713
rect 1358 9584 1376 9618
rect 1410 9584 1418 9618
rect 1358 9489 1418 9584
rect 1636 9618 1696 9713
rect 1636 9584 1644 9618
rect 1678 9584 1696 9618
rect 1636 9489 1696 9584
rect 1726 9618 1786 9713
rect 1726 9584 1744 9618
rect 1778 9584 1786 9618
rect 1726 9489 1786 9584
rect 2666 7250 2726 7345
rect 2666 7216 2674 7250
rect 2708 7216 2726 7250
rect 2666 7121 2726 7216
rect 2756 7250 2826 7345
rect 2756 7216 2774 7250
rect 2808 7216 2826 7250
rect 2756 7121 2826 7216
rect 2856 7250 2926 7345
rect 2856 7216 2874 7250
rect 2908 7216 2926 7250
rect 2856 7121 2926 7216
rect 2956 7250 3016 7345
rect 2956 7216 2974 7250
rect 3008 7216 3016 7250
rect 2956 7121 3016 7216
rect 3144 7338 3204 7521
rect 3144 7304 3152 7338
rect 3186 7304 3204 7338
rect 3144 7121 3204 7304
rect 3234 7338 3294 7521
rect 3234 7304 3252 7338
rect 3286 7304 3294 7338
rect 3234 7121 3294 7304
rect 2666 6924 2726 7019
rect 2666 6890 2674 6924
rect 2708 6890 2726 6924
rect 2666 6795 2726 6890
rect 2756 6924 2826 7019
rect 2756 6890 2774 6924
rect 2808 6890 2826 6924
rect 2756 6795 2826 6890
rect 2856 6924 2916 7019
rect 2856 6890 2874 6924
rect 2908 6890 2916 6924
rect 2856 6795 2916 6890
rect 3134 6924 3194 7019
rect 3134 6890 3142 6924
rect 3176 6890 3194 6924
rect 3134 6795 3194 6890
rect 3224 6924 3284 7019
rect 3224 6890 3242 6924
rect 3276 6890 3284 6924
rect 3224 6795 3284 6890
rect 3502 6924 3562 7019
rect 3502 6890 3510 6924
rect 3544 6890 3562 6924
rect 3502 6795 3562 6890
rect 3592 6924 3652 7019
rect 3592 6890 3610 6924
rect 3644 6890 3652 6924
rect 3592 6795 3652 6890
rect 3760 6836 3820 7019
rect 3760 6802 3768 6836
rect 3802 6802 3820 6836
rect 3760 6619 3820 6802
rect 3850 6836 3910 7019
rect 3850 6802 3868 6836
rect 3902 6802 3910 6836
rect 3850 6619 3910 6802
rect 4018 6836 4078 7019
rect 4018 6802 4026 6836
rect 4060 6802 4078 6836
rect 4018 6619 4078 6802
rect 4108 6836 4168 7019
rect 4108 6802 4126 6836
rect 4160 6802 4168 6836
rect 4108 6619 4168 6802
rect 2666 4422 2726 4517
rect 2666 4388 2674 4422
rect 2708 4388 2726 4422
rect 2666 4293 2726 4388
rect 2756 4422 2816 4517
rect 2756 4388 2774 4422
rect 2808 4388 2816 4422
rect 2756 4293 2816 4388
rect 3034 4422 3094 4517
rect 3034 4388 3042 4422
rect 3076 4388 3094 4422
rect 3034 4293 3094 4388
rect 3124 4422 3184 4517
rect 3124 4388 3142 4422
rect 3176 4388 3184 4422
rect 3124 4293 3184 4388
rect 3292 4422 3352 4517
rect 3292 4388 3300 4422
rect 3334 4388 3352 4422
rect 3292 4293 3352 4388
rect 3382 4422 3442 4517
rect 3382 4388 3400 4422
rect 3434 4388 3442 4422
rect 3382 4293 3442 4388
rect 3550 4510 3610 4693
rect 3550 4476 3558 4510
rect 3592 4476 3610 4510
rect 3550 4293 3610 4476
rect 3640 4510 3700 4693
rect 3640 4476 3658 4510
rect 3692 4476 3700 4510
rect 3640 4293 3700 4476
rect 3808 4510 3868 4693
rect 3808 4476 3816 4510
rect 3850 4476 3868 4510
rect 3808 4293 3868 4476
rect 3898 4510 3958 4693
rect 3898 4476 3916 4510
rect 3950 4476 3958 4510
rect 3898 4293 3958 4476
rect 4066 4510 4126 4693
rect 4066 4476 4074 4510
rect 4108 4476 4126 4510
rect 4066 4293 4126 4476
rect 4156 4510 4216 4693
rect 4156 4476 4174 4510
rect 4208 4476 4216 4510
rect 4156 4293 4216 4476
rect 2666 4096 2726 4191
rect 2666 4062 2674 4096
rect 2708 4062 2726 4096
rect 2666 3967 2726 4062
rect 2756 4096 2826 4191
rect 2756 4062 2774 4096
rect 2808 4062 2826 4096
rect 2756 3967 2826 4062
rect 2856 4096 2916 4191
rect 2856 4062 2874 4096
rect 2908 4062 2916 4096
rect 2856 3967 2916 4062
rect 3044 4008 3104 4191
rect 3044 3974 3052 4008
rect 3086 3974 3104 4008
rect 3044 3791 3104 3974
rect 3134 4008 3194 4191
rect 3134 3974 3152 4008
rect 3186 3974 3194 4008
rect 3134 3791 3194 3974
rect 2666 1594 2726 1689
rect 2666 1560 2674 1594
rect 2708 1560 2726 1594
rect 2666 1465 2726 1560
rect 2756 1594 2816 1689
rect 2756 1560 2774 1594
rect 2808 1560 2816 1594
rect 2756 1465 2816 1560
rect 3034 1594 3094 1689
rect 3034 1560 3042 1594
rect 3076 1560 3094 1594
rect 3034 1465 3094 1560
rect 3124 1594 3194 1689
rect 3124 1560 3142 1594
rect 3176 1560 3194 1594
rect 3124 1465 3194 1560
rect 3224 1594 3284 1689
rect 3224 1560 3242 1594
rect 3276 1560 3284 1594
rect 3224 1465 3284 1560
rect 3412 1682 3472 1865
rect 3412 1648 3420 1682
rect 3454 1648 3472 1682
rect 3412 1465 3472 1648
rect 3502 1682 3562 1865
rect 3502 1648 3520 1682
rect 3554 1648 3562 1682
rect 3502 1465 3562 1648
rect 28 1279 81 1312
rect 28 1245 36 1279
rect 70 1245 81 1279
rect 28 1211 81 1245
rect 28 1177 36 1211
rect 70 1177 81 1211
rect 28 1143 81 1177
rect 28 1109 36 1143
rect 70 1109 81 1143
rect 28 1075 81 1109
rect 28 1041 36 1075
rect 70 1041 81 1075
rect 28 1007 81 1041
rect 28 973 36 1007
rect 70 973 81 1007
rect 28 939 81 973
rect 28 905 36 939
rect 70 905 81 939
rect 28 871 81 905
rect 28 837 36 871
rect 70 837 81 871
rect 28 712 81 837
rect 111 1279 167 1312
rect 111 1245 122 1279
rect 156 1245 167 1279
rect 111 1211 167 1245
rect 111 1177 122 1211
rect 156 1177 167 1211
rect 111 1143 167 1177
rect 111 1109 122 1143
rect 156 1109 167 1143
rect 111 1075 167 1109
rect 111 1041 122 1075
rect 156 1041 167 1075
rect 111 1007 167 1041
rect 111 973 122 1007
rect 156 973 167 1007
rect 111 939 167 973
rect 111 905 122 939
rect 156 905 167 939
rect 111 871 167 905
rect 111 837 122 871
rect 156 837 167 871
rect 111 712 167 837
rect 197 712 239 1312
rect 269 1279 359 1312
rect 269 1245 297 1279
rect 331 1245 359 1279
rect 269 1211 359 1245
rect 269 1177 297 1211
rect 331 1177 359 1211
rect 269 1143 359 1177
rect 269 1109 297 1143
rect 331 1109 359 1143
rect 269 1075 359 1109
rect 269 1041 297 1075
rect 331 1041 359 1075
rect 269 1007 359 1041
rect 269 973 297 1007
rect 331 973 359 1007
rect 269 939 359 973
rect 269 905 297 939
rect 331 905 359 939
rect 269 871 359 905
rect 269 837 297 871
rect 331 837 359 871
rect 269 712 359 837
rect 389 712 431 1312
rect 461 1279 517 1312
rect 461 1245 472 1279
rect 506 1245 517 1279
rect 461 1211 517 1245
rect 461 1177 472 1211
rect 506 1177 517 1211
rect 461 1143 517 1177
rect 461 1109 472 1143
rect 506 1109 517 1143
rect 461 1075 517 1109
rect 461 1041 472 1075
rect 506 1041 517 1075
rect 461 1007 517 1041
rect 461 973 472 1007
rect 506 973 517 1007
rect 461 939 517 973
rect 461 905 472 939
rect 506 905 517 939
rect 461 871 517 905
rect 461 837 472 871
rect 506 837 517 871
rect 461 712 517 837
rect 547 712 589 1312
rect 619 1279 709 1312
rect 619 1245 647 1279
rect 681 1245 709 1279
rect 619 1211 709 1245
rect 619 1177 647 1211
rect 681 1177 709 1211
rect 619 1143 709 1177
rect 619 1109 647 1143
rect 681 1109 709 1143
rect 619 1075 709 1109
rect 619 1041 647 1075
rect 681 1041 709 1075
rect 619 1007 709 1041
rect 619 973 647 1007
rect 681 973 709 1007
rect 619 939 709 973
rect 619 905 647 939
rect 681 905 709 939
rect 619 871 709 905
rect 619 837 647 871
rect 681 837 709 871
rect 619 712 709 837
rect 739 712 781 1312
rect 811 1279 867 1312
rect 811 1245 822 1279
rect 856 1245 867 1279
rect 811 1211 867 1245
rect 811 1177 822 1211
rect 856 1177 867 1211
rect 811 1143 867 1177
rect 811 1109 822 1143
rect 856 1109 867 1143
rect 811 1075 867 1109
rect 811 1041 822 1075
rect 856 1041 867 1075
rect 811 1007 867 1041
rect 811 973 822 1007
rect 856 973 867 1007
rect 811 939 867 973
rect 811 905 822 939
rect 856 905 867 939
rect 811 871 867 905
rect 811 837 822 871
rect 856 837 867 871
rect 811 712 867 837
rect 897 1279 950 1312
rect 897 1245 908 1279
rect 942 1245 950 1279
rect 897 1211 950 1245
rect 897 1177 908 1211
rect 942 1177 950 1211
rect 897 1143 950 1177
rect 897 1109 908 1143
rect 942 1109 950 1143
rect 897 1075 950 1109
rect 897 1041 908 1075
rect 942 1041 950 1075
rect 897 1007 950 1041
rect 897 973 908 1007
rect 942 973 950 1007
rect 897 939 950 973
rect 897 905 908 939
rect 942 905 950 939
rect 897 871 950 905
rect 897 837 908 871
rect 942 837 950 871
rect 897 712 950 837
rect 1004 1279 1057 1312
rect 1004 1245 1012 1279
rect 1046 1245 1057 1279
rect 1004 1211 1057 1245
rect 1004 1177 1012 1211
rect 1046 1177 1057 1211
rect 1004 1143 1057 1177
rect 1004 1109 1012 1143
rect 1046 1109 1057 1143
rect 1004 1075 1057 1109
rect 1004 1041 1012 1075
rect 1046 1041 1057 1075
rect 1004 1007 1057 1041
rect 1004 973 1012 1007
rect 1046 973 1057 1007
rect 1004 939 1057 973
rect 1004 905 1012 939
rect 1046 905 1057 939
rect 1004 871 1057 905
rect 1004 837 1012 871
rect 1046 837 1057 871
rect 1004 712 1057 837
rect 1087 1279 1140 1312
rect 1087 1245 1098 1279
rect 1132 1245 1140 1279
rect 1087 1211 1140 1245
rect 1087 1177 1098 1211
rect 1132 1177 1140 1211
rect 1087 1143 1140 1177
rect 1087 1109 1098 1143
rect 1132 1109 1140 1143
rect 1258 1268 1318 1363
rect 1258 1234 1266 1268
rect 1300 1234 1318 1268
rect 1258 1139 1318 1234
rect 1348 1268 1408 1363
rect 1348 1234 1366 1268
rect 1400 1234 1408 1268
rect 1348 1139 1408 1234
rect 1626 1215 1686 1363
rect 1626 1181 1634 1215
rect 1668 1181 1686 1215
rect 1087 1075 1140 1109
rect 1087 1041 1098 1075
rect 1132 1041 1140 1075
rect 1087 1007 1140 1041
rect 1087 973 1098 1007
rect 1132 973 1140 1007
rect 1087 939 1140 973
rect 1087 905 1098 939
rect 1132 905 1140 939
rect 1087 871 1140 905
rect 1087 837 1098 871
rect 1132 837 1140 871
rect 1087 712 1140 837
rect 1626 1033 1686 1181
rect 1716 1215 1776 1363
rect 1716 1181 1734 1215
rect 1768 1181 1776 1215
rect 1716 1033 1776 1181
rect 2666 1268 2726 1363
rect 2666 1234 2674 1268
rect 2708 1234 2726 1268
rect 2666 1139 2726 1234
rect 2756 1268 2816 1363
rect 2756 1234 2774 1268
rect 2808 1234 2816 1268
rect 2756 1139 2816 1234
rect 3034 1268 3094 1363
rect 3034 1234 3042 1268
rect 3076 1234 3094 1268
rect 3034 1139 3094 1234
rect 3124 1268 3184 1363
rect 3124 1234 3142 1268
rect 3176 1234 3184 1268
rect 3124 1139 3184 1234
rect 3292 1215 3352 1363
rect 3292 1181 3300 1215
rect 3334 1181 3352 1215
rect 3292 1033 3352 1181
rect 3382 1215 3442 1363
rect 3382 1181 3400 1215
rect 3434 1181 3442 1215
rect 3382 1033 3442 1181
rect 3550 1180 3610 1363
rect 3550 1146 3558 1180
rect 3592 1146 3610 1180
rect 3550 963 3610 1146
rect 3640 1180 3700 1363
rect 3640 1146 3658 1180
rect 3692 1146 3700 1180
rect 3640 963 3700 1146
rect 3808 1180 3868 1363
rect 3808 1146 3816 1180
rect 3850 1146 3868 1180
rect 3808 963 3868 1146
rect 3898 1180 3958 1363
rect 3898 1146 3916 1180
rect 3950 1146 3958 1180
rect 3898 963 3958 1146
rect 4066 1180 4126 1363
rect 4066 1146 4074 1180
rect 4108 1146 4126 1180
rect 4066 963 4126 1146
rect 4156 1180 4216 1363
rect 4156 1146 4174 1180
rect 4208 1146 4216 1180
rect 4156 963 4216 1146
<< ndiffc >>
rect 172 17674 206 17708
rect 272 17674 306 17708
rect 540 17674 574 17708
rect 640 17674 674 17708
rect 908 17674 942 17708
rect 1008 17674 1042 17708
rect 1276 17674 1310 17708
rect 1376 17674 1410 17708
rect 1644 17674 1678 17708
rect 1744 17674 1778 17708
rect 172 17500 206 17534
rect 272 17500 306 17534
rect 540 17500 574 17534
rect 640 17500 674 17534
rect 908 17500 942 17534
rect 1008 17500 1042 17534
rect 1276 17500 1310 17534
rect 1376 17500 1410 17534
rect 1644 17500 1678 17534
rect 1744 17500 1778 17534
rect 172 15434 206 15468
rect 272 15434 306 15468
rect 540 15434 574 15468
rect 640 15434 674 15468
rect 908 15434 942 15468
rect 1008 15434 1042 15468
rect 1276 15434 1310 15468
rect 1376 15434 1410 15468
rect 1644 15434 1678 15468
rect 1744 15434 1778 15468
rect 172 15260 206 15294
rect 272 15260 306 15294
rect 540 15260 574 15294
rect 640 15260 674 15294
rect 908 15260 942 15294
rect 1008 15260 1042 15294
rect 1276 15260 1310 15294
rect 1376 15260 1410 15294
rect 1644 15260 1678 15294
rect 1744 15260 1778 15294
rect 172 13194 206 13228
rect 272 13194 306 13228
rect 540 13194 574 13228
rect 640 13194 674 13228
rect 908 13194 942 13228
rect 1008 13194 1042 13228
rect 1276 13194 1310 13228
rect 1376 13194 1410 13228
rect 1644 13194 1678 13228
rect 1744 13194 1778 13228
rect 172 13020 206 13054
rect 272 13020 306 13054
rect 540 13020 574 13054
rect 640 13020 674 13054
rect 908 13020 942 13054
rect 1008 13020 1042 13054
rect 1276 13020 1310 13054
rect 1376 13020 1410 13054
rect 1644 13020 1678 13054
rect 1744 13020 1778 13054
rect 172 10954 206 10988
rect 272 10954 306 10988
rect 540 10954 574 10988
rect 640 10954 674 10988
rect 908 10954 942 10988
rect 1008 10954 1042 10988
rect 1276 10954 1310 10988
rect 1376 10954 1410 10988
rect 1644 10954 1678 10988
rect 1744 10954 1778 10988
rect 172 10780 206 10814
rect 272 10780 306 10814
rect 540 10780 574 10814
rect 640 10780 674 10814
rect 908 10780 942 10814
rect 1008 10780 1042 10814
rect 1276 10780 1310 10814
rect 1376 10780 1410 10814
rect 1644 10780 1678 10814
rect 1744 10780 1778 10814
rect 172 8714 206 8748
rect 272 8714 306 8748
rect 540 8714 574 8748
rect 640 8714 674 8748
rect 908 8714 942 8748
rect 1008 8714 1042 8748
rect 1276 8714 1310 8748
rect 1376 8714 1410 8748
rect 1644 8714 1678 8748
rect 1744 8714 1778 8748
rect 2674 8342 2708 8376
rect 2974 8342 3008 8376
rect 3152 8216 3186 8250
rect 3252 8216 3286 8250
rect 2674 5764 2708 5798
rect 2874 5764 2908 5798
rect 3142 5726 3176 5760
rect 3242 5726 3276 5760
rect 3510 5764 3544 5798
rect 3610 5764 3644 5798
rect 3768 5816 3802 5850
rect 3868 5816 3902 5850
rect 4026 5890 4060 5924
rect 4126 5890 4160 5924
rect 2674 5552 2708 5586
rect 2774 5552 2808 5586
rect 3042 5476 3076 5510
rect 3142 5476 3176 5510
rect 3300 5514 3334 5548
rect 3400 5514 3434 5548
rect 3558 5388 3592 5422
rect 3658 5388 3692 5422
rect 3816 5420 3850 5454
rect 3916 5420 3950 5454
rect 4074 5388 4108 5422
rect 4174 5388 4208 5422
rect 3052 3030 3086 3064
rect 2674 2936 2708 2970
rect 2874 2936 2908 2970
rect 3152 3030 3186 3064
rect 2674 2724 2708 2758
rect 2774 2724 2808 2758
rect 3042 2686 3076 2720
rect 3242 2686 3276 2720
rect 3420 2592 3454 2626
rect 3520 2592 3554 2626
rect 36 203 70 237
rect 36 135 70 169
rect 122 203 156 237
rect 122 135 156 169
rect 297 203 331 237
rect 297 135 331 169
rect 472 203 506 237
rect 472 135 506 169
rect 647 203 681 237
rect 647 135 681 169
rect 822 203 856 237
rect 822 135 856 169
rect 908 203 942 237
rect 908 135 942 169
rect 1012 203 1046 237
rect 1012 135 1046 169
rect 1098 203 1132 237
rect 1634 202 1668 236
rect 1098 135 1132 169
rect 1266 108 1300 142
rect 1366 108 1400 142
rect 1734 202 1768 236
rect 2674 70 2708 104
rect 2774 70 2808 104
rect 3300 160 3334 194
rect 3042 70 3076 104
rect 3142 70 3176 104
rect 3400 160 3434 194
rect 3558 202 3592 236
rect 3658 202 3692 236
rect 3816 234 3850 268
rect 3916 234 3950 268
rect 4074 234 4108 268
rect 4174 234 4208 268
<< pdiffc >>
rect 172 18544 206 18578
rect 272 18544 306 18578
rect 540 18544 574 18578
rect 640 18544 674 18578
rect 908 18544 942 18578
rect 1008 18544 1042 18578
rect 1276 18544 1310 18578
rect 1376 18544 1410 18578
rect 1644 18544 1678 18578
rect 1744 18544 1778 18578
rect 172 16630 206 16664
rect 272 16630 306 16664
rect 540 16630 574 16664
rect 640 16630 674 16664
rect 908 16630 942 16664
rect 1008 16630 1042 16664
rect 1276 16630 1310 16664
rect 1376 16630 1410 16664
rect 1644 16630 1678 16664
rect 1744 16630 1778 16664
rect 172 16304 206 16338
rect 272 16304 306 16338
rect 540 16304 574 16338
rect 640 16304 674 16338
rect 908 16304 942 16338
rect 1008 16304 1042 16338
rect 1276 16304 1310 16338
rect 1376 16304 1410 16338
rect 1644 16304 1678 16338
rect 1744 16304 1778 16338
rect 172 14390 206 14424
rect 272 14390 306 14424
rect 540 14390 574 14424
rect 640 14390 674 14424
rect 908 14390 942 14424
rect 1008 14390 1042 14424
rect 1276 14390 1310 14424
rect 1376 14390 1410 14424
rect 1644 14390 1678 14424
rect 1744 14390 1778 14424
rect 172 14064 206 14098
rect 272 14064 306 14098
rect 540 14064 574 14098
rect 640 14064 674 14098
rect 908 14064 942 14098
rect 1008 14064 1042 14098
rect 1276 14064 1310 14098
rect 1376 14064 1410 14098
rect 1644 14064 1678 14098
rect 1744 14064 1778 14098
rect 172 12150 206 12184
rect 272 12150 306 12184
rect 540 12150 574 12184
rect 640 12150 674 12184
rect 908 12150 942 12184
rect 1008 12150 1042 12184
rect 1276 12150 1310 12184
rect 1376 12150 1410 12184
rect 1644 12150 1678 12184
rect 1744 12150 1778 12184
rect 172 11824 206 11858
rect 272 11824 306 11858
rect 540 11824 574 11858
rect 640 11824 674 11858
rect 908 11824 942 11858
rect 1008 11824 1042 11858
rect 1276 11824 1310 11858
rect 1376 11824 1410 11858
rect 1644 11824 1678 11858
rect 1744 11824 1778 11858
rect 172 9910 206 9944
rect 272 9910 306 9944
rect 540 9910 574 9944
rect 640 9910 674 9944
rect 908 9910 942 9944
rect 1008 9910 1042 9944
rect 1276 9910 1310 9944
rect 1376 9910 1410 9944
rect 1644 9910 1678 9944
rect 1744 9910 1778 9944
rect 172 9584 206 9618
rect 272 9584 306 9618
rect 540 9584 574 9618
rect 640 9584 674 9618
rect 908 9584 942 9618
rect 1008 9584 1042 9618
rect 1276 9584 1310 9618
rect 1376 9584 1410 9618
rect 1644 9584 1678 9618
rect 1744 9584 1778 9618
rect 2674 7216 2708 7250
rect 2774 7216 2808 7250
rect 2874 7216 2908 7250
rect 2974 7216 3008 7250
rect 3152 7304 3186 7338
rect 3252 7304 3286 7338
rect 2674 6890 2708 6924
rect 2774 6890 2808 6924
rect 2874 6890 2908 6924
rect 3142 6890 3176 6924
rect 3242 6890 3276 6924
rect 3510 6890 3544 6924
rect 3610 6890 3644 6924
rect 3768 6802 3802 6836
rect 3868 6802 3902 6836
rect 4026 6802 4060 6836
rect 4126 6802 4160 6836
rect 2674 4388 2708 4422
rect 2774 4388 2808 4422
rect 3042 4388 3076 4422
rect 3142 4388 3176 4422
rect 3300 4388 3334 4422
rect 3400 4388 3434 4422
rect 3558 4476 3592 4510
rect 3658 4476 3692 4510
rect 3816 4476 3850 4510
rect 3916 4476 3950 4510
rect 4074 4476 4108 4510
rect 4174 4476 4208 4510
rect 2674 4062 2708 4096
rect 2774 4062 2808 4096
rect 2874 4062 2908 4096
rect 3052 3974 3086 4008
rect 3152 3974 3186 4008
rect 2674 1560 2708 1594
rect 2774 1560 2808 1594
rect 3042 1560 3076 1594
rect 3142 1560 3176 1594
rect 3242 1560 3276 1594
rect 3420 1648 3454 1682
rect 3520 1648 3554 1682
rect 36 1245 70 1279
rect 36 1177 70 1211
rect 36 1109 70 1143
rect 36 1041 70 1075
rect 36 973 70 1007
rect 36 905 70 939
rect 36 837 70 871
rect 122 1245 156 1279
rect 122 1177 156 1211
rect 122 1109 156 1143
rect 122 1041 156 1075
rect 122 973 156 1007
rect 122 905 156 939
rect 122 837 156 871
rect 297 1245 331 1279
rect 297 1177 331 1211
rect 297 1109 331 1143
rect 297 1041 331 1075
rect 297 973 331 1007
rect 297 905 331 939
rect 297 837 331 871
rect 472 1245 506 1279
rect 472 1177 506 1211
rect 472 1109 506 1143
rect 472 1041 506 1075
rect 472 973 506 1007
rect 472 905 506 939
rect 472 837 506 871
rect 647 1245 681 1279
rect 647 1177 681 1211
rect 647 1109 681 1143
rect 647 1041 681 1075
rect 647 973 681 1007
rect 647 905 681 939
rect 647 837 681 871
rect 822 1245 856 1279
rect 822 1177 856 1211
rect 822 1109 856 1143
rect 822 1041 856 1075
rect 822 973 856 1007
rect 822 905 856 939
rect 822 837 856 871
rect 908 1245 942 1279
rect 908 1177 942 1211
rect 908 1109 942 1143
rect 908 1041 942 1075
rect 908 973 942 1007
rect 908 905 942 939
rect 908 837 942 871
rect 1012 1245 1046 1279
rect 1012 1177 1046 1211
rect 1012 1109 1046 1143
rect 1012 1041 1046 1075
rect 1012 973 1046 1007
rect 1012 905 1046 939
rect 1012 837 1046 871
rect 1098 1245 1132 1279
rect 1098 1177 1132 1211
rect 1098 1109 1132 1143
rect 1266 1234 1300 1268
rect 1366 1234 1400 1268
rect 1634 1181 1668 1215
rect 1098 1041 1132 1075
rect 1098 973 1132 1007
rect 1098 905 1132 939
rect 1098 837 1132 871
rect 1734 1181 1768 1215
rect 2674 1234 2708 1268
rect 2774 1234 2808 1268
rect 3042 1234 3076 1268
rect 3142 1234 3176 1268
rect 3300 1181 3334 1215
rect 3400 1181 3434 1215
rect 3558 1146 3592 1180
rect 3658 1146 3692 1180
rect 3816 1146 3850 1180
rect 3916 1146 3950 1180
rect 4074 1146 4108 1180
rect 4174 1146 4208 1180
<< psubdiff >>
rect 60 17713 110 17737
rect 60 17679 68 17713
rect 102 17679 110 17713
rect 60 17655 110 17679
rect 428 17713 478 17737
rect 428 17679 436 17713
rect 470 17679 478 17713
rect 428 17655 478 17679
rect 796 17713 846 17737
rect 796 17679 804 17713
rect 838 17679 846 17713
rect 796 17655 846 17679
rect 1164 17713 1214 17737
rect 1164 17679 1172 17713
rect 1206 17679 1214 17713
rect 1164 17655 1214 17679
rect 1532 17713 1582 17737
rect 1532 17679 1540 17713
rect 1574 17679 1582 17713
rect 1532 17655 1582 17679
rect 60 17529 110 17553
rect 60 17495 68 17529
rect 102 17495 110 17529
rect 60 17471 110 17495
rect 428 17529 478 17553
rect 428 17495 436 17529
rect 470 17495 478 17529
rect 428 17471 478 17495
rect 796 17529 846 17553
rect 796 17495 804 17529
rect 838 17495 846 17529
rect 796 17471 846 17495
rect 1164 17529 1214 17553
rect 1164 17495 1172 17529
rect 1206 17495 1214 17529
rect 1164 17471 1214 17495
rect 1532 17529 1582 17553
rect 1532 17495 1540 17529
rect 1574 17495 1582 17529
rect 1532 17471 1582 17495
rect 60 15473 110 15497
rect 60 15439 68 15473
rect 102 15439 110 15473
rect 60 15415 110 15439
rect 428 15473 478 15497
rect 428 15439 436 15473
rect 470 15439 478 15473
rect 428 15415 478 15439
rect 796 15473 846 15497
rect 796 15439 804 15473
rect 838 15439 846 15473
rect 796 15415 846 15439
rect 1164 15473 1214 15497
rect 1164 15439 1172 15473
rect 1206 15439 1214 15473
rect 1164 15415 1214 15439
rect 1532 15473 1582 15497
rect 1532 15439 1540 15473
rect 1574 15439 1582 15473
rect 1532 15415 1582 15439
rect 60 15289 110 15313
rect 60 15255 68 15289
rect 102 15255 110 15289
rect 60 15231 110 15255
rect 428 15289 478 15313
rect 428 15255 436 15289
rect 470 15255 478 15289
rect 428 15231 478 15255
rect 796 15289 846 15313
rect 796 15255 804 15289
rect 838 15255 846 15289
rect 796 15231 846 15255
rect 1164 15289 1214 15313
rect 1164 15255 1172 15289
rect 1206 15255 1214 15289
rect 1164 15231 1214 15255
rect 1532 15289 1582 15313
rect 1532 15255 1540 15289
rect 1574 15255 1582 15289
rect 1532 15231 1582 15255
rect 60 13233 110 13257
rect 60 13199 68 13233
rect 102 13199 110 13233
rect 60 13175 110 13199
rect 428 13233 478 13257
rect 428 13199 436 13233
rect 470 13199 478 13233
rect 428 13175 478 13199
rect 796 13233 846 13257
rect 796 13199 804 13233
rect 838 13199 846 13233
rect 796 13175 846 13199
rect 1164 13233 1214 13257
rect 1164 13199 1172 13233
rect 1206 13199 1214 13233
rect 1164 13175 1214 13199
rect 1532 13233 1582 13257
rect 1532 13199 1540 13233
rect 1574 13199 1582 13233
rect 1532 13175 1582 13199
rect 60 13049 110 13073
rect 60 13015 68 13049
rect 102 13015 110 13049
rect 60 12991 110 13015
rect 428 13049 478 13073
rect 428 13015 436 13049
rect 470 13015 478 13049
rect 428 12991 478 13015
rect 796 13049 846 13073
rect 796 13015 804 13049
rect 838 13015 846 13049
rect 796 12991 846 13015
rect 1164 13049 1214 13073
rect 1164 13015 1172 13049
rect 1206 13015 1214 13049
rect 1164 12991 1214 13015
rect 1532 13049 1582 13073
rect 1532 13015 1540 13049
rect 1574 13015 1582 13049
rect 1532 12991 1582 13015
rect 60 10993 110 11017
rect 60 10959 68 10993
rect 102 10959 110 10993
rect 60 10935 110 10959
rect 428 10993 478 11017
rect 428 10959 436 10993
rect 470 10959 478 10993
rect 428 10935 478 10959
rect 796 10993 846 11017
rect 796 10959 804 10993
rect 838 10959 846 10993
rect 796 10935 846 10959
rect 1164 10993 1214 11017
rect 1164 10959 1172 10993
rect 1206 10959 1214 10993
rect 1164 10935 1214 10959
rect 1532 10993 1582 11017
rect 1532 10959 1540 10993
rect 1574 10959 1582 10993
rect 1532 10935 1582 10959
rect 60 10809 110 10833
rect 60 10775 68 10809
rect 102 10775 110 10809
rect 60 10751 110 10775
rect 428 10809 478 10833
rect 428 10775 436 10809
rect 470 10775 478 10809
rect 428 10751 478 10775
rect 796 10809 846 10833
rect 796 10775 804 10809
rect 838 10775 846 10809
rect 796 10751 846 10775
rect 1164 10809 1214 10833
rect 1164 10775 1172 10809
rect 1206 10775 1214 10809
rect 1164 10751 1214 10775
rect 1532 10809 1582 10833
rect 1532 10775 1540 10809
rect 1574 10775 1582 10809
rect 1532 10751 1582 10775
rect 60 8753 110 8777
rect 60 8719 68 8753
rect 102 8719 110 8753
rect 60 8695 110 8719
rect 428 8753 478 8777
rect 428 8719 436 8753
rect 470 8719 478 8753
rect 428 8695 478 8719
rect 796 8753 846 8777
rect 796 8719 804 8753
rect 838 8719 846 8753
rect 796 8695 846 8719
rect 1164 8753 1214 8777
rect 1164 8719 1172 8753
rect 1206 8719 1214 8753
rect 1164 8695 1214 8719
rect 1532 8753 1582 8777
rect 1532 8719 1540 8753
rect 1574 8719 1582 8753
rect 1532 8695 1582 8719
rect 3348 8409 3398 8433
rect 3348 8375 3356 8409
rect 3390 8375 3398 8409
rect 3348 8351 3398 8375
rect 2970 5782 3020 5806
rect 2970 5748 2978 5782
rect 3012 5748 3020 5782
rect 2970 5724 3020 5748
rect 3338 5765 3388 5789
rect 3338 5731 3346 5765
rect 3380 5731 3388 5765
rect 3338 5707 3388 5731
rect 2870 5564 2920 5588
rect 2870 5530 2878 5564
rect 2912 5530 2920 5564
rect 2870 5506 2920 5530
rect 3248 2937 3298 2961
rect 3248 2903 3256 2937
rect 3290 2903 3298 2937
rect 3248 2879 3298 2903
rect 2870 2753 2920 2777
rect 2870 2719 2878 2753
rect 2912 2719 2920 2753
rect 2870 2695 2920 2719
rect 3616 2753 3666 2777
rect 3616 2719 3624 2753
rect 3658 2719 3666 2753
rect 3616 2695 3666 2719
rect 1462 109 1512 133
rect 1462 75 1470 109
rect 1504 75 1512 109
rect 1462 51 1512 75
rect 1830 109 1880 133
rect 1830 75 1838 109
rect 1872 75 1880 109
rect 1830 51 1880 75
rect 2870 109 2920 133
rect 2870 75 2878 109
rect 2912 75 2920 109
rect 2870 51 2920 75
rect 28 -17 52 17
rect 86 -17 110 17
rect 164 -17 188 17
rect 222 -17 246 17
rect 300 -17 324 17
rect 358 -17 382 17
rect 436 -17 460 17
rect 494 -17 518 17
rect 572 -17 596 17
rect 630 -17 654 17
rect 708 -17 732 17
rect 766 -17 790 17
rect 844 -17 868 17
rect 902 -17 926 17
rect 980 -17 1004 17
rect 1038 -17 1062 17
<< nsubdiff >>
rect 60 18649 110 18673
rect 60 18615 68 18649
rect 102 18615 110 18649
rect 60 18591 110 18615
rect 428 18649 478 18673
rect 428 18615 436 18649
rect 470 18615 478 18649
rect 428 18591 478 18615
rect 796 18649 846 18673
rect 796 18615 804 18649
rect 838 18615 846 18649
rect 796 18591 846 18615
rect 1164 18649 1214 18673
rect 1164 18615 1172 18649
rect 1206 18615 1214 18649
rect 1164 18591 1214 18615
rect 1532 18649 1582 18673
rect 1532 18615 1540 18649
rect 1574 18615 1582 18649
rect 1532 18591 1582 18615
rect 60 16593 110 16617
rect 60 16559 68 16593
rect 102 16559 110 16593
rect 60 16535 110 16559
rect 428 16593 478 16617
rect 428 16559 436 16593
rect 470 16559 478 16593
rect 428 16535 478 16559
rect 796 16593 846 16617
rect 796 16559 804 16593
rect 838 16559 846 16593
rect 796 16535 846 16559
rect 1164 16593 1214 16617
rect 1164 16559 1172 16593
rect 1206 16559 1214 16593
rect 1164 16535 1214 16559
rect 1532 16593 1582 16617
rect 1532 16559 1540 16593
rect 1574 16559 1582 16593
rect 1532 16535 1582 16559
rect 60 16409 110 16433
rect 60 16375 68 16409
rect 102 16375 110 16409
rect 60 16351 110 16375
rect 428 16409 478 16433
rect 428 16375 436 16409
rect 470 16375 478 16409
rect 428 16351 478 16375
rect 796 16409 846 16433
rect 796 16375 804 16409
rect 838 16375 846 16409
rect 796 16351 846 16375
rect 1164 16409 1214 16433
rect 1164 16375 1172 16409
rect 1206 16375 1214 16409
rect 1164 16351 1214 16375
rect 1532 16409 1582 16433
rect 1532 16375 1540 16409
rect 1574 16375 1582 16409
rect 1532 16351 1582 16375
rect 60 14353 110 14377
rect 60 14319 68 14353
rect 102 14319 110 14353
rect 60 14295 110 14319
rect 428 14353 478 14377
rect 428 14319 436 14353
rect 470 14319 478 14353
rect 428 14295 478 14319
rect 796 14353 846 14377
rect 796 14319 804 14353
rect 838 14319 846 14353
rect 796 14295 846 14319
rect 1164 14353 1214 14377
rect 1164 14319 1172 14353
rect 1206 14319 1214 14353
rect 1164 14295 1214 14319
rect 1532 14353 1582 14377
rect 1532 14319 1540 14353
rect 1574 14319 1582 14353
rect 1532 14295 1582 14319
rect 60 14169 110 14193
rect 60 14135 68 14169
rect 102 14135 110 14169
rect 60 14111 110 14135
rect 428 14169 478 14193
rect 428 14135 436 14169
rect 470 14135 478 14169
rect 428 14111 478 14135
rect 796 14169 846 14193
rect 796 14135 804 14169
rect 838 14135 846 14169
rect 796 14111 846 14135
rect 1164 14169 1214 14193
rect 1164 14135 1172 14169
rect 1206 14135 1214 14169
rect 1164 14111 1214 14135
rect 1532 14169 1582 14193
rect 1532 14135 1540 14169
rect 1574 14135 1582 14169
rect 1532 14111 1582 14135
rect 60 12113 110 12137
rect 60 12079 68 12113
rect 102 12079 110 12113
rect 60 12055 110 12079
rect 428 12113 478 12137
rect 428 12079 436 12113
rect 470 12079 478 12113
rect 428 12055 478 12079
rect 796 12113 846 12137
rect 796 12079 804 12113
rect 838 12079 846 12113
rect 796 12055 846 12079
rect 1164 12113 1214 12137
rect 1164 12079 1172 12113
rect 1206 12079 1214 12113
rect 1164 12055 1214 12079
rect 1532 12113 1582 12137
rect 1532 12079 1540 12113
rect 1574 12079 1582 12113
rect 1532 12055 1582 12079
rect 60 11929 110 11953
rect 60 11895 68 11929
rect 102 11895 110 11929
rect 60 11871 110 11895
rect 428 11929 478 11953
rect 428 11895 436 11929
rect 470 11895 478 11929
rect 428 11871 478 11895
rect 796 11929 846 11953
rect 796 11895 804 11929
rect 838 11895 846 11929
rect 796 11871 846 11895
rect 1164 11929 1214 11953
rect 1164 11895 1172 11929
rect 1206 11895 1214 11929
rect 1164 11871 1214 11895
rect 1532 11929 1582 11953
rect 1532 11895 1540 11929
rect 1574 11895 1582 11929
rect 1532 11871 1582 11895
rect 60 9873 110 9897
rect 60 9839 68 9873
rect 102 9839 110 9873
rect 60 9815 110 9839
rect 428 9873 478 9897
rect 428 9839 436 9873
rect 470 9839 478 9873
rect 428 9815 478 9839
rect 796 9873 846 9897
rect 796 9839 804 9873
rect 838 9839 846 9873
rect 796 9815 846 9839
rect 1164 9873 1214 9897
rect 1164 9839 1172 9873
rect 1206 9839 1214 9873
rect 1164 9815 1214 9839
rect 1532 9873 1582 9897
rect 1532 9839 1540 9873
rect 1574 9839 1582 9873
rect 1532 9815 1582 9839
rect 60 9689 110 9713
rect 60 9655 68 9689
rect 102 9655 110 9689
rect 60 9631 110 9655
rect 428 9689 478 9713
rect 428 9655 436 9689
rect 470 9655 478 9689
rect 428 9631 478 9655
rect 796 9689 846 9713
rect 796 9655 804 9689
rect 838 9655 846 9689
rect 796 9631 846 9655
rect 1164 9689 1214 9713
rect 1164 9655 1172 9689
rect 1206 9655 1214 9689
rect 1164 9631 1214 9655
rect 1532 9689 1582 9713
rect 1532 9655 1540 9689
rect 1574 9655 1582 9689
rect 1532 9631 1582 9655
rect 3348 7179 3398 7203
rect 3348 7145 3356 7179
rect 3390 7145 3398 7179
rect 3348 7121 3398 7145
rect 2970 6995 3020 7019
rect 2970 6961 2978 6995
rect 3012 6961 3020 6995
rect 2970 6937 3020 6961
rect 3338 6995 3388 7019
rect 3338 6961 3346 6995
rect 3380 6961 3388 6995
rect 3338 6937 3388 6961
rect 2870 4351 2920 4375
rect 2870 4317 2878 4351
rect 2912 4317 2920 4351
rect 2870 4293 2920 4317
rect 3248 4167 3298 4191
rect 3248 4133 3256 4167
rect 3290 4133 3298 4167
rect 3248 4109 3298 4133
rect 2870 1523 2920 1547
rect 2870 1489 2878 1523
rect 2912 1489 2920 1523
rect 2870 1465 2920 1489
rect 3616 1523 3666 1547
rect 3616 1489 3624 1523
rect 3658 1489 3666 1523
rect 3616 1465 3666 1489
rect 28 1397 52 1431
rect 86 1397 110 1431
rect 164 1397 188 1431
rect 222 1397 246 1431
rect 300 1397 324 1431
rect 358 1397 382 1431
rect 436 1397 460 1431
rect 494 1397 518 1431
rect 572 1397 596 1431
rect 630 1397 654 1431
rect 708 1397 732 1431
rect 766 1397 790 1431
rect 844 1397 868 1431
rect 902 1397 926 1431
rect 980 1397 1004 1431
rect 1038 1397 1062 1431
rect 1462 1339 1512 1363
rect 1462 1305 1470 1339
rect 1504 1305 1512 1339
rect 1462 1281 1512 1305
rect 1830 1339 1880 1363
rect 1830 1305 1838 1339
rect 1872 1305 1880 1339
rect 1830 1281 1880 1305
rect 2870 1339 2920 1363
rect 2870 1305 2878 1339
rect 2912 1305 2920 1339
rect 2870 1281 2920 1305
<< psubdiffcont >>
rect 68 17679 102 17713
rect 436 17679 470 17713
rect 804 17679 838 17713
rect 1172 17679 1206 17713
rect 1540 17679 1574 17713
rect 68 17495 102 17529
rect 436 17495 470 17529
rect 804 17495 838 17529
rect 1172 17495 1206 17529
rect 1540 17495 1574 17529
rect 68 15439 102 15473
rect 436 15439 470 15473
rect 804 15439 838 15473
rect 1172 15439 1206 15473
rect 1540 15439 1574 15473
rect 68 15255 102 15289
rect 436 15255 470 15289
rect 804 15255 838 15289
rect 1172 15255 1206 15289
rect 1540 15255 1574 15289
rect 68 13199 102 13233
rect 436 13199 470 13233
rect 804 13199 838 13233
rect 1172 13199 1206 13233
rect 1540 13199 1574 13233
rect 68 13015 102 13049
rect 436 13015 470 13049
rect 804 13015 838 13049
rect 1172 13015 1206 13049
rect 1540 13015 1574 13049
rect 68 10959 102 10993
rect 436 10959 470 10993
rect 804 10959 838 10993
rect 1172 10959 1206 10993
rect 1540 10959 1574 10993
rect 68 10775 102 10809
rect 436 10775 470 10809
rect 804 10775 838 10809
rect 1172 10775 1206 10809
rect 1540 10775 1574 10809
rect 68 8719 102 8753
rect 436 8719 470 8753
rect 804 8719 838 8753
rect 1172 8719 1206 8753
rect 1540 8719 1574 8753
rect 3356 8375 3390 8409
rect 2978 5748 3012 5782
rect 3346 5731 3380 5765
rect 2878 5530 2912 5564
rect 3256 2903 3290 2937
rect 2878 2719 2912 2753
rect 3624 2719 3658 2753
rect 1470 75 1504 109
rect 1838 75 1872 109
rect 2878 75 2912 109
rect 52 -17 86 17
rect 188 -17 222 17
rect 324 -17 358 17
rect 460 -17 494 17
rect 596 -17 630 17
rect 732 -17 766 17
rect 868 -17 902 17
rect 1004 -17 1038 17
<< nsubdiffcont >>
rect 68 18615 102 18649
rect 436 18615 470 18649
rect 804 18615 838 18649
rect 1172 18615 1206 18649
rect 1540 18615 1574 18649
rect 68 16559 102 16593
rect 436 16559 470 16593
rect 804 16559 838 16593
rect 1172 16559 1206 16593
rect 1540 16559 1574 16593
rect 68 16375 102 16409
rect 436 16375 470 16409
rect 804 16375 838 16409
rect 1172 16375 1206 16409
rect 1540 16375 1574 16409
rect 68 14319 102 14353
rect 436 14319 470 14353
rect 804 14319 838 14353
rect 1172 14319 1206 14353
rect 1540 14319 1574 14353
rect 68 14135 102 14169
rect 436 14135 470 14169
rect 804 14135 838 14169
rect 1172 14135 1206 14169
rect 1540 14135 1574 14169
rect 68 12079 102 12113
rect 436 12079 470 12113
rect 804 12079 838 12113
rect 1172 12079 1206 12113
rect 1540 12079 1574 12113
rect 68 11895 102 11929
rect 436 11895 470 11929
rect 804 11895 838 11929
rect 1172 11895 1206 11929
rect 1540 11895 1574 11929
rect 68 9839 102 9873
rect 436 9839 470 9873
rect 804 9839 838 9873
rect 1172 9839 1206 9873
rect 1540 9839 1574 9873
rect 68 9655 102 9689
rect 436 9655 470 9689
rect 804 9655 838 9689
rect 1172 9655 1206 9689
rect 1540 9655 1574 9689
rect 3356 7145 3390 7179
rect 2978 6961 3012 6995
rect 3346 6961 3380 6995
rect 2878 4317 2912 4351
rect 3256 4133 3290 4167
rect 2878 1489 2912 1523
rect 3624 1489 3658 1523
rect 52 1397 86 1431
rect 188 1397 222 1431
rect 324 1397 358 1431
rect 460 1397 494 1431
rect 596 1397 630 1431
rect 732 1397 766 1431
rect 868 1397 902 1431
rect 1004 1397 1038 1431
rect 1470 1305 1504 1339
rect 1838 1305 1872 1339
rect 2878 1305 2912 1339
<< poly >>
rect 224 18673 254 18699
rect 592 18673 622 18699
rect 960 18673 990 18699
rect 1328 18673 1358 18699
rect 1696 18673 1726 18699
rect 224 18159 254 18449
rect 592 18159 622 18449
rect 960 18159 990 18449
rect 1328 18159 1358 18449
rect 1696 18159 1726 18449
rect 224 18143 320 18159
rect 224 18109 270 18143
rect 304 18109 320 18143
rect 224 18093 320 18109
rect 592 18143 688 18159
rect 592 18109 638 18143
rect 672 18109 688 18143
rect 592 18093 688 18109
rect 960 18143 1056 18159
rect 960 18109 1006 18143
rect 1040 18109 1056 18143
rect 960 18093 1056 18109
rect 1328 18143 1424 18159
rect 1328 18109 1374 18143
rect 1408 18109 1424 18143
rect 1328 18093 1424 18109
rect 1696 18143 1792 18159
rect 1696 18109 1742 18143
rect 1776 18109 1792 18143
rect 1696 18093 1792 18109
rect 224 17727 254 18093
rect 592 17727 622 18093
rect 960 17727 990 18093
rect 1328 17727 1358 18093
rect 1696 17727 1726 18093
rect 224 17629 254 17655
rect 592 17629 622 17655
rect 960 17629 990 17655
rect 1328 17629 1358 17655
rect 1696 17629 1726 17655
rect 224 17553 254 17579
rect 592 17553 622 17579
rect 960 17553 990 17579
rect 1328 17553 1358 17579
rect 1696 17553 1726 17579
rect 224 17115 254 17481
rect 592 17115 622 17481
rect 960 17115 990 17481
rect 1328 17115 1358 17481
rect 1696 17115 1726 17481
rect 224 17099 320 17115
rect 224 17065 270 17099
rect 304 17065 320 17099
rect 224 17049 320 17065
rect 592 17099 688 17115
rect 592 17065 638 17099
rect 672 17065 688 17099
rect 592 17049 688 17065
rect 960 17099 1056 17115
rect 960 17065 1006 17099
rect 1040 17065 1056 17099
rect 960 17049 1056 17065
rect 1328 17099 1424 17115
rect 1328 17065 1374 17099
rect 1408 17065 1424 17099
rect 1328 17049 1424 17065
rect 1696 17099 1792 17115
rect 1696 17065 1742 17099
rect 1776 17065 1792 17099
rect 1696 17049 1792 17065
rect 224 16759 254 17049
rect 592 16759 622 17049
rect 960 16759 990 17049
rect 1328 16759 1358 17049
rect 1696 16759 1726 17049
rect 224 16509 254 16535
rect 592 16509 622 16535
rect 960 16509 990 16535
rect 1328 16509 1358 16535
rect 1696 16509 1726 16535
rect 224 16433 254 16459
rect 592 16433 622 16459
rect 960 16433 990 16459
rect 1328 16433 1358 16459
rect 1696 16433 1726 16459
rect 224 15919 254 16209
rect 592 15919 622 16209
rect 960 15919 990 16209
rect 1328 15919 1358 16209
rect 1696 15919 1726 16209
rect 224 15903 320 15919
rect 224 15869 270 15903
rect 304 15869 320 15903
rect 224 15853 320 15869
rect 592 15903 688 15919
rect 592 15869 638 15903
rect 672 15869 688 15903
rect 592 15853 688 15869
rect 960 15903 1056 15919
rect 960 15869 1006 15903
rect 1040 15869 1056 15903
rect 960 15853 1056 15869
rect 1328 15903 1424 15919
rect 1328 15869 1374 15903
rect 1408 15869 1424 15903
rect 1328 15853 1424 15869
rect 1696 15903 1792 15919
rect 1696 15869 1742 15903
rect 1776 15869 1792 15903
rect 1696 15853 1792 15869
rect 224 15487 254 15853
rect 592 15487 622 15853
rect 960 15487 990 15853
rect 1328 15487 1358 15853
rect 1696 15487 1726 15853
rect 224 15389 254 15415
rect 592 15389 622 15415
rect 960 15389 990 15415
rect 1328 15389 1358 15415
rect 1696 15389 1726 15415
rect 224 15313 254 15339
rect 592 15313 622 15339
rect 960 15313 990 15339
rect 1328 15313 1358 15339
rect 1696 15313 1726 15339
rect 224 14875 254 15241
rect 592 14875 622 15241
rect 960 14875 990 15241
rect 1328 14875 1358 15241
rect 1696 14875 1726 15241
rect 224 14859 320 14875
rect 224 14825 270 14859
rect 304 14825 320 14859
rect 224 14809 320 14825
rect 592 14859 688 14875
rect 592 14825 638 14859
rect 672 14825 688 14859
rect 592 14809 688 14825
rect 960 14859 1056 14875
rect 960 14825 1006 14859
rect 1040 14825 1056 14859
rect 960 14809 1056 14825
rect 1328 14859 1424 14875
rect 1328 14825 1374 14859
rect 1408 14825 1424 14859
rect 1328 14809 1424 14825
rect 1696 14859 1792 14875
rect 1696 14825 1742 14859
rect 1776 14825 1792 14859
rect 1696 14809 1792 14825
rect 224 14519 254 14809
rect 592 14519 622 14809
rect 960 14519 990 14809
rect 1328 14519 1358 14809
rect 1696 14519 1726 14809
rect 224 14269 254 14295
rect 592 14269 622 14295
rect 960 14269 990 14295
rect 1328 14269 1358 14295
rect 1696 14269 1726 14295
rect 224 14193 254 14219
rect 592 14193 622 14219
rect 960 14193 990 14219
rect 1328 14193 1358 14219
rect 1696 14193 1726 14219
rect 224 13679 254 13969
rect 592 13679 622 13969
rect 960 13679 990 13969
rect 1328 13679 1358 13969
rect 1696 13679 1726 13969
rect 224 13663 320 13679
rect 224 13629 270 13663
rect 304 13629 320 13663
rect 224 13613 320 13629
rect 592 13663 688 13679
rect 592 13629 638 13663
rect 672 13629 688 13663
rect 592 13613 688 13629
rect 960 13663 1056 13679
rect 960 13629 1006 13663
rect 1040 13629 1056 13663
rect 960 13613 1056 13629
rect 1328 13663 1424 13679
rect 1328 13629 1374 13663
rect 1408 13629 1424 13663
rect 1328 13613 1424 13629
rect 1696 13663 1792 13679
rect 1696 13629 1742 13663
rect 1776 13629 1792 13663
rect 1696 13613 1792 13629
rect 224 13247 254 13613
rect 592 13247 622 13613
rect 960 13247 990 13613
rect 1328 13247 1358 13613
rect 1696 13247 1726 13613
rect 224 13149 254 13175
rect 592 13149 622 13175
rect 960 13149 990 13175
rect 1328 13149 1358 13175
rect 1696 13149 1726 13175
rect 224 13073 254 13099
rect 592 13073 622 13099
rect 960 13073 990 13099
rect 1328 13073 1358 13099
rect 1696 13073 1726 13099
rect 224 12635 254 13001
rect 592 12635 622 13001
rect 960 12635 990 13001
rect 1328 12635 1358 13001
rect 1696 12635 1726 13001
rect 224 12619 320 12635
rect 224 12585 270 12619
rect 304 12585 320 12619
rect 224 12569 320 12585
rect 592 12619 688 12635
rect 592 12585 638 12619
rect 672 12585 688 12619
rect 592 12569 688 12585
rect 960 12619 1056 12635
rect 960 12585 1006 12619
rect 1040 12585 1056 12619
rect 960 12569 1056 12585
rect 1328 12619 1424 12635
rect 1328 12585 1374 12619
rect 1408 12585 1424 12619
rect 1328 12569 1424 12585
rect 1696 12619 1792 12635
rect 1696 12585 1742 12619
rect 1776 12585 1792 12619
rect 1696 12569 1792 12585
rect 224 12279 254 12569
rect 592 12279 622 12569
rect 960 12279 990 12569
rect 1328 12279 1358 12569
rect 1696 12279 1726 12569
rect 224 12029 254 12055
rect 592 12029 622 12055
rect 960 12029 990 12055
rect 1328 12029 1358 12055
rect 1696 12029 1726 12055
rect 224 11953 254 11979
rect 592 11953 622 11979
rect 960 11953 990 11979
rect 1328 11953 1358 11979
rect 1696 11953 1726 11979
rect 224 11439 254 11729
rect 592 11439 622 11729
rect 960 11439 990 11729
rect 1328 11439 1358 11729
rect 1696 11439 1726 11729
rect 224 11423 320 11439
rect 224 11389 270 11423
rect 304 11389 320 11423
rect 224 11373 320 11389
rect 592 11423 688 11439
rect 592 11389 638 11423
rect 672 11389 688 11423
rect 592 11373 688 11389
rect 960 11423 1056 11439
rect 960 11389 1006 11423
rect 1040 11389 1056 11423
rect 960 11373 1056 11389
rect 1328 11423 1424 11439
rect 1328 11389 1374 11423
rect 1408 11389 1424 11423
rect 1328 11373 1424 11389
rect 1696 11423 1792 11439
rect 1696 11389 1742 11423
rect 1776 11389 1792 11423
rect 1696 11373 1792 11389
rect 224 11007 254 11373
rect 592 11007 622 11373
rect 960 11007 990 11373
rect 1328 11007 1358 11373
rect 1696 11007 1726 11373
rect 224 10909 254 10935
rect 592 10909 622 10935
rect 960 10909 990 10935
rect 1328 10909 1358 10935
rect 1696 10909 1726 10935
rect 224 10833 254 10859
rect 592 10833 622 10859
rect 960 10833 990 10859
rect 1328 10833 1358 10859
rect 1696 10833 1726 10859
rect 224 10395 254 10761
rect 592 10395 622 10761
rect 960 10395 990 10761
rect 1328 10395 1358 10761
rect 1696 10395 1726 10761
rect 224 10379 320 10395
rect 224 10345 270 10379
rect 304 10345 320 10379
rect 224 10329 320 10345
rect 592 10379 688 10395
rect 592 10345 638 10379
rect 672 10345 688 10379
rect 592 10329 688 10345
rect 960 10379 1056 10395
rect 960 10345 1006 10379
rect 1040 10345 1056 10379
rect 960 10329 1056 10345
rect 1328 10379 1424 10395
rect 1328 10345 1374 10379
rect 1408 10345 1424 10379
rect 1328 10329 1424 10345
rect 1696 10379 1792 10395
rect 1696 10345 1742 10379
rect 1776 10345 1792 10379
rect 1696 10329 1792 10345
rect 224 10039 254 10329
rect 592 10039 622 10329
rect 960 10039 990 10329
rect 1328 10039 1358 10329
rect 1696 10039 1726 10329
rect 224 9789 254 9815
rect 592 9789 622 9815
rect 960 9789 990 9815
rect 1328 9789 1358 9815
rect 1696 9789 1726 9815
rect 224 9713 254 9739
rect 592 9713 622 9739
rect 960 9713 990 9739
rect 1328 9713 1358 9739
rect 1696 9713 1726 9739
rect 224 9199 254 9489
rect 592 9199 622 9489
rect 960 9199 990 9489
rect 1328 9199 1358 9489
rect 1696 9199 1726 9489
rect 224 9183 320 9199
rect 224 9149 270 9183
rect 304 9149 320 9183
rect 224 9133 320 9149
rect 592 9183 688 9199
rect 592 9149 638 9183
rect 672 9149 688 9183
rect 592 9133 688 9149
rect 960 9183 1056 9199
rect 960 9149 1006 9183
rect 1040 9149 1056 9183
rect 960 9133 1056 9149
rect 1328 9183 1424 9199
rect 1328 9149 1374 9183
rect 1408 9149 1424 9183
rect 1328 9133 1424 9149
rect 1696 9183 1792 9199
rect 1696 9149 1742 9183
rect 1776 9149 1792 9183
rect 1696 9133 1792 9149
rect 224 8767 254 9133
rect 592 8767 622 9133
rect 960 8767 990 9133
rect 1328 8767 1358 9133
rect 1696 8767 1726 9133
rect 224 8669 254 8695
rect 592 8669 622 8695
rect 960 8669 990 8695
rect 1328 8669 1358 8695
rect 1696 8669 1726 8695
rect 2726 8433 2756 8459
rect 2826 8433 2856 8459
rect 2926 8433 2956 8459
rect 3204 8433 3234 8459
rect 2726 8247 2756 8285
rect 2675 8231 2756 8247
rect 2675 8197 2691 8231
rect 2725 8197 2756 8231
rect 2675 8181 2756 8197
rect 2726 7345 2756 8181
rect 2826 8123 2856 8285
rect 2808 8107 2874 8123
rect 2808 8073 2824 8107
rect 2858 8073 2874 8107
rect 2808 8057 2874 8073
rect 2826 7345 2856 8057
rect 2926 7999 2956 8285
rect 2926 7983 3007 7999
rect 2926 7949 2957 7983
rect 2991 7949 3007 7983
rect 2926 7933 3007 7949
rect 2926 7345 2956 7933
rect 3204 7810 3234 8033
rect 3138 7794 3234 7810
rect 3138 7760 3154 7794
rect 3188 7760 3234 7794
rect 3138 7744 3234 7760
rect 3204 7521 3234 7744
rect 2726 7095 2756 7121
rect 2826 7095 2856 7121
rect 2926 7095 2956 7121
rect 3204 7095 3234 7121
rect 2726 7019 2756 7045
rect 2826 7019 2856 7045
rect 3194 7019 3224 7045
rect 3562 7019 3592 7045
rect 3820 7019 3850 7045
rect 4078 7019 4108 7045
rect 2726 5959 2756 6795
rect 2826 6207 2856 6795
rect 3194 6358 3224 6795
rect 3562 6377 3592 6795
rect 3128 6342 3224 6358
rect 3128 6308 3144 6342
rect 3178 6308 3224 6342
rect 3496 6361 3592 6377
rect 3496 6327 3512 6361
rect 3546 6327 3592 6361
rect 3820 6359 3850 6619
rect 4078 6396 4108 6619
rect 3496 6311 3592 6327
rect 3128 6292 3224 6308
rect 2808 6191 2874 6207
rect 2808 6157 2824 6191
rect 2858 6157 2874 6191
rect 2808 6141 2874 6157
rect 2708 5943 2774 5959
rect 2708 5909 2724 5943
rect 2758 5909 2774 5943
rect 2708 5893 2774 5909
rect 2726 5855 2756 5893
rect 2826 5855 2856 6141
rect 3194 5779 3224 6292
rect 3562 5855 3592 6311
rect 3754 6343 3850 6359
rect 3754 6309 3770 6343
rect 3804 6309 3850 6343
rect 4012 6380 4108 6396
rect 4012 6346 4028 6380
rect 4062 6346 4108 6380
rect 4012 6330 4108 6346
rect 3754 6293 3850 6309
rect 3820 5959 3850 6293
rect 4078 6107 4108 6330
rect 2726 5681 2756 5707
rect 2826 5681 2856 5707
rect 3194 5681 3224 5707
rect 3562 5681 3592 5707
rect 3820 5681 3850 5707
rect 4078 5681 4108 5707
rect 2726 5605 2756 5631
rect 3352 5605 3382 5631
rect 3610 5605 3640 5631
rect 3868 5605 3898 5631
rect 4126 5605 4156 5631
rect 2726 5020 2756 5533
rect 3094 5529 3124 5555
rect 3094 5020 3124 5457
rect 2660 5004 2756 5020
rect 2660 4970 2676 5004
rect 2710 4970 2756 5004
rect 2660 4954 2756 4970
rect 3028 5004 3124 5020
rect 3028 4970 3044 5004
rect 3078 4970 3124 5004
rect 3352 5001 3382 5457
rect 3028 4954 3124 4970
rect 2726 4517 2756 4954
rect 3094 4517 3124 4954
rect 3286 4985 3382 5001
rect 3286 4951 3302 4985
rect 3336 4951 3382 4985
rect 3610 4982 3640 5205
rect 3868 4998 3898 5269
rect 3286 4935 3382 4951
rect 3352 4517 3382 4935
rect 3544 4966 3640 4982
rect 3544 4932 3560 4966
rect 3594 4932 3640 4966
rect 3802 4982 3898 4998
rect 4126 4982 4156 5205
rect 3802 4948 3818 4982
rect 3852 4948 3898 4982
rect 3802 4932 3898 4948
rect 3544 4916 3640 4932
rect 3610 4693 3640 4916
rect 3868 4693 3898 4932
rect 4060 4966 4156 4982
rect 4060 4932 4076 4966
rect 4110 4932 4156 4966
rect 4060 4916 4156 4932
rect 4126 4693 4156 4916
rect 2726 4267 2756 4293
rect 3094 4267 3124 4293
rect 3352 4267 3382 4293
rect 3610 4267 3640 4293
rect 3868 4267 3898 4293
rect 4126 4267 4156 4293
rect 2726 4191 2756 4217
rect 2826 4191 2856 4217
rect 3104 4191 3134 4217
rect 2726 3131 2756 3967
rect 2826 3379 2856 3967
rect 3104 3552 3134 3791
rect 3038 3536 3134 3552
rect 3038 3502 3054 3536
rect 3088 3502 3134 3536
rect 3038 3486 3134 3502
rect 2808 3363 2874 3379
rect 2808 3329 2824 3363
rect 2858 3329 2874 3363
rect 2808 3313 2874 3329
rect 2708 3115 2774 3131
rect 2708 3081 2724 3115
rect 2758 3081 2774 3115
rect 2708 3065 2774 3081
rect 2726 3027 2756 3065
rect 2826 3027 2856 3313
rect 3104 3215 3134 3486
rect 2726 2853 2756 2879
rect 2826 2853 2856 2879
rect 3104 2853 3134 2879
rect 2726 2777 2756 2803
rect 3094 2777 3124 2803
rect 3194 2777 3224 2803
rect 3472 2777 3502 2803
rect 2726 2192 2756 2705
rect 3094 2591 3124 2629
rect 3076 2575 3142 2591
rect 3076 2541 3092 2575
rect 3126 2541 3142 2575
rect 3076 2525 3142 2541
rect 2660 2176 2756 2192
rect 2660 2142 2676 2176
rect 2710 2142 2756 2176
rect 2660 2126 2756 2142
rect 2726 1689 2756 2126
rect 3094 1689 3124 2525
rect 3194 2343 3224 2629
rect 3176 2327 3242 2343
rect 3176 2293 3192 2327
rect 3226 2293 3242 2327
rect 3176 2277 3242 2293
rect 3194 1689 3224 2277
rect 3472 2170 3502 2441
rect 3406 2154 3502 2170
rect 3406 2120 3422 2154
rect 3456 2120 3502 2154
rect 3406 2104 3502 2120
rect 3472 1865 3502 2104
rect 2726 1439 2756 1465
rect 3094 1439 3124 1465
rect 3194 1439 3224 1465
rect 3472 1439 3502 1465
rect 1318 1363 1348 1389
rect 1686 1363 1716 1389
rect 2726 1363 2756 1389
rect 3094 1363 3124 1389
rect 3352 1363 3382 1389
rect 3610 1363 3640 1389
rect 3868 1363 3898 1389
rect 4126 1363 4156 1389
rect 81 1312 111 1338
rect 167 1312 197 1338
rect 239 1312 269 1338
rect 359 1312 389 1338
rect 431 1312 461 1338
rect 517 1312 547 1338
rect 589 1312 619 1338
rect 709 1312 739 1338
rect 781 1312 811 1338
rect 867 1312 897 1338
rect 1057 1312 1087 1338
rect 1318 721 1348 1139
rect 1686 742 1716 1033
rect 81 697 111 712
rect 70 677 111 697
rect 47 667 111 677
rect 47 661 101 667
rect 47 627 57 661
rect 91 627 101 661
rect 47 611 101 627
rect 71 447 101 611
rect 167 597 197 712
rect 239 672 269 712
rect 239 656 293 672
rect 239 622 249 656
rect 283 622 293 656
rect 239 606 293 622
rect 143 581 197 597
rect 143 547 153 581
rect 187 547 197 581
rect 143 531 197 547
rect 359 531 389 712
rect 431 667 461 712
rect 517 667 547 712
rect 431 657 547 667
rect 431 623 472 657
rect 506 623 547 657
rect 431 613 547 623
rect 589 531 619 712
rect 709 672 739 712
rect 685 656 739 672
rect 685 622 695 656
rect 729 622 739 656
rect 685 606 739 622
rect 781 597 811 712
rect 867 677 897 712
rect 867 661 938 677
rect 867 647 894 661
rect 878 627 894 647
rect 928 627 938 661
rect 878 611 938 627
rect 781 581 835 597
rect 781 547 791 581
rect 825 547 835 581
rect 781 531 835 547
rect 71 417 111 447
rect 81 302 111 417
rect 167 302 197 531
rect 239 501 739 531
rect 239 302 269 501
rect 685 467 695 501
rect 729 467 739 501
rect 685 451 739 467
rect 335 421 389 437
rect 335 387 345 421
rect 379 387 389 421
rect 335 371 389 387
rect 359 302 389 371
rect 431 421 547 431
rect 431 387 472 421
rect 506 387 547 421
rect 431 377 547 387
rect 431 302 461 377
rect 517 302 547 377
rect 589 421 643 437
rect 589 387 599 421
rect 633 387 643 421
rect 589 371 643 387
rect 589 302 619 371
rect 709 302 739 451
rect 781 302 811 531
rect 878 481 908 611
rect 1057 517 1087 712
rect 1252 705 1348 721
rect 1252 671 1268 705
rect 1302 671 1348 705
rect 1620 726 1716 742
rect 1620 692 1636 726
rect 1670 692 1716 726
rect 2726 702 2756 1139
rect 3094 702 3124 1139
rect 3352 720 3382 1033
rect 3610 724 3640 963
rect 3868 740 3898 963
rect 4126 740 4156 963
rect 1620 676 1716 692
rect 1252 655 1348 671
rect 867 371 908 481
rect 1033 501 1087 517
rect 1033 467 1043 501
rect 1077 467 1087 501
rect 1033 451 1087 467
rect 867 302 897 371
rect 1057 302 1087 451
rect 1318 199 1348 655
rect 1686 387 1716 676
rect 2660 686 2756 702
rect 2660 652 2676 686
rect 2710 652 2756 686
rect 2660 636 2756 652
rect 3028 686 3124 702
rect 3028 652 3044 686
rect 3078 652 3124 686
rect 3286 704 3382 720
rect 3286 670 3302 704
rect 3336 670 3382 704
rect 3286 654 3382 670
rect 3544 708 3640 724
rect 3544 674 3560 708
rect 3594 674 3640 708
rect 3802 724 3898 740
rect 3802 690 3818 724
rect 3852 690 3898 724
rect 3802 674 3898 690
rect 4060 724 4156 740
rect 4060 690 4076 724
rect 4110 690 4156 724
rect 4060 674 4156 690
rect 3544 658 3640 674
rect 3028 636 3124 652
rect 81 76 111 102
rect 167 76 197 102
rect 239 76 269 102
rect 359 76 389 102
rect 431 76 461 102
rect 517 76 547 102
rect 589 76 619 102
rect 709 76 739 102
rect 781 76 811 102
rect 867 76 897 102
rect 1057 76 1087 102
rect 2726 123 2756 636
rect 3094 123 3124 636
rect 3352 303 3382 654
rect 3610 387 3640 658
rect 3868 451 3898 674
rect 4126 451 4156 674
rect 1318 25 1348 51
rect 1686 25 1716 51
rect 2726 25 2756 51
rect 3094 25 3124 51
rect 3352 25 3382 51
rect 3610 25 3640 51
rect 3868 25 3898 51
rect 4126 25 4156 51
<< polycont >>
rect 270 18109 304 18143
rect 638 18109 672 18143
rect 1006 18109 1040 18143
rect 1374 18109 1408 18143
rect 1742 18109 1776 18143
rect 270 17065 304 17099
rect 638 17065 672 17099
rect 1006 17065 1040 17099
rect 1374 17065 1408 17099
rect 1742 17065 1776 17099
rect 270 15869 304 15903
rect 638 15869 672 15903
rect 1006 15869 1040 15903
rect 1374 15869 1408 15903
rect 1742 15869 1776 15903
rect 270 14825 304 14859
rect 638 14825 672 14859
rect 1006 14825 1040 14859
rect 1374 14825 1408 14859
rect 1742 14825 1776 14859
rect 270 13629 304 13663
rect 638 13629 672 13663
rect 1006 13629 1040 13663
rect 1374 13629 1408 13663
rect 1742 13629 1776 13663
rect 270 12585 304 12619
rect 638 12585 672 12619
rect 1006 12585 1040 12619
rect 1374 12585 1408 12619
rect 1742 12585 1776 12619
rect 270 11389 304 11423
rect 638 11389 672 11423
rect 1006 11389 1040 11423
rect 1374 11389 1408 11423
rect 1742 11389 1776 11423
rect 270 10345 304 10379
rect 638 10345 672 10379
rect 1006 10345 1040 10379
rect 1374 10345 1408 10379
rect 1742 10345 1776 10379
rect 270 9149 304 9183
rect 638 9149 672 9183
rect 1006 9149 1040 9183
rect 1374 9149 1408 9183
rect 1742 9149 1776 9183
rect 2691 8197 2725 8231
rect 2824 8073 2858 8107
rect 2957 7949 2991 7983
rect 3154 7760 3188 7794
rect 3144 6308 3178 6342
rect 3512 6327 3546 6361
rect 2824 6157 2858 6191
rect 2724 5909 2758 5943
rect 3770 6309 3804 6343
rect 4028 6346 4062 6380
rect 2676 4970 2710 5004
rect 3044 4970 3078 5004
rect 3302 4951 3336 4985
rect 3560 4932 3594 4966
rect 3818 4948 3852 4982
rect 4076 4932 4110 4966
rect 3054 3502 3088 3536
rect 2824 3329 2858 3363
rect 2724 3081 2758 3115
rect 3092 2541 3126 2575
rect 2676 2142 2710 2176
rect 3192 2293 3226 2327
rect 3422 2120 3456 2154
rect 57 627 91 661
rect 249 622 283 656
rect 153 547 187 581
rect 472 623 506 657
rect 695 622 729 656
rect 894 627 928 661
rect 791 547 825 581
rect 695 467 729 501
rect 345 387 379 421
rect 472 387 506 421
rect 599 387 633 421
rect 1268 671 1302 705
rect 1636 692 1670 726
rect 1043 467 1077 501
rect 2676 652 2710 686
rect 3044 652 3078 686
rect 3302 670 3336 704
rect 3560 674 3594 708
rect 3818 690 3852 724
rect 4076 690 4110 724
<< locali >>
rect 431 18741 465 18757
rect 1167 18741 1201 18757
rect 0 18707 431 18741
rect 465 18707 1167 18741
rect 1201 18707 1840 18741
rect 68 18649 102 18707
rect 68 18599 102 18615
rect 172 18578 206 18594
rect 172 18143 206 18544
rect 272 18578 306 18707
rect 431 18691 470 18707
rect 436 18649 470 18691
rect 436 18599 470 18615
rect 272 18528 306 18544
rect 540 18578 574 18594
rect 155 18109 206 18143
rect 68 17713 102 17729
rect 68 17621 102 17679
rect 172 17708 206 18109
rect 270 18143 304 18159
rect 540 18143 574 18544
rect 640 18578 674 18707
rect 804 18649 838 18707
rect 804 18599 838 18615
rect 640 18528 674 18544
rect 908 18578 942 18594
rect 523 18109 574 18143
rect 270 18093 304 18109
rect 172 17658 206 17674
rect 272 17708 306 17724
rect 272 17621 306 17674
rect 436 17713 470 17729
rect 436 17637 470 17679
rect 540 17708 574 18109
rect 638 18143 672 18159
rect 908 18143 942 18544
rect 1008 18578 1042 18707
rect 1167 18691 1206 18707
rect 1172 18649 1206 18691
rect 1172 18599 1206 18615
rect 1008 18528 1042 18544
rect 1276 18578 1310 18594
rect 891 18109 942 18143
rect 638 18093 672 18109
rect 540 17658 574 17674
rect 640 17708 674 17724
rect 431 17621 470 17637
rect 640 17621 674 17674
rect 804 17713 838 17729
rect 804 17621 838 17679
rect 908 17708 942 18109
rect 1006 18143 1040 18159
rect 1276 18143 1310 18544
rect 1376 18578 1410 18707
rect 1540 18649 1574 18707
rect 1540 18599 1574 18615
rect 1376 18528 1410 18544
rect 1644 18578 1678 18594
rect 1644 18159 1678 18544
rect 1744 18578 1778 18707
rect 1744 18528 1778 18544
rect 1259 18109 1310 18143
rect 1006 18093 1040 18109
rect 908 17658 942 17674
rect 1008 17708 1042 17724
rect 1008 17621 1042 17674
rect 1172 17713 1206 17729
rect 1172 17637 1206 17679
rect 1276 17708 1310 18109
rect 1374 18143 1408 18159
rect 1374 18093 1408 18109
rect 1627 18143 1678 18159
rect 1661 18109 1678 18143
rect 1627 18093 1678 18109
rect 1742 18143 1776 18159
rect 1742 18093 1776 18109
rect 1276 17658 1310 17674
rect 1376 17708 1410 17724
rect 1167 17621 1206 17637
rect 1376 17621 1410 17674
rect 1540 17713 1574 17729
rect 1540 17621 1574 17679
rect 1644 17708 1678 18093
rect 1644 17658 1678 17674
rect 1744 17708 1778 17724
rect 1744 17621 1778 17674
rect 0 17587 431 17621
rect 465 17587 1167 17621
rect 1201 17587 1840 17621
rect 68 17529 102 17587
rect 68 17479 102 17495
rect 172 17534 206 17550
rect 172 17099 206 17500
rect 272 17534 306 17587
rect 431 17571 470 17587
rect 272 17484 306 17500
rect 436 17529 470 17571
rect 436 17479 470 17495
rect 540 17534 574 17550
rect 155 17065 206 17099
rect 172 16664 206 17065
rect 270 17099 304 17115
rect 540 17099 574 17500
rect 640 17534 674 17587
rect 640 17484 674 17500
rect 804 17529 838 17587
rect 804 17479 838 17495
rect 908 17534 942 17550
rect 523 17065 574 17099
rect 270 17049 304 17065
rect 172 16614 206 16630
rect 272 16664 306 16680
rect 68 16593 102 16609
rect 68 16501 102 16559
rect 272 16501 306 16630
rect 540 16664 574 17065
rect 638 17099 672 17115
rect 908 17099 942 17500
rect 1008 17534 1042 17587
rect 1167 17571 1206 17587
rect 1008 17484 1042 17500
rect 1172 17529 1206 17571
rect 1172 17479 1206 17495
rect 1276 17534 1310 17550
rect 891 17065 942 17099
rect 638 17049 672 17065
rect 540 16614 574 16630
rect 640 16664 674 16680
rect 436 16593 470 16609
rect 436 16517 470 16559
rect 431 16501 470 16517
rect 640 16501 674 16630
rect 908 16664 942 17065
rect 1006 17099 1040 17115
rect 1276 17099 1310 17500
rect 1376 17534 1410 17587
rect 1376 17484 1410 17500
rect 1540 17529 1574 17587
rect 1540 17479 1574 17495
rect 1644 17534 1678 17550
rect 1644 17115 1678 17500
rect 1744 17534 1778 17587
rect 1744 17484 1778 17500
rect 1259 17065 1310 17099
rect 1006 17049 1040 17065
rect 908 16614 942 16630
rect 1008 16664 1042 16680
rect 804 16593 838 16609
rect 804 16501 838 16559
rect 1008 16501 1042 16630
rect 1276 16664 1310 17065
rect 1374 17099 1408 17115
rect 1374 17049 1408 17065
rect 1627 17099 1678 17115
rect 1661 17065 1678 17099
rect 1627 17049 1678 17065
rect 1742 17099 1776 17115
rect 1742 17049 1776 17065
rect 1276 16614 1310 16630
rect 1376 16664 1410 16680
rect 1172 16593 1206 16609
rect 1172 16517 1206 16559
rect 1167 16501 1206 16517
rect 1376 16501 1410 16630
rect 1644 16664 1678 17049
rect 1644 16614 1678 16630
rect 1744 16664 1778 16680
rect 1540 16593 1574 16609
rect 1540 16501 1574 16559
rect 1744 16501 1778 16630
rect 0 16467 431 16501
rect 465 16467 1167 16501
rect 1201 16467 1840 16501
rect 68 16409 102 16467
rect 68 16359 102 16375
rect 172 16338 206 16354
rect 172 15903 206 16304
rect 272 16338 306 16467
rect 431 16451 470 16467
rect 436 16409 470 16451
rect 436 16359 470 16375
rect 272 16288 306 16304
rect 540 16338 574 16354
rect 155 15869 206 15903
rect 68 15473 102 15489
rect 68 15381 102 15439
rect 172 15468 206 15869
rect 270 15903 304 15919
rect 540 15903 574 16304
rect 640 16338 674 16467
rect 804 16409 838 16467
rect 804 16359 838 16375
rect 640 16288 674 16304
rect 908 16338 942 16354
rect 523 15869 574 15903
rect 270 15853 304 15869
rect 172 15418 206 15434
rect 272 15468 306 15484
rect 272 15381 306 15434
rect 436 15473 470 15489
rect 436 15397 470 15439
rect 540 15468 574 15869
rect 638 15903 672 15919
rect 908 15903 942 16304
rect 1008 16338 1042 16467
rect 1167 16451 1206 16467
rect 1172 16409 1206 16451
rect 1172 16359 1206 16375
rect 1008 16288 1042 16304
rect 1276 16338 1310 16354
rect 891 15869 942 15903
rect 638 15853 672 15869
rect 540 15418 574 15434
rect 640 15468 674 15484
rect 431 15381 470 15397
rect 640 15381 674 15434
rect 804 15473 838 15489
rect 804 15381 838 15439
rect 908 15468 942 15869
rect 1006 15903 1040 15919
rect 1276 15903 1310 16304
rect 1376 16338 1410 16467
rect 1540 16409 1574 16467
rect 1540 16359 1574 16375
rect 1376 16288 1410 16304
rect 1644 16338 1678 16354
rect 1644 15919 1678 16304
rect 1744 16338 1778 16467
rect 1744 16288 1778 16304
rect 1259 15869 1310 15903
rect 1006 15853 1040 15869
rect 908 15418 942 15434
rect 1008 15468 1042 15484
rect 1008 15381 1042 15434
rect 1172 15473 1206 15489
rect 1172 15397 1206 15439
rect 1276 15468 1310 15869
rect 1374 15903 1408 15919
rect 1374 15853 1408 15869
rect 1627 15903 1678 15919
rect 1661 15869 1678 15903
rect 1627 15853 1678 15869
rect 1742 15903 1776 15919
rect 1742 15853 1776 15869
rect 1276 15418 1310 15434
rect 1376 15468 1410 15484
rect 1167 15381 1206 15397
rect 1376 15381 1410 15434
rect 1540 15473 1574 15489
rect 1540 15381 1574 15439
rect 1644 15468 1678 15853
rect 1644 15418 1678 15434
rect 1744 15468 1778 15484
rect 1744 15381 1778 15434
rect 0 15347 431 15381
rect 465 15347 1167 15381
rect 1201 15347 1840 15381
rect 68 15289 102 15347
rect 68 15239 102 15255
rect 172 15294 206 15310
rect 172 14859 206 15260
rect 272 15294 306 15347
rect 431 15331 470 15347
rect 272 15244 306 15260
rect 436 15289 470 15331
rect 436 15239 470 15255
rect 540 15294 574 15310
rect 155 14825 206 14859
rect 172 14424 206 14825
rect 270 14859 304 14875
rect 540 14859 574 15260
rect 640 15294 674 15347
rect 640 15244 674 15260
rect 804 15289 838 15347
rect 804 15239 838 15255
rect 908 15294 942 15310
rect 523 14825 574 14859
rect 270 14809 304 14825
rect 172 14374 206 14390
rect 272 14424 306 14440
rect 68 14353 102 14369
rect 68 14261 102 14319
rect 272 14261 306 14390
rect 540 14424 574 14825
rect 638 14859 672 14875
rect 908 14859 942 15260
rect 1008 15294 1042 15347
rect 1167 15331 1206 15347
rect 1008 15244 1042 15260
rect 1172 15289 1206 15331
rect 1172 15239 1206 15255
rect 1276 15294 1310 15310
rect 891 14825 942 14859
rect 638 14809 672 14825
rect 540 14374 574 14390
rect 640 14424 674 14440
rect 436 14353 470 14369
rect 436 14277 470 14319
rect 431 14261 470 14277
rect 640 14261 674 14390
rect 908 14424 942 14825
rect 1006 14859 1040 14875
rect 1276 14859 1310 15260
rect 1376 15294 1410 15347
rect 1376 15244 1410 15260
rect 1540 15289 1574 15347
rect 1540 15239 1574 15255
rect 1644 15294 1678 15310
rect 1644 14875 1678 15260
rect 1744 15294 1778 15347
rect 1744 15244 1778 15260
rect 1259 14825 1310 14859
rect 1006 14809 1040 14825
rect 908 14374 942 14390
rect 1008 14424 1042 14440
rect 804 14353 838 14369
rect 804 14261 838 14319
rect 1008 14261 1042 14390
rect 1276 14424 1310 14825
rect 1374 14859 1408 14875
rect 1374 14809 1408 14825
rect 1627 14859 1678 14875
rect 1661 14825 1678 14859
rect 1627 14809 1678 14825
rect 1742 14859 1776 14875
rect 1742 14809 1776 14825
rect 1276 14374 1310 14390
rect 1376 14424 1410 14440
rect 1172 14353 1206 14369
rect 1172 14277 1206 14319
rect 1167 14261 1206 14277
rect 1376 14261 1410 14390
rect 1644 14424 1678 14809
rect 1644 14374 1678 14390
rect 1744 14424 1778 14440
rect 1540 14353 1574 14369
rect 1540 14261 1574 14319
rect 1744 14261 1778 14390
rect 0 14227 431 14261
rect 465 14227 1167 14261
rect 1201 14227 1840 14261
rect 68 14169 102 14227
rect 68 14119 102 14135
rect 172 14098 206 14114
rect 172 13663 206 14064
rect 272 14098 306 14227
rect 431 14211 470 14227
rect 436 14169 470 14211
rect 436 14119 470 14135
rect 272 14048 306 14064
rect 540 14098 574 14114
rect 155 13629 206 13663
rect 68 13233 102 13249
rect 68 13141 102 13199
rect 172 13228 206 13629
rect 270 13663 304 13679
rect 540 13663 574 14064
rect 640 14098 674 14227
rect 804 14169 838 14227
rect 804 14119 838 14135
rect 640 14048 674 14064
rect 908 14098 942 14114
rect 523 13629 574 13663
rect 270 13613 304 13629
rect 172 13178 206 13194
rect 272 13228 306 13244
rect 272 13141 306 13194
rect 436 13233 470 13249
rect 436 13157 470 13199
rect 540 13228 574 13629
rect 638 13663 672 13679
rect 908 13663 942 14064
rect 1008 14098 1042 14227
rect 1167 14211 1206 14227
rect 1172 14169 1206 14211
rect 1172 14119 1206 14135
rect 1008 14048 1042 14064
rect 1276 14098 1310 14114
rect 891 13629 942 13663
rect 638 13613 672 13629
rect 540 13178 574 13194
rect 640 13228 674 13244
rect 431 13141 470 13157
rect 640 13141 674 13194
rect 804 13233 838 13249
rect 804 13141 838 13199
rect 908 13228 942 13629
rect 1006 13663 1040 13679
rect 1276 13663 1310 14064
rect 1376 14098 1410 14227
rect 1540 14169 1574 14227
rect 1540 14119 1574 14135
rect 1376 14048 1410 14064
rect 1644 14098 1678 14114
rect 1644 13679 1678 14064
rect 1744 14098 1778 14227
rect 1744 14048 1778 14064
rect 1259 13629 1310 13663
rect 1006 13613 1040 13629
rect 908 13178 942 13194
rect 1008 13228 1042 13244
rect 1008 13141 1042 13194
rect 1172 13233 1206 13249
rect 1172 13157 1206 13199
rect 1276 13228 1310 13629
rect 1374 13663 1408 13679
rect 1374 13613 1408 13629
rect 1627 13663 1678 13679
rect 1661 13629 1678 13663
rect 1627 13613 1678 13629
rect 1742 13663 1776 13679
rect 1742 13613 1776 13629
rect 1276 13178 1310 13194
rect 1376 13228 1410 13244
rect 1167 13141 1206 13157
rect 1376 13141 1410 13194
rect 1540 13233 1574 13249
rect 1540 13141 1574 13199
rect 1644 13228 1678 13613
rect 1644 13178 1678 13194
rect 1744 13228 1778 13244
rect 1744 13141 1778 13194
rect 0 13107 431 13141
rect 465 13107 1167 13141
rect 1201 13107 1840 13141
rect 68 13049 102 13107
rect 68 12999 102 13015
rect 172 13054 206 13070
rect 172 12619 206 13020
rect 272 13054 306 13107
rect 431 13091 470 13107
rect 272 13004 306 13020
rect 436 13049 470 13091
rect 436 12999 470 13015
rect 540 13054 574 13070
rect 155 12585 206 12619
rect 172 12184 206 12585
rect 270 12619 304 12635
rect 540 12619 574 13020
rect 640 13054 674 13107
rect 640 13004 674 13020
rect 804 13049 838 13107
rect 804 12999 838 13015
rect 908 13054 942 13070
rect 523 12585 574 12619
rect 270 12569 304 12585
rect 172 12134 206 12150
rect 272 12184 306 12200
rect 68 12113 102 12129
rect 68 12021 102 12079
rect 272 12021 306 12150
rect 540 12184 574 12585
rect 638 12619 672 12635
rect 908 12619 942 13020
rect 1008 13054 1042 13107
rect 1167 13091 1206 13107
rect 1008 13004 1042 13020
rect 1172 13049 1206 13091
rect 1172 12999 1206 13015
rect 1276 13054 1310 13070
rect 891 12585 942 12619
rect 638 12569 672 12585
rect 540 12134 574 12150
rect 640 12184 674 12200
rect 436 12113 470 12129
rect 436 12037 470 12079
rect 431 12021 470 12037
rect 640 12021 674 12150
rect 908 12184 942 12585
rect 1006 12619 1040 12635
rect 1276 12619 1310 13020
rect 1376 13054 1410 13107
rect 1376 13004 1410 13020
rect 1540 13049 1574 13107
rect 1540 12999 1574 13015
rect 1644 13054 1678 13070
rect 1644 12635 1678 13020
rect 1744 13054 1778 13107
rect 1744 13004 1778 13020
rect 1259 12585 1310 12619
rect 1006 12569 1040 12585
rect 908 12134 942 12150
rect 1008 12184 1042 12200
rect 804 12113 838 12129
rect 804 12021 838 12079
rect 1008 12021 1042 12150
rect 1276 12184 1310 12585
rect 1374 12619 1408 12635
rect 1374 12569 1408 12585
rect 1627 12619 1678 12635
rect 1661 12585 1678 12619
rect 1627 12569 1678 12585
rect 1742 12619 1776 12635
rect 1742 12569 1776 12585
rect 1276 12134 1310 12150
rect 1376 12184 1410 12200
rect 1172 12113 1206 12129
rect 1172 12037 1206 12079
rect 1167 12021 1206 12037
rect 1376 12021 1410 12150
rect 1644 12184 1678 12569
rect 1644 12134 1678 12150
rect 1744 12184 1778 12200
rect 1540 12113 1574 12129
rect 1540 12021 1574 12079
rect 1744 12021 1778 12150
rect 0 11987 431 12021
rect 465 11987 1167 12021
rect 1201 11987 1840 12021
rect 68 11929 102 11987
rect 68 11879 102 11895
rect 172 11858 206 11874
rect 172 11423 206 11824
rect 272 11858 306 11987
rect 431 11971 470 11987
rect 436 11929 470 11971
rect 436 11879 470 11895
rect 272 11808 306 11824
rect 540 11858 574 11874
rect 155 11389 206 11423
rect 68 10993 102 11009
rect 68 10901 102 10959
rect 172 10988 206 11389
rect 270 11423 304 11439
rect 540 11423 574 11824
rect 640 11858 674 11987
rect 804 11929 838 11987
rect 804 11879 838 11895
rect 640 11808 674 11824
rect 908 11858 942 11874
rect 523 11389 574 11423
rect 270 11373 304 11389
rect 172 10938 206 10954
rect 272 10988 306 11004
rect 272 10901 306 10954
rect 436 10993 470 11009
rect 436 10917 470 10959
rect 540 10988 574 11389
rect 638 11423 672 11439
rect 908 11423 942 11824
rect 1008 11858 1042 11987
rect 1167 11971 1206 11987
rect 1172 11929 1206 11971
rect 1172 11879 1206 11895
rect 1008 11808 1042 11824
rect 1276 11858 1310 11874
rect 891 11389 942 11423
rect 638 11373 672 11389
rect 540 10938 574 10954
rect 640 10988 674 11004
rect 431 10901 470 10917
rect 640 10901 674 10954
rect 804 10993 838 11009
rect 804 10901 838 10959
rect 908 10988 942 11389
rect 1006 11423 1040 11439
rect 1276 11423 1310 11824
rect 1376 11858 1410 11987
rect 1540 11929 1574 11987
rect 1540 11879 1574 11895
rect 1376 11808 1410 11824
rect 1644 11858 1678 11874
rect 1644 11439 1678 11824
rect 1744 11858 1778 11987
rect 1744 11808 1778 11824
rect 1259 11389 1310 11423
rect 1006 11373 1040 11389
rect 908 10938 942 10954
rect 1008 10988 1042 11004
rect 1008 10901 1042 10954
rect 1172 10993 1206 11009
rect 1172 10917 1206 10959
rect 1276 10988 1310 11389
rect 1374 11423 1408 11439
rect 1374 11373 1408 11389
rect 1627 11423 1678 11439
rect 1661 11389 1678 11423
rect 1627 11373 1678 11389
rect 1742 11423 1776 11439
rect 1742 11373 1776 11389
rect 1276 10938 1310 10954
rect 1376 10988 1410 11004
rect 1167 10901 1206 10917
rect 1376 10901 1410 10954
rect 1540 10993 1574 11009
rect 1540 10901 1574 10959
rect 1644 10988 1678 11373
rect 1644 10938 1678 10954
rect 1744 10988 1778 11004
rect 1744 10901 1778 10954
rect 0 10867 431 10901
rect 465 10867 1167 10901
rect 1201 10867 1840 10901
rect 68 10809 102 10867
rect 68 10759 102 10775
rect 172 10814 206 10830
rect 172 10379 206 10780
rect 272 10814 306 10867
rect 431 10851 470 10867
rect 272 10764 306 10780
rect 436 10809 470 10851
rect 436 10759 470 10775
rect 540 10814 574 10830
rect 155 10345 206 10379
rect 172 9944 206 10345
rect 270 10379 304 10395
rect 540 10379 574 10780
rect 640 10814 674 10867
rect 640 10764 674 10780
rect 804 10809 838 10867
rect 804 10759 838 10775
rect 908 10814 942 10830
rect 523 10345 574 10379
rect 270 10329 304 10345
rect 172 9894 206 9910
rect 272 9944 306 9960
rect 68 9873 102 9889
rect 68 9781 102 9839
rect 272 9781 306 9910
rect 540 9944 574 10345
rect 638 10379 672 10395
rect 908 10379 942 10780
rect 1008 10814 1042 10867
rect 1167 10851 1206 10867
rect 1008 10764 1042 10780
rect 1172 10809 1206 10851
rect 1172 10759 1206 10775
rect 1276 10814 1310 10830
rect 891 10345 942 10379
rect 638 10329 672 10345
rect 540 9894 574 9910
rect 640 9944 674 9960
rect 436 9873 470 9889
rect 436 9797 470 9839
rect 431 9781 470 9797
rect 640 9781 674 9910
rect 908 9944 942 10345
rect 1006 10379 1040 10395
rect 1276 10379 1310 10780
rect 1376 10814 1410 10867
rect 1376 10764 1410 10780
rect 1540 10809 1574 10867
rect 1540 10759 1574 10775
rect 1644 10814 1678 10830
rect 1644 10395 1678 10780
rect 1744 10814 1778 10867
rect 1744 10764 1778 10780
rect 1259 10345 1310 10379
rect 1006 10329 1040 10345
rect 908 9894 942 9910
rect 1008 9944 1042 9960
rect 804 9873 838 9889
rect 804 9781 838 9839
rect 1008 9781 1042 9910
rect 1276 9944 1310 10345
rect 1374 10379 1408 10395
rect 1374 10329 1408 10345
rect 1627 10379 1678 10395
rect 1661 10345 1678 10379
rect 1627 10329 1678 10345
rect 1742 10379 1776 10395
rect 1742 10329 1776 10345
rect 1276 9894 1310 9910
rect 1376 9944 1410 9960
rect 1172 9873 1206 9889
rect 1172 9797 1206 9839
rect 1167 9781 1206 9797
rect 1376 9781 1410 9910
rect 1644 9944 1678 10329
rect 1644 9894 1678 9910
rect 1744 9944 1778 9960
rect 1540 9873 1574 9889
rect 1540 9781 1574 9839
rect 1744 9781 1778 9910
rect 0 9747 431 9781
rect 465 9747 1167 9781
rect 1201 9747 1840 9781
rect 68 9689 102 9747
rect 68 9639 102 9655
rect 172 9618 206 9634
rect 172 9183 206 9584
rect 272 9618 306 9747
rect 431 9731 470 9747
rect 436 9689 470 9731
rect 436 9639 470 9655
rect 272 9568 306 9584
rect 540 9618 574 9634
rect 155 9149 206 9183
rect 68 8753 102 8769
rect 68 8661 102 8719
rect 172 8748 206 9149
rect 270 9183 304 9199
rect 540 9183 574 9584
rect 640 9618 674 9747
rect 804 9689 838 9747
rect 804 9639 838 9655
rect 640 9568 674 9584
rect 908 9618 942 9634
rect 523 9149 574 9183
rect 270 9133 304 9149
rect 172 8698 206 8714
rect 272 8748 306 8764
rect 272 8661 306 8714
rect 436 8753 470 8769
rect 436 8677 470 8719
rect 540 8748 574 9149
rect 638 9183 672 9199
rect 908 9183 942 9584
rect 1008 9618 1042 9747
rect 1167 9731 1206 9747
rect 1172 9689 1206 9731
rect 1172 9639 1206 9655
rect 1008 9568 1042 9584
rect 1276 9618 1310 9634
rect 891 9149 942 9183
rect 638 9133 672 9149
rect 540 8698 574 8714
rect 640 8748 674 8764
rect 431 8661 470 8677
rect 640 8661 674 8714
rect 804 8753 838 8769
rect 804 8661 838 8719
rect 908 8748 942 9149
rect 1006 9183 1040 9199
rect 1276 9183 1310 9584
rect 1376 9618 1410 9747
rect 1540 9689 1574 9747
rect 1540 9639 1574 9655
rect 1376 9568 1410 9584
rect 1644 9618 1678 9634
rect 1644 9199 1678 9584
rect 1744 9618 1778 9747
rect 1744 9568 1778 9584
rect 1259 9149 1310 9183
rect 1006 9133 1040 9149
rect 908 8698 942 8714
rect 1008 8748 1042 8764
rect 1008 8661 1042 8714
rect 1172 8753 1206 8769
rect 1172 8677 1206 8719
rect 1276 8748 1310 9149
rect 1374 9183 1408 9199
rect 1374 9133 1408 9149
rect 1627 9183 1678 9199
rect 1661 9149 1678 9183
rect 1627 9133 1678 9149
rect 1742 9183 1776 9199
rect 1742 9133 1776 9149
rect 1276 8698 1310 8714
rect 1376 8748 1410 8764
rect 1167 8661 1206 8677
rect 1376 8661 1410 8714
rect 1540 8753 1574 8769
rect 1540 8661 1574 8719
rect 1644 8748 1678 9133
rect 1644 8698 1678 8714
rect 1744 8748 1778 8764
rect 1744 8661 1778 8714
rect 0 8627 431 8661
rect 465 8627 1167 8661
rect 1201 8627 1840 8661
rect 431 8611 465 8627
rect 1167 8611 1201 8627
rect 4253 8501 4287 8517
rect 2612 8467 4253 8501
rect 2674 8376 2708 8467
rect 2674 8326 2708 8342
rect 2974 8376 3076 8392
rect 3008 8342 3076 8376
rect 2974 8326 3076 8342
rect 2691 8231 2725 8247
rect 2691 8181 2725 8197
rect 2824 8107 2858 8123
rect 2824 8057 2858 8073
rect 2957 7983 2991 7999
rect 2957 7933 2991 7949
rect 3042 7794 3076 8326
rect 3152 8250 3186 8467
rect 3356 8409 3390 8467
rect 4253 8451 4287 8467
rect 3356 8359 3390 8375
rect 3152 8200 3186 8216
rect 3252 8250 3286 8266
rect 3252 7810 3286 8216
rect 3154 7794 3188 7810
rect 3042 7760 3154 7794
rect 3042 7334 3076 7760
rect 3154 7744 3188 7760
rect 3252 7794 3303 7810
rect 3252 7760 3269 7794
rect 3252 7744 3303 7760
rect 2774 7300 3076 7334
rect 3152 7338 3186 7354
rect 2674 7250 2708 7266
rect 2674 7087 2708 7216
rect 2774 7250 2808 7300
rect 2774 7200 2808 7216
rect 2874 7250 2908 7266
rect 2874 7087 2908 7216
rect 2974 7250 3008 7300
rect 2974 7200 3008 7216
rect 3152 7087 3186 7304
rect 3252 7338 3286 7744
rect 3252 7288 3286 7304
rect 3356 7179 3390 7195
rect 3356 7087 3390 7145
rect 4253 7087 4287 7103
rect 2612 7053 4253 7087
rect 2674 6924 2708 7053
rect 2674 6874 2708 6890
rect 2774 6924 2808 6940
rect 2774 6824 2808 6890
rect 2874 6924 2908 7053
rect 2978 6995 3012 7053
rect 2978 6945 3012 6961
rect 2874 6874 2908 6890
rect 3142 6924 3176 7053
rect 3346 6995 3380 7053
rect 3346 6945 3380 6961
rect 3142 6874 3176 6890
rect 3242 6924 3276 6940
rect 2774 6790 3178 6824
rect 2824 6191 2858 6207
rect 2824 6141 2858 6157
rect 2724 5943 2758 5959
rect 2724 5893 2758 5909
rect 2942 5899 2976 6790
rect 3144 6342 3178 6790
rect 3144 6292 3178 6308
rect 3242 6361 3276 6890
rect 3510 6924 3544 7053
rect 3510 6874 3544 6890
rect 3610 6924 3644 6940
rect 3512 6361 3546 6377
rect 3242 6327 3512 6361
rect 3242 6308 3293 6327
rect 3512 6311 3546 6327
rect 3610 6361 3644 6890
rect 3768 6836 3802 7053
rect 3768 6786 3802 6802
rect 3868 6836 3902 6852
rect 3868 6380 3902 6802
rect 4026 6836 4060 7053
rect 4253 7037 4287 7053
rect 4026 6786 4060 6802
rect 4126 6836 4160 6852
rect 4126 6396 4160 6802
rect 4028 6380 4062 6396
rect 3610 6343 3661 6361
rect 3770 6343 3804 6359
rect 3610 6309 3770 6343
rect 2874 5865 2976 5899
rect 2674 5798 2708 5814
rect 2674 5673 2708 5764
rect 2874 5798 2908 5865
rect 2874 5748 2908 5764
rect 2978 5782 3012 5798
rect 2978 5673 3012 5748
rect 3142 5760 3176 5776
rect 3142 5673 3176 5726
rect 3242 5760 3276 6308
rect 3510 5798 3544 5814
rect 3242 5710 3276 5726
rect 3346 5765 3380 5781
rect 3346 5673 3380 5731
rect 3510 5673 3544 5764
rect 3610 5798 3644 6309
rect 3770 6293 3804 6309
rect 3868 6346 4028 6380
rect 3868 6309 3919 6346
rect 4028 6330 4062 6346
rect 4126 6380 4177 6396
rect 4126 6346 4143 6380
rect 4126 6330 4177 6346
rect 3610 5748 3644 5764
rect 3768 5850 3802 5866
rect 3768 5673 3802 5816
rect 3868 5850 3902 6309
rect 3868 5800 3902 5816
rect 4026 5924 4060 5940
rect 4026 5673 4060 5890
rect 4126 5924 4160 6330
rect 4126 5874 4160 5890
rect 4253 5673 4287 5689
rect 2612 5639 4253 5673
rect 2674 5586 2708 5639
rect 2674 5536 2708 5552
rect 2774 5586 2808 5602
rect 2676 5004 2710 5020
rect 2676 4954 2710 4970
rect 2774 5004 2808 5552
rect 2878 5564 2912 5639
rect 2878 5514 2912 5530
rect 3042 5510 3076 5639
rect 3300 5548 3334 5639
rect 3042 5460 3076 5476
rect 3142 5510 3176 5526
rect 3300 5498 3334 5514
rect 3400 5548 3434 5564
rect 3044 5004 3078 5020
rect 2774 4970 3044 5004
rect 2674 4422 2708 4438
rect 2674 4259 2708 4388
rect 2774 4422 2808 4970
rect 3044 4954 3078 4970
rect 3142 5004 3176 5476
rect 3142 4985 3193 5004
rect 3302 4985 3336 5001
rect 3142 4951 3302 4985
rect 2774 4372 2808 4388
rect 3042 4422 3076 4438
rect 2878 4351 2912 4367
rect 2878 4259 2912 4317
rect 3042 4259 3076 4388
rect 3142 4422 3176 4951
rect 3302 4935 3336 4951
rect 3400 4985 3434 5514
rect 3558 5422 3592 5639
rect 3816 5454 3850 5639
rect 3558 5372 3592 5388
rect 3658 5422 3692 5438
rect 3816 5404 3850 5420
rect 3916 5454 3950 5470
rect 3400 4966 3451 4985
rect 3658 4982 3692 5388
rect 3818 4982 3852 4998
rect 3560 4966 3594 4982
rect 3400 4932 3560 4966
rect 3142 4370 3176 4388
rect 3300 4422 3334 4438
rect 3300 4259 3334 4388
rect 3400 4422 3434 4932
rect 3560 4916 3594 4932
rect 3658 4948 3818 4982
rect 3658 4932 3709 4948
rect 3818 4932 3852 4948
rect 3916 4982 3950 5420
rect 4074 5422 4108 5639
rect 4253 5623 4287 5639
rect 4074 5372 4108 5388
rect 4174 5422 4208 5438
rect 4174 4982 4208 5388
rect 3916 4966 3967 4982
rect 4076 4966 4110 4982
rect 3916 4932 4076 4966
rect 3400 4372 3434 4388
rect 3558 4510 3592 4526
rect 3558 4259 3592 4476
rect 3658 4510 3692 4932
rect 3658 4460 3692 4476
rect 3816 4510 3850 4526
rect 3816 4259 3850 4476
rect 3916 4510 3950 4932
rect 4076 4916 4110 4932
rect 4174 4966 4225 4982
rect 4174 4932 4191 4966
rect 4174 4916 4225 4932
rect 3916 4460 3950 4476
rect 4074 4510 4108 4526
rect 4074 4259 4108 4476
rect 4174 4510 4208 4916
rect 4174 4460 4208 4476
rect 4253 4259 4287 4275
rect 2612 4225 4253 4259
rect 2674 4096 2708 4225
rect 2674 4046 2708 4062
rect 2774 4096 2808 4112
rect 2774 3996 2808 4062
rect 2874 4096 2908 4225
rect 2874 4046 2908 4062
rect 3052 4008 3086 4225
rect 3256 4167 3290 4225
rect 4253 4209 4287 4225
rect 3256 4117 3290 4133
rect 2774 3962 2976 3996
rect 2942 3536 2976 3962
rect 3052 3958 3086 3974
rect 3152 4008 3186 4024
rect 3152 3552 3186 3974
rect 3054 3536 3088 3552
rect 2942 3502 3054 3536
rect 2824 3363 2858 3379
rect 2824 3313 2858 3329
rect 2724 3115 2758 3131
rect 2724 3065 2758 3081
rect 2942 3071 2976 3502
rect 3054 3486 3088 3502
rect 3152 3536 3203 3552
rect 3152 3502 3169 3536
rect 3152 3486 3203 3502
rect 2874 3037 2976 3071
rect 3052 3064 3086 3080
rect 2674 2970 2708 2986
rect 2674 2845 2708 2936
rect 2874 2970 2908 3037
rect 2874 2920 2908 2936
rect 3052 2845 3086 3030
rect 3152 3064 3186 3486
rect 3152 3014 3186 3030
rect 3256 2937 3290 2953
rect 3256 2845 3290 2903
rect 4253 2845 4287 2861
rect 2612 2811 4253 2845
rect 2674 2758 2708 2811
rect 2674 2708 2708 2724
rect 2774 2758 2808 2774
rect 2676 2176 2710 2192
rect 2676 2126 2710 2142
rect 2774 2176 2808 2724
rect 2878 2753 2912 2811
rect 2878 2703 2912 2719
rect 3042 2720 3076 2811
rect 3042 2670 3076 2686
rect 3242 2720 3276 2736
rect 3242 2619 3276 2686
rect 3420 2626 3454 2811
rect 3624 2753 3658 2811
rect 4253 2795 4287 2811
rect 3624 2703 3658 2719
rect 3092 2575 3126 2591
rect 3242 2585 3344 2619
rect 2941 2541 3092 2575
rect 2941 2176 2975 2541
rect 3092 2525 3126 2541
rect 3192 2327 3226 2343
rect 3192 2277 3226 2293
rect 2774 2142 2975 2176
rect 3310 2154 3344 2585
rect 3420 2576 3454 2592
rect 3520 2626 3554 2642
rect 3520 2170 3554 2592
rect 3422 2154 3456 2170
rect 2674 1594 2708 1610
rect -17 1432 17 1447
rect -17 1431 1940 1432
rect 2674 1431 2708 1560
rect 2774 1594 2808 2142
rect 3310 2120 3422 2154
rect 3310 1694 3344 2120
rect 3422 2104 3456 2120
rect 3520 2154 3571 2170
rect 3520 2120 3537 2154
rect 3520 2104 3571 2120
rect 3142 1660 3344 1694
rect 3420 1682 3454 1698
rect 2774 1544 2808 1560
rect 3042 1594 3076 1610
rect 2878 1523 2912 1539
rect 2878 1431 2912 1489
rect 3042 1431 3076 1560
rect 3142 1594 3176 1660
rect 3142 1544 3176 1560
rect 3242 1594 3276 1610
rect 3242 1431 3276 1560
rect 3420 1431 3454 1648
rect 3520 1682 3554 2104
rect 3520 1632 3554 1648
rect 3624 1523 3658 1539
rect 3624 1431 3658 1489
rect 4253 1431 4287 1447
rect 17 1397 52 1431
rect 86 1397 188 1431
rect 222 1397 324 1431
rect 358 1397 460 1431
rect 494 1397 596 1431
rect 630 1397 732 1431
rect 766 1397 868 1431
rect 902 1397 1004 1431
rect 1038 1397 1940 1431
rect 2612 1397 4253 1431
rect -17 1396 1940 1397
rect -17 1381 17 1396
rect 36 1279 70 1312
rect 36 1211 70 1245
rect 36 1143 70 1177
rect 36 1075 70 1109
rect 36 1007 70 1041
rect 36 939 70 973
rect 36 871 70 905
rect 36 821 70 837
rect 122 1279 156 1396
rect 122 1211 156 1245
rect 122 1143 156 1177
rect 122 1075 156 1109
rect 122 1007 156 1041
rect 122 939 156 973
rect 122 871 156 905
rect 122 804 156 837
rect 280 1279 348 1312
rect 280 1245 297 1279
rect 331 1245 348 1279
rect 280 1211 348 1245
rect 280 1177 297 1211
rect 331 1177 348 1211
rect 280 1143 348 1177
rect 280 1109 297 1143
rect 331 1109 348 1143
rect 280 1075 348 1109
rect 280 1041 297 1075
rect 331 1041 348 1075
rect 280 1007 348 1041
rect 280 973 297 1007
rect 331 973 348 1007
rect 280 939 348 973
rect 280 905 297 939
rect 331 905 348 939
rect 280 871 348 905
rect 280 837 297 871
rect 331 837 348 871
rect 280 821 348 837
rect 280 804 297 821
rect 331 804 348 821
rect 472 1279 506 1396
rect 472 1211 506 1245
rect 472 1143 506 1177
rect 472 1075 506 1109
rect 472 1007 506 1041
rect 472 939 506 973
rect 472 871 506 905
rect 472 804 506 837
rect 630 1279 698 1312
rect 630 1245 647 1279
rect 681 1245 698 1279
rect 630 1211 698 1245
rect 630 1177 647 1211
rect 681 1177 698 1211
rect 630 1143 698 1177
rect 630 1109 647 1143
rect 681 1109 698 1143
rect 630 1075 698 1109
rect 630 1041 647 1075
rect 681 1041 698 1075
rect 630 1007 698 1041
rect 630 973 647 1007
rect 681 973 698 1007
rect 630 939 698 973
rect 630 905 647 939
rect 681 905 698 939
rect 630 871 698 905
rect 630 837 647 871
rect 681 837 698 871
rect 630 821 698 837
rect 630 804 647 821
rect 681 804 698 821
rect 822 1279 856 1396
rect 822 1211 856 1245
rect 822 1143 856 1177
rect 822 1075 856 1109
rect 822 1007 856 1041
rect 822 939 856 973
rect 822 871 856 905
rect 822 804 856 837
rect 908 1279 942 1312
rect 908 1211 942 1245
rect 908 1143 942 1177
rect 908 1075 942 1109
rect 908 1007 942 1041
rect 908 939 942 973
rect 908 871 942 905
rect 908 821 942 837
rect 1012 1279 1046 1396
rect 1012 1211 1046 1245
rect 1012 1143 1046 1177
rect 1012 1075 1046 1109
rect 1012 1007 1046 1041
rect 1012 939 1046 973
rect 1012 871 1046 905
rect 1012 804 1046 837
rect 1098 1279 1132 1312
rect 1098 1211 1132 1245
rect 1266 1268 1300 1396
rect 1470 1339 1504 1396
rect 1470 1289 1504 1305
rect 1266 1218 1300 1234
rect 1366 1268 1400 1284
rect 1098 1143 1132 1177
rect 1098 1075 1132 1109
rect 1098 1007 1132 1041
rect 1098 939 1132 973
rect 1098 871 1132 905
rect 1098 821 1132 837
rect 41 707 379 741
rect 413 707 1132 741
rect 41 627 57 661
rect 91 627 113 661
rect 249 656 283 707
rect 456 623 472 657
rect 506 623 522 657
rect 249 606 283 622
rect 137 547 153 581
rect 187 547 203 581
rect 472 566 506 623
rect 239 532 506 566
rect 239 501 273 532
rect 70 467 273 501
rect 472 421 506 532
rect 599 421 633 707
rect 695 656 729 707
rect 894 661 928 707
rect 1268 705 1302 721
rect 878 627 894 661
rect 928 627 944 661
rect 1268 655 1302 671
rect 1366 705 1400 1234
rect 1634 1215 1668 1396
rect 1838 1339 1872 1396
rect 1838 1289 1872 1305
rect 2674 1268 2708 1397
rect 2878 1339 2912 1397
rect 2878 1289 2912 1305
rect 1634 1165 1668 1181
rect 1734 1215 1768 1231
rect 2674 1218 2708 1234
rect 2774 1268 2808 1284
rect 1510 909 1544 925
rect 1509 875 1510 892
rect 1509 859 1544 875
rect 1509 726 1543 859
rect 1636 726 1670 742
rect 1509 705 1636 726
rect 1366 692 1636 705
rect 1366 671 1543 692
rect 1636 676 1670 692
rect 1734 726 1768 1181
rect 1734 692 1887 726
rect 695 606 729 622
rect 1098 581 1132 618
rect 775 547 791 581
rect 825 547 1132 581
rect 679 467 695 501
rect 729 467 908 501
rect 1012 467 1020 501
rect 1077 467 1093 501
rect 328 387 345 421
rect 456 387 472 421
rect 506 387 522 421
rect 583 387 599 421
rect 633 387 649 421
rect 1012 341 1046 467
rect 647 307 1046 341
rect 647 270 681 307
rect 36 261 70 270
rect 36 169 70 203
rect 36 102 70 135
rect 122 237 156 270
rect 122 169 156 203
rect -17 20 17 31
rect 122 20 156 135
rect 280 261 348 270
rect 280 203 297 261
rect 331 203 348 261
rect 280 169 348 203
rect 280 135 297 169
rect 331 135 348 169
rect 280 102 348 135
rect 472 237 506 270
rect 472 169 506 203
rect 472 20 506 135
rect 630 261 698 270
rect 630 203 647 261
rect 681 203 698 261
rect 630 169 698 203
rect 630 135 647 169
rect 681 135 698 169
rect 630 102 698 135
rect 822 237 856 270
rect 822 169 856 203
rect 822 20 856 135
rect 908 261 942 271
rect 908 169 942 203
rect 908 102 942 135
rect 1012 237 1046 270
rect 1012 169 1046 203
rect 1012 20 1046 135
rect 1098 261 1132 271
rect 1098 169 1132 203
rect 1098 102 1132 135
rect 1266 142 1300 158
rect -17 17 1168 20
rect 1266 17 1300 108
rect 1366 142 1400 671
rect 1634 236 1668 252
rect 1366 92 1400 108
rect 1470 109 1504 125
rect 1470 17 1504 75
rect 1634 17 1668 202
rect 1734 236 1768 692
rect 1853 522 1887 692
rect 2676 686 2710 702
rect 2676 636 2710 652
rect 2774 686 2808 1234
rect 3042 1268 3076 1397
rect 3042 1218 3076 1234
rect 3142 1268 3176 1284
rect 3142 704 3176 1234
rect 3300 1215 3334 1397
rect 3300 1165 3334 1181
rect 3400 1215 3434 1231
rect 3302 704 3336 720
rect 3044 686 3078 702
rect 2774 652 3044 686
rect 1853 472 1887 488
rect 1734 186 1768 202
rect 1838 109 1872 125
rect 1838 17 1872 75
rect 2674 104 2708 120
rect 2674 17 2708 70
rect 2774 104 2808 652
rect 3044 636 3078 652
rect 3142 670 3302 704
rect 3142 652 3193 670
rect 3302 654 3336 670
rect 3400 708 3434 1181
rect 3558 1180 3592 1397
rect 3558 1130 3592 1146
rect 3658 1180 3692 1196
rect 3658 724 3692 1146
rect 3816 1180 3850 1397
rect 3816 1130 3850 1146
rect 3916 1180 3950 1196
rect 3818 724 3852 740
rect 3560 708 3594 724
rect 3400 674 3560 708
rect 3400 670 3451 674
rect 2774 54 2808 70
rect 2878 109 2912 125
rect 2878 17 2912 75
rect 3042 104 3076 120
rect 3042 17 3076 70
rect 3142 104 3176 652
rect 3142 54 3176 70
rect 3300 194 3334 210
rect 3300 17 3334 160
rect 3400 194 3434 670
rect 3560 658 3594 674
rect 3658 690 3818 724
rect 3658 674 3709 690
rect 3818 674 3852 690
rect 3916 724 3950 1146
rect 4074 1180 4108 1397
rect 4253 1381 4287 1397
rect 4074 1130 4108 1146
rect 4174 1180 4208 1196
rect 4174 740 4208 1146
rect 4076 724 4110 740
rect 3916 690 4076 724
rect 3400 144 3434 160
rect 3558 236 3592 252
rect 3558 17 3592 202
rect 3658 236 3692 674
rect 3658 186 3692 202
rect 3816 268 3850 284
rect 3816 17 3850 234
rect 3916 268 3950 690
rect 4076 674 4110 690
rect 4174 724 4225 740
rect 4174 690 4191 724
rect 4174 674 4225 690
rect 3916 218 3950 234
rect 4074 268 4108 284
rect 4074 17 4108 234
rect 4174 268 4208 674
rect 4174 218 4208 234
rect 4253 17 4287 33
rect -17 15 52 17
rect 17 -17 52 15
rect 86 -17 188 17
rect 222 -17 324 17
rect 358 -17 460 17
rect 494 -17 596 17
rect 630 -17 732 17
rect 766 -17 868 17
rect 902 -17 1004 17
rect 1038 16 1168 17
rect 1204 16 1940 17
rect 1038 -17 1940 16
rect 2612 -17 4253 17
rect 17 -19 1940 -17
rect -17 -20 1940 -19
rect -17 -35 17 -20
rect 4253 -33 4287 -17
<< viali >>
rect 431 18707 465 18741
rect 1167 18707 1201 18741
rect 270 18109 304 18143
rect 638 18109 672 18143
rect 1006 18109 1040 18143
rect 1374 18109 1408 18143
rect 1627 18109 1661 18143
rect 1742 18109 1776 18143
rect 431 17587 465 17621
rect 1167 17587 1201 17621
rect 270 17065 304 17099
rect 638 17065 672 17099
rect 1006 17065 1040 17099
rect 1374 17065 1408 17099
rect 1627 17065 1661 17099
rect 1742 17065 1776 17099
rect 431 16467 465 16501
rect 1167 16467 1201 16501
rect 270 15869 304 15903
rect 638 15869 672 15903
rect 1006 15869 1040 15903
rect 1374 15869 1408 15903
rect 1627 15869 1661 15903
rect 1742 15869 1776 15903
rect 431 15347 465 15381
rect 1167 15347 1201 15381
rect 270 14825 304 14859
rect 638 14825 672 14859
rect 1006 14825 1040 14859
rect 1374 14825 1408 14859
rect 1627 14825 1661 14859
rect 1742 14825 1776 14859
rect 431 14227 465 14261
rect 1167 14227 1201 14261
rect 270 13629 304 13663
rect 638 13629 672 13663
rect 1006 13629 1040 13663
rect 1374 13629 1408 13663
rect 1627 13629 1661 13663
rect 1742 13629 1776 13663
rect 431 13107 465 13141
rect 1167 13107 1201 13141
rect 270 12585 304 12619
rect 638 12585 672 12619
rect 1006 12585 1040 12619
rect 1374 12585 1408 12619
rect 1627 12585 1661 12619
rect 1742 12585 1776 12619
rect 431 11987 465 12021
rect 1167 11987 1201 12021
rect 270 11389 304 11423
rect 638 11389 672 11423
rect 1006 11389 1040 11423
rect 1374 11389 1408 11423
rect 1627 11389 1661 11423
rect 1742 11389 1776 11423
rect 431 10867 465 10901
rect 1167 10867 1201 10901
rect 270 10345 304 10379
rect 638 10345 672 10379
rect 1006 10345 1040 10379
rect 1374 10345 1408 10379
rect 1627 10345 1661 10379
rect 1742 10345 1776 10379
rect 431 9747 465 9781
rect 1167 9747 1201 9781
rect 270 9149 304 9183
rect 638 9149 672 9183
rect 1006 9149 1040 9183
rect 1374 9149 1408 9183
rect 1627 9149 1661 9183
rect 1742 9149 1776 9183
rect 431 8627 465 8661
rect 1167 8627 1201 8661
rect 4253 8467 4287 8501
rect 2691 8197 2725 8231
rect 2824 8073 2858 8107
rect 2957 7949 2991 7983
rect 3269 7760 3303 7794
rect 4253 7053 4287 7087
rect 2824 6157 2858 6191
rect 2724 5909 2758 5943
rect 4143 6346 4177 6380
rect 4253 5639 4287 5673
rect 2676 4970 2710 5004
rect 4191 4932 4225 4966
rect 4253 4225 4287 4259
rect 2824 3329 2858 3363
rect 2724 3081 2758 3115
rect 3169 3502 3203 3536
rect 4253 2811 4287 2845
rect 2676 2142 2710 2176
rect 3192 2293 3226 2327
rect 3537 2120 3571 2154
rect -17 1397 17 1431
rect 4253 1397 4287 1431
rect 36 787 70 821
rect 297 787 331 821
rect 647 787 681 821
rect 908 787 942 821
rect 1098 787 1132 821
rect 379 707 413 741
rect 113 627 147 661
rect 153 547 187 581
rect 36 467 70 501
rect 1268 671 1302 705
rect 1510 875 1544 909
rect 1098 618 1132 652
rect 908 467 942 501
rect 1020 467 1043 501
rect 1043 467 1054 501
rect 379 387 413 421
rect 36 237 70 261
rect 36 227 70 237
rect 297 237 331 261
rect 297 227 331 237
rect 647 237 681 261
rect 647 227 681 237
rect 908 237 942 261
rect 908 227 942 237
rect 1098 237 1132 261
rect 1098 227 1132 237
rect 2676 652 2710 686
rect 1853 488 1887 522
rect 4191 690 4225 724
rect -17 -19 17 15
rect 4253 -17 4287 17
<< metal1 >>
rect 416 18698 422 18750
rect 474 18698 480 18750
rect 1152 18698 1158 18750
rect 1210 18698 1216 18750
rect 255 18100 261 18152
rect 313 18100 319 18152
rect 623 18100 629 18152
rect 681 18100 687 18152
rect 991 18100 997 18152
rect 1049 18100 1055 18152
rect 1359 18100 1365 18152
rect 1417 18100 1423 18152
rect 1612 18100 1618 18152
rect 1670 18100 1676 18152
rect 1727 18100 1733 18152
rect 1785 18100 1791 18152
rect 416 17578 422 17630
rect 474 17578 480 17630
rect 1152 17578 1158 17630
rect 1210 17578 1216 17630
rect 255 17056 261 17108
rect 313 17056 319 17108
rect 623 17056 629 17108
rect 681 17056 687 17108
rect 991 17056 997 17108
rect 1049 17056 1055 17108
rect 1359 17056 1365 17108
rect 1417 17056 1423 17108
rect 1612 17056 1618 17108
rect 1670 17056 1676 17108
rect 1727 17056 1733 17108
rect 1785 17056 1791 17108
rect 416 16458 422 16510
rect 474 16458 480 16510
rect 1152 16458 1158 16510
rect 1210 16458 1216 16510
rect 255 15860 261 15912
rect 313 15860 319 15912
rect 623 15860 629 15912
rect 681 15860 687 15912
rect 991 15860 997 15912
rect 1049 15860 1055 15912
rect 1359 15860 1365 15912
rect 1417 15860 1423 15912
rect 1612 15860 1618 15912
rect 1670 15860 1676 15912
rect 1727 15860 1733 15912
rect 1785 15860 1791 15912
rect 416 15338 422 15390
rect 474 15338 480 15390
rect 1152 15338 1158 15390
rect 1210 15338 1216 15390
rect 255 14816 261 14868
rect 313 14816 319 14868
rect 623 14816 629 14868
rect 681 14816 687 14868
rect 991 14816 997 14868
rect 1049 14816 1055 14868
rect 1359 14816 1365 14868
rect 1417 14816 1423 14868
rect 1612 14816 1618 14868
rect 1670 14816 1676 14868
rect 1727 14816 1733 14868
rect 1785 14816 1791 14868
rect 416 14218 422 14270
rect 474 14218 480 14270
rect 1152 14218 1158 14270
rect 1210 14218 1216 14270
rect 255 13620 261 13672
rect 313 13620 319 13672
rect 623 13620 629 13672
rect 681 13620 687 13672
rect 991 13620 997 13672
rect 1049 13620 1055 13672
rect 1359 13620 1365 13672
rect 1417 13620 1423 13672
rect 1612 13620 1618 13672
rect 1670 13620 1676 13672
rect 1727 13620 1733 13672
rect 1785 13620 1791 13672
rect 416 13098 422 13150
rect 474 13098 480 13150
rect 1152 13098 1158 13150
rect 1210 13098 1216 13150
rect 255 12576 261 12628
rect 313 12576 319 12628
rect 623 12576 629 12628
rect 681 12576 687 12628
rect 991 12576 997 12628
rect 1049 12576 1055 12628
rect 1359 12576 1365 12628
rect 1417 12576 1423 12628
rect 1612 12576 1618 12628
rect 1670 12576 1676 12628
rect 1727 12576 1733 12628
rect 1785 12576 1791 12628
rect 416 11978 422 12030
rect 474 11978 480 12030
rect 1152 11978 1158 12030
rect 1210 11978 1216 12030
rect 255 11380 261 11432
rect 313 11380 319 11432
rect 623 11380 629 11432
rect 681 11380 687 11432
rect 991 11380 997 11432
rect 1049 11380 1055 11432
rect 1359 11380 1365 11432
rect 1417 11380 1423 11432
rect 1612 11380 1618 11432
rect 1670 11380 1676 11432
rect 1727 11380 1733 11432
rect 1785 11380 1791 11432
rect 416 10858 422 10910
rect 474 10858 480 10910
rect 1152 10858 1158 10910
rect 1210 10858 1216 10910
rect 255 10336 261 10388
rect 313 10336 319 10388
rect 623 10336 629 10388
rect 681 10336 687 10388
rect 991 10336 997 10388
rect 1049 10336 1055 10388
rect 1359 10336 1365 10388
rect 1417 10336 1423 10388
rect 1612 10336 1618 10388
rect 1670 10336 1676 10388
rect 1727 10336 1733 10388
rect 1785 10336 1791 10388
rect 416 9738 422 9790
rect 474 9738 480 9790
rect 1152 9738 1158 9790
rect 1210 9738 1216 9790
rect 255 9140 261 9192
rect 313 9140 319 9192
rect 623 9140 629 9192
rect 681 9140 687 9192
rect 991 9140 997 9192
rect 1049 9140 1055 9192
rect 1359 9140 1365 9192
rect 1417 9140 1423 9192
rect 1612 9140 1618 9192
rect 1670 9140 1676 9192
rect 1727 9140 1733 9192
rect 1785 9140 1791 9192
rect 416 8618 422 8670
rect 474 8618 480 8670
rect 1152 8618 1158 8670
rect 1210 8618 1216 8670
rect 4238 8458 4244 8510
rect 4296 8458 4302 8510
rect 2006 8188 2012 8240
rect 2064 8228 2070 8240
rect 2679 8231 2737 8237
rect 2679 8228 2691 8231
rect 2064 8200 2691 8228
rect 2064 8188 2070 8200
rect 2679 8197 2691 8200
rect 2725 8197 2737 8231
rect 2679 8191 2737 8197
rect 2090 8064 2096 8116
rect 2148 8104 2154 8116
rect 2812 8107 2870 8113
rect 2812 8104 2824 8107
rect 2148 8076 2824 8104
rect 2148 8064 2154 8076
rect 2812 8073 2824 8076
rect 2858 8073 2870 8107
rect 2812 8067 2870 8073
rect 2426 7940 2432 7992
rect 2484 7980 2490 7992
rect 2945 7983 3003 7989
rect 2945 7980 2957 7983
rect 2484 7952 2957 7980
rect 2484 7940 2490 7952
rect 2945 7949 2957 7952
rect 2991 7949 3003 7983
rect 2945 7943 3003 7949
rect 3254 7751 3260 7803
rect 3312 7751 3318 7803
rect 171 7027 177 7079
rect 229 7067 235 7079
rect 2006 7067 2012 7079
rect 229 7039 2012 7067
rect 229 7027 235 7039
rect 2006 7027 2012 7039
rect 2064 7027 2070 7079
rect 4238 7044 4244 7096
rect 4296 7044 4302 7096
rect 4128 6337 4134 6389
rect 4186 6337 4192 6389
rect 2006 6148 2012 6200
rect 2064 6188 2070 6200
rect 2812 6191 2870 6197
rect 2812 6188 2824 6191
rect 2064 6160 2824 6188
rect 2064 6148 2070 6160
rect 2812 6157 2824 6160
rect 2858 6157 2870 6191
rect 2812 6151 2870 6157
rect 2174 5900 2180 5952
rect 2232 5940 2238 5952
rect 2712 5943 2770 5949
rect 2712 5940 2724 5943
rect 2232 5912 2724 5940
rect 2232 5900 2238 5912
rect 2712 5909 2724 5912
rect 2758 5909 2770 5943
rect 2712 5903 2770 5909
rect 4238 5630 4244 5682
rect 4296 5630 4302 5682
rect 2090 4961 2096 5013
rect 2148 5001 2154 5013
rect 2664 5004 2722 5010
rect 2664 5001 2676 5004
rect 2148 4973 2676 5001
rect 2148 4961 2154 4973
rect 2664 4970 2676 4973
rect 2710 4970 2722 5004
rect 2664 4964 2722 4970
rect 4176 4923 4182 4975
rect 4234 4923 4240 4975
rect 4238 4216 4244 4268
rect 4296 4216 4302 4268
rect 3154 3493 3160 3545
rect 3212 3493 3218 3545
rect 2426 3320 2432 3372
rect 2484 3360 2490 3372
rect 2812 3363 2870 3369
rect 2812 3360 2824 3363
rect 2484 3332 2824 3360
rect 2484 3320 2490 3332
rect 2812 3329 2824 3332
rect 2858 3329 2870 3363
rect 2812 3323 2870 3329
rect 2258 3072 2264 3124
rect 2316 3112 2322 3124
rect 2712 3115 2770 3121
rect 2712 3112 2724 3115
rect 2316 3084 2724 3112
rect 2316 3072 2322 3084
rect 2712 3081 2724 3084
rect 2758 3081 2770 3115
rect 2712 3075 2770 3081
rect 351 2802 357 2854
rect 409 2842 415 2854
rect 2258 2842 2264 2854
rect 409 2814 2264 2842
rect 409 2802 415 2814
rect 2258 2802 2264 2814
rect 2316 2802 2322 2854
rect 4238 2802 4244 2854
rect 4296 2802 4302 2854
rect 3177 2284 3183 2336
rect 3235 2284 3241 2336
rect 2258 2133 2264 2185
rect 2316 2173 2322 2185
rect 2664 2176 2722 2182
rect 2664 2173 2676 2176
rect 2316 2145 2676 2173
rect 2316 2133 2322 2145
rect 2664 2142 2676 2145
rect 2710 2142 2722 2176
rect 2664 2136 2722 2142
rect 3522 2111 3528 2163
rect 3580 2111 3586 2163
rect -32 1388 -26 1440
rect 26 1388 32 1440
rect 4238 1388 4244 1440
rect 4296 1388 4302 1440
rect 1494 866 1500 918
rect 1552 866 1559 918
rect 24 821 82 827
rect 24 787 36 821
rect 70 787 82 821
rect 24 781 82 787
rect 285 821 343 827
rect 285 787 297 821
rect 331 787 343 821
rect 285 781 343 787
rect 635 821 693 827
rect 635 787 647 821
rect 681 787 693 821
rect 635 781 693 787
rect 896 821 954 827
rect 896 787 908 821
rect 942 787 954 821
rect 896 781 954 787
rect 1086 821 1144 827
rect 1086 787 1098 821
rect 1132 787 1144 821
rect 1086 781 1144 787
rect 36 507 70 781
rect 101 661 159 667
rect 297 661 331 781
rect 369 750 423 756
rect 369 747 370 750
rect 367 701 370 747
rect 422 747 423 750
rect 369 698 370 701
rect 422 701 425 747
rect 422 698 423 701
rect 369 692 423 698
rect 101 627 113 661
rect 147 627 331 661
rect 101 621 159 627
rect 137 538 144 590
rect 196 538 203 590
rect 24 501 82 507
rect 24 467 36 501
rect 70 467 82 501
rect 24 461 82 467
rect 36 267 70 461
rect 297 267 331 627
rect 379 436 413 692
rect 369 427 423 436
rect 367 421 425 427
rect 367 387 379 421
rect 413 387 425 421
rect 367 381 425 387
rect 369 372 423 381
rect 647 267 681 781
rect 908 507 942 781
rect 1098 661 1132 781
rect 1253 662 1259 714
rect 1311 662 1317 714
rect 1082 609 1089 661
rect 1141 609 1148 661
rect 2661 643 2667 695
rect 2719 643 2725 695
rect 4176 681 4182 733
rect 4234 681 4240 733
rect 896 501 954 507
rect 896 467 908 501
rect 942 467 954 501
rect 896 461 954 467
rect 908 267 942 461
rect 1004 458 1011 510
rect 1063 458 1070 510
rect 1098 267 1132 609
rect 1838 479 1844 531
rect 1896 479 1902 531
rect 24 261 82 267
rect 24 227 36 261
rect 70 227 82 261
rect 24 221 82 227
rect 285 261 343 267
rect 285 227 297 261
rect 331 227 343 261
rect 285 221 343 227
rect 635 261 693 267
rect 635 227 647 261
rect 681 227 693 261
rect 635 221 693 227
rect 896 261 954 267
rect 896 227 908 261
rect 942 227 954 261
rect 896 221 954 227
rect 1086 261 1144 267
rect 1086 227 1098 261
rect 1132 227 1144 261
rect 1086 221 1144 227
rect -32 -28 -26 24
rect 26 -28 32 24
rect 4238 -26 4244 26
rect 4296 -26 4302 26
<< via1 >>
rect 422 18741 474 18750
rect 422 18707 431 18741
rect 431 18707 465 18741
rect 465 18707 474 18741
rect 422 18698 474 18707
rect 1158 18741 1210 18750
rect 1158 18707 1167 18741
rect 1167 18707 1201 18741
rect 1201 18707 1210 18741
rect 1158 18698 1210 18707
rect 261 18143 313 18152
rect 261 18109 270 18143
rect 270 18109 304 18143
rect 304 18109 313 18143
rect 261 18100 313 18109
rect 629 18143 681 18152
rect 629 18109 638 18143
rect 638 18109 672 18143
rect 672 18109 681 18143
rect 629 18100 681 18109
rect 997 18143 1049 18152
rect 997 18109 1006 18143
rect 1006 18109 1040 18143
rect 1040 18109 1049 18143
rect 997 18100 1049 18109
rect 1365 18143 1417 18152
rect 1365 18109 1374 18143
rect 1374 18109 1408 18143
rect 1408 18109 1417 18143
rect 1365 18100 1417 18109
rect 1618 18143 1670 18152
rect 1618 18109 1627 18143
rect 1627 18109 1661 18143
rect 1661 18109 1670 18143
rect 1618 18100 1670 18109
rect 1733 18143 1785 18152
rect 1733 18109 1742 18143
rect 1742 18109 1776 18143
rect 1776 18109 1785 18143
rect 1733 18100 1785 18109
rect 422 17621 474 17630
rect 422 17587 431 17621
rect 431 17587 465 17621
rect 465 17587 474 17621
rect 422 17578 474 17587
rect 1158 17621 1210 17630
rect 1158 17587 1167 17621
rect 1167 17587 1201 17621
rect 1201 17587 1210 17621
rect 1158 17578 1210 17587
rect 261 17099 313 17108
rect 261 17065 270 17099
rect 270 17065 304 17099
rect 304 17065 313 17099
rect 261 17056 313 17065
rect 629 17099 681 17108
rect 629 17065 638 17099
rect 638 17065 672 17099
rect 672 17065 681 17099
rect 629 17056 681 17065
rect 997 17099 1049 17108
rect 997 17065 1006 17099
rect 1006 17065 1040 17099
rect 1040 17065 1049 17099
rect 997 17056 1049 17065
rect 1365 17099 1417 17108
rect 1365 17065 1374 17099
rect 1374 17065 1408 17099
rect 1408 17065 1417 17099
rect 1365 17056 1417 17065
rect 1618 17099 1670 17108
rect 1618 17065 1627 17099
rect 1627 17065 1661 17099
rect 1661 17065 1670 17099
rect 1618 17056 1670 17065
rect 1733 17099 1785 17108
rect 1733 17065 1742 17099
rect 1742 17065 1776 17099
rect 1776 17065 1785 17099
rect 1733 17056 1785 17065
rect 422 16501 474 16510
rect 422 16467 431 16501
rect 431 16467 465 16501
rect 465 16467 474 16501
rect 422 16458 474 16467
rect 1158 16501 1210 16510
rect 1158 16467 1167 16501
rect 1167 16467 1201 16501
rect 1201 16467 1210 16501
rect 1158 16458 1210 16467
rect 261 15903 313 15912
rect 261 15869 270 15903
rect 270 15869 304 15903
rect 304 15869 313 15903
rect 261 15860 313 15869
rect 629 15903 681 15912
rect 629 15869 638 15903
rect 638 15869 672 15903
rect 672 15869 681 15903
rect 629 15860 681 15869
rect 997 15903 1049 15912
rect 997 15869 1006 15903
rect 1006 15869 1040 15903
rect 1040 15869 1049 15903
rect 997 15860 1049 15869
rect 1365 15903 1417 15912
rect 1365 15869 1374 15903
rect 1374 15869 1408 15903
rect 1408 15869 1417 15903
rect 1365 15860 1417 15869
rect 1618 15903 1670 15912
rect 1618 15869 1627 15903
rect 1627 15869 1661 15903
rect 1661 15869 1670 15903
rect 1618 15860 1670 15869
rect 1733 15903 1785 15912
rect 1733 15869 1742 15903
rect 1742 15869 1776 15903
rect 1776 15869 1785 15903
rect 1733 15860 1785 15869
rect 422 15381 474 15390
rect 422 15347 431 15381
rect 431 15347 465 15381
rect 465 15347 474 15381
rect 422 15338 474 15347
rect 1158 15381 1210 15390
rect 1158 15347 1167 15381
rect 1167 15347 1201 15381
rect 1201 15347 1210 15381
rect 1158 15338 1210 15347
rect 261 14859 313 14868
rect 261 14825 270 14859
rect 270 14825 304 14859
rect 304 14825 313 14859
rect 261 14816 313 14825
rect 629 14859 681 14868
rect 629 14825 638 14859
rect 638 14825 672 14859
rect 672 14825 681 14859
rect 629 14816 681 14825
rect 997 14859 1049 14868
rect 997 14825 1006 14859
rect 1006 14825 1040 14859
rect 1040 14825 1049 14859
rect 997 14816 1049 14825
rect 1365 14859 1417 14868
rect 1365 14825 1374 14859
rect 1374 14825 1408 14859
rect 1408 14825 1417 14859
rect 1365 14816 1417 14825
rect 1618 14859 1670 14868
rect 1618 14825 1627 14859
rect 1627 14825 1661 14859
rect 1661 14825 1670 14859
rect 1618 14816 1670 14825
rect 1733 14859 1785 14868
rect 1733 14825 1742 14859
rect 1742 14825 1776 14859
rect 1776 14825 1785 14859
rect 1733 14816 1785 14825
rect 422 14261 474 14270
rect 422 14227 431 14261
rect 431 14227 465 14261
rect 465 14227 474 14261
rect 422 14218 474 14227
rect 1158 14261 1210 14270
rect 1158 14227 1167 14261
rect 1167 14227 1201 14261
rect 1201 14227 1210 14261
rect 1158 14218 1210 14227
rect 261 13663 313 13672
rect 261 13629 270 13663
rect 270 13629 304 13663
rect 304 13629 313 13663
rect 261 13620 313 13629
rect 629 13663 681 13672
rect 629 13629 638 13663
rect 638 13629 672 13663
rect 672 13629 681 13663
rect 629 13620 681 13629
rect 997 13663 1049 13672
rect 997 13629 1006 13663
rect 1006 13629 1040 13663
rect 1040 13629 1049 13663
rect 997 13620 1049 13629
rect 1365 13663 1417 13672
rect 1365 13629 1374 13663
rect 1374 13629 1408 13663
rect 1408 13629 1417 13663
rect 1365 13620 1417 13629
rect 1618 13663 1670 13672
rect 1618 13629 1627 13663
rect 1627 13629 1661 13663
rect 1661 13629 1670 13663
rect 1618 13620 1670 13629
rect 1733 13663 1785 13672
rect 1733 13629 1742 13663
rect 1742 13629 1776 13663
rect 1776 13629 1785 13663
rect 1733 13620 1785 13629
rect 422 13141 474 13150
rect 422 13107 431 13141
rect 431 13107 465 13141
rect 465 13107 474 13141
rect 422 13098 474 13107
rect 1158 13141 1210 13150
rect 1158 13107 1167 13141
rect 1167 13107 1201 13141
rect 1201 13107 1210 13141
rect 1158 13098 1210 13107
rect 261 12619 313 12628
rect 261 12585 270 12619
rect 270 12585 304 12619
rect 304 12585 313 12619
rect 261 12576 313 12585
rect 629 12619 681 12628
rect 629 12585 638 12619
rect 638 12585 672 12619
rect 672 12585 681 12619
rect 629 12576 681 12585
rect 997 12619 1049 12628
rect 997 12585 1006 12619
rect 1006 12585 1040 12619
rect 1040 12585 1049 12619
rect 997 12576 1049 12585
rect 1365 12619 1417 12628
rect 1365 12585 1374 12619
rect 1374 12585 1408 12619
rect 1408 12585 1417 12619
rect 1365 12576 1417 12585
rect 1618 12619 1670 12628
rect 1618 12585 1627 12619
rect 1627 12585 1661 12619
rect 1661 12585 1670 12619
rect 1618 12576 1670 12585
rect 1733 12619 1785 12628
rect 1733 12585 1742 12619
rect 1742 12585 1776 12619
rect 1776 12585 1785 12619
rect 1733 12576 1785 12585
rect 422 12021 474 12030
rect 422 11987 431 12021
rect 431 11987 465 12021
rect 465 11987 474 12021
rect 422 11978 474 11987
rect 1158 12021 1210 12030
rect 1158 11987 1167 12021
rect 1167 11987 1201 12021
rect 1201 11987 1210 12021
rect 1158 11978 1210 11987
rect 261 11423 313 11432
rect 261 11389 270 11423
rect 270 11389 304 11423
rect 304 11389 313 11423
rect 261 11380 313 11389
rect 629 11423 681 11432
rect 629 11389 638 11423
rect 638 11389 672 11423
rect 672 11389 681 11423
rect 629 11380 681 11389
rect 997 11423 1049 11432
rect 997 11389 1006 11423
rect 1006 11389 1040 11423
rect 1040 11389 1049 11423
rect 997 11380 1049 11389
rect 1365 11423 1417 11432
rect 1365 11389 1374 11423
rect 1374 11389 1408 11423
rect 1408 11389 1417 11423
rect 1365 11380 1417 11389
rect 1618 11423 1670 11432
rect 1618 11389 1627 11423
rect 1627 11389 1661 11423
rect 1661 11389 1670 11423
rect 1618 11380 1670 11389
rect 1733 11423 1785 11432
rect 1733 11389 1742 11423
rect 1742 11389 1776 11423
rect 1776 11389 1785 11423
rect 1733 11380 1785 11389
rect 422 10901 474 10910
rect 422 10867 431 10901
rect 431 10867 465 10901
rect 465 10867 474 10901
rect 422 10858 474 10867
rect 1158 10901 1210 10910
rect 1158 10867 1167 10901
rect 1167 10867 1201 10901
rect 1201 10867 1210 10901
rect 1158 10858 1210 10867
rect 261 10379 313 10388
rect 261 10345 270 10379
rect 270 10345 304 10379
rect 304 10345 313 10379
rect 261 10336 313 10345
rect 629 10379 681 10388
rect 629 10345 638 10379
rect 638 10345 672 10379
rect 672 10345 681 10379
rect 629 10336 681 10345
rect 997 10379 1049 10388
rect 997 10345 1006 10379
rect 1006 10345 1040 10379
rect 1040 10345 1049 10379
rect 997 10336 1049 10345
rect 1365 10379 1417 10388
rect 1365 10345 1374 10379
rect 1374 10345 1408 10379
rect 1408 10345 1417 10379
rect 1365 10336 1417 10345
rect 1618 10379 1670 10388
rect 1618 10345 1627 10379
rect 1627 10345 1661 10379
rect 1661 10345 1670 10379
rect 1618 10336 1670 10345
rect 1733 10379 1785 10388
rect 1733 10345 1742 10379
rect 1742 10345 1776 10379
rect 1776 10345 1785 10379
rect 1733 10336 1785 10345
rect 422 9781 474 9790
rect 422 9747 431 9781
rect 431 9747 465 9781
rect 465 9747 474 9781
rect 422 9738 474 9747
rect 1158 9781 1210 9790
rect 1158 9747 1167 9781
rect 1167 9747 1201 9781
rect 1201 9747 1210 9781
rect 1158 9738 1210 9747
rect 261 9183 313 9192
rect 261 9149 270 9183
rect 270 9149 304 9183
rect 304 9149 313 9183
rect 261 9140 313 9149
rect 629 9183 681 9192
rect 629 9149 638 9183
rect 638 9149 672 9183
rect 672 9149 681 9183
rect 629 9140 681 9149
rect 997 9183 1049 9192
rect 997 9149 1006 9183
rect 1006 9149 1040 9183
rect 1040 9149 1049 9183
rect 997 9140 1049 9149
rect 1365 9183 1417 9192
rect 1365 9149 1374 9183
rect 1374 9149 1408 9183
rect 1408 9149 1417 9183
rect 1365 9140 1417 9149
rect 1618 9183 1670 9192
rect 1618 9149 1627 9183
rect 1627 9149 1661 9183
rect 1661 9149 1670 9183
rect 1618 9140 1670 9149
rect 1733 9183 1785 9192
rect 1733 9149 1742 9183
rect 1742 9149 1776 9183
rect 1776 9149 1785 9183
rect 1733 9140 1785 9149
rect 422 8661 474 8670
rect 422 8627 431 8661
rect 431 8627 465 8661
rect 465 8627 474 8661
rect 422 8618 474 8627
rect 1158 8661 1210 8670
rect 1158 8627 1167 8661
rect 1167 8627 1201 8661
rect 1201 8627 1210 8661
rect 1158 8618 1210 8627
rect 4244 8501 4296 8510
rect 4244 8467 4253 8501
rect 4253 8467 4287 8501
rect 4287 8467 4296 8501
rect 4244 8458 4296 8467
rect 2012 8188 2064 8240
rect 2096 8064 2148 8116
rect 2432 7940 2484 7992
rect 3260 7794 3312 7803
rect 3260 7760 3269 7794
rect 3269 7760 3303 7794
rect 3303 7760 3312 7794
rect 3260 7751 3312 7760
rect 177 7027 229 7079
rect 2012 7027 2064 7079
rect 4244 7087 4296 7096
rect 4244 7053 4253 7087
rect 4253 7053 4287 7087
rect 4287 7053 4296 7087
rect 4244 7044 4296 7053
rect 4134 6380 4186 6389
rect 4134 6346 4143 6380
rect 4143 6346 4177 6380
rect 4177 6346 4186 6380
rect 4134 6337 4186 6346
rect 2012 6148 2064 6200
rect 2180 5900 2232 5952
rect 4244 5673 4296 5682
rect 4244 5639 4253 5673
rect 4253 5639 4287 5673
rect 4287 5639 4296 5673
rect 4244 5630 4296 5639
rect 2096 4961 2148 5013
rect 4182 4966 4234 4975
rect 4182 4932 4191 4966
rect 4191 4932 4225 4966
rect 4225 4932 4234 4966
rect 4182 4923 4234 4932
rect 4244 4259 4296 4268
rect 4244 4225 4253 4259
rect 4253 4225 4287 4259
rect 4287 4225 4296 4259
rect 4244 4216 4296 4225
rect 3160 3536 3212 3545
rect 3160 3502 3169 3536
rect 3169 3502 3203 3536
rect 3203 3502 3212 3536
rect 3160 3493 3212 3502
rect 2432 3320 2484 3372
rect 2264 3072 2316 3124
rect 357 2802 409 2854
rect 2264 2802 2316 2854
rect 4244 2845 4296 2854
rect 4244 2811 4253 2845
rect 4253 2811 4287 2845
rect 4287 2811 4296 2845
rect 4244 2802 4296 2811
rect 3183 2327 3235 2336
rect 3183 2293 3192 2327
rect 3192 2293 3226 2327
rect 3226 2293 3235 2327
rect 3183 2284 3235 2293
rect 2264 2133 2316 2185
rect 3528 2154 3580 2163
rect 3528 2120 3537 2154
rect 3537 2120 3571 2154
rect 3571 2120 3580 2154
rect 3528 2111 3580 2120
rect -26 1431 26 1440
rect -26 1397 -17 1431
rect -17 1397 17 1431
rect 17 1397 26 1431
rect -26 1388 26 1397
rect 4244 1431 4296 1440
rect 4244 1397 4253 1431
rect 4253 1397 4287 1431
rect 4287 1397 4296 1431
rect 4244 1388 4296 1397
rect 1500 909 1552 918
rect 1500 875 1510 909
rect 1510 875 1544 909
rect 1544 875 1552 909
rect 1500 866 1552 875
rect 370 741 422 750
rect 370 707 379 741
rect 379 707 413 741
rect 413 707 422 741
rect 370 698 422 707
rect 144 581 196 590
rect 144 547 153 581
rect 153 547 187 581
rect 187 547 196 581
rect 144 538 196 547
rect 1259 705 1311 714
rect 1259 671 1268 705
rect 1268 671 1302 705
rect 1302 671 1311 705
rect 1259 662 1311 671
rect 1089 652 1141 661
rect 1089 618 1098 652
rect 1098 618 1132 652
rect 1132 618 1141 652
rect 1089 609 1141 618
rect 2667 686 2719 695
rect 2667 652 2676 686
rect 2676 652 2710 686
rect 2710 652 2719 686
rect 2667 643 2719 652
rect 4182 724 4234 733
rect 4182 690 4191 724
rect 4191 690 4225 724
rect 4225 690 4234 724
rect 4182 681 4234 690
rect 1011 501 1063 510
rect 1011 467 1020 501
rect 1020 467 1054 501
rect 1054 467 1063 501
rect 1011 458 1063 467
rect 1844 522 1896 531
rect 1844 488 1853 522
rect 1853 488 1887 522
rect 1887 488 1896 522
rect 1844 479 1896 488
rect -26 15 26 24
rect -26 -19 -17 15
rect -17 -19 17 15
rect 17 -19 26 15
rect -26 -28 26 -19
rect 4244 17 4296 26
rect 4244 -17 4253 17
rect 4253 -17 4287 17
rect 4287 -17 4296 17
rect 4244 -26 4296 -17
<< metal2 >>
rect 420 18752 476 18761
rect 420 18687 476 18696
rect 1156 18752 1212 18761
rect 1156 18687 1212 18696
rect 259 18154 315 18163
rect 189 18112 259 18140
rect 189 7085 217 18112
rect 259 18089 315 18098
rect 627 18154 683 18163
rect 627 18089 683 18098
rect 995 18154 1051 18163
rect 995 18089 1051 18098
rect 1363 18154 1419 18163
rect 1363 18089 1419 18098
rect 1616 18154 1672 18163
rect 1616 18089 1672 18098
rect 1733 18152 1785 18158
rect 1733 18094 1785 18100
rect 420 17632 476 17641
rect 420 17567 476 17576
rect 1156 17632 1212 17641
rect 1745 17618 1773 18094
rect 1156 17567 1212 17576
rect 1630 17590 1773 17618
rect 1630 17119 1658 17590
rect 259 17110 315 17119
rect 259 17045 315 17054
rect 627 17110 683 17119
rect 627 17045 683 17054
rect 995 17110 1051 17119
rect 995 17045 1051 17054
rect 1363 17110 1419 17119
rect 1363 17045 1419 17054
rect 1616 17110 1672 17119
rect 1616 17045 1672 17054
rect 1733 17108 1785 17114
rect 1733 17050 1785 17056
rect 420 16512 476 16521
rect 420 16447 476 16456
rect 1156 16512 1212 16521
rect 1745 16498 1773 17050
rect 1156 16447 1212 16456
rect 1630 16470 1773 16498
rect 1630 15923 1658 16470
rect 259 15914 315 15923
rect 259 15849 315 15858
rect 627 15914 683 15923
rect 627 15849 683 15858
rect 995 15914 1051 15923
rect 995 15849 1051 15858
rect 1363 15914 1419 15923
rect 1363 15849 1419 15858
rect 1616 15914 1672 15923
rect 1616 15849 1672 15858
rect 1733 15912 1785 15918
rect 1733 15854 1785 15860
rect 420 15392 476 15401
rect 420 15327 476 15336
rect 1156 15392 1212 15401
rect 1745 15378 1773 15854
rect 1156 15327 1212 15336
rect 1630 15350 1773 15378
rect 1630 14879 1658 15350
rect 259 14870 315 14879
rect 259 14805 315 14814
rect 627 14870 683 14879
rect 627 14805 683 14814
rect 995 14870 1051 14879
rect 995 14805 1051 14814
rect 1363 14870 1419 14879
rect 1363 14805 1419 14814
rect 1616 14870 1672 14879
rect 1616 14805 1672 14814
rect 1733 14868 1785 14874
rect 1733 14810 1785 14816
rect 420 14272 476 14281
rect 420 14207 476 14216
rect 1156 14272 1212 14281
rect 1745 14258 1773 14810
rect 1156 14207 1212 14216
rect 1630 14230 1773 14258
rect 1630 13683 1658 14230
rect 259 13674 315 13683
rect 259 13609 315 13618
rect 627 13674 683 13683
rect 627 13609 683 13618
rect 995 13674 1051 13683
rect 995 13609 1051 13618
rect 1363 13674 1419 13683
rect 1363 13609 1419 13618
rect 1616 13674 1672 13683
rect 1616 13609 1672 13618
rect 1733 13672 1785 13678
rect 1733 13614 1785 13620
rect 420 13152 476 13161
rect 420 13087 476 13096
rect 1156 13152 1212 13161
rect 1745 13138 1773 13614
rect 1156 13087 1212 13096
rect 1630 13110 1773 13138
rect 1630 12639 1658 13110
rect 259 12630 315 12639
rect 259 12565 315 12574
rect 627 12630 683 12639
rect 627 12565 683 12574
rect 995 12630 1051 12639
rect 995 12565 1051 12574
rect 1363 12630 1419 12639
rect 1363 12565 1419 12574
rect 1616 12630 1672 12639
rect 1616 12565 1672 12574
rect 1733 12628 1785 12634
rect 1733 12570 1785 12576
rect 420 12032 476 12041
rect 420 11967 476 11976
rect 1156 12032 1212 12041
rect 1745 12018 1773 12570
rect 1156 11967 1212 11976
rect 1630 11990 1773 12018
rect 1630 11443 1658 11990
rect 259 11434 315 11443
rect 259 11369 315 11378
rect 627 11434 683 11443
rect 627 11369 683 11378
rect 995 11434 1051 11443
rect 995 11369 1051 11378
rect 1363 11434 1419 11443
rect 1363 11369 1419 11378
rect 1616 11434 1672 11443
rect 1616 11369 1672 11378
rect 1733 11432 1785 11438
rect 1733 11374 1785 11380
rect 420 10912 476 10921
rect 420 10847 476 10856
rect 1156 10912 1212 10921
rect 1745 10898 1773 11374
rect 1156 10847 1212 10856
rect 1630 10870 1773 10898
rect 1630 10399 1658 10870
rect 259 10390 315 10399
rect 259 10325 315 10334
rect 627 10390 683 10399
rect 627 10325 683 10334
rect 995 10390 1051 10399
rect 995 10325 1051 10334
rect 1363 10390 1419 10399
rect 1363 10325 1419 10334
rect 1616 10390 1672 10399
rect 1616 10325 1672 10334
rect 1733 10388 1785 10394
rect 1733 10330 1785 10336
rect 420 9792 476 9801
rect 420 9727 476 9736
rect 1156 9792 1212 9801
rect 1745 9778 1773 10330
rect 1156 9727 1212 9736
rect 1630 9750 1773 9778
rect 1630 9203 1658 9750
rect 259 9194 315 9203
rect 259 9129 315 9138
rect 627 9194 683 9203
rect 627 9129 683 9138
rect 995 9194 1051 9203
rect 995 9129 1051 9138
rect 1363 9194 1419 9203
rect 1363 9129 1419 9138
rect 1616 9194 1672 9203
rect 1616 9129 1672 9138
rect 1733 9192 1785 9198
rect 1733 9134 1785 9140
rect 420 8672 476 8681
rect 420 8607 476 8616
rect 1156 8672 1212 8681
rect 1748 8644 1776 9134
rect 1156 8607 1212 8616
rect 177 7079 229 7085
rect 177 7021 229 7027
rect 357 2854 409 2860
rect 357 2796 409 2802
rect -28 1442 28 1451
rect -28 1377 28 1386
rect 369 756 397 2796
rect 1498 920 1554 929
rect 1498 855 1554 864
rect 369 750 423 756
rect 369 698 370 750
rect 422 698 423 750
rect 369 692 423 698
rect 1259 714 1311 720
rect 137 538 144 590
rect 196 538 203 590
rect -28 26 28 35
rect 369 0 397 692
rect 1259 661 1311 662
rect 1082 609 1089 661
rect 1141 609 1311 661
rect 1842 533 1898 542
rect 1004 458 1011 510
rect 1063 458 1070 510
rect 1842 468 1898 477
rect 1940 0 1968 8560
rect 2024 8246 2052 8560
rect 2012 8240 2064 8246
rect 2012 8182 2064 8188
rect 2024 7085 2052 8182
rect 2108 8122 2136 8560
rect 2096 8116 2148 8122
rect 2096 8058 2148 8064
rect 2012 7079 2064 7085
rect 2012 7021 2064 7027
rect 2024 6206 2052 7021
rect 2012 6200 2064 6206
rect 2012 6142 2064 6148
rect 2024 0 2052 6142
rect 2108 5019 2136 8058
rect 2192 5958 2220 8560
rect 2180 5952 2232 5958
rect 2180 5894 2232 5900
rect 2096 5013 2148 5019
rect 2096 4955 2148 4961
rect 2108 1608 2136 4955
rect 2192 3556 2220 5894
rect 2178 3547 2234 3556
rect 2178 3482 2234 3491
rect 2094 1599 2150 1608
rect 2094 1534 2150 1543
rect 2108 0 2136 1534
rect 2192 0 2220 3482
rect 2276 3130 2304 8560
rect 2264 3124 2316 3130
rect 2264 3066 2316 3072
rect 2276 2860 2304 3066
rect 2264 2854 2316 2860
rect 2264 2796 2316 2802
rect 2276 2191 2304 2796
rect 2264 2185 2316 2191
rect 2264 2127 2316 2133
rect 2276 178 2304 2127
rect 2360 542 2388 8560
rect 2444 7998 2472 8560
rect 4242 8512 4298 8521
rect 4242 8447 4298 8456
rect 2432 7992 2484 7998
rect 2432 7934 2484 7940
rect 2444 3378 2472 7934
rect 3260 7803 3312 7809
rect 3312 7763 4354 7791
rect 3260 7745 3312 7751
rect 4242 7098 4298 7107
rect 4242 7033 4298 7042
rect 4134 6389 4186 6395
rect 4186 6349 4354 6377
rect 4134 6331 4186 6337
rect 4242 5684 4298 5693
rect 4242 5619 4298 5628
rect 4182 4975 4234 4981
rect 4234 4935 4354 4963
rect 4182 4917 4234 4923
rect 4242 4270 4298 4279
rect 4242 4205 4298 4214
rect 3158 3547 3214 3556
rect 3158 3482 3214 3491
rect 2432 3372 2484 3378
rect 2432 3314 2484 3320
rect 2444 2347 2472 3314
rect 4242 2856 4298 2865
rect 4242 2791 4298 2800
rect 2430 2338 2486 2347
rect 2430 2273 2486 2282
rect 3181 2338 3237 2347
rect 3181 2273 3237 2282
rect 2444 929 2472 2273
rect 3528 2163 3580 2169
rect 3528 2105 3580 2111
rect 3540 1608 3568 2105
rect 3526 1599 3582 1608
rect 3526 1534 3582 1543
rect 4242 1442 4298 1451
rect 4242 1377 4298 1386
rect 2430 920 2486 929
rect 2430 855 2486 864
rect 2346 533 2402 542
rect 2346 468 2402 477
rect 2262 169 2318 178
rect 2262 104 2318 113
rect 2276 0 2304 104
rect 2360 0 2388 468
rect 2444 0 2472 855
rect 4182 733 4234 739
rect 2667 695 2719 701
rect 4234 693 4354 721
rect 4182 675 4234 681
rect 2667 637 2719 643
rect 4194 178 4222 675
rect 4180 169 4236 178
rect 4180 104 4236 113
rect 4242 28 4298 37
rect -28 -39 28 -30
rect 4242 -37 4298 -28
<< via2 >>
rect 420 18750 476 18752
rect 420 18698 422 18750
rect 422 18698 474 18750
rect 474 18698 476 18750
rect 420 18696 476 18698
rect 1156 18750 1212 18752
rect 1156 18698 1158 18750
rect 1158 18698 1210 18750
rect 1210 18698 1212 18750
rect 1156 18696 1212 18698
rect 259 18152 315 18154
rect 259 18100 261 18152
rect 261 18100 313 18152
rect 313 18100 315 18152
rect 259 18098 315 18100
rect 627 18152 683 18154
rect 627 18100 629 18152
rect 629 18100 681 18152
rect 681 18100 683 18152
rect 627 18098 683 18100
rect 995 18152 1051 18154
rect 995 18100 997 18152
rect 997 18100 1049 18152
rect 1049 18100 1051 18152
rect 995 18098 1051 18100
rect 1363 18152 1419 18154
rect 1363 18100 1365 18152
rect 1365 18100 1417 18152
rect 1417 18100 1419 18152
rect 1363 18098 1419 18100
rect 1616 18152 1672 18154
rect 1616 18100 1618 18152
rect 1618 18100 1670 18152
rect 1670 18100 1672 18152
rect 1616 18098 1672 18100
rect 420 17630 476 17632
rect 420 17578 422 17630
rect 422 17578 474 17630
rect 474 17578 476 17630
rect 420 17576 476 17578
rect 1156 17630 1212 17632
rect 1156 17578 1158 17630
rect 1158 17578 1210 17630
rect 1210 17578 1212 17630
rect 1156 17576 1212 17578
rect 259 17108 315 17110
rect 259 17056 261 17108
rect 261 17056 313 17108
rect 313 17056 315 17108
rect 259 17054 315 17056
rect 627 17108 683 17110
rect 627 17056 629 17108
rect 629 17056 681 17108
rect 681 17056 683 17108
rect 627 17054 683 17056
rect 995 17108 1051 17110
rect 995 17056 997 17108
rect 997 17056 1049 17108
rect 1049 17056 1051 17108
rect 995 17054 1051 17056
rect 1363 17108 1419 17110
rect 1363 17056 1365 17108
rect 1365 17056 1417 17108
rect 1417 17056 1419 17108
rect 1363 17054 1419 17056
rect 1616 17108 1672 17110
rect 1616 17056 1618 17108
rect 1618 17056 1670 17108
rect 1670 17056 1672 17108
rect 1616 17054 1672 17056
rect 420 16510 476 16512
rect 420 16458 422 16510
rect 422 16458 474 16510
rect 474 16458 476 16510
rect 420 16456 476 16458
rect 1156 16510 1212 16512
rect 1156 16458 1158 16510
rect 1158 16458 1210 16510
rect 1210 16458 1212 16510
rect 1156 16456 1212 16458
rect 259 15912 315 15914
rect 259 15860 261 15912
rect 261 15860 313 15912
rect 313 15860 315 15912
rect 259 15858 315 15860
rect 627 15912 683 15914
rect 627 15860 629 15912
rect 629 15860 681 15912
rect 681 15860 683 15912
rect 627 15858 683 15860
rect 995 15912 1051 15914
rect 995 15860 997 15912
rect 997 15860 1049 15912
rect 1049 15860 1051 15912
rect 995 15858 1051 15860
rect 1363 15912 1419 15914
rect 1363 15860 1365 15912
rect 1365 15860 1417 15912
rect 1417 15860 1419 15912
rect 1363 15858 1419 15860
rect 1616 15912 1672 15914
rect 1616 15860 1618 15912
rect 1618 15860 1670 15912
rect 1670 15860 1672 15912
rect 1616 15858 1672 15860
rect 420 15390 476 15392
rect 420 15338 422 15390
rect 422 15338 474 15390
rect 474 15338 476 15390
rect 420 15336 476 15338
rect 1156 15390 1212 15392
rect 1156 15338 1158 15390
rect 1158 15338 1210 15390
rect 1210 15338 1212 15390
rect 1156 15336 1212 15338
rect 259 14868 315 14870
rect 259 14816 261 14868
rect 261 14816 313 14868
rect 313 14816 315 14868
rect 259 14814 315 14816
rect 627 14868 683 14870
rect 627 14816 629 14868
rect 629 14816 681 14868
rect 681 14816 683 14868
rect 627 14814 683 14816
rect 995 14868 1051 14870
rect 995 14816 997 14868
rect 997 14816 1049 14868
rect 1049 14816 1051 14868
rect 995 14814 1051 14816
rect 1363 14868 1419 14870
rect 1363 14816 1365 14868
rect 1365 14816 1417 14868
rect 1417 14816 1419 14868
rect 1363 14814 1419 14816
rect 1616 14868 1672 14870
rect 1616 14816 1618 14868
rect 1618 14816 1670 14868
rect 1670 14816 1672 14868
rect 1616 14814 1672 14816
rect 420 14270 476 14272
rect 420 14218 422 14270
rect 422 14218 474 14270
rect 474 14218 476 14270
rect 420 14216 476 14218
rect 1156 14270 1212 14272
rect 1156 14218 1158 14270
rect 1158 14218 1210 14270
rect 1210 14218 1212 14270
rect 1156 14216 1212 14218
rect 259 13672 315 13674
rect 259 13620 261 13672
rect 261 13620 313 13672
rect 313 13620 315 13672
rect 259 13618 315 13620
rect 627 13672 683 13674
rect 627 13620 629 13672
rect 629 13620 681 13672
rect 681 13620 683 13672
rect 627 13618 683 13620
rect 995 13672 1051 13674
rect 995 13620 997 13672
rect 997 13620 1049 13672
rect 1049 13620 1051 13672
rect 995 13618 1051 13620
rect 1363 13672 1419 13674
rect 1363 13620 1365 13672
rect 1365 13620 1417 13672
rect 1417 13620 1419 13672
rect 1363 13618 1419 13620
rect 1616 13672 1672 13674
rect 1616 13620 1618 13672
rect 1618 13620 1670 13672
rect 1670 13620 1672 13672
rect 1616 13618 1672 13620
rect 420 13150 476 13152
rect 420 13098 422 13150
rect 422 13098 474 13150
rect 474 13098 476 13150
rect 420 13096 476 13098
rect 1156 13150 1212 13152
rect 1156 13098 1158 13150
rect 1158 13098 1210 13150
rect 1210 13098 1212 13150
rect 1156 13096 1212 13098
rect 259 12628 315 12630
rect 259 12576 261 12628
rect 261 12576 313 12628
rect 313 12576 315 12628
rect 259 12574 315 12576
rect 627 12628 683 12630
rect 627 12576 629 12628
rect 629 12576 681 12628
rect 681 12576 683 12628
rect 627 12574 683 12576
rect 995 12628 1051 12630
rect 995 12576 997 12628
rect 997 12576 1049 12628
rect 1049 12576 1051 12628
rect 995 12574 1051 12576
rect 1363 12628 1419 12630
rect 1363 12576 1365 12628
rect 1365 12576 1417 12628
rect 1417 12576 1419 12628
rect 1363 12574 1419 12576
rect 1616 12628 1672 12630
rect 1616 12576 1618 12628
rect 1618 12576 1670 12628
rect 1670 12576 1672 12628
rect 1616 12574 1672 12576
rect 420 12030 476 12032
rect 420 11978 422 12030
rect 422 11978 474 12030
rect 474 11978 476 12030
rect 420 11976 476 11978
rect 1156 12030 1212 12032
rect 1156 11978 1158 12030
rect 1158 11978 1210 12030
rect 1210 11978 1212 12030
rect 1156 11976 1212 11978
rect 259 11432 315 11434
rect 259 11380 261 11432
rect 261 11380 313 11432
rect 313 11380 315 11432
rect 259 11378 315 11380
rect 627 11432 683 11434
rect 627 11380 629 11432
rect 629 11380 681 11432
rect 681 11380 683 11432
rect 627 11378 683 11380
rect 995 11432 1051 11434
rect 995 11380 997 11432
rect 997 11380 1049 11432
rect 1049 11380 1051 11432
rect 995 11378 1051 11380
rect 1363 11432 1419 11434
rect 1363 11380 1365 11432
rect 1365 11380 1417 11432
rect 1417 11380 1419 11432
rect 1363 11378 1419 11380
rect 1616 11432 1672 11434
rect 1616 11380 1618 11432
rect 1618 11380 1670 11432
rect 1670 11380 1672 11432
rect 1616 11378 1672 11380
rect 420 10910 476 10912
rect 420 10858 422 10910
rect 422 10858 474 10910
rect 474 10858 476 10910
rect 420 10856 476 10858
rect 1156 10910 1212 10912
rect 1156 10858 1158 10910
rect 1158 10858 1210 10910
rect 1210 10858 1212 10910
rect 1156 10856 1212 10858
rect 259 10388 315 10390
rect 259 10336 261 10388
rect 261 10336 313 10388
rect 313 10336 315 10388
rect 259 10334 315 10336
rect 627 10388 683 10390
rect 627 10336 629 10388
rect 629 10336 681 10388
rect 681 10336 683 10388
rect 627 10334 683 10336
rect 995 10388 1051 10390
rect 995 10336 997 10388
rect 997 10336 1049 10388
rect 1049 10336 1051 10388
rect 995 10334 1051 10336
rect 1363 10388 1419 10390
rect 1363 10336 1365 10388
rect 1365 10336 1417 10388
rect 1417 10336 1419 10388
rect 1363 10334 1419 10336
rect 1616 10388 1672 10390
rect 1616 10336 1618 10388
rect 1618 10336 1670 10388
rect 1670 10336 1672 10388
rect 1616 10334 1672 10336
rect 420 9790 476 9792
rect 420 9738 422 9790
rect 422 9738 474 9790
rect 474 9738 476 9790
rect 420 9736 476 9738
rect 1156 9790 1212 9792
rect 1156 9738 1158 9790
rect 1158 9738 1210 9790
rect 1210 9738 1212 9790
rect 1156 9736 1212 9738
rect 259 9192 315 9194
rect 259 9140 261 9192
rect 261 9140 313 9192
rect 313 9140 315 9192
rect 259 9138 315 9140
rect 627 9192 683 9194
rect 627 9140 629 9192
rect 629 9140 681 9192
rect 681 9140 683 9192
rect 627 9138 683 9140
rect 995 9192 1051 9194
rect 995 9140 997 9192
rect 997 9140 1049 9192
rect 1049 9140 1051 9192
rect 995 9138 1051 9140
rect 1363 9192 1419 9194
rect 1363 9140 1365 9192
rect 1365 9140 1417 9192
rect 1417 9140 1419 9192
rect 1363 9138 1419 9140
rect 1616 9192 1672 9194
rect 1616 9140 1618 9192
rect 1618 9140 1670 9192
rect 1670 9140 1672 9192
rect 1616 9138 1672 9140
rect 420 8670 476 8672
rect 420 8618 422 8670
rect 422 8618 474 8670
rect 474 8618 476 8670
rect 420 8616 476 8618
rect 1156 8670 1212 8672
rect 1156 8618 1158 8670
rect 1158 8618 1210 8670
rect 1210 8618 1212 8670
rect 1156 8616 1212 8618
rect -28 1440 28 1442
rect -28 1388 -26 1440
rect -26 1388 26 1440
rect 26 1388 28 1440
rect -28 1386 28 1388
rect 1498 918 1554 920
rect 1498 866 1500 918
rect 1500 866 1552 918
rect 1552 866 1554 918
rect 1498 864 1554 866
rect -28 24 28 26
rect -28 -28 -26 24
rect -26 -28 26 24
rect 26 -28 28 24
rect 1842 531 1898 533
rect 1842 479 1844 531
rect 1844 479 1896 531
rect 1896 479 1898 531
rect 1842 477 1898 479
rect 2178 3491 2234 3547
rect 2094 1543 2150 1599
rect 4242 8510 4298 8512
rect 4242 8458 4244 8510
rect 4244 8458 4296 8510
rect 4296 8458 4298 8510
rect 4242 8456 4298 8458
rect 4242 7096 4298 7098
rect 4242 7044 4244 7096
rect 4244 7044 4296 7096
rect 4296 7044 4298 7096
rect 4242 7042 4298 7044
rect 4242 5682 4298 5684
rect 4242 5630 4244 5682
rect 4244 5630 4296 5682
rect 4296 5630 4298 5682
rect 4242 5628 4298 5630
rect 4242 4268 4298 4270
rect 4242 4216 4244 4268
rect 4244 4216 4296 4268
rect 4296 4216 4298 4268
rect 4242 4214 4298 4216
rect 3158 3545 3214 3547
rect 3158 3493 3160 3545
rect 3160 3493 3212 3545
rect 3212 3493 3214 3545
rect 3158 3491 3214 3493
rect 4242 2854 4298 2856
rect 4242 2802 4244 2854
rect 4244 2802 4296 2854
rect 4296 2802 4298 2854
rect 4242 2800 4298 2802
rect 2430 2282 2486 2338
rect 3181 2336 3237 2338
rect 3181 2284 3183 2336
rect 3183 2284 3235 2336
rect 3235 2284 3237 2336
rect 3181 2282 3237 2284
rect 3526 1543 3582 1599
rect 4242 1440 4298 1442
rect 4242 1388 4244 1440
rect 4244 1388 4296 1440
rect 4296 1388 4298 1440
rect 4242 1386 4298 1388
rect 2430 864 2486 920
rect 2346 477 2402 533
rect 2262 113 2318 169
rect 4180 113 4236 169
rect 4242 26 4298 28
rect -28 -30 28 -28
rect 4242 -26 4244 26
rect 4244 -26 4296 26
rect 4296 -26 4298 26
rect 4242 -28 4298 -26
<< metal3 >>
rect 399 18752 497 18773
rect 399 18696 420 18752
rect 476 18696 497 18752
rect 399 18675 497 18696
rect 1135 18752 1233 18773
rect 1135 18696 1156 18752
rect 1212 18696 1233 18752
rect 1135 18675 1233 18696
rect 254 18156 320 18159
rect 622 18156 688 18159
rect 990 18156 1056 18159
rect 1358 18156 1424 18159
rect 1611 18156 1677 18159
rect 254 18154 1677 18156
rect 254 18098 259 18154
rect 315 18098 627 18154
rect 683 18098 995 18154
rect 1051 18098 1363 18154
rect 1419 18098 1616 18154
rect 1672 18098 1677 18154
rect 254 18096 1677 18098
rect 254 18093 320 18096
rect 622 18093 688 18096
rect 990 18093 1056 18096
rect 1358 18093 1424 18096
rect 1611 18093 1677 18096
rect 399 17632 497 17653
rect 399 17576 420 17632
rect 476 17576 497 17632
rect 399 17555 497 17576
rect 1135 17632 1233 17653
rect 1135 17576 1156 17632
rect 1212 17576 1233 17632
rect 1135 17555 1233 17576
rect 254 17112 320 17115
rect 622 17112 688 17115
rect 990 17112 1056 17115
rect 1358 17112 1424 17115
rect 1611 17112 1677 17115
rect 254 17110 1677 17112
rect 254 17054 259 17110
rect 315 17054 627 17110
rect 683 17054 995 17110
rect 1051 17054 1363 17110
rect 1419 17054 1616 17110
rect 1672 17054 1677 17110
rect 254 17052 1677 17054
rect 254 17049 320 17052
rect 622 17049 688 17052
rect 990 17049 1056 17052
rect 1358 17049 1424 17052
rect 1611 17049 1677 17052
rect 399 16512 497 16533
rect 399 16456 420 16512
rect 476 16456 497 16512
rect 399 16435 497 16456
rect 1135 16512 1233 16533
rect 1135 16456 1156 16512
rect 1212 16456 1233 16512
rect 1135 16435 1233 16456
rect 254 15916 320 15919
rect 622 15916 688 15919
rect 990 15916 1056 15919
rect 1358 15916 1424 15919
rect 1611 15916 1677 15919
rect 254 15914 1677 15916
rect 254 15858 259 15914
rect 315 15858 627 15914
rect 683 15858 995 15914
rect 1051 15858 1363 15914
rect 1419 15858 1616 15914
rect 1672 15858 1677 15914
rect 254 15856 1677 15858
rect 254 15853 320 15856
rect 622 15853 688 15856
rect 990 15853 1056 15856
rect 1358 15853 1424 15856
rect 1611 15853 1677 15856
rect 399 15392 497 15413
rect 399 15336 420 15392
rect 476 15336 497 15392
rect 399 15315 497 15336
rect 1135 15392 1233 15413
rect 1135 15336 1156 15392
rect 1212 15336 1233 15392
rect 1135 15315 1233 15336
rect 254 14872 320 14875
rect 622 14872 688 14875
rect 990 14872 1056 14875
rect 1358 14872 1424 14875
rect 1611 14872 1677 14875
rect 254 14870 1677 14872
rect 254 14814 259 14870
rect 315 14814 627 14870
rect 683 14814 995 14870
rect 1051 14814 1363 14870
rect 1419 14814 1616 14870
rect 1672 14814 1677 14870
rect 254 14812 1677 14814
rect 254 14809 320 14812
rect 622 14809 688 14812
rect 990 14809 1056 14812
rect 1358 14809 1424 14812
rect 1611 14809 1677 14812
rect 399 14272 497 14293
rect 399 14216 420 14272
rect 476 14216 497 14272
rect 399 14195 497 14216
rect 1135 14272 1233 14293
rect 1135 14216 1156 14272
rect 1212 14216 1233 14272
rect 1135 14195 1233 14216
rect 254 13676 320 13679
rect 622 13676 688 13679
rect 990 13676 1056 13679
rect 1358 13676 1424 13679
rect 1611 13676 1677 13679
rect 254 13674 1677 13676
rect 254 13618 259 13674
rect 315 13618 627 13674
rect 683 13618 995 13674
rect 1051 13618 1363 13674
rect 1419 13618 1616 13674
rect 1672 13618 1677 13674
rect 254 13616 1677 13618
rect 254 13613 320 13616
rect 622 13613 688 13616
rect 990 13613 1056 13616
rect 1358 13613 1424 13616
rect 1611 13613 1677 13616
rect 399 13152 497 13173
rect 399 13096 420 13152
rect 476 13096 497 13152
rect 399 13075 497 13096
rect 1135 13152 1233 13173
rect 1135 13096 1156 13152
rect 1212 13096 1233 13152
rect 1135 13075 1233 13096
rect 254 12632 320 12635
rect 622 12632 688 12635
rect 990 12632 1056 12635
rect 1358 12632 1424 12635
rect 1611 12632 1677 12635
rect 254 12630 1677 12632
rect 254 12574 259 12630
rect 315 12574 627 12630
rect 683 12574 995 12630
rect 1051 12574 1363 12630
rect 1419 12574 1616 12630
rect 1672 12574 1677 12630
rect 254 12572 1677 12574
rect 254 12569 320 12572
rect 622 12569 688 12572
rect 990 12569 1056 12572
rect 1358 12569 1424 12572
rect 1611 12569 1677 12572
rect 399 12032 497 12053
rect 399 11976 420 12032
rect 476 11976 497 12032
rect 399 11955 497 11976
rect 1135 12032 1233 12053
rect 1135 11976 1156 12032
rect 1212 11976 1233 12032
rect 1135 11955 1233 11976
rect 254 11436 320 11439
rect 622 11436 688 11439
rect 990 11436 1056 11439
rect 1358 11436 1424 11439
rect 1611 11436 1677 11439
rect 254 11434 1677 11436
rect 254 11378 259 11434
rect 315 11378 627 11434
rect 683 11378 995 11434
rect 1051 11378 1363 11434
rect 1419 11378 1616 11434
rect 1672 11378 1677 11434
rect 254 11376 1677 11378
rect 254 11373 320 11376
rect 622 11373 688 11376
rect 990 11373 1056 11376
rect 1358 11373 1424 11376
rect 1611 11373 1677 11376
rect 399 10912 497 10933
rect 399 10856 420 10912
rect 476 10856 497 10912
rect 399 10835 497 10856
rect 1135 10912 1233 10933
rect 1135 10856 1156 10912
rect 1212 10856 1233 10912
rect 1135 10835 1233 10856
rect 254 10392 320 10395
rect 622 10392 688 10395
rect 990 10392 1056 10395
rect 1358 10392 1424 10395
rect 1611 10392 1677 10395
rect 254 10390 1677 10392
rect 254 10334 259 10390
rect 315 10334 627 10390
rect 683 10334 995 10390
rect 1051 10334 1363 10390
rect 1419 10334 1616 10390
rect 1672 10334 1677 10390
rect 254 10332 1677 10334
rect 254 10329 320 10332
rect 622 10329 688 10332
rect 990 10329 1056 10332
rect 1358 10329 1424 10332
rect 1611 10329 1677 10332
rect 399 9792 497 9813
rect 399 9736 420 9792
rect 476 9736 497 9792
rect 399 9715 497 9736
rect 1135 9792 1233 9813
rect 1135 9736 1156 9792
rect 1212 9736 1233 9792
rect 1135 9715 1233 9736
rect 254 9196 320 9199
rect 622 9196 688 9199
rect 990 9196 1056 9199
rect 1358 9196 1424 9199
rect 1611 9196 1677 9199
rect 254 9194 1677 9196
rect 254 9138 259 9194
rect 315 9138 627 9194
rect 683 9138 995 9194
rect 1051 9138 1363 9194
rect 1419 9138 1616 9194
rect 1672 9138 1677 9194
rect 254 9136 1677 9138
rect 254 9133 320 9136
rect 622 9133 688 9136
rect 990 9133 1056 9136
rect 1358 9133 1424 9136
rect 1611 9133 1677 9136
rect 399 8672 497 8693
rect 399 8616 420 8672
rect 476 8616 497 8672
rect 399 8595 497 8616
rect 1135 8672 1233 8693
rect 1135 8616 1156 8672
rect 1212 8616 1233 8672
rect 1135 8595 1233 8616
rect 4221 8512 4319 8533
rect 4221 8456 4242 8512
rect 4298 8456 4319 8512
rect 4221 8435 4319 8456
rect 4221 7098 4319 7119
rect 4221 7042 4242 7098
rect 4298 7042 4319 7098
rect 4221 7021 4319 7042
rect 4221 5684 4319 5705
rect 4221 5628 4242 5684
rect 4298 5628 4319 5684
rect 4221 5607 4319 5628
rect 4221 4270 4319 4291
rect 4221 4214 4242 4270
rect 4298 4214 4319 4270
rect 4221 4193 4319 4214
rect 2173 3549 2239 3552
rect 3153 3549 3219 3552
rect 2173 3547 3219 3549
rect 2173 3491 2178 3547
rect 2234 3491 3158 3547
rect 3214 3491 3219 3547
rect 2173 3489 3219 3491
rect 2173 3486 2239 3489
rect 3153 3486 3219 3489
rect 4221 2856 4319 2877
rect 4221 2800 4242 2856
rect 4298 2800 4319 2856
rect 4221 2779 4319 2800
rect 2425 2340 2491 2343
rect 3176 2340 3242 2343
rect 2425 2338 3242 2340
rect 2425 2282 2430 2338
rect 2486 2282 3181 2338
rect 3237 2282 3242 2338
rect 2425 2280 3242 2282
rect 2425 2277 2491 2280
rect 3176 2277 3242 2280
rect 2089 1601 2155 1604
rect 3521 1601 3587 1604
rect 2089 1599 3587 1601
rect 2089 1543 2094 1599
rect 2150 1543 3526 1599
rect 3582 1543 3587 1599
rect 2089 1541 3587 1543
rect 2089 1538 2155 1541
rect 3521 1538 3587 1541
rect -49 1442 49 1463
rect -49 1386 -28 1442
rect 28 1386 49 1442
rect -49 1365 49 1386
rect 4221 1442 4319 1463
rect 4221 1386 4242 1442
rect 4298 1386 4319 1442
rect 4221 1365 4319 1386
rect 1493 922 1559 925
rect 2425 922 2491 925
rect 1493 920 2491 922
rect 1493 864 1498 920
rect 1554 864 2430 920
rect 2486 864 2491 920
rect 1493 862 2491 864
rect 1493 859 1559 862
rect 2425 859 2491 862
rect 1837 535 1903 538
rect 2341 535 2407 538
rect 1837 533 2407 535
rect 1837 477 1842 533
rect 1898 477 2346 533
rect 2402 477 2407 533
rect 1837 475 2407 477
rect 1837 472 1903 475
rect 2341 472 2407 475
rect 2257 171 2323 174
rect 4175 171 4241 174
rect 2257 169 4241 171
rect 2257 113 2262 169
rect 2318 113 4180 169
rect 4236 113 4241 169
rect 2257 111 4241 113
rect 2257 108 2323 111
rect 4175 108 4241 111
rect -49 26 49 47
rect 4237 31 4303 33
rect -49 -30 -28 26
rect 28 -30 49 26
rect -49 -51 49 -30
rect 4221 28 4319 31
rect 4221 -28 4242 28
rect 4298 -28 4319 28
rect 4221 -49 4319 -28
<< labels >>
rlabel locali 544 0 544 0 4 gnd
rlabel locali 548 1416 548 1416 4 vdd
rlabel locali s 1644 18126 1644 18126 4 Z
port 116 nsew
rlabel locali s 1759 18126 1759 18126 4 A
port 102 nsew
rlabel locali s 1656 18724 1656 18724 4 vdd
port 8 nsew
rlabel locali s 1656 17604 1656 17604 4 gnd
port 9 nsew
rlabel locali s 1661 18561 1661 18561 4 D
port 103 nsew
rlabel locali s 1761 18561 1761 18561 4 S
port 104 nsew
rlabel locali s 1661 17691 1661 17691 4 D
port 103 nsew
rlabel locali s 1761 17691 1761 17691 4 S
port 104 nsew
rlabel locali s 1276 18126 1276 18126 4 Z
port 116 nsew
rlabel locali s 1391 18126 1391 18126 4 A
port 102 nsew
rlabel locali s 1288 18724 1288 18724 4 vdd
port 8 nsew
rlabel locali s 1288 17604 1288 17604 4 gnd
port 9 nsew
rlabel locali s 1293 18561 1293 18561 4 D
port 103 nsew
rlabel locali s 1393 18561 1393 18561 4 S
port 104 nsew
rlabel locali s 1293 17691 1293 17691 4 D
port 103 nsew
rlabel locali s 1393 17691 1393 17691 4 S
port 104 nsew
rlabel locali s 1656 16484 1656 16484 4 vdd
port 8 nsew
rlabel locali s 1644 17082 1644 17082 4 Z
port 116 nsew
rlabel locali s 1759 17082 1759 17082 4 A
port 102 nsew
rlabel locali s 1656 16484 1656 16484 4 vdd
port 8 nsew
rlabel locali s 1656 17604 1656 17604 4 gnd
port 9 nsew
rlabel locali s 1661 16647 1661 16647 4 D
port 103 nsew
rlabel locali s 1761 16647 1761 16647 4 S
port 104 nsew
rlabel locali s 1661 17517 1661 17517 4 D
port 103 nsew
rlabel locali s 1761 17517 1761 17517 4 S
port 104 nsew
rlabel locali s 1276 17082 1276 17082 4 Z
port 116 nsew
rlabel locali s 1391 17082 1391 17082 4 A
port 102 nsew
rlabel locali s 1288 16484 1288 16484 4 vdd
port 8 nsew
rlabel locali s 1288 17604 1288 17604 4 gnd
port 9 nsew
rlabel locali s 1293 16647 1293 16647 4 D
port 103 nsew
rlabel locali s 1393 16647 1393 16647 4 S
port 104 nsew
rlabel locali s 1293 17517 1293 17517 4 D
port 103 nsew
rlabel locali s 1393 17517 1393 17517 4 S
port 104 nsew
rlabel locali s 1288 16484 1288 16484 4 vdd
port 8 nsew
rlabel locali s 920 16484 920 16484 4 vdd
port 8 nsew
rlabel locali s 908 17082 908 17082 4 Z
port 116 nsew
rlabel locali s 1023 17082 1023 17082 4 A
port 102 nsew
rlabel locali s 920 16484 920 16484 4 vdd
port 8 nsew
rlabel locali s 920 17604 920 17604 4 gnd
port 9 nsew
rlabel locali s 925 16647 925 16647 4 D
port 103 nsew
rlabel locali s 1025 16647 1025 16647 4 S
port 104 nsew
rlabel locali s 925 17517 925 17517 4 D
port 103 nsew
rlabel locali s 1025 17517 1025 17517 4 S
port 104 nsew
rlabel locali s 908 18126 908 18126 4 Z
port 116 nsew
rlabel locali s 1023 18126 1023 18126 4 A
port 102 nsew
rlabel locali s 920 18724 920 18724 4 vdd
port 8 nsew
rlabel locali s 920 17604 920 17604 4 gnd
port 9 nsew
rlabel locali s 925 18561 925 18561 4 D
port 103 nsew
rlabel locali s 1025 18561 1025 18561 4 S
port 104 nsew
rlabel locali s 925 17691 925 17691 4 D
port 103 nsew
rlabel locali s 1025 17691 1025 17691 4 S
port 104 nsew
rlabel locali s 655 18126 655 18126 4 A
port 102 nsew
rlabel locali s 552 18724 552 18724 4 vdd
port 8 nsew
rlabel locali s 552 17604 552 17604 4 gnd
port 9 nsew
rlabel locali s 557 18561 557 18561 4 D
port 103 nsew
rlabel locali s 657 18561 657 18561 4 S
port 104 nsew
rlabel locali s 557 17691 557 17691 4 D
port 103 nsew
rlabel locali s 657 17691 657 17691 4 S
port 104 nsew
rlabel locali s 287 18126 287 18126 4 A
port 102 nsew
rlabel locali s 184 18724 184 18724 4 vdd
port 8 nsew
rlabel locali s 184 17604 184 17604 4 gnd
port 9 nsew
rlabel locali s 189 18561 189 18561 4 D
port 103 nsew
rlabel locali s 289 18561 289 18561 4 S
port 104 nsew
rlabel locali s 189 17691 189 17691 4 D
port 103 nsew
rlabel locali s 289 17691 289 17691 4 S
port 104 nsew
rlabel locali s 540 17082 540 17082 4 Z
port 116 nsew
rlabel locali s 655 17082 655 17082 4 A
port 102 nsew
rlabel locali s 552 16484 552 16484 4 vdd
port 8 nsew
rlabel locali s 552 17604 552 17604 4 gnd
port 9 nsew
rlabel locali s 557 16647 557 16647 4 D
port 103 nsew
rlabel locali s 657 16647 657 16647 4 S
port 104 nsew
rlabel locali s 557 17517 557 17517 4 D
port 103 nsew
rlabel locali s 657 17517 657 17517 4 S
port 104 nsew
rlabel locali s 287 17082 287 17082 4 A
port 102 nsew
rlabel locali s 184 16484 184 16484 4 vdd
port 8 nsew
rlabel locali s 184 17604 184 17604 4 gnd
port 9 nsew
rlabel locali s 189 16647 189 16647 4 D
port 103 nsew
rlabel locali s 289 16647 289 16647 4 S
port 104 nsew
rlabel locali s 189 17517 189 17517 4 D
port 103 nsew
rlabel locali s 289 17517 289 17517 4 S
port 104 nsew
rlabel locali s 540 18126 540 18126 4 Z
port 116 nsew
rlabel locali s 552 16484 552 16484 4 vdd
port 8 nsew
rlabel locali s 184 16484 184 16484 4 vdd
port 8 nsew
rlabel locali s 655 14842 655 14842 4 A
port 102 nsew
rlabel locali s 552 14244 552 14244 4 vdd
port 8 nsew
rlabel locali s 552 15364 552 15364 4 gnd
port 9 nsew
rlabel locali s 557 14407 557 14407 4 D
port 103 nsew
rlabel locali s 657 14407 657 14407 4 S
port 104 nsew
rlabel locali s 552 14244 552 14244 4 vdd
port 8 nsew
rlabel locali s 557 14081 557 14081 4 D
port 103 nsew
rlabel locali s 657 14081 657 14081 4 S
port 104 nsew
rlabel locali s 184 14244 184 14244 4 vdd
port 8 nsew
rlabel locali s 189 14081 189 14081 4 D
port 103 nsew
rlabel locali s 289 14081 289 14081 4 S
port 104 nsew
rlabel locali s 557 15277 557 15277 4 D
port 103 nsew
rlabel locali s 657 15277 657 15277 4 S
port 104 nsew
rlabel locali s 540 15886 540 15886 4 Z
port 116 nsew
rlabel locali s 655 15886 655 15886 4 A
port 102 nsew
rlabel locali s 289 15277 289 15277 4 S
port 104 nsew
rlabel locali s 552 15364 552 15364 4 gnd
port 9 nsew
rlabel locali s 557 16321 557 16321 4 D
port 103 nsew
rlabel locali s 657 16321 657 16321 4 S
port 104 nsew
rlabel locali s 557 15451 557 15451 4 D
port 103 nsew
rlabel locali s 657 15451 657 15451 4 S
port 104 nsew
rlabel locali s 287 15886 287 15886 4 A
port 102 nsew
rlabel locali s 540 14842 540 14842 4 Z
port 116 nsew
rlabel locali s 184 15364 184 15364 4 gnd
port 9 nsew
rlabel locali s 189 16321 189 16321 4 D
port 103 nsew
rlabel locali s 289 16321 289 16321 4 S
port 104 nsew
rlabel locali s 189 15451 189 15451 4 D
port 103 nsew
rlabel locali s 289 15451 289 15451 4 S
port 104 nsew
rlabel locali s 287 14842 287 14842 4 A
port 102 nsew
rlabel locali s 184 14244 184 14244 4 vdd
port 8 nsew
rlabel locali s 184 15364 184 15364 4 gnd
port 9 nsew
rlabel locali s 189 14407 189 14407 4 D
port 103 nsew
rlabel locali s 289 14407 289 14407 4 S
port 104 nsew
rlabel locali s 189 15277 189 15277 4 D
port 103 nsew
rlabel locali s 1023 14842 1023 14842 4 A
port 102 nsew
rlabel locali s 920 14244 920 14244 4 vdd
port 8 nsew
rlabel locali s 920 15364 920 15364 4 gnd
port 9 nsew
rlabel locali s 925 14407 925 14407 4 D
port 103 nsew
rlabel locali s 1025 14407 1025 14407 4 S
port 104 nsew
rlabel locali s 925 15277 925 15277 4 D
port 103 nsew
rlabel locali s 1025 15277 1025 15277 4 S
port 104 nsew
rlabel locali s 908 15886 908 15886 4 Z
port 116 nsew
rlabel locali s 1023 15886 1023 15886 4 A
port 102 nsew
rlabel locali s 920 14244 920 14244 4 vdd
port 8 nsew
rlabel locali s 920 15364 920 15364 4 gnd
port 9 nsew
rlabel locali s 925 16321 925 16321 4 D
port 103 nsew
rlabel locali s 1025 16321 1025 16321 4 S
port 104 nsew
rlabel locali s 925 15451 925 15451 4 D
port 103 nsew
rlabel locali s 1025 15451 1025 15451 4 S
port 104 nsew
rlabel locali s 925 14081 925 14081 4 D
port 103 nsew
rlabel locali s 1025 14081 1025 14081 4 S
port 104 nsew
rlabel locali s 908 14842 908 14842 4 Z
port 116 nsew
rlabel locali s 1759 14842 1759 14842 4 A
port 102 nsew
rlabel locali s 1656 14244 1656 14244 4 vdd
port 8 nsew
rlabel locali s 1656 15364 1656 15364 4 gnd
port 9 nsew
rlabel locali s 1661 14407 1661 14407 4 D
port 103 nsew
rlabel locali s 1761 14407 1761 14407 4 S
port 104 nsew
rlabel locali s 1661 15277 1661 15277 4 D
port 103 nsew
rlabel locali s 1761 15277 1761 15277 4 S
port 104 nsew
rlabel locali s 1288 14244 1288 14244 4 vdd
port 8 nsew
rlabel locali s 1644 15886 1644 15886 4 Z
port 116 nsew
rlabel locali s 1759 15886 1759 15886 4 A
port 102 nsew
rlabel locali s 1293 14081 1293 14081 4 D
port 103 nsew
rlabel locali s 1656 15364 1656 15364 4 gnd
port 9 nsew
rlabel locali s 1661 16321 1661 16321 4 D
port 103 nsew
rlabel locali s 1761 16321 1761 16321 4 S
port 104 nsew
rlabel locali s 1661 15451 1661 15451 4 D
port 103 nsew
rlabel locali s 1761 15451 1761 15451 4 S
port 104 nsew
rlabel locali s 1393 14081 1393 14081 4 S
port 104 nsew
rlabel locali s 1656 14244 1656 14244 4 vdd
port 8 nsew
rlabel locali s 1661 14081 1661 14081 4 D
port 103 nsew
rlabel locali s 1276 15886 1276 15886 4 Z
port 116 nsew
rlabel locali s 1391 15886 1391 15886 4 A
port 102 nsew
rlabel locali s 1761 14081 1761 14081 4 S
port 104 nsew
rlabel locali s 1288 15364 1288 15364 4 gnd
port 9 nsew
rlabel locali s 1293 16321 1293 16321 4 D
port 103 nsew
rlabel locali s 1393 16321 1393 16321 4 S
port 104 nsew
rlabel locali s 1293 15451 1293 15451 4 D
port 103 nsew
rlabel locali s 1393 15451 1393 15451 4 S
port 104 nsew
rlabel locali s 1276 14842 1276 14842 4 Z
port 116 nsew
rlabel locali s 1391 14842 1391 14842 4 A
port 102 nsew
rlabel locali s 1288 14244 1288 14244 4 vdd
port 8 nsew
rlabel locali s 1288 15364 1288 15364 4 gnd
port 9 nsew
rlabel locali s 1293 14407 1293 14407 4 D
port 103 nsew
rlabel locali s 1393 14407 1393 14407 4 S
port 104 nsew
rlabel locali s 1293 15277 1293 15277 4 D
port 103 nsew
rlabel locali s 1393 15277 1393 15277 4 S
port 104 nsew
rlabel locali s 1644 14842 1644 14842 4 Z
port 116 nsew
rlabel locali s 1656 13124 1656 13124 4 gnd
port 9 nsew
rlabel locali s 1288 13124 1288 13124 4 gnd
port 9 nsew
rlabel locali s 1759 13646 1759 13646 4 A
port 102 nsew
rlabel locali s 1644 13646 1644 13646 4 Z
port 116 nsew
rlabel locali s 1293 13211 1293 13211 4 D
port 103 nsew
rlabel locali s 1393 13211 1393 13211 4 S
port 104 nsew
rlabel locali s 1661 13211 1661 13211 4 D
port 103 nsew
rlabel locali s 1761 13211 1761 13211 4 S
port 104 nsew
rlabel locali s 1276 13646 1276 13646 4 Z
port 116 nsew
rlabel locali s 1391 13646 1391 13646 4 A
port 102 nsew
rlabel locali s 1656 12004 1656 12004 4 vdd
port 8 nsew
rlabel locali s 1661 11841 1661 11841 4 D
port 103 nsew
rlabel locali s 1761 11841 1761 11841 4 S
port 104 nsew
rlabel locali s 1288 12004 1288 12004 4 vdd
port 8 nsew
rlabel locali s 1293 11841 1293 11841 4 D
port 103 nsew
rlabel locali s 1393 11841 1393 11841 4 S
port 104 nsew
rlabel locali s 1644 12602 1644 12602 4 Z
port 116 nsew
rlabel locali s 1759 12602 1759 12602 4 A
port 102 nsew
rlabel locali s 1656 12004 1656 12004 4 vdd
port 8 nsew
rlabel locali s 1656 13124 1656 13124 4 gnd
port 9 nsew
rlabel locali s 1661 12167 1661 12167 4 D
port 103 nsew
rlabel locali s 1761 12167 1761 12167 4 S
port 104 nsew
rlabel locali s 1661 13037 1661 13037 4 D
port 103 nsew
rlabel locali s 1761 13037 1761 13037 4 S
port 104 nsew
rlabel locali s 1276 12602 1276 12602 4 Z
port 116 nsew
rlabel locali s 1391 12602 1391 12602 4 A
port 102 nsew
rlabel locali s 1288 12004 1288 12004 4 vdd
port 8 nsew
rlabel locali s 1288 13124 1288 13124 4 gnd
port 9 nsew
rlabel locali s 1293 12167 1293 12167 4 D
port 103 nsew
rlabel locali s 1393 12167 1393 12167 4 S
port 104 nsew
rlabel locali s 1293 13037 1293 13037 4 D
port 103 nsew
rlabel locali s 1393 13037 1393 13037 4 S
port 104 nsew
rlabel locali s 552 12004 552 12004 4 vdd
port 8 nsew
rlabel locali s 557 11841 557 11841 4 D
port 103 nsew
rlabel locali s 657 11841 657 11841 4 S
port 104 nsew
rlabel locali s 184 12004 184 12004 4 vdd
port 8 nsew
rlabel locali s 189 11841 189 11841 4 D
port 103 nsew
rlabel locali s 289 11841 289 11841 4 S
port 104 nsew
rlabel locali s 540 12602 540 12602 4 Z
port 116 nsew
rlabel locali s 655 12602 655 12602 4 A
port 102 nsew
rlabel locali s 552 12004 552 12004 4 vdd
port 8 nsew
rlabel locali s 552 13124 552 13124 4 gnd
port 9 nsew
rlabel locali s 557 12167 557 12167 4 D
port 103 nsew
rlabel locali s 657 12167 657 12167 4 S
port 104 nsew
rlabel locali s 557 13037 557 13037 4 D
port 103 nsew
rlabel locali s 657 13037 657 13037 4 S
port 104 nsew
rlabel locali s 287 13646 287 13646 4 A
port 102 nsew
rlabel locali s 184 13124 184 13124 4 gnd
port 9 nsew
rlabel locali s 920 12004 920 12004 4 vdd
port 8 nsew
rlabel locali s 189 13211 189 13211 4 D
port 103 nsew
rlabel locali s 289 13211 289 13211 4 S
port 104 nsew
rlabel locali s 925 11841 925 11841 4 D
port 103 nsew
rlabel locali s 1025 11841 1025 11841 4 S
port 104 nsew
rlabel locali s 908 12602 908 12602 4 Z
port 116 nsew
rlabel locali s 1023 12602 1023 12602 4 A
port 102 nsew
rlabel locali s 920 12004 920 12004 4 vdd
port 8 nsew
rlabel locali s 920 13124 920 13124 4 gnd
port 9 nsew
rlabel locali s 925 12167 925 12167 4 D
port 103 nsew
rlabel locali s 1025 12167 1025 12167 4 S
port 104 nsew
rlabel locali s 925 13037 925 13037 4 D
port 103 nsew
rlabel locali s 1025 13037 1025 13037 4 S
port 104 nsew
rlabel locali s 908 13646 908 13646 4 Z
port 116 nsew
rlabel locali s 1023 13646 1023 13646 4 A
port 102 nsew
rlabel locali s 920 13124 920 13124 4 gnd
port 9 nsew
rlabel locali s 925 13211 925 13211 4 D
port 103 nsew
rlabel locali s 1025 13211 1025 13211 4 S
port 104 nsew
rlabel locali s 540 13646 540 13646 4 Z
port 116 nsew
rlabel locali s 655 13646 655 13646 4 A
port 102 nsew
rlabel locali s 552 13124 552 13124 4 gnd
port 9 nsew
rlabel locali s 557 13211 557 13211 4 D
port 103 nsew
rlabel locali s 657 13211 657 13211 4 S
port 104 nsew
rlabel locali s 287 12602 287 12602 4 A
port 102 nsew
rlabel locali s 184 12004 184 12004 4 vdd
port 8 nsew
rlabel locali s 184 13124 184 13124 4 gnd
port 9 nsew
rlabel locali s 189 12167 189 12167 4 D
port 103 nsew
rlabel locali s 289 12167 289 12167 4 S
port 104 nsew
rlabel locali s 189 13037 189 13037 4 D
port 103 nsew
rlabel locali s 289 13037 289 13037 4 S
port 104 nsew
rlabel locali s 184 9764 184 9764 4 vdd
port 8 nsew
rlabel locali s 189 9601 189 9601 4 D
port 103 nsew
rlabel locali s 289 9601 289 9601 4 S
port 104 nsew
rlabel locali s 552 9764 552 9764 4 vdd
port 8 nsew
rlabel locali s 557 9601 557 9601 4 D
port 103 nsew
rlabel locali s 657 9601 657 9601 4 S
port 104 nsew
rlabel locali s 908 11406 908 11406 4 Z
port 116 nsew
rlabel locali s 1023 10362 1023 10362 4 A
port 102 nsew
rlabel locali s 920 9764 920 9764 4 vdd
port 8 nsew
rlabel locali s 1023 11406 1023 11406 4 A
port 102 nsew
rlabel locali s 920 10884 920 10884 4 gnd
port 9 nsew
rlabel locali s 920 10884 920 10884 4 gnd
port 9 nsew
rlabel locali s 925 10971 925 10971 4 D
port 103 nsew
rlabel locali s 925 9927 925 9927 4 D
port 103 nsew
rlabel locali s 1025 9927 1025 9927 4 S
port 104 nsew
rlabel locali s 1025 10971 1025 10971 4 S
port 104 nsew
rlabel locali s 540 10362 540 10362 4 Z
port 116 nsew
rlabel locali s 655 10362 655 10362 4 A
port 102 nsew
rlabel locali s 552 9764 552 9764 4 vdd
port 8 nsew
rlabel locali s 552 10884 552 10884 4 gnd
port 9 nsew
rlabel locali s 557 9927 557 9927 4 D
port 103 nsew
rlabel locali s 657 9927 657 9927 4 S
port 104 nsew
rlabel locali s 557 10797 557 10797 4 D
port 103 nsew
rlabel locali s 657 10797 657 10797 4 S
port 104 nsew
rlabel locali s 540 11406 540 11406 4 Z
port 116 nsew
rlabel locali s 655 11406 655 11406 4 A
port 102 nsew
rlabel locali s 920 9764 920 9764 4 vdd
port 8 nsew
rlabel locali s 552 10884 552 10884 4 gnd
port 9 nsew
rlabel locali s 925 9601 925 9601 4 D
port 103 nsew
rlabel locali s 1025 9601 1025 9601 4 S
port 104 nsew
rlabel locali s 557 10971 557 10971 4 D
port 103 nsew
rlabel locali s 657 10971 657 10971 4 S
port 104 nsew
rlabel locali s 287 11406 287 11406 4 A
port 102 nsew
rlabel locali s 925 10797 925 10797 4 D
port 103 nsew
rlabel locali s 184 10884 184 10884 4 gnd
port 9 nsew
rlabel locali s 908 10362 908 10362 4 Z
port 116 nsew
rlabel locali s 1025 10797 1025 10797 4 S
port 104 nsew
rlabel locali s 189 10971 189 10971 4 D
port 103 nsew
rlabel locali s 289 10971 289 10971 4 S
port 104 nsew
rlabel locali s 287 10362 287 10362 4 A
port 102 nsew
rlabel locali s 184 9764 184 9764 4 vdd
port 8 nsew
rlabel locali s 184 10884 184 10884 4 gnd
port 9 nsew
rlabel locali s 189 9927 189 9927 4 D
port 103 nsew
rlabel locali s 289 9927 289 9927 4 S
port 104 nsew
rlabel locali s 189 10797 189 10797 4 D
port 103 nsew
rlabel locali s 289 10797 289 10797 4 S
port 104 nsew
rlabel locali s 1391 11406 1391 11406 4 A
port 102 nsew
rlabel locali s 1391 10362 1391 10362 4 A
port 102 nsew
rlabel locali s 1288 10884 1288 10884 4 gnd
port 9 nsew
rlabel locali s 1288 9764 1288 9764 4 vdd
port 8 nsew
rlabel locali s 1288 10884 1288 10884 4 gnd
port 9 nsew
rlabel locali s 1293 10971 1293 10971 4 D
port 103 nsew
rlabel locali s 1393 10971 1393 10971 4 S
port 104 nsew
rlabel locali s 1656 9764 1656 9764 4 vdd
port 8 nsew
rlabel locali s 1661 9601 1661 9601 4 D
port 103 nsew
rlabel locali s 1761 9601 1761 9601 4 S
port 104 nsew
rlabel locali s 1293 9927 1293 9927 4 D
port 103 nsew
rlabel locali s 1393 9927 1393 9927 4 S
port 104 nsew
rlabel locali s 1293 10797 1293 10797 4 D
port 103 nsew
rlabel locali s 1393 10797 1393 10797 4 S
port 104 nsew
rlabel locali s 1288 9764 1288 9764 4 vdd
port 8 nsew
rlabel locali s 1293 9601 1293 9601 4 D
port 103 nsew
rlabel locali s 1393 9601 1393 9601 4 S
port 104 nsew
rlabel locali s 1644 11406 1644 11406 4 Z
port 116 nsew
rlabel locali s 1759 11406 1759 11406 4 A
port 102 nsew
rlabel locali s 1661 10797 1661 10797 4 D
port 103 nsew
rlabel locali s 1656 10884 1656 10884 4 gnd
port 9 nsew
rlabel locali s 1761 10797 1761 10797 4 S
port 104 nsew
rlabel locali s 1276 10362 1276 10362 4 Z
port 116 nsew
rlabel locali s 1661 10971 1661 10971 4 D
port 103 nsew
rlabel locali s 1761 10971 1761 10971 4 S
port 104 nsew
rlabel locali s 1276 11406 1276 11406 4 Z
port 116 nsew
rlabel locali s 1644 10362 1644 10362 4 Z
port 116 nsew
rlabel locali s 1759 10362 1759 10362 4 A
port 102 nsew
rlabel locali s 1656 9764 1656 9764 4 vdd
port 8 nsew
rlabel locali s 1656 10884 1656 10884 4 gnd
port 9 nsew
rlabel locali s 1661 9927 1661 9927 4 D
port 103 nsew
rlabel locali s 1761 9927 1761 9927 4 S
port 104 nsew
rlabel locali s 172 18126 172 18126 4 Z
port 116 nsew
rlabel locali s 172 11406 172 11406 4 Z
port 116 nsew
rlabel locali s 172 10362 172 10362 4 Z
port 116 nsew
rlabel locali s 172 12602 172 12602 4 Z
port 116 nsew
rlabel locali s 172 15886 172 15886 4 Z
port 116 nsew
rlabel locali s 172 17082 172 17082 4 Z
port 116 nsew
rlabel locali s 172 14842 172 14842 4 Z
port 116 nsew
rlabel locali s 172 13646 172 13646 4 Z
port 116 nsew
rlabel locali s 172 9166 172 9166 4 Z
port 116 nsew
rlabel locali s 3286 7777 3286 7777 4 Z
port 116 nsew
rlabel locali s 3286 7777 3286 7777 4 Z
port 116 nsew
rlabel locali s 3274 7070 3274 7070 4 vdd
port 8 nsew
rlabel locali s 3274 8484 3274 8484 4 gnd
port 9 nsew
rlabel locali s 3286 7777 3286 7777 4 Z
port 116 nsew
rlabel locali s 3274 7070 3274 7070 4 vdd
port 8 nsew
rlabel locali s 3274 8484 3274 8484 4 gnd
port 9 nsew
rlabel locali s 3269 7321 3269 7321 4 D
port 103 nsew
rlabel locali s 3269 8233 3269 8233 4 D
port 103 nsew
rlabel locali s 3651 7070 3651 7070 4 vdd
port 8 nsew
rlabel locali s 3264 7070 3264 7070 4 vdd
port 8 nsew
rlabel locali s 3577 7070 3577 7070 4 vdd
port 8 nsew
rlabel locali s 3835 7070 3835 7070 4 vdd
port 8 nsew
rlabel locali s 4093 7070 4093 7070 4 vdd
port 8 nsew
rlabel locali s 3169 8233 3169 8233 4 S
port 104 nsew
rlabel locali s 2846 7070 2846 7070 4 vdd
port 8 nsew
rlabel locali s 3035 7070 3035 7070 4 vdd
port 8 nsew
rlabel locali s 3035 8484 3035 8484 4 gnd
port 9 nsew
rlabel locali s 2708 8214 2708 8214 4 A
port 102 nsew
rlabel locali s 2974 7966 2974 7966 4 C
port 105 nsew
rlabel locali s 2841 8090 2841 8090 4 B
port 106 nsew
rlabel locali s 3059 7317 3059 7317 4 Z
port 116 nsew
rlabel locali s 2851 7070 2851 7070 4 vdd
port 8 nsew
rlabel locali s 2851 8484 2851 8484 4 gnd
port 9 nsew
rlabel locali s 2708 8214 2708 8214 4 A
port 102 nsew
rlabel locali s 2974 7966 2974 7966 4 C
port 105 nsew
rlabel locali s 2841 8090 2841 8090 4 B
port 106 nsew
rlabel locali s 2791 7233 2791 7233 4 D
port 103 nsew
rlabel locali s 2691 7233 2691 7233 4 S
port 104 nsew
rlabel locali s 2891 7233 2891 7233 4 D
port 103 nsew
rlabel locali s 2791 7233 2791 7233 4 S
port 104 nsew
rlabel locali s 2991 7233 2991 7233 4 D
port 103 nsew
rlabel locali s 2891 7233 2891 7233 4 S
port 104 nsew
rlabel locali s 2691 8359 2691 8359 4 S
port 104 nsew
rlabel locali s 2991 8359 2991 8359 4 D
port 103 nsew
rlabel locali s 3171 7777 3171 7777 4 A
port 102 nsew
rlabel locali s 3171 7777 3171 7777 4 A
port 102 nsew
rlabel locali s 3169 7321 3169 7321 4 S
port 104 nsew
rlabel locali s 2846 5656 2846 5656 4 gnd
port 9 nsew
rlabel locali s 3159 5743 3159 5743 4 S
port 104 nsew
rlabel locali s 3109 5580 3109 5580 4 gnd
port 9 nsew
rlabel locali s 2841 6174 2841 6174 4 B
port 106 nsew
rlabel locali s 2741 5926 2741 5926 4 A
port 102 nsew
rlabel locali s 2791 6907 2791 6907 4 D
port 103 nsew
rlabel locali s 2691 6907 2691 6907 4 S
port 104 nsew
rlabel locali s 2891 6907 2891 6907 4 D
port 103 nsew
rlabel locali s 2791 6907 2791 6907 4 S
port 104 nsew
rlabel locali s 2691 5781 2691 5781 4 S
port 104 nsew
rlabel locali s 2891 5781 2891 5781 4 D
port 103 nsew
rlabel locali s 3061 4987 3061 4987 4 A
port 102 nsew
rlabel locali s 3161 6325 3161 6325 4 A
port 102 nsew
rlabel locali s 3159 5493 3159 5493 4 D
port 103 nsew
rlabel locali s 3161 6325 3161 6325 4 A
port 102 nsew
rlabel locali s 3176 4987 3176 4987 4 Z
port 116 nsew
rlabel locali s 3059 5493 3059 5493 4 S
port 104 nsew
rlabel locali s 2693 4987 2693 4987 4 A
port 102 nsew
rlabel locali s 2808 4987 2808 4987 4 Z
port 116 nsew
rlabel locali s 2693 4987 2693 4987 4 A
port 102 nsew
rlabel locali s 2959 6807 2959 6807 4 Z
port 116 nsew
rlabel locali s 2796 5656 2796 5656 4 gnd
port 9 nsew
rlabel locali s 2791 5569 2791 5569 4 D
port 103 nsew
rlabel locali s 2691 5569 2691 5569 4 S
port 104 nsew
rlabel locali s 3159 6907 3159 6907 4 S
port 104 nsew
rlabel locali s 3883 5656 3883 5656 4 gnd
port 9 nsew
rlabel locali s 3933 5437 3933 5437 4 D
port 103 nsew
rlabel locali s 3833 5437 3833 5437 4 S
port 104 nsew
rlabel locali s 4208 4949 4208 4949 4 Z
port 116 nsew
rlabel locali s 4093 4949 4093 4949 4 A
port 102 nsew
rlabel locali s 4141 5656 4141 5656 4 gnd
port 9 nsew
rlabel locali s 4191 5405 4191 5405 4 D
port 103 nsew
rlabel locali s 4091 5405 4091 5405 4 S
port 104 nsew
rlabel locali s 4208 4949 4208 4949 4 Z
port 116 nsew
rlabel locali s 3441 5656 3441 5656 4 gnd
port 9 nsew
rlabel locali s 3434 4968 3434 4968 4 Z
port 116 nsew
rlabel locali s 3319 4968 3319 4968 4 A
port 102 nsew
rlabel locali s 3367 5656 3367 5656 4 gnd
port 9 nsew
rlabel locali s 3417 5531 3417 5531 4 D
port 103 nsew
rlabel locali s 3317 5531 3317 5531 4 S
port 104 nsew
rlabel locali s 3692 4949 3692 4949 4 Z
port 116 nsew
rlabel locali s 3577 4949 3577 4949 4 A
port 102 nsew
rlabel locali s 4160 6363 4160 6363 4 Z
port 116 nsew
rlabel locali s 3625 5656 3625 5656 4 gnd
port 9 nsew
rlabel locali s 3651 5656 3651 5656 4 gnd
port 9 nsew
rlabel locali s 3276 6325 3276 6325 4 Z
port 116 nsew
rlabel locali s 3675 5405 3675 5405 4 D
port 103 nsew
rlabel locali s 3264 5656 3264 5656 4 gnd
port 9 nsew
rlabel locali s 3259 6907 3259 6907 4 D
port 103 nsew
rlabel locali s 3259 5743 3259 5743 4 D
port 103 nsew
rlabel locali s 3644 6344 3644 6344 4 Z
port 116 nsew
rlabel locali s 3529 6344 3529 6344 4 A
port 102 nsew
rlabel locali s 3575 5405 3575 5405 4 S
port 104 nsew
rlabel locali s 3577 5656 3577 5656 4 gnd
port 9 nsew
rlabel locali s 3627 6907 3627 6907 4 D
port 103 nsew
rlabel locali s 3527 6907 3527 6907 4 S
port 104 nsew
rlabel locali s 3627 5781 3627 5781 4 D
port 103 nsew
rlabel locali s 3527 5781 3527 5781 4 S
port 104 nsew
rlabel locali s 3902 6326 3902 6326 4 Z
port 116 nsew
rlabel locali s 3787 6326 3787 6326 4 A
port 102 nsew
rlabel locali s 3950 4965 3950 4965 4 Z
port 116 nsew
rlabel locali s 3835 5656 3835 5656 4 gnd
port 9 nsew
rlabel locali s 3885 6819 3885 6819 4 D
port 103 nsew
rlabel locali s 3785 6819 3785 6819 4 S
port 104 nsew
rlabel locali s 3885 5833 3885 5833 4 D
port 103 nsew
rlabel locali s 3785 5833 3785 5833 4 S
port 104 nsew
rlabel locali s 4160 6363 4160 6363 4 Z
port 116 nsew
rlabel locali s 4045 6363 4045 6363 4 A
port 102 nsew
rlabel locali s 3835 4965 3835 4965 4 A
port 102 nsew
rlabel locali s 4093 5656 4093 5656 4 gnd
port 9 nsew
rlabel locali s 4143 6819 4143 6819 4 D
port 103 nsew
rlabel locali s 4043 6819 4043 6819 4 S
port 104 nsew
rlabel locali s 4143 5907 4143 5907 4 D
port 103 nsew
rlabel locali s 4043 5907 4043 5907 4 S
port 104 nsew
rlabel locali s 1276 9166 1276 9166 4 Z
port 116 nsew
rlabel locali s 1391 9166 1391 9166 4 A
port 102 nsew
rlabel locali s 1025 8731 1025 8731 4 S
port 104 nsew
rlabel locali s 1288 8644 1288 8644 4 gnd
port 9 nsew
rlabel locali s 1644 9166 1644 9166 4 Z
port 116 nsew
rlabel locali s 1759 9166 1759 9166 4 A
port 102 nsew
rlabel locali s 920 8644 920 8644 4 gnd
port 9 nsew
rlabel locali s 1656 8644 1656 8644 4 gnd
port 9 nsew
rlabel locali s 1023 9166 1023 9166 4 A
port 102 nsew
rlabel locali s 287 9166 287 9166 4 A
port 102 nsew
rlabel locali s 1293 8731 1293 8731 4 D
port 103 nsew
rlabel locali s 184 8644 184 8644 4 gnd
port 9 nsew
rlabel locali s 1661 8731 1661 8731 4 D
port 103 nsew
rlabel locali s 1761 8731 1761 8731 4 S
port 104 nsew
rlabel locali s 189 8731 189 8731 4 D
port 103 nsew
rlabel locali s 289 8731 289 8731 4 S
port 104 nsew
rlabel locali s 540 9166 540 9166 4 Z
port 116 nsew
rlabel locali s 655 9166 655 9166 4 A
port 102 nsew
rlabel locali s 1393 8731 1393 8731 4 S
port 104 nsew
rlabel locali s 552 8644 552 8644 4 gnd
port 9 nsew
rlabel locali s 908 9166 908 9166 4 Z
port 116 nsew
rlabel locali s 925 8731 925 8731 4 D
port 103 nsew
rlabel locali s 557 8731 557 8731 4 D
port 103 nsew
rlabel locali s 657 8731 657 8731 4 S
port 104 nsew
rlabel locali s 1768 709 1768 709 4 Z
port 116 nsew
rlabel locali s 1653 709 1653 709 4 A
port 102 nsew
rlabel locali s 1756 1414 1756 1414 4 vdd
port 8 nsew
rlabel locali s 1756 0 1756 0 4 gnd
port 9 nsew
rlabel locali s 1751 1198 1751 1198 4 D
port 103 nsew
rlabel locali s 1651 1198 1651 1198 4 S
port 104 nsew
rlabel locali s 1751 219 1751 219 4 D
port 103 nsew
rlabel locali s 1651 219 1651 219 4 S
port 104 nsew
rlabel locali s 970 1414 970 1414 4 vdd
port 8 nsew
rlabel locali s 970 -2 970 -2 4 gnd
port 9 nsew
rlabel locali s 584 1414 584 1414 4 vdd
port 8 nsew
rlabel locali s 584 0 584 0 4 gnd
port 9 nsew
rlabel locali s 1400 688 1400 688 4 Z
port 116 nsew
rlabel locali s 1285 688 1285 688 4 A
port 102 nsew
rlabel locali s 1388 1414 1388 1414 4 vdd
port 8 nsew
rlabel locali s 1388 0 1388 0 4 gnd
port 9 nsew
rlabel locali s 1383 1251 1383 1251 4 D
port 103 nsew
rlabel locali s 1283 1251 1283 1251 4 S
port 104 nsew
rlabel locali s 1383 125 1383 125 4 D
port 103 nsew
rlabel locali s 1283 125 1283 125 4 S
port 104 nsew
rlabel locali s 3542 2828 3542 2828 4 gnd
port 9 nsew
rlabel locali s 3883 4242 3883 4242 4 vdd
port 8 nsew
rlabel locali s 3537 2609 3537 2609 4 D
port 103 nsew
rlabel locali s 3933 4493 3933 4493 4 D
port 103 nsew
rlabel locali s 3833 4493 3833 4493 4 S
port 104 nsew
rlabel locali s 3437 2609 3437 2609 4 S
port 104 nsew
rlabel locali s 3353 2828 3353 2828 4 gnd
port 9 nsew
rlabel locali s 4141 4242 4141 4242 4 vdd
port 8 nsew
rlabel locali s 4191 4493 4191 4493 4 D
port 103 nsew
rlabel locali s 4091 4493 4091 4493 4 S
port 104 nsew
rlabel locali s 3259 2703 3259 2703 4 D
port 103 nsew
rlabel locali s 3367 4242 3367 4242 4 vdd
port 8 nsew
rlabel locali s 3417 4405 3417 4405 4 D
port 103 nsew
rlabel locali s 3317 4405 3317 4405 4 S
port 104 nsew
rlabel locali s 3441 4242 3441 4242 4 vdd
port 8 nsew
rlabel locali s 3542 2828 3542 2828 4 gnd
port 9 nsew
rlabel locali s 3625 4242 3625 4242 4 vdd
port 8 nsew
rlabel locali s 3675 4493 3675 4493 4 D
port 103 nsew
rlabel locali s 3575 4493 3575 4493 4 S
port 104 nsew
rlabel locali s 3059 2703 3059 2703 4 S
port 104 nsew
rlabel locali s 3186 3519 3186 3519 4 Z
port 116 nsew
rlabel locali s 2741 3098 2741 3098 4 A
port 102 nsew
rlabel locali s 3109 4242 3109 4242 4 vdd
port 8 nsew
rlabel locali s 2985 4242 2985 4242 4 vdd
port 8 nsew
rlabel locali s 3159 4405 3159 4405 4 D
port 103 nsew
rlabel locali s 3059 4405 3059 4405 4 S
port 104 nsew
rlabel locali s 2985 2828 2985 2828 4 gnd
port 9 nsew
rlabel locali s 2841 3346 2841 3346 4 B
port 106 nsew
rlabel locali s 2959 3979 2959 3979 4 Z
port 116 nsew
rlabel locali s 2801 2828 2801 2828 4 gnd
port 9 nsew
rlabel locali s 2801 4242 2801 4242 4 vdd
port 8 nsew
rlabel locali s 2841 3346 2841 3346 4 B
port 106 nsew
rlabel locali s 2741 3098 2741 3098 4 A
port 102 nsew
rlabel locali s 2791 4079 2791 4079 4 D
port 103 nsew
rlabel locali s 2691 4079 2691 4079 4 S
port 104 nsew
rlabel locali s 2891 4079 2891 4079 4 D
port 103 nsew
rlabel locali s 2791 4079 2791 4079 4 S
port 104 nsew
rlabel locali s 2691 2953 2691 2953 4 S
port 104 nsew
rlabel locali s 2796 2828 2796 2828 4 gnd
port 9 nsew
rlabel locali s 2791 2741 2791 2741 4 D
port 103 nsew
rlabel locali s 2691 2741 2691 2741 4 S
port 104 nsew
rlabel locali s 2891 2953 2891 2953 4 D
port 103 nsew
rlabel locali s 3186 3519 3186 3519 4 Z
port 116 nsew
rlabel locali s 3071 3519 3071 3519 4 A
port 102 nsew
rlabel locali s 3174 4242 3174 4242 4 vdd
port 8 nsew
rlabel locali s 3174 2828 3174 2828 4 gnd
port 9 nsew
rlabel locali s 3186 3519 3186 3519 4 Z
port 116 nsew
rlabel locali s 3071 3519 3071 3519 4 A
port 102 nsew
rlabel locali s 3174 4242 3174 4242 4 vdd
port 8 nsew
rlabel locali s 3174 2828 3174 2828 4 gnd
port 9 nsew
rlabel locali s 3169 3991 3169 3991 4 D
port 103 nsew
rlabel locali s 3069 3991 3069 3991 4 S
port 104 nsew
rlabel locali s 3169 3047 3169 3047 4 D
port 103 nsew
rlabel locali s 3069 3047 3069 3047 4 S
port 104 nsew
rlabel locali s 3109 2558 3109 2558 4 A
port 102 nsew
rlabel locali s 3169 2828 3169 2828 4 gnd
port 9 nsew
rlabel locali s 3109 2558 3109 2558 4 A
port 102 nsew
rlabel locali s 2796 4242 2796 4242 4 vdd
port 8 nsew
rlabel locali s 2791 4405 2791 4405 4 D
port 103 nsew
rlabel locali s 2691 4405 2691 4405 4 S
port 104 nsew
rlabel locali s 2693 2159 2693 2159 4 A
port 102 nsew
rlabel locali s 2796 1414 2796 1414 4 vdd
port 8 nsew
rlabel locali s 3159 87 3159 87 4 D
port 103 nsew
rlabel locali s 2791 1577 2791 1577 4 D
port 103 nsew
rlabel locali s 2691 1577 2691 1577 4 S
port 104 nsew
rlabel locali s 3059 87 3059 87 4 S
port 104 nsew
rlabel locali s 2791 1251 2791 1251 4 D
port 103 nsew
rlabel locali s 2691 1251 2691 1251 4 S
port 104 nsew
rlabel locali s 2791 87 2791 87 4 D
port 103 nsew
rlabel locali s 3169 1414 3169 1414 4 vdd
port 8 nsew
rlabel locali s 2691 87 2691 87 4 S
port 104 nsew
rlabel locali s 3159 1577 3159 1577 4 D
port 103 nsew
rlabel locali s 3176 669 3176 669 4 Z
port 116 nsew
rlabel locali s 3059 1577 3059 1577 4 S
port 104 nsew
rlabel locali s 3061 669 3061 669 4 A
port 102 nsew
rlabel locali s 3109 1414 3109 1414 4 vdd
port 8 nsew
rlabel locali s 3159 1577 3159 1577 4 S
port 104 nsew
rlabel locali s 3109 0 3109 0 4 gnd
port 9 nsew
rlabel locali s 3159 1251 3159 1251 4 D
port 103 nsew
rlabel locali s 3059 1251 3059 1251 4 S
port 104 nsew
rlabel locali s 2693 669 2693 669 4 A
port 102 nsew
rlabel locali s 2808 669 2808 669 4 Z
port 116 nsew
rlabel locali s 2693 669 2693 669 4 A
port 102 nsew
rlabel locali s 2796 1414 2796 1414 4 vdd
port 8 nsew
rlabel locali s 2796 0 2796 0 4 gnd
port 9 nsew
rlabel locali s 2808 2159 2808 2159 4 Z
port 116 nsew
rlabel locali s 3833 251 3833 251 4 S
port 104 nsew
rlabel locali s 4208 707 4208 707 4 Z
port 116 nsew
rlabel locali s 3209 2310 3209 2310 4 B
port 106 nsew
rlabel locali s 4093 707 4093 707 4 A
port 102 nsew
rlabel locali s 3209 2310 3209 2310 4 B
port 106 nsew
rlabel locali s 4141 1414 4141 1414 4 vdd
port 8 nsew
rlabel locali s 3327 1677 3327 1677 4 Z
port 116 nsew
rlabel locali s 4141 0 4141 0 4 gnd
port 9 nsew
rlabel locali s 4191 1163 4191 1163 4 D
port 103 nsew
rlabel locali s 3259 1577 3259 1577 4 D
port 103 nsew
rlabel locali s 4208 707 4208 707 4 Z
port 116 nsew
rlabel locali s 3554 2137 3554 2137 4 Z
port 116 nsew
rlabel locali s 3441 1414 3441 1414 4 vdd
port 8 nsew
rlabel locali s 3441 0 3441 0 4 gnd
port 9 nsew
rlabel locali s 3353 1414 3353 1414 4 vdd
port 8 nsew
rlabel locali s 4091 1163 4091 1163 4 S
port 104 nsew
rlabel locali s 3554 2137 3554 2137 4 Z
port 116 nsew
rlabel locali s 4191 251 4191 251 4 D
port 103 nsew
rlabel locali s 3439 2137 3439 2137 4 A
port 102 nsew
rlabel locali s 4091 251 4091 251 4 S
port 104 nsew
rlabel locali s 3883 0 3883 0 4 gnd
port 9 nsew
rlabel locali s 3537 1665 3537 1665 4 D
port 103 nsew
rlabel locali s 3542 1414 3542 1414 4 vdd
port 8 nsew
rlabel locali s 3437 1665 3437 1665 4 S
port 104 nsew
rlabel locali s 3554 2137 3554 2137 4 Z
port 116 nsew
rlabel locali s 3933 1163 3933 1163 4 D
port 103 nsew
rlabel locali s 3439 2137 3439 2137 4 A
port 102 nsew
rlabel locali s 3833 1163 3833 1163 4 S
port 104 nsew
rlabel locali s 3933 251 3933 251 4 D
port 103 nsew
rlabel locali s 3542 1414 3542 1414 4 vdd
port 8 nsew
rlabel locali s 3434 687 3434 687 4 Z
port 116 nsew
rlabel locali s 3319 687 3319 687 4 A
port 102 nsew
rlabel locali s 3367 1414 3367 1414 4 vdd
port 8 nsew
rlabel locali s 3367 0 3367 0 4 gnd
port 9 nsew
rlabel locali s 3417 1198 3417 1198 4 D
port 103 nsew
rlabel locali s 3317 1198 3317 1198 4 S
port 104 nsew
rlabel locali s 3417 177 3417 177 4 D
port 103 nsew
rlabel locali s 3317 177 3317 177 4 S
port 104 nsew
rlabel locali s 3692 691 3692 691 4 Z
port 116 nsew
rlabel locali s 3577 691 3577 691 4 A
port 102 nsew
rlabel locali s 3625 1414 3625 1414 4 vdd
port 8 nsew
rlabel locali s 3625 0 3625 0 4 gnd
port 9 nsew
rlabel locali s 3675 1163 3675 1163 4 D
port 103 nsew
rlabel locali s 3575 1163 3575 1163 4 S
port 104 nsew
rlabel locali s 3675 219 3675 219 4 D
port 103 nsew
rlabel locali s 3575 219 3575 219 4 S
port 104 nsew
rlabel locali s 3950 707 3950 707 4 Z
port 116 nsew
rlabel locali s 3835 707 3835 707 4 A
port 102 nsew
rlabel locali s 3883 1414 3883 1414 4 vdd
port 8 nsew
rlabel poly s 975 9601 975 9601 4 G
port 107 nsew
rlabel poly s 975 9927 975 9927 4 G
port 107 nsew
rlabel poly s 975 10797 975 10797 4 G
port 107 nsew
rlabel poly s 975 11841 975 11841 4 G
port 107 nsew
rlabel poly s 975 10971 975 10971 4 G
port 107 nsew
rlabel poly s 975 12167 975 12167 4 G
port 107 nsew
rlabel poly s 975 13037 975 13037 4 G
port 107 nsew
rlabel poly s 1711 14081 1711 14081 4 G
port 107 nsew
rlabel poly s 1711 13211 1711 13211 4 G
port 107 nsew
rlabel poly s 1343 14081 1343 14081 4 G
port 107 nsew
rlabel poly s 1343 13211 1343 13211 4 G
port 107 nsew
rlabel poly s 975 14081 975 14081 4 G
port 107 nsew
rlabel poly s 975 13211 975 13211 4 G
port 107 nsew
rlabel poly s 607 14081 607 14081 4 G
port 107 nsew
rlabel poly s 607 13211 607 13211 4 G
port 107 nsew
rlabel poly s 975 14407 975 14407 4 G
port 107 nsew
rlabel poly s 975 15277 975 15277 4 G
port 107 nsew
rlabel poly s 975 16321 975 16321 4 G
port 107 nsew
rlabel poly s 975 15451 975 15451 4 G
port 107 nsew
rlabel poly s 975 16647 975 16647 4 G
port 107 nsew
rlabel poly s 975 17517 975 17517 4 G
port 107 nsew
rlabel poly s 975 18561 975 18561 4 G
port 107 nsew
rlabel poly s 975 17691 975 17691 4 G
port 107 nsew
rlabel poly s 607 16321 607 16321 4 G
port 107 nsew
rlabel poly s 607 15451 607 15451 4 G
port 107 nsew
rlabel poly s 607 16647 607 16647 4 G
port 107 nsew
rlabel poly s 607 17517 607 17517 4 G
port 107 nsew
rlabel poly s 607 14407 607 14407 4 G
port 107 nsew
rlabel poly s 607 15277 607 15277 4 G
port 107 nsew
rlabel poly s 607 18561 607 18561 4 G
port 107 nsew
rlabel poly s 607 17691 607 17691 4 G
port 107 nsew
rlabel poly s 1711 18561 1711 18561 4 G
port 107 nsew
rlabel poly s 1711 17691 1711 17691 4 G
port 107 nsew
rlabel poly s 1343 18561 1343 18561 4 G
port 107 nsew
rlabel poly s 1343 17691 1343 17691 4 G
port 107 nsew
rlabel poly s 1711 16321 1711 16321 4 G
port 107 nsew
rlabel poly s 1711 15451 1711 15451 4 G
port 107 nsew
rlabel poly s 1711 16647 1711 16647 4 G
port 107 nsew
rlabel poly s 1711 17517 1711 17517 4 G
port 107 nsew
rlabel poly s 1343 16647 1343 16647 4 G
port 107 nsew
rlabel poly s 1343 17517 1343 17517 4 G
port 107 nsew
rlabel poly s 1343 16321 1343 16321 4 G
port 107 nsew
rlabel poly s 1343 15451 1343 15451 4 G
port 107 nsew
rlabel poly s 1343 14407 1343 14407 4 G
port 107 nsew
rlabel poly s 1343 15277 1343 15277 4 G
port 107 nsew
rlabel poly s 1711 14407 1711 14407 4 G
port 107 nsew
rlabel poly s 1711 15277 1711 15277 4 G
port 107 nsew
rlabel poly s 1343 9601 1343 9601 4 G
port 107 nsew
rlabel poly s 1711 11841 1711 11841 4 G
port 107 nsew
rlabel poly s 1711 10971 1711 10971 4 G
port 107 nsew
rlabel poly s 1343 11841 1343 11841 4 G
port 107 nsew
rlabel poly s 1343 10971 1343 10971 4 G
port 107 nsew
rlabel poly s 1711 9601 1711 9601 4 G
port 107 nsew
rlabel poly s 1711 12167 1711 12167 4 G
port 107 nsew
rlabel poly s 1711 13037 1711 13037 4 G
port 107 nsew
rlabel poly s 1343 12167 1343 12167 4 G
port 107 nsew
rlabel poly s 1343 13037 1343 13037 4 G
port 107 nsew
rlabel poly s 1711 9927 1711 9927 4 G
port 107 nsew
rlabel poly s 1711 10797 1711 10797 4 G
port 107 nsew
rlabel poly s 1343 9927 1343 9927 4 G
port 107 nsew
rlabel poly s 1343 10797 1343 10797 4 G
port 107 nsew
rlabel poly s 607 9927 607 9927 4 G
port 107 nsew
rlabel poly s 607 10797 607 10797 4 G
port 107 nsew
rlabel poly s 607 11841 607 11841 4 G
port 107 nsew
rlabel poly s 607 10971 607 10971 4 G
port 107 nsew
rlabel poly s 607 9601 607 9601 4 G
port 107 nsew
rlabel poly s 607 12167 607 12167 4 G
port 107 nsew
rlabel poly s 607 13037 607 13037 4 G
port 107 nsew
rlabel poly s 239 15277 239 15277 4 G
port 107 nsew
rlabel poly s 239 18561 239 18561 4 G
port 107 nsew
rlabel poly s 239 17691 239 17691 4 G
port 107 nsew
rlabel poly s 239 12167 239 12167 4 G
port 107 nsew
rlabel poly s 239 13037 239 13037 4 G
port 107 nsew
rlabel poly s 239 14081 239 14081 4 G
port 107 nsew
rlabel poly s 239 13211 239 13211 4 G
port 107 nsew
rlabel poly s 239 16647 239 16647 4 G
port 107 nsew
rlabel poly s 239 17517 239 17517 4 G
port 107 nsew
rlabel poly s 239 11841 239 11841 4 G
port 107 nsew
rlabel poly s 239 10971 239 10971 4 G
port 107 nsew
rlabel poly s 239 9927 239 9927 4 G
port 107 nsew
rlabel poly s 239 10797 239 10797 4 G
port 107 nsew
rlabel poly s 239 9601 239 9601 4 G
port 107 nsew
rlabel poly s 239 16321 239 16321 4 G
port 107 nsew
rlabel poly s 239 15451 239 15451 4 G
port 107 nsew
rlabel poly s 239 14407 239 14407 4 G
port 107 nsew
rlabel poly s 239 8731 239 8731 4 G
port 107 nsew
rlabel poly s 975 8731 975 8731 4 G
port 107 nsew
rlabel poly s 607 8731 607 8731 4 G
port 107 nsew
rlabel poly s 1711 8731 1711 8731 4 G
port 107 nsew
rlabel poly s 1343 8731 1343 8731 4 G
port 107 nsew
rlabel poly s 1333 1251 1333 1251 4 G
port 107 nsew
rlabel poly s 1333 125 1333 125 4 G
port 107 nsew
rlabel poly s 1701 1198 1701 1198 4 G
port 107 nsew
rlabel poly s 1701 219 1701 219 4 G
port 107 nsew
rlabel poly s 3109 5493 3109 5493 4 G
port 107 nsew
rlabel poly s 3109 1577 3109 1577 4 G
port 107 nsew
rlabel poly s 3209 1577 3209 1577 4 G
port 107 nsew
rlabel poly s 3109 2703 3109 2703 4 G
port 107 nsew
rlabel poly s 3209 2703 3209 2703 4 G
port 107 nsew
rlabel poly s 3487 1665 3487 1665 4 G
port 107 nsew
rlabel poly s 3487 2609 3487 2609 4 G
port 107 nsew
rlabel poly s 2741 4079 2741 4079 4 G
port 107 nsew
rlabel poly s 2841 4079 2841 4079 4 G
port 107 nsew
rlabel poly s 2741 2953 2741 2953 4 G
port 107 nsew
rlabel poly s 2841 2953 2841 2953 4 G
port 107 nsew
rlabel poly s 3119 3991 3119 3991 4 G
port 107 nsew
rlabel poly s 3119 3047 3119 3047 4 G
port 107 nsew
rlabel poly s 2741 4405 2741 4405 4 G
port 107 nsew
rlabel poly s 2741 5569 2741 5569 4 G
port 107 nsew
rlabel poly s 3109 4405 3109 4405 4 G
port 107 nsew
rlabel poly s 3367 4405 3367 4405 4 G
port 107 nsew
rlabel poly s 3367 5531 3367 5531 4 G
port 107 nsew
rlabel poly s 3625 4493 3625 4493 4 G
port 107 nsew
rlabel poly s 3625 5405 3625 5405 4 G
port 107 nsew
rlabel poly s 3883 4493 3883 4493 4 G
port 107 nsew
rlabel poly s 3883 5437 3883 5437 4 G
port 107 nsew
rlabel poly s 4141 4493 4141 4493 4 G
port 107 nsew
rlabel poly s 4141 5405 4141 5405 4 G
port 107 nsew
rlabel poly s 2741 7233 2741 7233 4 G
port 107 nsew
rlabel poly s 2841 7233 2841 7233 4 G
port 107 nsew
rlabel poly s 2941 7233 2941 7233 4 G
port 107 nsew
rlabel poly s 2741 8359 2741 8359 4 G
port 107 nsew
rlabel poly s 2841 8359 2841 8359 4 G
port 107 nsew
rlabel poly s 2941 8359 2941 8359 4 G
port 107 nsew
rlabel poly s 3219 7321 3219 7321 4 G
port 107 nsew
rlabel poly s 3219 8233 3219 8233 4 G
port 107 nsew
rlabel poly s 2741 1251 2741 1251 4 G
port 107 nsew
rlabel poly s 2741 87 2741 87 4 G
port 107 nsew
rlabel poly s 3109 1251 3109 1251 4 G
port 107 nsew
rlabel poly s 3109 87 3109 87 4 G
port 107 nsew
rlabel poly s 3367 1198 3367 1198 4 G
port 107 nsew
rlabel poly s 3367 177 3367 177 4 G
port 107 nsew
rlabel poly s 3625 1163 3625 1163 4 G
port 107 nsew
rlabel poly s 3625 219 3625 219 4 G
port 107 nsew
rlabel poly s 3883 1163 3883 1163 4 G
port 107 nsew
rlabel poly s 3883 251 3883 251 4 G
port 107 nsew
rlabel poly s 4141 1163 4141 1163 4 G
port 107 nsew
rlabel poly s 4141 251 4141 251 4 G
port 107 nsew
rlabel poly s 2741 6907 2741 6907 4 G
port 107 nsew
rlabel poly s 2841 6907 2841 6907 4 G
port 107 nsew
rlabel poly s 2741 5781 2741 5781 4 G
port 107 nsew
rlabel poly s 2841 5781 2841 5781 4 G
port 107 nsew
rlabel poly s 3209 6907 3209 6907 4 G
port 107 nsew
rlabel poly s 3209 5743 3209 5743 4 G
port 107 nsew
rlabel poly s 3577 6907 3577 6907 4 G
port 107 nsew
rlabel poly s 3577 5781 3577 5781 4 G
port 107 nsew
rlabel poly s 3835 6819 3835 6819 4 G
port 107 nsew
rlabel poly s 3835 5833 3835 5833 4 G
port 107 nsew
rlabel poly s 4093 6819 4093 6819 4 G
port 107 nsew
rlabel poly s 4093 5907 4093 5907 4 G
port 107 nsew
rlabel poly s 2741 1577 2741 1577 4 G
port 107 nsew
rlabel poly s 2741 2741 2741 2741 4 G
port 107 nsew
rlabel mvpdiff s 3159 2703 3159 2703 4 D
port 103 nsew
rlabel mvpdiff s 3159 2703 3159 2703 4 S
port 104 nsew
rlabel mvpdiff s 2791 2953 2791 2953 4 D
port 103 nsew
rlabel mvpdiff s 2791 2953 2791 2953 4 S
port 104 nsew
rlabel mvpdiff s 2791 8359 2791 8359 4 D
port 103 nsew
rlabel mvpdiff s 2891 8359 2891 8359 4 D
port 103 nsew
rlabel mvpdiff s 2791 8359 2791 8359 4 S
port 104 nsew
rlabel mvpdiff s 2891 8359 2891 8359 4 S
port 104 nsew
rlabel mvpdiff s 2791 5781 2791 5781 4 D
port 103 nsew
rlabel mvpdiff s 2791 5781 2791 5781 4 S
port 104 nsew
rlabel metal2 s 1762 8905 1762 8905 4 in
port 108 nsew
rlabel metal2 s 203 13385 203 13385 4 out
port 109 nsew
rlabel metal2 s 170 564 170 564 4 din_0
port 110 nsew
rlabel metal2 s 1870 505 1870 505 4 dout_0
port 111 nsew
rlabel metal2 s 1526 892 1526 892 4 dout_bar_0
port 112 nsew
rlabel metal2 s 383 707 383 707 4 clk
port 2 nsew
rlabel metal2 s 170 564 170 564 4 D
port 103 nsew
rlabel metal2 s 1870 505 1870 505 4 Q
port 113 nsew
rlabel metal2 s 1526 892 1526 892 4 Qb
port 114 nsew
rlabel metal2 s 396 724 396 724 4 clk
port 2 nsew
rlabel metal2 s 1146 659 1146 659 4 Q
port 113 nsew
rlabel metal2 s 419 753 419 753 4 clk
port 2 nsew
rlabel metal2 s 1007 504 1007 504 4 ON
port 115 nsew
rlabel metal2 s 139 586 139 586 4 D
port 103 nsew
rlabel metal2 s 170 564 170 564 4 D
port 103 nsew
rlabel metal2 s 1115 635 1115 635 4 Q
port 113 nsew
rlabel metal2 s 396 724 396 724 4 clk
port 2 nsew
rlabel metal2 s 1762 8905 1762 8905 4 rbl_bl
port 3 nsew
rlabel metal2 s 4257 6363 4257 6363 4 p_en_bar
port 5 nsew
rlabel metal2 s 170 564 170 564 4 csb
port 1 nsew
rlabel metal2 s 3820 7777 3820 7777 4 s_en
port 4 nsew
rlabel metal2 s 4281 707 4281 707 4 clk_buf
port 7 nsew
rlabel metal2 s 2693 669 2693 669 4 clk
port 2 nsew
rlabel metal2 s 4281 4949 4281 4949 4 wl_en
port 6 nsew
rlabel metal3 s 1184 10884 1184 10884 4 gnd
port 9 nsew
rlabel metal3 s 448 13124 448 13124 4 gnd
port 9 nsew
rlabel metal3 s 1184 13124 1184 13124 4 gnd
port 9 nsew
rlabel metal3 s 448 10884 448 10884 4 gnd
port 9 nsew
rlabel metal3 s 1184 15364 1184 15364 4 gnd
port 9 nsew
rlabel metal3 s 1184 17604 1184 17604 4 gnd
port 9 nsew
rlabel metal3 s 448 8644 448 8644 4 gnd
port 9 nsew
rlabel metal3 s 448 15364 448 15364 4 gnd
port 9 nsew
rlabel metal3 s 448 17604 448 17604 4 gnd
port 9 nsew
rlabel metal3 s 1184 8644 1184 8644 4 gnd
port 9 nsew
rlabel metal3 s 1184 18724 1184 18724 4 vdd
port 8 nsew
rlabel metal3 s 1184 16484 1184 16484 4 vdd
port 8 nsew
rlabel metal3 s 1184 12004 1184 12004 4 vdd
port 8 nsew
rlabel metal3 s 1184 12004 1184 12004 4 vdd
port 8 nsew
rlabel metal3 s 448 12004 448 12004 4 vdd
port 8 nsew
rlabel metal3 s 448 12004 448 12004 4 vdd
port 8 nsew
rlabel metal3 s 448 16484 448 16484 4 vdd
port 8 nsew
rlabel metal3 s 1184 9764 1184 9764 4 vdd
port 8 nsew
rlabel metal3 s 448 9764 448 9764 4 vdd
port 8 nsew
rlabel metal3 s 448 9764 448 9764 4 vdd
port 8 nsew
rlabel metal3 s 1184 9764 1184 9764 4 vdd
port 8 nsew
rlabel metal3 s 1184 14244 1184 14244 4 vdd
port 8 nsew
rlabel metal3 s 448 14244 448 14244 4 vdd
port 8 nsew
rlabel metal3 s 448 18724 448 18724 4 vdd
port 8 nsew
rlabel metal3 s 0 1414 0 1414 4 vdd
port 8 nsew
rlabel metal3 s 0 -2 0 -2 4 gnd
port 9 nsew
rlabel metal3 s 448 14244 448 14244 4 vdd
port 8 nsew
rlabel metal3 s 4270 7070 4270 7070 4 vdd
port 8 nsew
rlabel metal3 s 4270 4242 4270 4242 4 vdd
port 8 nsew
rlabel metal3 s 448 16484 448 16484 4 vdd
port 8 nsew
rlabel metal3 s 448 18724 448 18724 4 vdd
port 8 nsew
rlabel metal3 s 4270 1414 4270 1414 4 vdd
port 8 nsew
rlabel metal3 s 1184 12004 1184 12004 4 vdd
port 8 nsew
rlabel metal3 s 448 9764 448 9764 4 vdd
port 8 nsew
rlabel metal3 s 1184 14244 1184 14244 4 vdd
port 8 nsew
rlabel metal3 s 0 1414 0 1414 4 vdd
port 8 nsew
rlabel metal3 s 1184 9764 1184 9764 4 vdd
port 8 nsew
rlabel metal3 s 1184 18724 1184 18724 4 vdd
port 8 nsew
rlabel metal3 s 1184 16484 1184 16484 4 vdd
port 8 nsew
rlabel metal3 s 448 12004 448 12004 4 vdd
port 8 nsew
rlabel metal3 s 1184 15364 1184 15364 4 gnd
port 9 nsew
rlabel metal3 s 1184 8644 1184 8644 4 gnd
port 9 nsew
rlabel metal3 s 0 -2 0 -2 4 gnd
port 9 nsew
rlabel metal3 s 1184 17604 1184 17604 4 gnd
port 9 nsew
rlabel metal3 s 4270 2828 4270 2828 4 gnd
port 9 nsew
rlabel metal3 s 1184 10884 1184 10884 4 gnd
port 9 nsew
rlabel metal3 s 448 10884 448 10884 4 gnd
port 9 nsew
rlabel metal3 s 4270 8484 4270 8484 4 gnd
port 9 nsew
rlabel metal3 s 448 13124 448 13124 4 gnd
port 9 nsew
rlabel metal3 s 448 8644 448 8644 4 gnd
port 9 nsew
rlabel metal3 s 4270 0 4270 0 4 gnd
port 9 nsew
rlabel metal3 s 1184 13124 1184 13124 4 gnd
port 9 nsew
rlabel metal3 s 4270 5656 4270 5656 4 gnd
port 9 nsew
rlabel metal3 s 448 15364 448 15364 4 gnd
port 9 nsew
rlabel metal3 s 448 17604 448 17604 4 gnd
port 9 nsew
<< properties >>
string FIXED_BBOX 4237 -37 4303 0
string GDS_END 5901490
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 5302732
<< end >>
