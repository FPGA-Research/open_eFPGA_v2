magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< dnwell >>
rect -2090 7579 -629 14487
<< nwell >>
rect -735 14583 -431 16959
rect -2175 14281 -431 14583
rect -2175 7785 -1873 14281
rect -735 7785 -431 14281
rect -2175 7483 -431 7785
rect -735 7121 -431 7483
rect -1715 2165 -778 2897
rect -1715 1359 -1221 2091
rect -118 -451 20038 3045
<< pwell >>
rect -1813 14067 -1035 14221
rect -1813 12413 -1659 14067
rect -1189 12413 -1035 14067
rect -1813 10297 -1035 12413
rect -1813 8020 -1659 10297
rect -1189 8020 -1035 10297
rect -1813 7866 -1035 8020
<< mvnmos >>
rect -1552 11787 -1452 12387
rect -1396 11787 -1296 12387
rect -1552 11055 -1452 11655
rect -1396 11055 -1296 11655
rect -1552 10323 -1452 10923
rect -1396 10323 -1296 10923
<< mvpmos >>
rect -1596 2231 -1496 2831
rect -1440 2231 -1340 2831
rect -1153 2231 -1053 2831
rect -997 2231 -897 2831
rect -1596 1425 -1496 2025
rect -1440 1425 -1340 2025
<< mvpmosesd >>
tri 264 1436 284 1456 sw
tri 3344 1436 3364 1456 se
rect 264 1326 3364 1436
tri 3506 1436 3526 1456 sw
tri 6586 1436 6606 1456 se
tri 264 1306 284 1326 nw
tri 3344 1306 3364 1326 ne
rect 3506 1326 6606 1436
tri 3506 1306 3526 1326 nw
tri 6586 1306 6606 1326 ne
tri 6748 1436 6768 1456 sw
tri 9828 1436 9848 1456 se
rect 6748 1326 9848 1436
tri 9990 1436 10010 1456 sw
tri 13070 1436 13090 1456 se
tri 6748 1306 6768 1326 nw
tri 9828 1306 9848 1326 ne
rect 9990 1326 13090 1436
tri 9990 1306 10010 1326 nw
tri 13070 1306 13090 1326 ne
tri 13232 1436 13252 1456 sw
tri 16312 1436 16332 1456 se
rect 13232 1326 16332 1436
tri 16474 1436 16494 1456 sw
tri 19554 1436 19574 1456 se
tri 13232 1306 13252 1326 nw
tri 16312 1306 16332 1326 ne
rect 16474 1326 19574 1436
tri 16474 1306 16494 1326 nw
tri 19554 1306 19574 1326 ne
tri 264 1024 284 1044 sw
tri 3344 1024 3364 1044 se
rect 264 914 3364 1024
tri 3506 1024 3526 1044 sw
tri 6586 1024 6606 1044 se
tri 264 894 284 914 nw
tri 3344 894 3364 914 ne
rect 3506 914 6606 1024
tri 6748 1024 6768 1044 sw
tri 9828 1024 9848 1044 se
tri 3506 894 3526 914 nw
tri 6586 894 6606 914 ne
rect 6748 914 9848 1024
tri 9990 1024 10010 1044 sw
tri 13070 1024 13090 1044 se
tri 6748 894 6768 914 nw
tri 9828 894 9848 914 ne
rect 9990 914 13090 1024
tri 13232 1024 13252 1044 sw
tri 16312 1024 16332 1044 se
tri 9990 894 10010 914 nw
tri 13070 894 13090 914 ne
rect 13232 914 16332 1024
tri 13232 894 13252 914 nw
tri 16312 894 16332 914 ne
tri 16474 1024 16494 1044 sw
tri 19554 1024 19574 1044 se
rect 16474 914 19574 1024
tri 16474 894 16494 914 nw
tri 19554 894 19574 914 ne
tri 264 612 284 632 sw
tri 3344 612 3364 632 se
rect 264 502 3364 612
tri 3506 612 3526 632 sw
tri 6586 612 6606 632 se
tri 264 482 284 502 nw
tri 3344 482 3364 502 ne
rect 3506 502 6606 612
tri 6748 612 6768 632 sw
tri 9828 612 9848 632 se
tri 3506 482 3526 502 nw
tri 6586 482 6606 502 ne
rect 6748 502 9848 612
tri 9990 612 10010 632 sw
tri 13070 612 13090 632 se
tri 6748 482 6768 502 nw
tri 9828 482 9848 502 ne
rect 9990 502 13090 612
tri 13232 612 13252 632 sw
tri 16312 612 16332 632 se
tri 9990 482 10010 502 nw
tri 13070 482 13090 502 ne
rect 13232 502 16332 612
tri 16474 612 16494 632 sw
tri 19554 612 19574 632 se
tri 13232 482 13252 502 nw
tri 16312 482 16332 502 ne
rect 16474 502 19574 612
tri 16474 482 16494 502 nw
tri 19554 482 19574 502 ne
tri 264 200 284 220 sw
tri 3344 200 3364 220 se
rect 264 90 3364 200
tri 3506 200 3526 220 sw
tri 6586 200 6606 220 se
tri 264 70 284 90 nw
tri 3344 70 3364 90 ne
rect 3506 90 6606 200
tri 3506 70 3526 90 nw
tri 6586 70 6606 90 ne
tri 6748 200 6768 220 sw
tri 9828 200 9848 220 se
rect 6748 90 9848 200
tri 9990 200 10010 220 sw
tri 13070 200 13090 220 se
tri 6748 70 6768 90 nw
tri 9828 70 9848 90 ne
rect 9990 90 13090 200
tri 9990 70 10010 90 nw
tri 13070 70 13090 90 ne
tri 13232 200 13252 220 sw
tri 16312 200 16332 220 se
rect 13232 90 16332 200
tri 16474 200 16494 220 sw
tri 19554 200 19574 220 se
tri 13232 70 13252 90 nw
tri 16312 70 16332 90 ne
rect 16474 90 19574 200
tri 16474 70 16494 90 nw
tri 19554 70 19574 90 ne
<< mvndiff >>
rect -1605 12309 -1552 12387
rect -1605 12275 -1597 12309
rect -1563 12275 -1552 12309
rect -1605 12241 -1552 12275
rect -1605 12207 -1597 12241
rect -1563 12207 -1552 12241
rect -1605 12173 -1552 12207
rect -1605 12139 -1597 12173
rect -1563 12139 -1552 12173
rect -1605 12105 -1552 12139
rect -1605 12071 -1597 12105
rect -1563 12071 -1552 12105
rect -1605 12037 -1552 12071
rect -1605 12003 -1597 12037
rect -1563 12003 -1552 12037
rect -1605 11969 -1552 12003
rect -1605 11935 -1597 11969
rect -1563 11935 -1552 11969
rect -1605 11901 -1552 11935
rect -1605 11867 -1597 11901
rect -1563 11867 -1552 11901
rect -1605 11833 -1552 11867
rect -1605 11799 -1597 11833
rect -1563 11799 -1552 11833
rect -1605 11787 -1552 11799
rect -1452 12309 -1396 12387
rect -1452 12275 -1441 12309
rect -1407 12275 -1396 12309
rect -1452 12241 -1396 12275
rect -1452 12207 -1441 12241
rect -1407 12207 -1396 12241
rect -1452 12173 -1396 12207
rect -1452 12139 -1441 12173
rect -1407 12139 -1396 12173
rect -1452 12105 -1396 12139
rect -1452 12071 -1441 12105
rect -1407 12071 -1396 12105
rect -1452 12037 -1396 12071
rect -1452 12003 -1441 12037
rect -1407 12003 -1396 12037
rect -1452 11969 -1396 12003
rect -1452 11935 -1441 11969
rect -1407 11935 -1396 11969
rect -1452 11901 -1396 11935
rect -1452 11867 -1441 11901
rect -1407 11867 -1396 11901
rect -1452 11833 -1396 11867
rect -1452 11799 -1441 11833
rect -1407 11799 -1396 11833
rect -1452 11787 -1396 11799
rect -1296 12309 -1243 12387
rect -1296 12275 -1285 12309
rect -1251 12275 -1243 12309
rect -1296 12241 -1243 12275
rect -1296 12207 -1285 12241
rect -1251 12207 -1243 12241
rect -1296 12173 -1243 12207
rect -1296 12139 -1285 12173
rect -1251 12139 -1243 12173
rect -1296 12105 -1243 12139
rect -1296 12071 -1285 12105
rect -1251 12071 -1243 12105
rect -1296 12037 -1243 12071
rect -1296 12003 -1285 12037
rect -1251 12003 -1243 12037
rect -1296 11969 -1243 12003
rect -1296 11935 -1285 11969
rect -1251 11935 -1243 11969
rect -1296 11901 -1243 11935
rect -1296 11867 -1285 11901
rect -1251 11867 -1243 11901
rect -1296 11833 -1243 11867
rect -1296 11799 -1285 11833
rect -1251 11799 -1243 11833
rect -1296 11787 -1243 11799
rect -1605 11643 -1552 11655
rect -1605 11609 -1597 11643
rect -1563 11609 -1552 11643
rect -1605 11575 -1552 11609
rect -1605 11541 -1597 11575
rect -1563 11541 -1552 11575
rect -1605 11507 -1552 11541
rect -1605 11473 -1597 11507
rect -1563 11473 -1552 11507
rect -1605 11439 -1552 11473
rect -1605 11405 -1597 11439
rect -1563 11405 -1552 11439
rect -1605 11371 -1552 11405
rect -1605 11337 -1597 11371
rect -1563 11337 -1552 11371
rect -1605 11303 -1552 11337
rect -1605 11269 -1597 11303
rect -1563 11269 -1552 11303
rect -1605 11235 -1552 11269
rect -1605 11201 -1597 11235
rect -1563 11201 -1552 11235
rect -1605 11167 -1552 11201
rect -1605 11133 -1597 11167
rect -1563 11133 -1552 11167
rect -1605 11055 -1552 11133
rect -1452 11643 -1396 11655
rect -1452 11609 -1441 11643
rect -1407 11609 -1396 11643
rect -1452 11575 -1396 11609
rect -1452 11541 -1441 11575
rect -1407 11541 -1396 11575
rect -1452 11507 -1396 11541
rect -1452 11473 -1441 11507
rect -1407 11473 -1396 11507
rect -1452 11439 -1396 11473
rect -1452 11405 -1441 11439
rect -1407 11405 -1396 11439
rect -1452 11371 -1396 11405
rect -1452 11337 -1441 11371
rect -1407 11337 -1396 11371
rect -1452 11303 -1396 11337
rect -1452 11269 -1441 11303
rect -1407 11269 -1396 11303
rect -1452 11235 -1396 11269
rect -1452 11201 -1441 11235
rect -1407 11201 -1396 11235
rect -1452 11167 -1396 11201
rect -1452 11133 -1441 11167
rect -1407 11133 -1396 11167
rect -1452 11055 -1396 11133
rect -1296 11643 -1243 11655
rect -1296 11609 -1285 11643
rect -1251 11609 -1243 11643
rect -1296 11575 -1243 11609
rect -1296 11541 -1285 11575
rect -1251 11541 -1243 11575
rect -1296 11507 -1243 11541
rect -1296 11473 -1285 11507
rect -1251 11473 -1243 11507
rect -1296 11439 -1243 11473
rect -1296 11405 -1285 11439
rect -1251 11405 -1243 11439
rect -1296 11371 -1243 11405
rect -1296 11337 -1285 11371
rect -1251 11337 -1243 11371
rect -1296 11303 -1243 11337
rect -1296 11269 -1285 11303
rect -1251 11269 -1243 11303
rect -1296 11235 -1243 11269
rect -1296 11201 -1285 11235
rect -1251 11201 -1243 11235
rect -1296 11167 -1243 11201
rect -1296 11133 -1285 11167
rect -1251 11133 -1243 11167
rect -1296 11055 -1243 11133
rect -1605 10845 -1552 10923
rect -1605 10811 -1597 10845
rect -1563 10811 -1552 10845
rect -1605 10777 -1552 10811
rect -1605 10743 -1597 10777
rect -1563 10743 -1552 10777
rect -1605 10709 -1552 10743
rect -1605 10675 -1597 10709
rect -1563 10675 -1552 10709
rect -1605 10641 -1552 10675
rect -1605 10607 -1597 10641
rect -1563 10607 -1552 10641
rect -1605 10573 -1552 10607
rect -1605 10539 -1597 10573
rect -1563 10539 -1552 10573
rect -1605 10505 -1552 10539
rect -1605 10471 -1597 10505
rect -1563 10471 -1552 10505
rect -1605 10437 -1552 10471
rect -1605 10403 -1597 10437
rect -1563 10403 -1552 10437
rect -1605 10369 -1552 10403
rect -1605 10335 -1597 10369
rect -1563 10335 -1552 10369
rect -1605 10323 -1552 10335
rect -1452 10845 -1396 10923
rect -1452 10811 -1441 10845
rect -1407 10811 -1396 10845
rect -1452 10777 -1396 10811
rect -1452 10743 -1441 10777
rect -1407 10743 -1396 10777
rect -1452 10709 -1396 10743
rect -1452 10675 -1441 10709
rect -1407 10675 -1396 10709
rect -1452 10641 -1396 10675
rect -1452 10607 -1441 10641
rect -1407 10607 -1396 10641
rect -1452 10573 -1396 10607
rect -1452 10539 -1441 10573
rect -1407 10539 -1396 10573
rect -1452 10505 -1396 10539
rect -1452 10471 -1441 10505
rect -1407 10471 -1396 10505
rect -1452 10437 -1396 10471
rect -1452 10403 -1441 10437
rect -1407 10403 -1396 10437
rect -1452 10369 -1396 10403
rect -1452 10335 -1441 10369
rect -1407 10335 -1396 10369
rect -1452 10323 -1396 10335
rect -1296 10845 -1243 10923
rect -1296 10811 -1285 10845
rect -1251 10811 -1243 10845
rect -1296 10777 -1243 10811
rect -1296 10743 -1285 10777
rect -1251 10743 -1243 10777
rect -1296 10709 -1243 10743
rect -1296 10675 -1285 10709
rect -1251 10675 -1243 10709
rect -1296 10641 -1243 10675
rect -1296 10607 -1285 10641
rect -1251 10607 -1243 10641
rect -1296 10573 -1243 10607
rect -1296 10539 -1285 10573
rect -1251 10539 -1243 10573
rect -1296 10505 -1243 10539
rect -1296 10471 -1285 10505
rect -1251 10471 -1243 10505
rect -1296 10437 -1243 10471
rect -1296 10403 -1285 10437
rect -1251 10403 -1243 10437
rect -1296 10369 -1243 10403
rect -1296 10335 -1285 10369
rect -1251 10335 -1243 10369
rect -1296 10323 -1243 10335
<< mvpdiff >>
rect -1649 2819 -1596 2831
rect -1649 2785 -1641 2819
rect -1607 2785 -1596 2819
rect -1649 2751 -1596 2785
rect -1649 2717 -1641 2751
rect -1607 2717 -1596 2751
rect -1649 2683 -1596 2717
rect -1649 2649 -1641 2683
rect -1607 2649 -1596 2683
rect -1649 2615 -1596 2649
rect -1649 2581 -1641 2615
rect -1607 2581 -1596 2615
rect -1649 2547 -1596 2581
rect -1649 2513 -1641 2547
rect -1607 2513 -1596 2547
rect -1649 2479 -1596 2513
rect -1649 2445 -1641 2479
rect -1607 2445 -1596 2479
rect -1649 2411 -1596 2445
rect -1649 2377 -1641 2411
rect -1607 2377 -1596 2411
rect -1649 2343 -1596 2377
rect -1649 2309 -1641 2343
rect -1607 2309 -1596 2343
rect -1649 2231 -1596 2309
rect -1496 2819 -1440 2831
rect -1496 2785 -1485 2819
rect -1451 2785 -1440 2819
rect -1496 2751 -1440 2785
rect -1496 2717 -1485 2751
rect -1451 2717 -1440 2751
rect -1496 2683 -1440 2717
rect -1496 2649 -1485 2683
rect -1451 2649 -1440 2683
rect -1496 2615 -1440 2649
rect -1496 2581 -1485 2615
rect -1451 2581 -1440 2615
rect -1496 2547 -1440 2581
rect -1496 2513 -1485 2547
rect -1451 2513 -1440 2547
rect -1496 2479 -1440 2513
rect -1496 2445 -1485 2479
rect -1451 2445 -1440 2479
rect -1496 2411 -1440 2445
rect -1496 2377 -1485 2411
rect -1451 2377 -1440 2411
rect -1496 2343 -1440 2377
rect -1496 2309 -1485 2343
rect -1451 2309 -1440 2343
rect -1496 2231 -1440 2309
rect -1340 2819 -1287 2831
rect -1340 2785 -1329 2819
rect -1295 2785 -1287 2819
rect -1340 2751 -1287 2785
rect -1340 2717 -1329 2751
rect -1295 2717 -1287 2751
rect -1340 2683 -1287 2717
rect -1340 2649 -1329 2683
rect -1295 2649 -1287 2683
rect -1340 2615 -1287 2649
rect -1340 2581 -1329 2615
rect -1295 2581 -1287 2615
rect -1340 2547 -1287 2581
rect -1340 2513 -1329 2547
rect -1295 2513 -1287 2547
rect -1340 2479 -1287 2513
rect -1340 2445 -1329 2479
rect -1295 2445 -1287 2479
rect -1340 2411 -1287 2445
rect -1340 2377 -1329 2411
rect -1295 2377 -1287 2411
rect -1340 2343 -1287 2377
rect -1340 2309 -1329 2343
rect -1295 2309 -1287 2343
rect -1340 2231 -1287 2309
rect -1206 2819 -1153 2831
rect -1206 2785 -1198 2819
rect -1164 2785 -1153 2819
rect -1206 2751 -1153 2785
rect -1206 2717 -1198 2751
rect -1164 2717 -1153 2751
rect -1206 2683 -1153 2717
rect -1206 2649 -1198 2683
rect -1164 2649 -1153 2683
rect -1206 2615 -1153 2649
rect -1206 2581 -1198 2615
rect -1164 2581 -1153 2615
rect -1206 2547 -1153 2581
rect -1206 2513 -1198 2547
rect -1164 2513 -1153 2547
rect -1206 2479 -1153 2513
rect -1206 2445 -1198 2479
rect -1164 2445 -1153 2479
rect -1206 2411 -1153 2445
rect -1206 2377 -1198 2411
rect -1164 2377 -1153 2411
rect -1206 2343 -1153 2377
rect -1206 2309 -1198 2343
rect -1164 2309 -1153 2343
rect -1206 2231 -1153 2309
rect -1053 2819 -997 2831
rect -1053 2785 -1042 2819
rect -1008 2785 -997 2819
rect -1053 2751 -997 2785
rect -1053 2717 -1042 2751
rect -1008 2717 -997 2751
rect -1053 2683 -997 2717
rect -1053 2649 -1042 2683
rect -1008 2649 -997 2683
rect -1053 2615 -997 2649
rect -1053 2581 -1042 2615
rect -1008 2581 -997 2615
rect -1053 2547 -997 2581
rect -1053 2513 -1042 2547
rect -1008 2513 -997 2547
rect -1053 2479 -997 2513
rect -1053 2445 -1042 2479
rect -1008 2445 -997 2479
rect -1053 2411 -997 2445
rect -1053 2377 -1042 2411
rect -1008 2377 -997 2411
rect -1053 2343 -997 2377
rect -1053 2309 -1042 2343
rect -1008 2309 -997 2343
rect -1053 2231 -997 2309
rect -897 2819 -844 2831
rect -897 2785 -886 2819
rect -852 2785 -844 2819
rect -897 2751 -844 2785
rect -897 2717 -886 2751
rect -852 2717 -844 2751
rect -897 2683 -844 2717
rect -897 2649 -886 2683
rect -852 2649 -844 2683
rect -897 2615 -844 2649
rect -897 2581 -886 2615
rect -852 2581 -844 2615
rect -897 2547 -844 2581
rect -897 2513 -886 2547
rect -852 2513 -844 2547
rect -897 2479 -844 2513
rect -897 2445 -886 2479
rect -852 2445 -844 2479
rect -897 2411 -844 2445
rect -897 2377 -886 2411
rect -852 2377 -844 2411
rect -897 2343 -844 2377
rect -897 2309 -886 2343
rect -852 2309 -844 2343
rect -897 2231 -844 2309
rect -1649 2013 -1596 2025
rect -1649 1979 -1641 2013
rect -1607 1979 -1596 2013
rect -1649 1945 -1596 1979
rect -1649 1911 -1641 1945
rect -1607 1911 -1596 1945
rect -1649 1877 -1596 1911
rect -1649 1843 -1641 1877
rect -1607 1843 -1596 1877
rect -1649 1809 -1596 1843
rect -1649 1775 -1641 1809
rect -1607 1775 -1596 1809
rect -1649 1741 -1596 1775
rect -1649 1707 -1641 1741
rect -1607 1707 -1596 1741
rect -1649 1673 -1596 1707
rect -1649 1639 -1641 1673
rect -1607 1639 -1596 1673
rect -1649 1605 -1596 1639
rect -1649 1571 -1641 1605
rect -1607 1571 -1596 1605
rect -1649 1537 -1596 1571
rect -1649 1503 -1641 1537
rect -1607 1503 -1596 1537
rect -1649 1425 -1596 1503
rect -1496 2013 -1440 2025
rect -1496 1979 -1485 2013
rect -1451 1979 -1440 2013
rect -1496 1945 -1440 1979
rect -1496 1911 -1485 1945
rect -1451 1911 -1440 1945
rect -1496 1877 -1440 1911
rect -1496 1843 -1485 1877
rect -1451 1843 -1440 1877
rect -1496 1809 -1440 1843
rect -1496 1775 -1485 1809
rect -1451 1775 -1440 1809
rect -1496 1741 -1440 1775
rect -1496 1707 -1485 1741
rect -1451 1707 -1440 1741
rect -1496 1673 -1440 1707
rect -1496 1639 -1485 1673
rect -1451 1639 -1440 1673
rect -1496 1605 -1440 1639
rect -1496 1571 -1485 1605
rect -1451 1571 -1440 1605
rect -1496 1537 -1440 1571
rect -1496 1503 -1485 1537
rect -1451 1503 -1440 1537
rect -1496 1425 -1440 1503
rect -1340 2013 -1287 2025
rect -1340 1979 -1329 2013
rect -1295 1979 -1287 2013
rect -1340 1945 -1287 1979
rect -1340 1911 -1329 1945
rect -1295 1911 -1287 1945
rect -1340 1877 -1287 1911
rect -1340 1843 -1329 1877
rect -1295 1843 -1287 1877
rect -1340 1809 -1287 1843
rect -1340 1775 -1329 1809
rect -1295 1775 -1287 1809
rect -1340 1741 -1287 1775
rect -1340 1707 -1329 1741
rect -1295 1707 -1287 1741
rect -1340 1673 -1287 1707
rect -1340 1639 -1329 1673
rect -1295 1639 -1287 1673
rect -1340 1605 -1287 1639
rect -1340 1571 -1329 1605
rect -1295 1571 -1287 1605
rect -1340 1537 -1287 1571
rect -1340 1503 -1329 1537
rect -1295 1503 -1287 1537
rect -1340 1425 -1287 1503
rect 264 1638 3364 1668
rect 264 1536 364 1638
rect 2574 1604 2609 1638
rect 2643 1604 2678 1638
rect 2712 1604 2747 1638
rect 2781 1604 2816 1638
rect 2850 1604 2885 1638
rect 2919 1604 2954 1638
rect 2988 1604 3023 1638
rect 3057 1604 3092 1638
rect 3126 1604 3161 1638
rect 3195 1604 3230 1638
rect 3264 1604 3364 1638
rect 2574 1570 3364 1604
rect 2574 1536 2609 1570
rect 2643 1536 2678 1570
rect 2712 1536 2747 1570
rect 2781 1536 2816 1570
rect 2850 1536 2885 1570
rect 2919 1536 2954 1570
rect 2988 1536 3023 1570
rect 3057 1536 3092 1570
rect 3126 1536 3161 1570
rect 3195 1536 3230 1570
rect 3264 1536 3364 1570
rect 264 1456 3364 1536
rect 3506 1638 6606 1668
rect 3506 1604 3606 1638
rect 3640 1604 3675 1638
rect 3709 1604 3744 1638
rect 3778 1604 3813 1638
rect 3847 1604 3882 1638
rect 3916 1604 3951 1638
rect 3985 1604 4020 1638
rect 4054 1604 4089 1638
rect 4123 1604 4158 1638
rect 4192 1604 4227 1638
rect 4261 1604 4296 1638
rect 3506 1570 4296 1604
rect 3506 1536 3606 1570
rect 3640 1536 3675 1570
rect 3709 1536 3744 1570
rect 3778 1536 3813 1570
rect 3847 1536 3882 1570
rect 3916 1536 3951 1570
rect 3985 1536 4020 1570
rect 4054 1536 4089 1570
rect 4123 1536 4158 1570
rect 4192 1536 4227 1570
rect 4261 1536 4296 1570
rect 6506 1536 6606 1638
rect 3506 1456 6606 1536
rect 6748 1638 9848 1668
rect 6748 1536 6848 1638
rect 9058 1604 9093 1638
rect 9127 1604 9162 1638
rect 9196 1604 9231 1638
rect 9265 1604 9300 1638
rect 9334 1604 9369 1638
rect 9403 1604 9438 1638
rect 9472 1604 9507 1638
rect 9541 1604 9576 1638
rect 9610 1604 9645 1638
rect 9679 1604 9714 1638
rect 9748 1604 9848 1638
rect 9058 1570 9848 1604
rect 9058 1536 9093 1570
rect 9127 1536 9162 1570
rect 9196 1536 9231 1570
rect 9265 1536 9300 1570
rect 9334 1536 9369 1570
rect 9403 1536 9438 1570
rect 9472 1536 9507 1570
rect 9541 1536 9576 1570
rect 9610 1536 9645 1570
rect 9679 1536 9714 1570
rect 9748 1536 9848 1570
tri 264 1436 284 1456 ne
rect 284 1436 3344 1456
tri 3344 1436 3364 1456 nw
tri 3506 1436 3526 1456 ne
rect 3526 1436 6586 1456
tri 6586 1436 6606 1456 nw
tri 264 1306 284 1326 se
rect 284 1306 3344 1326
tri 3344 1306 3364 1326 sw
tri 3506 1306 3526 1326 se
rect 3526 1306 6586 1326
tri 6586 1306 6606 1326 sw
rect 264 1226 3364 1306
rect 264 1124 364 1226
rect 2574 1192 2609 1226
rect 2643 1192 2678 1226
rect 2712 1192 2747 1226
rect 2781 1192 2816 1226
rect 2850 1192 2885 1226
rect 2919 1192 2954 1226
rect 2988 1192 3023 1226
rect 3057 1192 3092 1226
rect 3126 1192 3161 1226
rect 3195 1192 3230 1226
rect 3264 1192 3364 1226
rect 2574 1158 3364 1192
rect 2574 1124 2609 1158
rect 2643 1124 2678 1158
rect 2712 1124 2747 1158
rect 2781 1124 2816 1158
rect 2850 1124 2885 1158
rect 2919 1124 2954 1158
rect 2988 1124 3023 1158
rect 3057 1124 3092 1158
rect 3126 1124 3161 1158
rect 3195 1124 3230 1158
rect 3264 1124 3364 1158
rect 264 1044 3364 1124
rect 3506 1226 6606 1306
rect 6748 1456 9848 1536
rect 9990 1638 13090 1668
rect 9990 1604 10090 1638
rect 10124 1604 10159 1638
rect 10193 1604 10228 1638
rect 10262 1604 10297 1638
rect 10331 1604 10366 1638
rect 10400 1604 10435 1638
rect 10469 1604 10504 1638
rect 10538 1604 10573 1638
rect 10607 1604 10642 1638
rect 10676 1604 10711 1638
rect 10745 1604 10780 1638
rect 9990 1570 10780 1604
rect 9990 1536 10090 1570
rect 10124 1536 10159 1570
rect 10193 1536 10228 1570
rect 10262 1536 10297 1570
rect 10331 1536 10366 1570
rect 10400 1536 10435 1570
rect 10469 1536 10504 1570
rect 10538 1536 10573 1570
rect 10607 1536 10642 1570
rect 10676 1536 10711 1570
rect 10745 1536 10780 1570
rect 12990 1536 13090 1638
rect 9990 1456 13090 1536
rect 13232 1638 16332 1668
rect 13232 1536 13332 1638
rect 15542 1604 15577 1638
rect 15611 1604 15646 1638
rect 15680 1604 15715 1638
rect 15749 1604 15784 1638
rect 15818 1604 15853 1638
rect 15887 1604 15922 1638
rect 15956 1604 15991 1638
rect 16025 1604 16060 1638
rect 16094 1604 16129 1638
rect 16163 1604 16198 1638
rect 16232 1604 16332 1638
rect 15542 1570 16332 1604
rect 15542 1536 15577 1570
rect 15611 1536 15646 1570
rect 15680 1536 15715 1570
rect 15749 1536 15784 1570
rect 15818 1536 15853 1570
rect 15887 1536 15922 1570
rect 15956 1536 15991 1570
rect 16025 1536 16060 1570
rect 16094 1536 16129 1570
rect 16163 1536 16198 1570
rect 16232 1536 16332 1570
tri 6748 1436 6768 1456 ne
rect 6768 1436 9828 1456
tri 9828 1436 9848 1456 nw
tri 9990 1436 10010 1456 ne
rect 10010 1436 13070 1456
tri 13070 1436 13090 1456 nw
tri 6748 1306 6768 1326 se
rect 6768 1306 9828 1326
tri 9828 1306 9848 1326 sw
tri 9990 1306 10010 1326 se
rect 10010 1306 13070 1326
tri 13070 1306 13090 1326 sw
rect 3506 1192 3606 1226
rect 3640 1192 3675 1226
rect 3709 1192 3744 1226
rect 3778 1192 3813 1226
rect 3847 1192 3882 1226
rect 3916 1192 3951 1226
rect 3985 1192 4020 1226
rect 4054 1192 4089 1226
rect 4123 1192 4158 1226
rect 4192 1192 4227 1226
rect 4261 1192 4296 1226
rect 3506 1158 4296 1192
rect 3506 1124 3606 1158
rect 3640 1124 3675 1158
rect 3709 1124 3744 1158
rect 3778 1124 3813 1158
rect 3847 1124 3882 1158
rect 3916 1124 3951 1158
rect 3985 1124 4020 1158
rect 4054 1124 4089 1158
rect 4123 1124 4158 1158
rect 4192 1124 4227 1158
rect 4261 1124 4296 1158
rect 6506 1124 6606 1226
rect 3506 1044 6606 1124
rect 6748 1226 9848 1306
rect 6748 1124 6848 1226
rect 9058 1192 9093 1226
rect 9127 1192 9162 1226
rect 9196 1192 9231 1226
rect 9265 1192 9300 1226
rect 9334 1192 9369 1226
rect 9403 1192 9438 1226
rect 9472 1192 9507 1226
rect 9541 1192 9576 1226
rect 9610 1192 9645 1226
rect 9679 1192 9714 1226
rect 9748 1192 9848 1226
rect 9058 1158 9848 1192
rect 9058 1124 9093 1158
rect 9127 1124 9162 1158
rect 9196 1124 9231 1158
rect 9265 1124 9300 1158
rect 9334 1124 9369 1158
rect 9403 1124 9438 1158
rect 9472 1124 9507 1158
rect 9541 1124 9576 1158
rect 9610 1124 9645 1158
rect 9679 1124 9714 1158
rect 9748 1124 9848 1158
rect 6748 1044 9848 1124
rect 9990 1226 13090 1306
rect 13232 1456 16332 1536
rect 16474 1638 19574 1668
rect 16474 1604 16574 1638
rect 16608 1604 16643 1638
rect 16677 1604 16712 1638
rect 16746 1604 16781 1638
rect 16815 1604 16850 1638
rect 16884 1604 16919 1638
rect 16953 1604 16988 1638
rect 17022 1604 17057 1638
rect 17091 1604 17126 1638
rect 17160 1604 17195 1638
rect 17229 1604 17264 1638
rect 16474 1570 17264 1604
rect 16474 1536 16574 1570
rect 16608 1536 16643 1570
rect 16677 1536 16712 1570
rect 16746 1536 16781 1570
rect 16815 1536 16850 1570
rect 16884 1536 16919 1570
rect 16953 1536 16988 1570
rect 17022 1536 17057 1570
rect 17091 1536 17126 1570
rect 17160 1536 17195 1570
rect 17229 1536 17264 1570
rect 19474 1536 19574 1638
rect 16474 1456 19574 1536
tri 13232 1436 13252 1456 ne
rect 13252 1436 16312 1456
tri 16312 1436 16332 1456 nw
tri 16474 1436 16494 1456 ne
rect 16494 1436 19554 1456
tri 19554 1436 19574 1456 nw
tri 13232 1306 13252 1326 se
rect 13252 1306 16312 1326
tri 16312 1306 16332 1326 sw
tri 16474 1306 16494 1326 se
rect 16494 1306 19554 1326
tri 19554 1306 19574 1326 sw
rect 9990 1192 10090 1226
rect 10124 1192 10159 1226
rect 10193 1192 10228 1226
rect 10262 1192 10297 1226
rect 10331 1192 10366 1226
rect 10400 1192 10435 1226
rect 10469 1192 10504 1226
rect 10538 1192 10573 1226
rect 10607 1192 10642 1226
rect 10676 1192 10711 1226
rect 10745 1192 10780 1226
rect 9990 1158 10780 1192
rect 9990 1124 10090 1158
rect 10124 1124 10159 1158
rect 10193 1124 10228 1158
rect 10262 1124 10297 1158
rect 10331 1124 10366 1158
rect 10400 1124 10435 1158
rect 10469 1124 10504 1158
rect 10538 1124 10573 1158
rect 10607 1124 10642 1158
rect 10676 1124 10711 1158
rect 10745 1124 10780 1158
rect 12990 1124 13090 1226
rect 9990 1044 13090 1124
rect 13232 1226 16332 1306
rect 13232 1124 13332 1226
rect 15542 1192 15577 1226
rect 15611 1192 15646 1226
rect 15680 1192 15715 1226
rect 15749 1192 15784 1226
rect 15818 1192 15853 1226
rect 15887 1192 15922 1226
rect 15956 1192 15991 1226
rect 16025 1192 16060 1226
rect 16094 1192 16129 1226
rect 16163 1192 16198 1226
rect 16232 1192 16332 1226
rect 15542 1158 16332 1192
rect 15542 1124 15577 1158
rect 15611 1124 15646 1158
rect 15680 1124 15715 1158
rect 15749 1124 15784 1158
rect 15818 1124 15853 1158
rect 15887 1124 15922 1158
rect 15956 1124 15991 1158
rect 16025 1124 16060 1158
rect 16094 1124 16129 1158
rect 16163 1124 16198 1158
rect 16232 1124 16332 1158
rect 13232 1044 16332 1124
rect 16474 1226 19574 1306
rect 16474 1192 16574 1226
rect 16608 1192 16643 1226
rect 16677 1192 16712 1226
rect 16746 1192 16781 1226
rect 16815 1192 16850 1226
rect 16884 1192 16919 1226
rect 16953 1192 16988 1226
rect 17022 1192 17057 1226
rect 17091 1192 17126 1226
rect 17160 1192 17195 1226
rect 17229 1192 17264 1226
rect 16474 1158 17264 1192
rect 16474 1124 16574 1158
rect 16608 1124 16643 1158
rect 16677 1124 16712 1158
rect 16746 1124 16781 1158
rect 16815 1124 16850 1158
rect 16884 1124 16919 1158
rect 16953 1124 16988 1158
rect 17022 1124 17057 1158
rect 17091 1124 17126 1158
rect 17160 1124 17195 1158
rect 17229 1124 17264 1158
rect 19474 1124 19574 1226
tri 264 1024 284 1044 ne
rect 284 1024 3344 1044
tri 3344 1024 3364 1044 nw
tri 3506 1024 3526 1044 ne
rect 3526 1024 6586 1044
tri 6586 1024 6606 1044 nw
tri 264 894 284 914 se
rect 284 894 3344 914
tri 3344 894 3364 914 sw
tri 6748 1024 6768 1044 ne
rect 6768 1024 9828 1044
tri 9828 1024 9848 1044 nw
tri 3506 894 3526 914 se
rect 3526 894 6586 914
tri 6586 894 6606 914 sw
tri 9990 1024 10010 1044 ne
rect 10010 1024 13070 1044
tri 13070 1024 13090 1044 nw
tri 6748 894 6768 914 se
rect 6768 894 9828 914
tri 9828 894 9848 914 sw
tri 13232 1024 13252 1044 ne
rect 13252 1024 16312 1044
tri 16312 1024 16332 1044 nw
tri 9990 894 10010 914 se
rect 10010 894 13070 914
tri 13070 894 13090 914 sw
tri 13232 894 13252 914 se
rect 13252 894 16312 914
tri 16312 894 16332 914 sw
rect 264 814 3364 894
rect 264 712 364 814
rect 2574 780 2609 814
rect 2643 780 2678 814
rect 2712 780 2747 814
rect 2781 780 2816 814
rect 2850 780 2885 814
rect 2919 780 2954 814
rect 2988 780 3023 814
rect 3057 780 3092 814
rect 3126 780 3161 814
rect 3195 780 3230 814
rect 3264 780 3364 814
rect 2574 746 3364 780
rect 2574 712 2609 746
rect 2643 712 2678 746
rect 2712 712 2747 746
rect 2781 712 2816 746
rect 2850 712 2885 746
rect 2919 712 2954 746
rect 2988 712 3023 746
rect 3057 712 3092 746
rect 3126 712 3161 746
rect 3195 712 3230 746
rect 3264 712 3364 746
rect 264 632 3364 712
rect 3506 814 6606 894
rect 3506 780 3606 814
rect 3640 780 3675 814
rect 3709 780 3744 814
rect 3778 780 3813 814
rect 3847 780 3882 814
rect 3916 780 3951 814
rect 3985 780 4020 814
rect 4054 780 4089 814
rect 4123 780 4158 814
rect 4192 780 4227 814
rect 4261 780 4296 814
rect 3506 746 4296 780
rect 3506 712 3606 746
rect 3640 712 3675 746
rect 3709 712 3744 746
rect 3778 712 3813 746
rect 3847 712 3882 746
rect 3916 712 3951 746
rect 3985 712 4020 746
rect 4054 712 4089 746
rect 4123 712 4158 746
rect 4192 712 4227 746
rect 4261 712 4296 746
rect 6506 712 6606 814
rect 3506 632 6606 712
rect 6748 814 9848 894
rect 6748 712 6848 814
rect 9058 780 9093 814
rect 9127 780 9162 814
rect 9196 780 9231 814
rect 9265 780 9300 814
rect 9334 780 9369 814
rect 9403 780 9438 814
rect 9472 780 9507 814
rect 9541 780 9576 814
rect 9610 780 9645 814
rect 9679 780 9714 814
rect 9748 780 9848 814
rect 9058 746 9848 780
rect 9058 712 9093 746
rect 9127 712 9162 746
rect 9196 712 9231 746
rect 9265 712 9300 746
rect 9334 712 9369 746
rect 9403 712 9438 746
rect 9472 712 9507 746
rect 9541 712 9576 746
rect 9610 712 9645 746
rect 9679 712 9714 746
rect 9748 712 9848 746
rect 6748 632 9848 712
rect 9990 814 13090 894
rect 9990 780 10090 814
rect 10124 780 10159 814
rect 10193 780 10228 814
rect 10262 780 10297 814
rect 10331 780 10366 814
rect 10400 780 10435 814
rect 10469 780 10504 814
rect 10538 780 10573 814
rect 10607 780 10642 814
rect 10676 780 10711 814
rect 10745 780 10780 814
rect 9990 746 10780 780
rect 9990 712 10090 746
rect 10124 712 10159 746
rect 10193 712 10228 746
rect 10262 712 10297 746
rect 10331 712 10366 746
rect 10400 712 10435 746
rect 10469 712 10504 746
rect 10538 712 10573 746
rect 10607 712 10642 746
rect 10676 712 10711 746
rect 10745 712 10780 746
rect 12990 712 13090 814
rect 9990 632 13090 712
rect 13232 814 16332 894
rect 16474 1044 19574 1124
tri 16474 1024 16494 1044 ne
rect 16494 1024 19554 1044
tri 19554 1024 19574 1044 nw
tri 16474 894 16494 914 se
rect 16494 894 19554 914
tri 19554 894 19574 914 sw
rect 13232 712 13332 814
rect 15542 780 15577 814
rect 15611 780 15646 814
rect 15680 780 15715 814
rect 15749 780 15784 814
rect 15818 780 15853 814
rect 15887 780 15922 814
rect 15956 780 15991 814
rect 16025 780 16060 814
rect 16094 780 16129 814
rect 16163 780 16198 814
rect 16232 780 16332 814
rect 15542 746 16332 780
rect 15542 712 15577 746
rect 15611 712 15646 746
rect 15680 712 15715 746
rect 15749 712 15784 746
rect 15818 712 15853 746
rect 15887 712 15922 746
rect 15956 712 15991 746
rect 16025 712 16060 746
rect 16094 712 16129 746
rect 16163 712 16198 746
rect 16232 712 16332 746
rect 13232 632 16332 712
rect 16474 814 19574 894
rect 16474 780 16574 814
rect 16608 780 16643 814
rect 16677 780 16712 814
rect 16746 780 16781 814
rect 16815 780 16850 814
rect 16884 780 16919 814
rect 16953 780 16988 814
rect 17022 780 17057 814
rect 17091 780 17126 814
rect 17160 780 17195 814
rect 17229 780 17264 814
rect 16474 746 17264 780
rect 16474 712 16574 746
rect 16608 712 16643 746
rect 16677 712 16712 746
rect 16746 712 16781 746
rect 16815 712 16850 746
rect 16884 712 16919 746
rect 16953 712 16988 746
rect 17022 712 17057 746
rect 17091 712 17126 746
rect 17160 712 17195 746
rect 17229 712 17264 746
rect 19474 712 19574 814
rect 16474 632 19574 712
tri 264 612 284 632 ne
rect 284 612 3344 632
tri 3344 612 3364 632 nw
tri 3506 612 3526 632 ne
rect 3526 612 6586 632
tri 6586 612 6606 632 nw
tri 264 482 284 502 se
rect 284 482 3344 502
tri 3344 482 3364 502 sw
tri 6748 612 6768 632 ne
rect 6768 612 9828 632
tri 9828 612 9848 632 nw
tri 3506 482 3526 502 se
rect 3526 482 6586 502
tri 6586 482 6606 502 sw
tri 9990 612 10010 632 ne
rect 10010 612 13070 632
tri 13070 612 13090 632 nw
tri 6748 482 6768 502 se
rect 6768 482 9828 502
tri 9828 482 9848 502 sw
tri 13232 612 13252 632 ne
rect 13252 612 16312 632
tri 16312 612 16332 632 nw
tri 9990 482 10010 502 se
rect 10010 482 13070 502
tri 13070 482 13090 502 sw
tri 16474 612 16494 632 ne
rect 16494 612 19554 632
tri 19554 612 19574 632 nw
tri 13232 482 13252 502 se
rect 13252 482 16312 502
tri 16312 482 16332 502 sw
tri 16474 482 16494 502 se
rect 16494 482 19554 502
tri 19554 482 19574 502 sw
rect 264 402 3364 482
rect 264 300 364 402
rect 2574 368 2609 402
rect 2643 368 2678 402
rect 2712 368 2747 402
rect 2781 368 2816 402
rect 2850 368 2885 402
rect 2919 368 2954 402
rect 2988 368 3023 402
rect 3057 368 3092 402
rect 3126 368 3161 402
rect 3195 368 3230 402
rect 3264 368 3364 402
rect 2574 334 3364 368
rect 2574 300 2609 334
rect 2643 300 2678 334
rect 2712 300 2747 334
rect 2781 300 2816 334
rect 2850 300 2885 334
rect 2919 300 2954 334
rect 2988 300 3023 334
rect 3057 300 3092 334
rect 3126 300 3161 334
rect 3195 300 3230 334
rect 3264 300 3364 334
rect 264 220 3364 300
rect 3506 402 6606 482
rect 3506 368 3606 402
rect 3640 368 3675 402
rect 3709 368 3744 402
rect 3778 368 3813 402
rect 3847 368 3882 402
rect 3916 368 3951 402
rect 3985 368 4020 402
rect 4054 368 4089 402
rect 4123 368 4158 402
rect 4192 368 4227 402
rect 4261 368 4296 402
rect 3506 334 4296 368
rect 3506 300 3606 334
rect 3640 300 3675 334
rect 3709 300 3744 334
rect 3778 300 3813 334
rect 3847 300 3882 334
rect 3916 300 3951 334
rect 3985 300 4020 334
rect 4054 300 4089 334
rect 4123 300 4158 334
rect 4192 300 4227 334
rect 4261 300 4296 334
rect 6506 300 6606 402
rect 3506 220 6606 300
rect 6748 402 9848 482
rect 6748 300 6848 402
rect 9058 368 9093 402
rect 9127 368 9162 402
rect 9196 368 9231 402
rect 9265 368 9300 402
rect 9334 368 9369 402
rect 9403 368 9438 402
rect 9472 368 9507 402
rect 9541 368 9576 402
rect 9610 368 9645 402
rect 9679 368 9714 402
rect 9748 368 9848 402
rect 9058 334 9848 368
rect 9058 300 9093 334
rect 9127 300 9162 334
rect 9196 300 9231 334
rect 9265 300 9300 334
rect 9334 300 9369 334
rect 9403 300 9438 334
rect 9472 300 9507 334
rect 9541 300 9576 334
rect 9610 300 9645 334
rect 9679 300 9714 334
rect 9748 300 9848 334
rect 6748 220 9848 300
rect 9990 402 13090 482
rect 9990 368 10090 402
rect 10124 368 10159 402
rect 10193 368 10228 402
rect 10262 368 10297 402
rect 10331 368 10366 402
rect 10400 368 10435 402
rect 10469 368 10504 402
rect 10538 368 10573 402
rect 10607 368 10642 402
rect 10676 368 10711 402
rect 10745 368 10780 402
rect 9990 334 10780 368
rect 9990 300 10090 334
rect 10124 300 10159 334
rect 10193 300 10228 334
rect 10262 300 10297 334
rect 10331 300 10366 334
rect 10400 300 10435 334
rect 10469 300 10504 334
rect 10538 300 10573 334
rect 10607 300 10642 334
rect 10676 300 10711 334
rect 10745 300 10780 334
rect 12990 300 13090 402
rect 9990 220 13090 300
rect 13232 402 16332 482
rect 13232 300 13332 402
rect 15542 368 15577 402
rect 15611 368 15646 402
rect 15680 368 15715 402
rect 15749 368 15784 402
rect 15818 368 15853 402
rect 15887 368 15922 402
rect 15956 368 15991 402
rect 16025 368 16060 402
rect 16094 368 16129 402
rect 16163 368 16198 402
rect 16232 368 16332 402
rect 15542 334 16332 368
rect 15542 300 15577 334
rect 15611 300 15646 334
rect 15680 300 15715 334
rect 15749 300 15784 334
rect 15818 300 15853 334
rect 15887 300 15922 334
rect 15956 300 15991 334
rect 16025 300 16060 334
rect 16094 300 16129 334
rect 16163 300 16198 334
rect 16232 300 16332 334
tri 264 200 284 220 ne
rect 284 200 3344 220
tri 3344 200 3364 220 nw
tri 3506 200 3526 220 ne
rect 3526 200 6586 220
tri 6586 200 6606 220 nw
tri 264 70 284 90 se
rect 284 70 3344 90
tri 3344 70 3364 90 sw
tri 3506 70 3526 90 se
rect 3526 70 6586 90
tri 6586 70 6606 90 sw
tri 6748 200 6768 220 ne
rect 6768 200 9828 220
tri 9828 200 9848 220 nw
tri 9990 200 10010 220 ne
rect 10010 200 13070 220
tri 13070 200 13090 220 nw
tri 6748 70 6768 90 se
rect 6768 70 9828 90
tri 9828 70 9848 90 sw
tri 9990 70 10010 90 se
rect 10010 70 13070 90
tri 13070 70 13090 90 sw
rect 264 -10 3364 70
rect 264 -112 364 -10
rect 2574 -44 2609 -10
rect 2643 -44 2678 -10
rect 2712 -44 2747 -10
rect 2781 -44 2816 -10
rect 2850 -44 2885 -10
rect 2919 -44 2954 -10
rect 2988 -44 3023 -10
rect 3057 -44 3092 -10
rect 3126 -44 3161 -10
rect 3195 -44 3230 -10
rect 3264 -44 3364 -10
rect 2574 -78 3364 -44
rect 2574 -112 2609 -78
rect 2643 -112 2678 -78
rect 2712 -112 2747 -78
rect 2781 -112 2816 -78
rect 2850 -112 2885 -78
rect 2919 -112 2954 -78
rect 2988 -112 3023 -78
rect 3057 -112 3092 -78
rect 3126 -112 3161 -78
rect 3195 -112 3230 -78
rect 3264 -112 3364 -78
rect 264 -142 3364 -112
rect 3506 -10 6606 70
rect 3506 -44 3606 -10
rect 3640 -44 3675 -10
rect 3709 -44 3744 -10
rect 3778 -44 3813 -10
rect 3847 -44 3882 -10
rect 3916 -44 3951 -10
rect 3985 -44 4020 -10
rect 4054 -44 4089 -10
rect 4123 -44 4158 -10
rect 4192 -44 4227 -10
rect 4261 -44 4296 -10
rect 3506 -78 4296 -44
rect 3506 -112 3606 -78
rect 3640 -112 3675 -78
rect 3709 -112 3744 -78
rect 3778 -112 3813 -78
rect 3847 -112 3882 -78
rect 3916 -112 3951 -78
rect 3985 -112 4020 -78
rect 4054 -112 4089 -78
rect 4123 -112 4158 -78
rect 4192 -112 4227 -78
rect 4261 -112 4296 -78
rect 6506 -112 6606 -10
rect 3506 -142 6606 -112
rect 6748 -10 9848 70
rect 6748 -112 6848 -10
rect 9058 -44 9093 -10
rect 9127 -44 9162 -10
rect 9196 -44 9231 -10
rect 9265 -44 9300 -10
rect 9334 -44 9369 -10
rect 9403 -44 9438 -10
rect 9472 -44 9507 -10
rect 9541 -44 9576 -10
rect 9610 -44 9645 -10
rect 9679 -44 9714 -10
rect 9748 -44 9848 -10
rect 9058 -78 9848 -44
rect 9058 -112 9093 -78
rect 9127 -112 9162 -78
rect 9196 -112 9231 -78
rect 9265 -112 9300 -78
rect 9334 -112 9369 -78
rect 9403 -112 9438 -78
rect 9472 -112 9507 -78
rect 9541 -112 9576 -78
rect 9610 -112 9645 -78
rect 9679 -112 9714 -78
rect 9748 -112 9848 -78
rect 6748 -142 9848 -112
rect 9990 -10 13090 70
rect 13232 220 16332 300
rect 16474 402 19574 482
rect 16474 368 16574 402
rect 16608 368 16643 402
rect 16677 368 16712 402
rect 16746 368 16781 402
rect 16815 368 16850 402
rect 16884 368 16919 402
rect 16953 368 16988 402
rect 17022 368 17057 402
rect 17091 368 17126 402
rect 17160 368 17195 402
rect 17229 368 17264 402
rect 16474 334 17264 368
rect 16474 300 16574 334
rect 16608 300 16643 334
rect 16677 300 16712 334
rect 16746 300 16781 334
rect 16815 300 16850 334
rect 16884 300 16919 334
rect 16953 300 16988 334
rect 17022 300 17057 334
rect 17091 300 17126 334
rect 17160 300 17195 334
rect 17229 300 17264 334
rect 19474 300 19574 402
rect 16474 220 19574 300
tri 13232 200 13252 220 ne
rect 13252 200 16312 220
tri 16312 200 16332 220 nw
tri 16474 200 16494 220 ne
rect 16494 200 19554 220
tri 19554 200 19574 220 nw
tri 13232 70 13252 90 se
rect 13252 70 16312 90
tri 16312 70 16332 90 sw
tri 16474 70 16494 90 se
rect 16494 70 19554 90
tri 19554 70 19574 90 sw
rect 9990 -44 10090 -10
rect 10124 -44 10159 -10
rect 10193 -44 10228 -10
rect 10262 -44 10297 -10
rect 10331 -44 10366 -10
rect 10400 -44 10435 -10
rect 10469 -44 10504 -10
rect 10538 -44 10573 -10
rect 10607 -44 10642 -10
rect 10676 -44 10711 -10
rect 10745 -44 10780 -10
rect 9990 -78 10780 -44
rect 9990 -112 10090 -78
rect 10124 -112 10159 -78
rect 10193 -112 10228 -78
rect 10262 -112 10297 -78
rect 10331 -112 10366 -78
rect 10400 -112 10435 -78
rect 10469 -112 10504 -78
rect 10538 -112 10573 -78
rect 10607 -112 10642 -78
rect 10676 -112 10711 -78
rect 10745 -112 10780 -78
rect 12990 -112 13090 -10
rect 9990 -142 13090 -112
rect 13232 -10 16332 70
rect 13232 -112 13332 -10
rect 15542 -44 15577 -10
rect 15611 -44 15646 -10
rect 15680 -44 15715 -10
rect 15749 -44 15784 -10
rect 15818 -44 15853 -10
rect 15887 -44 15922 -10
rect 15956 -44 15991 -10
rect 16025 -44 16060 -10
rect 16094 -44 16129 -10
rect 16163 -44 16198 -10
rect 16232 -44 16332 -10
rect 15542 -78 16332 -44
rect 15542 -112 15577 -78
rect 15611 -112 15646 -78
rect 15680 -112 15715 -78
rect 15749 -112 15784 -78
rect 15818 -112 15853 -78
rect 15887 -112 15922 -78
rect 15956 -112 15991 -78
rect 16025 -112 16060 -78
rect 16094 -112 16129 -78
rect 16163 -112 16198 -78
rect 16232 -112 16332 -78
rect 13232 -142 16332 -112
rect 16474 -10 19574 70
rect 16474 -44 16574 -10
rect 16608 -44 16643 -10
rect 16677 -44 16712 -10
rect 16746 -44 16781 -10
rect 16815 -44 16850 -10
rect 16884 -44 16919 -10
rect 16953 -44 16988 -10
rect 17022 -44 17057 -10
rect 17091 -44 17126 -10
rect 17160 -44 17195 -10
rect 17229 -44 17264 -10
rect 16474 -78 17264 -44
rect 16474 -112 16574 -78
rect 16608 -112 16643 -78
rect 16677 -112 16712 -78
rect 16746 -112 16781 -78
rect 16815 -112 16850 -78
rect 16884 -112 16919 -78
rect 16953 -112 16988 -78
rect 17022 -112 17057 -78
rect 17091 -112 17126 -78
rect 17160 -112 17195 -78
rect 17229 -112 17264 -78
rect 19474 -112 19574 -10
rect 16474 -142 19574 -112
<< mvndiffc >>
rect -1597 12275 -1563 12309
rect -1597 12207 -1563 12241
rect -1597 12139 -1563 12173
rect -1597 12071 -1563 12105
rect -1597 12003 -1563 12037
rect -1597 11935 -1563 11969
rect -1597 11867 -1563 11901
rect -1597 11799 -1563 11833
rect -1441 12275 -1407 12309
rect -1441 12207 -1407 12241
rect -1441 12139 -1407 12173
rect -1441 12071 -1407 12105
rect -1441 12003 -1407 12037
rect -1441 11935 -1407 11969
rect -1441 11867 -1407 11901
rect -1441 11799 -1407 11833
rect -1285 12275 -1251 12309
rect -1285 12207 -1251 12241
rect -1285 12139 -1251 12173
rect -1285 12071 -1251 12105
rect -1285 12003 -1251 12037
rect -1285 11935 -1251 11969
rect -1285 11867 -1251 11901
rect -1285 11799 -1251 11833
rect -1597 11609 -1563 11643
rect -1597 11541 -1563 11575
rect -1597 11473 -1563 11507
rect -1597 11405 -1563 11439
rect -1597 11337 -1563 11371
rect -1597 11269 -1563 11303
rect -1597 11201 -1563 11235
rect -1597 11133 -1563 11167
rect -1441 11609 -1407 11643
rect -1441 11541 -1407 11575
rect -1441 11473 -1407 11507
rect -1441 11405 -1407 11439
rect -1441 11337 -1407 11371
rect -1441 11269 -1407 11303
rect -1441 11201 -1407 11235
rect -1441 11133 -1407 11167
rect -1285 11609 -1251 11643
rect -1285 11541 -1251 11575
rect -1285 11473 -1251 11507
rect -1285 11405 -1251 11439
rect -1285 11337 -1251 11371
rect -1285 11269 -1251 11303
rect -1285 11201 -1251 11235
rect -1285 11133 -1251 11167
rect -1597 10811 -1563 10845
rect -1597 10743 -1563 10777
rect -1597 10675 -1563 10709
rect -1597 10607 -1563 10641
rect -1597 10539 -1563 10573
rect -1597 10471 -1563 10505
rect -1597 10403 -1563 10437
rect -1597 10335 -1563 10369
rect -1441 10811 -1407 10845
rect -1441 10743 -1407 10777
rect -1441 10675 -1407 10709
rect -1441 10607 -1407 10641
rect -1441 10539 -1407 10573
rect -1441 10471 -1407 10505
rect -1441 10403 -1407 10437
rect -1441 10335 -1407 10369
rect -1285 10811 -1251 10845
rect -1285 10743 -1251 10777
rect -1285 10675 -1251 10709
rect -1285 10607 -1251 10641
rect -1285 10539 -1251 10573
rect -1285 10471 -1251 10505
rect -1285 10403 -1251 10437
rect -1285 10335 -1251 10369
<< mvpdiffc >>
rect -1641 2785 -1607 2819
rect -1641 2717 -1607 2751
rect -1641 2649 -1607 2683
rect -1641 2581 -1607 2615
rect -1641 2513 -1607 2547
rect -1641 2445 -1607 2479
rect -1641 2377 -1607 2411
rect -1641 2309 -1607 2343
rect -1485 2785 -1451 2819
rect -1485 2717 -1451 2751
rect -1485 2649 -1451 2683
rect -1485 2581 -1451 2615
rect -1485 2513 -1451 2547
rect -1485 2445 -1451 2479
rect -1485 2377 -1451 2411
rect -1485 2309 -1451 2343
rect -1329 2785 -1295 2819
rect -1329 2717 -1295 2751
rect -1329 2649 -1295 2683
rect -1329 2581 -1295 2615
rect -1329 2513 -1295 2547
rect -1329 2445 -1295 2479
rect -1329 2377 -1295 2411
rect -1329 2309 -1295 2343
rect -1198 2785 -1164 2819
rect -1198 2717 -1164 2751
rect -1198 2649 -1164 2683
rect -1198 2581 -1164 2615
rect -1198 2513 -1164 2547
rect -1198 2445 -1164 2479
rect -1198 2377 -1164 2411
rect -1198 2309 -1164 2343
rect -1042 2785 -1008 2819
rect -1042 2717 -1008 2751
rect -1042 2649 -1008 2683
rect -1042 2581 -1008 2615
rect -1042 2513 -1008 2547
rect -1042 2445 -1008 2479
rect -1042 2377 -1008 2411
rect -1042 2309 -1008 2343
rect -886 2785 -852 2819
rect -886 2717 -852 2751
rect -886 2649 -852 2683
rect -886 2581 -852 2615
rect -886 2513 -852 2547
rect -886 2445 -852 2479
rect -886 2377 -852 2411
rect -886 2309 -852 2343
rect -1641 1979 -1607 2013
rect -1641 1911 -1607 1945
rect -1641 1843 -1607 1877
rect -1641 1775 -1607 1809
rect -1641 1707 -1607 1741
rect -1641 1639 -1607 1673
rect -1641 1571 -1607 1605
rect -1641 1503 -1607 1537
rect -1485 1979 -1451 2013
rect -1485 1911 -1451 1945
rect -1485 1843 -1451 1877
rect -1485 1775 -1451 1809
rect -1485 1707 -1451 1741
rect -1485 1639 -1451 1673
rect -1485 1571 -1451 1605
rect -1485 1503 -1451 1537
rect -1329 1979 -1295 2013
rect -1329 1911 -1295 1945
rect -1329 1843 -1295 1877
rect -1329 1775 -1295 1809
rect -1329 1707 -1295 1741
rect -1329 1639 -1295 1673
rect -1329 1571 -1295 1605
rect -1329 1503 -1295 1537
rect 364 1536 2574 1638
rect 2609 1604 2643 1638
rect 2678 1604 2712 1638
rect 2747 1604 2781 1638
rect 2816 1604 2850 1638
rect 2885 1604 2919 1638
rect 2954 1604 2988 1638
rect 3023 1604 3057 1638
rect 3092 1604 3126 1638
rect 3161 1604 3195 1638
rect 3230 1604 3264 1638
rect 2609 1536 2643 1570
rect 2678 1536 2712 1570
rect 2747 1536 2781 1570
rect 2816 1536 2850 1570
rect 2885 1536 2919 1570
rect 2954 1536 2988 1570
rect 3023 1536 3057 1570
rect 3092 1536 3126 1570
rect 3161 1536 3195 1570
rect 3230 1536 3264 1570
rect 3606 1604 3640 1638
rect 3675 1604 3709 1638
rect 3744 1604 3778 1638
rect 3813 1604 3847 1638
rect 3882 1604 3916 1638
rect 3951 1604 3985 1638
rect 4020 1604 4054 1638
rect 4089 1604 4123 1638
rect 4158 1604 4192 1638
rect 4227 1604 4261 1638
rect 3606 1536 3640 1570
rect 3675 1536 3709 1570
rect 3744 1536 3778 1570
rect 3813 1536 3847 1570
rect 3882 1536 3916 1570
rect 3951 1536 3985 1570
rect 4020 1536 4054 1570
rect 4089 1536 4123 1570
rect 4158 1536 4192 1570
rect 4227 1536 4261 1570
rect 4296 1536 6506 1638
rect 6848 1536 9058 1638
rect 9093 1604 9127 1638
rect 9162 1604 9196 1638
rect 9231 1604 9265 1638
rect 9300 1604 9334 1638
rect 9369 1604 9403 1638
rect 9438 1604 9472 1638
rect 9507 1604 9541 1638
rect 9576 1604 9610 1638
rect 9645 1604 9679 1638
rect 9714 1604 9748 1638
rect 9093 1536 9127 1570
rect 9162 1536 9196 1570
rect 9231 1536 9265 1570
rect 9300 1536 9334 1570
rect 9369 1536 9403 1570
rect 9438 1536 9472 1570
rect 9507 1536 9541 1570
rect 9576 1536 9610 1570
rect 9645 1536 9679 1570
rect 9714 1536 9748 1570
rect 364 1124 2574 1226
rect 2609 1192 2643 1226
rect 2678 1192 2712 1226
rect 2747 1192 2781 1226
rect 2816 1192 2850 1226
rect 2885 1192 2919 1226
rect 2954 1192 2988 1226
rect 3023 1192 3057 1226
rect 3092 1192 3126 1226
rect 3161 1192 3195 1226
rect 3230 1192 3264 1226
rect 2609 1124 2643 1158
rect 2678 1124 2712 1158
rect 2747 1124 2781 1158
rect 2816 1124 2850 1158
rect 2885 1124 2919 1158
rect 2954 1124 2988 1158
rect 3023 1124 3057 1158
rect 3092 1124 3126 1158
rect 3161 1124 3195 1158
rect 3230 1124 3264 1158
rect 10090 1604 10124 1638
rect 10159 1604 10193 1638
rect 10228 1604 10262 1638
rect 10297 1604 10331 1638
rect 10366 1604 10400 1638
rect 10435 1604 10469 1638
rect 10504 1604 10538 1638
rect 10573 1604 10607 1638
rect 10642 1604 10676 1638
rect 10711 1604 10745 1638
rect 10090 1536 10124 1570
rect 10159 1536 10193 1570
rect 10228 1536 10262 1570
rect 10297 1536 10331 1570
rect 10366 1536 10400 1570
rect 10435 1536 10469 1570
rect 10504 1536 10538 1570
rect 10573 1536 10607 1570
rect 10642 1536 10676 1570
rect 10711 1536 10745 1570
rect 10780 1536 12990 1638
rect 13332 1536 15542 1638
rect 15577 1604 15611 1638
rect 15646 1604 15680 1638
rect 15715 1604 15749 1638
rect 15784 1604 15818 1638
rect 15853 1604 15887 1638
rect 15922 1604 15956 1638
rect 15991 1604 16025 1638
rect 16060 1604 16094 1638
rect 16129 1604 16163 1638
rect 16198 1604 16232 1638
rect 15577 1536 15611 1570
rect 15646 1536 15680 1570
rect 15715 1536 15749 1570
rect 15784 1536 15818 1570
rect 15853 1536 15887 1570
rect 15922 1536 15956 1570
rect 15991 1536 16025 1570
rect 16060 1536 16094 1570
rect 16129 1536 16163 1570
rect 16198 1536 16232 1570
rect 3606 1192 3640 1226
rect 3675 1192 3709 1226
rect 3744 1192 3778 1226
rect 3813 1192 3847 1226
rect 3882 1192 3916 1226
rect 3951 1192 3985 1226
rect 4020 1192 4054 1226
rect 4089 1192 4123 1226
rect 4158 1192 4192 1226
rect 4227 1192 4261 1226
rect 3606 1124 3640 1158
rect 3675 1124 3709 1158
rect 3744 1124 3778 1158
rect 3813 1124 3847 1158
rect 3882 1124 3916 1158
rect 3951 1124 3985 1158
rect 4020 1124 4054 1158
rect 4089 1124 4123 1158
rect 4158 1124 4192 1158
rect 4227 1124 4261 1158
rect 4296 1124 6506 1226
rect 6848 1124 9058 1226
rect 9093 1192 9127 1226
rect 9162 1192 9196 1226
rect 9231 1192 9265 1226
rect 9300 1192 9334 1226
rect 9369 1192 9403 1226
rect 9438 1192 9472 1226
rect 9507 1192 9541 1226
rect 9576 1192 9610 1226
rect 9645 1192 9679 1226
rect 9714 1192 9748 1226
rect 9093 1124 9127 1158
rect 9162 1124 9196 1158
rect 9231 1124 9265 1158
rect 9300 1124 9334 1158
rect 9369 1124 9403 1158
rect 9438 1124 9472 1158
rect 9507 1124 9541 1158
rect 9576 1124 9610 1158
rect 9645 1124 9679 1158
rect 9714 1124 9748 1158
rect 16574 1604 16608 1638
rect 16643 1604 16677 1638
rect 16712 1604 16746 1638
rect 16781 1604 16815 1638
rect 16850 1604 16884 1638
rect 16919 1604 16953 1638
rect 16988 1604 17022 1638
rect 17057 1604 17091 1638
rect 17126 1604 17160 1638
rect 17195 1604 17229 1638
rect 16574 1536 16608 1570
rect 16643 1536 16677 1570
rect 16712 1536 16746 1570
rect 16781 1536 16815 1570
rect 16850 1536 16884 1570
rect 16919 1536 16953 1570
rect 16988 1536 17022 1570
rect 17057 1536 17091 1570
rect 17126 1536 17160 1570
rect 17195 1536 17229 1570
rect 17264 1536 19474 1638
rect 10090 1192 10124 1226
rect 10159 1192 10193 1226
rect 10228 1192 10262 1226
rect 10297 1192 10331 1226
rect 10366 1192 10400 1226
rect 10435 1192 10469 1226
rect 10504 1192 10538 1226
rect 10573 1192 10607 1226
rect 10642 1192 10676 1226
rect 10711 1192 10745 1226
rect 10090 1124 10124 1158
rect 10159 1124 10193 1158
rect 10228 1124 10262 1158
rect 10297 1124 10331 1158
rect 10366 1124 10400 1158
rect 10435 1124 10469 1158
rect 10504 1124 10538 1158
rect 10573 1124 10607 1158
rect 10642 1124 10676 1158
rect 10711 1124 10745 1158
rect 10780 1124 12990 1226
rect 13332 1124 15542 1226
rect 15577 1192 15611 1226
rect 15646 1192 15680 1226
rect 15715 1192 15749 1226
rect 15784 1192 15818 1226
rect 15853 1192 15887 1226
rect 15922 1192 15956 1226
rect 15991 1192 16025 1226
rect 16060 1192 16094 1226
rect 16129 1192 16163 1226
rect 16198 1192 16232 1226
rect 15577 1124 15611 1158
rect 15646 1124 15680 1158
rect 15715 1124 15749 1158
rect 15784 1124 15818 1158
rect 15853 1124 15887 1158
rect 15922 1124 15956 1158
rect 15991 1124 16025 1158
rect 16060 1124 16094 1158
rect 16129 1124 16163 1158
rect 16198 1124 16232 1158
rect 16574 1192 16608 1226
rect 16643 1192 16677 1226
rect 16712 1192 16746 1226
rect 16781 1192 16815 1226
rect 16850 1192 16884 1226
rect 16919 1192 16953 1226
rect 16988 1192 17022 1226
rect 17057 1192 17091 1226
rect 17126 1192 17160 1226
rect 17195 1192 17229 1226
rect 16574 1124 16608 1158
rect 16643 1124 16677 1158
rect 16712 1124 16746 1158
rect 16781 1124 16815 1158
rect 16850 1124 16884 1158
rect 16919 1124 16953 1158
rect 16988 1124 17022 1158
rect 17057 1124 17091 1158
rect 17126 1124 17160 1158
rect 17195 1124 17229 1158
rect 17264 1124 19474 1226
rect 364 712 2574 814
rect 2609 780 2643 814
rect 2678 780 2712 814
rect 2747 780 2781 814
rect 2816 780 2850 814
rect 2885 780 2919 814
rect 2954 780 2988 814
rect 3023 780 3057 814
rect 3092 780 3126 814
rect 3161 780 3195 814
rect 3230 780 3264 814
rect 2609 712 2643 746
rect 2678 712 2712 746
rect 2747 712 2781 746
rect 2816 712 2850 746
rect 2885 712 2919 746
rect 2954 712 2988 746
rect 3023 712 3057 746
rect 3092 712 3126 746
rect 3161 712 3195 746
rect 3230 712 3264 746
rect 3606 780 3640 814
rect 3675 780 3709 814
rect 3744 780 3778 814
rect 3813 780 3847 814
rect 3882 780 3916 814
rect 3951 780 3985 814
rect 4020 780 4054 814
rect 4089 780 4123 814
rect 4158 780 4192 814
rect 4227 780 4261 814
rect 3606 712 3640 746
rect 3675 712 3709 746
rect 3744 712 3778 746
rect 3813 712 3847 746
rect 3882 712 3916 746
rect 3951 712 3985 746
rect 4020 712 4054 746
rect 4089 712 4123 746
rect 4158 712 4192 746
rect 4227 712 4261 746
rect 4296 712 6506 814
rect 6848 712 9058 814
rect 9093 780 9127 814
rect 9162 780 9196 814
rect 9231 780 9265 814
rect 9300 780 9334 814
rect 9369 780 9403 814
rect 9438 780 9472 814
rect 9507 780 9541 814
rect 9576 780 9610 814
rect 9645 780 9679 814
rect 9714 780 9748 814
rect 9093 712 9127 746
rect 9162 712 9196 746
rect 9231 712 9265 746
rect 9300 712 9334 746
rect 9369 712 9403 746
rect 9438 712 9472 746
rect 9507 712 9541 746
rect 9576 712 9610 746
rect 9645 712 9679 746
rect 9714 712 9748 746
rect 10090 780 10124 814
rect 10159 780 10193 814
rect 10228 780 10262 814
rect 10297 780 10331 814
rect 10366 780 10400 814
rect 10435 780 10469 814
rect 10504 780 10538 814
rect 10573 780 10607 814
rect 10642 780 10676 814
rect 10711 780 10745 814
rect 10090 712 10124 746
rect 10159 712 10193 746
rect 10228 712 10262 746
rect 10297 712 10331 746
rect 10366 712 10400 746
rect 10435 712 10469 746
rect 10504 712 10538 746
rect 10573 712 10607 746
rect 10642 712 10676 746
rect 10711 712 10745 746
rect 10780 712 12990 814
rect 13332 712 15542 814
rect 15577 780 15611 814
rect 15646 780 15680 814
rect 15715 780 15749 814
rect 15784 780 15818 814
rect 15853 780 15887 814
rect 15922 780 15956 814
rect 15991 780 16025 814
rect 16060 780 16094 814
rect 16129 780 16163 814
rect 16198 780 16232 814
rect 15577 712 15611 746
rect 15646 712 15680 746
rect 15715 712 15749 746
rect 15784 712 15818 746
rect 15853 712 15887 746
rect 15922 712 15956 746
rect 15991 712 16025 746
rect 16060 712 16094 746
rect 16129 712 16163 746
rect 16198 712 16232 746
rect 16574 780 16608 814
rect 16643 780 16677 814
rect 16712 780 16746 814
rect 16781 780 16815 814
rect 16850 780 16884 814
rect 16919 780 16953 814
rect 16988 780 17022 814
rect 17057 780 17091 814
rect 17126 780 17160 814
rect 17195 780 17229 814
rect 16574 712 16608 746
rect 16643 712 16677 746
rect 16712 712 16746 746
rect 16781 712 16815 746
rect 16850 712 16884 746
rect 16919 712 16953 746
rect 16988 712 17022 746
rect 17057 712 17091 746
rect 17126 712 17160 746
rect 17195 712 17229 746
rect 17264 712 19474 814
rect 364 300 2574 402
rect 2609 368 2643 402
rect 2678 368 2712 402
rect 2747 368 2781 402
rect 2816 368 2850 402
rect 2885 368 2919 402
rect 2954 368 2988 402
rect 3023 368 3057 402
rect 3092 368 3126 402
rect 3161 368 3195 402
rect 3230 368 3264 402
rect 2609 300 2643 334
rect 2678 300 2712 334
rect 2747 300 2781 334
rect 2816 300 2850 334
rect 2885 300 2919 334
rect 2954 300 2988 334
rect 3023 300 3057 334
rect 3092 300 3126 334
rect 3161 300 3195 334
rect 3230 300 3264 334
rect 3606 368 3640 402
rect 3675 368 3709 402
rect 3744 368 3778 402
rect 3813 368 3847 402
rect 3882 368 3916 402
rect 3951 368 3985 402
rect 4020 368 4054 402
rect 4089 368 4123 402
rect 4158 368 4192 402
rect 4227 368 4261 402
rect 3606 300 3640 334
rect 3675 300 3709 334
rect 3744 300 3778 334
rect 3813 300 3847 334
rect 3882 300 3916 334
rect 3951 300 3985 334
rect 4020 300 4054 334
rect 4089 300 4123 334
rect 4158 300 4192 334
rect 4227 300 4261 334
rect 4296 300 6506 402
rect 6848 300 9058 402
rect 9093 368 9127 402
rect 9162 368 9196 402
rect 9231 368 9265 402
rect 9300 368 9334 402
rect 9369 368 9403 402
rect 9438 368 9472 402
rect 9507 368 9541 402
rect 9576 368 9610 402
rect 9645 368 9679 402
rect 9714 368 9748 402
rect 9093 300 9127 334
rect 9162 300 9196 334
rect 9231 300 9265 334
rect 9300 300 9334 334
rect 9369 300 9403 334
rect 9438 300 9472 334
rect 9507 300 9541 334
rect 9576 300 9610 334
rect 9645 300 9679 334
rect 9714 300 9748 334
rect 10090 368 10124 402
rect 10159 368 10193 402
rect 10228 368 10262 402
rect 10297 368 10331 402
rect 10366 368 10400 402
rect 10435 368 10469 402
rect 10504 368 10538 402
rect 10573 368 10607 402
rect 10642 368 10676 402
rect 10711 368 10745 402
rect 10090 300 10124 334
rect 10159 300 10193 334
rect 10228 300 10262 334
rect 10297 300 10331 334
rect 10366 300 10400 334
rect 10435 300 10469 334
rect 10504 300 10538 334
rect 10573 300 10607 334
rect 10642 300 10676 334
rect 10711 300 10745 334
rect 10780 300 12990 402
rect 13332 300 15542 402
rect 15577 368 15611 402
rect 15646 368 15680 402
rect 15715 368 15749 402
rect 15784 368 15818 402
rect 15853 368 15887 402
rect 15922 368 15956 402
rect 15991 368 16025 402
rect 16060 368 16094 402
rect 16129 368 16163 402
rect 16198 368 16232 402
rect 15577 300 15611 334
rect 15646 300 15680 334
rect 15715 300 15749 334
rect 15784 300 15818 334
rect 15853 300 15887 334
rect 15922 300 15956 334
rect 15991 300 16025 334
rect 16060 300 16094 334
rect 16129 300 16163 334
rect 16198 300 16232 334
rect 364 -112 2574 -10
rect 2609 -44 2643 -10
rect 2678 -44 2712 -10
rect 2747 -44 2781 -10
rect 2816 -44 2850 -10
rect 2885 -44 2919 -10
rect 2954 -44 2988 -10
rect 3023 -44 3057 -10
rect 3092 -44 3126 -10
rect 3161 -44 3195 -10
rect 3230 -44 3264 -10
rect 2609 -112 2643 -78
rect 2678 -112 2712 -78
rect 2747 -112 2781 -78
rect 2816 -112 2850 -78
rect 2885 -112 2919 -78
rect 2954 -112 2988 -78
rect 3023 -112 3057 -78
rect 3092 -112 3126 -78
rect 3161 -112 3195 -78
rect 3230 -112 3264 -78
rect 3606 -44 3640 -10
rect 3675 -44 3709 -10
rect 3744 -44 3778 -10
rect 3813 -44 3847 -10
rect 3882 -44 3916 -10
rect 3951 -44 3985 -10
rect 4020 -44 4054 -10
rect 4089 -44 4123 -10
rect 4158 -44 4192 -10
rect 4227 -44 4261 -10
rect 3606 -112 3640 -78
rect 3675 -112 3709 -78
rect 3744 -112 3778 -78
rect 3813 -112 3847 -78
rect 3882 -112 3916 -78
rect 3951 -112 3985 -78
rect 4020 -112 4054 -78
rect 4089 -112 4123 -78
rect 4158 -112 4192 -78
rect 4227 -112 4261 -78
rect 4296 -112 6506 -10
rect 6848 -112 9058 -10
rect 9093 -44 9127 -10
rect 9162 -44 9196 -10
rect 9231 -44 9265 -10
rect 9300 -44 9334 -10
rect 9369 -44 9403 -10
rect 9438 -44 9472 -10
rect 9507 -44 9541 -10
rect 9576 -44 9610 -10
rect 9645 -44 9679 -10
rect 9714 -44 9748 -10
rect 9093 -112 9127 -78
rect 9162 -112 9196 -78
rect 9231 -112 9265 -78
rect 9300 -112 9334 -78
rect 9369 -112 9403 -78
rect 9438 -112 9472 -78
rect 9507 -112 9541 -78
rect 9576 -112 9610 -78
rect 9645 -112 9679 -78
rect 9714 -112 9748 -78
rect 16574 368 16608 402
rect 16643 368 16677 402
rect 16712 368 16746 402
rect 16781 368 16815 402
rect 16850 368 16884 402
rect 16919 368 16953 402
rect 16988 368 17022 402
rect 17057 368 17091 402
rect 17126 368 17160 402
rect 17195 368 17229 402
rect 16574 300 16608 334
rect 16643 300 16677 334
rect 16712 300 16746 334
rect 16781 300 16815 334
rect 16850 300 16884 334
rect 16919 300 16953 334
rect 16988 300 17022 334
rect 17057 300 17091 334
rect 17126 300 17160 334
rect 17195 300 17229 334
rect 17264 300 19474 402
rect 10090 -44 10124 -10
rect 10159 -44 10193 -10
rect 10228 -44 10262 -10
rect 10297 -44 10331 -10
rect 10366 -44 10400 -10
rect 10435 -44 10469 -10
rect 10504 -44 10538 -10
rect 10573 -44 10607 -10
rect 10642 -44 10676 -10
rect 10711 -44 10745 -10
rect 10090 -112 10124 -78
rect 10159 -112 10193 -78
rect 10228 -112 10262 -78
rect 10297 -112 10331 -78
rect 10366 -112 10400 -78
rect 10435 -112 10469 -78
rect 10504 -112 10538 -78
rect 10573 -112 10607 -78
rect 10642 -112 10676 -78
rect 10711 -112 10745 -78
rect 10780 -112 12990 -10
rect 13332 -112 15542 -10
rect 15577 -44 15611 -10
rect 15646 -44 15680 -10
rect 15715 -44 15749 -10
rect 15784 -44 15818 -10
rect 15853 -44 15887 -10
rect 15922 -44 15956 -10
rect 15991 -44 16025 -10
rect 16060 -44 16094 -10
rect 16129 -44 16163 -10
rect 16198 -44 16232 -10
rect 15577 -112 15611 -78
rect 15646 -112 15680 -78
rect 15715 -112 15749 -78
rect 15784 -112 15818 -78
rect 15853 -112 15887 -78
rect 15922 -112 15956 -78
rect 15991 -112 16025 -78
rect 16060 -112 16094 -78
rect 16129 -112 16163 -78
rect 16198 -112 16232 -78
rect 16574 -44 16608 -10
rect 16643 -44 16677 -10
rect 16712 -44 16746 -10
rect 16781 -44 16815 -10
rect 16850 -44 16884 -10
rect 16919 -44 16953 -10
rect 16988 -44 17022 -10
rect 17057 -44 17091 -10
rect 17126 -44 17160 -10
rect 17195 -44 17229 -10
rect 16574 -112 16608 -78
rect 16643 -112 16677 -78
rect 16712 -112 16746 -78
rect 16781 -112 16815 -78
rect 16850 -112 16884 -78
rect 16919 -112 16953 -78
rect 16988 -112 17022 -78
rect 17057 -112 17091 -78
rect 17126 -112 17160 -78
rect 17195 -112 17229 -78
rect 17264 -112 19474 -10
<< psubdiff >>
rect -1787 14161 -1711 14195
rect -1677 14161 -1571 14195
rect -1787 14127 -1571 14161
rect -1685 14093 -1571 14127
rect -1129 14114 -1061 14195
rect -1129 14093 -1095 14114
rect -1163 14080 -1095 14093
rect -1163 14046 -1061 14080
rect -1787 8007 -1685 8041
rect -1753 7994 -1685 8007
rect -1753 7973 -1719 7994
rect -1787 7892 -1719 7973
rect -1209 7960 -1163 7994
rect -1209 7926 -1061 7960
rect -1209 7892 -1175 7926
rect -1141 7892 -1061 7926
<< mvnsubdiff >>
rect -668 16925 -498 16959
rect -2109 14449 -2041 14517
rect -2075 14415 -2041 14449
rect -1599 14483 -1564 14517
rect -1530 14483 -1495 14517
rect -1461 14483 -1426 14517
rect -1392 14483 -1357 14517
rect -1323 14483 -1288 14517
rect -1254 14483 -1219 14517
rect -1185 14483 -1150 14517
rect -1116 14483 -1081 14517
rect -1047 14483 -1012 14517
rect -978 14483 -943 14517
rect -909 14483 -874 14517
rect -840 14483 -805 14517
rect -771 14483 -736 14517
rect -1599 14449 -736 14483
rect -1599 14415 -1564 14449
rect -1530 14415 -1495 14449
rect -1461 14415 -1426 14449
rect -1392 14415 -1357 14449
rect -1323 14415 -1288 14449
rect -1254 14415 -1219 14449
rect -1185 14415 -1150 14449
rect -1116 14415 -1081 14449
rect -1047 14415 -1012 14449
rect -978 14415 -943 14449
rect -909 14415 -874 14449
rect -840 14415 -805 14449
rect -771 14415 -736 14449
rect -2109 14380 -1973 14415
rect -2075 14346 -2041 14380
rect -2007 14347 -1973 14380
rect -1599 14381 -736 14415
rect -1599 14347 -1564 14381
rect -1530 14347 -1495 14381
rect -1461 14347 -1426 14381
rect -1392 14347 -1357 14381
rect -1323 14347 -1288 14381
rect -1254 14347 -1219 14381
rect -1185 14347 -1150 14381
rect -1116 14347 -1081 14381
rect -1047 14347 -1012 14381
rect -978 14347 -943 14381
rect -909 14347 -874 14381
rect -840 14347 -805 14381
rect -771 14347 -736 14381
rect -2007 14346 -1939 14347
rect -2109 14312 -1939 14346
rect -2109 14311 -1973 14312
rect -2075 14277 -2041 14311
rect -2007 14278 -1973 14311
rect -2007 14277 -1939 14278
rect -2109 14243 -1939 14277
rect -2109 14242 -1973 14243
rect -2075 14208 -2041 14242
rect -2007 14209 -1973 14242
rect -2007 14208 -1939 14209
rect -2109 14174 -1939 14208
rect -2109 14173 -1973 14174
rect -2075 14139 -2041 14173
rect -2007 14140 -1973 14173
rect -2007 14139 -1939 14140
rect -2109 14105 -1939 14139
rect -2109 14104 -1973 14105
rect -2075 14070 -2041 14104
rect -2007 14071 -1973 14104
rect -2007 14070 -1939 14071
rect -2109 14036 -1939 14070
rect -2109 14035 -1973 14036
rect -2075 14001 -2041 14035
rect -2007 14002 -1973 14035
rect -2007 14001 -1939 14002
rect -2109 13967 -1939 14001
rect -2109 13966 -1973 13967
rect -2075 13932 -2041 13966
rect -2007 13933 -1973 13966
rect -2007 13932 -1939 13933
rect -2109 13898 -1939 13932
rect -2109 13897 -1973 13898
rect -2075 13863 -2041 13897
rect -2007 13864 -1973 13897
rect -2007 13863 -1939 13864
rect -2109 13829 -1939 13863
rect -2109 13828 -1973 13829
rect -2075 13794 -2041 13828
rect -2007 13795 -1973 13828
rect -2007 13794 -1939 13795
rect -2109 13760 -1939 13794
rect -2109 13759 -1973 13760
rect -2075 13725 -2041 13759
rect -2007 13726 -1973 13759
rect -2007 13725 -1939 13726
rect -2109 13691 -1939 13725
rect -2109 13690 -1973 13691
rect -2075 13656 -2041 13690
rect -2007 13657 -1973 13690
rect -2007 13656 -1939 13657
rect -2109 13622 -1939 13656
rect -2109 13621 -1973 13622
rect -2075 13587 -2041 13621
rect -2007 13588 -1973 13621
rect -2007 13587 -1939 13588
rect -2109 13553 -1939 13587
rect -2109 13552 -1973 13553
rect -2075 13518 -2041 13552
rect -2007 13519 -1973 13552
rect -2007 13518 -1939 13519
rect -2109 13484 -1939 13518
rect -2109 13483 -1973 13484
rect -2075 13449 -2041 13483
rect -2007 13450 -1973 13483
rect -2007 13449 -1939 13450
rect -2109 13415 -1939 13449
rect -2109 13414 -1973 13415
rect -2075 13380 -2041 13414
rect -2007 13381 -1973 13414
rect -2007 13380 -1939 13381
rect -2109 13346 -1939 13380
rect -2109 13345 -1973 13346
rect -2075 13311 -2041 13345
rect -2007 13312 -1973 13345
rect -2007 13311 -1939 13312
rect -2109 13277 -1939 13311
rect -2109 13276 -1973 13277
rect -2075 13242 -2041 13276
rect -2007 13243 -1973 13276
rect -2007 13242 -1939 13243
rect -2109 13208 -1939 13242
rect -2109 13207 -1973 13208
rect -2075 13173 -2041 13207
rect -2007 13174 -1973 13207
rect -2007 13173 -1939 13174
rect -2109 13139 -1939 13173
rect -2109 13138 -1973 13139
rect -2075 13104 -2041 13138
rect -2007 13105 -1973 13138
rect -2007 13104 -1939 13105
rect -2109 13070 -1939 13104
rect -2109 13069 -1973 13070
rect -2075 13035 -2041 13069
rect -2007 13036 -1973 13069
rect -2007 13035 -1939 13036
rect -2109 13001 -1939 13035
rect -2109 13000 -1973 13001
rect -2075 12966 -2041 13000
rect -2007 12967 -1973 13000
rect -2007 12966 -1939 12967
rect -2109 12932 -1939 12966
rect -2109 12931 -1973 12932
rect -2075 12897 -2041 12931
rect -2007 12898 -1973 12931
rect -2007 12897 -1939 12898
rect -2109 12863 -1939 12897
rect -2109 12862 -1973 12863
rect -2075 12828 -2041 12862
rect -2007 12829 -1973 12862
rect -2007 12828 -1939 12829
rect -2109 12794 -1939 12828
rect -2109 12793 -1973 12794
rect -2075 12759 -2041 12793
rect -2007 12760 -1973 12793
rect -2007 12759 -1939 12760
rect -2109 12725 -1939 12759
rect -2109 12724 -1973 12725
rect -2075 12690 -2041 12724
rect -2007 12691 -1973 12724
rect -2007 12690 -1939 12691
rect -2109 12656 -1939 12690
rect -2109 12655 -1973 12656
rect -2075 12621 -2041 12655
rect -2007 12622 -1973 12655
rect -2007 12621 -1939 12622
rect -2109 12587 -1939 12621
rect -2109 12586 -1973 12587
rect -2075 12552 -2041 12586
rect -2007 12553 -1973 12586
rect -2007 12552 -1939 12553
rect -2109 12518 -1939 12552
rect -2109 12517 -1973 12518
rect -2075 12483 -2041 12517
rect -2007 12484 -1973 12517
rect -2007 12483 -1939 12484
rect -2109 12449 -1939 12483
rect -2109 12448 -1973 12449
rect -2075 12414 -2041 12448
rect -2007 12415 -1973 12448
rect -2007 12414 -1939 12415
rect -2109 12380 -1939 12414
rect -2109 12379 -1973 12380
rect -2075 12345 -2041 12379
rect -2007 12346 -1973 12379
rect -2007 12345 -1939 12346
rect -2109 12311 -1939 12345
rect -2109 12310 -1973 12311
rect -2075 12276 -2041 12310
rect -2007 12277 -1973 12310
rect -2007 12276 -1939 12277
rect -2109 12242 -1939 12276
rect -2109 12241 -1973 12242
rect -2075 12207 -2041 12241
rect -2007 12208 -1973 12241
rect -2007 12207 -1939 12208
rect -2109 12173 -1939 12207
rect -2109 12172 -1973 12173
rect -2075 12138 -2041 12172
rect -2007 12139 -1973 12172
rect -2007 12138 -1939 12139
rect -2109 12104 -1939 12138
rect -2109 12103 -1973 12104
rect -2075 12069 -2041 12103
rect -2007 12070 -1973 12103
rect -2007 12069 -1939 12070
rect -2109 12035 -1939 12069
rect -2109 12034 -1973 12035
rect -2075 12000 -2041 12034
rect -2007 12001 -1973 12034
rect -2007 12000 -1939 12001
rect -2109 11966 -1939 12000
rect -2109 11965 -1973 11966
rect -2075 11931 -2041 11965
rect -2007 11932 -1973 11965
rect -2007 11931 -1939 11932
rect -2109 11897 -1939 11931
rect -2109 11896 -1973 11897
rect -2075 11862 -2041 11896
rect -2007 11863 -1973 11896
rect -2007 11862 -1939 11863
rect -2109 11828 -1939 11862
rect -2109 11827 -1973 11828
rect -2075 11793 -2041 11827
rect -2007 11794 -1973 11827
rect -2007 11793 -1939 11794
rect -2109 11759 -1939 11793
rect -2109 11758 -1973 11759
rect -2075 11724 -2041 11758
rect -2007 11725 -1973 11758
rect -2007 11724 -1939 11725
rect -2109 11690 -1939 11724
rect -2109 11689 -1973 11690
rect -2075 11655 -2041 11689
rect -2007 11656 -1973 11689
rect -2007 11655 -1939 11656
rect -2109 11621 -1939 11655
rect -2109 11620 -1973 11621
rect -2075 11586 -2041 11620
rect -2007 11587 -1973 11620
rect -2007 11586 -1939 11587
rect -2109 11552 -1939 11586
rect -2109 11551 -1973 11552
rect -2075 11517 -2041 11551
rect -2007 11518 -1973 11551
rect -2007 11517 -1939 11518
rect -2109 11483 -1939 11517
rect -2109 11482 -1973 11483
rect -2075 11448 -2041 11482
rect -2007 11449 -1973 11482
rect -2007 11448 -1939 11449
rect -2109 11414 -1939 11448
rect -2109 11413 -1973 11414
rect -2075 11379 -2041 11413
rect -2007 11380 -1973 11413
rect -2007 11379 -1939 11380
rect -2109 11345 -1939 11379
rect -2109 11344 -1973 11345
rect -2075 11310 -2041 11344
rect -2007 11311 -1973 11344
rect -2007 11310 -1939 11311
rect -2109 11276 -1939 11310
rect -2109 11275 -1973 11276
rect -2075 11241 -2041 11275
rect -2007 11242 -1973 11275
rect -2007 11241 -1939 11242
rect -2109 11207 -1939 11241
rect -2109 11206 -1973 11207
rect -2075 11172 -2041 11206
rect -2007 11173 -1973 11206
rect -2007 11172 -1939 11173
rect -2109 11138 -1939 11172
rect -2109 11137 -1973 11138
rect -2075 11103 -2041 11137
rect -2007 11104 -1973 11137
rect -2007 11103 -1939 11104
rect -2109 11069 -1939 11103
rect -2109 11068 -1973 11069
rect -2075 11034 -2041 11068
rect -2007 11035 -1973 11068
rect -2007 11034 -1939 11035
rect -2109 11000 -1939 11034
rect -2109 10999 -1973 11000
rect -2075 10965 -2041 10999
rect -2007 10966 -1973 10999
rect -2007 10965 -1939 10966
rect -2109 10931 -1939 10965
rect -2109 10930 -1973 10931
rect -2075 10896 -2041 10930
rect -2007 10897 -1973 10930
rect -2007 10896 -1939 10897
rect -2109 10862 -1939 10896
rect -2109 10861 -1973 10862
rect -2075 10827 -2041 10861
rect -2007 10828 -1973 10861
rect -2007 10827 -1939 10828
rect -2109 10793 -1939 10827
rect -2109 10792 -1973 10793
rect -2075 10758 -2041 10792
rect -2007 10759 -1973 10792
rect -2007 10758 -1939 10759
rect -2109 10724 -1939 10758
rect -2109 10723 -1973 10724
rect -2075 10689 -2041 10723
rect -2007 10690 -1973 10723
rect -2007 10689 -1939 10690
rect -2109 10655 -1939 10689
rect -2109 10654 -1973 10655
rect -2075 10620 -2041 10654
rect -2007 10621 -1973 10654
rect -2007 10620 -1939 10621
rect -2109 10586 -1939 10620
rect -2109 10585 -1973 10586
rect -2075 10551 -2041 10585
rect -2007 10552 -1973 10585
rect -2007 10551 -1939 10552
rect -2109 10517 -1939 10551
rect -2109 10516 -1973 10517
rect -2075 10482 -2041 10516
rect -2007 10483 -1973 10516
rect -2007 10482 -1939 10483
rect -2109 10448 -1939 10482
rect -2109 10447 -1973 10448
rect -2075 10413 -2041 10447
rect -2007 10414 -1973 10447
rect -2007 10413 -1939 10414
rect -2109 10379 -1939 10413
rect -2109 10378 -1973 10379
rect -2075 10344 -2041 10378
rect -2007 10345 -1973 10378
rect -2007 10344 -1939 10345
rect -2109 10310 -1939 10344
rect -2109 10309 -1973 10310
rect -2075 10275 -2041 10309
rect -2007 10276 -1973 10309
rect -2007 10275 -1939 10276
rect -2109 10241 -1939 10275
rect -2109 10240 -1973 10241
rect -2075 10206 -2041 10240
rect -2007 10207 -1973 10240
rect -2007 10206 -1939 10207
rect -2109 10172 -1939 10206
rect -2109 10171 -1973 10172
rect -2075 10137 -2041 10171
rect -2007 10138 -1973 10171
rect -2007 10137 -1939 10138
rect -2109 10103 -1939 10137
rect -2109 10102 -1973 10103
rect -2075 10068 -2041 10102
rect -2007 10069 -1973 10102
rect -2007 10068 -1939 10069
rect -2109 10034 -1939 10068
rect -2109 10033 -1973 10034
rect -2075 9999 -2041 10033
rect -2007 10000 -1973 10033
rect -2007 9999 -1939 10000
rect -2109 9965 -1939 9999
rect -2109 9964 -1973 9965
rect -2075 9930 -2041 9964
rect -2007 9931 -1973 9964
rect -2007 9930 -1939 9931
rect -2109 9896 -1939 9930
rect -2109 9895 -1973 9896
rect -2007 9862 -1973 9895
rect -2007 9827 -1939 9862
rect -668 7948 -498 7983
rect -634 7914 -600 7948
rect -566 7914 -532 7948
rect -668 7879 -498 7914
rect -634 7845 -600 7879
rect -566 7845 -532 7879
rect -668 7810 -498 7845
rect -634 7776 -600 7810
rect -566 7776 -532 7810
rect -668 7741 -498 7776
rect -1939 7685 -1904 7719
rect -1870 7685 -1835 7719
rect -1801 7685 -1766 7719
rect -1732 7685 -1697 7719
rect -1663 7685 -1628 7719
rect -1594 7685 -1559 7719
rect -1525 7685 -1490 7719
rect -1456 7685 -1421 7719
rect -1387 7685 -1352 7719
rect -1318 7685 -1283 7719
rect -1249 7685 -1214 7719
rect -1180 7685 -1145 7719
rect -1111 7685 -1076 7719
rect -2007 7651 -1076 7685
rect -702 7707 -668 7719
rect -634 7707 -600 7741
rect -566 7707 -532 7741
rect -702 7672 -498 7707
rect -2007 7617 -1972 7651
rect -1938 7617 -1903 7651
rect -1869 7617 -1834 7651
rect -1800 7617 -1765 7651
rect -1731 7617 -1696 7651
rect -1662 7617 -1627 7651
rect -1593 7617 -1558 7651
rect -1524 7617 -1489 7651
rect -1455 7617 -1420 7651
rect -1386 7617 -1351 7651
rect -1317 7617 -1282 7651
rect -1248 7617 -1213 7651
rect -1179 7617 -1144 7651
rect -2109 7583 -1144 7617
rect -2109 7549 -2041 7583
rect -2007 7549 -1972 7583
rect -1938 7549 -1903 7583
rect -1869 7549 -1834 7583
rect -1800 7549 -1765 7583
rect -1731 7549 -1696 7583
rect -1662 7549 -1627 7583
rect -1593 7549 -1558 7583
rect -1524 7549 -1489 7583
rect -1455 7549 -1420 7583
rect -1386 7549 -1351 7583
rect -1317 7549 -1282 7583
rect -1248 7549 -1213 7583
rect -1179 7549 -1144 7583
rect -702 7638 -668 7672
rect -634 7638 -600 7672
rect -566 7638 -532 7672
rect -702 7603 -498 7638
rect -702 7569 -668 7603
rect -634 7569 -600 7603
rect -566 7569 -532 7603
rect -702 7549 -498 7569
rect -668 7534 -498 7549
rect -634 7500 -600 7534
rect -566 7500 -532 7534
rect -668 7465 -498 7500
rect -634 7431 -600 7465
rect -566 7431 -532 7465
rect -668 7396 -498 7431
rect -634 7362 -600 7396
rect -566 7362 -532 7396
rect -668 7327 -498 7362
rect -634 7293 -600 7327
rect -566 7293 -532 7327
rect -668 7258 -498 7293
rect -634 7224 -600 7258
rect -566 7224 -532 7258
rect -668 7189 -498 7224
rect -634 7155 -600 7189
rect -566 7155 -532 7189
rect -668 7121 -498 7155
rect -52 2808 48 2978
rect 19938 2808 19972 2978
rect -52 2774 82 2808
rect -52 2740 -2 2774
rect 32 2740 82 2774
rect -52 2705 82 2740
rect -52 2671 -2 2705
rect 32 2671 82 2705
rect -52 2636 82 2671
rect -52 2602 -2 2636
rect 32 2602 82 2636
rect -52 2567 82 2602
rect -52 2533 -2 2567
rect 32 2533 82 2567
rect -52 2498 82 2533
rect -52 2464 -2 2498
rect 32 2464 82 2498
rect -52 2429 82 2464
rect -52 2395 -2 2429
rect 32 2395 82 2429
rect -52 2360 82 2395
rect -52 2326 -2 2360
rect 32 2326 82 2360
rect -52 2291 82 2326
rect -52 2257 -2 2291
rect 32 2257 82 2291
rect -52 2222 82 2257
rect -52 2188 -2 2222
rect 32 2188 82 2222
rect -52 2153 82 2188
rect -52 2119 -2 2153
rect 32 2119 82 2153
rect -52 2084 82 2119
rect -52 2050 -2 2084
rect 32 2050 82 2084
rect -52 2015 82 2050
rect -52 1981 -2 2015
rect 32 1981 82 2015
rect -52 1946 82 1981
rect -52 1912 -2 1946
rect 32 1912 82 1946
rect -52 1877 82 1912
rect -52 1843 -2 1877
rect 32 1843 82 1877
rect -52 1808 82 1843
rect -52 1774 -2 1808
rect 32 1774 82 1808
rect -52 1739 82 1774
rect -52 1705 -2 1739
rect 32 1705 82 1739
rect -52 1670 82 1705
rect -52 1636 -2 1670
rect 32 1636 82 1670
rect 19838 2558 19972 2592
rect 19838 2524 19888 2558
rect 19922 2524 19972 2558
rect 19838 2489 19972 2524
rect 19838 2455 19888 2489
rect 19922 2455 19972 2489
rect 19838 2420 19972 2455
rect 19838 2386 19888 2420
rect 19922 2386 19972 2420
rect 19838 2351 19972 2386
rect 19838 2317 19888 2351
rect 19922 2317 19972 2351
rect 19838 2282 19972 2317
rect 19838 2248 19888 2282
rect 19922 2248 19972 2282
rect 19838 2213 19972 2248
rect 19838 2179 19888 2213
rect 19922 2179 19972 2213
rect 19838 2144 19972 2179
rect 19838 2110 19888 2144
rect 19922 2110 19972 2144
rect 19838 2075 19972 2110
rect 19838 2041 19888 2075
rect 19922 2041 19972 2075
rect 19838 2006 19972 2041
rect 19838 1972 19888 2006
rect 19922 1972 19972 2006
rect 19838 1937 19972 1972
rect 19838 1903 19888 1937
rect 19922 1903 19972 1937
rect 19838 1868 19972 1903
rect 19838 1834 19888 1868
rect 19922 1834 19972 1868
rect 19838 1799 19972 1834
rect 19838 1765 19888 1799
rect 19922 1765 19972 1799
rect 19838 1730 19972 1765
rect 19838 1696 19888 1730
rect 19922 1696 19972 1730
rect -52 1601 82 1636
rect -52 1567 -2 1601
rect 32 1567 82 1601
rect -52 1532 82 1567
rect -52 1498 -2 1532
rect 32 1498 82 1532
rect -52 1463 82 1498
rect -52 1429 -2 1463
rect 32 1429 82 1463
rect -52 1393 82 1429
rect -52 1359 -2 1393
rect 32 1359 82 1393
rect -52 1323 82 1359
rect -52 1289 -2 1323
rect 32 1289 82 1323
rect -52 1253 82 1289
rect -52 1219 -2 1253
rect 32 1219 82 1253
rect -52 1183 82 1219
rect -52 1149 -2 1183
rect 32 1149 82 1183
rect -52 1113 82 1149
rect -52 1079 -2 1113
rect 32 1079 82 1113
rect -52 1043 82 1079
rect -52 1009 -2 1043
rect 32 1009 82 1043
rect -52 973 82 1009
rect -52 939 -2 973
rect 32 939 82 973
rect -52 903 82 939
rect -52 869 -2 903
rect 32 869 82 903
rect 19838 1661 19972 1696
rect 19838 1627 19888 1661
rect 19922 1627 19972 1661
rect 19838 1592 19972 1627
rect 19838 1558 19888 1592
rect 19922 1558 19972 1592
rect 19838 1523 19972 1558
rect 19838 1489 19888 1523
rect 19922 1489 19972 1523
rect 19838 1454 19972 1489
rect 19838 1420 19888 1454
rect 19922 1420 19972 1454
rect 19838 1385 19972 1420
rect 19838 1351 19888 1385
rect 19922 1351 19972 1385
rect 19838 1316 19972 1351
rect -52 833 82 869
rect -52 799 -2 833
rect 32 799 82 833
rect -52 763 82 799
rect -52 729 -2 763
rect 32 729 82 763
rect -52 693 82 729
rect -52 659 -2 693
rect 32 659 82 693
rect -52 623 82 659
rect -52 589 -2 623
rect 32 589 82 623
rect -52 553 82 589
rect -52 519 -2 553
rect 32 519 82 553
rect -52 483 82 519
rect -52 449 -2 483
rect 32 449 82 483
rect 19838 1282 19888 1316
rect 19922 1282 19972 1316
rect 19838 1247 19972 1282
rect 19838 1213 19888 1247
rect 19922 1213 19972 1247
rect 19838 1178 19972 1213
rect 19838 1144 19888 1178
rect 19922 1144 19972 1178
rect 19838 1109 19972 1144
rect 19838 1075 19888 1109
rect 19922 1075 19972 1109
rect 19838 1040 19972 1075
rect 19838 1006 19888 1040
rect 19922 1006 19972 1040
rect 19838 971 19972 1006
rect 19838 937 19888 971
rect 19922 937 19972 971
rect 19838 902 19972 937
rect 19838 868 19888 902
rect 19922 868 19972 902
rect 19838 833 19972 868
rect 19838 799 19888 833
rect 19922 799 19972 833
rect 19838 763 19972 799
rect 19838 729 19888 763
rect 19922 729 19972 763
rect 19838 693 19972 729
rect 19838 659 19888 693
rect 19922 659 19972 693
rect -52 413 82 449
rect -52 379 -2 413
rect 32 379 82 413
rect -52 343 82 379
rect -52 309 -2 343
rect 32 309 82 343
rect -52 273 82 309
rect -52 239 -2 273
rect 32 239 82 273
rect -52 203 82 239
rect -52 169 -2 203
rect 32 169 82 203
rect -52 133 82 169
rect -52 99 -2 133
rect 32 99 82 133
rect -52 63 82 99
rect -52 29 -2 63
rect 32 29 82 63
rect -52 -7 82 29
rect -52 -41 -2 -7
rect 32 -41 82 -7
rect -52 -77 82 -41
rect -52 -111 -2 -77
rect 32 -111 82 -77
rect -52 -147 82 -111
rect 19838 623 19972 659
rect 19838 589 19888 623
rect 19922 589 19972 623
rect 19838 553 19972 589
rect 19838 519 19888 553
rect 19922 519 19972 553
rect 19838 483 19972 519
rect 19838 449 19888 483
rect 19922 449 19972 483
rect 19838 413 19972 449
rect 19838 379 19888 413
rect 19922 379 19972 413
rect 19838 343 19972 379
rect 19838 309 19888 343
rect 19922 309 19972 343
rect 19838 273 19972 309
rect 19838 239 19888 273
rect 19922 239 19972 273
rect 19838 203 19972 239
rect 19838 169 19888 203
rect 19922 169 19972 203
rect 19838 133 19972 169
rect 19838 99 19888 133
rect 19922 99 19972 133
rect 19838 63 19972 99
rect 19838 29 19888 63
rect 19922 29 19972 63
rect 19838 -7 19972 29
rect 19838 -41 19888 -7
rect 19922 -41 19972 -7
rect 19838 -77 19972 -41
rect 19838 -111 19888 -77
rect 19922 -111 19972 -77
rect -52 -181 -2 -147
rect 32 -181 82 -147
rect -52 -215 82 -181
rect 19838 -147 19972 -111
rect 19838 -181 19888 -147
rect 19922 -181 19972 -147
rect 19838 -215 19972 -181
rect -52 -238 19972 -215
rect -52 -272 48 -238
rect 82 -272 116 -238
rect 150 -272 184 -238
rect 218 -272 252 -238
rect 286 -272 320 -238
rect 354 -272 388 -238
rect 422 -272 456 -238
rect 490 -272 524 -238
rect 558 -272 592 -238
rect 626 -272 660 -238
rect 694 -272 728 -238
rect 762 -272 796 -238
rect 830 -272 864 -238
rect 898 -272 932 -238
rect 966 -272 1000 -238
rect 1034 -272 1068 -238
rect 1102 -272 1136 -238
rect 1170 -272 1204 -238
rect 1238 -272 1272 -238
rect 1306 -272 1340 -238
rect 1374 -272 1408 -238
rect 1442 -272 1476 -238
rect 1510 -272 1544 -238
rect 1578 -272 1612 -238
rect 1646 -272 1680 -238
rect 1714 -272 1748 -238
rect 1782 -272 1816 -238
rect 1850 -272 1884 -238
rect 1918 -272 1952 -238
rect 1986 -272 2020 -238
rect 2054 -272 2088 -238
rect 2122 -272 2156 -238
rect 2190 -272 2224 -238
rect 2258 -272 2292 -238
rect 2326 -272 2360 -238
rect 2394 -272 2428 -238
rect 2462 -272 2496 -238
rect 2530 -272 2564 -238
rect 2598 -272 2632 -238
rect 2666 -272 2700 -238
rect 2734 -272 2768 -238
rect 2802 -272 2836 -238
rect 2870 -272 2904 -238
rect 2938 -272 2972 -238
rect 3006 -272 3040 -238
rect 3074 -272 3108 -238
rect 3142 -272 3176 -238
rect 3210 -272 3244 -238
rect 3278 -272 3312 -238
rect 3346 -272 3380 -238
rect 3414 -272 3448 -238
rect 3482 -272 3516 -238
rect 3550 -272 3584 -238
rect 3618 -272 3652 -238
rect 3686 -272 3720 -238
rect 3754 -272 3788 -238
rect 3822 -272 3856 -238
rect 3890 -272 3924 -238
rect 3958 -272 3992 -238
rect 4026 -272 4060 -238
rect 4094 -272 4128 -238
rect 4162 -272 4196 -238
rect 4230 -272 4264 -238
rect 4298 -272 4332 -238
rect 4366 -272 4400 -238
rect 4434 -272 4468 -238
rect 4502 -272 4536 -238
rect 4570 -272 4604 -238
rect 4638 -272 4672 -238
rect 4706 -272 4740 -238
rect 4774 -272 4808 -238
rect 4842 -272 4876 -238
rect 4910 -272 4944 -238
rect 4978 -272 5012 -238
rect 5046 -272 5080 -238
rect 5114 -272 5148 -238
rect 5182 -272 5216 -238
rect 5250 -272 5284 -238
rect 5318 -272 5352 -238
rect 5386 -272 5420 -238
rect 5454 -272 5488 -238
rect 5522 -272 5556 -238
rect 5590 -272 5624 -238
rect 5658 -272 5692 -238
rect 5726 -272 5760 -238
rect 5794 -272 5828 -238
rect 5862 -272 5896 -238
rect 5930 -272 5964 -238
rect 5998 -272 6032 -238
rect 6066 -272 6100 -238
rect 6134 -272 6168 -238
rect 6202 -272 6236 -238
rect 6270 -272 6304 -238
rect 6338 -272 6372 -238
rect 6406 -272 6440 -238
rect 6474 -272 6508 -238
rect 6542 -272 6576 -238
rect 6610 -272 6644 -238
rect 6678 -272 6712 -238
rect 6746 -272 6780 -238
rect 6814 -272 6848 -238
rect 6882 -272 6916 -238
rect 6950 -272 6984 -238
rect 7018 -272 7052 -238
rect 7086 -272 7120 -238
rect 7154 -272 7188 -238
rect 7222 -272 7256 -238
rect 7290 -272 7324 -238
rect 7358 -272 7392 -238
rect 7426 -272 7460 -238
rect 7494 -272 7528 -238
rect 7562 -272 7596 -238
rect 7630 -272 7664 -238
rect 7698 -272 7732 -238
rect 7766 -272 7800 -238
rect 7834 -272 7868 -238
rect 7902 -272 7936 -238
rect 7970 -272 8004 -238
rect 8038 -272 8072 -238
rect 8106 -272 8140 -238
rect 8174 -272 8208 -238
rect 8242 -272 8276 -238
rect 8310 -272 8344 -238
rect 8378 -272 8412 -238
rect 8446 -272 8480 -238
rect 8514 -272 8548 -238
rect 8582 -272 8616 -238
rect 8650 -272 8684 -238
rect 8718 -272 8752 -238
rect 8786 -272 8820 -238
rect 8854 -272 8888 -238
rect 8922 -272 8956 -238
rect 8990 -272 9024 -238
rect 9058 -272 9092 -238
rect 9126 -272 9160 -238
rect 9194 -272 9228 -238
rect 9262 -272 9296 -238
rect 9330 -272 9364 -238
rect 9398 -272 9432 -238
rect 9466 -272 9500 -238
rect 9534 -272 9568 -238
rect 9602 -272 9636 -238
rect 9670 -272 9704 -238
rect 9738 -272 9772 -238
rect 9806 -272 9840 -238
rect 9874 -272 9908 -238
rect 9942 -272 9976 -238
rect 10010 -272 10044 -238
rect 10078 -272 10112 -238
rect 10146 -272 10180 -238
rect 10214 -272 10248 -238
rect 10282 -272 10316 -238
rect 10350 -272 10384 -238
rect 10418 -272 10452 -238
rect 10486 -272 10520 -238
rect 10554 -272 10588 -238
rect 10622 -272 10656 -238
rect 10690 -272 10724 -238
rect 10758 -272 10792 -238
rect 10826 -272 10860 -238
rect 10894 -272 10928 -238
rect 10962 -272 10996 -238
rect 11030 -272 11064 -238
rect 11098 -272 11132 -238
rect 11166 -272 11200 -238
rect 11234 -272 11268 -238
rect 11302 -272 11336 -238
rect 11370 -272 11404 -238
rect 11438 -272 11472 -238
rect 11506 -272 11540 -238
rect 11574 -272 11608 -238
rect 11642 -272 11676 -238
rect 11710 -272 11744 -238
rect 11778 -272 11812 -238
rect 11846 -272 11880 -238
rect 11914 -272 11948 -238
rect 11982 -272 12016 -238
rect 12050 -272 12084 -238
rect 12118 -272 12152 -238
rect 12186 -272 12220 -238
rect 12254 -272 12288 -238
rect 12322 -272 12356 -238
rect 12390 -272 12424 -238
rect 12458 -272 12492 -238
rect 12526 -272 12560 -238
rect 12594 -272 12628 -238
rect 12662 -272 12696 -238
rect 12730 -272 12764 -238
rect 12798 -272 12832 -238
rect 12866 -272 12900 -238
rect 12934 -272 12968 -238
rect 13002 -272 13036 -238
rect 13070 -272 13104 -238
rect 13138 -272 13172 -238
rect 13206 -272 13240 -238
rect 13274 -272 13308 -238
rect 13342 -272 13376 -238
rect 13410 -272 13444 -238
rect 13478 -272 13512 -238
rect 13546 -272 13580 -238
rect 13614 -272 13648 -238
rect 13682 -272 13716 -238
rect 13750 -272 13784 -238
rect 13818 -272 13852 -238
rect 13886 -272 13920 -238
rect 13954 -272 13988 -238
rect 14022 -272 14056 -238
rect 14090 -272 14124 -238
rect 14158 -272 14192 -238
rect 14226 -272 14260 -238
rect 14294 -272 14328 -238
rect 14362 -272 14396 -238
rect 14430 -272 14464 -238
rect 14498 -272 14532 -238
rect 14566 -272 14600 -238
rect 14634 -272 14668 -238
rect 14702 -272 14736 -238
rect 14770 -272 14804 -238
rect 14838 -272 14872 -238
rect 14906 -272 14940 -238
rect 14974 -272 15008 -238
rect 15042 -272 15076 -238
rect 15110 -272 15144 -238
rect 15178 -272 15212 -238
rect 15246 -272 15280 -238
rect 15314 -272 15348 -238
rect 15382 -272 15416 -238
rect 15450 -272 15484 -238
rect 15518 -272 15552 -238
rect 15586 -272 15620 -238
rect 15654 -272 15688 -238
rect 15722 -272 15756 -238
rect 15790 -272 15824 -238
rect 15858 -272 15892 -238
rect 15926 -272 15960 -238
rect 15994 -272 16028 -238
rect 16062 -272 16096 -238
rect 16130 -272 16164 -238
rect 16198 -272 16232 -238
rect 16266 -272 16300 -238
rect 16334 -272 16368 -238
rect 16402 -272 16436 -238
rect 16470 -272 16504 -238
rect 16538 -272 16572 -238
rect 16606 -272 16640 -238
rect 16674 -272 16708 -238
rect 16742 -272 16776 -238
rect 16810 -272 16844 -238
rect 16878 -272 16912 -238
rect 16946 -272 16980 -238
rect 17014 -272 17048 -238
rect 17082 -272 17116 -238
rect 17150 -272 17184 -238
rect 17218 -272 17252 -238
rect 17286 -272 17320 -238
rect 17354 -272 17388 -238
rect 17422 -272 17456 -238
rect 17490 -272 17524 -238
rect 17558 -272 17592 -238
rect 17626 -272 17660 -238
rect 17694 -272 17728 -238
rect 17762 -272 17796 -238
rect 17830 -272 17864 -238
rect 17898 -272 17932 -238
rect 17966 -272 18000 -238
rect 18034 -272 18068 -238
rect 18102 -272 18136 -238
rect 18170 -272 18204 -238
rect 18238 -272 18272 -238
rect 18306 -272 18340 -238
rect 18374 -272 18408 -238
rect 18442 -272 18476 -238
rect 18510 -272 18544 -238
rect 18578 -272 18612 -238
rect 18646 -272 18680 -238
rect 18714 -272 18748 -238
rect 18782 -272 18816 -238
rect 18850 -272 18884 -238
rect 18918 -272 18952 -238
rect 18986 -272 19020 -238
rect 19054 -272 19088 -238
rect 19122 -272 19156 -238
rect 19190 -272 19224 -238
rect 19258 -272 19292 -238
rect 19326 -272 19360 -238
rect 19394 -272 19428 -238
rect 19462 -272 19496 -238
rect 19530 -272 19564 -238
rect 19598 -272 19632 -238
rect 19666 -272 19700 -238
rect 19734 -272 19768 -238
rect 19802 -272 19836 -238
rect 19870 -272 19904 -238
rect 19938 -272 19972 -238
rect -52 -295 19972 -272
<< psubdiffcont >>
rect -1711 14161 -1677 14195
rect -1787 8041 -1685 14127
rect -1571 14093 -1129 14195
rect -1095 14080 -1061 14114
rect -1787 7973 -1753 8007
rect -1719 7892 -1209 7994
rect -1163 7960 -1061 14046
rect -1175 7892 -1141 7926
<< mvnsubdiffcont >>
rect -668 14517 -498 16925
rect -2109 14415 -2075 14449
rect -2041 14415 -1599 14517
rect -1564 14483 -1530 14517
rect -1495 14483 -1461 14517
rect -1426 14483 -1392 14517
rect -1357 14483 -1323 14517
rect -1288 14483 -1254 14517
rect -1219 14483 -1185 14517
rect -1150 14483 -1116 14517
rect -1081 14483 -1047 14517
rect -1012 14483 -978 14517
rect -943 14483 -909 14517
rect -874 14483 -840 14517
rect -805 14483 -771 14517
rect -1564 14415 -1530 14449
rect -1495 14415 -1461 14449
rect -1426 14415 -1392 14449
rect -1357 14415 -1323 14449
rect -1288 14415 -1254 14449
rect -1219 14415 -1185 14449
rect -1150 14415 -1116 14449
rect -1081 14415 -1047 14449
rect -1012 14415 -978 14449
rect -943 14415 -909 14449
rect -874 14415 -840 14449
rect -805 14415 -771 14449
rect -2109 14346 -2075 14380
rect -2041 14346 -2007 14380
rect -1973 14347 -1599 14415
rect -1564 14347 -1530 14381
rect -1495 14347 -1461 14381
rect -1426 14347 -1392 14381
rect -1357 14347 -1323 14381
rect -1288 14347 -1254 14381
rect -1219 14347 -1185 14381
rect -1150 14347 -1116 14381
rect -1081 14347 -1047 14381
rect -1012 14347 -978 14381
rect -943 14347 -909 14381
rect -874 14347 -840 14381
rect -805 14347 -771 14381
rect -736 14347 -498 14517
rect -2109 14277 -2075 14311
rect -2041 14277 -2007 14311
rect -1973 14278 -1939 14312
rect -2109 14208 -2075 14242
rect -2041 14208 -2007 14242
rect -1973 14209 -1939 14243
rect -2109 14139 -2075 14173
rect -2041 14139 -2007 14173
rect -1973 14140 -1939 14174
rect -2109 14070 -2075 14104
rect -2041 14070 -2007 14104
rect -1973 14071 -1939 14105
rect -2109 14001 -2075 14035
rect -2041 14001 -2007 14035
rect -1973 14002 -1939 14036
rect -2109 13932 -2075 13966
rect -2041 13932 -2007 13966
rect -1973 13933 -1939 13967
rect -2109 13863 -2075 13897
rect -2041 13863 -2007 13897
rect -1973 13864 -1939 13898
rect -2109 13794 -2075 13828
rect -2041 13794 -2007 13828
rect -1973 13795 -1939 13829
rect -2109 13725 -2075 13759
rect -2041 13725 -2007 13759
rect -1973 13726 -1939 13760
rect -2109 13656 -2075 13690
rect -2041 13656 -2007 13690
rect -1973 13657 -1939 13691
rect -2109 13587 -2075 13621
rect -2041 13587 -2007 13621
rect -1973 13588 -1939 13622
rect -2109 13518 -2075 13552
rect -2041 13518 -2007 13552
rect -1973 13519 -1939 13553
rect -2109 13449 -2075 13483
rect -2041 13449 -2007 13483
rect -1973 13450 -1939 13484
rect -2109 13380 -2075 13414
rect -2041 13380 -2007 13414
rect -1973 13381 -1939 13415
rect -2109 13311 -2075 13345
rect -2041 13311 -2007 13345
rect -1973 13312 -1939 13346
rect -2109 13242 -2075 13276
rect -2041 13242 -2007 13276
rect -1973 13243 -1939 13277
rect -2109 13173 -2075 13207
rect -2041 13173 -2007 13207
rect -1973 13174 -1939 13208
rect -2109 13104 -2075 13138
rect -2041 13104 -2007 13138
rect -1973 13105 -1939 13139
rect -2109 13035 -2075 13069
rect -2041 13035 -2007 13069
rect -1973 13036 -1939 13070
rect -2109 12966 -2075 13000
rect -2041 12966 -2007 13000
rect -1973 12967 -1939 13001
rect -2109 12897 -2075 12931
rect -2041 12897 -2007 12931
rect -1973 12898 -1939 12932
rect -2109 12828 -2075 12862
rect -2041 12828 -2007 12862
rect -1973 12829 -1939 12863
rect -2109 12759 -2075 12793
rect -2041 12759 -2007 12793
rect -1973 12760 -1939 12794
rect -2109 12690 -2075 12724
rect -2041 12690 -2007 12724
rect -1973 12691 -1939 12725
rect -2109 12621 -2075 12655
rect -2041 12621 -2007 12655
rect -1973 12622 -1939 12656
rect -2109 12552 -2075 12586
rect -2041 12552 -2007 12586
rect -1973 12553 -1939 12587
rect -2109 12483 -2075 12517
rect -2041 12483 -2007 12517
rect -1973 12484 -1939 12518
rect -2109 12414 -2075 12448
rect -2041 12414 -2007 12448
rect -1973 12415 -1939 12449
rect -2109 12345 -2075 12379
rect -2041 12345 -2007 12379
rect -1973 12346 -1939 12380
rect -2109 12276 -2075 12310
rect -2041 12276 -2007 12310
rect -1973 12277 -1939 12311
rect -2109 12207 -2075 12241
rect -2041 12207 -2007 12241
rect -1973 12208 -1939 12242
rect -2109 12138 -2075 12172
rect -2041 12138 -2007 12172
rect -1973 12139 -1939 12173
rect -2109 12069 -2075 12103
rect -2041 12069 -2007 12103
rect -1973 12070 -1939 12104
rect -2109 12000 -2075 12034
rect -2041 12000 -2007 12034
rect -1973 12001 -1939 12035
rect -2109 11931 -2075 11965
rect -2041 11931 -2007 11965
rect -1973 11932 -1939 11966
rect -2109 11862 -2075 11896
rect -2041 11862 -2007 11896
rect -1973 11863 -1939 11897
rect -2109 11793 -2075 11827
rect -2041 11793 -2007 11827
rect -1973 11794 -1939 11828
rect -2109 11724 -2075 11758
rect -2041 11724 -2007 11758
rect -1973 11725 -1939 11759
rect -2109 11655 -2075 11689
rect -2041 11655 -2007 11689
rect -1973 11656 -1939 11690
rect -2109 11586 -2075 11620
rect -2041 11586 -2007 11620
rect -1973 11587 -1939 11621
rect -2109 11517 -2075 11551
rect -2041 11517 -2007 11551
rect -1973 11518 -1939 11552
rect -2109 11448 -2075 11482
rect -2041 11448 -2007 11482
rect -1973 11449 -1939 11483
rect -2109 11379 -2075 11413
rect -2041 11379 -2007 11413
rect -1973 11380 -1939 11414
rect -2109 11310 -2075 11344
rect -2041 11310 -2007 11344
rect -1973 11311 -1939 11345
rect -2109 11241 -2075 11275
rect -2041 11241 -2007 11275
rect -1973 11242 -1939 11276
rect -2109 11172 -2075 11206
rect -2041 11172 -2007 11206
rect -1973 11173 -1939 11207
rect -2109 11103 -2075 11137
rect -2041 11103 -2007 11137
rect -1973 11104 -1939 11138
rect -2109 11034 -2075 11068
rect -2041 11034 -2007 11068
rect -1973 11035 -1939 11069
rect -2109 10965 -2075 10999
rect -2041 10965 -2007 10999
rect -1973 10966 -1939 11000
rect -2109 10896 -2075 10930
rect -2041 10896 -2007 10930
rect -1973 10897 -1939 10931
rect -2109 10827 -2075 10861
rect -2041 10827 -2007 10861
rect -1973 10828 -1939 10862
rect -2109 10758 -2075 10792
rect -2041 10758 -2007 10792
rect -1973 10759 -1939 10793
rect -2109 10689 -2075 10723
rect -2041 10689 -2007 10723
rect -1973 10690 -1939 10724
rect -2109 10620 -2075 10654
rect -2041 10620 -2007 10654
rect -1973 10621 -1939 10655
rect -2109 10551 -2075 10585
rect -2041 10551 -2007 10585
rect -1973 10552 -1939 10586
rect -2109 10482 -2075 10516
rect -2041 10482 -2007 10516
rect -1973 10483 -1939 10517
rect -2109 10413 -2075 10447
rect -2041 10413 -2007 10447
rect -1973 10414 -1939 10448
rect -2109 10344 -2075 10378
rect -2041 10344 -2007 10378
rect -1973 10345 -1939 10379
rect -2109 10275 -2075 10309
rect -2041 10275 -2007 10309
rect -1973 10276 -1939 10310
rect -2109 10206 -2075 10240
rect -2041 10206 -2007 10240
rect -1973 10207 -1939 10241
rect -2109 10137 -2075 10171
rect -2041 10137 -2007 10171
rect -1973 10138 -1939 10172
rect -2109 10068 -2075 10102
rect -2041 10068 -2007 10102
rect -1973 10069 -1939 10103
rect -2109 9999 -2075 10033
rect -2041 9999 -2007 10033
rect -1973 10000 -1939 10034
rect -2109 9930 -2075 9964
rect -2041 9930 -2007 9964
rect -1973 9931 -1939 9965
rect -2109 9827 -2007 9895
rect -1973 9862 -1939 9896
rect -2109 7685 -1939 9827
rect -668 7983 -498 14347
rect -668 7914 -634 7948
rect -600 7914 -566 7948
rect -532 7914 -498 7948
rect -668 7845 -634 7879
rect -600 7845 -566 7879
rect -532 7845 -498 7879
rect -668 7776 -634 7810
rect -600 7776 -566 7810
rect -532 7776 -498 7810
rect -1904 7685 -1870 7719
rect -1835 7685 -1801 7719
rect -1766 7685 -1732 7719
rect -1697 7685 -1663 7719
rect -1628 7685 -1594 7719
rect -1559 7685 -1525 7719
rect -1490 7685 -1456 7719
rect -1421 7685 -1387 7719
rect -1352 7685 -1318 7719
rect -1283 7685 -1249 7719
rect -1214 7685 -1180 7719
rect -1145 7685 -1111 7719
rect -2109 7617 -2007 7685
rect -1076 7651 -702 7719
rect -668 7707 -634 7741
rect -600 7707 -566 7741
rect -532 7707 -498 7741
rect -1972 7617 -1938 7651
rect -1903 7617 -1869 7651
rect -1834 7617 -1800 7651
rect -1765 7617 -1731 7651
rect -1696 7617 -1662 7651
rect -1627 7617 -1593 7651
rect -1558 7617 -1524 7651
rect -1489 7617 -1455 7651
rect -1420 7617 -1386 7651
rect -1351 7617 -1317 7651
rect -1282 7617 -1248 7651
rect -1213 7617 -1179 7651
rect -2041 7549 -2007 7583
rect -1972 7549 -1938 7583
rect -1903 7549 -1869 7583
rect -1834 7549 -1800 7583
rect -1765 7549 -1731 7583
rect -1696 7549 -1662 7583
rect -1627 7549 -1593 7583
rect -1558 7549 -1524 7583
rect -1489 7549 -1455 7583
rect -1420 7549 -1386 7583
rect -1351 7549 -1317 7583
rect -1282 7549 -1248 7583
rect -1213 7549 -1179 7583
rect -1144 7549 -702 7651
rect -668 7638 -634 7672
rect -600 7638 -566 7672
rect -532 7638 -498 7672
rect -668 7569 -634 7603
rect -600 7569 -566 7603
rect -532 7569 -498 7603
rect -668 7500 -634 7534
rect -600 7500 -566 7534
rect -532 7500 -498 7534
rect -668 7431 -634 7465
rect -600 7431 -566 7465
rect -532 7431 -498 7465
rect -668 7362 -634 7396
rect -600 7362 -566 7396
rect -532 7362 -498 7396
rect -668 7293 -634 7327
rect -600 7293 -566 7327
rect -532 7293 -498 7327
rect -668 7224 -634 7258
rect -600 7224 -566 7258
rect -532 7224 -498 7258
rect -668 7155 -634 7189
rect -600 7155 -566 7189
rect -532 7155 -498 7189
rect 48 2808 19938 2978
rect -2 2740 32 2774
rect -2 2671 32 2705
rect -2 2602 32 2636
rect -2 2533 32 2567
rect -2 2464 32 2498
rect -2 2395 32 2429
rect -2 2326 32 2360
rect -2 2257 32 2291
rect -2 2188 32 2222
rect -2 2119 32 2153
rect -2 2050 32 2084
rect -2 1981 32 2015
rect -2 1912 32 1946
rect -2 1843 32 1877
rect -2 1774 32 1808
rect -2 1705 32 1739
rect -2 1636 32 1670
rect 19888 2524 19922 2558
rect 19888 2455 19922 2489
rect 19888 2386 19922 2420
rect 19888 2317 19922 2351
rect 19888 2248 19922 2282
rect 19888 2179 19922 2213
rect 19888 2110 19922 2144
rect 19888 2041 19922 2075
rect 19888 1972 19922 2006
rect 19888 1903 19922 1937
rect 19888 1834 19922 1868
rect 19888 1765 19922 1799
rect 19888 1696 19922 1730
rect -2 1567 32 1601
rect -2 1498 32 1532
rect -2 1429 32 1463
rect -2 1359 32 1393
rect -2 1289 32 1323
rect -2 1219 32 1253
rect -2 1149 32 1183
rect -2 1079 32 1113
rect -2 1009 32 1043
rect -2 939 32 973
rect -2 869 32 903
rect 19888 1627 19922 1661
rect 19888 1558 19922 1592
rect 19888 1489 19922 1523
rect 19888 1420 19922 1454
rect 19888 1351 19922 1385
rect -2 799 32 833
rect -2 729 32 763
rect -2 659 32 693
rect -2 589 32 623
rect -2 519 32 553
rect -2 449 32 483
rect 19888 1282 19922 1316
rect 19888 1213 19922 1247
rect 19888 1144 19922 1178
rect 19888 1075 19922 1109
rect 19888 1006 19922 1040
rect 19888 937 19922 971
rect 19888 868 19922 902
rect 19888 799 19922 833
rect 19888 729 19922 763
rect 19888 659 19922 693
rect -2 379 32 413
rect -2 309 32 343
rect -2 239 32 273
rect -2 169 32 203
rect -2 99 32 133
rect -2 29 32 63
rect -2 -41 32 -7
rect -2 -111 32 -77
rect 19888 589 19922 623
rect 19888 519 19922 553
rect 19888 449 19922 483
rect 19888 379 19922 413
rect 19888 309 19922 343
rect 19888 239 19922 273
rect 19888 169 19922 203
rect 19888 99 19922 133
rect 19888 29 19922 63
rect 19888 -41 19922 -7
rect 19888 -111 19922 -77
rect -2 -181 32 -147
rect 19888 -181 19922 -147
rect 48 -272 82 -238
rect 116 -272 150 -238
rect 184 -272 218 -238
rect 252 -272 286 -238
rect 320 -272 354 -238
rect 388 -272 422 -238
rect 456 -272 490 -238
rect 524 -272 558 -238
rect 592 -272 626 -238
rect 660 -272 694 -238
rect 728 -272 762 -238
rect 796 -272 830 -238
rect 864 -272 898 -238
rect 932 -272 966 -238
rect 1000 -272 1034 -238
rect 1068 -272 1102 -238
rect 1136 -272 1170 -238
rect 1204 -272 1238 -238
rect 1272 -272 1306 -238
rect 1340 -272 1374 -238
rect 1408 -272 1442 -238
rect 1476 -272 1510 -238
rect 1544 -272 1578 -238
rect 1612 -272 1646 -238
rect 1680 -272 1714 -238
rect 1748 -272 1782 -238
rect 1816 -272 1850 -238
rect 1884 -272 1918 -238
rect 1952 -272 1986 -238
rect 2020 -272 2054 -238
rect 2088 -272 2122 -238
rect 2156 -272 2190 -238
rect 2224 -272 2258 -238
rect 2292 -272 2326 -238
rect 2360 -272 2394 -238
rect 2428 -272 2462 -238
rect 2496 -272 2530 -238
rect 2564 -272 2598 -238
rect 2632 -272 2666 -238
rect 2700 -272 2734 -238
rect 2768 -272 2802 -238
rect 2836 -272 2870 -238
rect 2904 -272 2938 -238
rect 2972 -272 3006 -238
rect 3040 -272 3074 -238
rect 3108 -272 3142 -238
rect 3176 -272 3210 -238
rect 3244 -272 3278 -238
rect 3312 -272 3346 -238
rect 3380 -272 3414 -238
rect 3448 -272 3482 -238
rect 3516 -272 3550 -238
rect 3584 -272 3618 -238
rect 3652 -272 3686 -238
rect 3720 -272 3754 -238
rect 3788 -272 3822 -238
rect 3856 -272 3890 -238
rect 3924 -272 3958 -238
rect 3992 -272 4026 -238
rect 4060 -272 4094 -238
rect 4128 -272 4162 -238
rect 4196 -272 4230 -238
rect 4264 -272 4298 -238
rect 4332 -272 4366 -238
rect 4400 -272 4434 -238
rect 4468 -272 4502 -238
rect 4536 -272 4570 -238
rect 4604 -272 4638 -238
rect 4672 -272 4706 -238
rect 4740 -272 4774 -238
rect 4808 -272 4842 -238
rect 4876 -272 4910 -238
rect 4944 -272 4978 -238
rect 5012 -272 5046 -238
rect 5080 -272 5114 -238
rect 5148 -272 5182 -238
rect 5216 -272 5250 -238
rect 5284 -272 5318 -238
rect 5352 -272 5386 -238
rect 5420 -272 5454 -238
rect 5488 -272 5522 -238
rect 5556 -272 5590 -238
rect 5624 -272 5658 -238
rect 5692 -272 5726 -238
rect 5760 -272 5794 -238
rect 5828 -272 5862 -238
rect 5896 -272 5930 -238
rect 5964 -272 5998 -238
rect 6032 -272 6066 -238
rect 6100 -272 6134 -238
rect 6168 -272 6202 -238
rect 6236 -272 6270 -238
rect 6304 -272 6338 -238
rect 6372 -272 6406 -238
rect 6440 -272 6474 -238
rect 6508 -272 6542 -238
rect 6576 -272 6610 -238
rect 6644 -272 6678 -238
rect 6712 -272 6746 -238
rect 6780 -272 6814 -238
rect 6848 -272 6882 -238
rect 6916 -272 6950 -238
rect 6984 -272 7018 -238
rect 7052 -272 7086 -238
rect 7120 -272 7154 -238
rect 7188 -272 7222 -238
rect 7256 -272 7290 -238
rect 7324 -272 7358 -238
rect 7392 -272 7426 -238
rect 7460 -272 7494 -238
rect 7528 -272 7562 -238
rect 7596 -272 7630 -238
rect 7664 -272 7698 -238
rect 7732 -272 7766 -238
rect 7800 -272 7834 -238
rect 7868 -272 7902 -238
rect 7936 -272 7970 -238
rect 8004 -272 8038 -238
rect 8072 -272 8106 -238
rect 8140 -272 8174 -238
rect 8208 -272 8242 -238
rect 8276 -272 8310 -238
rect 8344 -272 8378 -238
rect 8412 -272 8446 -238
rect 8480 -272 8514 -238
rect 8548 -272 8582 -238
rect 8616 -272 8650 -238
rect 8684 -272 8718 -238
rect 8752 -272 8786 -238
rect 8820 -272 8854 -238
rect 8888 -272 8922 -238
rect 8956 -272 8990 -238
rect 9024 -272 9058 -238
rect 9092 -272 9126 -238
rect 9160 -272 9194 -238
rect 9228 -272 9262 -238
rect 9296 -272 9330 -238
rect 9364 -272 9398 -238
rect 9432 -272 9466 -238
rect 9500 -272 9534 -238
rect 9568 -272 9602 -238
rect 9636 -272 9670 -238
rect 9704 -272 9738 -238
rect 9772 -272 9806 -238
rect 9840 -272 9874 -238
rect 9908 -272 9942 -238
rect 9976 -272 10010 -238
rect 10044 -272 10078 -238
rect 10112 -272 10146 -238
rect 10180 -272 10214 -238
rect 10248 -272 10282 -238
rect 10316 -272 10350 -238
rect 10384 -272 10418 -238
rect 10452 -272 10486 -238
rect 10520 -272 10554 -238
rect 10588 -272 10622 -238
rect 10656 -272 10690 -238
rect 10724 -272 10758 -238
rect 10792 -272 10826 -238
rect 10860 -272 10894 -238
rect 10928 -272 10962 -238
rect 10996 -272 11030 -238
rect 11064 -272 11098 -238
rect 11132 -272 11166 -238
rect 11200 -272 11234 -238
rect 11268 -272 11302 -238
rect 11336 -272 11370 -238
rect 11404 -272 11438 -238
rect 11472 -272 11506 -238
rect 11540 -272 11574 -238
rect 11608 -272 11642 -238
rect 11676 -272 11710 -238
rect 11744 -272 11778 -238
rect 11812 -272 11846 -238
rect 11880 -272 11914 -238
rect 11948 -272 11982 -238
rect 12016 -272 12050 -238
rect 12084 -272 12118 -238
rect 12152 -272 12186 -238
rect 12220 -272 12254 -238
rect 12288 -272 12322 -238
rect 12356 -272 12390 -238
rect 12424 -272 12458 -238
rect 12492 -272 12526 -238
rect 12560 -272 12594 -238
rect 12628 -272 12662 -238
rect 12696 -272 12730 -238
rect 12764 -272 12798 -238
rect 12832 -272 12866 -238
rect 12900 -272 12934 -238
rect 12968 -272 13002 -238
rect 13036 -272 13070 -238
rect 13104 -272 13138 -238
rect 13172 -272 13206 -238
rect 13240 -272 13274 -238
rect 13308 -272 13342 -238
rect 13376 -272 13410 -238
rect 13444 -272 13478 -238
rect 13512 -272 13546 -238
rect 13580 -272 13614 -238
rect 13648 -272 13682 -238
rect 13716 -272 13750 -238
rect 13784 -272 13818 -238
rect 13852 -272 13886 -238
rect 13920 -272 13954 -238
rect 13988 -272 14022 -238
rect 14056 -272 14090 -238
rect 14124 -272 14158 -238
rect 14192 -272 14226 -238
rect 14260 -272 14294 -238
rect 14328 -272 14362 -238
rect 14396 -272 14430 -238
rect 14464 -272 14498 -238
rect 14532 -272 14566 -238
rect 14600 -272 14634 -238
rect 14668 -272 14702 -238
rect 14736 -272 14770 -238
rect 14804 -272 14838 -238
rect 14872 -272 14906 -238
rect 14940 -272 14974 -238
rect 15008 -272 15042 -238
rect 15076 -272 15110 -238
rect 15144 -272 15178 -238
rect 15212 -272 15246 -238
rect 15280 -272 15314 -238
rect 15348 -272 15382 -238
rect 15416 -272 15450 -238
rect 15484 -272 15518 -238
rect 15552 -272 15586 -238
rect 15620 -272 15654 -238
rect 15688 -272 15722 -238
rect 15756 -272 15790 -238
rect 15824 -272 15858 -238
rect 15892 -272 15926 -238
rect 15960 -272 15994 -238
rect 16028 -272 16062 -238
rect 16096 -272 16130 -238
rect 16164 -272 16198 -238
rect 16232 -272 16266 -238
rect 16300 -272 16334 -238
rect 16368 -272 16402 -238
rect 16436 -272 16470 -238
rect 16504 -272 16538 -238
rect 16572 -272 16606 -238
rect 16640 -272 16674 -238
rect 16708 -272 16742 -238
rect 16776 -272 16810 -238
rect 16844 -272 16878 -238
rect 16912 -272 16946 -238
rect 16980 -272 17014 -238
rect 17048 -272 17082 -238
rect 17116 -272 17150 -238
rect 17184 -272 17218 -238
rect 17252 -272 17286 -238
rect 17320 -272 17354 -238
rect 17388 -272 17422 -238
rect 17456 -272 17490 -238
rect 17524 -272 17558 -238
rect 17592 -272 17626 -238
rect 17660 -272 17694 -238
rect 17728 -272 17762 -238
rect 17796 -272 17830 -238
rect 17864 -272 17898 -238
rect 17932 -272 17966 -238
rect 18000 -272 18034 -238
rect 18068 -272 18102 -238
rect 18136 -272 18170 -238
rect 18204 -272 18238 -238
rect 18272 -272 18306 -238
rect 18340 -272 18374 -238
rect 18408 -272 18442 -238
rect 18476 -272 18510 -238
rect 18544 -272 18578 -238
rect 18612 -272 18646 -238
rect 18680 -272 18714 -238
rect 18748 -272 18782 -238
rect 18816 -272 18850 -238
rect 18884 -272 18918 -238
rect 18952 -272 18986 -238
rect 19020 -272 19054 -238
rect 19088 -272 19122 -238
rect 19156 -272 19190 -238
rect 19224 -272 19258 -238
rect 19292 -272 19326 -238
rect 19360 -272 19394 -238
rect 19428 -272 19462 -238
rect 19496 -272 19530 -238
rect 19564 -272 19598 -238
rect 19632 -272 19666 -238
rect 19700 -272 19734 -238
rect 19768 -272 19802 -238
rect 19836 -272 19870 -238
rect 19904 -272 19938 -238
<< poly >>
rect -1552 12470 -1452 12493
rect -1552 12436 -1519 12470
rect -1485 12436 -1452 12470
rect -1552 12387 -1452 12436
rect -1396 12470 -1296 12493
rect -1396 12436 -1363 12470
rect -1329 12436 -1296 12470
rect -1396 12387 -1296 12436
rect -1552 11761 -1452 11787
rect -1396 11761 -1296 11787
rect -1552 11738 -1452 11755
rect -1552 11704 -1519 11738
rect -1485 11704 -1452 11738
rect -1552 11655 -1452 11704
rect -1396 11738 -1296 11755
rect -1396 11704 -1363 11738
rect -1329 11704 -1296 11738
rect -1396 11655 -1296 11704
rect -1552 11029 -1452 11055
rect -1396 11029 -1296 11055
rect -1552 11006 -1452 11023
rect -1552 10972 -1519 11006
rect -1485 10972 -1452 11006
rect -1552 10923 -1452 10972
rect -1396 11006 -1296 11023
rect -1396 10972 -1363 11006
rect -1329 10972 -1296 11006
rect -1396 10923 -1296 10972
rect -1552 10297 -1452 10323
rect -1396 10297 -1296 10323
rect 19638 6118 19756 6151
rect 19638 6084 19654 6118
rect 19688 6084 19722 6118
rect 19638 6051 19756 6084
rect 21796 6118 21914 6151
rect 21830 6084 21864 6118
rect 21898 6084 21914 6118
rect 21796 6051 21914 6084
rect 19647 5934 19715 5951
rect 21855 5934 21923 5951
rect 19647 5918 19781 5934
rect 19647 5884 19663 5918
rect 19697 5884 19731 5918
rect 19765 5884 19781 5918
rect 19647 5868 19781 5884
rect 21789 5918 21923 5934
rect 21789 5884 21805 5918
rect 21839 5884 21873 5918
rect 21907 5884 21923 5918
rect 21789 5868 21923 5884
rect 19647 5851 19715 5868
rect 21855 5851 21923 5868
rect 19638 5708 19706 5725
rect 21846 5708 21914 5725
rect 19638 5692 19772 5708
rect 19638 5658 19654 5692
rect 19688 5658 19722 5692
rect 19756 5658 19772 5692
rect 19638 5642 19772 5658
rect 21780 5692 21914 5708
rect 21780 5658 21796 5692
rect 21830 5658 21864 5692
rect 21898 5658 21914 5692
rect 21780 5642 21914 5658
rect 19638 5625 19706 5642
rect 21846 5625 21914 5642
rect 19681 5491 19799 5524
rect 19681 5457 19697 5491
rect 19731 5457 19765 5491
rect 19681 5424 19799 5457
rect 21839 5491 21957 5524
rect 21873 5457 21907 5491
rect 21941 5457 21957 5491
rect 21839 5424 21957 5457
rect -1596 2920 -1340 2943
rect -1596 2886 -1580 2920
rect -1546 2886 -1485 2920
rect -1451 2886 -1390 2920
rect -1356 2886 -1340 2920
rect -1596 2863 -1340 2886
rect -1596 2831 -1496 2863
rect -1440 2831 -1340 2863
rect -1153 2920 -897 2943
rect -1153 2886 -1137 2920
rect -1103 2886 -1042 2920
rect -1008 2886 -947 2920
rect -913 2886 -897 2920
rect -1153 2863 -897 2886
rect -1153 2831 -1053 2863
rect -997 2831 -897 2863
rect -1596 2199 -1496 2231
rect -1440 2199 -1340 2231
rect -1153 2199 -1053 2231
rect -997 2199 -897 2231
rect -1596 2114 -1340 2137
rect -1596 2080 -1580 2114
rect -1546 2080 -1485 2114
rect -1451 2080 -1390 2114
rect -1356 2080 -1340 2114
rect -1596 2057 -1340 2080
rect -1596 2025 -1496 2057
rect -1440 2025 -1340 2057
rect -1596 1393 -1496 1425
rect -1440 1393 -1340 1425
rect 166 1456 244 1476
tri 244 1456 264 1476 sw
tri 3364 1456 3384 1476 se
rect 3384 1456 3486 1476
tri 3486 1456 3506 1476 sw
tri 6606 1456 6626 1476 se
rect 6626 1456 6656 1476
rect 166 1432 264 1456
rect 166 1398 182 1432
rect 216 1398 264 1432
rect 166 1364 264 1398
rect 166 1330 182 1364
rect 216 1330 264 1364
rect 166 1306 264 1330
rect 3364 1432 3506 1456
rect 3364 1398 3423 1432
rect 3457 1398 3506 1432
rect 3364 1364 3506 1398
rect 3364 1330 3423 1364
rect 3457 1330 3506 1364
rect 3364 1306 3506 1330
rect 6606 1306 6656 1456
rect 166 1286 244 1306
tri 244 1286 264 1306 nw
tri 3364 1286 3384 1306 ne
rect 3384 1286 3486 1306
tri 3486 1286 3506 1306 nw
rect 166 1044 244 1064
tri 244 1044 264 1064 sw
tri 6606 1286 6626 1306 ne
rect 6626 1286 6656 1306
rect 6698 1456 6728 1476
tri 6728 1456 6748 1476 sw
tri 9848 1456 9868 1476 se
rect 9868 1456 9970 1476
tri 9970 1456 9990 1476 sw
tri 13090 1456 13110 1476 se
rect 13110 1456 13140 1476
rect 6698 1306 6748 1456
rect 9848 1432 9990 1456
rect 9848 1398 9907 1432
rect 9941 1398 9990 1432
rect 9848 1364 9990 1398
rect 9848 1330 9907 1364
rect 9941 1330 9990 1364
rect 9848 1306 9990 1330
rect 13090 1306 13140 1456
rect 6698 1286 6728 1306
tri 6728 1286 6748 1306 nw
tri 3364 1044 3384 1064 se
rect 3384 1044 3486 1064
tri 3486 1044 3506 1064 sw
tri 9848 1286 9868 1306 ne
rect 9868 1286 9970 1306
tri 9970 1286 9990 1306 nw
tri 6606 1044 6626 1064 se
rect 6626 1044 6728 1064
tri 6728 1044 6748 1064 sw
tri 13090 1286 13110 1306 ne
rect 13110 1286 13140 1306
rect 13182 1456 13212 1476
tri 13212 1456 13232 1476 sw
tri 16332 1456 16352 1476 se
rect 16352 1456 16454 1476
tri 16454 1456 16474 1476 sw
tri 19574 1456 19594 1476 se
rect 19594 1456 19672 1476
rect 13182 1306 13232 1456
rect 16332 1432 16474 1456
rect 16332 1398 16392 1432
rect 16426 1398 16474 1432
rect 16332 1364 16474 1398
rect 16332 1330 16392 1364
rect 16426 1330 16474 1364
rect 16332 1306 16474 1330
rect 19574 1432 19672 1456
rect 19574 1398 19622 1432
rect 19656 1398 19672 1432
rect 19574 1364 19672 1398
rect 19574 1330 19622 1364
rect 19656 1330 19672 1364
rect 19574 1306 19672 1330
rect 13182 1286 13212 1306
tri 13212 1286 13232 1306 nw
tri 9848 1044 9868 1064 se
rect 9868 1044 9970 1064
tri 9970 1044 9990 1064 sw
tri 16332 1286 16352 1306 ne
rect 16352 1286 16454 1306
tri 16454 1286 16474 1306 nw
tri 13090 1044 13110 1064 se
rect 13110 1044 13212 1064
tri 13212 1044 13232 1064 sw
tri 19574 1286 19594 1306 ne
rect 19594 1286 19672 1306
tri 16332 1044 16352 1064 se
rect 16352 1044 16382 1064
rect 166 1020 264 1044
rect 166 986 182 1020
rect 216 986 264 1020
rect 166 952 264 986
rect 166 918 182 952
rect 216 918 264 952
rect 166 894 264 918
rect 3364 1020 3506 1044
rect 3364 986 3423 1020
rect 3457 986 3506 1020
rect 3364 952 3506 986
rect 3364 918 3423 952
rect 3457 918 3506 952
rect 3364 894 3506 918
rect 6606 1020 6748 1044
rect 6606 986 6665 1020
rect 6699 986 6748 1020
rect 6606 952 6748 986
rect 6606 918 6665 952
rect 6699 918 6748 952
rect 6606 894 6748 918
rect 9848 1020 9990 1044
rect 9848 986 9907 1020
rect 9941 986 9990 1020
rect 9848 952 9990 986
rect 9848 918 9907 952
rect 9941 918 9990 952
rect 9848 894 9990 918
rect 13090 1020 13232 1044
rect 13090 986 13150 1020
rect 13184 986 13232 1020
rect 13090 952 13232 986
rect 13090 918 13150 952
rect 13184 918 13232 952
rect 13090 894 13232 918
rect 16332 894 16382 1044
rect 166 874 244 894
tri 244 874 264 894 nw
tri 3364 874 3384 894 ne
rect 3384 874 3486 894
tri 3486 874 3506 894 nw
rect 166 632 244 652
tri 244 632 264 652 sw
tri 6606 874 6626 894 ne
rect 6626 874 6728 894
tri 6728 874 6748 894 nw
tri 3364 632 3384 652 se
rect 3384 632 3486 652
tri 3486 632 3506 652 sw
tri 9848 874 9868 894 ne
rect 9868 874 9970 894
tri 9970 874 9990 894 nw
tri 6606 632 6626 652 se
rect 6626 632 6728 652
tri 6728 632 6748 652 sw
tri 13090 874 13110 894 ne
rect 13110 874 13212 894
tri 13212 874 13232 894 nw
tri 9848 632 9868 652 se
rect 9868 632 9970 652
tri 9970 632 9990 652 sw
tri 16332 874 16352 894 ne
rect 16352 874 16382 894
rect 16424 1044 16454 1064
tri 16454 1044 16474 1064 sw
tri 19574 1044 19594 1064 se
rect 19594 1044 19672 1064
rect 16424 894 16474 1044
rect 19574 1020 19672 1044
rect 19574 986 19622 1020
rect 19656 986 19672 1020
rect 19574 952 19672 986
rect 19574 918 19622 952
rect 19656 918 19672 952
rect 19574 894 19672 918
rect 16424 874 16454 894
tri 16454 874 16474 894 nw
tri 13090 632 13110 652 se
rect 13110 632 13212 652
tri 13212 632 13232 652 sw
tri 19574 874 19594 894 ne
rect 19594 874 19672 894
tri 16332 632 16352 652 se
rect 16352 632 16454 652
tri 16454 632 16474 652 sw
tri 19574 632 19594 652 se
rect 19594 632 19672 652
rect 166 608 264 632
rect 166 574 182 608
rect 216 574 264 608
rect 166 540 264 574
rect 166 506 182 540
rect 216 506 264 540
rect 166 482 264 506
rect 3364 608 3506 632
rect 3364 574 3423 608
rect 3457 574 3506 608
rect 3364 540 3506 574
rect 3364 506 3423 540
rect 3457 506 3506 540
rect 3364 482 3506 506
rect 6606 608 6748 632
rect 6606 574 6665 608
rect 6699 574 6748 608
rect 6606 540 6748 574
rect 6606 506 6665 540
rect 6699 506 6748 540
rect 6606 482 6748 506
rect 9848 608 9990 632
rect 9848 574 9907 608
rect 9941 574 9990 608
rect 9848 540 9990 574
rect 9848 506 9907 540
rect 9941 506 9990 540
rect 9848 482 9990 506
rect 13090 608 13232 632
rect 13090 574 13149 608
rect 13183 574 13232 608
rect 13090 540 13232 574
rect 13090 506 13149 540
rect 13183 506 13232 540
rect 13090 482 13232 506
rect 16332 608 16474 632
rect 16332 574 16391 608
rect 16425 574 16474 608
rect 16332 540 16474 574
rect 16332 506 16391 540
rect 16425 506 16474 540
rect 16332 482 16474 506
rect 19574 608 19672 632
rect 19574 574 19622 608
rect 19656 574 19672 608
rect 19574 540 19672 574
rect 19574 506 19622 540
rect 19656 506 19672 540
rect 19574 482 19672 506
rect 166 462 244 482
tri 244 462 264 482 nw
tri 3364 462 3384 482 ne
rect 3384 462 3486 482
tri 3486 462 3506 482 nw
rect 166 220 244 240
tri 244 220 264 240 sw
tri 6606 462 6626 482 ne
rect 6626 462 6728 482
tri 6728 462 6748 482 nw
tri 3364 220 3384 240 se
rect 3384 220 3486 240
tri 3486 220 3506 240 sw
tri 9848 462 9868 482 ne
rect 9868 462 9970 482
tri 9970 462 9990 482 nw
tri 6606 220 6626 240 se
rect 6626 220 6728 240
tri 6728 220 6748 240 sw
tri 13090 462 13110 482 ne
rect 13110 462 13212 482
tri 13212 462 13232 482 nw
tri 9848 220 9868 240 se
rect 9868 220 9970 240
tri 9970 220 9990 240 sw
tri 16332 462 16352 482 ne
rect 16352 462 16454 482
tri 16454 462 16474 482 nw
tri 13090 220 13110 240 se
rect 13110 220 13140 240
rect 166 196 264 220
rect 166 162 182 196
rect 216 162 264 196
rect 166 128 264 162
rect 166 94 182 128
rect 216 94 264 128
rect 166 70 264 94
rect 3364 196 3506 220
rect 3364 162 3423 196
rect 3457 162 3506 196
rect 3364 128 3506 162
rect 3364 94 3423 128
rect 3457 94 3506 128
rect 3364 70 3506 94
rect 6606 70 6748 220
rect 9848 196 9990 220
rect 9848 162 9907 196
rect 9941 162 9990 196
rect 9848 128 9990 162
rect 9848 94 9907 128
rect 9941 94 9990 128
rect 9848 70 9990 94
rect 13090 70 13140 220
rect 166 50 244 70
tri 244 50 264 70 nw
tri 3364 50 3384 70 ne
rect 3384 50 3486 70
tri 3486 50 3506 70 nw
tri 6606 50 6626 70 ne
rect 6626 50 6728 70
tri 6728 50 6748 70 nw
tri 9848 50 9868 70 ne
rect 9868 50 9970 70
tri 9970 50 9990 70 nw
tri 13090 50 13110 70 ne
rect 13110 50 13140 70
rect 13182 220 13212 240
tri 13212 220 13232 240 sw
tri 19574 462 19594 482 ne
rect 19594 462 19672 482
tri 16332 220 16352 240 se
rect 16352 220 16454 240
tri 16454 220 16474 240 sw
tri 19574 220 19594 240 se
rect 19594 220 19672 240
rect 13182 70 13232 220
rect 16332 196 16474 220
rect 16332 162 16391 196
rect 16425 162 16474 196
rect 16332 128 16474 162
rect 16332 94 16391 128
rect 16425 94 16474 128
rect 16332 70 16474 94
rect 19574 196 19672 220
rect 19574 162 19622 196
rect 19656 162 19672 196
rect 19574 128 19672 162
rect 19574 94 19622 128
rect 19656 94 19672 128
rect 19574 70 19672 94
rect 13182 50 13212 70
tri 13212 50 13232 70 nw
tri 16332 50 16352 70 ne
rect 16352 50 16454 70
tri 16454 50 16474 70 nw
tri 19574 50 19594 70 ne
rect 19594 50 19672 70
<< polycont >>
rect -1519 12436 -1485 12470
rect -1363 12436 -1329 12470
rect -1519 11704 -1485 11738
rect -1363 11704 -1329 11738
rect -1519 10972 -1485 11006
rect -1363 10972 -1329 11006
rect 19654 6084 19688 6118
rect 19722 6084 19756 6118
rect 21796 6084 21830 6118
rect 21864 6084 21898 6118
rect 19663 5884 19697 5918
rect 19731 5884 19765 5918
rect 21805 5884 21839 5918
rect 21873 5884 21907 5918
rect 19654 5658 19688 5692
rect 19722 5658 19756 5692
rect 21796 5658 21830 5692
rect 21864 5658 21898 5692
rect 19697 5457 19731 5491
rect 19765 5457 19799 5491
rect 21839 5457 21873 5491
rect 21907 5457 21941 5491
rect -1580 2886 -1546 2920
rect -1485 2886 -1451 2920
rect -1390 2886 -1356 2920
rect -1137 2886 -1103 2920
rect -1042 2886 -1008 2920
rect -947 2886 -913 2920
rect -1580 2080 -1546 2114
rect -1485 2080 -1451 2114
rect -1390 2080 -1356 2114
rect 182 1398 216 1432
rect 182 1330 216 1364
rect 3423 1398 3457 1432
rect 3423 1330 3457 1364
rect 9907 1398 9941 1432
rect 9907 1330 9941 1364
rect 16392 1398 16426 1432
rect 16392 1330 16426 1364
rect 19622 1398 19656 1432
rect 19622 1330 19656 1364
rect 182 986 216 1020
rect 182 918 216 952
rect 3423 986 3457 1020
rect 3423 918 3457 952
rect 6665 986 6699 1020
rect 6665 918 6699 952
rect 9907 986 9941 1020
rect 9907 918 9941 952
rect 13150 986 13184 1020
rect 13150 918 13184 952
rect 19622 986 19656 1020
rect 19622 918 19656 952
rect 182 574 216 608
rect 182 506 216 540
rect 3423 574 3457 608
rect 3423 506 3457 540
rect 6665 574 6699 608
rect 6665 506 6699 540
rect 9907 574 9941 608
rect 9907 506 9941 540
rect 13149 574 13183 608
rect 13149 506 13183 540
rect 16391 574 16425 608
rect 16391 506 16425 540
rect 19622 574 19656 608
rect 19622 506 19656 540
rect 182 162 216 196
rect 182 94 216 128
rect 3423 162 3457 196
rect 3423 94 3457 128
rect 9907 162 9941 196
rect 9907 94 9941 128
rect 16391 162 16425 196
rect 16391 94 16425 128
rect 19622 162 19656 196
rect 19622 94 19656 128
<< npolyres >>
rect 19756 6051 21796 6151
rect 19799 5424 21839 5524
<< locali >>
rect -668 16925 -498 16959
rect -2119 14521 -668 14527
rect -2119 14517 -2040 14521
rect -2006 14517 -1967 14521
rect -1933 14517 -1894 14521
rect -1860 14517 -1821 14521
rect -1787 14517 -1748 14521
rect -1714 14517 -1675 14521
rect -1641 14517 -1601 14521
rect -1567 14517 -1527 14521
rect -1493 14517 -1453 14521
rect -1419 14517 -1379 14521
rect -1345 14517 -1305 14521
rect -1271 14517 -1231 14521
rect -1197 14517 -1157 14521
rect -1123 14517 -1083 14521
rect -1049 14517 -1009 14521
rect -975 14517 -935 14521
rect -901 14517 -861 14521
rect -827 14517 -787 14521
rect -753 14517 -713 14521
rect -679 14517 -668 14521
rect -2119 14449 -2041 14517
rect -1567 14487 -1564 14517
rect -1599 14483 -1564 14487
rect -1530 14487 -1527 14517
rect -1461 14487 -1453 14517
rect -1392 14487 -1379 14517
rect -1323 14487 -1305 14517
rect -1254 14487 -1231 14517
rect -1185 14487 -1157 14517
rect -1116 14487 -1083 14517
rect -1530 14483 -1495 14487
rect -1461 14483 -1426 14487
rect -1392 14483 -1357 14487
rect -1323 14483 -1288 14487
rect -1254 14483 -1219 14487
rect -1185 14483 -1150 14487
rect -1116 14483 -1081 14487
rect -1047 14483 -1012 14517
rect -975 14487 -943 14517
rect -901 14487 -874 14517
rect -827 14487 -805 14517
rect -753 14487 -736 14517
rect -978 14483 -943 14487
rect -909 14483 -874 14487
rect -840 14483 -805 14487
rect -771 14483 -736 14487
rect -1599 14449 -736 14483
rect -2119 14415 -2113 14449
rect -2075 14415 -2041 14449
rect -1567 14415 -1564 14449
rect -1530 14415 -1527 14449
rect -1461 14415 -1453 14449
rect -1392 14415 -1379 14449
rect -1323 14415 -1305 14449
rect -1254 14415 -1231 14449
rect -1185 14415 -1157 14449
rect -1116 14415 -1083 14449
rect -1047 14415 -1012 14449
rect -975 14415 -943 14449
rect -901 14415 -874 14449
rect -827 14415 -805 14449
rect -753 14415 -736 14449
rect -2119 14380 -1973 14415
rect -2119 14376 -2109 14380
rect -2119 14342 -2113 14376
rect -2075 14346 -2041 14380
rect -2007 14347 -1973 14380
rect -1599 14381 -736 14415
rect -1599 14377 -1564 14381
rect -1567 14347 -1564 14377
rect -1530 14377 -1495 14381
rect -1461 14377 -1426 14381
rect -1392 14377 -1357 14381
rect -1323 14377 -1288 14381
rect -1254 14377 -1219 14381
rect -1185 14377 -1150 14381
rect -1116 14377 -1081 14381
rect -1530 14347 -1527 14377
rect -1461 14347 -1453 14377
rect -1392 14347 -1379 14377
rect -1323 14347 -1305 14377
rect -1254 14347 -1231 14377
rect -1185 14347 -1157 14377
rect -1116 14347 -1083 14377
rect -1047 14347 -1012 14381
rect -978 14377 -943 14381
rect -909 14377 -874 14381
rect -840 14377 -805 14381
rect -771 14377 -736 14381
rect -975 14347 -943 14377
rect -901 14347 -874 14377
rect -827 14347 -805 14377
rect -753 14347 -736 14377
rect -2079 14342 -2041 14346
rect -2007 14343 -1969 14347
rect -1935 14343 -1896 14347
rect -1862 14343 -1823 14347
rect -1789 14343 -1749 14347
rect -1715 14343 -1675 14347
rect -1641 14343 -1601 14347
rect -1567 14343 -1527 14347
rect -1493 14343 -1453 14347
rect -1419 14343 -1379 14347
rect -1345 14343 -1305 14347
rect -1271 14343 -1231 14347
rect -1197 14343 -1157 14347
rect -1123 14343 -1083 14347
rect -1049 14343 -1009 14347
rect -975 14343 -935 14347
rect -901 14343 -861 14347
rect -827 14343 -787 14347
rect -753 14343 -713 14347
rect -679 14343 -668 14347
rect -2007 14342 -668 14343
rect -2119 14337 -668 14342
rect -2119 14312 -1929 14337
rect -2119 14311 -1973 14312
rect -2119 14303 -2109 14311
rect -2119 14269 -2113 14303
rect -2075 14277 -2041 14311
rect -2007 14278 -1973 14311
rect -1939 14304 -1929 14312
rect -2079 14269 -2041 14277
rect -2007 14270 -1969 14278
rect -1935 14270 -1929 14304
rect -2007 14269 -1929 14270
rect -2119 14243 -1929 14269
rect -2119 14242 -1973 14243
rect -2119 14230 -2109 14242
rect -2119 14196 -2113 14230
rect -2075 14208 -2041 14242
rect -2007 14209 -1973 14242
rect -1939 14231 -1929 14243
rect -2079 14196 -2041 14208
rect -2007 14197 -1969 14209
rect -1935 14197 -1929 14231
rect -2007 14196 -1929 14197
rect -2119 14174 -1929 14196
rect -2119 14173 -1973 14174
rect -2119 14157 -2109 14173
rect -2119 14123 -2113 14157
rect -2075 14139 -2041 14173
rect -2007 14140 -1973 14173
rect -1939 14158 -1929 14174
rect -2079 14123 -2041 14139
rect -2007 14124 -1969 14140
rect -1935 14124 -1929 14158
rect -2007 14123 -1929 14124
rect -2119 14105 -1929 14123
rect -2119 14104 -1973 14105
rect -2119 14084 -2109 14104
rect -2119 14050 -2113 14084
rect -2075 14070 -2041 14104
rect -2007 14071 -1973 14104
rect -1939 14085 -1929 14105
rect -2079 14050 -2041 14070
rect -2007 14051 -1969 14071
rect -1935 14051 -1929 14085
rect -2007 14050 -1929 14051
rect -2119 14036 -1929 14050
rect -2119 14035 -1973 14036
rect -2119 14011 -2109 14035
rect -2119 13977 -2113 14011
rect -2075 14001 -2041 14035
rect -2007 14002 -1973 14035
rect -1939 14012 -1929 14036
rect -2079 13977 -2041 14001
rect -2007 13978 -1969 14002
rect -1935 13978 -1929 14012
rect -2007 13977 -1929 13978
rect -2119 13967 -1929 13977
rect -2119 13966 -1973 13967
rect -2119 13938 -2109 13966
rect -2119 13904 -2113 13938
rect -2075 13932 -2041 13966
rect -2007 13933 -1973 13966
rect -1939 13939 -1929 13967
rect -2079 13904 -2041 13932
rect -2007 13905 -1969 13933
rect -1935 13905 -1929 13939
rect -2007 13904 -1929 13905
rect -2119 13898 -1929 13904
rect -2119 13897 -1973 13898
rect -2119 13865 -2109 13897
rect -2119 13831 -2113 13865
rect -2075 13863 -2041 13897
rect -2007 13864 -1973 13897
rect -1939 13866 -1929 13898
rect -2079 13831 -2041 13863
rect -2007 13832 -1969 13864
rect -1935 13832 -1929 13866
rect -2007 13831 -1929 13832
rect -2119 13829 -1929 13831
rect -2119 13828 -1973 13829
rect -2119 13794 -2109 13828
rect -2075 13794 -2041 13828
rect -2007 13795 -1973 13828
rect -1939 13795 -1929 13829
rect -2007 13794 -1929 13795
rect -2119 13793 -1929 13794
rect -2119 13792 -1969 13793
rect -2119 13758 -2113 13792
rect -2079 13759 -2041 13792
rect -2007 13760 -1969 13792
rect -2119 13725 -2109 13758
rect -2075 13725 -2041 13759
rect -2007 13726 -1973 13760
rect -1935 13759 -1929 13793
rect -1939 13726 -1929 13759
rect -2007 13725 -1929 13726
rect -2119 13720 -1929 13725
rect -2119 13719 -1969 13720
rect -2119 13685 -2113 13719
rect -2079 13690 -2041 13719
rect -2007 13691 -1969 13719
rect -2119 13656 -2109 13685
rect -2075 13656 -2041 13690
rect -2007 13657 -1973 13691
rect -1935 13686 -1929 13720
rect -1939 13657 -1929 13686
rect -2007 13656 -1929 13657
rect -2119 13647 -1929 13656
rect -2119 13646 -1969 13647
rect -2119 13612 -2113 13646
rect -2079 13621 -2041 13646
rect -2007 13622 -1969 13646
rect -2119 13587 -2109 13612
rect -2075 13587 -2041 13621
rect -2007 13588 -1973 13622
rect -1935 13613 -1929 13647
rect -1939 13588 -1929 13613
rect -2007 13587 -1929 13588
rect -2119 13574 -1929 13587
rect -2119 13573 -1969 13574
rect -2119 13539 -2113 13573
rect -2079 13552 -2041 13573
rect -2007 13553 -1969 13573
rect -2119 13518 -2109 13539
rect -2075 13518 -2041 13552
rect -2007 13519 -1973 13553
rect -1935 13540 -1929 13574
rect -1939 13519 -1929 13540
rect -2007 13518 -1929 13519
rect -2119 13501 -1929 13518
rect -2119 13500 -1969 13501
rect -2119 13466 -2113 13500
rect -2079 13483 -2041 13500
rect -2007 13484 -1969 13500
rect -2119 13449 -2109 13466
rect -2075 13449 -2041 13483
rect -2007 13450 -1973 13484
rect -1935 13467 -1929 13501
rect -1939 13450 -1929 13467
rect -2007 13449 -1929 13450
rect -2119 13428 -1929 13449
rect -2119 13427 -1969 13428
rect -2119 13393 -2113 13427
rect -2079 13414 -2041 13427
rect -2007 13415 -1969 13427
rect -2119 13380 -2109 13393
rect -2075 13380 -2041 13414
rect -2007 13381 -1973 13415
rect -1935 13394 -1929 13428
rect -1939 13381 -1929 13394
rect -2007 13380 -1929 13381
rect -2119 13355 -1929 13380
rect -2119 13354 -1969 13355
rect -2119 13320 -2113 13354
rect -2079 13345 -2041 13354
rect -2007 13346 -1969 13354
rect -2119 13311 -2109 13320
rect -2075 13311 -2041 13345
rect -2007 13312 -1973 13346
rect -1935 13321 -1929 13355
rect -1939 13312 -1929 13321
rect -2007 13311 -1929 13312
rect -2119 13282 -1929 13311
rect -2119 13281 -1969 13282
rect -2119 13247 -2113 13281
rect -2079 13276 -2041 13281
rect -2007 13277 -1969 13281
rect -2119 13242 -2109 13247
rect -2075 13242 -2041 13276
rect -2007 13243 -1973 13277
rect -1935 13248 -1929 13282
rect -1939 13243 -1929 13248
rect -2007 13242 -1929 13243
rect -2119 13209 -1929 13242
rect -2119 13208 -1969 13209
rect -2119 13174 -2113 13208
rect -2079 13207 -2041 13208
rect -2119 13173 -2109 13174
rect -2075 13173 -2041 13207
rect -2007 13174 -1973 13208
rect -1935 13175 -1929 13209
rect -1939 13174 -1929 13175
rect -2007 13173 -1929 13174
rect -2119 13139 -1929 13173
rect -2119 13138 -1973 13139
rect -2119 13135 -2109 13138
rect -2119 13101 -2113 13135
rect -2075 13104 -2041 13138
rect -2007 13105 -1973 13138
rect -1939 13136 -1929 13139
rect -2079 13101 -2041 13104
rect -2007 13102 -1969 13105
rect -1935 13102 -1929 13136
rect -2007 13101 -1929 13102
rect -2119 13070 -1929 13101
rect -2119 13069 -1973 13070
rect -2119 13062 -2109 13069
rect -2119 13028 -2113 13062
rect -2075 13035 -2041 13069
rect -2007 13036 -1973 13069
rect -1939 13063 -1929 13070
rect -2079 13028 -2041 13035
rect -2007 13029 -1969 13036
rect -1935 13029 -1929 13063
rect -2007 13028 -1929 13029
rect -2119 13001 -1929 13028
rect -2119 13000 -1973 13001
rect -2119 12989 -2109 13000
rect -2119 12955 -2113 12989
rect -2075 12966 -2041 13000
rect -2007 12967 -1973 13000
rect -1939 12990 -1929 13001
rect -2079 12955 -2041 12966
rect -2007 12956 -1969 12967
rect -1935 12956 -1929 12990
rect -2007 12955 -1929 12956
rect -2119 12932 -1929 12955
rect -2119 12931 -1973 12932
rect -2119 12916 -2109 12931
rect -2119 12882 -2113 12916
rect -2075 12897 -2041 12931
rect -2007 12898 -1973 12931
rect -1939 12917 -1929 12932
rect -2079 12882 -2041 12897
rect -2007 12883 -1969 12898
rect -1935 12883 -1929 12917
rect -2007 12882 -1929 12883
rect -2119 12863 -1929 12882
rect -2119 12862 -1973 12863
rect -2119 12843 -2109 12862
rect -2119 12809 -2113 12843
rect -2075 12828 -2041 12862
rect -2007 12829 -1973 12862
rect -1939 12844 -1929 12863
rect -2079 12809 -2041 12828
rect -2007 12810 -1969 12829
rect -1935 12810 -1929 12844
rect -2007 12809 -1929 12810
rect -2119 12794 -1929 12809
rect -2119 12793 -1973 12794
rect -2119 12770 -2109 12793
rect -2119 12736 -2113 12770
rect -2075 12759 -2041 12793
rect -2007 12760 -1973 12793
rect -1939 12771 -1929 12794
rect -2079 12736 -2041 12759
rect -2007 12737 -1969 12760
rect -1935 12737 -1929 12771
rect -2007 12736 -1929 12737
rect -2119 12725 -1929 12736
rect -2119 12724 -1973 12725
rect -2119 12697 -2109 12724
rect -2119 12663 -2113 12697
rect -2075 12690 -2041 12724
rect -2007 12691 -1973 12724
rect -1939 12698 -1929 12725
rect -2079 12663 -2041 12690
rect -2007 12664 -1969 12691
rect -1935 12664 -1929 12698
rect -2007 12663 -1929 12664
rect -2119 12656 -1929 12663
rect -2119 12655 -1973 12656
rect -2119 12624 -2109 12655
rect -2119 12590 -2113 12624
rect -2075 12621 -2041 12655
rect -2007 12622 -1973 12655
rect -1939 12625 -1929 12656
rect -2079 12590 -2041 12621
rect -2007 12591 -1969 12622
rect -1935 12591 -1929 12625
rect -2007 12590 -1929 12591
rect -2119 12587 -1929 12590
rect -2119 12586 -1973 12587
rect -2119 12552 -2109 12586
rect -2075 12552 -2041 12586
rect -2007 12553 -1973 12586
rect -1939 12553 -1929 12587
rect -2007 12552 -1929 12553
rect -2119 12551 -1969 12552
rect -2119 12517 -2113 12551
rect -2079 12517 -2041 12551
rect -2007 12518 -1969 12551
rect -1935 12518 -1929 12552
rect -2119 12483 -2109 12517
rect -2075 12483 -2041 12517
rect -2007 12484 -1973 12518
rect -1939 12484 -1929 12518
rect -2007 12483 -1929 12484
rect -2119 12479 -1929 12483
rect -2119 12478 -1969 12479
rect -2119 12444 -2113 12478
rect -2079 12448 -2041 12478
rect -2007 12449 -1969 12478
rect -2119 12414 -2109 12444
rect -2075 12414 -2041 12448
rect -2007 12415 -1973 12449
rect -1935 12445 -1929 12479
rect -1939 12415 -1929 12445
rect -2007 12414 -1929 12415
rect -2119 12406 -1929 12414
rect -2119 12405 -1969 12406
rect -2119 12371 -2113 12405
rect -2079 12379 -2041 12405
rect -2007 12380 -1969 12405
rect -2119 12345 -2109 12371
rect -2075 12345 -2041 12379
rect -2007 12346 -1973 12380
rect -1935 12372 -1929 12406
rect -1939 12346 -1929 12372
rect -2007 12345 -1929 12346
rect -2119 12333 -1929 12345
rect -2119 12332 -1969 12333
rect -2119 12298 -2113 12332
rect -2079 12310 -2041 12332
rect -2007 12311 -1969 12332
rect -2119 12276 -2109 12298
rect -2075 12276 -2041 12310
rect -2007 12277 -1973 12311
rect -1935 12299 -1929 12333
rect -1939 12277 -1929 12299
rect -2007 12276 -1929 12277
rect -2119 12260 -1929 12276
rect -2119 12259 -1969 12260
rect -2119 12225 -2113 12259
rect -2079 12241 -2041 12259
rect -2007 12242 -1969 12259
rect -2119 12207 -2109 12225
rect -2075 12207 -2041 12241
rect -2007 12208 -1973 12242
rect -1935 12226 -1929 12260
rect -1939 12208 -1929 12226
rect -2007 12207 -1929 12208
rect -2119 12187 -1929 12207
rect -2119 12186 -1969 12187
rect -2119 7616 -2113 12186
rect -2007 12173 -1969 12186
rect -2007 12139 -1973 12173
rect -1935 12153 -1929 12187
rect -1939 12139 -1929 12153
rect -2007 12114 -1929 12139
rect -1935 7728 -1929 12114
rect -1795 14197 -1053 14203
rect -1795 14161 -1711 14197
rect -1677 14163 -1633 14197
rect -1599 14195 -1555 14197
rect -1521 14195 -1477 14197
rect -1443 14195 -1399 14197
rect -1365 14195 -1321 14197
rect -1287 14195 -1243 14197
rect -1209 14195 -1165 14197
rect -1131 14195 -1053 14197
rect -1599 14163 -1571 14195
rect -1677 14161 -1571 14163
rect -1795 14127 -1571 14161
rect -1795 14125 -1787 14127
rect -1685 14125 -1571 14127
rect -1129 14125 -1053 14195
rect -1795 14091 -1789 14125
rect -1683 14091 -1633 14125
rect -1599 14093 -1571 14125
rect -1599 14091 -1555 14093
rect -1521 14091 -1477 14093
rect -1443 14091 -1399 14093
rect -1365 14091 -1321 14093
rect -1287 14091 -1243 14093
rect -1209 14091 -1165 14093
rect -1795 14052 -1787 14091
rect -1685 14085 -1165 14091
rect -1685 14052 -1677 14085
rect -1795 14018 -1789 14052
rect -1683 14018 -1677 14052
rect -1795 13979 -1787 14018
rect -1685 13979 -1677 14018
rect -1795 13945 -1789 13979
rect -1683 13945 -1677 13979
rect -1795 13906 -1787 13945
rect -1685 13906 -1677 13945
rect -1795 13872 -1789 13906
rect -1683 13872 -1677 13906
rect -1795 13833 -1787 13872
rect -1685 13833 -1677 13872
rect -1795 13799 -1789 13833
rect -1683 13799 -1677 13833
rect -1795 13760 -1787 13799
rect -1685 13760 -1677 13799
rect -1795 13726 -1789 13760
rect -1683 13726 -1677 13760
rect -1795 13687 -1787 13726
rect -1685 13687 -1677 13726
rect -1795 13653 -1789 13687
rect -1683 13653 -1677 13687
rect -1795 13614 -1787 13653
rect -1685 13614 -1677 13653
rect -1795 13580 -1789 13614
rect -1683 13580 -1677 13614
rect -1795 13541 -1787 13580
rect -1685 13541 -1677 13580
rect -1795 13507 -1789 13541
rect -1683 13507 -1677 13541
rect -1795 13468 -1787 13507
rect -1685 13468 -1677 13507
rect -1795 7962 -1789 13468
rect -1683 8002 -1677 13468
rect -1171 14019 -1165 14085
rect -1059 14019 -1053 14125
rect -1171 13980 -1163 14019
rect -1061 13980 -1053 14019
rect -1171 13946 -1165 13980
rect -1059 13946 -1053 13980
rect -1171 13907 -1163 13946
rect -1061 13907 -1053 13946
rect -1171 13873 -1165 13907
rect -1059 13873 -1053 13907
rect -1171 13834 -1163 13873
rect -1061 13834 -1053 13873
rect -1171 13800 -1165 13834
rect -1059 13800 -1053 13834
rect -1171 13761 -1163 13800
rect -1061 13761 -1053 13800
rect -1171 13727 -1165 13761
rect -1059 13727 -1053 13761
rect -1171 13688 -1163 13727
rect -1061 13688 -1053 13727
rect -1171 13654 -1165 13688
rect -1059 13654 -1053 13688
rect -1171 13615 -1163 13654
rect -1061 13615 -1053 13654
rect -1171 13581 -1165 13615
rect -1059 13581 -1053 13615
rect -1171 13542 -1163 13581
rect -1061 13542 -1053 13581
rect -1171 13508 -1165 13542
rect -1059 13508 -1053 13542
rect -1171 13469 -1163 13508
rect -1061 13469 -1053 13508
rect -1171 13435 -1165 13469
rect -1059 13435 -1053 13469
rect -1171 13396 -1163 13435
rect -1061 13396 -1053 13435
rect -1171 13362 -1165 13396
rect -1059 13362 -1053 13396
rect -1171 13323 -1163 13362
rect -1061 13323 -1053 13362
rect -1171 13289 -1165 13323
rect -1059 13289 -1053 13323
rect -1171 13250 -1163 13289
rect -1061 13250 -1053 13289
rect -1171 13216 -1165 13250
rect -1059 13216 -1053 13250
rect -1171 13177 -1163 13216
rect -1061 13177 -1053 13216
rect -1171 13143 -1165 13177
rect -1059 13143 -1053 13177
rect -1171 13104 -1163 13143
rect -1061 13104 -1053 13143
rect -1171 13070 -1165 13104
rect -1059 13070 -1053 13104
rect -1171 13031 -1163 13070
rect -1061 13031 -1053 13070
rect -1171 12997 -1165 13031
rect -1059 12997 -1053 13031
rect -1171 12958 -1163 12997
rect -1061 12958 -1053 12997
rect -1171 12924 -1165 12958
rect -1059 12924 -1053 12958
rect -1171 12885 -1163 12924
rect -1061 12885 -1053 12924
rect -1171 12851 -1165 12885
rect -1059 12851 -1053 12885
rect -1171 12812 -1163 12851
rect -1061 12812 -1053 12851
rect -1171 12778 -1165 12812
rect -1059 12778 -1053 12812
rect -1171 12739 -1163 12778
rect -1061 12739 -1053 12778
rect -1171 12705 -1165 12739
rect -1059 12705 -1053 12739
rect -1171 12666 -1163 12705
rect -1061 12666 -1053 12705
rect -1171 12632 -1165 12666
rect -1059 12632 -1053 12666
rect -1171 12568 -1163 12632
rect -1061 12568 -1053 12632
rect -1171 12534 -1165 12568
rect -1059 12534 -1053 12568
rect -1526 12472 -1519 12487
rect -1485 12477 -1478 12487
rect -1370 12477 -1363 12487
rect -1485 12472 -1363 12477
rect -1171 12495 -1163 12534
rect -1061 12495 -1053 12534
rect -1329 12472 -1322 12487
rect -1526 12470 -1322 12472
rect -1526 12436 -1519 12470
rect -1485 12436 -1363 12470
rect -1329 12436 -1322 12470
rect -1526 12434 -1322 12436
rect -1526 12420 -1519 12434
rect -1485 12429 -1363 12434
rect -1485 12420 -1478 12429
rect -1370 12420 -1363 12429
rect -1329 12420 -1322 12434
rect -1171 12461 -1165 12495
rect -1059 12461 -1053 12495
rect -1171 12422 -1163 12461
rect -1061 12422 -1053 12461
rect -1171 12388 -1165 12422
rect -1059 12388 -1053 12422
rect -1171 12349 -1163 12388
rect -1061 12349 -1053 12388
rect -1597 12321 -1563 12325
rect -1597 12249 -1563 12275
rect -1597 12177 -1563 12207
rect -1597 12105 -1563 12139
rect -1597 12037 -1563 12071
rect -1597 11969 -1563 11999
rect -1597 11901 -1563 11927
rect -1597 11833 -1563 11855
rect -1441 12321 -1407 12325
rect -1441 12249 -1407 12275
rect -1441 12177 -1407 12207
rect -1441 12105 -1407 12139
rect -1441 12037 -1407 12071
rect -1441 11969 -1407 11999
rect -1441 11901 -1407 11927
rect -1441 11833 -1407 11855
rect -1285 12321 -1251 12325
rect -1285 12249 -1251 12275
rect -1285 12177 -1251 12207
rect -1285 12105 -1251 12139
rect -1285 12037 -1251 12071
rect -1285 11969 -1251 11999
rect -1285 11901 -1251 11927
rect -1285 11833 -1251 11855
rect -1171 12315 -1165 12349
rect -1059 12315 -1053 12349
rect -1171 12276 -1163 12315
rect -1061 12276 -1053 12315
rect -1171 12242 -1165 12276
rect -1059 12242 -1053 12276
rect -1171 12203 -1163 12242
rect -1061 12203 -1053 12242
rect -1171 12169 -1165 12203
rect -1059 12169 -1053 12203
rect -1171 12130 -1163 12169
rect -1061 12130 -1053 12169
rect -1171 12096 -1165 12130
rect -1059 12096 -1053 12130
rect -1171 12057 -1163 12096
rect -1061 12057 -1053 12096
rect -1171 12023 -1165 12057
rect -1059 12023 -1053 12057
rect -1171 11984 -1163 12023
rect -1061 11984 -1053 12023
rect -1171 11950 -1165 11984
rect -1059 11950 -1053 11984
rect -1171 11911 -1163 11950
rect -1061 11911 -1053 11950
rect -1171 11877 -1165 11911
rect -1059 11877 -1053 11911
rect -1171 11838 -1163 11877
rect -1061 11838 -1053 11877
rect -1171 11804 -1165 11838
rect -1059 11804 -1053 11838
rect -1526 11740 -1519 11755
rect -1485 11745 -1478 11755
rect -1370 11745 -1363 11755
rect -1485 11740 -1363 11745
rect -1171 11765 -1163 11804
rect -1061 11765 -1053 11804
rect -1329 11740 -1322 11755
rect -1526 11738 -1322 11740
rect -1526 11704 -1519 11738
rect -1485 11704 -1363 11738
rect -1329 11704 -1322 11738
rect -1526 11702 -1322 11704
rect -1526 11688 -1519 11702
rect -1485 11697 -1363 11702
rect -1485 11688 -1478 11697
rect -1370 11688 -1363 11697
rect -1329 11688 -1322 11702
rect -1171 11731 -1165 11765
rect -1059 11731 -1053 11765
rect -1171 11692 -1163 11731
rect -1061 11692 -1053 11731
rect -1597 11587 -1563 11609
rect -1597 11515 -1563 11541
rect -1597 11443 -1563 11473
rect -1597 11371 -1563 11405
rect -1597 11303 -1563 11337
rect -1597 11235 -1563 11265
rect -1597 11167 -1563 11193
rect -1597 11117 -1563 11121
rect -1441 11587 -1407 11609
rect -1441 11515 -1407 11541
rect -1441 11443 -1407 11473
rect -1441 11371 -1407 11405
rect -1441 11303 -1407 11337
rect -1441 11235 -1407 11265
rect -1441 11167 -1407 11193
rect -1441 11117 -1407 11121
rect -1285 11587 -1251 11609
rect -1285 11515 -1251 11541
rect -1285 11443 -1251 11473
rect -1285 11371 -1251 11405
rect -1285 11303 -1251 11337
rect -1285 11235 -1251 11265
rect -1285 11167 -1251 11193
rect -1285 11117 -1251 11121
rect -1171 11658 -1165 11692
rect -1059 11658 -1053 11692
rect -1171 11619 -1163 11658
rect -1061 11619 -1053 11658
rect -1171 11585 -1165 11619
rect -1059 11585 -1053 11619
rect -1171 11546 -1163 11585
rect -1061 11546 -1053 11585
rect -1171 11512 -1165 11546
rect -1059 11512 -1053 11546
rect -1171 11473 -1163 11512
rect -1061 11473 -1053 11512
rect -1171 11439 -1165 11473
rect -1059 11439 -1053 11473
rect -1171 11400 -1163 11439
rect -1061 11400 -1053 11439
rect -1171 11366 -1165 11400
rect -1059 11366 -1053 11400
rect -1171 11327 -1163 11366
rect -1061 11327 -1053 11366
rect -1171 11293 -1165 11327
rect -1059 11293 -1053 11327
rect -1171 11254 -1163 11293
rect -1061 11254 -1053 11293
rect -1171 11220 -1165 11254
rect -1059 11220 -1053 11254
rect -1171 11181 -1163 11220
rect -1061 11181 -1053 11220
rect -1171 11147 -1165 11181
rect -1059 11147 -1053 11181
rect -1171 11108 -1163 11147
rect -1061 11108 -1053 11147
rect -1171 11074 -1165 11108
rect -1059 11074 -1053 11108
rect -1526 11008 -1519 11023
rect -1485 11013 -1478 11023
rect -1370 11013 -1363 11023
rect -1485 11008 -1363 11013
rect -1171 11035 -1163 11074
rect -1061 11035 -1053 11074
rect -1329 11008 -1322 11023
rect -1526 11006 -1322 11008
rect -1526 10972 -1519 11006
rect -1485 10972 -1363 11006
rect -1329 10972 -1322 11006
rect -1526 10970 -1322 10972
rect -1526 10956 -1519 10970
rect -1485 10965 -1363 10970
rect -1485 10956 -1478 10965
rect -1370 10956 -1363 10965
rect -1329 10956 -1322 10970
rect -1171 11001 -1165 11035
rect -1059 11001 -1053 11035
rect -1171 10962 -1163 11001
rect -1061 10962 -1053 11001
rect -1171 10928 -1165 10962
rect -1059 10928 -1053 10962
rect -1171 10889 -1163 10928
rect -1061 10889 -1053 10928
rect -1597 10857 -1563 10861
rect -1597 10785 -1563 10811
rect -1597 10713 -1563 10743
rect -1597 10641 -1563 10675
rect -1597 10573 -1563 10607
rect -1597 10505 -1563 10535
rect -1597 10437 -1563 10463
rect -1597 10369 -1563 10391
rect -1441 10857 -1407 10861
rect -1441 10785 -1407 10811
rect -1441 10713 -1407 10743
rect -1441 10641 -1407 10675
rect -1441 10573 -1407 10607
rect -1441 10505 -1407 10535
rect -1441 10437 -1407 10463
rect -1441 10369 -1407 10391
rect -1285 10857 -1251 10861
rect -1285 10785 -1251 10811
rect -1285 10713 -1251 10743
rect -1285 10641 -1251 10675
rect -1285 10573 -1251 10607
rect -1285 10505 -1251 10535
rect -1285 10437 -1251 10463
rect -1285 10369 -1251 10391
rect -1171 10855 -1165 10889
rect -1059 10855 -1053 10889
rect -1171 10816 -1163 10855
rect -1061 10816 -1053 10855
rect -1171 10782 -1165 10816
rect -1059 10782 -1053 10816
rect -1171 10743 -1163 10782
rect -1061 10743 -1053 10782
rect -1171 10709 -1165 10743
rect -1059 10709 -1053 10743
rect -1171 10670 -1163 10709
rect -1061 10670 -1053 10709
rect -1171 10636 -1165 10670
rect -1059 10636 -1053 10670
rect -1171 10597 -1163 10636
rect -1061 10597 -1053 10636
rect -1171 10563 -1165 10597
rect -1059 10563 -1053 10597
rect -1171 10524 -1163 10563
rect -1061 10524 -1053 10563
rect -1171 10490 -1165 10524
rect -1059 10490 -1053 10524
rect -1171 10451 -1163 10490
rect -1061 10451 -1053 10490
rect -1171 10417 -1165 10451
rect -1059 10417 -1053 10451
rect -1171 10378 -1163 10417
rect -1061 10378 -1053 10417
rect -1171 10344 -1165 10378
rect -1059 10344 -1053 10378
rect -1171 10305 -1163 10344
rect -1061 10305 -1053 10344
rect -1171 10271 -1165 10305
rect -1059 10271 -1053 10305
rect -1171 10232 -1163 10271
rect -1061 10232 -1053 10271
rect -1171 10198 -1165 10232
rect -1059 10198 -1053 10232
rect -1171 10159 -1163 10198
rect -1061 10159 -1053 10198
rect -1171 10125 -1165 10159
rect -1059 10125 -1053 10159
rect -1171 10086 -1163 10125
rect -1061 10086 -1053 10125
rect -1171 10052 -1165 10086
rect -1059 10052 -1053 10086
rect -1171 10013 -1163 10052
rect -1061 10013 -1053 10052
rect -1171 8035 -1165 10013
rect -1059 8035 -1053 10013
rect -1171 8002 -1163 8035
rect -1683 7996 -1163 8002
rect -1683 7994 -1641 7996
rect -1607 7994 -1565 7996
rect -1531 7994 -1490 7996
rect -1456 7994 -1415 7996
rect -1381 7994 -1340 7996
rect -1306 7994 -1265 7996
rect -1231 7994 -1190 7996
rect -1209 7962 -1190 7994
rect -1795 7892 -1719 7962
rect -1209 7960 -1163 7962
rect -1061 7960 -1053 8035
rect -1209 7947 -1053 7960
rect -1209 7926 -1093 7947
rect -1209 7892 -1175 7926
rect -1141 7924 -1093 7926
rect -1137 7913 -1093 7924
rect -1059 7913 -1053 7947
rect -1795 7890 -1717 7892
rect -1683 7890 -1639 7892
rect -1605 7890 -1561 7892
rect -1527 7890 -1483 7892
rect -1449 7890 -1405 7892
rect -1371 7890 -1327 7892
rect -1293 7890 -1249 7892
rect -1215 7890 -1171 7892
rect -1137 7890 -1053 7913
rect -1795 7884 -1053 7890
rect -668 7948 -498 7983
rect -634 7914 -600 7948
rect -566 7914 -532 7948
rect -668 7879 -498 7914
rect -634 7845 -600 7879
rect -566 7845 -532 7879
rect -668 7810 -498 7845
rect -634 7776 -600 7810
rect -566 7776 -532 7810
rect -668 7741 -498 7776
rect -1935 7722 -668 7728
rect -1935 7719 -1895 7722
rect -1861 7719 -1821 7722
rect -1787 7719 -1747 7722
rect -1713 7719 -1673 7722
rect -1639 7719 -1599 7722
rect -1565 7719 -1525 7722
rect -1935 7688 -1904 7719
rect -1861 7688 -1835 7719
rect -1787 7688 -1766 7719
rect -1713 7688 -1697 7719
rect -1639 7688 -1628 7719
rect -1565 7688 -1559 7719
rect -1939 7685 -1904 7688
rect -1870 7685 -1835 7688
rect -1801 7685 -1766 7688
rect -1732 7685 -1697 7688
rect -1663 7685 -1628 7688
rect -1594 7685 -1559 7688
rect -1491 7719 -1451 7722
rect -1417 7719 -1377 7722
rect -1343 7719 -1303 7722
rect -1269 7719 -1229 7722
rect -1195 7719 -1155 7722
rect -1121 7719 -1081 7722
rect -1047 7719 -1007 7722
rect -973 7719 -933 7722
rect -899 7719 -859 7722
rect -825 7719 -786 7722
rect -752 7719 -713 7722
rect -1491 7688 -1490 7719
rect -1525 7685 -1490 7688
rect -1456 7688 -1451 7719
rect -1387 7688 -1377 7719
rect -1318 7688 -1303 7719
rect -1249 7688 -1229 7719
rect -1180 7688 -1155 7719
rect -1111 7688 -1081 7719
rect -679 7707 -668 7722
rect -634 7707 -600 7741
rect -566 7707 -532 7741
rect -679 7688 -498 7707
rect -1456 7685 -1421 7688
rect -1387 7685 -1352 7688
rect -1318 7685 -1283 7688
rect -1249 7685 -1214 7688
rect -1180 7685 -1145 7688
rect -1111 7685 -1076 7688
rect -2007 7651 -1076 7685
rect -702 7672 -498 7688
rect -2007 7617 -1972 7651
rect -1938 7650 -1903 7651
rect -1869 7650 -1834 7651
rect -1800 7650 -1765 7651
rect -1731 7650 -1696 7651
rect -1662 7650 -1627 7651
rect -1593 7650 -1558 7651
rect -1933 7617 -1903 7650
rect -1859 7617 -1834 7650
rect -1785 7617 -1765 7650
rect -1711 7617 -1696 7650
rect -1637 7617 -1627 7650
rect -1563 7617 -1558 7650
rect -1524 7650 -1489 7651
rect -1524 7617 -1523 7650
rect -2007 7616 -1967 7617
rect -1933 7616 -1893 7617
rect -1859 7616 -1819 7617
rect -1785 7616 -1745 7617
rect -1711 7616 -1671 7617
rect -1637 7616 -1597 7617
rect -1563 7616 -1523 7617
rect -1455 7650 -1420 7651
rect -1386 7650 -1351 7651
rect -1317 7650 -1282 7651
rect -1248 7650 -1213 7651
rect -1179 7650 -1144 7651
rect -702 7650 -668 7672
rect -1455 7617 -1449 7650
rect -1386 7617 -1375 7650
rect -1317 7617 -1301 7650
rect -1248 7617 -1227 7650
rect -1179 7617 -1153 7650
rect -1489 7616 -1449 7617
rect -1415 7616 -1375 7617
rect -1341 7616 -1301 7617
rect -1267 7616 -1227 7617
rect -1193 7616 -1153 7617
rect -679 7638 -668 7650
rect -634 7638 -600 7672
rect -566 7638 -532 7672
rect -679 7616 -498 7638
rect -2119 7583 -1144 7616
rect -2119 7544 -2041 7583
rect -2007 7549 -1972 7583
rect -1938 7578 -1903 7583
rect -1869 7578 -1834 7583
rect -1800 7578 -1765 7583
rect -1731 7578 -1696 7583
rect -1662 7578 -1627 7583
rect -1593 7578 -1558 7583
rect -1933 7549 -1903 7578
rect -1859 7549 -1834 7578
rect -1785 7549 -1765 7578
rect -1711 7549 -1696 7578
rect -1637 7549 -1627 7578
rect -1563 7549 -1558 7578
rect -1524 7578 -1489 7583
rect -1524 7549 -1523 7578
rect -2007 7544 -1967 7549
rect -1933 7544 -1893 7549
rect -1859 7544 -1819 7549
rect -1785 7544 -1745 7549
rect -1711 7544 -1671 7549
rect -1637 7544 -1597 7549
rect -1563 7544 -1523 7549
rect -1455 7578 -1420 7583
rect -1386 7578 -1351 7583
rect -1317 7578 -1282 7583
rect -1248 7578 -1213 7583
rect -1179 7578 -1144 7583
rect -702 7603 -498 7616
rect -702 7578 -668 7603
rect -1455 7549 -1449 7578
rect -1386 7549 -1375 7578
rect -1317 7549 -1301 7578
rect -1248 7549 -1227 7578
rect -1179 7549 -1153 7578
rect -679 7569 -668 7578
rect -634 7569 -600 7603
rect -566 7569 -532 7603
rect -1489 7544 -1449 7549
rect -1415 7544 -1375 7549
rect -1341 7544 -1301 7549
rect -1267 7544 -1227 7549
rect -1193 7544 -1153 7549
rect -1119 7544 -1079 7549
rect -1045 7544 -1005 7549
rect -971 7544 -932 7549
rect -898 7544 -859 7549
rect -825 7544 -786 7549
rect -752 7544 -713 7549
rect -679 7544 -498 7569
rect -2119 7538 -498 7544
rect -668 7534 -498 7538
rect -634 7500 -600 7534
rect -566 7500 -532 7534
rect -668 7465 -498 7500
rect -634 7431 -600 7465
rect -566 7431 -532 7465
rect -668 7396 -498 7431
rect -634 7362 -600 7396
rect -566 7362 -532 7396
rect -668 7327 -498 7362
rect -634 7293 -600 7327
rect -566 7293 -532 7327
rect -668 7258 -498 7293
rect -634 7224 -600 7258
rect -566 7224 -532 7258
rect -668 7189 -498 7224
rect -634 7155 -600 7189
rect -566 7155 -532 7189
rect -668 7121 -498 7155
rect 19654 6118 19756 6134
rect 19688 6117 19722 6118
rect 21895 6118 21898 6134
rect 19688 6084 19693 6117
rect 19756 6084 19765 6117
rect 19654 6083 19693 6084
rect 19727 6083 19765 6084
rect 19654 6068 19756 6083
rect 21895 6068 21898 6084
rect 19663 5918 19765 5934
rect 19697 5884 19731 5918
rect 19663 5868 19765 5884
rect 21805 5918 21907 5934
rect 21839 5884 21873 5918
rect 21805 5868 21907 5884
rect 19654 5692 19756 5708
rect 19688 5658 19722 5692
rect 19654 5642 19756 5658
rect 21796 5692 21898 5708
rect 21830 5658 21864 5692
rect 21796 5642 21898 5658
rect 19697 5491 19799 5507
rect 19731 5457 19765 5491
rect 19727 5456 19765 5457
rect 19697 5441 19799 5456
rect 21878 5491 21941 5507
rect 21878 5457 21907 5491
rect 21878 5441 21941 5457
rect 19832 2978 19972 2980
rect -52 2928 48 2978
rect -1596 2920 -1340 2927
rect -1596 2886 -1580 2920
rect -1546 2886 -1485 2920
rect -1451 2886 -1390 2920
rect -1356 2886 -1340 2920
rect -1596 2879 -1340 2886
rect -1153 2920 -897 2927
rect -1153 2886 -1137 2920
rect -1103 2886 -1042 2920
rect -1008 2886 -947 2920
rect -913 2886 -897 2920
rect -1153 2879 -897 2886
rect -52 2894 -20 2928
rect 14 2894 48 2928
rect -1641 2823 -1607 2835
rect -1641 2751 -1607 2785
rect -1641 2683 -1607 2716
rect -1641 2615 -1607 2642
rect -1641 2547 -1607 2581
rect -1641 2479 -1607 2513
rect -1641 2411 -1607 2445
rect -1641 2343 -1607 2377
rect -1641 2293 -1607 2309
rect -1485 2819 -1451 2835
rect -1485 2751 -1451 2785
rect -1485 2683 -1451 2717
rect -1485 2615 -1451 2649
rect -1485 2561 -1451 2581
rect -1485 2489 -1451 2513
rect -1485 2411 -1451 2445
rect -1485 2343 -1451 2377
rect -1485 2293 -1451 2309
rect -1329 2823 -1295 2835
rect -1329 2751 -1295 2785
rect -1329 2683 -1295 2716
rect -1329 2615 -1295 2642
rect -1329 2547 -1295 2581
rect -1329 2479 -1295 2513
rect -1329 2411 -1295 2445
rect -1329 2343 -1295 2377
rect -1329 2293 -1295 2309
rect -1198 2823 -1164 2835
rect -1198 2751 -1164 2785
rect -1198 2683 -1164 2716
rect -1198 2615 -1164 2642
rect -1198 2547 -1164 2581
rect -1198 2479 -1164 2513
rect -1198 2411 -1164 2445
rect -1198 2343 -1164 2377
rect -1198 2293 -1164 2309
rect -1042 2819 -1008 2835
rect -1042 2751 -1008 2785
rect -1042 2683 -1008 2717
rect -1042 2615 -1008 2649
rect -1042 2547 -1008 2581
rect -1042 2479 -1008 2513
rect -1042 2411 -1008 2441
rect -1042 2343 -1008 2369
rect -1042 2293 -1008 2309
rect -886 2823 -852 2835
rect -886 2751 -852 2785
rect -886 2683 -852 2716
rect -886 2615 -852 2642
rect -886 2547 -852 2581
rect -886 2479 -852 2513
rect -886 2411 -852 2445
rect -886 2343 -852 2377
rect -886 2293 -852 2309
rect -52 2808 48 2894
rect 19938 2808 19972 2978
rect -52 2794 82 2808
rect -52 2760 -46 2794
rect -12 2774 42 2794
rect -12 2760 -2 2774
rect -52 2740 -2 2760
rect 32 2760 42 2774
rect 76 2760 82 2794
rect 32 2740 82 2760
rect -52 2721 82 2740
rect -52 2687 -46 2721
rect -12 2705 42 2721
rect -12 2687 -2 2705
rect -52 2671 -2 2687
rect 32 2687 42 2705
rect 76 2687 82 2721
rect 32 2671 82 2687
rect -52 2648 82 2671
rect -52 2614 -46 2648
rect -12 2636 42 2648
rect -12 2614 -2 2636
rect -52 2602 -2 2614
rect 32 2614 42 2636
rect 76 2614 82 2648
rect 32 2602 82 2614
rect -52 2575 82 2602
rect 19859 2800 19939 2808
rect 19859 2766 19882 2800
rect 19916 2766 19939 2800
rect 19859 2727 19939 2766
rect 19859 2693 19882 2727
rect 19916 2693 19939 2727
rect 19859 2654 19939 2693
rect 19859 2620 19882 2654
rect 19916 2620 19939 2654
rect 19859 2592 19939 2620
rect -52 2541 -46 2575
rect -12 2567 42 2575
rect -12 2541 -2 2567
rect -52 2533 -2 2541
rect 32 2541 42 2567
rect 76 2541 82 2575
rect 32 2533 82 2541
rect -52 2502 82 2533
rect -52 2468 -46 2502
rect -12 2498 42 2502
rect -12 2468 -2 2498
rect -52 2464 -2 2468
rect 32 2468 42 2498
rect 76 2468 82 2502
rect 32 2464 82 2468
rect -52 2429 82 2464
rect -52 2395 -46 2429
rect -12 2395 -2 2429
rect 32 2395 42 2429
rect 76 2395 82 2429
rect -52 2360 82 2395
rect -52 2356 -2 2360
rect -52 2322 -46 2356
rect -12 2326 -2 2356
rect 32 2356 82 2360
rect 32 2326 42 2356
rect -12 2322 42 2326
rect 76 2322 82 2356
rect -52 2291 82 2322
rect -52 2283 -2 2291
rect -52 2249 -46 2283
rect -12 2257 -2 2283
rect 32 2283 82 2291
rect 32 2257 42 2283
rect -12 2249 42 2257
rect 76 2249 82 2283
rect -52 2222 82 2249
rect -52 2210 -2 2222
rect -52 2176 -46 2210
rect -12 2188 -2 2210
rect 32 2210 82 2222
rect 32 2188 42 2210
rect -12 2176 42 2188
rect 76 2176 82 2210
rect -52 2153 82 2176
rect -52 2137 -2 2153
rect -1596 2114 -1340 2121
rect -1596 2080 -1584 2114
rect -1546 2080 -1503 2114
rect -1451 2080 -1423 2114
rect -1356 2080 -1343 2114
rect -1309 2080 -1263 2114
rect -1229 2080 -1183 2114
rect -1149 2080 -1103 2114
rect -1069 2080 -1023 2114
rect -989 2080 -943 2114
rect -52 2103 -46 2137
rect -12 2119 -2 2137
rect 32 2137 82 2153
rect 32 2119 42 2137
rect -12 2103 42 2119
rect 76 2103 82 2137
rect -52 2084 82 2103
rect -1596 2073 -1340 2080
rect -52 2064 -2 2084
rect -52 2030 -46 2064
rect -12 2050 -2 2064
rect 32 2064 82 2084
rect 32 2050 42 2064
rect -12 2030 42 2050
rect 76 2030 82 2064
rect -1641 1956 -1607 1979
rect -1641 1882 -1607 1911
rect -1641 1809 -1607 1843
rect -1641 1741 -1607 1775
rect -1641 1673 -1607 1707
rect -1641 1605 -1607 1639
rect -1641 1537 -1607 1571
rect -1641 1487 -1607 1503
rect -1485 2013 -1451 2029
rect -1485 1945 -1451 1979
rect -1485 1877 -1451 1911
rect -1485 1809 -1451 1843
rect -1485 1765 -1451 1775
rect -1485 1693 -1451 1707
rect -1485 1605 -1451 1639
rect -1485 1537 -1451 1571
rect -1485 1487 -1451 1503
rect -1329 1956 -1295 1979
rect -1329 1882 -1295 1911
rect -1329 1809 -1295 1843
rect -1329 1741 -1295 1775
rect -1329 1673 -1295 1707
rect -1329 1605 -1295 1639
rect -1329 1537 -1295 1571
rect -1329 1487 -1295 1503
rect -52 2015 82 2030
rect -52 1991 -2 2015
rect -52 1957 -46 1991
rect -12 1981 -2 1991
rect 32 1991 82 2015
rect 32 1981 42 1991
rect -12 1957 42 1981
rect 76 1957 82 1991
rect -52 1946 82 1957
rect -52 1918 -2 1946
rect -52 1884 -46 1918
rect -12 1912 -2 1918
rect 32 1918 82 1946
rect 32 1912 42 1918
rect -12 1884 42 1912
rect 76 1884 82 1918
rect -52 1877 82 1884
rect -52 1845 -2 1877
rect -52 1811 -46 1845
rect -12 1843 -2 1845
rect 32 1845 82 1877
rect 32 1843 42 1845
rect -12 1811 42 1843
rect 76 1811 82 1845
rect -52 1808 82 1811
rect -52 1774 -2 1808
rect 32 1774 82 1808
rect -52 1772 82 1774
rect -52 1738 -46 1772
rect -12 1739 42 1772
rect -12 1738 -2 1739
rect -52 1705 -2 1738
rect 32 1738 42 1739
rect 76 1738 82 1772
rect 32 1705 82 1738
rect -52 1699 82 1705
rect -52 1665 -46 1699
rect -12 1670 42 1699
rect -12 1665 -2 1670
rect -52 1636 -2 1665
rect 32 1665 42 1670
rect 76 1665 82 1699
rect 32 1636 82 1665
rect 19838 2581 19972 2592
rect 19838 2547 19882 2581
rect 19916 2558 19972 2581
rect 19838 2524 19888 2547
rect 19922 2524 19972 2558
rect 19838 2508 19972 2524
rect 19838 2474 19882 2508
rect 19916 2489 19972 2508
rect 19838 2455 19888 2474
rect 19922 2455 19972 2489
rect 19838 2435 19972 2455
rect 19838 2401 19882 2435
rect 19916 2420 19972 2435
rect 19838 2386 19888 2401
rect 19922 2386 19972 2420
rect 19838 2362 19972 2386
rect 19838 2328 19882 2362
rect 19916 2351 19972 2362
rect 19838 2317 19888 2328
rect 19922 2317 19972 2351
rect 19838 2289 19972 2317
rect 19838 2255 19882 2289
rect 19916 2282 19972 2289
rect 19838 2248 19888 2255
rect 19922 2248 19972 2282
rect 19838 2216 19972 2248
rect 19838 2182 19882 2216
rect 19916 2213 19972 2216
rect 19838 2179 19888 2182
rect 19922 2179 19972 2213
rect 19838 2144 19972 2179
rect 19838 2143 19888 2144
rect 19838 2109 19882 2143
rect 19922 2110 19972 2144
rect 19916 2109 19972 2110
rect 19838 2075 19972 2109
rect 19838 2070 19888 2075
rect 19838 2036 19882 2070
rect 19922 2041 19972 2075
rect 19916 2036 19972 2041
rect 19838 2006 19972 2036
rect 19838 1997 19888 2006
rect 19838 1963 19882 1997
rect 19922 1972 19972 2006
rect 19916 1963 19972 1972
rect 19838 1937 19972 1963
rect 19838 1924 19888 1937
rect 19838 1890 19882 1924
rect 19922 1903 19972 1937
rect 19916 1890 19972 1903
rect 19838 1868 19972 1890
rect 19838 1851 19888 1868
rect 19838 1817 19882 1851
rect 19922 1834 19972 1868
rect 19916 1817 19972 1834
rect 19838 1799 19972 1817
rect 19838 1778 19888 1799
rect 19838 1744 19882 1778
rect 19922 1765 19972 1799
rect 19916 1744 19972 1765
rect 19838 1730 19972 1744
rect 19838 1705 19888 1730
rect 19838 1671 19882 1705
rect 19922 1696 19972 1730
rect 19916 1671 19972 1696
rect 19838 1661 19972 1671
rect -52 1626 82 1636
rect -52 1592 -46 1626
rect -12 1601 42 1626
rect -12 1592 -2 1601
rect -52 1567 -2 1592
rect 32 1592 42 1601
rect 76 1592 82 1626
rect 32 1567 82 1592
rect -52 1553 82 1567
rect -52 1519 -46 1553
rect -12 1532 42 1553
rect -12 1519 -2 1532
rect -52 1498 -2 1519
rect 32 1519 42 1532
rect 76 1519 82 1553
rect 264 1534 364 1640
rect 398 1638 437 1640
rect 471 1638 510 1640
rect 544 1638 583 1640
rect 617 1638 656 1640
rect 690 1638 729 1640
rect 763 1638 802 1640
rect 836 1638 875 1640
rect 909 1638 948 1640
rect 982 1638 1021 1640
rect 1055 1638 1094 1640
rect 1128 1638 1167 1640
rect 1201 1638 1240 1640
rect 1274 1638 1313 1640
rect 1347 1638 1386 1640
rect 1420 1638 1459 1640
rect 1493 1638 1532 1640
rect 1566 1638 1605 1640
rect 1639 1638 1678 1640
rect 1712 1638 1751 1640
rect 1785 1638 1824 1640
rect 1858 1638 1898 1640
rect 1932 1638 1972 1640
rect 2006 1638 2046 1640
rect 2080 1638 2120 1640
rect 2154 1638 2194 1640
rect 2228 1638 2268 1640
rect 2302 1638 2342 1640
rect 2376 1638 2416 1640
rect 2450 1638 2490 1640
rect 2524 1638 2564 1640
rect 2598 1638 2638 1640
rect 2672 1638 2712 1640
rect 2598 1606 2609 1638
rect 2672 1606 2678 1638
rect 2574 1604 2609 1606
rect 2643 1604 2678 1606
rect 2746 1638 2786 1640
rect 2820 1638 2860 1640
rect 2894 1638 2934 1640
rect 2968 1638 3008 1640
rect 3042 1638 3082 1640
rect 3116 1638 3156 1640
rect 3190 1638 3230 1640
rect 2746 1606 2747 1638
rect 2712 1604 2747 1606
rect 2781 1606 2786 1638
rect 2850 1606 2860 1638
rect 2919 1606 2934 1638
rect 2988 1606 3008 1638
rect 3057 1606 3082 1638
rect 3126 1606 3156 1638
rect 2781 1604 2816 1606
rect 2850 1604 2885 1606
rect 2919 1604 2954 1606
rect 2988 1604 3023 1606
rect 3057 1604 3092 1606
rect 3126 1604 3161 1606
rect 3195 1604 3230 1638
rect 3264 1604 3364 1640
rect 2574 1570 3364 1604
rect 2574 1568 2609 1570
rect 2643 1568 2678 1570
rect 2598 1536 2609 1568
rect 2672 1536 2678 1568
rect 2712 1568 2747 1570
rect 398 1534 437 1536
rect 471 1534 510 1536
rect 544 1534 583 1536
rect 617 1534 656 1536
rect 690 1534 729 1536
rect 763 1534 802 1536
rect 836 1534 875 1536
rect 909 1534 948 1536
rect 982 1534 1021 1536
rect 1055 1534 1094 1536
rect 1128 1534 1167 1536
rect 1201 1534 1240 1536
rect 1274 1534 1313 1536
rect 1347 1534 1386 1536
rect 1420 1534 1459 1536
rect 1493 1534 1532 1536
rect 1566 1534 1605 1536
rect 1639 1534 1678 1536
rect 1712 1534 1751 1536
rect 1785 1534 1824 1536
rect 1858 1534 1898 1536
rect 1932 1534 1972 1536
rect 2006 1534 2046 1536
rect 2080 1534 2120 1536
rect 2154 1534 2194 1536
rect 2228 1534 2268 1536
rect 2302 1534 2342 1536
rect 2376 1534 2416 1536
rect 2450 1534 2490 1536
rect 2524 1534 2564 1536
rect 2598 1534 2638 1536
rect 2672 1534 2712 1536
rect 2746 1536 2747 1568
rect 2781 1568 2816 1570
rect 2850 1568 2885 1570
rect 2919 1568 2954 1570
rect 2988 1568 3023 1570
rect 3057 1568 3092 1570
rect 3126 1568 3161 1570
rect 2781 1536 2786 1568
rect 2850 1536 2860 1568
rect 2919 1536 2934 1568
rect 2988 1536 3008 1568
rect 3057 1536 3082 1568
rect 3126 1536 3156 1568
rect 3195 1536 3230 1570
rect 2746 1534 2786 1536
rect 2820 1534 2860 1536
rect 2894 1534 2934 1536
rect 2968 1534 3008 1536
rect 3042 1534 3082 1536
rect 3116 1534 3156 1536
rect 3190 1534 3230 1536
rect 3264 1534 3364 1570
rect 3506 1604 3606 1640
rect 3640 1638 3680 1640
rect 3714 1638 3754 1640
rect 3788 1638 3828 1640
rect 3862 1638 3902 1640
rect 3936 1638 3976 1640
rect 4010 1638 4050 1640
rect 4084 1638 4124 1640
rect 3640 1604 3675 1638
rect 3714 1606 3744 1638
rect 3788 1606 3813 1638
rect 3862 1606 3882 1638
rect 3936 1606 3951 1638
rect 4010 1606 4020 1638
rect 4084 1606 4089 1638
rect 3709 1604 3744 1606
rect 3778 1604 3813 1606
rect 3847 1604 3882 1606
rect 3916 1604 3951 1606
rect 3985 1604 4020 1606
rect 4054 1604 4089 1606
rect 4123 1606 4124 1638
rect 4158 1638 4198 1640
rect 4232 1638 4272 1640
rect 4306 1638 4346 1640
rect 4380 1638 4420 1640
rect 4454 1638 4494 1640
rect 4528 1638 4568 1640
rect 4602 1638 4642 1640
rect 4676 1638 4716 1640
rect 4750 1638 4790 1640
rect 4824 1638 4864 1640
rect 4898 1638 4938 1640
rect 4972 1638 5012 1640
rect 5046 1638 5085 1640
rect 5119 1638 5158 1640
rect 5192 1638 5231 1640
rect 5265 1638 5304 1640
rect 5338 1638 5377 1640
rect 5411 1638 5450 1640
rect 5484 1638 5523 1640
rect 5557 1638 5596 1640
rect 5630 1638 5669 1640
rect 5703 1638 5742 1640
rect 5776 1638 5815 1640
rect 5849 1638 5888 1640
rect 5922 1638 5961 1640
rect 5995 1638 6034 1640
rect 6068 1638 6107 1640
rect 6141 1638 6180 1640
rect 6214 1638 6253 1640
rect 6287 1638 6326 1640
rect 6360 1638 6399 1640
rect 6433 1638 6472 1640
rect 4123 1604 4158 1606
rect 4192 1606 4198 1638
rect 4261 1606 4272 1638
rect 4192 1604 4227 1606
rect 4261 1604 4296 1606
rect 3506 1570 4296 1604
rect 3506 1534 3606 1570
rect 3640 1536 3675 1570
rect 3709 1568 3744 1570
rect 3778 1568 3813 1570
rect 3847 1568 3882 1570
rect 3916 1568 3951 1570
rect 3985 1568 4020 1570
rect 4054 1568 4089 1570
rect 3714 1536 3744 1568
rect 3788 1536 3813 1568
rect 3862 1536 3882 1568
rect 3936 1536 3951 1568
rect 4010 1536 4020 1568
rect 4084 1536 4089 1568
rect 4123 1568 4158 1570
rect 4123 1536 4124 1568
rect 3640 1534 3680 1536
rect 3714 1534 3754 1536
rect 3788 1534 3828 1536
rect 3862 1534 3902 1536
rect 3936 1534 3976 1536
rect 4010 1534 4050 1536
rect 4084 1534 4124 1536
rect 4192 1568 4227 1570
rect 4261 1568 4296 1570
rect 4192 1536 4198 1568
rect 4261 1536 4272 1568
rect 4158 1534 4198 1536
rect 4232 1534 4272 1536
rect 4306 1534 4346 1536
rect 4380 1534 4420 1536
rect 4454 1534 4494 1536
rect 4528 1534 4568 1536
rect 4602 1534 4642 1536
rect 4676 1534 4716 1536
rect 4750 1534 4790 1536
rect 4824 1534 4864 1536
rect 4898 1534 4938 1536
rect 4972 1534 5012 1536
rect 5046 1534 5085 1536
rect 5119 1534 5158 1536
rect 5192 1534 5231 1536
rect 5265 1534 5304 1536
rect 5338 1534 5377 1536
rect 5411 1534 5450 1536
rect 5484 1534 5523 1536
rect 5557 1534 5596 1536
rect 5630 1534 5669 1536
rect 5703 1534 5742 1536
rect 5776 1534 5815 1536
rect 5849 1534 5888 1536
rect 5922 1534 5961 1536
rect 5995 1534 6034 1536
rect 6068 1534 6107 1536
rect 6141 1534 6180 1536
rect 6214 1534 6253 1536
rect 6287 1534 6326 1536
rect 6360 1534 6399 1536
rect 6433 1534 6472 1536
rect 6506 1534 6606 1640
rect 6748 1534 6848 1640
rect 6882 1638 6921 1640
rect 6955 1638 6994 1640
rect 7028 1638 7067 1640
rect 7101 1638 7140 1640
rect 7174 1638 7213 1640
rect 7247 1638 7286 1640
rect 7320 1638 7359 1640
rect 7393 1638 7432 1640
rect 7466 1638 7505 1640
rect 7539 1638 7578 1640
rect 7612 1638 7651 1640
rect 7685 1638 7724 1640
rect 7758 1638 7797 1640
rect 7831 1638 7870 1640
rect 7904 1638 7943 1640
rect 7977 1638 8016 1640
rect 8050 1638 8089 1640
rect 8123 1638 8162 1640
rect 8196 1638 8235 1640
rect 8269 1638 8308 1640
rect 8342 1638 8382 1640
rect 8416 1638 8456 1640
rect 8490 1638 8530 1640
rect 8564 1638 8604 1640
rect 8638 1638 8678 1640
rect 8712 1638 8752 1640
rect 8786 1638 8826 1640
rect 8860 1638 8900 1640
rect 8934 1638 8974 1640
rect 9008 1638 9048 1640
rect 9082 1638 9122 1640
rect 9156 1638 9196 1640
rect 9082 1606 9093 1638
rect 9156 1606 9162 1638
rect 9058 1604 9093 1606
rect 9127 1604 9162 1606
rect 9230 1638 9270 1640
rect 9304 1638 9344 1640
rect 9378 1638 9418 1640
rect 9452 1638 9492 1640
rect 9526 1638 9566 1640
rect 9600 1638 9640 1640
rect 9674 1638 9714 1640
rect 9230 1606 9231 1638
rect 9196 1604 9231 1606
rect 9265 1606 9270 1638
rect 9334 1606 9344 1638
rect 9403 1606 9418 1638
rect 9472 1606 9492 1638
rect 9541 1606 9566 1638
rect 9610 1606 9640 1638
rect 9265 1604 9300 1606
rect 9334 1604 9369 1606
rect 9403 1604 9438 1606
rect 9472 1604 9507 1606
rect 9541 1604 9576 1606
rect 9610 1604 9645 1606
rect 9679 1604 9714 1638
rect 9748 1604 9848 1640
rect 9058 1570 9848 1604
rect 9058 1568 9093 1570
rect 9127 1568 9162 1570
rect 9082 1536 9093 1568
rect 9156 1536 9162 1568
rect 9196 1568 9231 1570
rect 6882 1534 6921 1536
rect 6955 1534 6994 1536
rect 7028 1534 7067 1536
rect 7101 1534 7140 1536
rect 7174 1534 7213 1536
rect 7247 1534 7286 1536
rect 7320 1534 7359 1536
rect 7393 1534 7432 1536
rect 7466 1534 7505 1536
rect 7539 1534 7578 1536
rect 7612 1534 7651 1536
rect 7685 1534 7724 1536
rect 7758 1534 7797 1536
rect 7831 1534 7870 1536
rect 7904 1534 7943 1536
rect 7977 1534 8016 1536
rect 8050 1534 8089 1536
rect 8123 1534 8162 1536
rect 8196 1534 8235 1536
rect 8269 1534 8308 1536
rect 8342 1534 8382 1536
rect 8416 1534 8456 1536
rect 8490 1534 8530 1536
rect 8564 1534 8604 1536
rect 8638 1534 8678 1536
rect 8712 1534 8752 1536
rect 8786 1534 8826 1536
rect 8860 1534 8900 1536
rect 8934 1534 8974 1536
rect 9008 1534 9048 1536
rect 9082 1534 9122 1536
rect 9156 1534 9196 1536
rect 9230 1536 9231 1568
rect 9265 1568 9300 1570
rect 9334 1568 9369 1570
rect 9403 1568 9438 1570
rect 9472 1568 9507 1570
rect 9541 1568 9576 1570
rect 9610 1568 9645 1570
rect 9265 1536 9270 1568
rect 9334 1536 9344 1568
rect 9403 1536 9418 1568
rect 9472 1536 9492 1568
rect 9541 1536 9566 1568
rect 9610 1536 9640 1568
rect 9679 1536 9714 1570
rect 9230 1534 9270 1536
rect 9304 1534 9344 1536
rect 9378 1534 9418 1536
rect 9452 1534 9492 1536
rect 9526 1534 9566 1536
rect 9600 1534 9640 1536
rect 9674 1534 9714 1536
rect 9748 1534 9848 1570
rect 9990 1604 10090 1640
rect 10124 1638 10164 1640
rect 10198 1638 10238 1640
rect 10272 1638 10312 1640
rect 10346 1638 10386 1640
rect 10420 1638 10460 1640
rect 10494 1638 10534 1640
rect 10568 1638 10608 1640
rect 10124 1604 10159 1638
rect 10198 1606 10228 1638
rect 10272 1606 10297 1638
rect 10346 1606 10366 1638
rect 10420 1606 10435 1638
rect 10494 1606 10504 1638
rect 10568 1606 10573 1638
rect 10193 1604 10228 1606
rect 10262 1604 10297 1606
rect 10331 1604 10366 1606
rect 10400 1604 10435 1606
rect 10469 1604 10504 1606
rect 10538 1604 10573 1606
rect 10607 1606 10608 1638
rect 10642 1638 10682 1640
rect 10716 1638 10756 1640
rect 10790 1638 10830 1640
rect 10864 1638 10904 1640
rect 10938 1638 10978 1640
rect 11012 1638 11052 1640
rect 11086 1638 11126 1640
rect 11160 1638 11200 1640
rect 11234 1638 11274 1640
rect 11308 1638 11348 1640
rect 11382 1638 11422 1640
rect 11456 1638 11496 1640
rect 11530 1638 11569 1640
rect 11603 1638 11642 1640
rect 11676 1638 11715 1640
rect 11749 1638 11788 1640
rect 11822 1638 11861 1640
rect 11895 1638 11934 1640
rect 11968 1638 12007 1640
rect 12041 1638 12080 1640
rect 12114 1638 12153 1640
rect 12187 1638 12226 1640
rect 12260 1638 12299 1640
rect 12333 1638 12372 1640
rect 12406 1638 12445 1640
rect 12479 1638 12518 1640
rect 12552 1638 12591 1640
rect 12625 1638 12664 1640
rect 12698 1638 12737 1640
rect 12771 1638 12810 1640
rect 12844 1638 12883 1640
rect 12917 1638 12956 1640
rect 10607 1604 10642 1606
rect 10676 1606 10682 1638
rect 10745 1606 10756 1638
rect 10676 1604 10711 1606
rect 10745 1604 10780 1606
rect 9990 1570 10780 1604
rect 9990 1534 10090 1570
rect 10124 1536 10159 1570
rect 10193 1568 10228 1570
rect 10262 1568 10297 1570
rect 10331 1568 10366 1570
rect 10400 1568 10435 1570
rect 10469 1568 10504 1570
rect 10538 1568 10573 1570
rect 10198 1536 10228 1568
rect 10272 1536 10297 1568
rect 10346 1536 10366 1568
rect 10420 1536 10435 1568
rect 10494 1536 10504 1568
rect 10568 1536 10573 1568
rect 10607 1568 10642 1570
rect 10607 1536 10608 1568
rect 10124 1534 10164 1536
rect 10198 1534 10238 1536
rect 10272 1534 10312 1536
rect 10346 1534 10386 1536
rect 10420 1534 10460 1536
rect 10494 1534 10534 1536
rect 10568 1534 10608 1536
rect 10676 1568 10711 1570
rect 10745 1568 10780 1570
rect 10676 1536 10682 1568
rect 10745 1536 10756 1568
rect 10642 1534 10682 1536
rect 10716 1534 10756 1536
rect 10790 1534 10830 1536
rect 10864 1534 10904 1536
rect 10938 1534 10978 1536
rect 11012 1534 11052 1536
rect 11086 1534 11126 1536
rect 11160 1534 11200 1536
rect 11234 1534 11274 1536
rect 11308 1534 11348 1536
rect 11382 1534 11422 1536
rect 11456 1534 11496 1536
rect 11530 1534 11569 1536
rect 11603 1534 11642 1536
rect 11676 1534 11715 1536
rect 11749 1534 11788 1536
rect 11822 1534 11861 1536
rect 11895 1534 11934 1536
rect 11968 1534 12007 1536
rect 12041 1534 12080 1536
rect 12114 1534 12153 1536
rect 12187 1534 12226 1536
rect 12260 1534 12299 1536
rect 12333 1534 12372 1536
rect 12406 1534 12445 1536
rect 12479 1534 12518 1536
rect 12552 1534 12591 1536
rect 12625 1534 12664 1536
rect 12698 1534 12737 1536
rect 12771 1534 12810 1536
rect 12844 1534 12883 1536
rect 12917 1534 12956 1536
rect 12990 1534 13090 1640
rect 13232 1534 13332 1640
rect 13366 1638 13405 1640
rect 13439 1638 13478 1640
rect 13512 1638 13551 1640
rect 13585 1638 13624 1640
rect 13658 1638 13697 1640
rect 13731 1638 13770 1640
rect 13804 1638 13843 1640
rect 13877 1638 13916 1640
rect 13950 1638 13989 1640
rect 14023 1638 14062 1640
rect 14096 1638 14135 1640
rect 14169 1638 14208 1640
rect 14242 1638 14281 1640
rect 14315 1638 14354 1640
rect 14388 1638 14427 1640
rect 14461 1638 14500 1640
rect 14534 1638 14573 1640
rect 14607 1638 14646 1640
rect 14680 1638 14719 1640
rect 14753 1638 14792 1640
rect 14826 1638 14866 1640
rect 14900 1638 14940 1640
rect 14974 1638 15014 1640
rect 15048 1638 15088 1640
rect 15122 1638 15162 1640
rect 15196 1638 15236 1640
rect 15270 1638 15310 1640
rect 15344 1638 15384 1640
rect 15418 1638 15458 1640
rect 15492 1638 15532 1640
rect 15566 1638 15606 1640
rect 15640 1638 15680 1640
rect 15566 1606 15577 1638
rect 15640 1606 15646 1638
rect 15542 1604 15577 1606
rect 15611 1604 15646 1606
rect 15714 1638 15754 1640
rect 15788 1638 15828 1640
rect 15862 1638 15902 1640
rect 15936 1638 15976 1640
rect 16010 1638 16050 1640
rect 16084 1638 16124 1640
rect 16158 1638 16198 1640
rect 15714 1606 15715 1638
rect 15680 1604 15715 1606
rect 15749 1606 15754 1638
rect 15818 1606 15828 1638
rect 15887 1606 15902 1638
rect 15956 1606 15976 1638
rect 16025 1606 16050 1638
rect 16094 1606 16124 1638
rect 15749 1604 15784 1606
rect 15818 1604 15853 1606
rect 15887 1604 15922 1606
rect 15956 1604 15991 1606
rect 16025 1604 16060 1606
rect 16094 1604 16129 1606
rect 16163 1604 16198 1638
rect 16232 1604 16332 1640
rect 15542 1570 16332 1604
rect 15542 1568 15577 1570
rect 15611 1568 15646 1570
rect 15566 1536 15577 1568
rect 15640 1536 15646 1568
rect 15680 1568 15715 1570
rect 13366 1534 13405 1536
rect 13439 1534 13478 1536
rect 13512 1534 13551 1536
rect 13585 1534 13624 1536
rect 13658 1534 13697 1536
rect 13731 1534 13770 1536
rect 13804 1534 13843 1536
rect 13877 1534 13916 1536
rect 13950 1534 13989 1536
rect 14023 1534 14062 1536
rect 14096 1534 14135 1536
rect 14169 1534 14208 1536
rect 14242 1534 14281 1536
rect 14315 1534 14354 1536
rect 14388 1534 14427 1536
rect 14461 1534 14500 1536
rect 14534 1534 14573 1536
rect 14607 1534 14646 1536
rect 14680 1534 14719 1536
rect 14753 1534 14792 1536
rect 14826 1534 14866 1536
rect 14900 1534 14940 1536
rect 14974 1534 15014 1536
rect 15048 1534 15088 1536
rect 15122 1534 15162 1536
rect 15196 1534 15236 1536
rect 15270 1534 15310 1536
rect 15344 1534 15384 1536
rect 15418 1534 15458 1536
rect 15492 1534 15532 1536
rect 15566 1534 15606 1536
rect 15640 1534 15680 1536
rect 15714 1536 15715 1568
rect 15749 1568 15784 1570
rect 15818 1568 15853 1570
rect 15887 1568 15922 1570
rect 15956 1568 15991 1570
rect 16025 1568 16060 1570
rect 16094 1568 16129 1570
rect 15749 1536 15754 1568
rect 15818 1536 15828 1568
rect 15887 1536 15902 1568
rect 15956 1536 15976 1568
rect 16025 1536 16050 1568
rect 16094 1536 16124 1568
rect 16163 1536 16198 1570
rect 15714 1534 15754 1536
rect 15788 1534 15828 1536
rect 15862 1534 15902 1536
rect 15936 1534 15976 1536
rect 16010 1534 16050 1536
rect 16084 1534 16124 1536
rect 16158 1534 16198 1536
rect 16232 1534 16332 1570
rect 16474 1604 16574 1640
rect 16608 1638 16648 1640
rect 16682 1638 16722 1640
rect 16756 1638 16796 1640
rect 16830 1638 16870 1640
rect 16904 1638 16944 1640
rect 16978 1638 17018 1640
rect 17052 1638 17092 1640
rect 16608 1604 16643 1638
rect 16682 1606 16712 1638
rect 16756 1606 16781 1638
rect 16830 1606 16850 1638
rect 16904 1606 16919 1638
rect 16978 1606 16988 1638
rect 17052 1606 17057 1638
rect 16677 1604 16712 1606
rect 16746 1604 16781 1606
rect 16815 1604 16850 1606
rect 16884 1604 16919 1606
rect 16953 1604 16988 1606
rect 17022 1604 17057 1606
rect 17091 1606 17092 1638
rect 17126 1638 17166 1640
rect 17200 1638 17240 1640
rect 17274 1638 17314 1640
rect 17348 1638 17388 1640
rect 17422 1638 17462 1640
rect 17496 1638 17536 1640
rect 17570 1638 17610 1640
rect 17644 1638 17684 1640
rect 17718 1638 17758 1640
rect 17792 1638 17832 1640
rect 17866 1638 17906 1640
rect 17940 1638 17980 1640
rect 18014 1638 18053 1640
rect 18087 1638 18126 1640
rect 18160 1638 18199 1640
rect 18233 1638 18272 1640
rect 18306 1638 18345 1640
rect 18379 1638 18418 1640
rect 18452 1638 18491 1640
rect 18525 1638 18564 1640
rect 18598 1638 18637 1640
rect 18671 1638 18710 1640
rect 18744 1638 18783 1640
rect 18817 1638 18856 1640
rect 18890 1638 18929 1640
rect 18963 1638 19002 1640
rect 19036 1638 19075 1640
rect 19109 1638 19148 1640
rect 19182 1638 19221 1640
rect 19255 1638 19294 1640
rect 19328 1638 19367 1640
rect 19401 1638 19440 1640
rect 17091 1604 17126 1606
rect 17160 1606 17166 1638
rect 17229 1606 17240 1638
rect 17160 1604 17195 1606
rect 17229 1604 17264 1606
rect 16474 1570 17264 1604
rect 16474 1534 16574 1570
rect 16608 1536 16643 1570
rect 16677 1568 16712 1570
rect 16746 1568 16781 1570
rect 16815 1568 16850 1570
rect 16884 1568 16919 1570
rect 16953 1568 16988 1570
rect 17022 1568 17057 1570
rect 16682 1536 16712 1568
rect 16756 1536 16781 1568
rect 16830 1536 16850 1568
rect 16904 1536 16919 1568
rect 16978 1536 16988 1568
rect 17052 1536 17057 1568
rect 17091 1568 17126 1570
rect 17091 1536 17092 1568
rect 16608 1534 16648 1536
rect 16682 1534 16722 1536
rect 16756 1534 16796 1536
rect 16830 1534 16870 1536
rect 16904 1534 16944 1536
rect 16978 1534 17018 1536
rect 17052 1534 17092 1536
rect 17160 1568 17195 1570
rect 17229 1568 17264 1570
rect 17160 1536 17166 1568
rect 17229 1536 17240 1568
rect 17126 1534 17166 1536
rect 17200 1534 17240 1536
rect 17274 1534 17314 1536
rect 17348 1534 17388 1536
rect 17422 1534 17462 1536
rect 17496 1534 17536 1536
rect 17570 1534 17610 1536
rect 17644 1534 17684 1536
rect 17718 1534 17758 1536
rect 17792 1534 17832 1536
rect 17866 1534 17906 1536
rect 17940 1534 17980 1536
rect 18014 1534 18053 1536
rect 18087 1534 18126 1536
rect 18160 1534 18199 1536
rect 18233 1534 18272 1536
rect 18306 1534 18345 1536
rect 18379 1534 18418 1536
rect 18452 1534 18491 1536
rect 18525 1534 18564 1536
rect 18598 1534 18637 1536
rect 18671 1534 18710 1536
rect 18744 1534 18783 1536
rect 18817 1534 18856 1536
rect 18890 1534 18929 1536
rect 18963 1534 19002 1536
rect 19036 1534 19075 1536
rect 19109 1534 19148 1536
rect 19182 1534 19221 1536
rect 19255 1534 19294 1536
rect 19328 1534 19367 1536
rect 19401 1534 19440 1536
rect 19474 1534 19574 1640
rect 19838 1632 19888 1661
rect 19838 1598 19882 1632
rect 19922 1627 19972 1661
rect 19916 1598 19972 1627
rect 19838 1592 19972 1598
rect 19838 1559 19888 1592
rect 32 1498 82 1519
rect -52 1479 82 1498
rect -52 1445 -46 1479
rect -12 1463 42 1479
rect -12 1445 -2 1463
rect -52 1429 -2 1445
rect 32 1445 42 1463
rect 76 1445 82 1479
rect 19838 1525 19882 1559
rect 19922 1558 19972 1592
rect 19916 1525 19972 1558
rect 19838 1523 19972 1525
rect 19838 1489 19888 1523
rect 19922 1489 19972 1523
rect 19838 1486 19972 1489
rect 19838 1452 19882 1486
rect 19916 1454 19972 1486
rect 182 1446 216 1448
rect 3423 1446 3457 1448
rect 9907 1446 9941 1448
rect 16392 1446 16426 1448
rect 19622 1446 19656 1448
rect 32 1429 82 1445
rect -52 1405 82 1429
rect 202 1432 240 1446
rect 216 1412 240 1432
rect 3420 1432 3458 1446
rect 3420 1412 3423 1432
rect -52 1371 -46 1405
rect -12 1393 42 1405
rect -12 1371 -2 1393
rect -52 1359 -2 1371
rect 32 1371 42 1393
rect 76 1371 82 1405
rect 32 1359 82 1371
rect -52 1331 82 1359
rect -52 1297 -46 1331
rect -12 1323 42 1331
rect -12 1297 -2 1323
rect -52 1289 -2 1297
rect 32 1297 42 1323
rect 76 1297 82 1331
rect 182 1364 216 1398
rect 182 1314 216 1330
rect 3457 1412 3458 1432
rect 9904 1432 9942 1446
rect 9904 1412 9907 1432
rect 3423 1364 3457 1398
rect 3423 1314 3457 1330
rect 9941 1412 9942 1432
rect 16388 1432 16426 1446
rect 16388 1412 16392 1432
rect 9907 1364 9941 1398
rect 9907 1314 9941 1330
rect 19598 1432 19636 1446
rect 19598 1412 19622 1432
rect 19838 1420 19888 1452
rect 19922 1420 19972 1454
rect 19838 1413 19972 1420
rect 16392 1364 16426 1398
rect 16392 1314 16426 1330
rect 19622 1364 19656 1398
rect 19622 1314 19656 1330
rect 19838 1379 19882 1413
rect 19916 1385 19972 1413
rect 19838 1351 19888 1379
rect 19922 1351 19972 1385
rect 19838 1340 19972 1351
rect 32 1289 82 1297
rect -52 1257 82 1289
rect -52 1223 -46 1257
rect -12 1253 42 1257
rect -12 1223 -2 1253
rect -52 1219 -2 1223
rect 32 1223 42 1253
rect 76 1223 82 1257
rect 19838 1306 19882 1340
rect 19916 1316 19972 1340
rect 19838 1282 19888 1306
rect 19922 1282 19972 1316
rect 19838 1267 19972 1282
rect 19838 1233 19882 1267
rect 19916 1247 19972 1267
rect 32 1219 82 1223
rect -52 1183 82 1219
rect -52 1149 -46 1183
rect -12 1149 -2 1183
rect 32 1149 42 1183
rect 76 1149 82 1183
rect -52 1113 82 1149
rect 264 1122 364 1228
rect 398 1226 437 1228
rect 471 1226 510 1228
rect 544 1226 583 1228
rect 617 1226 656 1228
rect 690 1226 729 1228
rect 763 1226 802 1228
rect 836 1226 875 1228
rect 909 1226 948 1228
rect 982 1226 1021 1228
rect 1055 1226 1094 1228
rect 1128 1226 1167 1228
rect 1201 1226 1240 1228
rect 1274 1226 1313 1228
rect 1347 1226 1386 1228
rect 1420 1226 1459 1228
rect 1493 1226 1532 1228
rect 1566 1226 1605 1228
rect 1639 1226 1678 1228
rect 1712 1226 1751 1228
rect 1785 1226 1824 1228
rect 1858 1226 1898 1228
rect 1932 1226 1972 1228
rect 2006 1226 2046 1228
rect 2080 1226 2120 1228
rect 2154 1226 2194 1228
rect 2228 1226 2268 1228
rect 2302 1226 2342 1228
rect 2376 1226 2416 1228
rect 2450 1226 2490 1228
rect 2524 1226 2564 1228
rect 2598 1226 2638 1228
rect 2672 1226 2712 1228
rect 2598 1194 2609 1226
rect 2672 1194 2678 1226
rect 2574 1192 2609 1194
rect 2643 1192 2678 1194
rect 2746 1226 2786 1228
rect 2820 1226 2860 1228
rect 2894 1226 2934 1228
rect 2968 1226 3008 1228
rect 3042 1226 3082 1228
rect 3116 1226 3156 1228
rect 3190 1226 3230 1228
rect 2746 1194 2747 1226
rect 2712 1192 2747 1194
rect 2781 1194 2786 1226
rect 2850 1194 2860 1226
rect 2919 1194 2934 1226
rect 2988 1194 3008 1226
rect 3057 1194 3082 1226
rect 3126 1194 3156 1226
rect 2781 1192 2816 1194
rect 2850 1192 2885 1194
rect 2919 1192 2954 1194
rect 2988 1192 3023 1194
rect 3057 1192 3092 1194
rect 3126 1192 3161 1194
rect 3195 1192 3230 1226
rect 3264 1192 3364 1228
rect 2574 1158 3364 1192
rect 2574 1156 2609 1158
rect 2643 1156 2678 1158
rect 2598 1124 2609 1156
rect 2672 1124 2678 1156
rect 2712 1156 2747 1158
rect 398 1122 437 1124
rect 471 1122 510 1124
rect 544 1122 583 1124
rect 617 1122 656 1124
rect 690 1122 729 1124
rect 763 1122 802 1124
rect 836 1122 875 1124
rect 909 1122 948 1124
rect 982 1122 1021 1124
rect 1055 1122 1094 1124
rect 1128 1122 1167 1124
rect 1201 1122 1240 1124
rect 1274 1122 1313 1124
rect 1347 1122 1386 1124
rect 1420 1122 1459 1124
rect 1493 1122 1532 1124
rect 1566 1122 1605 1124
rect 1639 1122 1678 1124
rect 1712 1122 1751 1124
rect 1785 1122 1824 1124
rect 1858 1122 1898 1124
rect 1932 1122 1972 1124
rect 2006 1122 2046 1124
rect 2080 1122 2120 1124
rect 2154 1122 2194 1124
rect 2228 1122 2268 1124
rect 2302 1122 2342 1124
rect 2376 1122 2416 1124
rect 2450 1122 2490 1124
rect 2524 1122 2564 1124
rect 2598 1122 2638 1124
rect 2672 1122 2712 1124
rect 2746 1124 2747 1156
rect 2781 1156 2816 1158
rect 2850 1156 2885 1158
rect 2919 1156 2954 1158
rect 2988 1156 3023 1158
rect 3057 1156 3092 1158
rect 3126 1156 3161 1158
rect 2781 1124 2786 1156
rect 2850 1124 2860 1156
rect 2919 1124 2934 1156
rect 2988 1124 3008 1156
rect 3057 1124 3082 1156
rect 3126 1124 3156 1156
rect 3195 1124 3230 1158
rect 2746 1122 2786 1124
rect 2820 1122 2860 1124
rect 2894 1122 2934 1124
rect 2968 1122 3008 1124
rect 3042 1122 3082 1124
rect 3116 1122 3156 1124
rect 3190 1122 3230 1124
rect 3264 1122 3364 1158
rect 3506 1192 3606 1228
rect 3640 1226 3680 1228
rect 3714 1226 3754 1228
rect 3788 1226 3828 1228
rect 3862 1226 3902 1228
rect 3936 1226 3976 1228
rect 4010 1226 4050 1228
rect 4084 1226 4124 1228
rect 3640 1192 3675 1226
rect 3714 1194 3744 1226
rect 3788 1194 3813 1226
rect 3862 1194 3882 1226
rect 3936 1194 3951 1226
rect 4010 1194 4020 1226
rect 4084 1194 4089 1226
rect 3709 1192 3744 1194
rect 3778 1192 3813 1194
rect 3847 1192 3882 1194
rect 3916 1192 3951 1194
rect 3985 1192 4020 1194
rect 4054 1192 4089 1194
rect 4123 1194 4124 1226
rect 4158 1226 4198 1228
rect 4232 1226 4272 1228
rect 4306 1226 4346 1228
rect 4380 1226 4420 1228
rect 4454 1226 4494 1228
rect 4528 1226 4568 1228
rect 4602 1226 4642 1228
rect 4676 1226 4716 1228
rect 4750 1226 4790 1228
rect 4824 1226 4864 1228
rect 4898 1226 4938 1228
rect 4972 1226 5012 1228
rect 5046 1226 5085 1228
rect 5119 1226 5158 1228
rect 5192 1226 5231 1228
rect 5265 1226 5304 1228
rect 5338 1226 5377 1228
rect 5411 1226 5450 1228
rect 5484 1226 5523 1228
rect 5557 1226 5596 1228
rect 5630 1226 5669 1228
rect 5703 1226 5742 1228
rect 5776 1226 5815 1228
rect 5849 1226 5888 1228
rect 5922 1226 5961 1228
rect 5995 1226 6034 1228
rect 6068 1226 6107 1228
rect 6141 1226 6180 1228
rect 6214 1226 6253 1228
rect 6287 1226 6326 1228
rect 6360 1226 6399 1228
rect 6433 1226 6472 1228
rect 4123 1192 4158 1194
rect 4192 1194 4198 1226
rect 4261 1194 4272 1226
rect 4192 1192 4227 1194
rect 4261 1192 4296 1194
rect 3506 1158 4296 1192
rect 3506 1122 3606 1158
rect 3640 1124 3675 1158
rect 3709 1156 3744 1158
rect 3778 1156 3813 1158
rect 3847 1156 3882 1158
rect 3916 1156 3951 1158
rect 3985 1156 4020 1158
rect 4054 1156 4089 1158
rect 3714 1124 3744 1156
rect 3788 1124 3813 1156
rect 3862 1124 3882 1156
rect 3936 1124 3951 1156
rect 4010 1124 4020 1156
rect 4084 1124 4089 1156
rect 4123 1156 4158 1158
rect 4123 1124 4124 1156
rect 3640 1122 3680 1124
rect 3714 1122 3754 1124
rect 3788 1122 3828 1124
rect 3862 1122 3902 1124
rect 3936 1122 3976 1124
rect 4010 1122 4050 1124
rect 4084 1122 4124 1124
rect 4192 1156 4227 1158
rect 4261 1156 4296 1158
rect 4192 1124 4198 1156
rect 4261 1124 4272 1156
rect 4158 1122 4198 1124
rect 4232 1122 4272 1124
rect 4306 1122 4346 1124
rect 4380 1122 4420 1124
rect 4454 1122 4494 1124
rect 4528 1122 4568 1124
rect 4602 1122 4642 1124
rect 4676 1122 4716 1124
rect 4750 1122 4790 1124
rect 4824 1122 4864 1124
rect 4898 1122 4938 1124
rect 4972 1122 5012 1124
rect 5046 1122 5085 1124
rect 5119 1122 5158 1124
rect 5192 1122 5231 1124
rect 5265 1122 5304 1124
rect 5338 1122 5377 1124
rect 5411 1122 5450 1124
rect 5484 1122 5523 1124
rect 5557 1122 5596 1124
rect 5630 1122 5669 1124
rect 5703 1122 5742 1124
rect 5776 1122 5815 1124
rect 5849 1122 5888 1124
rect 5922 1122 5961 1124
rect 5995 1122 6034 1124
rect 6068 1122 6107 1124
rect 6141 1122 6180 1124
rect 6214 1122 6253 1124
rect 6287 1122 6326 1124
rect 6360 1122 6399 1124
rect 6433 1122 6472 1124
rect 6506 1122 6606 1228
rect 6748 1122 6848 1228
rect 6882 1226 6921 1228
rect 6955 1226 6994 1228
rect 7028 1226 7067 1228
rect 7101 1226 7140 1228
rect 7174 1226 7213 1228
rect 7247 1226 7286 1228
rect 7320 1226 7359 1228
rect 7393 1226 7432 1228
rect 7466 1226 7505 1228
rect 7539 1226 7578 1228
rect 7612 1226 7651 1228
rect 7685 1226 7724 1228
rect 7758 1226 7797 1228
rect 7831 1226 7870 1228
rect 7904 1226 7943 1228
rect 7977 1226 8016 1228
rect 8050 1226 8089 1228
rect 8123 1226 8162 1228
rect 8196 1226 8235 1228
rect 8269 1226 8308 1228
rect 8342 1226 8382 1228
rect 8416 1226 8456 1228
rect 8490 1226 8530 1228
rect 8564 1226 8604 1228
rect 8638 1226 8678 1228
rect 8712 1226 8752 1228
rect 8786 1226 8826 1228
rect 8860 1226 8900 1228
rect 8934 1226 8974 1228
rect 9008 1226 9048 1228
rect 9082 1226 9122 1228
rect 9156 1226 9196 1228
rect 9082 1194 9093 1226
rect 9156 1194 9162 1226
rect 9058 1192 9093 1194
rect 9127 1192 9162 1194
rect 9230 1226 9270 1228
rect 9304 1226 9344 1228
rect 9378 1226 9418 1228
rect 9452 1226 9492 1228
rect 9526 1226 9566 1228
rect 9600 1226 9640 1228
rect 9674 1226 9714 1228
rect 9230 1194 9231 1226
rect 9196 1192 9231 1194
rect 9265 1194 9270 1226
rect 9334 1194 9344 1226
rect 9403 1194 9418 1226
rect 9472 1194 9492 1226
rect 9541 1194 9566 1226
rect 9610 1194 9640 1226
rect 9265 1192 9300 1194
rect 9334 1192 9369 1194
rect 9403 1192 9438 1194
rect 9472 1192 9507 1194
rect 9541 1192 9576 1194
rect 9610 1192 9645 1194
rect 9679 1192 9714 1226
rect 9748 1192 9848 1228
rect 9058 1158 9848 1192
rect 9058 1156 9093 1158
rect 9127 1156 9162 1158
rect 9082 1124 9093 1156
rect 9156 1124 9162 1156
rect 9196 1156 9231 1158
rect 6882 1122 6921 1124
rect 6955 1122 6994 1124
rect 7028 1122 7067 1124
rect 7101 1122 7140 1124
rect 7174 1122 7213 1124
rect 7247 1122 7286 1124
rect 7320 1122 7359 1124
rect 7393 1122 7432 1124
rect 7466 1122 7505 1124
rect 7539 1122 7578 1124
rect 7612 1122 7651 1124
rect 7685 1122 7724 1124
rect 7758 1122 7797 1124
rect 7831 1122 7870 1124
rect 7904 1122 7943 1124
rect 7977 1122 8016 1124
rect 8050 1122 8089 1124
rect 8123 1122 8162 1124
rect 8196 1122 8235 1124
rect 8269 1122 8308 1124
rect 8342 1122 8382 1124
rect 8416 1122 8456 1124
rect 8490 1122 8530 1124
rect 8564 1122 8604 1124
rect 8638 1122 8678 1124
rect 8712 1122 8752 1124
rect 8786 1122 8826 1124
rect 8860 1122 8900 1124
rect 8934 1122 8974 1124
rect 9008 1122 9048 1124
rect 9082 1122 9122 1124
rect 9156 1122 9196 1124
rect 9230 1124 9231 1156
rect 9265 1156 9300 1158
rect 9334 1156 9369 1158
rect 9403 1156 9438 1158
rect 9472 1156 9507 1158
rect 9541 1156 9576 1158
rect 9610 1156 9645 1158
rect 9265 1124 9270 1156
rect 9334 1124 9344 1156
rect 9403 1124 9418 1156
rect 9472 1124 9492 1156
rect 9541 1124 9566 1156
rect 9610 1124 9640 1156
rect 9679 1124 9714 1158
rect 9230 1122 9270 1124
rect 9304 1122 9344 1124
rect 9378 1122 9418 1124
rect 9452 1122 9492 1124
rect 9526 1122 9566 1124
rect 9600 1122 9640 1124
rect 9674 1122 9714 1124
rect 9748 1122 9848 1158
rect 9990 1192 10090 1228
rect 10124 1226 10164 1228
rect 10198 1226 10238 1228
rect 10272 1226 10312 1228
rect 10346 1226 10386 1228
rect 10420 1226 10460 1228
rect 10494 1226 10534 1228
rect 10568 1226 10608 1228
rect 10124 1192 10159 1226
rect 10198 1194 10228 1226
rect 10272 1194 10297 1226
rect 10346 1194 10366 1226
rect 10420 1194 10435 1226
rect 10494 1194 10504 1226
rect 10568 1194 10573 1226
rect 10193 1192 10228 1194
rect 10262 1192 10297 1194
rect 10331 1192 10366 1194
rect 10400 1192 10435 1194
rect 10469 1192 10504 1194
rect 10538 1192 10573 1194
rect 10607 1194 10608 1226
rect 10642 1226 10682 1228
rect 10716 1226 10756 1228
rect 10790 1226 10830 1228
rect 10864 1226 10904 1228
rect 10938 1226 10978 1228
rect 11012 1226 11052 1228
rect 11086 1226 11126 1228
rect 11160 1226 11200 1228
rect 11234 1226 11274 1228
rect 11308 1226 11348 1228
rect 11382 1226 11422 1228
rect 11456 1226 11496 1228
rect 11530 1226 11569 1228
rect 11603 1226 11642 1228
rect 11676 1226 11715 1228
rect 11749 1226 11788 1228
rect 11822 1226 11861 1228
rect 11895 1226 11934 1228
rect 11968 1226 12007 1228
rect 12041 1226 12080 1228
rect 12114 1226 12153 1228
rect 12187 1226 12226 1228
rect 12260 1226 12299 1228
rect 12333 1226 12372 1228
rect 12406 1226 12445 1228
rect 12479 1226 12518 1228
rect 12552 1226 12591 1228
rect 12625 1226 12664 1228
rect 12698 1226 12737 1228
rect 12771 1226 12810 1228
rect 12844 1226 12883 1228
rect 12917 1226 12956 1228
rect 10607 1192 10642 1194
rect 10676 1194 10682 1226
rect 10745 1194 10756 1226
rect 10676 1192 10711 1194
rect 10745 1192 10780 1194
rect 9990 1158 10780 1192
rect 9990 1122 10090 1158
rect 10124 1124 10159 1158
rect 10193 1156 10228 1158
rect 10262 1156 10297 1158
rect 10331 1156 10366 1158
rect 10400 1156 10435 1158
rect 10469 1156 10504 1158
rect 10538 1156 10573 1158
rect 10198 1124 10228 1156
rect 10272 1124 10297 1156
rect 10346 1124 10366 1156
rect 10420 1124 10435 1156
rect 10494 1124 10504 1156
rect 10568 1124 10573 1156
rect 10607 1156 10642 1158
rect 10607 1124 10608 1156
rect 10124 1122 10164 1124
rect 10198 1122 10238 1124
rect 10272 1122 10312 1124
rect 10346 1122 10386 1124
rect 10420 1122 10460 1124
rect 10494 1122 10534 1124
rect 10568 1122 10608 1124
rect 10676 1156 10711 1158
rect 10745 1156 10780 1158
rect 10676 1124 10682 1156
rect 10745 1124 10756 1156
rect 10642 1122 10682 1124
rect 10716 1122 10756 1124
rect 10790 1122 10830 1124
rect 10864 1122 10904 1124
rect 10938 1122 10978 1124
rect 11012 1122 11052 1124
rect 11086 1122 11126 1124
rect 11160 1122 11200 1124
rect 11234 1122 11274 1124
rect 11308 1122 11348 1124
rect 11382 1122 11422 1124
rect 11456 1122 11496 1124
rect 11530 1122 11569 1124
rect 11603 1122 11642 1124
rect 11676 1122 11715 1124
rect 11749 1122 11788 1124
rect 11822 1122 11861 1124
rect 11895 1122 11934 1124
rect 11968 1122 12007 1124
rect 12041 1122 12080 1124
rect 12114 1122 12153 1124
rect 12187 1122 12226 1124
rect 12260 1122 12299 1124
rect 12333 1122 12372 1124
rect 12406 1122 12445 1124
rect 12479 1122 12518 1124
rect 12552 1122 12591 1124
rect 12625 1122 12664 1124
rect 12698 1122 12737 1124
rect 12771 1122 12810 1124
rect 12844 1122 12883 1124
rect 12917 1122 12956 1124
rect 12990 1122 13090 1228
rect 13232 1122 13332 1228
rect 13366 1226 13405 1228
rect 13439 1226 13478 1228
rect 13512 1226 13551 1228
rect 13585 1226 13624 1228
rect 13658 1226 13697 1228
rect 13731 1226 13770 1228
rect 13804 1226 13843 1228
rect 13877 1226 13916 1228
rect 13950 1226 13989 1228
rect 14023 1226 14062 1228
rect 14096 1226 14135 1228
rect 14169 1226 14208 1228
rect 14242 1226 14281 1228
rect 14315 1226 14354 1228
rect 14388 1226 14427 1228
rect 14461 1226 14500 1228
rect 14534 1226 14573 1228
rect 14607 1226 14646 1228
rect 14680 1226 14719 1228
rect 14753 1226 14792 1228
rect 14826 1226 14866 1228
rect 14900 1226 14940 1228
rect 14974 1226 15014 1228
rect 15048 1226 15088 1228
rect 15122 1226 15162 1228
rect 15196 1226 15236 1228
rect 15270 1226 15310 1228
rect 15344 1226 15384 1228
rect 15418 1226 15458 1228
rect 15492 1226 15532 1228
rect 15566 1226 15606 1228
rect 15640 1226 15680 1228
rect 15566 1194 15577 1226
rect 15640 1194 15646 1226
rect 15542 1192 15577 1194
rect 15611 1192 15646 1194
rect 15714 1226 15754 1228
rect 15788 1226 15828 1228
rect 15862 1226 15902 1228
rect 15936 1226 15976 1228
rect 16010 1226 16050 1228
rect 16084 1226 16124 1228
rect 16158 1226 16198 1228
rect 15714 1194 15715 1226
rect 15680 1192 15715 1194
rect 15749 1194 15754 1226
rect 15818 1194 15828 1226
rect 15887 1194 15902 1226
rect 15956 1194 15976 1226
rect 16025 1194 16050 1226
rect 16094 1194 16124 1226
rect 15749 1192 15784 1194
rect 15818 1192 15853 1194
rect 15887 1192 15922 1194
rect 15956 1192 15991 1194
rect 16025 1192 16060 1194
rect 16094 1192 16129 1194
rect 16163 1192 16198 1226
rect 16232 1192 16332 1228
rect 15542 1158 16332 1192
rect 15542 1156 15577 1158
rect 15611 1156 15646 1158
rect 15566 1124 15577 1156
rect 15640 1124 15646 1156
rect 15680 1156 15715 1158
rect 13366 1122 13405 1124
rect 13439 1122 13478 1124
rect 13512 1122 13551 1124
rect 13585 1122 13624 1124
rect 13658 1122 13697 1124
rect 13731 1122 13770 1124
rect 13804 1122 13843 1124
rect 13877 1122 13916 1124
rect 13950 1122 13989 1124
rect 14023 1122 14062 1124
rect 14096 1122 14135 1124
rect 14169 1122 14208 1124
rect 14242 1122 14281 1124
rect 14315 1122 14354 1124
rect 14388 1122 14427 1124
rect 14461 1122 14500 1124
rect 14534 1122 14573 1124
rect 14607 1122 14646 1124
rect 14680 1122 14719 1124
rect 14753 1122 14792 1124
rect 14826 1122 14866 1124
rect 14900 1122 14940 1124
rect 14974 1122 15014 1124
rect 15048 1122 15088 1124
rect 15122 1122 15162 1124
rect 15196 1122 15236 1124
rect 15270 1122 15310 1124
rect 15344 1122 15384 1124
rect 15418 1122 15458 1124
rect 15492 1122 15532 1124
rect 15566 1122 15606 1124
rect 15640 1122 15680 1124
rect 15714 1124 15715 1156
rect 15749 1156 15784 1158
rect 15818 1156 15853 1158
rect 15887 1156 15922 1158
rect 15956 1156 15991 1158
rect 16025 1156 16060 1158
rect 16094 1156 16129 1158
rect 15749 1124 15754 1156
rect 15818 1124 15828 1156
rect 15887 1124 15902 1156
rect 15956 1124 15976 1156
rect 16025 1124 16050 1156
rect 16094 1124 16124 1156
rect 16163 1124 16198 1158
rect 15714 1122 15754 1124
rect 15788 1122 15828 1124
rect 15862 1122 15902 1124
rect 15936 1122 15976 1124
rect 16010 1122 16050 1124
rect 16084 1122 16124 1124
rect 16158 1122 16198 1124
rect 16232 1122 16332 1158
rect 16474 1192 16574 1228
rect 16608 1226 16648 1228
rect 16682 1226 16722 1228
rect 16756 1226 16796 1228
rect 16830 1226 16870 1228
rect 16904 1226 16944 1228
rect 16978 1226 17018 1228
rect 17052 1226 17092 1228
rect 16608 1192 16643 1226
rect 16682 1194 16712 1226
rect 16756 1194 16781 1226
rect 16830 1194 16850 1226
rect 16904 1194 16919 1226
rect 16978 1194 16988 1226
rect 17052 1194 17057 1226
rect 16677 1192 16712 1194
rect 16746 1192 16781 1194
rect 16815 1192 16850 1194
rect 16884 1192 16919 1194
rect 16953 1192 16988 1194
rect 17022 1192 17057 1194
rect 17091 1194 17092 1226
rect 17126 1226 17166 1228
rect 17200 1226 17240 1228
rect 17274 1226 17314 1228
rect 17348 1226 17388 1228
rect 17422 1226 17462 1228
rect 17496 1226 17536 1228
rect 17570 1226 17610 1228
rect 17644 1226 17684 1228
rect 17718 1226 17758 1228
rect 17792 1226 17832 1228
rect 17866 1226 17906 1228
rect 17940 1226 17980 1228
rect 18014 1226 18053 1228
rect 18087 1226 18126 1228
rect 18160 1226 18199 1228
rect 18233 1226 18272 1228
rect 18306 1226 18345 1228
rect 18379 1226 18418 1228
rect 18452 1226 18491 1228
rect 18525 1226 18564 1228
rect 18598 1226 18637 1228
rect 18671 1226 18710 1228
rect 18744 1226 18783 1228
rect 18817 1226 18856 1228
rect 18890 1226 18929 1228
rect 18963 1226 19002 1228
rect 19036 1226 19075 1228
rect 19109 1226 19148 1228
rect 19182 1226 19221 1228
rect 19255 1226 19294 1228
rect 19328 1226 19367 1228
rect 19401 1226 19440 1228
rect 17091 1192 17126 1194
rect 17160 1194 17166 1226
rect 17229 1194 17240 1226
rect 17160 1192 17195 1194
rect 17229 1192 17264 1194
rect 16474 1158 17264 1192
rect 16474 1122 16574 1158
rect 16608 1124 16643 1158
rect 16677 1156 16712 1158
rect 16746 1156 16781 1158
rect 16815 1156 16850 1158
rect 16884 1156 16919 1158
rect 16953 1156 16988 1158
rect 17022 1156 17057 1158
rect 16682 1124 16712 1156
rect 16756 1124 16781 1156
rect 16830 1124 16850 1156
rect 16904 1124 16919 1156
rect 16978 1124 16988 1156
rect 17052 1124 17057 1156
rect 17091 1156 17126 1158
rect 17091 1124 17092 1156
rect 16608 1122 16648 1124
rect 16682 1122 16722 1124
rect 16756 1122 16796 1124
rect 16830 1122 16870 1124
rect 16904 1122 16944 1124
rect 16978 1122 17018 1124
rect 17052 1122 17092 1124
rect 17160 1156 17195 1158
rect 17229 1156 17264 1158
rect 17160 1124 17166 1156
rect 17229 1124 17240 1156
rect 17126 1122 17166 1124
rect 17200 1122 17240 1124
rect 17274 1122 17314 1124
rect 17348 1122 17388 1124
rect 17422 1122 17462 1124
rect 17496 1122 17536 1124
rect 17570 1122 17610 1124
rect 17644 1122 17684 1124
rect 17718 1122 17758 1124
rect 17792 1122 17832 1124
rect 17866 1122 17906 1124
rect 17940 1122 17980 1124
rect 18014 1122 18053 1124
rect 18087 1122 18126 1124
rect 18160 1122 18199 1124
rect 18233 1122 18272 1124
rect 18306 1122 18345 1124
rect 18379 1122 18418 1124
rect 18452 1122 18491 1124
rect 18525 1122 18564 1124
rect 18598 1122 18637 1124
rect 18671 1122 18710 1124
rect 18744 1122 18783 1124
rect 18817 1122 18856 1124
rect 18890 1122 18929 1124
rect 18963 1122 19002 1124
rect 19036 1122 19075 1124
rect 19109 1122 19148 1124
rect 19182 1122 19221 1124
rect 19255 1122 19294 1124
rect 19328 1122 19367 1124
rect 19401 1122 19440 1124
rect 19474 1122 19574 1228
rect 19838 1213 19888 1233
rect 19922 1213 19972 1247
rect 19838 1194 19972 1213
rect 19838 1160 19882 1194
rect 19916 1178 19972 1194
rect 19838 1144 19888 1160
rect 19922 1144 19972 1178
rect -52 1109 -2 1113
rect -52 1075 -46 1109
rect -12 1079 -2 1109
rect 32 1109 82 1113
rect 32 1079 42 1109
rect -12 1075 42 1079
rect 76 1075 82 1109
rect -52 1043 82 1075
rect -52 1035 -2 1043
rect -52 1001 -46 1035
rect -12 1009 -2 1035
rect 32 1035 82 1043
rect 19838 1121 19972 1144
rect 19838 1087 19882 1121
rect 19916 1109 19972 1121
rect 19838 1075 19888 1087
rect 19922 1075 19972 1109
rect 19838 1048 19972 1075
rect 32 1009 42 1035
rect -12 1001 42 1009
rect 76 1001 82 1035
rect -52 973 82 1001
rect -52 961 -2 973
rect -52 927 -46 961
rect -12 939 -2 961
rect 32 961 82 973
rect 32 939 42 961
rect -12 927 42 939
rect 76 927 82 961
rect 182 1020 216 1036
rect 182 952 216 986
rect 3423 1020 3457 1036
rect 3423 952 3457 986
rect -52 903 82 927
rect 216 918 240 938
rect 202 904 240 918
rect 3420 918 3423 938
rect 6665 1020 6699 1036
rect 6665 952 6699 986
rect 3457 918 3458 938
rect 3420 904 3458 918
rect 6662 918 6665 938
rect 9907 1020 9941 1036
rect 9907 952 9941 986
rect 6699 918 6700 938
rect 6662 904 6700 918
rect 9904 918 9907 938
rect 13150 1020 13184 1036
rect 13150 952 13184 986
rect 19622 1020 19656 1036
rect 19622 952 19656 986
rect 9941 918 9942 938
rect 9904 904 9942 918
rect 13184 918 13208 938
rect 13170 904 13208 918
rect 19838 1014 19882 1048
rect 19916 1040 19972 1048
rect 19838 1006 19888 1014
rect 19922 1006 19972 1040
rect 19838 975 19972 1006
rect 19838 941 19882 975
rect 19916 971 19972 975
rect 19656 918 19660 938
rect 19622 904 19660 918
rect 19838 937 19888 941
rect 19922 937 19972 971
rect -52 887 -2 903
rect -52 853 -46 887
rect -12 869 -2 887
rect 32 887 82 903
rect 182 902 216 904
rect 3423 902 3457 904
rect 6665 902 6699 904
rect 9907 902 9941 904
rect 13150 902 13184 904
rect 19622 902 19656 904
rect 19838 902 19972 937
rect 32 869 42 887
rect -12 853 42 869
rect 76 853 82 887
rect -52 833 82 853
rect -52 813 -2 833
rect -52 779 -46 813
rect -12 799 -2 813
rect 32 813 82 833
rect 19838 868 19882 902
rect 19922 868 19972 902
rect 19838 833 19972 868
rect 19838 829 19888 833
rect 32 799 42 813
rect -12 779 42 799
rect 76 779 82 813
rect -52 763 82 779
rect -52 739 -2 763
rect -52 705 -46 739
rect -12 729 -2 739
rect 32 739 82 763
rect 32 729 42 739
rect -12 705 42 729
rect 76 705 82 739
rect 264 710 364 816
rect 398 814 437 816
rect 471 814 510 816
rect 544 814 583 816
rect 617 814 656 816
rect 690 814 729 816
rect 763 814 802 816
rect 836 814 875 816
rect 909 814 948 816
rect 982 814 1021 816
rect 1055 814 1094 816
rect 1128 814 1167 816
rect 1201 814 1240 816
rect 1274 814 1313 816
rect 1347 814 1386 816
rect 1420 814 1459 816
rect 1493 814 1532 816
rect 1566 814 1605 816
rect 1639 814 1678 816
rect 1712 814 1751 816
rect 1785 814 1824 816
rect 1858 814 1898 816
rect 1932 814 1972 816
rect 2006 814 2046 816
rect 2080 814 2120 816
rect 2154 814 2194 816
rect 2228 814 2268 816
rect 2302 814 2342 816
rect 2376 814 2416 816
rect 2450 814 2490 816
rect 2524 814 2564 816
rect 2598 814 2638 816
rect 2672 814 2712 816
rect 2598 782 2609 814
rect 2672 782 2678 814
rect 2574 780 2609 782
rect 2643 780 2678 782
rect 2746 814 2786 816
rect 2820 814 2860 816
rect 2894 814 2934 816
rect 2968 814 3008 816
rect 3042 814 3082 816
rect 3116 814 3156 816
rect 3190 814 3230 816
rect 2746 782 2747 814
rect 2712 780 2747 782
rect 2781 782 2786 814
rect 2850 782 2860 814
rect 2919 782 2934 814
rect 2988 782 3008 814
rect 3057 782 3082 814
rect 3126 782 3156 814
rect 2781 780 2816 782
rect 2850 780 2885 782
rect 2919 780 2954 782
rect 2988 780 3023 782
rect 3057 780 3092 782
rect 3126 780 3161 782
rect 3195 780 3230 814
rect 3264 780 3364 816
rect 2574 746 3364 780
rect 2574 744 2609 746
rect 2643 744 2678 746
rect 2598 712 2609 744
rect 2672 712 2678 744
rect 2712 744 2747 746
rect 398 710 437 712
rect 471 710 510 712
rect 544 710 583 712
rect 617 710 656 712
rect 690 710 729 712
rect 763 710 802 712
rect 836 710 875 712
rect 909 710 948 712
rect 982 710 1021 712
rect 1055 710 1094 712
rect 1128 710 1167 712
rect 1201 710 1240 712
rect 1274 710 1313 712
rect 1347 710 1386 712
rect 1420 710 1459 712
rect 1493 710 1532 712
rect 1566 710 1605 712
rect 1639 710 1678 712
rect 1712 710 1751 712
rect 1785 710 1824 712
rect 1858 710 1898 712
rect 1932 710 1972 712
rect 2006 710 2046 712
rect 2080 710 2120 712
rect 2154 710 2194 712
rect 2228 710 2268 712
rect 2302 710 2342 712
rect 2376 710 2416 712
rect 2450 710 2490 712
rect 2524 710 2564 712
rect 2598 710 2638 712
rect 2672 710 2712 712
rect 2746 712 2747 744
rect 2781 744 2816 746
rect 2850 744 2885 746
rect 2919 744 2954 746
rect 2988 744 3023 746
rect 3057 744 3092 746
rect 3126 744 3161 746
rect 2781 712 2786 744
rect 2850 712 2860 744
rect 2919 712 2934 744
rect 2988 712 3008 744
rect 3057 712 3082 744
rect 3126 712 3156 744
rect 3195 712 3230 746
rect 2746 710 2786 712
rect 2820 710 2860 712
rect 2894 710 2934 712
rect 2968 710 3008 712
rect 3042 710 3082 712
rect 3116 710 3156 712
rect 3190 710 3230 712
rect 3264 710 3364 746
rect 3506 780 3606 816
rect 3640 814 3680 816
rect 3714 814 3754 816
rect 3788 814 3828 816
rect 3862 814 3902 816
rect 3936 814 3976 816
rect 4010 814 4050 816
rect 4084 814 4124 816
rect 3640 780 3675 814
rect 3714 782 3744 814
rect 3788 782 3813 814
rect 3862 782 3882 814
rect 3936 782 3951 814
rect 4010 782 4020 814
rect 4084 782 4089 814
rect 3709 780 3744 782
rect 3778 780 3813 782
rect 3847 780 3882 782
rect 3916 780 3951 782
rect 3985 780 4020 782
rect 4054 780 4089 782
rect 4123 782 4124 814
rect 4158 814 4198 816
rect 4232 814 4272 816
rect 4306 814 4346 816
rect 4380 814 4420 816
rect 4454 814 4494 816
rect 4528 814 4568 816
rect 4602 814 4642 816
rect 4676 814 4716 816
rect 4750 814 4790 816
rect 4824 814 4864 816
rect 4898 814 4938 816
rect 4972 814 5012 816
rect 5046 814 5085 816
rect 5119 814 5158 816
rect 5192 814 5231 816
rect 5265 814 5304 816
rect 5338 814 5377 816
rect 5411 814 5450 816
rect 5484 814 5523 816
rect 5557 814 5596 816
rect 5630 814 5669 816
rect 5703 814 5742 816
rect 5776 814 5815 816
rect 5849 814 5888 816
rect 5922 814 5961 816
rect 5995 814 6034 816
rect 6068 814 6107 816
rect 6141 814 6180 816
rect 6214 814 6253 816
rect 6287 814 6326 816
rect 6360 814 6399 816
rect 6433 814 6472 816
rect 4123 780 4158 782
rect 4192 782 4198 814
rect 4261 782 4272 814
rect 4192 780 4227 782
rect 4261 780 4296 782
rect 3506 746 4296 780
rect 3506 710 3606 746
rect 3640 712 3675 746
rect 3709 744 3744 746
rect 3778 744 3813 746
rect 3847 744 3882 746
rect 3916 744 3951 746
rect 3985 744 4020 746
rect 4054 744 4089 746
rect 3714 712 3744 744
rect 3788 712 3813 744
rect 3862 712 3882 744
rect 3936 712 3951 744
rect 4010 712 4020 744
rect 4084 712 4089 744
rect 4123 744 4158 746
rect 4123 712 4124 744
rect 3640 710 3680 712
rect 3714 710 3754 712
rect 3788 710 3828 712
rect 3862 710 3902 712
rect 3936 710 3976 712
rect 4010 710 4050 712
rect 4084 710 4124 712
rect 4192 744 4227 746
rect 4261 744 4296 746
rect 4192 712 4198 744
rect 4261 712 4272 744
rect 4158 710 4198 712
rect 4232 710 4272 712
rect 4306 710 4346 712
rect 4380 710 4420 712
rect 4454 710 4494 712
rect 4528 710 4568 712
rect 4602 710 4642 712
rect 4676 710 4716 712
rect 4750 710 4790 712
rect 4824 710 4864 712
rect 4898 710 4938 712
rect 4972 710 5012 712
rect 5046 710 5085 712
rect 5119 710 5158 712
rect 5192 710 5231 712
rect 5265 710 5304 712
rect 5338 710 5377 712
rect 5411 710 5450 712
rect 5484 710 5523 712
rect 5557 710 5596 712
rect 5630 710 5669 712
rect 5703 710 5742 712
rect 5776 710 5815 712
rect 5849 710 5888 712
rect 5922 710 5961 712
rect 5995 710 6034 712
rect 6068 710 6107 712
rect 6141 710 6180 712
rect 6214 710 6253 712
rect 6287 710 6326 712
rect 6360 710 6399 712
rect 6433 710 6472 712
rect 6506 710 6606 816
rect 6748 710 6848 816
rect 6882 814 6921 816
rect 6955 814 6994 816
rect 7028 814 7067 816
rect 7101 814 7140 816
rect 7174 814 7213 816
rect 7247 814 7286 816
rect 7320 814 7359 816
rect 7393 814 7432 816
rect 7466 814 7505 816
rect 7539 814 7578 816
rect 7612 814 7651 816
rect 7685 814 7724 816
rect 7758 814 7797 816
rect 7831 814 7870 816
rect 7904 814 7943 816
rect 7977 814 8016 816
rect 8050 814 8089 816
rect 8123 814 8162 816
rect 8196 814 8235 816
rect 8269 814 8308 816
rect 8342 814 8382 816
rect 8416 814 8456 816
rect 8490 814 8530 816
rect 8564 814 8604 816
rect 8638 814 8678 816
rect 8712 814 8752 816
rect 8786 814 8826 816
rect 8860 814 8900 816
rect 8934 814 8974 816
rect 9008 814 9048 816
rect 9082 814 9122 816
rect 9156 814 9196 816
rect 9082 782 9093 814
rect 9156 782 9162 814
rect 9058 780 9093 782
rect 9127 780 9162 782
rect 9230 814 9270 816
rect 9304 814 9344 816
rect 9378 814 9418 816
rect 9452 814 9492 816
rect 9526 814 9566 816
rect 9600 814 9640 816
rect 9674 814 9714 816
rect 9230 782 9231 814
rect 9196 780 9231 782
rect 9265 782 9270 814
rect 9334 782 9344 814
rect 9403 782 9418 814
rect 9472 782 9492 814
rect 9541 782 9566 814
rect 9610 782 9640 814
rect 9265 780 9300 782
rect 9334 780 9369 782
rect 9403 780 9438 782
rect 9472 780 9507 782
rect 9541 780 9576 782
rect 9610 780 9645 782
rect 9679 780 9714 814
rect 9748 780 9848 816
rect 9058 746 9848 780
rect 9058 744 9093 746
rect 9127 744 9162 746
rect 9082 712 9093 744
rect 9156 712 9162 744
rect 9196 744 9231 746
rect 6882 710 6921 712
rect 6955 710 6994 712
rect 7028 710 7067 712
rect 7101 710 7140 712
rect 7174 710 7213 712
rect 7247 710 7286 712
rect 7320 710 7359 712
rect 7393 710 7432 712
rect 7466 710 7505 712
rect 7539 710 7578 712
rect 7612 710 7651 712
rect 7685 710 7724 712
rect 7758 710 7797 712
rect 7831 710 7870 712
rect 7904 710 7943 712
rect 7977 710 8016 712
rect 8050 710 8089 712
rect 8123 710 8162 712
rect 8196 710 8235 712
rect 8269 710 8308 712
rect 8342 710 8382 712
rect 8416 710 8456 712
rect 8490 710 8530 712
rect 8564 710 8604 712
rect 8638 710 8678 712
rect 8712 710 8752 712
rect 8786 710 8826 712
rect 8860 710 8900 712
rect 8934 710 8974 712
rect 9008 710 9048 712
rect 9082 710 9122 712
rect 9156 710 9196 712
rect 9230 712 9231 744
rect 9265 744 9300 746
rect 9334 744 9369 746
rect 9403 744 9438 746
rect 9472 744 9507 746
rect 9541 744 9576 746
rect 9610 744 9645 746
rect 9265 712 9270 744
rect 9334 712 9344 744
rect 9403 712 9418 744
rect 9472 712 9492 744
rect 9541 712 9566 744
rect 9610 712 9640 744
rect 9679 712 9714 746
rect 9230 710 9270 712
rect 9304 710 9344 712
rect 9378 710 9418 712
rect 9452 710 9492 712
rect 9526 710 9566 712
rect 9600 710 9640 712
rect 9674 710 9714 712
rect 9748 710 9848 746
rect 9990 780 10090 816
rect 10124 814 10164 816
rect 10198 814 10238 816
rect 10272 814 10312 816
rect 10346 814 10386 816
rect 10420 814 10460 816
rect 10494 814 10534 816
rect 10568 814 10608 816
rect 10124 780 10159 814
rect 10198 782 10228 814
rect 10272 782 10297 814
rect 10346 782 10366 814
rect 10420 782 10435 814
rect 10494 782 10504 814
rect 10568 782 10573 814
rect 10193 780 10228 782
rect 10262 780 10297 782
rect 10331 780 10366 782
rect 10400 780 10435 782
rect 10469 780 10504 782
rect 10538 780 10573 782
rect 10607 782 10608 814
rect 10642 814 10682 816
rect 10716 814 10756 816
rect 10790 814 10830 816
rect 10864 814 10904 816
rect 10938 814 10978 816
rect 11012 814 11052 816
rect 11086 814 11126 816
rect 11160 814 11200 816
rect 11234 814 11274 816
rect 11308 814 11348 816
rect 11382 814 11422 816
rect 11456 814 11496 816
rect 11530 814 11569 816
rect 11603 814 11642 816
rect 11676 814 11715 816
rect 11749 814 11788 816
rect 11822 814 11861 816
rect 11895 814 11934 816
rect 11968 814 12007 816
rect 12041 814 12080 816
rect 12114 814 12153 816
rect 12187 814 12226 816
rect 12260 814 12299 816
rect 12333 814 12372 816
rect 12406 814 12445 816
rect 12479 814 12518 816
rect 12552 814 12591 816
rect 12625 814 12664 816
rect 12698 814 12737 816
rect 12771 814 12810 816
rect 12844 814 12883 816
rect 12917 814 12956 816
rect 10607 780 10642 782
rect 10676 782 10682 814
rect 10745 782 10756 814
rect 10676 780 10711 782
rect 10745 780 10780 782
rect 9990 746 10780 780
rect 9990 710 10090 746
rect 10124 712 10159 746
rect 10193 744 10228 746
rect 10262 744 10297 746
rect 10331 744 10366 746
rect 10400 744 10435 746
rect 10469 744 10504 746
rect 10538 744 10573 746
rect 10198 712 10228 744
rect 10272 712 10297 744
rect 10346 712 10366 744
rect 10420 712 10435 744
rect 10494 712 10504 744
rect 10568 712 10573 744
rect 10607 744 10642 746
rect 10607 712 10608 744
rect 10124 710 10164 712
rect 10198 710 10238 712
rect 10272 710 10312 712
rect 10346 710 10386 712
rect 10420 710 10460 712
rect 10494 710 10534 712
rect 10568 710 10608 712
rect 10676 744 10711 746
rect 10745 744 10780 746
rect 10676 712 10682 744
rect 10745 712 10756 744
rect 10642 710 10682 712
rect 10716 710 10756 712
rect 10790 710 10830 712
rect 10864 710 10904 712
rect 10938 710 10978 712
rect 11012 710 11052 712
rect 11086 710 11126 712
rect 11160 710 11200 712
rect 11234 710 11274 712
rect 11308 710 11348 712
rect 11382 710 11422 712
rect 11456 710 11496 712
rect 11530 710 11569 712
rect 11603 710 11642 712
rect 11676 710 11715 712
rect 11749 710 11788 712
rect 11822 710 11861 712
rect 11895 710 11934 712
rect 11968 710 12007 712
rect 12041 710 12080 712
rect 12114 710 12153 712
rect 12187 710 12226 712
rect 12260 710 12299 712
rect 12333 710 12372 712
rect 12406 710 12445 712
rect 12479 710 12518 712
rect 12552 710 12591 712
rect 12625 710 12664 712
rect 12698 710 12737 712
rect 12771 710 12810 712
rect 12844 710 12883 712
rect 12917 710 12956 712
rect 12990 710 13090 816
rect 13232 710 13332 816
rect 13366 814 13405 816
rect 13439 814 13478 816
rect 13512 814 13551 816
rect 13585 814 13624 816
rect 13658 814 13697 816
rect 13731 814 13770 816
rect 13804 814 13843 816
rect 13877 814 13916 816
rect 13950 814 13989 816
rect 14023 814 14062 816
rect 14096 814 14135 816
rect 14169 814 14208 816
rect 14242 814 14281 816
rect 14315 814 14354 816
rect 14388 814 14427 816
rect 14461 814 14500 816
rect 14534 814 14573 816
rect 14607 814 14646 816
rect 14680 814 14719 816
rect 14753 814 14792 816
rect 14826 814 14866 816
rect 14900 814 14940 816
rect 14974 814 15014 816
rect 15048 814 15088 816
rect 15122 814 15162 816
rect 15196 814 15236 816
rect 15270 814 15310 816
rect 15344 814 15384 816
rect 15418 814 15458 816
rect 15492 814 15532 816
rect 15566 814 15606 816
rect 15640 814 15680 816
rect 15566 782 15577 814
rect 15640 782 15646 814
rect 15542 780 15577 782
rect 15611 780 15646 782
rect 15714 814 15754 816
rect 15788 814 15828 816
rect 15862 814 15902 816
rect 15936 814 15976 816
rect 16010 814 16050 816
rect 16084 814 16124 816
rect 16158 814 16198 816
rect 15714 782 15715 814
rect 15680 780 15715 782
rect 15749 782 15754 814
rect 15818 782 15828 814
rect 15887 782 15902 814
rect 15956 782 15976 814
rect 16025 782 16050 814
rect 16094 782 16124 814
rect 15749 780 15784 782
rect 15818 780 15853 782
rect 15887 780 15922 782
rect 15956 780 15991 782
rect 16025 780 16060 782
rect 16094 780 16129 782
rect 16163 780 16198 814
rect 16232 780 16332 816
rect 15542 746 16332 780
rect 15542 744 15577 746
rect 15611 744 15646 746
rect 15566 712 15577 744
rect 15640 712 15646 744
rect 15680 744 15715 746
rect 13366 710 13405 712
rect 13439 710 13478 712
rect 13512 710 13551 712
rect 13585 710 13624 712
rect 13658 710 13697 712
rect 13731 710 13770 712
rect 13804 710 13843 712
rect 13877 710 13916 712
rect 13950 710 13989 712
rect 14023 710 14062 712
rect 14096 710 14135 712
rect 14169 710 14208 712
rect 14242 710 14281 712
rect 14315 710 14354 712
rect 14388 710 14427 712
rect 14461 710 14500 712
rect 14534 710 14573 712
rect 14607 710 14646 712
rect 14680 710 14719 712
rect 14753 710 14792 712
rect 14826 710 14866 712
rect 14900 710 14940 712
rect 14974 710 15014 712
rect 15048 710 15088 712
rect 15122 710 15162 712
rect 15196 710 15236 712
rect 15270 710 15310 712
rect 15344 710 15384 712
rect 15418 710 15458 712
rect 15492 710 15532 712
rect 15566 710 15606 712
rect 15640 710 15680 712
rect 15714 712 15715 744
rect 15749 744 15784 746
rect 15818 744 15853 746
rect 15887 744 15922 746
rect 15956 744 15991 746
rect 16025 744 16060 746
rect 16094 744 16129 746
rect 15749 712 15754 744
rect 15818 712 15828 744
rect 15887 712 15902 744
rect 15956 712 15976 744
rect 16025 712 16050 744
rect 16094 712 16124 744
rect 16163 712 16198 746
rect 15714 710 15754 712
rect 15788 710 15828 712
rect 15862 710 15902 712
rect 15936 710 15976 712
rect 16010 710 16050 712
rect 16084 710 16124 712
rect 16158 710 16198 712
rect 16232 710 16332 746
rect 16474 780 16574 816
rect 16608 814 16648 816
rect 16682 814 16722 816
rect 16756 814 16796 816
rect 16830 814 16870 816
rect 16904 814 16944 816
rect 16978 814 17018 816
rect 17052 814 17092 816
rect 16608 780 16643 814
rect 16682 782 16712 814
rect 16756 782 16781 814
rect 16830 782 16850 814
rect 16904 782 16919 814
rect 16978 782 16988 814
rect 17052 782 17057 814
rect 16677 780 16712 782
rect 16746 780 16781 782
rect 16815 780 16850 782
rect 16884 780 16919 782
rect 16953 780 16988 782
rect 17022 780 17057 782
rect 17091 782 17092 814
rect 17126 814 17166 816
rect 17200 814 17240 816
rect 17274 814 17314 816
rect 17348 814 17388 816
rect 17422 814 17462 816
rect 17496 814 17536 816
rect 17570 814 17610 816
rect 17644 814 17684 816
rect 17718 814 17758 816
rect 17792 814 17832 816
rect 17866 814 17906 816
rect 17940 814 17980 816
rect 18014 814 18053 816
rect 18087 814 18126 816
rect 18160 814 18199 816
rect 18233 814 18272 816
rect 18306 814 18345 816
rect 18379 814 18418 816
rect 18452 814 18491 816
rect 18525 814 18564 816
rect 18598 814 18637 816
rect 18671 814 18710 816
rect 18744 814 18783 816
rect 18817 814 18856 816
rect 18890 814 18929 816
rect 18963 814 19002 816
rect 19036 814 19075 816
rect 19109 814 19148 816
rect 19182 814 19221 816
rect 19255 814 19294 816
rect 19328 814 19367 816
rect 19401 814 19440 816
rect 17091 780 17126 782
rect 17160 782 17166 814
rect 17229 782 17240 814
rect 17160 780 17195 782
rect 17229 780 17264 782
rect 16474 746 17264 780
rect 16474 710 16574 746
rect 16608 712 16643 746
rect 16677 744 16712 746
rect 16746 744 16781 746
rect 16815 744 16850 746
rect 16884 744 16919 746
rect 16953 744 16988 746
rect 17022 744 17057 746
rect 16682 712 16712 744
rect 16756 712 16781 744
rect 16830 712 16850 744
rect 16904 712 16919 744
rect 16978 712 16988 744
rect 17052 712 17057 744
rect 17091 744 17126 746
rect 17091 712 17092 744
rect 16608 710 16648 712
rect 16682 710 16722 712
rect 16756 710 16796 712
rect 16830 710 16870 712
rect 16904 710 16944 712
rect 16978 710 17018 712
rect 17052 710 17092 712
rect 17160 744 17195 746
rect 17229 744 17264 746
rect 17160 712 17166 744
rect 17229 712 17240 744
rect 17126 710 17166 712
rect 17200 710 17240 712
rect 17274 710 17314 712
rect 17348 710 17388 712
rect 17422 710 17462 712
rect 17496 710 17536 712
rect 17570 710 17610 712
rect 17644 710 17684 712
rect 17718 710 17758 712
rect 17792 710 17832 712
rect 17866 710 17906 712
rect 17940 710 17980 712
rect 18014 710 18053 712
rect 18087 710 18126 712
rect 18160 710 18199 712
rect 18233 710 18272 712
rect 18306 710 18345 712
rect 18379 710 18418 712
rect 18452 710 18491 712
rect 18525 710 18564 712
rect 18598 710 18637 712
rect 18671 710 18710 712
rect 18744 710 18783 712
rect 18817 710 18856 712
rect 18890 710 18929 712
rect 18963 710 19002 712
rect 19036 710 19075 712
rect 19109 710 19148 712
rect 19182 710 19221 712
rect 19255 710 19294 712
rect 19328 710 19367 712
rect 19401 710 19440 712
rect 19474 710 19574 816
rect 19838 795 19882 829
rect 19922 799 19972 833
rect 19916 795 19972 799
rect 19838 763 19972 795
rect 19838 756 19888 763
rect 19838 722 19882 756
rect 19922 729 19972 763
rect 19916 722 19972 729
rect -52 693 82 705
rect -52 665 -2 693
rect -52 631 -46 665
rect -12 659 -2 665
rect 32 665 82 693
rect 32 659 42 665
rect -12 631 42 659
rect 76 631 82 665
rect -52 623 82 631
rect 19838 693 19972 722
rect 19838 683 19888 693
rect 19838 649 19882 683
rect 19922 659 19972 693
rect 19916 649 19972 659
rect -52 591 -2 623
rect -52 557 -46 591
rect -12 589 -2 591
rect 32 591 82 623
rect 182 622 216 624
rect 3423 622 3457 624
rect 6665 622 6699 624
rect 9907 622 9941 624
rect 13149 622 13183 624
rect 16391 622 16425 624
rect 19622 622 19656 624
rect 19838 623 19972 649
rect 32 589 42 591
rect -12 557 42 589
rect 76 557 82 591
rect 178 608 216 622
rect 178 588 182 608
rect -52 553 82 557
rect -52 519 -2 553
rect 32 519 82 553
rect -52 517 82 519
rect -52 483 -46 517
rect -12 483 42 517
rect 76 483 82 517
rect 3420 608 3458 622
rect 3420 588 3423 608
rect 182 540 216 574
rect 182 490 216 506
rect 3457 588 3458 608
rect 6662 608 6700 622
rect 6662 588 6665 608
rect 3423 540 3457 574
rect 3423 490 3457 506
rect 6699 588 6700 608
rect 9904 608 9942 622
rect 9904 588 9907 608
rect 6665 540 6699 574
rect 6665 490 6699 506
rect 9941 588 9942 608
rect 13146 608 13184 622
rect 13146 588 13149 608
rect 9907 540 9941 574
rect 9907 490 9941 506
rect 13183 588 13184 608
rect 16388 608 16426 622
rect 16388 588 16391 608
rect 13149 540 13183 574
rect 13149 490 13183 506
rect 16425 588 16426 608
rect 19598 608 19636 622
rect 19598 588 19622 608
rect 19838 610 19888 623
rect 16391 540 16425 574
rect 16391 490 16425 506
rect 19622 540 19656 574
rect 19622 490 19656 506
rect 19838 576 19882 610
rect 19922 589 19972 623
rect 19916 576 19972 589
rect 19838 553 19972 576
rect 19838 537 19888 553
rect 19838 503 19882 537
rect 19922 519 19972 553
rect 19916 503 19972 519
rect -52 449 -2 483
rect 32 449 82 483
rect -52 443 82 449
rect -52 409 -46 443
rect -12 413 42 443
rect -12 409 -2 413
rect -52 379 -2 409
rect 32 409 42 413
rect 76 409 82 443
rect 32 379 82 409
rect 19838 483 19972 503
rect 19838 465 19888 483
rect 19838 431 19882 465
rect 19922 449 19972 483
rect 19916 431 19972 449
rect 19838 413 19972 431
rect -52 369 82 379
rect -52 335 -46 369
rect -12 343 42 369
rect -12 335 -2 343
rect -52 309 -2 335
rect 32 335 42 343
rect 76 335 82 369
rect 32 309 82 335
rect -52 295 82 309
rect 264 298 364 404
rect 398 402 437 404
rect 471 402 510 404
rect 544 402 583 404
rect 617 402 656 404
rect 690 402 729 404
rect 763 402 802 404
rect 836 402 875 404
rect 909 402 948 404
rect 982 402 1021 404
rect 1055 402 1094 404
rect 1128 402 1167 404
rect 1201 402 1240 404
rect 1274 402 1313 404
rect 1347 402 1386 404
rect 1420 402 1459 404
rect 1493 402 1532 404
rect 1566 402 1605 404
rect 1639 402 1678 404
rect 1712 402 1751 404
rect 1785 402 1824 404
rect 1858 402 1898 404
rect 1932 402 1972 404
rect 2006 402 2046 404
rect 2080 402 2120 404
rect 2154 402 2194 404
rect 2228 402 2268 404
rect 2302 402 2342 404
rect 2376 402 2416 404
rect 2450 402 2490 404
rect 2524 402 2564 404
rect 2598 402 2638 404
rect 2672 402 2712 404
rect 2598 370 2609 402
rect 2672 370 2678 402
rect 2574 368 2609 370
rect 2643 368 2678 370
rect 2746 402 2786 404
rect 2820 402 2860 404
rect 2894 402 2934 404
rect 2968 402 3008 404
rect 3042 402 3082 404
rect 3116 402 3156 404
rect 3190 402 3230 404
rect 2746 370 2747 402
rect 2712 368 2747 370
rect 2781 370 2786 402
rect 2850 370 2860 402
rect 2919 370 2934 402
rect 2988 370 3008 402
rect 3057 370 3082 402
rect 3126 370 3156 402
rect 2781 368 2816 370
rect 2850 368 2885 370
rect 2919 368 2954 370
rect 2988 368 3023 370
rect 3057 368 3092 370
rect 3126 368 3161 370
rect 3195 368 3230 402
rect 3264 368 3364 404
rect 2574 334 3364 368
rect 2574 332 2609 334
rect 2643 332 2678 334
rect 2598 300 2609 332
rect 2672 300 2678 332
rect 2712 332 2747 334
rect 398 298 437 300
rect 471 298 510 300
rect 544 298 583 300
rect 617 298 656 300
rect 690 298 729 300
rect 763 298 802 300
rect 836 298 875 300
rect 909 298 948 300
rect 982 298 1021 300
rect 1055 298 1094 300
rect 1128 298 1167 300
rect 1201 298 1240 300
rect 1274 298 1313 300
rect 1347 298 1386 300
rect 1420 298 1459 300
rect 1493 298 1532 300
rect 1566 298 1605 300
rect 1639 298 1678 300
rect 1712 298 1751 300
rect 1785 298 1824 300
rect 1858 298 1898 300
rect 1932 298 1972 300
rect 2006 298 2046 300
rect 2080 298 2120 300
rect 2154 298 2194 300
rect 2228 298 2268 300
rect 2302 298 2342 300
rect 2376 298 2416 300
rect 2450 298 2490 300
rect 2524 298 2564 300
rect 2598 298 2638 300
rect 2672 298 2712 300
rect 2746 300 2747 332
rect 2781 332 2816 334
rect 2850 332 2885 334
rect 2919 332 2954 334
rect 2988 332 3023 334
rect 3057 332 3092 334
rect 3126 332 3161 334
rect 2781 300 2786 332
rect 2850 300 2860 332
rect 2919 300 2934 332
rect 2988 300 3008 332
rect 3057 300 3082 332
rect 3126 300 3156 332
rect 3195 300 3230 334
rect 2746 298 2786 300
rect 2820 298 2860 300
rect 2894 298 2934 300
rect 2968 298 3008 300
rect 3042 298 3082 300
rect 3116 298 3156 300
rect 3190 298 3230 300
rect 3264 298 3364 334
rect 3506 368 3606 404
rect 3640 402 3680 404
rect 3714 402 3754 404
rect 3788 402 3828 404
rect 3862 402 3902 404
rect 3936 402 3976 404
rect 4010 402 4050 404
rect 4084 402 4124 404
rect 3640 368 3675 402
rect 3714 370 3744 402
rect 3788 370 3813 402
rect 3862 370 3882 402
rect 3936 370 3951 402
rect 4010 370 4020 402
rect 4084 370 4089 402
rect 3709 368 3744 370
rect 3778 368 3813 370
rect 3847 368 3882 370
rect 3916 368 3951 370
rect 3985 368 4020 370
rect 4054 368 4089 370
rect 4123 370 4124 402
rect 4158 402 4198 404
rect 4232 402 4272 404
rect 4306 402 4346 404
rect 4380 402 4420 404
rect 4454 402 4494 404
rect 4528 402 4568 404
rect 4602 402 4642 404
rect 4676 402 4716 404
rect 4750 402 4790 404
rect 4824 402 4864 404
rect 4898 402 4938 404
rect 4972 402 5012 404
rect 5046 402 5085 404
rect 5119 402 5158 404
rect 5192 402 5231 404
rect 5265 402 5304 404
rect 5338 402 5377 404
rect 5411 402 5450 404
rect 5484 402 5523 404
rect 5557 402 5596 404
rect 5630 402 5669 404
rect 5703 402 5742 404
rect 5776 402 5815 404
rect 5849 402 5888 404
rect 5922 402 5961 404
rect 5995 402 6034 404
rect 6068 402 6107 404
rect 6141 402 6180 404
rect 6214 402 6253 404
rect 6287 402 6326 404
rect 6360 402 6399 404
rect 6433 402 6472 404
rect 4123 368 4158 370
rect 4192 370 4198 402
rect 4261 370 4272 402
rect 4192 368 4227 370
rect 4261 368 4296 370
rect 3506 334 4296 368
rect 3506 298 3606 334
rect 3640 300 3675 334
rect 3709 332 3744 334
rect 3778 332 3813 334
rect 3847 332 3882 334
rect 3916 332 3951 334
rect 3985 332 4020 334
rect 4054 332 4089 334
rect 3714 300 3744 332
rect 3788 300 3813 332
rect 3862 300 3882 332
rect 3936 300 3951 332
rect 4010 300 4020 332
rect 4084 300 4089 332
rect 4123 332 4158 334
rect 4123 300 4124 332
rect 3640 298 3680 300
rect 3714 298 3754 300
rect 3788 298 3828 300
rect 3862 298 3902 300
rect 3936 298 3976 300
rect 4010 298 4050 300
rect 4084 298 4124 300
rect 4192 332 4227 334
rect 4261 332 4296 334
rect 4192 300 4198 332
rect 4261 300 4272 332
rect 4158 298 4198 300
rect 4232 298 4272 300
rect 4306 298 4346 300
rect 4380 298 4420 300
rect 4454 298 4494 300
rect 4528 298 4568 300
rect 4602 298 4642 300
rect 4676 298 4716 300
rect 4750 298 4790 300
rect 4824 298 4864 300
rect 4898 298 4938 300
rect 4972 298 5012 300
rect 5046 298 5085 300
rect 5119 298 5158 300
rect 5192 298 5231 300
rect 5265 298 5304 300
rect 5338 298 5377 300
rect 5411 298 5450 300
rect 5484 298 5523 300
rect 5557 298 5596 300
rect 5630 298 5669 300
rect 5703 298 5742 300
rect 5776 298 5815 300
rect 5849 298 5888 300
rect 5922 298 5961 300
rect 5995 298 6034 300
rect 6068 298 6107 300
rect 6141 298 6180 300
rect 6214 298 6253 300
rect 6287 298 6326 300
rect 6360 298 6399 300
rect 6433 298 6472 300
rect 6506 298 6606 404
rect 6748 298 6848 404
rect 6882 402 6921 404
rect 6955 402 6994 404
rect 7028 402 7067 404
rect 7101 402 7140 404
rect 7174 402 7213 404
rect 7247 402 7286 404
rect 7320 402 7359 404
rect 7393 402 7432 404
rect 7466 402 7505 404
rect 7539 402 7578 404
rect 7612 402 7651 404
rect 7685 402 7724 404
rect 7758 402 7797 404
rect 7831 402 7870 404
rect 7904 402 7943 404
rect 7977 402 8016 404
rect 8050 402 8089 404
rect 8123 402 8162 404
rect 8196 402 8235 404
rect 8269 402 8308 404
rect 8342 402 8382 404
rect 8416 402 8456 404
rect 8490 402 8530 404
rect 8564 402 8604 404
rect 8638 402 8678 404
rect 8712 402 8752 404
rect 8786 402 8826 404
rect 8860 402 8900 404
rect 8934 402 8974 404
rect 9008 402 9048 404
rect 9082 402 9122 404
rect 9156 402 9196 404
rect 9082 370 9093 402
rect 9156 370 9162 402
rect 9058 368 9093 370
rect 9127 368 9162 370
rect 9230 402 9270 404
rect 9304 402 9344 404
rect 9378 402 9418 404
rect 9452 402 9492 404
rect 9526 402 9566 404
rect 9600 402 9640 404
rect 9674 402 9714 404
rect 9230 370 9231 402
rect 9196 368 9231 370
rect 9265 370 9270 402
rect 9334 370 9344 402
rect 9403 370 9418 402
rect 9472 370 9492 402
rect 9541 370 9566 402
rect 9610 370 9640 402
rect 9265 368 9300 370
rect 9334 368 9369 370
rect 9403 368 9438 370
rect 9472 368 9507 370
rect 9541 368 9576 370
rect 9610 368 9645 370
rect 9679 368 9714 402
rect 9748 368 9848 404
rect 9058 334 9848 368
rect 9058 332 9093 334
rect 9127 332 9162 334
rect 9082 300 9093 332
rect 9156 300 9162 332
rect 9196 332 9231 334
rect 6882 298 6921 300
rect 6955 298 6994 300
rect 7028 298 7067 300
rect 7101 298 7140 300
rect 7174 298 7213 300
rect 7247 298 7286 300
rect 7320 298 7359 300
rect 7393 298 7432 300
rect 7466 298 7505 300
rect 7539 298 7578 300
rect 7612 298 7651 300
rect 7685 298 7724 300
rect 7758 298 7797 300
rect 7831 298 7870 300
rect 7904 298 7943 300
rect 7977 298 8016 300
rect 8050 298 8089 300
rect 8123 298 8162 300
rect 8196 298 8235 300
rect 8269 298 8308 300
rect 8342 298 8382 300
rect 8416 298 8456 300
rect 8490 298 8530 300
rect 8564 298 8604 300
rect 8638 298 8678 300
rect 8712 298 8752 300
rect 8786 298 8826 300
rect 8860 298 8900 300
rect 8934 298 8974 300
rect 9008 298 9048 300
rect 9082 298 9122 300
rect 9156 298 9196 300
rect 9230 300 9231 332
rect 9265 332 9300 334
rect 9334 332 9369 334
rect 9403 332 9438 334
rect 9472 332 9507 334
rect 9541 332 9576 334
rect 9610 332 9645 334
rect 9265 300 9270 332
rect 9334 300 9344 332
rect 9403 300 9418 332
rect 9472 300 9492 332
rect 9541 300 9566 332
rect 9610 300 9640 332
rect 9679 300 9714 334
rect 9230 298 9270 300
rect 9304 298 9344 300
rect 9378 298 9418 300
rect 9452 298 9492 300
rect 9526 298 9566 300
rect 9600 298 9640 300
rect 9674 298 9714 300
rect 9748 298 9848 334
rect 9990 368 10090 404
rect 10124 402 10164 404
rect 10198 402 10238 404
rect 10272 402 10312 404
rect 10346 402 10386 404
rect 10420 402 10460 404
rect 10494 402 10534 404
rect 10568 402 10608 404
rect 10124 368 10159 402
rect 10198 370 10228 402
rect 10272 370 10297 402
rect 10346 370 10366 402
rect 10420 370 10435 402
rect 10494 370 10504 402
rect 10568 370 10573 402
rect 10193 368 10228 370
rect 10262 368 10297 370
rect 10331 368 10366 370
rect 10400 368 10435 370
rect 10469 368 10504 370
rect 10538 368 10573 370
rect 10607 370 10608 402
rect 10642 402 10682 404
rect 10716 402 10756 404
rect 10790 402 10830 404
rect 10864 402 10904 404
rect 10938 402 10978 404
rect 11012 402 11052 404
rect 11086 402 11126 404
rect 11160 402 11200 404
rect 11234 402 11274 404
rect 11308 402 11348 404
rect 11382 402 11422 404
rect 11456 402 11496 404
rect 11530 402 11569 404
rect 11603 402 11642 404
rect 11676 402 11715 404
rect 11749 402 11788 404
rect 11822 402 11861 404
rect 11895 402 11934 404
rect 11968 402 12007 404
rect 12041 402 12080 404
rect 12114 402 12153 404
rect 12187 402 12226 404
rect 12260 402 12299 404
rect 12333 402 12372 404
rect 12406 402 12445 404
rect 12479 402 12518 404
rect 12552 402 12591 404
rect 12625 402 12664 404
rect 12698 402 12737 404
rect 12771 402 12810 404
rect 12844 402 12883 404
rect 12917 402 12956 404
rect 10607 368 10642 370
rect 10676 370 10682 402
rect 10745 370 10756 402
rect 10676 368 10711 370
rect 10745 368 10780 370
rect 9990 334 10780 368
rect 9990 298 10090 334
rect 10124 300 10159 334
rect 10193 332 10228 334
rect 10262 332 10297 334
rect 10331 332 10366 334
rect 10400 332 10435 334
rect 10469 332 10504 334
rect 10538 332 10573 334
rect 10198 300 10228 332
rect 10272 300 10297 332
rect 10346 300 10366 332
rect 10420 300 10435 332
rect 10494 300 10504 332
rect 10568 300 10573 332
rect 10607 332 10642 334
rect 10607 300 10608 332
rect 10124 298 10164 300
rect 10198 298 10238 300
rect 10272 298 10312 300
rect 10346 298 10386 300
rect 10420 298 10460 300
rect 10494 298 10534 300
rect 10568 298 10608 300
rect 10676 332 10711 334
rect 10745 332 10780 334
rect 10676 300 10682 332
rect 10745 300 10756 332
rect 10642 298 10682 300
rect 10716 298 10756 300
rect 10790 298 10830 300
rect 10864 298 10904 300
rect 10938 298 10978 300
rect 11012 298 11052 300
rect 11086 298 11126 300
rect 11160 298 11200 300
rect 11234 298 11274 300
rect 11308 298 11348 300
rect 11382 298 11422 300
rect 11456 298 11496 300
rect 11530 298 11569 300
rect 11603 298 11642 300
rect 11676 298 11715 300
rect 11749 298 11788 300
rect 11822 298 11861 300
rect 11895 298 11934 300
rect 11968 298 12007 300
rect 12041 298 12080 300
rect 12114 298 12153 300
rect 12187 298 12226 300
rect 12260 298 12299 300
rect 12333 298 12372 300
rect 12406 298 12445 300
rect 12479 298 12518 300
rect 12552 298 12591 300
rect 12625 298 12664 300
rect 12698 298 12737 300
rect 12771 298 12810 300
rect 12844 298 12883 300
rect 12917 298 12956 300
rect 12990 298 13090 404
rect 13232 298 13332 404
rect 13366 402 13405 404
rect 13439 402 13478 404
rect 13512 402 13551 404
rect 13585 402 13624 404
rect 13658 402 13697 404
rect 13731 402 13770 404
rect 13804 402 13843 404
rect 13877 402 13916 404
rect 13950 402 13989 404
rect 14023 402 14062 404
rect 14096 402 14135 404
rect 14169 402 14208 404
rect 14242 402 14281 404
rect 14315 402 14354 404
rect 14388 402 14427 404
rect 14461 402 14500 404
rect 14534 402 14573 404
rect 14607 402 14646 404
rect 14680 402 14719 404
rect 14753 402 14792 404
rect 14826 402 14866 404
rect 14900 402 14940 404
rect 14974 402 15014 404
rect 15048 402 15088 404
rect 15122 402 15162 404
rect 15196 402 15236 404
rect 15270 402 15310 404
rect 15344 402 15384 404
rect 15418 402 15458 404
rect 15492 402 15532 404
rect 15566 402 15606 404
rect 15640 402 15680 404
rect 15566 370 15577 402
rect 15640 370 15646 402
rect 15542 368 15577 370
rect 15611 368 15646 370
rect 15714 402 15754 404
rect 15788 402 15828 404
rect 15862 402 15902 404
rect 15936 402 15976 404
rect 16010 402 16050 404
rect 16084 402 16124 404
rect 16158 402 16198 404
rect 15714 370 15715 402
rect 15680 368 15715 370
rect 15749 370 15754 402
rect 15818 370 15828 402
rect 15887 370 15902 402
rect 15956 370 15976 402
rect 16025 370 16050 402
rect 16094 370 16124 402
rect 15749 368 15784 370
rect 15818 368 15853 370
rect 15887 368 15922 370
rect 15956 368 15991 370
rect 16025 368 16060 370
rect 16094 368 16129 370
rect 16163 368 16198 402
rect 16232 368 16332 404
rect 15542 334 16332 368
rect 15542 332 15577 334
rect 15611 332 15646 334
rect 15566 300 15577 332
rect 15640 300 15646 332
rect 15680 332 15715 334
rect 13366 298 13405 300
rect 13439 298 13478 300
rect 13512 298 13551 300
rect 13585 298 13624 300
rect 13658 298 13697 300
rect 13731 298 13770 300
rect 13804 298 13843 300
rect 13877 298 13916 300
rect 13950 298 13989 300
rect 14023 298 14062 300
rect 14096 298 14135 300
rect 14169 298 14208 300
rect 14242 298 14281 300
rect 14315 298 14354 300
rect 14388 298 14427 300
rect 14461 298 14500 300
rect 14534 298 14573 300
rect 14607 298 14646 300
rect 14680 298 14719 300
rect 14753 298 14792 300
rect 14826 298 14866 300
rect 14900 298 14940 300
rect 14974 298 15014 300
rect 15048 298 15088 300
rect 15122 298 15162 300
rect 15196 298 15236 300
rect 15270 298 15310 300
rect 15344 298 15384 300
rect 15418 298 15458 300
rect 15492 298 15532 300
rect 15566 298 15606 300
rect 15640 298 15680 300
rect 15714 300 15715 332
rect 15749 332 15784 334
rect 15818 332 15853 334
rect 15887 332 15922 334
rect 15956 332 15991 334
rect 16025 332 16060 334
rect 16094 332 16129 334
rect 15749 300 15754 332
rect 15818 300 15828 332
rect 15887 300 15902 332
rect 15956 300 15976 332
rect 16025 300 16050 332
rect 16094 300 16124 332
rect 16163 300 16198 334
rect 15714 298 15754 300
rect 15788 298 15828 300
rect 15862 298 15902 300
rect 15936 298 15976 300
rect 16010 298 16050 300
rect 16084 298 16124 300
rect 16158 298 16198 300
rect 16232 298 16332 334
rect 16474 368 16574 404
rect 16608 402 16648 404
rect 16682 402 16722 404
rect 16756 402 16796 404
rect 16830 402 16870 404
rect 16904 402 16944 404
rect 16978 402 17018 404
rect 17052 402 17092 404
rect 16608 368 16643 402
rect 16682 370 16712 402
rect 16756 370 16781 402
rect 16830 370 16850 402
rect 16904 370 16919 402
rect 16978 370 16988 402
rect 17052 370 17057 402
rect 16677 368 16712 370
rect 16746 368 16781 370
rect 16815 368 16850 370
rect 16884 368 16919 370
rect 16953 368 16988 370
rect 17022 368 17057 370
rect 17091 370 17092 402
rect 17126 402 17166 404
rect 17200 402 17240 404
rect 17274 402 17314 404
rect 17348 402 17388 404
rect 17422 402 17462 404
rect 17496 402 17536 404
rect 17570 402 17610 404
rect 17644 402 17684 404
rect 17718 402 17758 404
rect 17792 402 17832 404
rect 17866 402 17906 404
rect 17940 402 17980 404
rect 18014 402 18053 404
rect 18087 402 18126 404
rect 18160 402 18199 404
rect 18233 402 18272 404
rect 18306 402 18345 404
rect 18379 402 18418 404
rect 18452 402 18491 404
rect 18525 402 18564 404
rect 18598 402 18637 404
rect 18671 402 18710 404
rect 18744 402 18783 404
rect 18817 402 18856 404
rect 18890 402 18929 404
rect 18963 402 19002 404
rect 19036 402 19075 404
rect 19109 402 19148 404
rect 19182 402 19221 404
rect 19255 402 19294 404
rect 19328 402 19367 404
rect 19401 402 19440 404
rect 17091 368 17126 370
rect 17160 370 17166 402
rect 17229 370 17240 402
rect 17160 368 17195 370
rect 17229 368 17264 370
rect 16474 334 17264 368
rect 16474 298 16574 334
rect 16608 300 16643 334
rect 16677 332 16712 334
rect 16746 332 16781 334
rect 16815 332 16850 334
rect 16884 332 16919 334
rect 16953 332 16988 334
rect 17022 332 17057 334
rect 16682 300 16712 332
rect 16756 300 16781 332
rect 16830 300 16850 332
rect 16904 300 16919 332
rect 16978 300 16988 332
rect 17052 300 17057 332
rect 17091 332 17126 334
rect 17091 300 17092 332
rect 16608 298 16648 300
rect 16682 298 16722 300
rect 16756 298 16796 300
rect 16830 298 16870 300
rect 16904 298 16944 300
rect 16978 298 17018 300
rect 17052 298 17092 300
rect 17160 332 17195 334
rect 17229 332 17264 334
rect 17160 300 17166 332
rect 17229 300 17240 332
rect 17126 298 17166 300
rect 17200 298 17240 300
rect 17274 298 17314 300
rect 17348 298 17388 300
rect 17422 298 17462 300
rect 17496 298 17536 300
rect 17570 298 17610 300
rect 17644 298 17684 300
rect 17718 298 17758 300
rect 17792 298 17832 300
rect 17866 298 17906 300
rect 17940 298 17980 300
rect 18014 298 18053 300
rect 18087 298 18126 300
rect 18160 298 18199 300
rect 18233 298 18272 300
rect 18306 298 18345 300
rect 18379 298 18418 300
rect 18452 298 18491 300
rect 18525 298 18564 300
rect 18598 298 18637 300
rect 18671 298 18710 300
rect 18744 298 18783 300
rect 18817 298 18856 300
rect 18890 298 18929 300
rect 18963 298 19002 300
rect 19036 298 19075 300
rect 19109 298 19148 300
rect 19182 298 19221 300
rect 19255 298 19294 300
rect 19328 298 19367 300
rect 19401 298 19440 300
rect 19474 298 19574 404
rect 19838 393 19888 413
rect 19838 359 19882 393
rect 19922 379 19972 413
rect 19916 359 19972 379
rect 19838 343 19972 359
rect 19838 321 19888 343
rect -52 261 -46 295
rect -12 273 42 295
rect -12 261 -2 273
rect -52 239 -2 261
rect 32 261 42 273
rect 76 261 82 295
rect 32 239 82 261
rect -52 221 82 239
rect -52 187 -46 221
rect -12 203 42 221
rect -12 187 -2 203
rect -52 169 -2 187
rect 32 187 42 203
rect 76 187 82 221
rect 19838 287 19882 321
rect 19922 309 19972 343
rect 19916 287 19972 309
rect 19838 273 19972 287
rect 19838 249 19888 273
rect 19838 215 19882 249
rect 19922 239 19972 273
rect 19916 215 19972 239
rect 32 169 82 187
rect -52 147 82 169
rect -52 113 -46 147
rect -12 133 42 147
rect -12 113 -2 133
rect -52 99 -2 113
rect 32 113 42 133
rect 76 113 82 147
rect 182 196 216 212
rect 182 128 216 162
rect 3423 196 3457 212
rect 3423 128 3457 162
rect 32 99 82 113
rect -52 73 82 99
rect 216 94 240 114
rect 202 80 240 94
rect 3420 94 3423 114
rect 9907 196 9941 212
rect 9907 128 9941 162
rect 3457 94 3458 114
rect 3420 80 3458 94
rect 9904 94 9907 114
rect 16391 196 16425 212
rect 16391 128 16425 162
rect 9941 94 9942 114
rect 9904 80 9942 94
rect 16388 94 16391 114
rect 19622 196 19656 212
rect 19622 128 19656 162
rect 16425 94 16426 114
rect 16388 80 16426 94
rect 19838 203 19972 215
rect 19838 177 19888 203
rect 19838 143 19882 177
rect 19922 169 19972 203
rect 19916 143 19972 169
rect 19838 133 19972 143
rect 19656 94 19660 114
rect 19622 80 19660 94
rect 19838 105 19888 133
rect 182 78 216 80
rect 3423 78 3457 80
rect 9907 78 9941 80
rect 16391 78 16425 80
rect 19622 78 19656 80
rect -52 39 -46 73
rect -12 63 42 73
rect -12 39 -2 63
rect -52 29 -2 39
rect 32 39 42 63
rect 76 39 82 73
rect 32 29 82 39
rect -52 -1 82 29
rect -52 -35 -46 -1
rect -12 -7 42 -1
rect -12 -35 -2 -7
rect -52 -41 -2 -35
rect 32 -35 42 -7
rect 76 -35 82 -1
rect 19838 71 19882 105
rect 19922 99 19972 133
rect 19916 71 19972 99
rect 19838 63 19972 71
rect 19838 33 19888 63
rect 19838 -1 19882 33
rect 19922 29 19972 63
rect 19916 -1 19972 29
rect 19838 -7 19972 -1
rect 32 -41 82 -35
rect -52 -75 82 -41
rect -52 -109 -46 -75
rect -12 -77 42 -75
rect -12 -109 -2 -77
rect -52 -111 -2 -109
rect 32 -109 42 -77
rect 76 -109 82 -75
rect 32 -111 82 -109
rect -52 -147 82 -111
rect 264 -114 364 -8
rect 398 -10 437 -8
rect 471 -10 510 -8
rect 544 -10 583 -8
rect 617 -10 656 -8
rect 690 -10 729 -8
rect 763 -10 802 -8
rect 836 -10 875 -8
rect 909 -10 948 -8
rect 982 -10 1021 -8
rect 1055 -10 1094 -8
rect 1128 -10 1167 -8
rect 1201 -10 1240 -8
rect 1274 -10 1313 -8
rect 1347 -10 1386 -8
rect 1420 -10 1459 -8
rect 1493 -10 1532 -8
rect 1566 -10 1605 -8
rect 1639 -10 1678 -8
rect 1712 -10 1751 -8
rect 1785 -10 1824 -8
rect 1858 -10 1898 -8
rect 1932 -10 1972 -8
rect 2006 -10 2046 -8
rect 2080 -10 2120 -8
rect 2154 -10 2194 -8
rect 2228 -10 2268 -8
rect 2302 -10 2342 -8
rect 2376 -10 2416 -8
rect 2450 -10 2490 -8
rect 2524 -10 2564 -8
rect 2598 -10 2638 -8
rect 2672 -10 2712 -8
rect 2598 -42 2609 -10
rect 2672 -42 2678 -10
rect 2574 -44 2609 -42
rect 2643 -44 2678 -42
rect 2746 -10 2786 -8
rect 2820 -10 2860 -8
rect 2894 -10 2934 -8
rect 2968 -10 3008 -8
rect 3042 -10 3082 -8
rect 3116 -10 3156 -8
rect 3190 -10 3230 -8
rect 2746 -42 2747 -10
rect 2712 -44 2747 -42
rect 2781 -42 2786 -10
rect 2850 -42 2860 -10
rect 2919 -42 2934 -10
rect 2988 -42 3008 -10
rect 3057 -42 3082 -10
rect 3126 -42 3156 -10
rect 2781 -44 2816 -42
rect 2850 -44 2885 -42
rect 2919 -44 2954 -42
rect 2988 -44 3023 -42
rect 3057 -44 3092 -42
rect 3126 -44 3161 -42
rect 3195 -44 3230 -10
rect 3264 -44 3364 -8
rect 2574 -78 3364 -44
rect 2574 -80 2609 -78
rect 2643 -80 2678 -78
rect 2598 -112 2609 -80
rect 2672 -112 2678 -80
rect 2712 -80 2747 -78
rect 398 -114 437 -112
rect 471 -114 510 -112
rect 544 -114 583 -112
rect 617 -114 656 -112
rect 690 -114 729 -112
rect 763 -114 802 -112
rect 836 -114 875 -112
rect 909 -114 948 -112
rect 982 -114 1021 -112
rect 1055 -114 1094 -112
rect 1128 -114 1167 -112
rect 1201 -114 1240 -112
rect 1274 -114 1313 -112
rect 1347 -114 1386 -112
rect 1420 -114 1459 -112
rect 1493 -114 1532 -112
rect 1566 -114 1605 -112
rect 1639 -114 1678 -112
rect 1712 -114 1751 -112
rect 1785 -114 1824 -112
rect 1858 -114 1898 -112
rect 1932 -114 1972 -112
rect 2006 -114 2046 -112
rect 2080 -114 2120 -112
rect 2154 -114 2194 -112
rect 2228 -114 2268 -112
rect 2302 -114 2342 -112
rect 2376 -114 2416 -112
rect 2450 -114 2490 -112
rect 2524 -114 2564 -112
rect 2598 -114 2638 -112
rect 2672 -114 2712 -112
rect 2746 -112 2747 -80
rect 2781 -80 2816 -78
rect 2850 -80 2885 -78
rect 2919 -80 2954 -78
rect 2988 -80 3023 -78
rect 3057 -80 3092 -78
rect 3126 -80 3161 -78
rect 2781 -112 2786 -80
rect 2850 -112 2860 -80
rect 2919 -112 2934 -80
rect 2988 -112 3008 -80
rect 3057 -112 3082 -80
rect 3126 -112 3156 -80
rect 3195 -112 3230 -78
rect 2746 -114 2786 -112
rect 2820 -114 2860 -112
rect 2894 -114 2934 -112
rect 2968 -114 3008 -112
rect 3042 -114 3082 -112
rect 3116 -114 3156 -112
rect 3190 -114 3230 -112
rect 3264 -114 3364 -78
rect 3506 -44 3606 -8
rect 3640 -10 3680 -8
rect 3714 -10 3754 -8
rect 3788 -10 3828 -8
rect 3862 -10 3902 -8
rect 3936 -10 3976 -8
rect 4010 -10 4050 -8
rect 4084 -10 4124 -8
rect 3640 -44 3675 -10
rect 3714 -42 3744 -10
rect 3788 -42 3813 -10
rect 3862 -42 3882 -10
rect 3936 -42 3951 -10
rect 4010 -42 4020 -10
rect 4084 -42 4089 -10
rect 3709 -44 3744 -42
rect 3778 -44 3813 -42
rect 3847 -44 3882 -42
rect 3916 -44 3951 -42
rect 3985 -44 4020 -42
rect 4054 -44 4089 -42
rect 4123 -42 4124 -10
rect 4158 -10 4198 -8
rect 4232 -10 4272 -8
rect 4306 -10 4346 -8
rect 4380 -10 4420 -8
rect 4454 -10 4494 -8
rect 4528 -10 4568 -8
rect 4602 -10 4642 -8
rect 4676 -10 4716 -8
rect 4750 -10 4790 -8
rect 4824 -10 4864 -8
rect 4898 -10 4938 -8
rect 4972 -10 5012 -8
rect 5046 -10 5085 -8
rect 5119 -10 5158 -8
rect 5192 -10 5231 -8
rect 5265 -10 5304 -8
rect 5338 -10 5377 -8
rect 5411 -10 5450 -8
rect 5484 -10 5523 -8
rect 5557 -10 5596 -8
rect 5630 -10 5669 -8
rect 5703 -10 5742 -8
rect 5776 -10 5815 -8
rect 5849 -10 5888 -8
rect 5922 -10 5961 -8
rect 5995 -10 6034 -8
rect 6068 -10 6107 -8
rect 6141 -10 6180 -8
rect 6214 -10 6253 -8
rect 6287 -10 6326 -8
rect 6360 -10 6399 -8
rect 6433 -10 6472 -8
rect 4123 -44 4158 -42
rect 4192 -42 4198 -10
rect 4261 -42 4272 -10
rect 4192 -44 4227 -42
rect 4261 -44 4296 -42
rect 3506 -78 4296 -44
rect 3506 -114 3606 -78
rect 3640 -112 3675 -78
rect 3709 -80 3744 -78
rect 3778 -80 3813 -78
rect 3847 -80 3882 -78
rect 3916 -80 3951 -78
rect 3985 -80 4020 -78
rect 4054 -80 4089 -78
rect 3714 -112 3744 -80
rect 3788 -112 3813 -80
rect 3862 -112 3882 -80
rect 3936 -112 3951 -80
rect 4010 -112 4020 -80
rect 4084 -112 4089 -80
rect 4123 -80 4158 -78
rect 4123 -112 4124 -80
rect 3640 -114 3680 -112
rect 3714 -114 3754 -112
rect 3788 -114 3828 -112
rect 3862 -114 3902 -112
rect 3936 -114 3976 -112
rect 4010 -114 4050 -112
rect 4084 -114 4124 -112
rect 4192 -80 4227 -78
rect 4261 -80 4296 -78
rect 4192 -112 4198 -80
rect 4261 -112 4272 -80
rect 4158 -114 4198 -112
rect 4232 -114 4272 -112
rect 4306 -114 4346 -112
rect 4380 -114 4420 -112
rect 4454 -114 4494 -112
rect 4528 -114 4568 -112
rect 4602 -114 4642 -112
rect 4676 -114 4716 -112
rect 4750 -114 4790 -112
rect 4824 -114 4864 -112
rect 4898 -114 4938 -112
rect 4972 -114 5012 -112
rect 5046 -114 5085 -112
rect 5119 -114 5158 -112
rect 5192 -114 5231 -112
rect 5265 -114 5304 -112
rect 5338 -114 5377 -112
rect 5411 -114 5450 -112
rect 5484 -114 5523 -112
rect 5557 -114 5596 -112
rect 5630 -114 5669 -112
rect 5703 -114 5742 -112
rect 5776 -114 5815 -112
rect 5849 -114 5888 -112
rect 5922 -114 5961 -112
rect 5995 -114 6034 -112
rect 6068 -114 6107 -112
rect 6141 -114 6180 -112
rect 6214 -114 6253 -112
rect 6287 -114 6326 -112
rect 6360 -114 6399 -112
rect 6433 -114 6472 -112
rect 6506 -114 6606 -8
rect 6748 -114 6848 -8
rect 6882 -10 6921 -8
rect 6955 -10 6994 -8
rect 7028 -10 7067 -8
rect 7101 -10 7140 -8
rect 7174 -10 7213 -8
rect 7247 -10 7286 -8
rect 7320 -10 7359 -8
rect 7393 -10 7432 -8
rect 7466 -10 7505 -8
rect 7539 -10 7578 -8
rect 7612 -10 7651 -8
rect 7685 -10 7724 -8
rect 7758 -10 7797 -8
rect 7831 -10 7870 -8
rect 7904 -10 7943 -8
rect 7977 -10 8016 -8
rect 8050 -10 8089 -8
rect 8123 -10 8162 -8
rect 8196 -10 8235 -8
rect 8269 -10 8308 -8
rect 8342 -10 8382 -8
rect 8416 -10 8456 -8
rect 8490 -10 8530 -8
rect 8564 -10 8604 -8
rect 8638 -10 8678 -8
rect 8712 -10 8752 -8
rect 8786 -10 8826 -8
rect 8860 -10 8900 -8
rect 8934 -10 8974 -8
rect 9008 -10 9048 -8
rect 9082 -10 9122 -8
rect 9156 -10 9196 -8
rect 9082 -42 9093 -10
rect 9156 -42 9162 -10
rect 9058 -44 9093 -42
rect 9127 -44 9162 -42
rect 9230 -10 9270 -8
rect 9304 -10 9344 -8
rect 9378 -10 9418 -8
rect 9452 -10 9492 -8
rect 9526 -10 9566 -8
rect 9600 -10 9640 -8
rect 9674 -10 9714 -8
rect 9230 -42 9231 -10
rect 9196 -44 9231 -42
rect 9265 -42 9270 -10
rect 9334 -42 9344 -10
rect 9403 -42 9418 -10
rect 9472 -42 9492 -10
rect 9541 -42 9566 -10
rect 9610 -42 9640 -10
rect 9265 -44 9300 -42
rect 9334 -44 9369 -42
rect 9403 -44 9438 -42
rect 9472 -44 9507 -42
rect 9541 -44 9576 -42
rect 9610 -44 9645 -42
rect 9679 -44 9714 -10
rect 9748 -44 9848 -8
rect 9058 -78 9848 -44
rect 9058 -80 9093 -78
rect 9127 -80 9162 -78
rect 9082 -112 9093 -80
rect 9156 -112 9162 -80
rect 9196 -80 9231 -78
rect 6882 -114 6921 -112
rect 6955 -114 6994 -112
rect 7028 -114 7067 -112
rect 7101 -114 7140 -112
rect 7174 -114 7213 -112
rect 7247 -114 7286 -112
rect 7320 -114 7359 -112
rect 7393 -114 7432 -112
rect 7466 -114 7505 -112
rect 7539 -114 7578 -112
rect 7612 -114 7651 -112
rect 7685 -114 7724 -112
rect 7758 -114 7797 -112
rect 7831 -114 7870 -112
rect 7904 -114 7943 -112
rect 7977 -114 8016 -112
rect 8050 -114 8089 -112
rect 8123 -114 8162 -112
rect 8196 -114 8235 -112
rect 8269 -114 8308 -112
rect 8342 -114 8382 -112
rect 8416 -114 8456 -112
rect 8490 -114 8530 -112
rect 8564 -114 8604 -112
rect 8638 -114 8678 -112
rect 8712 -114 8752 -112
rect 8786 -114 8826 -112
rect 8860 -114 8900 -112
rect 8934 -114 8974 -112
rect 9008 -114 9048 -112
rect 9082 -114 9122 -112
rect 9156 -114 9196 -112
rect 9230 -112 9231 -80
rect 9265 -80 9300 -78
rect 9334 -80 9369 -78
rect 9403 -80 9438 -78
rect 9472 -80 9507 -78
rect 9541 -80 9576 -78
rect 9610 -80 9645 -78
rect 9265 -112 9270 -80
rect 9334 -112 9344 -80
rect 9403 -112 9418 -80
rect 9472 -112 9492 -80
rect 9541 -112 9566 -80
rect 9610 -112 9640 -80
rect 9679 -112 9714 -78
rect 9230 -114 9270 -112
rect 9304 -114 9344 -112
rect 9378 -114 9418 -112
rect 9452 -114 9492 -112
rect 9526 -114 9566 -112
rect 9600 -114 9640 -112
rect 9674 -114 9714 -112
rect 9748 -114 9848 -78
rect 9990 -44 10090 -8
rect 10124 -10 10164 -8
rect 10198 -10 10238 -8
rect 10272 -10 10312 -8
rect 10346 -10 10386 -8
rect 10420 -10 10460 -8
rect 10494 -10 10534 -8
rect 10568 -10 10608 -8
rect 10124 -44 10159 -10
rect 10198 -42 10228 -10
rect 10272 -42 10297 -10
rect 10346 -42 10366 -10
rect 10420 -42 10435 -10
rect 10494 -42 10504 -10
rect 10568 -42 10573 -10
rect 10193 -44 10228 -42
rect 10262 -44 10297 -42
rect 10331 -44 10366 -42
rect 10400 -44 10435 -42
rect 10469 -44 10504 -42
rect 10538 -44 10573 -42
rect 10607 -42 10608 -10
rect 10642 -10 10682 -8
rect 10716 -10 10756 -8
rect 10790 -10 10830 -8
rect 10864 -10 10904 -8
rect 10938 -10 10978 -8
rect 11012 -10 11052 -8
rect 11086 -10 11126 -8
rect 11160 -10 11200 -8
rect 11234 -10 11274 -8
rect 11308 -10 11348 -8
rect 11382 -10 11422 -8
rect 11456 -10 11496 -8
rect 11530 -10 11569 -8
rect 11603 -10 11642 -8
rect 11676 -10 11715 -8
rect 11749 -10 11788 -8
rect 11822 -10 11861 -8
rect 11895 -10 11934 -8
rect 11968 -10 12007 -8
rect 12041 -10 12080 -8
rect 12114 -10 12153 -8
rect 12187 -10 12226 -8
rect 12260 -10 12299 -8
rect 12333 -10 12372 -8
rect 12406 -10 12445 -8
rect 12479 -10 12518 -8
rect 12552 -10 12591 -8
rect 12625 -10 12664 -8
rect 12698 -10 12737 -8
rect 12771 -10 12810 -8
rect 12844 -10 12883 -8
rect 12917 -10 12956 -8
rect 10607 -44 10642 -42
rect 10676 -42 10682 -10
rect 10745 -42 10756 -10
rect 10676 -44 10711 -42
rect 10745 -44 10780 -42
rect 9990 -78 10780 -44
rect 9990 -114 10090 -78
rect 10124 -112 10159 -78
rect 10193 -80 10228 -78
rect 10262 -80 10297 -78
rect 10331 -80 10366 -78
rect 10400 -80 10435 -78
rect 10469 -80 10504 -78
rect 10538 -80 10573 -78
rect 10198 -112 10228 -80
rect 10272 -112 10297 -80
rect 10346 -112 10366 -80
rect 10420 -112 10435 -80
rect 10494 -112 10504 -80
rect 10568 -112 10573 -80
rect 10607 -80 10642 -78
rect 10607 -112 10608 -80
rect 10124 -114 10164 -112
rect 10198 -114 10238 -112
rect 10272 -114 10312 -112
rect 10346 -114 10386 -112
rect 10420 -114 10460 -112
rect 10494 -114 10534 -112
rect 10568 -114 10608 -112
rect 10676 -80 10711 -78
rect 10745 -80 10780 -78
rect 10676 -112 10682 -80
rect 10745 -112 10756 -80
rect 10642 -114 10682 -112
rect 10716 -114 10756 -112
rect 10790 -114 10830 -112
rect 10864 -114 10904 -112
rect 10938 -114 10978 -112
rect 11012 -114 11052 -112
rect 11086 -114 11126 -112
rect 11160 -114 11200 -112
rect 11234 -114 11274 -112
rect 11308 -114 11348 -112
rect 11382 -114 11422 -112
rect 11456 -114 11496 -112
rect 11530 -114 11569 -112
rect 11603 -114 11642 -112
rect 11676 -114 11715 -112
rect 11749 -114 11788 -112
rect 11822 -114 11861 -112
rect 11895 -114 11934 -112
rect 11968 -114 12007 -112
rect 12041 -114 12080 -112
rect 12114 -114 12153 -112
rect 12187 -114 12226 -112
rect 12260 -114 12299 -112
rect 12333 -114 12372 -112
rect 12406 -114 12445 -112
rect 12479 -114 12518 -112
rect 12552 -114 12591 -112
rect 12625 -114 12664 -112
rect 12698 -114 12737 -112
rect 12771 -114 12810 -112
rect 12844 -114 12883 -112
rect 12917 -114 12956 -112
rect 12990 -114 13090 -8
rect 13232 -114 13332 -8
rect 13366 -10 13405 -8
rect 13439 -10 13478 -8
rect 13512 -10 13551 -8
rect 13585 -10 13624 -8
rect 13658 -10 13697 -8
rect 13731 -10 13770 -8
rect 13804 -10 13843 -8
rect 13877 -10 13916 -8
rect 13950 -10 13989 -8
rect 14023 -10 14062 -8
rect 14096 -10 14135 -8
rect 14169 -10 14208 -8
rect 14242 -10 14281 -8
rect 14315 -10 14354 -8
rect 14388 -10 14427 -8
rect 14461 -10 14500 -8
rect 14534 -10 14573 -8
rect 14607 -10 14646 -8
rect 14680 -10 14719 -8
rect 14753 -10 14792 -8
rect 14826 -10 14866 -8
rect 14900 -10 14940 -8
rect 14974 -10 15014 -8
rect 15048 -10 15088 -8
rect 15122 -10 15162 -8
rect 15196 -10 15236 -8
rect 15270 -10 15310 -8
rect 15344 -10 15384 -8
rect 15418 -10 15458 -8
rect 15492 -10 15532 -8
rect 15566 -10 15606 -8
rect 15640 -10 15680 -8
rect 15566 -42 15577 -10
rect 15640 -42 15646 -10
rect 15542 -44 15577 -42
rect 15611 -44 15646 -42
rect 15714 -10 15754 -8
rect 15788 -10 15828 -8
rect 15862 -10 15902 -8
rect 15936 -10 15976 -8
rect 16010 -10 16050 -8
rect 16084 -10 16124 -8
rect 16158 -10 16198 -8
rect 15714 -42 15715 -10
rect 15680 -44 15715 -42
rect 15749 -42 15754 -10
rect 15818 -42 15828 -10
rect 15887 -42 15902 -10
rect 15956 -42 15976 -10
rect 16025 -42 16050 -10
rect 16094 -42 16124 -10
rect 15749 -44 15784 -42
rect 15818 -44 15853 -42
rect 15887 -44 15922 -42
rect 15956 -44 15991 -42
rect 16025 -44 16060 -42
rect 16094 -44 16129 -42
rect 16163 -44 16198 -10
rect 16232 -44 16332 -8
rect 15542 -78 16332 -44
rect 15542 -80 15577 -78
rect 15611 -80 15646 -78
rect 15566 -112 15577 -80
rect 15640 -112 15646 -80
rect 15680 -80 15715 -78
rect 13366 -114 13405 -112
rect 13439 -114 13478 -112
rect 13512 -114 13551 -112
rect 13585 -114 13624 -112
rect 13658 -114 13697 -112
rect 13731 -114 13770 -112
rect 13804 -114 13843 -112
rect 13877 -114 13916 -112
rect 13950 -114 13989 -112
rect 14023 -114 14062 -112
rect 14096 -114 14135 -112
rect 14169 -114 14208 -112
rect 14242 -114 14281 -112
rect 14315 -114 14354 -112
rect 14388 -114 14427 -112
rect 14461 -114 14500 -112
rect 14534 -114 14573 -112
rect 14607 -114 14646 -112
rect 14680 -114 14719 -112
rect 14753 -114 14792 -112
rect 14826 -114 14866 -112
rect 14900 -114 14940 -112
rect 14974 -114 15014 -112
rect 15048 -114 15088 -112
rect 15122 -114 15162 -112
rect 15196 -114 15236 -112
rect 15270 -114 15310 -112
rect 15344 -114 15384 -112
rect 15418 -114 15458 -112
rect 15492 -114 15532 -112
rect 15566 -114 15606 -112
rect 15640 -114 15680 -112
rect 15714 -112 15715 -80
rect 15749 -80 15784 -78
rect 15818 -80 15853 -78
rect 15887 -80 15922 -78
rect 15956 -80 15991 -78
rect 16025 -80 16060 -78
rect 16094 -80 16129 -78
rect 15749 -112 15754 -80
rect 15818 -112 15828 -80
rect 15887 -112 15902 -80
rect 15956 -112 15976 -80
rect 16025 -112 16050 -80
rect 16094 -112 16124 -80
rect 16163 -112 16198 -78
rect 15714 -114 15754 -112
rect 15788 -114 15828 -112
rect 15862 -114 15902 -112
rect 15936 -114 15976 -112
rect 16010 -114 16050 -112
rect 16084 -114 16124 -112
rect 16158 -114 16198 -112
rect 16232 -114 16332 -78
rect 16474 -44 16574 -8
rect 16608 -10 16648 -8
rect 16682 -10 16722 -8
rect 16756 -10 16796 -8
rect 16830 -10 16870 -8
rect 16904 -10 16944 -8
rect 16978 -10 17018 -8
rect 17052 -10 17092 -8
rect 16608 -44 16643 -10
rect 16682 -42 16712 -10
rect 16756 -42 16781 -10
rect 16830 -42 16850 -10
rect 16904 -42 16919 -10
rect 16978 -42 16988 -10
rect 17052 -42 17057 -10
rect 16677 -44 16712 -42
rect 16746 -44 16781 -42
rect 16815 -44 16850 -42
rect 16884 -44 16919 -42
rect 16953 -44 16988 -42
rect 17022 -44 17057 -42
rect 17091 -42 17092 -10
rect 17126 -10 17166 -8
rect 17200 -10 17240 -8
rect 17274 -10 17314 -8
rect 17348 -10 17388 -8
rect 17422 -10 17462 -8
rect 17496 -10 17536 -8
rect 17570 -10 17610 -8
rect 17644 -10 17684 -8
rect 17718 -10 17758 -8
rect 17792 -10 17832 -8
rect 17866 -10 17906 -8
rect 17940 -10 17980 -8
rect 18014 -10 18053 -8
rect 18087 -10 18126 -8
rect 18160 -10 18199 -8
rect 18233 -10 18272 -8
rect 18306 -10 18345 -8
rect 18379 -10 18418 -8
rect 18452 -10 18491 -8
rect 18525 -10 18564 -8
rect 18598 -10 18637 -8
rect 18671 -10 18710 -8
rect 18744 -10 18783 -8
rect 18817 -10 18856 -8
rect 18890 -10 18929 -8
rect 18963 -10 19002 -8
rect 19036 -10 19075 -8
rect 19109 -10 19148 -8
rect 19182 -10 19221 -8
rect 19255 -10 19294 -8
rect 19328 -10 19367 -8
rect 19401 -10 19440 -8
rect 17091 -44 17126 -42
rect 17160 -42 17166 -10
rect 17229 -42 17240 -10
rect 17160 -44 17195 -42
rect 17229 -44 17264 -42
rect 16474 -78 17264 -44
rect 16474 -114 16574 -78
rect 16608 -112 16643 -78
rect 16677 -80 16712 -78
rect 16746 -80 16781 -78
rect 16815 -80 16850 -78
rect 16884 -80 16919 -78
rect 16953 -80 16988 -78
rect 17022 -80 17057 -78
rect 16682 -112 16712 -80
rect 16756 -112 16781 -80
rect 16830 -112 16850 -80
rect 16904 -112 16919 -80
rect 16978 -112 16988 -80
rect 17052 -112 17057 -80
rect 17091 -80 17126 -78
rect 17091 -112 17092 -80
rect 16608 -114 16648 -112
rect 16682 -114 16722 -112
rect 16756 -114 16796 -112
rect 16830 -114 16870 -112
rect 16904 -114 16944 -112
rect 16978 -114 17018 -112
rect 17052 -114 17092 -112
rect 17160 -80 17195 -78
rect 17229 -80 17264 -78
rect 17160 -112 17166 -80
rect 17229 -112 17240 -80
rect 17126 -114 17166 -112
rect 17200 -114 17240 -112
rect 17274 -114 17314 -112
rect 17348 -114 17388 -112
rect 17422 -114 17462 -112
rect 17496 -114 17536 -112
rect 17570 -114 17610 -112
rect 17644 -114 17684 -112
rect 17718 -114 17758 -112
rect 17792 -114 17832 -112
rect 17866 -114 17906 -112
rect 17940 -114 17980 -112
rect 18014 -114 18053 -112
rect 18087 -114 18126 -112
rect 18160 -114 18199 -112
rect 18233 -114 18272 -112
rect 18306 -114 18345 -112
rect 18379 -114 18418 -112
rect 18452 -114 18491 -112
rect 18525 -114 18564 -112
rect 18598 -114 18637 -112
rect 18671 -114 18710 -112
rect 18744 -114 18783 -112
rect 18817 -114 18856 -112
rect 18890 -114 18929 -112
rect 18963 -114 19002 -112
rect 19036 -114 19075 -112
rect 19109 -114 19148 -112
rect 19182 -114 19221 -112
rect 19255 -114 19294 -112
rect 19328 -114 19367 -112
rect 19401 -114 19440 -112
rect 19474 -114 19574 -8
rect 19838 -39 19888 -7
rect 19838 -73 19882 -39
rect 19922 -41 19972 -7
rect 19916 -73 19972 -41
rect 19838 -77 19972 -73
rect 19838 -111 19888 -77
rect 19922 -111 19972 -77
rect -52 -149 -2 -147
rect -52 -183 -46 -149
rect -12 -181 -2 -149
rect 32 -149 82 -147
rect 32 -181 42 -149
rect -12 -183 42 -181
rect 76 -183 82 -149
rect -52 -209 82 -183
rect 19838 -145 19882 -111
rect 19916 -145 19972 -111
rect 19838 -147 19972 -145
rect 19838 -181 19888 -147
rect 19922 -181 19972 -147
rect 19838 -209 19972 -181
rect -415 -238 20466 -209
rect -415 -272 8 -238
rect 42 -272 48 -238
rect 114 -272 116 -238
rect 150 -272 152 -238
rect 218 -272 224 -238
rect 286 -272 296 -238
rect 354 -272 368 -238
rect 422 -272 440 -238
rect 490 -272 512 -238
rect 558 -272 584 -238
rect 626 -272 656 -238
rect 694 -272 728 -238
rect 762 -272 796 -238
rect 834 -272 864 -238
rect 906 -272 932 -238
rect 978 -272 1000 -238
rect 1050 -272 1068 -238
rect 1122 -272 1136 -238
rect 1194 -272 1204 -238
rect 1266 -272 1272 -238
rect 1338 -272 1340 -238
rect 1374 -272 1376 -238
rect 1442 -272 1448 -238
rect 1510 -272 1520 -238
rect 1578 -272 1592 -238
rect 1646 -272 1664 -238
rect 1714 -272 1736 -238
rect 1782 -272 1808 -238
rect 1850 -272 1880 -238
rect 1918 -272 1952 -238
rect 1986 -272 2020 -238
rect 2058 -272 2088 -238
rect 2130 -272 2156 -238
rect 2202 -272 2224 -238
rect 2274 -272 2292 -238
rect 2346 -272 2360 -238
rect 2418 -272 2428 -238
rect 2490 -272 2496 -238
rect 2562 -272 2564 -238
rect 2598 -272 2600 -238
rect 2666 -272 2672 -238
rect 2734 -272 2744 -238
rect 2802 -272 2816 -238
rect 2870 -272 2888 -238
rect 2938 -272 2960 -238
rect 3006 -272 3032 -238
rect 3074 -272 3104 -238
rect 3142 -272 3176 -238
rect 3210 -272 3244 -238
rect 3282 -272 3312 -238
rect 3354 -272 3380 -238
rect 3426 -272 3448 -238
rect 3498 -272 3516 -238
rect 3570 -272 3584 -238
rect 3642 -272 3652 -238
rect 3714 -272 3720 -238
rect 3786 -272 3788 -238
rect 3822 -272 3824 -238
rect 3890 -272 3896 -238
rect 3958 -272 3968 -238
rect 4026 -272 4040 -238
rect 4094 -272 4112 -238
rect 4162 -272 4184 -238
rect 4230 -272 4256 -238
rect 4298 -272 4328 -238
rect 4366 -272 4400 -238
rect 4434 -272 4468 -238
rect 4506 -272 4536 -238
rect 4578 -272 4604 -238
rect 4650 -272 4672 -238
rect 4722 -272 4740 -238
rect 4794 -272 4808 -238
rect 4866 -272 4876 -238
rect 4938 -272 4944 -238
rect 5010 -272 5012 -238
rect 5046 -272 5048 -238
rect 5114 -272 5120 -238
rect 5182 -272 5192 -238
rect 5250 -272 5264 -238
rect 5318 -272 5336 -238
rect 5386 -272 5408 -238
rect 5454 -272 5480 -238
rect 5522 -272 5552 -238
rect 5590 -272 5624 -238
rect 5658 -272 5692 -238
rect 5730 -272 5760 -238
rect 5802 -272 5828 -238
rect 5874 -272 5896 -238
rect 5946 -272 5964 -238
rect 6018 -272 6032 -238
rect 6090 -272 6100 -238
rect 6162 -272 6168 -238
rect 6234 -272 6236 -238
rect 6270 -272 6272 -238
rect 6338 -272 6344 -238
rect 6406 -272 6416 -238
rect 6474 -272 6488 -238
rect 6542 -272 6560 -238
rect 6610 -272 6632 -238
rect 6678 -272 6704 -238
rect 6746 -272 6776 -238
rect 6814 -272 6848 -238
rect 6882 -272 6916 -238
rect 6954 -272 6984 -238
rect 7026 -272 7052 -238
rect 7098 -272 7120 -238
rect 7170 -272 7188 -238
rect 7242 -272 7256 -238
rect 7314 -272 7324 -238
rect 7386 -272 7392 -238
rect 7458 -272 7460 -238
rect 7494 -272 7496 -238
rect 7562 -272 7568 -238
rect 7630 -272 7640 -238
rect 7698 -272 7712 -238
rect 7766 -272 7784 -238
rect 7834 -272 7856 -238
rect 7902 -272 7928 -238
rect 7970 -272 8000 -238
rect 8038 -272 8072 -238
rect 8106 -272 8140 -238
rect 8178 -272 8208 -238
rect 8250 -272 8276 -238
rect 8322 -272 8344 -238
rect 8394 -272 8412 -238
rect 8466 -272 8480 -238
rect 8538 -272 8548 -238
rect 8610 -272 8616 -238
rect 8682 -272 8684 -238
rect 8718 -272 8720 -238
rect 8786 -272 8792 -238
rect 8854 -272 8864 -238
rect 8922 -272 8936 -238
rect 8990 -272 9008 -238
rect 9058 -272 9080 -238
rect 9126 -272 9152 -238
rect 9194 -272 9224 -238
rect 9262 -272 9296 -238
rect 9330 -272 9364 -238
rect 9402 -272 9432 -238
rect 9474 -272 9500 -238
rect 9546 -272 9568 -238
rect 9618 -272 9636 -238
rect 9690 -272 9704 -238
rect 9762 -272 9772 -238
rect 9834 -272 9840 -238
rect 9906 -272 9908 -238
rect 9942 -272 9944 -238
rect 10010 -272 10016 -238
rect 10078 -272 10088 -238
rect 10146 -272 10160 -238
rect 10214 -272 10232 -238
rect 10282 -272 10304 -238
rect 10350 -272 10376 -238
rect 10418 -272 10448 -238
rect 10486 -272 10520 -238
rect 10554 -272 10588 -238
rect 10626 -272 10656 -238
rect 10698 -272 10724 -238
rect 10770 -272 10792 -238
rect 10842 -272 10860 -238
rect 10914 -272 10928 -238
rect 10986 -272 10996 -238
rect 11058 -272 11064 -238
rect 11130 -272 11132 -238
rect 11166 -272 11168 -238
rect 11234 -272 11240 -238
rect 11302 -272 11312 -238
rect 11370 -272 11384 -238
rect 11438 -272 11456 -238
rect 11506 -272 11528 -238
rect 11574 -272 11600 -238
rect 11642 -272 11672 -238
rect 11710 -272 11744 -238
rect 11778 -272 11812 -238
rect 11850 -272 11880 -238
rect 11922 -272 11948 -238
rect 11994 -272 12016 -238
rect 12066 -272 12084 -238
rect 12138 -272 12152 -238
rect 12210 -272 12220 -238
rect 12282 -272 12288 -238
rect 12354 -272 12356 -238
rect 12390 -272 12392 -238
rect 12458 -272 12464 -238
rect 12526 -272 12536 -238
rect 12594 -272 12608 -238
rect 12662 -272 12680 -238
rect 12730 -272 12752 -238
rect 12798 -272 12824 -238
rect 12866 -272 12896 -238
rect 12934 -272 12968 -238
rect 13002 -272 13036 -238
rect 13074 -272 13104 -238
rect 13146 -272 13172 -238
rect 13218 -272 13240 -238
rect 13290 -272 13308 -238
rect 13362 -272 13376 -238
rect 13434 -272 13444 -238
rect 13506 -272 13512 -238
rect 13578 -272 13580 -238
rect 13614 -272 13616 -238
rect 13682 -272 13688 -238
rect 13750 -272 13760 -238
rect 13818 -272 13832 -238
rect 13886 -272 13904 -238
rect 13954 -272 13976 -238
rect 14022 -272 14048 -238
rect 14090 -272 14120 -238
rect 14158 -272 14192 -238
rect 14226 -272 14260 -238
rect 14298 -272 14328 -238
rect 14370 -272 14396 -238
rect 14442 -272 14464 -238
rect 14514 -272 14532 -238
rect 14586 -272 14600 -238
rect 14658 -272 14668 -238
rect 14730 -272 14736 -238
rect 14802 -272 14804 -238
rect 14838 -272 14840 -238
rect 14906 -272 14912 -238
rect 14974 -272 14984 -238
rect 15042 -272 15056 -238
rect 15110 -272 15128 -238
rect 15178 -272 15200 -238
rect 15246 -272 15272 -238
rect 15314 -272 15344 -238
rect 15382 -272 15416 -238
rect 15450 -272 15484 -238
rect 15522 -272 15552 -238
rect 15594 -272 15620 -238
rect 15666 -272 15688 -238
rect 15738 -272 15756 -238
rect 15810 -272 15824 -238
rect 15882 -272 15892 -238
rect 15954 -272 15960 -238
rect 16026 -272 16028 -238
rect 16062 -272 16064 -238
rect 16130 -272 16136 -238
rect 16198 -272 16208 -238
rect 16266 -272 16280 -238
rect 16334 -272 16352 -238
rect 16402 -272 16424 -238
rect 16470 -272 16496 -238
rect 16538 -272 16568 -238
rect 16606 -272 16640 -238
rect 16674 -272 16708 -238
rect 16746 -272 16776 -238
rect 16818 -272 16844 -238
rect 16890 -272 16912 -238
rect 16962 -272 16980 -238
rect 17034 -272 17048 -238
rect 17106 -272 17116 -238
rect 17178 -272 17184 -238
rect 17250 -272 17252 -238
rect 17286 -272 17288 -238
rect 17354 -272 17360 -238
rect 17422 -272 17432 -238
rect 17490 -272 17504 -238
rect 17558 -272 17576 -238
rect 17626 -272 17648 -238
rect 17694 -272 17720 -238
rect 17762 -272 17792 -238
rect 17830 -272 17864 -238
rect 17898 -272 17932 -238
rect 17970 -272 18000 -238
rect 18042 -272 18068 -238
rect 18114 -272 18136 -238
rect 18186 -272 18204 -238
rect 18258 -272 18272 -238
rect 18330 -272 18340 -238
rect 18402 -272 18408 -238
rect 18474 -272 18476 -238
rect 18510 -272 18513 -238
rect 18578 -272 18586 -238
rect 18646 -272 18659 -238
rect 18714 -272 18732 -238
rect 18782 -272 18805 -238
rect 18850 -272 18878 -238
rect 18918 -272 18951 -238
rect 18986 -272 19020 -238
rect 19058 -272 19088 -238
rect 19131 -272 19156 -238
rect 19204 -272 19224 -238
rect 19277 -272 19292 -238
rect 19350 -272 19360 -238
rect 19423 -272 19428 -238
rect 19530 -272 19535 -238
rect 19598 -272 19608 -238
rect 19666 -272 19681 -238
rect 19734 -272 19754 -238
rect 19802 -272 19827 -238
rect 19870 -272 19904 -238
rect 19938 -272 20466 -238
rect -415 -379 20466 -272
<< viali >>
rect -2040 14517 -2006 14521
rect -1967 14517 -1933 14521
rect -1894 14517 -1860 14521
rect -1821 14517 -1787 14521
rect -1748 14517 -1714 14521
rect -1675 14517 -1641 14521
rect -1601 14517 -1567 14521
rect -1527 14517 -1493 14521
rect -1453 14517 -1419 14521
rect -1379 14517 -1345 14521
rect -1305 14517 -1271 14521
rect -1231 14517 -1197 14521
rect -1157 14517 -1123 14521
rect -1083 14517 -1049 14521
rect -1009 14517 -975 14521
rect -935 14517 -901 14521
rect -861 14517 -827 14521
rect -787 14517 -753 14521
rect -713 14517 -679 14521
rect -2040 14487 -2006 14517
rect -1967 14487 -1933 14517
rect -1894 14487 -1860 14517
rect -1821 14487 -1787 14517
rect -1748 14487 -1714 14517
rect -1675 14487 -1641 14517
rect -1601 14487 -1599 14517
rect -1599 14487 -1567 14517
rect -1527 14487 -1495 14517
rect -1495 14487 -1493 14517
rect -1453 14487 -1426 14517
rect -1426 14487 -1419 14517
rect -1379 14487 -1357 14517
rect -1357 14487 -1345 14517
rect -1305 14487 -1288 14517
rect -1288 14487 -1271 14517
rect -1231 14487 -1219 14517
rect -1219 14487 -1197 14517
rect -1157 14487 -1150 14517
rect -1150 14487 -1123 14517
rect -1083 14487 -1081 14517
rect -1081 14487 -1049 14517
rect -1009 14487 -978 14517
rect -978 14487 -975 14517
rect -935 14487 -909 14517
rect -909 14487 -901 14517
rect -861 14487 -840 14517
rect -840 14487 -827 14517
rect -787 14487 -771 14517
rect -771 14487 -753 14517
rect -713 14487 -679 14517
rect -2113 14415 -2109 14449
rect -2109 14415 -2079 14449
rect -2041 14415 -2007 14449
rect -1967 14415 -1933 14449
rect -1894 14415 -1860 14449
rect -1821 14415 -1787 14449
rect -1748 14415 -1714 14449
rect -1675 14415 -1641 14449
rect -1601 14415 -1599 14449
rect -1599 14415 -1567 14449
rect -1527 14415 -1495 14449
rect -1495 14415 -1493 14449
rect -1453 14415 -1426 14449
rect -1426 14415 -1419 14449
rect -1379 14415 -1357 14449
rect -1357 14415 -1345 14449
rect -1305 14415 -1288 14449
rect -1288 14415 -1271 14449
rect -1231 14415 -1219 14449
rect -1219 14415 -1197 14449
rect -1157 14415 -1150 14449
rect -1150 14415 -1123 14449
rect -1083 14415 -1081 14449
rect -1081 14415 -1049 14449
rect -1009 14415 -978 14449
rect -978 14415 -975 14449
rect -935 14415 -909 14449
rect -909 14415 -901 14449
rect -861 14415 -840 14449
rect -840 14415 -827 14449
rect -787 14415 -771 14449
rect -771 14415 -753 14449
rect -713 14415 -679 14449
rect -2113 14346 -2109 14376
rect -2109 14346 -2079 14376
rect -2041 14346 -2007 14376
rect -1969 14347 -1935 14377
rect -1896 14347 -1862 14377
rect -1823 14347 -1789 14377
rect -1749 14347 -1715 14377
rect -1675 14347 -1641 14377
rect -1601 14347 -1599 14377
rect -1599 14347 -1567 14377
rect -1527 14347 -1495 14377
rect -1495 14347 -1493 14377
rect -1453 14347 -1426 14377
rect -1426 14347 -1419 14377
rect -1379 14347 -1357 14377
rect -1357 14347 -1345 14377
rect -1305 14347 -1288 14377
rect -1288 14347 -1271 14377
rect -1231 14347 -1219 14377
rect -1219 14347 -1197 14377
rect -1157 14347 -1150 14377
rect -1150 14347 -1123 14377
rect -1083 14347 -1081 14377
rect -1081 14347 -1049 14377
rect -1009 14347 -978 14377
rect -978 14347 -975 14377
rect -935 14347 -909 14377
rect -909 14347 -901 14377
rect -861 14347 -840 14377
rect -840 14347 -827 14377
rect -787 14347 -771 14377
rect -771 14347 -753 14377
rect -713 14347 -679 14377
rect -2113 14342 -2079 14346
rect -2041 14342 -2007 14346
rect -1969 14343 -1935 14347
rect -1896 14343 -1862 14347
rect -1823 14343 -1789 14347
rect -1749 14343 -1715 14347
rect -1675 14343 -1641 14347
rect -1601 14343 -1567 14347
rect -1527 14343 -1493 14347
rect -1453 14343 -1419 14347
rect -1379 14343 -1345 14347
rect -1305 14343 -1271 14347
rect -1231 14343 -1197 14347
rect -1157 14343 -1123 14347
rect -1083 14343 -1049 14347
rect -1009 14343 -975 14347
rect -935 14343 -901 14347
rect -861 14343 -827 14347
rect -787 14343 -753 14347
rect -713 14343 -679 14347
rect -2113 14277 -2109 14303
rect -2109 14277 -2079 14303
rect -2041 14277 -2007 14303
rect -1969 14278 -1939 14304
rect -1939 14278 -1935 14304
rect -2113 14269 -2079 14277
rect -2041 14269 -2007 14277
rect -1969 14270 -1935 14278
rect -2113 14208 -2109 14230
rect -2109 14208 -2079 14230
rect -2041 14208 -2007 14230
rect -1969 14209 -1939 14231
rect -1939 14209 -1935 14231
rect -2113 14196 -2079 14208
rect -2041 14196 -2007 14208
rect -1969 14197 -1935 14209
rect -2113 14139 -2109 14157
rect -2109 14139 -2079 14157
rect -2041 14139 -2007 14157
rect -1969 14140 -1939 14158
rect -1939 14140 -1935 14158
rect -2113 14123 -2079 14139
rect -2041 14123 -2007 14139
rect -1969 14124 -1935 14140
rect -2113 14070 -2109 14084
rect -2109 14070 -2079 14084
rect -2041 14070 -2007 14084
rect -1969 14071 -1939 14085
rect -1939 14071 -1935 14085
rect -2113 14050 -2079 14070
rect -2041 14050 -2007 14070
rect -1969 14051 -1935 14071
rect -2113 14001 -2109 14011
rect -2109 14001 -2079 14011
rect -2041 14001 -2007 14011
rect -1969 14002 -1939 14012
rect -1939 14002 -1935 14012
rect -2113 13977 -2079 14001
rect -2041 13977 -2007 14001
rect -1969 13978 -1935 14002
rect -2113 13932 -2109 13938
rect -2109 13932 -2079 13938
rect -2041 13932 -2007 13938
rect -1969 13933 -1939 13939
rect -1939 13933 -1935 13939
rect -2113 13904 -2079 13932
rect -2041 13904 -2007 13932
rect -1969 13905 -1935 13933
rect -2113 13863 -2109 13865
rect -2109 13863 -2079 13865
rect -2041 13863 -2007 13865
rect -1969 13864 -1939 13866
rect -1939 13864 -1935 13866
rect -2113 13831 -2079 13863
rect -2041 13831 -2007 13863
rect -1969 13832 -1935 13864
rect -2113 13759 -2079 13792
rect -2041 13759 -2007 13792
rect -1969 13760 -1935 13793
rect -2113 13758 -2109 13759
rect -2109 13758 -2079 13759
rect -2041 13758 -2007 13759
rect -1969 13759 -1939 13760
rect -1939 13759 -1935 13760
rect -2113 13690 -2079 13719
rect -2041 13690 -2007 13719
rect -1969 13691 -1935 13720
rect -2113 13685 -2109 13690
rect -2109 13685 -2079 13690
rect -2041 13685 -2007 13690
rect -1969 13686 -1939 13691
rect -1939 13686 -1935 13691
rect -2113 13621 -2079 13646
rect -2041 13621 -2007 13646
rect -1969 13622 -1935 13647
rect -2113 13612 -2109 13621
rect -2109 13612 -2079 13621
rect -2041 13612 -2007 13621
rect -1969 13613 -1939 13622
rect -1939 13613 -1935 13622
rect -2113 13552 -2079 13573
rect -2041 13552 -2007 13573
rect -1969 13553 -1935 13574
rect -2113 13539 -2109 13552
rect -2109 13539 -2079 13552
rect -2041 13539 -2007 13552
rect -1969 13540 -1939 13553
rect -1939 13540 -1935 13553
rect -2113 13483 -2079 13500
rect -2041 13483 -2007 13500
rect -1969 13484 -1935 13501
rect -2113 13466 -2109 13483
rect -2109 13466 -2079 13483
rect -2041 13466 -2007 13483
rect -1969 13467 -1939 13484
rect -1939 13467 -1935 13484
rect -2113 13414 -2079 13427
rect -2041 13414 -2007 13427
rect -1969 13415 -1935 13428
rect -2113 13393 -2109 13414
rect -2109 13393 -2079 13414
rect -2041 13393 -2007 13414
rect -1969 13394 -1939 13415
rect -1939 13394 -1935 13415
rect -2113 13345 -2079 13354
rect -2041 13345 -2007 13354
rect -1969 13346 -1935 13355
rect -2113 13320 -2109 13345
rect -2109 13320 -2079 13345
rect -2041 13320 -2007 13345
rect -1969 13321 -1939 13346
rect -1939 13321 -1935 13346
rect -2113 13276 -2079 13281
rect -2041 13276 -2007 13281
rect -1969 13277 -1935 13282
rect -2113 13247 -2109 13276
rect -2109 13247 -2079 13276
rect -2041 13247 -2007 13276
rect -1969 13248 -1939 13277
rect -1939 13248 -1935 13277
rect -1969 13208 -1935 13209
rect -2113 13207 -2079 13208
rect -2041 13207 -2007 13208
rect -2113 13174 -2109 13207
rect -2109 13174 -2079 13207
rect -2041 13174 -2007 13207
rect -1969 13175 -1939 13208
rect -1939 13175 -1935 13208
rect -2113 13104 -2109 13135
rect -2109 13104 -2079 13135
rect -2041 13104 -2007 13135
rect -1969 13105 -1939 13136
rect -1939 13105 -1935 13136
rect -2113 13101 -2079 13104
rect -2041 13101 -2007 13104
rect -1969 13102 -1935 13105
rect -2113 13035 -2109 13062
rect -2109 13035 -2079 13062
rect -2041 13035 -2007 13062
rect -1969 13036 -1939 13063
rect -1939 13036 -1935 13063
rect -2113 13028 -2079 13035
rect -2041 13028 -2007 13035
rect -1969 13029 -1935 13036
rect -2113 12966 -2109 12989
rect -2109 12966 -2079 12989
rect -2041 12966 -2007 12989
rect -1969 12967 -1939 12990
rect -1939 12967 -1935 12990
rect -2113 12955 -2079 12966
rect -2041 12955 -2007 12966
rect -1969 12956 -1935 12967
rect -2113 12897 -2109 12916
rect -2109 12897 -2079 12916
rect -2041 12897 -2007 12916
rect -1969 12898 -1939 12917
rect -1939 12898 -1935 12917
rect -2113 12882 -2079 12897
rect -2041 12882 -2007 12897
rect -1969 12883 -1935 12898
rect -2113 12828 -2109 12843
rect -2109 12828 -2079 12843
rect -2041 12828 -2007 12843
rect -1969 12829 -1939 12844
rect -1939 12829 -1935 12844
rect -2113 12809 -2079 12828
rect -2041 12809 -2007 12828
rect -1969 12810 -1935 12829
rect -2113 12759 -2109 12770
rect -2109 12759 -2079 12770
rect -2041 12759 -2007 12770
rect -1969 12760 -1939 12771
rect -1939 12760 -1935 12771
rect -2113 12736 -2079 12759
rect -2041 12736 -2007 12759
rect -1969 12737 -1935 12760
rect -2113 12690 -2109 12697
rect -2109 12690 -2079 12697
rect -2041 12690 -2007 12697
rect -1969 12691 -1939 12698
rect -1939 12691 -1935 12698
rect -2113 12663 -2079 12690
rect -2041 12663 -2007 12690
rect -1969 12664 -1935 12691
rect -2113 12621 -2109 12624
rect -2109 12621 -2079 12624
rect -2041 12621 -2007 12624
rect -1969 12622 -1939 12625
rect -1939 12622 -1935 12625
rect -2113 12590 -2079 12621
rect -2041 12590 -2007 12621
rect -1969 12591 -1935 12622
rect -2113 12517 -2079 12551
rect -2041 12517 -2007 12551
rect -1969 12518 -1935 12552
rect -2113 12448 -2079 12478
rect -2041 12448 -2007 12478
rect -1969 12449 -1935 12479
rect -2113 12444 -2109 12448
rect -2109 12444 -2079 12448
rect -2041 12444 -2007 12448
rect -1969 12445 -1939 12449
rect -1939 12445 -1935 12449
rect -2113 12379 -2079 12405
rect -2041 12379 -2007 12405
rect -1969 12380 -1935 12406
rect -2113 12371 -2109 12379
rect -2109 12371 -2079 12379
rect -2041 12371 -2007 12379
rect -1969 12372 -1939 12380
rect -1939 12372 -1935 12380
rect -2113 12310 -2079 12332
rect -2041 12310 -2007 12332
rect -1969 12311 -1935 12333
rect -2113 12298 -2109 12310
rect -2109 12298 -2079 12310
rect -2041 12298 -2007 12310
rect -1969 12299 -1939 12311
rect -1939 12299 -1935 12311
rect -2113 12241 -2079 12259
rect -2041 12241 -2007 12259
rect -1969 12242 -1935 12260
rect -2113 12225 -2109 12241
rect -2109 12225 -2079 12241
rect -2041 12225 -2007 12241
rect -1969 12226 -1939 12242
rect -1939 12226 -1935 12242
rect -2113 12172 -2007 12186
rect -1969 12173 -1935 12187
rect -2113 12138 -2109 12172
rect -2109 12138 -2075 12172
rect -2075 12138 -2041 12172
rect -2041 12138 -2007 12172
rect -1969 12153 -1939 12173
rect -1939 12153 -1935 12173
rect -2113 12114 -2007 12138
rect -2113 12104 -1935 12114
rect -2113 12103 -1973 12104
rect -2113 12069 -2109 12103
rect -2109 12069 -2075 12103
rect -2075 12069 -2041 12103
rect -2041 12069 -2007 12103
rect -2007 12070 -1973 12103
rect -1973 12070 -1939 12104
rect -1939 12070 -1935 12104
rect -2007 12069 -1935 12070
rect -2113 12035 -1935 12069
rect -2113 12034 -1973 12035
rect -2113 12000 -2109 12034
rect -2109 12000 -2075 12034
rect -2075 12000 -2041 12034
rect -2041 12000 -2007 12034
rect -2007 12001 -1973 12034
rect -1973 12001 -1939 12035
rect -1939 12001 -1935 12035
rect -2007 12000 -1935 12001
rect -2113 11966 -1935 12000
rect -2113 11965 -1973 11966
rect -2113 11931 -2109 11965
rect -2109 11931 -2075 11965
rect -2075 11931 -2041 11965
rect -2041 11931 -2007 11965
rect -2007 11932 -1973 11965
rect -1973 11932 -1939 11966
rect -1939 11932 -1935 11966
rect -2007 11931 -1935 11932
rect -2113 11897 -1935 11931
rect -2113 11896 -1973 11897
rect -2113 11862 -2109 11896
rect -2109 11862 -2075 11896
rect -2075 11862 -2041 11896
rect -2041 11862 -2007 11896
rect -2007 11863 -1973 11896
rect -1973 11863 -1939 11897
rect -1939 11863 -1935 11897
rect -2007 11862 -1935 11863
rect -2113 11828 -1935 11862
rect -2113 11827 -1973 11828
rect -2113 11793 -2109 11827
rect -2109 11793 -2075 11827
rect -2075 11793 -2041 11827
rect -2041 11793 -2007 11827
rect -2007 11794 -1973 11827
rect -1973 11794 -1939 11828
rect -1939 11794 -1935 11828
rect -2007 11793 -1935 11794
rect -2113 11759 -1935 11793
rect -2113 11758 -1973 11759
rect -2113 11724 -2109 11758
rect -2109 11724 -2075 11758
rect -2075 11724 -2041 11758
rect -2041 11724 -2007 11758
rect -2007 11725 -1973 11758
rect -1973 11725 -1939 11759
rect -1939 11725 -1935 11759
rect -2007 11724 -1935 11725
rect -2113 11690 -1935 11724
rect -2113 11689 -1973 11690
rect -2113 11655 -2109 11689
rect -2109 11655 -2075 11689
rect -2075 11655 -2041 11689
rect -2041 11655 -2007 11689
rect -2007 11656 -1973 11689
rect -1973 11656 -1939 11690
rect -1939 11656 -1935 11690
rect -2007 11655 -1935 11656
rect -2113 11621 -1935 11655
rect -2113 11620 -1973 11621
rect -2113 11586 -2109 11620
rect -2109 11586 -2075 11620
rect -2075 11586 -2041 11620
rect -2041 11586 -2007 11620
rect -2007 11587 -1973 11620
rect -1973 11587 -1939 11621
rect -1939 11587 -1935 11621
rect -2007 11586 -1935 11587
rect -2113 11552 -1935 11586
rect -2113 11551 -1973 11552
rect -2113 11517 -2109 11551
rect -2109 11517 -2075 11551
rect -2075 11517 -2041 11551
rect -2041 11517 -2007 11551
rect -2007 11518 -1973 11551
rect -1973 11518 -1939 11552
rect -1939 11518 -1935 11552
rect -2007 11517 -1935 11518
rect -2113 11483 -1935 11517
rect -2113 11482 -1973 11483
rect -2113 11448 -2109 11482
rect -2109 11448 -2075 11482
rect -2075 11448 -2041 11482
rect -2041 11448 -2007 11482
rect -2007 11449 -1973 11482
rect -1973 11449 -1939 11483
rect -1939 11449 -1935 11483
rect -2007 11448 -1935 11449
rect -2113 11414 -1935 11448
rect -2113 11413 -1973 11414
rect -2113 11379 -2109 11413
rect -2109 11379 -2075 11413
rect -2075 11379 -2041 11413
rect -2041 11379 -2007 11413
rect -2007 11380 -1973 11413
rect -1973 11380 -1939 11414
rect -1939 11380 -1935 11414
rect -2007 11379 -1935 11380
rect -2113 11345 -1935 11379
rect -2113 11344 -1973 11345
rect -2113 11310 -2109 11344
rect -2109 11310 -2075 11344
rect -2075 11310 -2041 11344
rect -2041 11310 -2007 11344
rect -2007 11311 -1973 11344
rect -1973 11311 -1939 11345
rect -1939 11311 -1935 11345
rect -2007 11310 -1935 11311
rect -2113 11276 -1935 11310
rect -2113 11275 -1973 11276
rect -2113 11241 -2109 11275
rect -2109 11241 -2075 11275
rect -2075 11241 -2041 11275
rect -2041 11241 -2007 11275
rect -2007 11242 -1973 11275
rect -1973 11242 -1939 11276
rect -1939 11242 -1935 11276
rect -2007 11241 -1935 11242
rect -2113 11207 -1935 11241
rect -2113 11206 -1973 11207
rect -2113 11172 -2109 11206
rect -2109 11172 -2075 11206
rect -2075 11172 -2041 11206
rect -2041 11172 -2007 11206
rect -2007 11173 -1973 11206
rect -1973 11173 -1939 11207
rect -1939 11173 -1935 11207
rect -2007 11172 -1935 11173
rect -2113 11138 -1935 11172
rect -2113 11137 -1973 11138
rect -2113 11103 -2109 11137
rect -2109 11103 -2075 11137
rect -2075 11103 -2041 11137
rect -2041 11103 -2007 11137
rect -2007 11104 -1973 11137
rect -1973 11104 -1939 11138
rect -1939 11104 -1935 11138
rect -2007 11103 -1935 11104
rect -2113 11069 -1935 11103
rect -2113 11068 -1973 11069
rect -2113 11034 -2109 11068
rect -2109 11034 -2075 11068
rect -2075 11034 -2041 11068
rect -2041 11034 -2007 11068
rect -2007 11035 -1973 11068
rect -1973 11035 -1939 11069
rect -1939 11035 -1935 11069
rect -2007 11034 -1935 11035
rect -2113 11000 -1935 11034
rect -2113 10999 -1973 11000
rect -2113 10965 -2109 10999
rect -2109 10965 -2075 10999
rect -2075 10965 -2041 10999
rect -2041 10965 -2007 10999
rect -2007 10966 -1973 10999
rect -1973 10966 -1939 11000
rect -1939 10966 -1935 11000
rect -2007 10965 -1935 10966
rect -2113 10931 -1935 10965
rect -2113 10930 -1973 10931
rect -2113 10896 -2109 10930
rect -2109 10896 -2075 10930
rect -2075 10896 -2041 10930
rect -2041 10896 -2007 10930
rect -2007 10897 -1973 10930
rect -1973 10897 -1939 10931
rect -1939 10897 -1935 10931
rect -2007 10896 -1935 10897
rect -2113 10862 -1935 10896
rect -2113 10861 -1973 10862
rect -2113 10827 -2109 10861
rect -2109 10827 -2075 10861
rect -2075 10827 -2041 10861
rect -2041 10827 -2007 10861
rect -2007 10828 -1973 10861
rect -1973 10828 -1939 10862
rect -1939 10828 -1935 10862
rect -2007 10827 -1935 10828
rect -2113 10793 -1935 10827
rect -2113 10792 -1973 10793
rect -2113 10758 -2109 10792
rect -2109 10758 -2075 10792
rect -2075 10758 -2041 10792
rect -2041 10758 -2007 10792
rect -2007 10759 -1973 10792
rect -1973 10759 -1939 10793
rect -1939 10759 -1935 10793
rect -2007 10758 -1935 10759
rect -2113 10724 -1935 10758
rect -2113 10723 -1973 10724
rect -2113 10689 -2109 10723
rect -2109 10689 -2075 10723
rect -2075 10689 -2041 10723
rect -2041 10689 -2007 10723
rect -2007 10690 -1973 10723
rect -1973 10690 -1939 10724
rect -1939 10690 -1935 10724
rect -2007 10689 -1935 10690
rect -2113 10655 -1935 10689
rect -2113 10654 -1973 10655
rect -2113 10620 -2109 10654
rect -2109 10620 -2075 10654
rect -2075 10620 -2041 10654
rect -2041 10620 -2007 10654
rect -2007 10621 -1973 10654
rect -1973 10621 -1939 10655
rect -1939 10621 -1935 10655
rect -2007 10620 -1935 10621
rect -2113 10586 -1935 10620
rect -2113 10585 -1973 10586
rect -2113 10551 -2109 10585
rect -2109 10551 -2075 10585
rect -2075 10551 -2041 10585
rect -2041 10551 -2007 10585
rect -2007 10552 -1973 10585
rect -1973 10552 -1939 10586
rect -1939 10552 -1935 10586
rect -2007 10551 -1935 10552
rect -2113 10517 -1935 10551
rect -2113 10516 -1973 10517
rect -2113 10482 -2109 10516
rect -2109 10482 -2075 10516
rect -2075 10482 -2041 10516
rect -2041 10482 -2007 10516
rect -2007 10483 -1973 10516
rect -1973 10483 -1939 10517
rect -1939 10483 -1935 10517
rect -2007 10482 -1935 10483
rect -2113 10448 -1935 10482
rect -2113 10447 -1973 10448
rect -2113 10413 -2109 10447
rect -2109 10413 -2075 10447
rect -2075 10413 -2041 10447
rect -2041 10413 -2007 10447
rect -2007 10414 -1973 10447
rect -1973 10414 -1939 10448
rect -1939 10414 -1935 10448
rect -2007 10413 -1935 10414
rect -2113 10379 -1935 10413
rect -2113 10378 -1973 10379
rect -2113 10344 -2109 10378
rect -2109 10344 -2075 10378
rect -2075 10344 -2041 10378
rect -2041 10344 -2007 10378
rect -2007 10345 -1973 10378
rect -1973 10345 -1939 10379
rect -1939 10345 -1935 10379
rect -2007 10344 -1935 10345
rect -2113 10310 -1935 10344
rect -2113 10309 -1973 10310
rect -2113 10275 -2109 10309
rect -2109 10275 -2075 10309
rect -2075 10275 -2041 10309
rect -2041 10275 -2007 10309
rect -2007 10276 -1973 10309
rect -1973 10276 -1939 10310
rect -1939 10276 -1935 10310
rect -2007 10275 -1935 10276
rect -2113 10241 -1935 10275
rect -2113 10240 -1973 10241
rect -2113 10206 -2109 10240
rect -2109 10206 -2075 10240
rect -2075 10206 -2041 10240
rect -2041 10206 -2007 10240
rect -2007 10207 -1973 10240
rect -1973 10207 -1939 10241
rect -1939 10207 -1935 10241
rect -2007 10206 -1935 10207
rect -2113 10172 -1935 10206
rect -2113 10171 -1973 10172
rect -2113 10137 -2109 10171
rect -2109 10137 -2075 10171
rect -2075 10137 -2041 10171
rect -2041 10137 -2007 10171
rect -2007 10138 -1973 10171
rect -1973 10138 -1939 10172
rect -1939 10138 -1935 10172
rect -2007 10137 -1935 10138
rect -2113 10103 -1935 10137
rect -2113 10102 -1973 10103
rect -2113 10068 -2109 10102
rect -2109 10068 -2075 10102
rect -2075 10068 -2041 10102
rect -2041 10068 -2007 10102
rect -2007 10069 -1973 10102
rect -1973 10069 -1939 10103
rect -1939 10069 -1935 10103
rect -2007 10068 -1935 10069
rect -2113 10034 -1935 10068
rect -2113 10033 -1973 10034
rect -2113 9999 -2109 10033
rect -2109 9999 -2075 10033
rect -2075 9999 -2041 10033
rect -2041 9999 -2007 10033
rect -2007 10000 -1973 10033
rect -1973 10000 -1939 10034
rect -1939 10000 -1935 10034
rect -2007 9999 -1935 10000
rect -2113 9965 -1935 9999
rect -2113 9964 -1973 9965
rect -2113 9930 -2109 9964
rect -2109 9930 -2075 9964
rect -2075 9930 -2041 9964
rect -2041 9930 -2007 9964
rect -2007 9931 -1973 9964
rect -1973 9931 -1939 9965
rect -1939 9931 -1935 9965
rect -2007 9930 -1935 9931
rect -2113 9896 -1935 9930
rect -2113 9895 -1973 9896
rect -2113 7617 -2109 9895
rect -2109 9827 -2007 9895
rect -2007 9862 -1973 9895
rect -1973 9862 -1939 9896
rect -1939 9862 -1935 9896
rect -2007 9827 -1935 9862
rect -2109 7688 -1939 9827
rect -1939 7688 -1935 9827
rect -1711 14195 -1677 14197
rect -1711 14163 -1677 14195
rect -1633 14163 -1599 14197
rect -1555 14195 -1521 14197
rect -1477 14195 -1443 14197
rect -1399 14195 -1365 14197
rect -1321 14195 -1287 14197
rect -1243 14195 -1209 14197
rect -1165 14195 -1131 14197
rect -1555 14163 -1521 14195
rect -1477 14163 -1443 14195
rect -1399 14163 -1365 14195
rect -1321 14163 -1287 14195
rect -1243 14163 -1209 14195
rect -1165 14163 -1131 14195
rect -1789 14091 -1787 14125
rect -1787 14091 -1755 14125
rect -1717 14091 -1685 14125
rect -1685 14091 -1683 14125
rect -1633 14091 -1599 14125
rect -1555 14093 -1521 14125
rect -1477 14093 -1443 14125
rect -1399 14093 -1365 14125
rect -1321 14093 -1287 14125
rect -1243 14093 -1209 14125
rect -1165 14093 -1129 14125
rect -1129 14114 -1059 14125
rect -1129 14093 -1095 14114
rect -1555 14091 -1521 14093
rect -1477 14091 -1443 14093
rect -1399 14091 -1365 14093
rect -1321 14091 -1287 14093
rect -1243 14091 -1209 14093
rect -1789 14018 -1787 14052
rect -1787 14018 -1755 14052
rect -1717 14018 -1685 14052
rect -1685 14018 -1683 14052
rect -1789 13945 -1787 13979
rect -1787 13945 -1755 13979
rect -1717 13945 -1685 13979
rect -1685 13945 -1683 13979
rect -1789 13872 -1787 13906
rect -1787 13872 -1755 13906
rect -1717 13872 -1685 13906
rect -1685 13872 -1683 13906
rect -1789 13799 -1787 13833
rect -1787 13799 -1755 13833
rect -1717 13799 -1685 13833
rect -1685 13799 -1683 13833
rect -1789 13726 -1787 13760
rect -1787 13726 -1755 13760
rect -1717 13726 -1685 13760
rect -1685 13726 -1683 13760
rect -1789 13653 -1787 13687
rect -1787 13653 -1755 13687
rect -1717 13653 -1685 13687
rect -1685 13653 -1683 13687
rect -1789 13580 -1787 13614
rect -1787 13580 -1755 13614
rect -1717 13580 -1685 13614
rect -1685 13580 -1683 13614
rect -1789 13507 -1787 13541
rect -1787 13507 -1755 13541
rect -1717 13507 -1685 13541
rect -1685 13507 -1683 13541
rect -1789 8041 -1787 13468
rect -1787 8041 -1685 13468
rect -1685 8041 -1683 13468
rect -1789 8007 -1683 8041
rect -1789 7973 -1787 8007
rect -1787 7973 -1753 8007
rect -1753 7994 -1683 8007
rect -1165 14080 -1095 14093
rect -1095 14080 -1061 14114
rect -1061 14080 -1059 14114
rect -1165 14046 -1059 14080
rect -1165 14019 -1163 14046
rect -1163 14019 -1061 14046
rect -1061 14019 -1059 14046
rect -1165 13946 -1163 13980
rect -1163 13946 -1131 13980
rect -1093 13946 -1061 13980
rect -1061 13946 -1059 13980
rect -1165 13873 -1163 13907
rect -1163 13873 -1131 13907
rect -1093 13873 -1061 13907
rect -1061 13873 -1059 13907
rect -1165 13800 -1163 13834
rect -1163 13800 -1131 13834
rect -1093 13800 -1061 13834
rect -1061 13800 -1059 13834
rect -1165 13727 -1163 13761
rect -1163 13727 -1131 13761
rect -1093 13727 -1061 13761
rect -1061 13727 -1059 13761
rect -1165 13654 -1163 13688
rect -1163 13654 -1131 13688
rect -1093 13654 -1061 13688
rect -1061 13654 -1059 13688
rect -1165 13581 -1163 13615
rect -1163 13581 -1131 13615
rect -1093 13581 -1061 13615
rect -1061 13581 -1059 13615
rect -1165 13508 -1163 13542
rect -1163 13508 -1131 13542
rect -1093 13508 -1061 13542
rect -1061 13508 -1059 13542
rect -1165 13435 -1163 13469
rect -1163 13435 -1131 13469
rect -1093 13435 -1061 13469
rect -1061 13435 -1059 13469
rect -1165 13362 -1163 13396
rect -1163 13362 -1131 13396
rect -1093 13362 -1061 13396
rect -1061 13362 -1059 13396
rect -1165 13289 -1163 13323
rect -1163 13289 -1131 13323
rect -1093 13289 -1061 13323
rect -1061 13289 -1059 13323
rect -1165 13216 -1163 13250
rect -1163 13216 -1131 13250
rect -1093 13216 -1061 13250
rect -1061 13216 -1059 13250
rect -1165 13143 -1163 13177
rect -1163 13143 -1131 13177
rect -1093 13143 -1061 13177
rect -1061 13143 -1059 13177
rect -1165 13070 -1163 13104
rect -1163 13070 -1131 13104
rect -1093 13070 -1061 13104
rect -1061 13070 -1059 13104
rect -1165 12997 -1163 13031
rect -1163 12997 -1131 13031
rect -1093 12997 -1061 13031
rect -1061 12997 -1059 13031
rect -1165 12924 -1163 12958
rect -1163 12924 -1131 12958
rect -1093 12924 -1061 12958
rect -1061 12924 -1059 12958
rect -1165 12851 -1163 12885
rect -1163 12851 -1131 12885
rect -1093 12851 -1061 12885
rect -1061 12851 -1059 12885
rect -1165 12778 -1163 12812
rect -1163 12778 -1131 12812
rect -1093 12778 -1061 12812
rect -1061 12778 -1059 12812
rect -1165 12705 -1163 12739
rect -1163 12705 -1131 12739
rect -1093 12705 -1061 12739
rect -1061 12705 -1059 12739
rect -1165 12632 -1163 12666
rect -1163 12632 -1131 12666
rect -1093 12632 -1061 12666
rect -1061 12632 -1059 12666
rect -1165 12534 -1163 12568
rect -1163 12534 -1131 12568
rect -1093 12534 -1061 12568
rect -1061 12534 -1059 12568
rect -1519 12472 -1485 12506
rect -1363 12472 -1329 12506
rect -1519 12400 -1485 12434
rect -1363 12400 -1329 12434
rect -1165 12461 -1163 12495
rect -1163 12461 -1131 12495
rect -1093 12461 -1061 12495
rect -1061 12461 -1059 12495
rect -1165 12388 -1163 12422
rect -1163 12388 -1131 12422
rect -1093 12388 -1061 12422
rect -1061 12388 -1059 12422
rect -1597 12309 -1563 12321
rect -1597 12287 -1563 12309
rect -1597 12241 -1563 12249
rect -1597 12215 -1563 12241
rect -1597 12173 -1563 12177
rect -1597 12143 -1563 12173
rect -1597 12071 -1563 12105
rect -1597 12003 -1563 12033
rect -1597 11999 -1563 12003
rect -1597 11935 -1563 11961
rect -1597 11927 -1563 11935
rect -1597 11867 -1563 11889
rect -1597 11855 -1563 11867
rect -1597 11799 -1563 11817
rect -1597 11783 -1563 11799
rect -1441 12309 -1407 12321
rect -1441 12287 -1407 12309
rect -1441 12241 -1407 12249
rect -1441 12215 -1407 12241
rect -1441 12173 -1407 12177
rect -1441 12143 -1407 12173
rect -1441 12071 -1407 12105
rect -1441 12003 -1407 12033
rect -1441 11999 -1407 12003
rect -1441 11935 -1407 11961
rect -1441 11927 -1407 11935
rect -1441 11867 -1407 11889
rect -1441 11855 -1407 11867
rect -1441 11799 -1407 11817
rect -1441 11783 -1407 11799
rect -1285 12309 -1251 12321
rect -1285 12287 -1251 12309
rect -1285 12241 -1251 12249
rect -1285 12215 -1251 12241
rect -1285 12173 -1251 12177
rect -1285 12143 -1251 12173
rect -1285 12071 -1251 12105
rect -1285 12003 -1251 12033
rect -1285 11999 -1251 12003
rect -1285 11935 -1251 11961
rect -1285 11927 -1251 11935
rect -1285 11867 -1251 11889
rect -1285 11855 -1251 11867
rect -1285 11799 -1251 11817
rect -1285 11783 -1251 11799
rect -1165 12315 -1163 12349
rect -1163 12315 -1131 12349
rect -1093 12315 -1061 12349
rect -1061 12315 -1059 12349
rect -1165 12242 -1163 12276
rect -1163 12242 -1131 12276
rect -1093 12242 -1061 12276
rect -1061 12242 -1059 12276
rect -1165 12169 -1163 12203
rect -1163 12169 -1131 12203
rect -1093 12169 -1061 12203
rect -1061 12169 -1059 12203
rect -1165 12096 -1163 12130
rect -1163 12096 -1131 12130
rect -1093 12096 -1061 12130
rect -1061 12096 -1059 12130
rect -1165 12023 -1163 12057
rect -1163 12023 -1131 12057
rect -1093 12023 -1061 12057
rect -1061 12023 -1059 12057
rect -1165 11950 -1163 11984
rect -1163 11950 -1131 11984
rect -1093 11950 -1061 11984
rect -1061 11950 -1059 11984
rect -1165 11877 -1163 11911
rect -1163 11877 -1131 11911
rect -1093 11877 -1061 11911
rect -1061 11877 -1059 11911
rect -1165 11804 -1163 11838
rect -1163 11804 -1131 11838
rect -1093 11804 -1061 11838
rect -1061 11804 -1059 11838
rect -1519 11740 -1485 11774
rect -1363 11740 -1329 11774
rect -1519 11668 -1485 11702
rect -1363 11668 -1329 11702
rect -1165 11731 -1163 11765
rect -1163 11731 -1131 11765
rect -1093 11731 -1061 11765
rect -1061 11731 -1059 11765
rect -1597 11643 -1563 11659
rect -1597 11625 -1563 11643
rect -1597 11575 -1563 11587
rect -1597 11553 -1563 11575
rect -1597 11507 -1563 11515
rect -1597 11481 -1563 11507
rect -1597 11439 -1563 11443
rect -1597 11409 -1563 11439
rect -1597 11337 -1563 11371
rect -1597 11269 -1563 11299
rect -1597 11265 -1563 11269
rect -1597 11201 -1563 11227
rect -1597 11193 -1563 11201
rect -1597 11133 -1563 11155
rect -1597 11121 -1563 11133
rect -1441 11643 -1407 11659
rect -1441 11625 -1407 11643
rect -1441 11575 -1407 11587
rect -1441 11553 -1407 11575
rect -1441 11507 -1407 11515
rect -1441 11481 -1407 11507
rect -1441 11439 -1407 11443
rect -1441 11409 -1407 11439
rect -1441 11337 -1407 11371
rect -1441 11269 -1407 11299
rect -1441 11265 -1407 11269
rect -1441 11201 -1407 11227
rect -1441 11193 -1407 11201
rect -1441 11133 -1407 11155
rect -1441 11121 -1407 11133
rect -1285 11643 -1251 11659
rect -1285 11625 -1251 11643
rect -1285 11575 -1251 11587
rect -1285 11553 -1251 11575
rect -1285 11507 -1251 11515
rect -1285 11481 -1251 11507
rect -1285 11439 -1251 11443
rect -1285 11409 -1251 11439
rect -1285 11337 -1251 11371
rect -1285 11269 -1251 11299
rect -1285 11265 -1251 11269
rect -1285 11201 -1251 11227
rect -1285 11193 -1251 11201
rect -1285 11133 -1251 11155
rect -1285 11121 -1251 11133
rect -1165 11658 -1163 11692
rect -1163 11658 -1131 11692
rect -1093 11658 -1061 11692
rect -1061 11658 -1059 11692
rect -1165 11585 -1163 11619
rect -1163 11585 -1131 11619
rect -1093 11585 -1061 11619
rect -1061 11585 -1059 11619
rect -1165 11512 -1163 11546
rect -1163 11512 -1131 11546
rect -1093 11512 -1061 11546
rect -1061 11512 -1059 11546
rect -1165 11439 -1163 11473
rect -1163 11439 -1131 11473
rect -1093 11439 -1061 11473
rect -1061 11439 -1059 11473
rect -1165 11366 -1163 11400
rect -1163 11366 -1131 11400
rect -1093 11366 -1061 11400
rect -1061 11366 -1059 11400
rect -1165 11293 -1163 11327
rect -1163 11293 -1131 11327
rect -1093 11293 -1061 11327
rect -1061 11293 -1059 11327
rect -1165 11220 -1163 11254
rect -1163 11220 -1131 11254
rect -1093 11220 -1061 11254
rect -1061 11220 -1059 11254
rect -1165 11147 -1163 11181
rect -1163 11147 -1131 11181
rect -1093 11147 -1061 11181
rect -1061 11147 -1059 11181
rect -1165 11074 -1163 11108
rect -1163 11074 -1131 11108
rect -1093 11074 -1061 11108
rect -1061 11074 -1059 11108
rect -1519 11008 -1485 11042
rect -1363 11008 -1329 11042
rect -1519 10936 -1485 10970
rect -1363 10936 -1329 10970
rect -1165 11001 -1163 11035
rect -1163 11001 -1131 11035
rect -1093 11001 -1061 11035
rect -1061 11001 -1059 11035
rect -1165 10928 -1163 10962
rect -1163 10928 -1131 10962
rect -1093 10928 -1061 10962
rect -1061 10928 -1059 10962
rect -1597 10845 -1563 10857
rect -1597 10823 -1563 10845
rect -1597 10777 -1563 10785
rect -1597 10751 -1563 10777
rect -1597 10709 -1563 10713
rect -1597 10679 -1563 10709
rect -1597 10607 -1563 10641
rect -1597 10539 -1563 10569
rect -1597 10535 -1563 10539
rect -1597 10471 -1563 10497
rect -1597 10463 -1563 10471
rect -1597 10403 -1563 10425
rect -1597 10391 -1563 10403
rect -1597 10335 -1563 10353
rect -1597 10319 -1563 10335
rect -1441 10845 -1407 10857
rect -1441 10823 -1407 10845
rect -1441 10777 -1407 10785
rect -1441 10751 -1407 10777
rect -1441 10709 -1407 10713
rect -1441 10679 -1407 10709
rect -1441 10607 -1407 10641
rect -1441 10539 -1407 10569
rect -1441 10535 -1407 10539
rect -1441 10471 -1407 10497
rect -1441 10463 -1407 10471
rect -1441 10403 -1407 10425
rect -1441 10391 -1407 10403
rect -1441 10335 -1407 10353
rect -1441 10319 -1407 10335
rect -1285 10845 -1251 10857
rect -1285 10823 -1251 10845
rect -1285 10777 -1251 10785
rect -1285 10751 -1251 10777
rect -1285 10709 -1251 10713
rect -1285 10679 -1251 10709
rect -1285 10607 -1251 10641
rect -1285 10539 -1251 10569
rect -1285 10535 -1251 10539
rect -1285 10471 -1251 10497
rect -1285 10463 -1251 10471
rect -1285 10403 -1251 10425
rect -1285 10391 -1251 10403
rect -1285 10335 -1251 10353
rect -1285 10319 -1251 10335
rect -1165 10855 -1163 10889
rect -1163 10855 -1131 10889
rect -1093 10855 -1061 10889
rect -1061 10855 -1059 10889
rect -1165 10782 -1163 10816
rect -1163 10782 -1131 10816
rect -1093 10782 -1061 10816
rect -1061 10782 -1059 10816
rect -1165 10709 -1163 10743
rect -1163 10709 -1131 10743
rect -1093 10709 -1061 10743
rect -1061 10709 -1059 10743
rect -1165 10636 -1163 10670
rect -1163 10636 -1131 10670
rect -1093 10636 -1061 10670
rect -1061 10636 -1059 10670
rect -1165 10563 -1163 10597
rect -1163 10563 -1131 10597
rect -1093 10563 -1061 10597
rect -1061 10563 -1059 10597
rect -1165 10490 -1163 10524
rect -1163 10490 -1131 10524
rect -1093 10490 -1061 10524
rect -1061 10490 -1059 10524
rect -1165 10417 -1163 10451
rect -1163 10417 -1131 10451
rect -1093 10417 -1061 10451
rect -1061 10417 -1059 10451
rect -1165 10344 -1163 10378
rect -1163 10344 -1131 10378
rect -1093 10344 -1061 10378
rect -1061 10344 -1059 10378
rect -1165 10271 -1163 10305
rect -1163 10271 -1131 10305
rect -1093 10271 -1061 10305
rect -1061 10271 -1059 10305
rect -1165 10198 -1163 10232
rect -1163 10198 -1131 10232
rect -1093 10198 -1061 10232
rect -1061 10198 -1059 10232
rect -1165 10125 -1163 10159
rect -1163 10125 -1131 10159
rect -1093 10125 -1061 10159
rect -1061 10125 -1059 10159
rect -1165 10052 -1163 10086
rect -1163 10052 -1131 10086
rect -1093 10052 -1061 10086
rect -1061 10052 -1059 10086
rect -1165 8035 -1163 10013
rect -1163 8035 -1061 10013
rect -1061 8035 -1059 10013
rect -1641 7994 -1607 7996
rect -1565 7994 -1531 7996
rect -1490 7994 -1456 7996
rect -1415 7994 -1381 7996
rect -1340 7994 -1306 7996
rect -1265 7994 -1231 7996
rect -1753 7973 -1719 7994
rect -1789 7962 -1719 7973
rect -1719 7962 -1683 7994
rect -1641 7962 -1607 7994
rect -1565 7962 -1531 7994
rect -1490 7962 -1456 7994
rect -1415 7962 -1381 7994
rect -1340 7962 -1306 7994
rect -1265 7962 -1231 7994
rect -1190 7962 -1163 7996
rect -1163 7962 -1156 7996
rect -1717 7892 -1683 7924
rect -1639 7892 -1605 7924
rect -1561 7892 -1527 7924
rect -1483 7892 -1449 7924
rect -1405 7892 -1371 7924
rect -1327 7892 -1293 7924
rect -1249 7892 -1215 7924
rect -1171 7892 -1141 7924
rect -1141 7892 -1137 7924
rect -1093 7913 -1059 7947
rect -1717 7890 -1683 7892
rect -1639 7890 -1605 7892
rect -1561 7890 -1527 7892
rect -1483 7890 -1449 7892
rect -1405 7890 -1371 7892
rect -1327 7890 -1293 7892
rect -1249 7890 -1215 7892
rect -1171 7890 -1137 7892
rect -1895 7719 -1861 7722
rect -1821 7719 -1787 7722
rect -1747 7719 -1713 7722
rect -1673 7719 -1639 7722
rect -1599 7719 -1565 7722
rect -1895 7688 -1870 7719
rect -1870 7688 -1861 7719
rect -1821 7688 -1801 7719
rect -1801 7688 -1787 7719
rect -1747 7688 -1732 7719
rect -1732 7688 -1713 7719
rect -1673 7688 -1663 7719
rect -1663 7688 -1639 7719
rect -1599 7688 -1594 7719
rect -1594 7688 -1565 7719
rect -2109 7617 -2007 7688
rect -1525 7688 -1491 7722
rect -1451 7719 -1417 7722
rect -1377 7719 -1343 7722
rect -1303 7719 -1269 7722
rect -1229 7719 -1195 7722
rect -1155 7719 -1121 7722
rect -1081 7719 -1047 7722
rect -1007 7719 -973 7722
rect -933 7719 -899 7722
rect -859 7719 -825 7722
rect -786 7719 -752 7722
rect -713 7719 -679 7722
rect -1451 7688 -1421 7719
rect -1421 7688 -1417 7719
rect -1377 7688 -1352 7719
rect -1352 7688 -1343 7719
rect -1303 7688 -1283 7719
rect -1283 7688 -1269 7719
rect -1229 7688 -1214 7719
rect -1214 7688 -1195 7719
rect -1155 7688 -1145 7719
rect -1145 7688 -1121 7719
rect -1081 7688 -1076 7719
rect -1076 7688 -1047 7719
rect -1007 7688 -973 7719
rect -933 7688 -899 7719
rect -859 7688 -825 7719
rect -786 7688 -752 7719
rect -713 7688 -702 7719
rect -702 7688 -679 7719
rect -1967 7617 -1938 7650
rect -1938 7617 -1933 7650
rect -1893 7617 -1869 7650
rect -1869 7617 -1859 7650
rect -1819 7617 -1800 7650
rect -1800 7617 -1785 7650
rect -1745 7617 -1731 7650
rect -1731 7617 -1711 7650
rect -1671 7617 -1662 7650
rect -1662 7617 -1637 7650
rect -1597 7617 -1593 7650
rect -1593 7617 -1563 7650
rect -2113 7616 -2007 7617
rect -1967 7616 -1933 7617
rect -1893 7616 -1859 7617
rect -1819 7616 -1785 7617
rect -1745 7616 -1711 7617
rect -1671 7616 -1637 7617
rect -1597 7616 -1563 7617
rect -1523 7616 -1489 7650
rect -1449 7617 -1420 7650
rect -1420 7617 -1415 7650
rect -1375 7617 -1351 7650
rect -1351 7617 -1341 7650
rect -1301 7617 -1282 7650
rect -1282 7617 -1267 7650
rect -1227 7617 -1213 7650
rect -1213 7617 -1193 7650
rect -1449 7616 -1415 7617
rect -1375 7616 -1341 7617
rect -1301 7616 -1267 7617
rect -1227 7616 -1193 7617
rect -1153 7616 -1144 7650
rect -1144 7616 -1119 7650
rect -1079 7616 -1045 7650
rect -1005 7616 -971 7650
rect -932 7616 -898 7650
rect -859 7616 -825 7650
rect -786 7616 -752 7650
rect -713 7616 -702 7650
rect -702 7616 -679 7650
rect -2041 7549 -2007 7578
rect -1967 7549 -1938 7578
rect -1938 7549 -1933 7578
rect -1893 7549 -1869 7578
rect -1869 7549 -1859 7578
rect -1819 7549 -1800 7578
rect -1800 7549 -1785 7578
rect -1745 7549 -1731 7578
rect -1731 7549 -1711 7578
rect -1671 7549 -1662 7578
rect -1662 7549 -1637 7578
rect -1597 7549 -1593 7578
rect -1593 7549 -1563 7578
rect -2041 7544 -2007 7549
rect -1967 7544 -1933 7549
rect -1893 7544 -1859 7549
rect -1819 7544 -1785 7549
rect -1745 7544 -1711 7549
rect -1671 7544 -1637 7549
rect -1597 7544 -1563 7549
rect -1523 7544 -1489 7578
rect -1449 7549 -1420 7578
rect -1420 7549 -1415 7578
rect -1375 7549 -1351 7578
rect -1351 7549 -1341 7578
rect -1301 7549 -1282 7578
rect -1282 7549 -1267 7578
rect -1227 7549 -1213 7578
rect -1213 7549 -1193 7578
rect -1153 7549 -1144 7578
rect -1144 7549 -1119 7578
rect -1079 7549 -1045 7578
rect -1005 7549 -971 7578
rect -932 7549 -898 7578
rect -859 7549 -825 7578
rect -786 7549 -752 7578
rect -713 7549 -702 7578
rect -702 7549 -679 7578
rect -1449 7544 -1415 7549
rect -1375 7544 -1341 7549
rect -1301 7544 -1267 7549
rect -1227 7544 -1193 7549
rect -1153 7544 -1119 7549
rect -1079 7544 -1045 7549
rect -1005 7544 -971 7549
rect -932 7544 -898 7549
rect -859 7544 -825 7549
rect -786 7544 -752 7549
rect -713 7544 -679 7549
rect 21789 6118 21895 6165
rect 19693 6084 19722 6117
rect 19722 6084 19727 6117
rect 19693 6083 19727 6084
rect 19765 6083 19799 6117
rect 21789 6084 21796 6118
rect 21796 6084 21830 6118
rect 21830 6084 21864 6118
rect 21864 6084 21895 6118
rect 21789 6059 21895 6084
rect 19693 5457 19697 5490
rect 19697 5457 19727 5490
rect 19765 5457 19799 5490
rect 19693 5456 19727 5457
rect 19765 5456 19799 5457
rect 21772 5491 21878 5526
rect 21772 5457 21839 5491
rect 21839 5457 21873 5491
rect 21873 5457 21878 5491
rect 21772 5420 21878 5457
rect -20 2894 14 2928
rect 53 2894 87 2928
rect 126 2894 160 2928
rect 199 2894 233 2928
rect 272 2894 306 2928
rect 345 2894 379 2928
rect 418 2894 452 2928
rect 491 2894 525 2928
rect 564 2894 598 2928
rect 637 2894 671 2928
rect 710 2894 744 2928
rect 783 2894 817 2928
rect 856 2894 890 2928
rect 929 2894 963 2928
rect 1002 2894 1036 2928
rect 1075 2894 1109 2928
rect 1148 2894 1182 2928
rect 1221 2894 1255 2928
rect 1294 2894 1328 2928
rect 1367 2894 1401 2928
rect 1440 2894 1474 2928
rect 1513 2894 1547 2928
rect 1586 2894 1620 2928
rect 1659 2894 1693 2928
rect 1732 2894 1766 2928
rect 1805 2894 1839 2928
rect 1878 2894 1912 2928
rect 1951 2894 1985 2928
rect 2024 2894 2058 2928
rect 2097 2894 2131 2928
rect 2170 2894 2204 2928
rect 2243 2894 2277 2928
rect 2316 2894 2350 2928
rect 2389 2894 2423 2928
rect 2462 2894 2496 2928
rect 2535 2894 2569 2928
rect 2608 2894 2642 2928
rect 2681 2894 2715 2928
rect 2754 2894 2788 2928
rect 2827 2894 2861 2928
rect 2900 2894 2934 2928
rect 2973 2894 3007 2928
rect 3046 2894 3080 2928
rect 3119 2894 3153 2928
rect 3192 2894 3226 2928
rect 3265 2894 3299 2928
rect 3338 2894 3372 2928
rect 3411 2894 3445 2928
rect 3483 2894 3517 2928
rect 3555 2894 3589 2928
rect 3627 2894 3661 2928
rect 3699 2894 3733 2928
rect 3771 2894 3805 2928
rect 3843 2894 3877 2928
rect 3915 2894 3949 2928
rect 3987 2894 4021 2928
rect 4059 2894 4093 2928
rect 4131 2894 4165 2928
rect 4203 2894 4237 2928
rect 4275 2894 4309 2928
rect 4347 2894 4381 2928
rect 4419 2894 4453 2928
rect 4491 2894 4525 2928
rect 4563 2894 4597 2928
rect 4635 2894 4669 2928
rect 4707 2894 4741 2928
rect 4779 2894 4813 2928
rect 4851 2894 4885 2928
rect 4923 2894 4957 2928
rect 4995 2894 5029 2928
rect 5067 2894 5101 2928
rect 5139 2894 5173 2928
rect 5211 2894 5245 2928
rect 5283 2894 5317 2928
rect 5355 2894 5389 2928
rect 5427 2894 5461 2928
rect 5499 2894 5533 2928
rect 5571 2894 5605 2928
rect 5643 2894 5677 2928
rect 5715 2894 5749 2928
rect 5787 2894 5821 2928
rect 5859 2894 5893 2928
rect 5931 2894 5965 2928
rect 6003 2894 6037 2928
rect 6075 2894 6109 2928
rect 6147 2894 6181 2928
rect 6219 2894 6253 2928
rect 6291 2894 6325 2928
rect 6363 2894 6397 2928
rect 6435 2894 6469 2928
rect 6507 2894 6541 2928
rect 6579 2894 6613 2928
rect 6651 2894 6685 2928
rect 6723 2894 6757 2928
rect 6795 2894 6829 2928
rect 6867 2894 6901 2928
rect 6939 2894 6973 2928
rect 7011 2894 7045 2928
rect 7083 2894 7117 2928
rect 7155 2894 7189 2928
rect 7227 2894 7261 2928
rect 7299 2894 7333 2928
rect 7371 2894 7405 2928
rect 7443 2894 7477 2928
rect 7515 2894 7549 2928
rect 7587 2894 7621 2928
rect 7659 2894 7693 2928
rect 7731 2894 7765 2928
rect 7803 2894 7837 2928
rect 7875 2894 7909 2928
rect 7947 2894 7981 2928
rect 8019 2894 8053 2928
rect 8091 2894 8125 2928
rect 8163 2894 8197 2928
rect 8235 2894 8269 2928
rect 8307 2894 8341 2928
rect 8379 2894 8413 2928
rect 8451 2894 8485 2928
rect 8523 2894 8557 2928
rect 8595 2894 8629 2928
rect 8667 2894 8701 2928
rect 8739 2894 8773 2928
rect 8811 2894 8845 2928
rect 8883 2894 8917 2928
rect 8955 2894 8989 2928
rect 9027 2894 9061 2928
rect 9099 2894 9133 2928
rect 9171 2894 9205 2928
rect 9243 2894 9277 2928
rect 9315 2894 9349 2928
rect 9387 2894 9421 2928
rect 9459 2894 9493 2928
rect 9531 2894 9565 2928
rect 9603 2894 9637 2928
rect 9675 2894 9709 2928
rect 9747 2894 9781 2928
rect 9819 2894 9853 2928
rect 9891 2894 9925 2928
rect 9963 2894 9997 2928
rect 10035 2894 10069 2928
rect 10107 2894 10141 2928
rect 10179 2894 10213 2928
rect 10251 2894 10285 2928
rect 10323 2894 10357 2928
rect 10395 2894 10429 2928
rect 10467 2894 10501 2928
rect 10539 2894 10573 2928
rect 10611 2894 10645 2928
rect 10683 2894 10717 2928
rect 10755 2894 10789 2928
rect 10827 2894 10861 2928
rect 10899 2894 10933 2928
rect 10971 2894 11005 2928
rect 11043 2894 11077 2928
rect 11115 2894 11149 2928
rect 11187 2894 11221 2928
rect 11259 2894 11293 2928
rect 11331 2894 11365 2928
rect 11403 2894 11437 2928
rect 11475 2894 11509 2928
rect 11547 2894 11581 2928
rect 11619 2894 11653 2928
rect 11691 2894 11725 2928
rect 11763 2894 11797 2928
rect 11835 2894 11869 2928
rect 11907 2894 11941 2928
rect 11979 2894 12013 2928
rect 12051 2894 12085 2928
rect 12123 2894 12157 2928
rect 12195 2894 12229 2928
rect 12267 2894 12301 2928
rect 12339 2894 12373 2928
rect 12411 2894 12445 2928
rect 12483 2894 12517 2928
rect 12555 2894 12589 2928
rect 12627 2894 12661 2928
rect 12699 2894 12733 2928
rect 12771 2894 12805 2928
rect 12843 2894 12877 2928
rect 12915 2894 12949 2928
rect 12987 2894 13021 2928
rect 13059 2894 13093 2928
rect 13131 2894 13165 2928
rect 13203 2894 13237 2928
rect 13275 2894 13309 2928
rect 13347 2894 13381 2928
rect 13419 2894 13453 2928
rect 13491 2894 13525 2928
rect 13563 2894 13597 2928
rect 13635 2894 13669 2928
rect 13707 2894 13741 2928
rect 13779 2894 13813 2928
rect 13851 2894 13885 2928
rect 13923 2894 13957 2928
rect 13995 2894 14029 2928
rect 14067 2894 14101 2928
rect 14139 2894 14173 2928
rect 14211 2894 14245 2928
rect 14283 2894 14317 2928
rect 14355 2894 14389 2928
rect 14427 2894 14461 2928
rect 14499 2894 14533 2928
rect 14571 2894 14605 2928
rect 14643 2894 14677 2928
rect 14715 2894 14749 2928
rect 14787 2894 14821 2928
rect 14859 2894 14893 2928
rect 14931 2894 14965 2928
rect 15003 2894 15037 2928
rect 15075 2894 15109 2928
rect 15147 2894 15181 2928
rect 15219 2894 15253 2928
rect 15291 2894 15325 2928
rect 15363 2894 15397 2928
rect 15435 2894 15469 2928
rect 15507 2894 15541 2928
rect 15579 2894 15613 2928
rect 15651 2894 15685 2928
rect 15723 2894 15757 2928
rect 15795 2894 15829 2928
rect 15867 2894 15901 2928
rect 15939 2894 15973 2928
rect 16011 2894 16045 2928
rect 16083 2894 16117 2928
rect 16155 2894 16189 2928
rect 16227 2894 16261 2928
rect 16299 2894 16333 2928
rect 16371 2894 16405 2928
rect 16443 2894 16477 2928
rect 16515 2894 16549 2928
rect 16587 2894 16621 2928
rect 16659 2894 16693 2928
rect 16731 2894 16765 2928
rect 16803 2894 16837 2928
rect 16875 2894 16909 2928
rect 16947 2894 16981 2928
rect 17019 2894 17053 2928
rect 17091 2894 17125 2928
rect 17163 2894 17197 2928
rect 17235 2894 17269 2928
rect 17307 2894 17341 2928
rect 17379 2894 17413 2928
rect 17451 2894 17485 2928
rect 17523 2894 17557 2928
rect 17595 2894 17629 2928
rect 17667 2894 17701 2928
rect 17739 2894 17773 2928
rect 17811 2894 17845 2928
rect 17883 2894 17917 2928
rect 17955 2894 17989 2928
rect 18027 2894 18061 2928
rect 18099 2894 18133 2928
rect 18171 2894 18205 2928
rect 18243 2894 18277 2928
rect 18315 2894 18349 2928
rect 18387 2894 18421 2928
rect 18459 2894 18493 2928
rect 18531 2894 18565 2928
rect 18603 2894 18637 2928
rect 18675 2894 18709 2928
rect 18747 2894 18781 2928
rect 18819 2894 18853 2928
rect 18891 2894 18925 2928
rect 18963 2894 18997 2928
rect 19035 2894 19069 2928
rect 19107 2894 19141 2928
rect 19179 2894 19213 2928
rect 19251 2894 19285 2928
rect 19323 2894 19357 2928
rect 19395 2894 19429 2928
rect 19467 2894 19501 2928
rect 19539 2894 19573 2928
rect 19611 2894 19645 2928
rect 19683 2894 19717 2928
rect 19755 2894 19789 2928
rect -1641 2819 -1607 2823
rect -1641 2789 -1607 2819
rect -1641 2717 -1607 2750
rect -1641 2716 -1607 2717
rect -1641 2649 -1607 2676
rect -1641 2642 -1607 2649
rect -1485 2547 -1451 2561
rect -1485 2527 -1451 2547
rect -1485 2479 -1451 2489
rect -1485 2455 -1451 2479
rect -1329 2819 -1295 2823
rect -1329 2789 -1295 2819
rect -1329 2717 -1295 2750
rect -1329 2716 -1295 2717
rect -1329 2649 -1295 2676
rect -1329 2642 -1295 2649
rect -1198 2819 -1164 2823
rect -1198 2789 -1164 2819
rect -1198 2717 -1164 2750
rect -1198 2716 -1164 2717
rect -1198 2649 -1164 2676
rect -1198 2642 -1164 2649
rect -1042 2445 -1008 2475
rect -1042 2441 -1008 2445
rect -1042 2377 -1008 2403
rect -1042 2369 -1008 2377
rect -886 2819 -852 2823
rect -886 2789 -852 2819
rect -886 2717 -852 2750
rect -886 2716 -852 2717
rect -886 2649 -852 2676
rect -886 2642 -852 2649
rect 19882 2839 19916 2873
rect -46 2760 -12 2794
rect 42 2760 76 2794
rect -46 2687 -12 2721
rect 42 2687 76 2721
rect -46 2614 -12 2648
rect 42 2614 76 2648
rect 19882 2766 19916 2800
rect 19882 2693 19916 2727
rect 19882 2620 19916 2654
rect -46 2541 -12 2575
rect 42 2541 76 2575
rect -46 2468 -12 2502
rect 42 2468 76 2502
rect -46 2395 -12 2429
rect 42 2395 76 2429
rect -46 2322 -12 2356
rect 42 2322 76 2356
rect -46 2249 -12 2283
rect 42 2249 76 2283
rect -46 2176 -12 2210
rect 42 2176 76 2210
rect -1584 2080 -1580 2114
rect -1580 2080 -1550 2114
rect -1503 2080 -1485 2114
rect -1485 2080 -1469 2114
rect -1423 2080 -1390 2114
rect -1390 2080 -1389 2114
rect -1343 2080 -1309 2114
rect -1263 2080 -1229 2114
rect -1183 2080 -1149 2114
rect -1103 2080 -1069 2114
rect -1023 2080 -989 2114
rect -943 2080 -909 2114
rect -46 2103 -12 2137
rect 42 2103 76 2137
rect -46 2030 -12 2064
rect 42 2030 76 2064
rect -1641 2013 -1607 2029
rect -1641 1995 -1607 2013
rect -1641 1945 -1607 1956
rect -1641 1922 -1607 1945
rect -1641 1877 -1607 1882
rect -1641 1848 -1607 1877
rect -1485 1741 -1451 1765
rect -1485 1731 -1451 1741
rect -1485 1673 -1451 1693
rect -1485 1659 -1451 1673
rect -1329 2013 -1295 2029
rect -1329 1995 -1295 2013
rect -1329 1945 -1295 1956
rect -1329 1922 -1295 1945
rect -1329 1877 -1295 1882
rect -1329 1848 -1295 1877
rect -46 1957 -12 1991
rect 42 1957 76 1991
rect -46 1884 -12 1918
rect 42 1884 76 1918
rect -46 1811 -12 1845
rect 42 1811 76 1845
rect -46 1738 -12 1772
rect 42 1738 76 1772
rect -46 1665 -12 1699
rect 42 1665 76 1699
rect 19882 2558 19916 2581
rect 19882 2547 19888 2558
rect 19888 2547 19916 2558
rect 19882 2489 19916 2508
rect 19882 2474 19888 2489
rect 19888 2474 19916 2489
rect 19882 2420 19916 2435
rect 19882 2401 19888 2420
rect 19888 2401 19916 2420
rect 19882 2351 19916 2362
rect 19882 2328 19888 2351
rect 19888 2328 19916 2351
rect 19882 2282 19916 2289
rect 19882 2255 19888 2282
rect 19888 2255 19916 2282
rect 19882 2213 19916 2216
rect 19882 2182 19888 2213
rect 19888 2182 19916 2213
rect 19882 2110 19888 2143
rect 19888 2110 19916 2143
rect 19882 2109 19916 2110
rect 19882 2041 19888 2070
rect 19888 2041 19916 2070
rect 19882 2036 19916 2041
rect 19882 1972 19888 1997
rect 19888 1972 19916 1997
rect 19882 1963 19916 1972
rect 19882 1903 19888 1924
rect 19888 1903 19916 1924
rect 19882 1890 19916 1903
rect 19882 1834 19888 1851
rect 19888 1834 19916 1851
rect 19882 1817 19916 1834
rect 19882 1765 19888 1778
rect 19888 1765 19916 1778
rect 19882 1744 19916 1765
rect 19882 1696 19888 1705
rect 19888 1696 19916 1705
rect 19882 1671 19916 1696
rect -46 1592 -12 1626
rect 42 1592 76 1626
rect -46 1519 -12 1553
rect 42 1519 76 1553
rect 364 1638 398 1640
rect 437 1638 471 1640
rect 510 1638 544 1640
rect 583 1638 617 1640
rect 656 1638 690 1640
rect 729 1638 763 1640
rect 802 1638 836 1640
rect 875 1638 909 1640
rect 948 1638 982 1640
rect 1021 1638 1055 1640
rect 1094 1638 1128 1640
rect 1167 1638 1201 1640
rect 1240 1638 1274 1640
rect 1313 1638 1347 1640
rect 1386 1638 1420 1640
rect 1459 1638 1493 1640
rect 1532 1638 1566 1640
rect 1605 1638 1639 1640
rect 1678 1638 1712 1640
rect 1751 1638 1785 1640
rect 1824 1638 1858 1640
rect 1898 1638 1932 1640
rect 1972 1638 2006 1640
rect 2046 1638 2080 1640
rect 2120 1638 2154 1640
rect 2194 1638 2228 1640
rect 2268 1638 2302 1640
rect 2342 1638 2376 1640
rect 2416 1638 2450 1640
rect 2490 1638 2524 1640
rect 2564 1638 2598 1640
rect 2638 1638 2672 1640
rect 364 1606 398 1638
rect 437 1606 471 1638
rect 510 1606 544 1638
rect 583 1606 617 1638
rect 656 1606 690 1638
rect 729 1606 763 1638
rect 802 1606 836 1638
rect 875 1606 909 1638
rect 948 1606 982 1638
rect 1021 1606 1055 1638
rect 1094 1606 1128 1638
rect 1167 1606 1201 1638
rect 1240 1606 1274 1638
rect 1313 1606 1347 1638
rect 1386 1606 1420 1638
rect 1459 1606 1493 1638
rect 1532 1606 1566 1638
rect 1605 1606 1639 1638
rect 1678 1606 1712 1638
rect 1751 1606 1785 1638
rect 1824 1606 1858 1638
rect 1898 1606 1932 1638
rect 1972 1606 2006 1638
rect 2046 1606 2080 1638
rect 2120 1606 2154 1638
rect 2194 1606 2228 1638
rect 2268 1606 2302 1638
rect 2342 1606 2376 1638
rect 2416 1606 2450 1638
rect 2490 1606 2524 1638
rect 2564 1606 2574 1638
rect 2574 1606 2598 1638
rect 2638 1606 2643 1638
rect 2643 1606 2672 1638
rect 2712 1606 2746 1640
rect 2786 1638 2820 1640
rect 2860 1638 2894 1640
rect 2934 1638 2968 1640
rect 3008 1638 3042 1640
rect 3082 1638 3116 1640
rect 3156 1638 3190 1640
rect 3230 1638 3264 1640
rect 2786 1606 2816 1638
rect 2816 1606 2820 1638
rect 2860 1606 2885 1638
rect 2885 1606 2894 1638
rect 2934 1606 2954 1638
rect 2954 1606 2968 1638
rect 3008 1606 3023 1638
rect 3023 1606 3042 1638
rect 3082 1606 3092 1638
rect 3092 1606 3116 1638
rect 3156 1606 3161 1638
rect 3161 1606 3190 1638
rect 3230 1606 3264 1638
rect 364 1536 398 1568
rect 437 1536 471 1568
rect 510 1536 544 1568
rect 583 1536 617 1568
rect 656 1536 690 1568
rect 729 1536 763 1568
rect 802 1536 836 1568
rect 875 1536 909 1568
rect 948 1536 982 1568
rect 1021 1536 1055 1568
rect 1094 1536 1128 1568
rect 1167 1536 1201 1568
rect 1240 1536 1274 1568
rect 1313 1536 1347 1568
rect 1386 1536 1420 1568
rect 1459 1536 1493 1568
rect 1532 1536 1566 1568
rect 1605 1536 1639 1568
rect 1678 1536 1712 1568
rect 1751 1536 1785 1568
rect 1824 1536 1858 1568
rect 1898 1536 1932 1568
rect 1972 1536 2006 1568
rect 2046 1536 2080 1568
rect 2120 1536 2154 1568
rect 2194 1536 2228 1568
rect 2268 1536 2302 1568
rect 2342 1536 2376 1568
rect 2416 1536 2450 1568
rect 2490 1536 2524 1568
rect 2564 1536 2574 1568
rect 2574 1536 2598 1568
rect 2638 1536 2643 1568
rect 2643 1536 2672 1568
rect 364 1534 398 1536
rect 437 1534 471 1536
rect 510 1534 544 1536
rect 583 1534 617 1536
rect 656 1534 690 1536
rect 729 1534 763 1536
rect 802 1534 836 1536
rect 875 1534 909 1536
rect 948 1534 982 1536
rect 1021 1534 1055 1536
rect 1094 1534 1128 1536
rect 1167 1534 1201 1536
rect 1240 1534 1274 1536
rect 1313 1534 1347 1536
rect 1386 1534 1420 1536
rect 1459 1534 1493 1536
rect 1532 1534 1566 1536
rect 1605 1534 1639 1536
rect 1678 1534 1712 1536
rect 1751 1534 1785 1536
rect 1824 1534 1858 1536
rect 1898 1534 1932 1536
rect 1972 1534 2006 1536
rect 2046 1534 2080 1536
rect 2120 1534 2154 1536
rect 2194 1534 2228 1536
rect 2268 1534 2302 1536
rect 2342 1534 2376 1536
rect 2416 1534 2450 1536
rect 2490 1534 2524 1536
rect 2564 1534 2598 1536
rect 2638 1534 2672 1536
rect 2712 1534 2746 1568
rect 2786 1536 2816 1568
rect 2816 1536 2820 1568
rect 2860 1536 2885 1568
rect 2885 1536 2894 1568
rect 2934 1536 2954 1568
rect 2954 1536 2968 1568
rect 3008 1536 3023 1568
rect 3023 1536 3042 1568
rect 3082 1536 3092 1568
rect 3092 1536 3116 1568
rect 3156 1536 3161 1568
rect 3161 1536 3190 1568
rect 3230 1536 3264 1568
rect 2786 1534 2820 1536
rect 2860 1534 2894 1536
rect 2934 1534 2968 1536
rect 3008 1534 3042 1536
rect 3082 1534 3116 1536
rect 3156 1534 3190 1536
rect 3230 1534 3264 1536
rect 3606 1638 3640 1640
rect 3680 1638 3714 1640
rect 3754 1638 3788 1640
rect 3828 1638 3862 1640
rect 3902 1638 3936 1640
rect 3976 1638 4010 1640
rect 4050 1638 4084 1640
rect 3606 1606 3640 1638
rect 3680 1606 3709 1638
rect 3709 1606 3714 1638
rect 3754 1606 3778 1638
rect 3778 1606 3788 1638
rect 3828 1606 3847 1638
rect 3847 1606 3862 1638
rect 3902 1606 3916 1638
rect 3916 1606 3936 1638
rect 3976 1606 3985 1638
rect 3985 1606 4010 1638
rect 4050 1606 4054 1638
rect 4054 1606 4084 1638
rect 4124 1606 4158 1640
rect 4198 1638 4232 1640
rect 4272 1638 4306 1640
rect 4346 1638 4380 1640
rect 4420 1638 4454 1640
rect 4494 1638 4528 1640
rect 4568 1638 4602 1640
rect 4642 1638 4676 1640
rect 4716 1638 4750 1640
rect 4790 1638 4824 1640
rect 4864 1638 4898 1640
rect 4938 1638 4972 1640
rect 5012 1638 5046 1640
rect 5085 1638 5119 1640
rect 5158 1638 5192 1640
rect 5231 1638 5265 1640
rect 5304 1638 5338 1640
rect 5377 1638 5411 1640
rect 5450 1638 5484 1640
rect 5523 1638 5557 1640
rect 5596 1638 5630 1640
rect 5669 1638 5703 1640
rect 5742 1638 5776 1640
rect 5815 1638 5849 1640
rect 5888 1638 5922 1640
rect 5961 1638 5995 1640
rect 6034 1638 6068 1640
rect 6107 1638 6141 1640
rect 6180 1638 6214 1640
rect 6253 1638 6287 1640
rect 6326 1638 6360 1640
rect 6399 1638 6433 1640
rect 6472 1638 6506 1640
rect 4198 1606 4227 1638
rect 4227 1606 4232 1638
rect 4272 1606 4296 1638
rect 4296 1606 4306 1638
rect 4346 1606 4380 1638
rect 4420 1606 4454 1638
rect 4494 1606 4528 1638
rect 4568 1606 4602 1638
rect 4642 1606 4676 1638
rect 4716 1606 4750 1638
rect 4790 1606 4824 1638
rect 4864 1606 4898 1638
rect 4938 1606 4972 1638
rect 5012 1606 5046 1638
rect 5085 1606 5119 1638
rect 5158 1606 5192 1638
rect 5231 1606 5265 1638
rect 5304 1606 5338 1638
rect 5377 1606 5411 1638
rect 5450 1606 5484 1638
rect 5523 1606 5557 1638
rect 5596 1606 5630 1638
rect 5669 1606 5703 1638
rect 5742 1606 5776 1638
rect 5815 1606 5849 1638
rect 5888 1606 5922 1638
rect 5961 1606 5995 1638
rect 6034 1606 6068 1638
rect 6107 1606 6141 1638
rect 6180 1606 6214 1638
rect 6253 1606 6287 1638
rect 6326 1606 6360 1638
rect 6399 1606 6433 1638
rect 6472 1606 6506 1638
rect 3606 1536 3640 1568
rect 3680 1536 3709 1568
rect 3709 1536 3714 1568
rect 3754 1536 3778 1568
rect 3778 1536 3788 1568
rect 3828 1536 3847 1568
rect 3847 1536 3862 1568
rect 3902 1536 3916 1568
rect 3916 1536 3936 1568
rect 3976 1536 3985 1568
rect 3985 1536 4010 1568
rect 4050 1536 4054 1568
rect 4054 1536 4084 1568
rect 3606 1534 3640 1536
rect 3680 1534 3714 1536
rect 3754 1534 3788 1536
rect 3828 1534 3862 1536
rect 3902 1534 3936 1536
rect 3976 1534 4010 1536
rect 4050 1534 4084 1536
rect 4124 1534 4158 1568
rect 4198 1536 4227 1568
rect 4227 1536 4232 1568
rect 4272 1536 4296 1568
rect 4296 1536 4306 1568
rect 4346 1536 4380 1568
rect 4420 1536 4454 1568
rect 4494 1536 4528 1568
rect 4568 1536 4602 1568
rect 4642 1536 4676 1568
rect 4716 1536 4750 1568
rect 4790 1536 4824 1568
rect 4864 1536 4898 1568
rect 4938 1536 4972 1568
rect 5012 1536 5046 1568
rect 5085 1536 5119 1568
rect 5158 1536 5192 1568
rect 5231 1536 5265 1568
rect 5304 1536 5338 1568
rect 5377 1536 5411 1568
rect 5450 1536 5484 1568
rect 5523 1536 5557 1568
rect 5596 1536 5630 1568
rect 5669 1536 5703 1568
rect 5742 1536 5776 1568
rect 5815 1536 5849 1568
rect 5888 1536 5922 1568
rect 5961 1536 5995 1568
rect 6034 1536 6068 1568
rect 6107 1536 6141 1568
rect 6180 1536 6214 1568
rect 6253 1536 6287 1568
rect 6326 1536 6360 1568
rect 6399 1536 6433 1568
rect 6472 1536 6506 1568
rect 4198 1534 4232 1536
rect 4272 1534 4306 1536
rect 4346 1534 4380 1536
rect 4420 1534 4454 1536
rect 4494 1534 4528 1536
rect 4568 1534 4602 1536
rect 4642 1534 4676 1536
rect 4716 1534 4750 1536
rect 4790 1534 4824 1536
rect 4864 1534 4898 1536
rect 4938 1534 4972 1536
rect 5012 1534 5046 1536
rect 5085 1534 5119 1536
rect 5158 1534 5192 1536
rect 5231 1534 5265 1536
rect 5304 1534 5338 1536
rect 5377 1534 5411 1536
rect 5450 1534 5484 1536
rect 5523 1534 5557 1536
rect 5596 1534 5630 1536
rect 5669 1534 5703 1536
rect 5742 1534 5776 1536
rect 5815 1534 5849 1536
rect 5888 1534 5922 1536
rect 5961 1534 5995 1536
rect 6034 1534 6068 1536
rect 6107 1534 6141 1536
rect 6180 1534 6214 1536
rect 6253 1534 6287 1536
rect 6326 1534 6360 1536
rect 6399 1534 6433 1536
rect 6472 1534 6506 1536
rect 6848 1638 6882 1640
rect 6921 1638 6955 1640
rect 6994 1638 7028 1640
rect 7067 1638 7101 1640
rect 7140 1638 7174 1640
rect 7213 1638 7247 1640
rect 7286 1638 7320 1640
rect 7359 1638 7393 1640
rect 7432 1638 7466 1640
rect 7505 1638 7539 1640
rect 7578 1638 7612 1640
rect 7651 1638 7685 1640
rect 7724 1638 7758 1640
rect 7797 1638 7831 1640
rect 7870 1638 7904 1640
rect 7943 1638 7977 1640
rect 8016 1638 8050 1640
rect 8089 1638 8123 1640
rect 8162 1638 8196 1640
rect 8235 1638 8269 1640
rect 8308 1638 8342 1640
rect 8382 1638 8416 1640
rect 8456 1638 8490 1640
rect 8530 1638 8564 1640
rect 8604 1638 8638 1640
rect 8678 1638 8712 1640
rect 8752 1638 8786 1640
rect 8826 1638 8860 1640
rect 8900 1638 8934 1640
rect 8974 1638 9008 1640
rect 9048 1638 9082 1640
rect 9122 1638 9156 1640
rect 6848 1606 6882 1638
rect 6921 1606 6955 1638
rect 6994 1606 7028 1638
rect 7067 1606 7101 1638
rect 7140 1606 7174 1638
rect 7213 1606 7247 1638
rect 7286 1606 7320 1638
rect 7359 1606 7393 1638
rect 7432 1606 7466 1638
rect 7505 1606 7539 1638
rect 7578 1606 7612 1638
rect 7651 1606 7685 1638
rect 7724 1606 7758 1638
rect 7797 1606 7831 1638
rect 7870 1606 7904 1638
rect 7943 1606 7977 1638
rect 8016 1606 8050 1638
rect 8089 1606 8123 1638
rect 8162 1606 8196 1638
rect 8235 1606 8269 1638
rect 8308 1606 8342 1638
rect 8382 1606 8416 1638
rect 8456 1606 8490 1638
rect 8530 1606 8564 1638
rect 8604 1606 8638 1638
rect 8678 1606 8712 1638
rect 8752 1606 8786 1638
rect 8826 1606 8860 1638
rect 8900 1606 8934 1638
rect 8974 1606 9008 1638
rect 9048 1606 9058 1638
rect 9058 1606 9082 1638
rect 9122 1606 9127 1638
rect 9127 1606 9156 1638
rect 9196 1606 9230 1640
rect 9270 1638 9304 1640
rect 9344 1638 9378 1640
rect 9418 1638 9452 1640
rect 9492 1638 9526 1640
rect 9566 1638 9600 1640
rect 9640 1638 9674 1640
rect 9714 1638 9748 1640
rect 9270 1606 9300 1638
rect 9300 1606 9304 1638
rect 9344 1606 9369 1638
rect 9369 1606 9378 1638
rect 9418 1606 9438 1638
rect 9438 1606 9452 1638
rect 9492 1606 9507 1638
rect 9507 1606 9526 1638
rect 9566 1606 9576 1638
rect 9576 1606 9600 1638
rect 9640 1606 9645 1638
rect 9645 1606 9674 1638
rect 9714 1606 9748 1638
rect 6848 1536 6882 1568
rect 6921 1536 6955 1568
rect 6994 1536 7028 1568
rect 7067 1536 7101 1568
rect 7140 1536 7174 1568
rect 7213 1536 7247 1568
rect 7286 1536 7320 1568
rect 7359 1536 7393 1568
rect 7432 1536 7466 1568
rect 7505 1536 7539 1568
rect 7578 1536 7612 1568
rect 7651 1536 7685 1568
rect 7724 1536 7758 1568
rect 7797 1536 7831 1568
rect 7870 1536 7904 1568
rect 7943 1536 7977 1568
rect 8016 1536 8050 1568
rect 8089 1536 8123 1568
rect 8162 1536 8196 1568
rect 8235 1536 8269 1568
rect 8308 1536 8342 1568
rect 8382 1536 8416 1568
rect 8456 1536 8490 1568
rect 8530 1536 8564 1568
rect 8604 1536 8638 1568
rect 8678 1536 8712 1568
rect 8752 1536 8786 1568
rect 8826 1536 8860 1568
rect 8900 1536 8934 1568
rect 8974 1536 9008 1568
rect 9048 1536 9058 1568
rect 9058 1536 9082 1568
rect 9122 1536 9127 1568
rect 9127 1536 9156 1568
rect 6848 1534 6882 1536
rect 6921 1534 6955 1536
rect 6994 1534 7028 1536
rect 7067 1534 7101 1536
rect 7140 1534 7174 1536
rect 7213 1534 7247 1536
rect 7286 1534 7320 1536
rect 7359 1534 7393 1536
rect 7432 1534 7466 1536
rect 7505 1534 7539 1536
rect 7578 1534 7612 1536
rect 7651 1534 7685 1536
rect 7724 1534 7758 1536
rect 7797 1534 7831 1536
rect 7870 1534 7904 1536
rect 7943 1534 7977 1536
rect 8016 1534 8050 1536
rect 8089 1534 8123 1536
rect 8162 1534 8196 1536
rect 8235 1534 8269 1536
rect 8308 1534 8342 1536
rect 8382 1534 8416 1536
rect 8456 1534 8490 1536
rect 8530 1534 8564 1536
rect 8604 1534 8638 1536
rect 8678 1534 8712 1536
rect 8752 1534 8786 1536
rect 8826 1534 8860 1536
rect 8900 1534 8934 1536
rect 8974 1534 9008 1536
rect 9048 1534 9082 1536
rect 9122 1534 9156 1536
rect 9196 1534 9230 1568
rect 9270 1536 9300 1568
rect 9300 1536 9304 1568
rect 9344 1536 9369 1568
rect 9369 1536 9378 1568
rect 9418 1536 9438 1568
rect 9438 1536 9452 1568
rect 9492 1536 9507 1568
rect 9507 1536 9526 1568
rect 9566 1536 9576 1568
rect 9576 1536 9600 1568
rect 9640 1536 9645 1568
rect 9645 1536 9674 1568
rect 9714 1536 9748 1568
rect 9270 1534 9304 1536
rect 9344 1534 9378 1536
rect 9418 1534 9452 1536
rect 9492 1534 9526 1536
rect 9566 1534 9600 1536
rect 9640 1534 9674 1536
rect 9714 1534 9748 1536
rect 10090 1638 10124 1640
rect 10164 1638 10198 1640
rect 10238 1638 10272 1640
rect 10312 1638 10346 1640
rect 10386 1638 10420 1640
rect 10460 1638 10494 1640
rect 10534 1638 10568 1640
rect 10090 1606 10124 1638
rect 10164 1606 10193 1638
rect 10193 1606 10198 1638
rect 10238 1606 10262 1638
rect 10262 1606 10272 1638
rect 10312 1606 10331 1638
rect 10331 1606 10346 1638
rect 10386 1606 10400 1638
rect 10400 1606 10420 1638
rect 10460 1606 10469 1638
rect 10469 1606 10494 1638
rect 10534 1606 10538 1638
rect 10538 1606 10568 1638
rect 10608 1606 10642 1640
rect 10682 1638 10716 1640
rect 10756 1638 10790 1640
rect 10830 1638 10864 1640
rect 10904 1638 10938 1640
rect 10978 1638 11012 1640
rect 11052 1638 11086 1640
rect 11126 1638 11160 1640
rect 11200 1638 11234 1640
rect 11274 1638 11308 1640
rect 11348 1638 11382 1640
rect 11422 1638 11456 1640
rect 11496 1638 11530 1640
rect 11569 1638 11603 1640
rect 11642 1638 11676 1640
rect 11715 1638 11749 1640
rect 11788 1638 11822 1640
rect 11861 1638 11895 1640
rect 11934 1638 11968 1640
rect 12007 1638 12041 1640
rect 12080 1638 12114 1640
rect 12153 1638 12187 1640
rect 12226 1638 12260 1640
rect 12299 1638 12333 1640
rect 12372 1638 12406 1640
rect 12445 1638 12479 1640
rect 12518 1638 12552 1640
rect 12591 1638 12625 1640
rect 12664 1638 12698 1640
rect 12737 1638 12771 1640
rect 12810 1638 12844 1640
rect 12883 1638 12917 1640
rect 12956 1638 12990 1640
rect 10682 1606 10711 1638
rect 10711 1606 10716 1638
rect 10756 1606 10780 1638
rect 10780 1606 10790 1638
rect 10830 1606 10864 1638
rect 10904 1606 10938 1638
rect 10978 1606 11012 1638
rect 11052 1606 11086 1638
rect 11126 1606 11160 1638
rect 11200 1606 11234 1638
rect 11274 1606 11308 1638
rect 11348 1606 11382 1638
rect 11422 1606 11456 1638
rect 11496 1606 11530 1638
rect 11569 1606 11603 1638
rect 11642 1606 11676 1638
rect 11715 1606 11749 1638
rect 11788 1606 11822 1638
rect 11861 1606 11895 1638
rect 11934 1606 11968 1638
rect 12007 1606 12041 1638
rect 12080 1606 12114 1638
rect 12153 1606 12187 1638
rect 12226 1606 12260 1638
rect 12299 1606 12333 1638
rect 12372 1606 12406 1638
rect 12445 1606 12479 1638
rect 12518 1606 12552 1638
rect 12591 1606 12625 1638
rect 12664 1606 12698 1638
rect 12737 1606 12771 1638
rect 12810 1606 12844 1638
rect 12883 1606 12917 1638
rect 12956 1606 12990 1638
rect 10090 1536 10124 1568
rect 10164 1536 10193 1568
rect 10193 1536 10198 1568
rect 10238 1536 10262 1568
rect 10262 1536 10272 1568
rect 10312 1536 10331 1568
rect 10331 1536 10346 1568
rect 10386 1536 10400 1568
rect 10400 1536 10420 1568
rect 10460 1536 10469 1568
rect 10469 1536 10494 1568
rect 10534 1536 10538 1568
rect 10538 1536 10568 1568
rect 10090 1534 10124 1536
rect 10164 1534 10198 1536
rect 10238 1534 10272 1536
rect 10312 1534 10346 1536
rect 10386 1534 10420 1536
rect 10460 1534 10494 1536
rect 10534 1534 10568 1536
rect 10608 1534 10642 1568
rect 10682 1536 10711 1568
rect 10711 1536 10716 1568
rect 10756 1536 10780 1568
rect 10780 1536 10790 1568
rect 10830 1536 10864 1568
rect 10904 1536 10938 1568
rect 10978 1536 11012 1568
rect 11052 1536 11086 1568
rect 11126 1536 11160 1568
rect 11200 1536 11234 1568
rect 11274 1536 11308 1568
rect 11348 1536 11382 1568
rect 11422 1536 11456 1568
rect 11496 1536 11530 1568
rect 11569 1536 11603 1568
rect 11642 1536 11676 1568
rect 11715 1536 11749 1568
rect 11788 1536 11822 1568
rect 11861 1536 11895 1568
rect 11934 1536 11968 1568
rect 12007 1536 12041 1568
rect 12080 1536 12114 1568
rect 12153 1536 12187 1568
rect 12226 1536 12260 1568
rect 12299 1536 12333 1568
rect 12372 1536 12406 1568
rect 12445 1536 12479 1568
rect 12518 1536 12552 1568
rect 12591 1536 12625 1568
rect 12664 1536 12698 1568
rect 12737 1536 12771 1568
rect 12810 1536 12844 1568
rect 12883 1536 12917 1568
rect 12956 1536 12990 1568
rect 10682 1534 10716 1536
rect 10756 1534 10790 1536
rect 10830 1534 10864 1536
rect 10904 1534 10938 1536
rect 10978 1534 11012 1536
rect 11052 1534 11086 1536
rect 11126 1534 11160 1536
rect 11200 1534 11234 1536
rect 11274 1534 11308 1536
rect 11348 1534 11382 1536
rect 11422 1534 11456 1536
rect 11496 1534 11530 1536
rect 11569 1534 11603 1536
rect 11642 1534 11676 1536
rect 11715 1534 11749 1536
rect 11788 1534 11822 1536
rect 11861 1534 11895 1536
rect 11934 1534 11968 1536
rect 12007 1534 12041 1536
rect 12080 1534 12114 1536
rect 12153 1534 12187 1536
rect 12226 1534 12260 1536
rect 12299 1534 12333 1536
rect 12372 1534 12406 1536
rect 12445 1534 12479 1536
rect 12518 1534 12552 1536
rect 12591 1534 12625 1536
rect 12664 1534 12698 1536
rect 12737 1534 12771 1536
rect 12810 1534 12844 1536
rect 12883 1534 12917 1536
rect 12956 1534 12990 1536
rect 13332 1638 13366 1640
rect 13405 1638 13439 1640
rect 13478 1638 13512 1640
rect 13551 1638 13585 1640
rect 13624 1638 13658 1640
rect 13697 1638 13731 1640
rect 13770 1638 13804 1640
rect 13843 1638 13877 1640
rect 13916 1638 13950 1640
rect 13989 1638 14023 1640
rect 14062 1638 14096 1640
rect 14135 1638 14169 1640
rect 14208 1638 14242 1640
rect 14281 1638 14315 1640
rect 14354 1638 14388 1640
rect 14427 1638 14461 1640
rect 14500 1638 14534 1640
rect 14573 1638 14607 1640
rect 14646 1638 14680 1640
rect 14719 1638 14753 1640
rect 14792 1638 14826 1640
rect 14866 1638 14900 1640
rect 14940 1638 14974 1640
rect 15014 1638 15048 1640
rect 15088 1638 15122 1640
rect 15162 1638 15196 1640
rect 15236 1638 15270 1640
rect 15310 1638 15344 1640
rect 15384 1638 15418 1640
rect 15458 1638 15492 1640
rect 15532 1638 15566 1640
rect 15606 1638 15640 1640
rect 13332 1606 13366 1638
rect 13405 1606 13439 1638
rect 13478 1606 13512 1638
rect 13551 1606 13585 1638
rect 13624 1606 13658 1638
rect 13697 1606 13731 1638
rect 13770 1606 13804 1638
rect 13843 1606 13877 1638
rect 13916 1606 13950 1638
rect 13989 1606 14023 1638
rect 14062 1606 14096 1638
rect 14135 1606 14169 1638
rect 14208 1606 14242 1638
rect 14281 1606 14315 1638
rect 14354 1606 14388 1638
rect 14427 1606 14461 1638
rect 14500 1606 14534 1638
rect 14573 1606 14607 1638
rect 14646 1606 14680 1638
rect 14719 1606 14753 1638
rect 14792 1606 14826 1638
rect 14866 1606 14900 1638
rect 14940 1606 14974 1638
rect 15014 1606 15048 1638
rect 15088 1606 15122 1638
rect 15162 1606 15196 1638
rect 15236 1606 15270 1638
rect 15310 1606 15344 1638
rect 15384 1606 15418 1638
rect 15458 1606 15492 1638
rect 15532 1606 15542 1638
rect 15542 1606 15566 1638
rect 15606 1606 15611 1638
rect 15611 1606 15640 1638
rect 15680 1606 15714 1640
rect 15754 1638 15788 1640
rect 15828 1638 15862 1640
rect 15902 1638 15936 1640
rect 15976 1638 16010 1640
rect 16050 1638 16084 1640
rect 16124 1638 16158 1640
rect 16198 1638 16232 1640
rect 15754 1606 15784 1638
rect 15784 1606 15788 1638
rect 15828 1606 15853 1638
rect 15853 1606 15862 1638
rect 15902 1606 15922 1638
rect 15922 1606 15936 1638
rect 15976 1606 15991 1638
rect 15991 1606 16010 1638
rect 16050 1606 16060 1638
rect 16060 1606 16084 1638
rect 16124 1606 16129 1638
rect 16129 1606 16158 1638
rect 16198 1606 16232 1638
rect 13332 1536 13366 1568
rect 13405 1536 13439 1568
rect 13478 1536 13512 1568
rect 13551 1536 13585 1568
rect 13624 1536 13658 1568
rect 13697 1536 13731 1568
rect 13770 1536 13804 1568
rect 13843 1536 13877 1568
rect 13916 1536 13950 1568
rect 13989 1536 14023 1568
rect 14062 1536 14096 1568
rect 14135 1536 14169 1568
rect 14208 1536 14242 1568
rect 14281 1536 14315 1568
rect 14354 1536 14388 1568
rect 14427 1536 14461 1568
rect 14500 1536 14534 1568
rect 14573 1536 14607 1568
rect 14646 1536 14680 1568
rect 14719 1536 14753 1568
rect 14792 1536 14826 1568
rect 14866 1536 14900 1568
rect 14940 1536 14974 1568
rect 15014 1536 15048 1568
rect 15088 1536 15122 1568
rect 15162 1536 15196 1568
rect 15236 1536 15270 1568
rect 15310 1536 15344 1568
rect 15384 1536 15418 1568
rect 15458 1536 15492 1568
rect 15532 1536 15542 1568
rect 15542 1536 15566 1568
rect 15606 1536 15611 1568
rect 15611 1536 15640 1568
rect 13332 1534 13366 1536
rect 13405 1534 13439 1536
rect 13478 1534 13512 1536
rect 13551 1534 13585 1536
rect 13624 1534 13658 1536
rect 13697 1534 13731 1536
rect 13770 1534 13804 1536
rect 13843 1534 13877 1536
rect 13916 1534 13950 1536
rect 13989 1534 14023 1536
rect 14062 1534 14096 1536
rect 14135 1534 14169 1536
rect 14208 1534 14242 1536
rect 14281 1534 14315 1536
rect 14354 1534 14388 1536
rect 14427 1534 14461 1536
rect 14500 1534 14534 1536
rect 14573 1534 14607 1536
rect 14646 1534 14680 1536
rect 14719 1534 14753 1536
rect 14792 1534 14826 1536
rect 14866 1534 14900 1536
rect 14940 1534 14974 1536
rect 15014 1534 15048 1536
rect 15088 1534 15122 1536
rect 15162 1534 15196 1536
rect 15236 1534 15270 1536
rect 15310 1534 15344 1536
rect 15384 1534 15418 1536
rect 15458 1534 15492 1536
rect 15532 1534 15566 1536
rect 15606 1534 15640 1536
rect 15680 1534 15714 1568
rect 15754 1536 15784 1568
rect 15784 1536 15788 1568
rect 15828 1536 15853 1568
rect 15853 1536 15862 1568
rect 15902 1536 15922 1568
rect 15922 1536 15936 1568
rect 15976 1536 15991 1568
rect 15991 1536 16010 1568
rect 16050 1536 16060 1568
rect 16060 1536 16084 1568
rect 16124 1536 16129 1568
rect 16129 1536 16158 1568
rect 16198 1536 16232 1568
rect 15754 1534 15788 1536
rect 15828 1534 15862 1536
rect 15902 1534 15936 1536
rect 15976 1534 16010 1536
rect 16050 1534 16084 1536
rect 16124 1534 16158 1536
rect 16198 1534 16232 1536
rect 16574 1638 16608 1640
rect 16648 1638 16682 1640
rect 16722 1638 16756 1640
rect 16796 1638 16830 1640
rect 16870 1638 16904 1640
rect 16944 1638 16978 1640
rect 17018 1638 17052 1640
rect 16574 1606 16608 1638
rect 16648 1606 16677 1638
rect 16677 1606 16682 1638
rect 16722 1606 16746 1638
rect 16746 1606 16756 1638
rect 16796 1606 16815 1638
rect 16815 1606 16830 1638
rect 16870 1606 16884 1638
rect 16884 1606 16904 1638
rect 16944 1606 16953 1638
rect 16953 1606 16978 1638
rect 17018 1606 17022 1638
rect 17022 1606 17052 1638
rect 17092 1606 17126 1640
rect 17166 1638 17200 1640
rect 17240 1638 17274 1640
rect 17314 1638 17348 1640
rect 17388 1638 17422 1640
rect 17462 1638 17496 1640
rect 17536 1638 17570 1640
rect 17610 1638 17644 1640
rect 17684 1638 17718 1640
rect 17758 1638 17792 1640
rect 17832 1638 17866 1640
rect 17906 1638 17940 1640
rect 17980 1638 18014 1640
rect 18053 1638 18087 1640
rect 18126 1638 18160 1640
rect 18199 1638 18233 1640
rect 18272 1638 18306 1640
rect 18345 1638 18379 1640
rect 18418 1638 18452 1640
rect 18491 1638 18525 1640
rect 18564 1638 18598 1640
rect 18637 1638 18671 1640
rect 18710 1638 18744 1640
rect 18783 1638 18817 1640
rect 18856 1638 18890 1640
rect 18929 1638 18963 1640
rect 19002 1638 19036 1640
rect 19075 1638 19109 1640
rect 19148 1638 19182 1640
rect 19221 1638 19255 1640
rect 19294 1638 19328 1640
rect 19367 1638 19401 1640
rect 19440 1638 19474 1640
rect 17166 1606 17195 1638
rect 17195 1606 17200 1638
rect 17240 1606 17264 1638
rect 17264 1606 17274 1638
rect 17314 1606 17348 1638
rect 17388 1606 17422 1638
rect 17462 1606 17496 1638
rect 17536 1606 17570 1638
rect 17610 1606 17644 1638
rect 17684 1606 17718 1638
rect 17758 1606 17792 1638
rect 17832 1606 17866 1638
rect 17906 1606 17940 1638
rect 17980 1606 18014 1638
rect 18053 1606 18087 1638
rect 18126 1606 18160 1638
rect 18199 1606 18233 1638
rect 18272 1606 18306 1638
rect 18345 1606 18379 1638
rect 18418 1606 18452 1638
rect 18491 1606 18525 1638
rect 18564 1606 18598 1638
rect 18637 1606 18671 1638
rect 18710 1606 18744 1638
rect 18783 1606 18817 1638
rect 18856 1606 18890 1638
rect 18929 1606 18963 1638
rect 19002 1606 19036 1638
rect 19075 1606 19109 1638
rect 19148 1606 19182 1638
rect 19221 1606 19255 1638
rect 19294 1606 19328 1638
rect 19367 1606 19401 1638
rect 19440 1606 19474 1638
rect 16574 1536 16608 1568
rect 16648 1536 16677 1568
rect 16677 1536 16682 1568
rect 16722 1536 16746 1568
rect 16746 1536 16756 1568
rect 16796 1536 16815 1568
rect 16815 1536 16830 1568
rect 16870 1536 16884 1568
rect 16884 1536 16904 1568
rect 16944 1536 16953 1568
rect 16953 1536 16978 1568
rect 17018 1536 17022 1568
rect 17022 1536 17052 1568
rect 16574 1534 16608 1536
rect 16648 1534 16682 1536
rect 16722 1534 16756 1536
rect 16796 1534 16830 1536
rect 16870 1534 16904 1536
rect 16944 1534 16978 1536
rect 17018 1534 17052 1536
rect 17092 1534 17126 1568
rect 17166 1536 17195 1568
rect 17195 1536 17200 1568
rect 17240 1536 17264 1568
rect 17264 1536 17274 1568
rect 17314 1536 17348 1568
rect 17388 1536 17422 1568
rect 17462 1536 17496 1568
rect 17536 1536 17570 1568
rect 17610 1536 17644 1568
rect 17684 1536 17718 1568
rect 17758 1536 17792 1568
rect 17832 1536 17866 1568
rect 17906 1536 17940 1568
rect 17980 1536 18014 1568
rect 18053 1536 18087 1568
rect 18126 1536 18160 1568
rect 18199 1536 18233 1568
rect 18272 1536 18306 1568
rect 18345 1536 18379 1568
rect 18418 1536 18452 1568
rect 18491 1536 18525 1568
rect 18564 1536 18598 1568
rect 18637 1536 18671 1568
rect 18710 1536 18744 1568
rect 18783 1536 18817 1568
rect 18856 1536 18890 1568
rect 18929 1536 18963 1568
rect 19002 1536 19036 1568
rect 19075 1536 19109 1568
rect 19148 1536 19182 1568
rect 19221 1536 19255 1568
rect 19294 1536 19328 1568
rect 19367 1536 19401 1568
rect 19440 1536 19474 1568
rect 17166 1534 17200 1536
rect 17240 1534 17274 1536
rect 17314 1534 17348 1536
rect 17388 1534 17422 1536
rect 17462 1534 17496 1536
rect 17536 1534 17570 1536
rect 17610 1534 17644 1536
rect 17684 1534 17718 1536
rect 17758 1534 17792 1536
rect 17832 1534 17866 1536
rect 17906 1534 17940 1536
rect 17980 1534 18014 1536
rect 18053 1534 18087 1536
rect 18126 1534 18160 1536
rect 18199 1534 18233 1536
rect 18272 1534 18306 1536
rect 18345 1534 18379 1536
rect 18418 1534 18452 1536
rect 18491 1534 18525 1536
rect 18564 1534 18598 1536
rect 18637 1534 18671 1536
rect 18710 1534 18744 1536
rect 18783 1534 18817 1536
rect 18856 1534 18890 1536
rect 18929 1534 18963 1536
rect 19002 1534 19036 1536
rect 19075 1534 19109 1536
rect 19148 1534 19182 1536
rect 19221 1534 19255 1536
rect 19294 1534 19328 1536
rect 19367 1534 19401 1536
rect 19440 1534 19474 1536
rect 19882 1627 19888 1632
rect 19888 1627 19916 1632
rect 19882 1598 19916 1627
rect -46 1445 -12 1479
rect 42 1445 76 1479
rect 19882 1558 19888 1559
rect 19888 1558 19916 1559
rect 19882 1525 19916 1558
rect 19882 1454 19916 1486
rect 19882 1452 19888 1454
rect 19888 1452 19916 1454
rect 168 1432 202 1446
rect 168 1412 182 1432
rect 182 1412 202 1432
rect 240 1412 274 1446
rect 3386 1412 3420 1446
rect -46 1371 -12 1405
rect 42 1371 76 1405
rect -46 1297 -12 1331
rect 42 1297 76 1331
rect 3458 1412 3492 1446
rect 9870 1412 9904 1446
rect 9942 1412 9976 1446
rect 16354 1412 16388 1446
rect 16426 1412 16460 1446
rect 19564 1412 19598 1446
rect 19636 1432 19670 1446
rect 19636 1412 19656 1432
rect 19656 1412 19670 1432
rect 19882 1385 19916 1413
rect 19882 1379 19888 1385
rect 19888 1379 19916 1385
rect -46 1223 -12 1257
rect 42 1223 76 1257
rect 19882 1316 19916 1340
rect 19882 1306 19888 1316
rect 19888 1306 19916 1316
rect 19882 1247 19916 1267
rect 19882 1233 19888 1247
rect 19888 1233 19916 1247
rect -46 1149 -12 1183
rect 42 1149 76 1183
rect 364 1226 398 1228
rect 437 1226 471 1228
rect 510 1226 544 1228
rect 583 1226 617 1228
rect 656 1226 690 1228
rect 729 1226 763 1228
rect 802 1226 836 1228
rect 875 1226 909 1228
rect 948 1226 982 1228
rect 1021 1226 1055 1228
rect 1094 1226 1128 1228
rect 1167 1226 1201 1228
rect 1240 1226 1274 1228
rect 1313 1226 1347 1228
rect 1386 1226 1420 1228
rect 1459 1226 1493 1228
rect 1532 1226 1566 1228
rect 1605 1226 1639 1228
rect 1678 1226 1712 1228
rect 1751 1226 1785 1228
rect 1824 1226 1858 1228
rect 1898 1226 1932 1228
rect 1972 1226 2006 1228
rect 2046 1226 2080 1228
rect 2120 1226 2154 1228
rect 2194 1226 2228 1228
rect 2268 1226 2302 1228
rect 2342 1226 2376 1228
rect 2416 1226 2450 1228
rect 2490 1226 2524 1228
rect 2564 1226 2598 1228
rect 2638 1226 2672 1228
rect 364 1194 398 1226
rect 437 1194 471 1226
rect 510 1194 544 1226
rect 583 1194 617 1226
rect 656 1194 690 1226
rect 729 1194 763 1226
rect 802 1194 836 1226
rect 875 1194 909 1226
rect 948 1194 982 1226
rect 1021 1194 1055 1226
rect 1094 1194 1128 1226
rect 1167 1194 1201 1226
rect 1240 1194 1274 1226
rect 1313 1194 1347 1226
rect 1386 1194 1420 1226
rect 1459 1194 1493 1226
rect 1532 1194 1566 1226
rect 1605 1194 1639 1226
rect 1678 1194 1712 1226
rect 1751 1194 1785 1226
rect 1824 1194 1858 1226
rect 1898 1194 1932 1226
rect 1972 1194 2006 1226
rect 2046 1194 2080 1226
rect 2120 1194 2154 1226
rect 2194 1194 2228 1226
rect 2268 1194 2302 1226
rect 2342 1194 2376 1226
rect 2416 1194 2450 1226
rect 2490 1194 2524 1226
rect 2564 1194 2574 1226
rect 2574 1194 2598 1226
rect 2638 1194 2643 1226
rect 2643 1194 2672 1226
rect 2712 1194 2746 1228
rect 2786 1226 2820 1228
rect 2860 1226 2894 1228
rect 2934 1226 2968 1228
rect 3008 1226 3042 1228
rect 3082 1226 3116 1228
rect 3156 1226 3190 1228
rect 3230 1226 3264 1228
rect 2786 1194 2816 1226
rect 2816 1194 2820 1226
rect 2860 1194 2885 1226
rect 2885 1194 2894 1226
rect 2934 1194 2954 1226
rect 2954 1194 2968 1226
rect 3008 1194 3023 1226
rect 3023 1194 3042 1226
rect 3082 1194 3092 1226
rect 3092 1194 3116 1226
rect 3156 1194 3161 1226
rect 3161 1194 3190 1226
rect 3230 1194 3264 1226
rect 364 1124 398 1156
rect 437 1124 471 1156
rect 510 1124 544 1156
rect 583 1124 617 1156
rect 656 1124 690 1156
rect 729 1124 763 1156
rect 802 1124 836 1156
rect 875 1124 909 1156
rect 948 1124 982 1156
rect 1021 1124 1055 1156
rect 1094 1124 1128 1156
rect 1167 1124 1201 1156
rect 1240 1124 1274 1156
rect 1313 1124 1347 1156
rect 1386 1124 1420 1156
rect 1459 1124 1493 1156
rect 1532 1124 1566 1156
rect 1605 1124 1639 1156
rect 1678 1124 1712 1156
rect 1751 1124 1785 1156
rect 1824 1124 1858 1156
rect 1898 1124 1932 1156
rect 1972 1124 2006 1156
rect 2046 1124 2080 1156
rect 2120 1124 2154 1156
rect 2194 1124 2228 1156
rect 2268 1124 2302 1156
rect 2342 1124 2376 1156
rect 2416 1124 2450 1156
rect 2490 1124 2524 1156
rect 2564 1124 2574 1156
rect 2574 1124 2598 1156
rect 2638 1124 2643 1156
rect 2643 1124 2672 1156
rect 364 1122 398 1124
rect 437 1122 471 1124
rect 510 1122 544 1124
rect 583 1122 617 1124
rect 656 1122 690 1124
rect 729 1122 763 1124
rect 802 1122 836 1124
rect 875 1122 909 1124
rect 948 1122 982 1124
rect 1021 1122 1055 1124
rect 1094 1122 1128 1124
rect 1167 1122 1201 1124
rect 1240 1122 1274 1124
rect 1313 1122 1347 1124
rect 1386 1122 1420 1124
rect 1459 1122 1493 1124
rect 1532 1122 1566 1124
rect 1605 1122 1639 1124
rect 1678 1122 1712 1124
rect 1751 1122 1785 1124
rect 1824 1122 1858 1124
rect 1898 1122 1932 1124
rect 1972 1122 2006 1124
rect 2046 1122 2080 1124
rect 2120 1122 2154 1124
rect 2194 1122 2228 1124
rect 2268 1122 2302 1124
rect 2342 1122 2376 1124
rect 2416 1122 2450 1124
rect 2490 1122 2524 1124
rect 2564 1122 2598 1124
rect 2638 1122 2672 1124
rect 2712 1122 2746 1156
rect 2786 1124 2816 1156
rect 2816 1124 2820 1156
rect 2860 1124 2885 1156
rect 2885 1124 2894 1156
rect 2934 1124 2954 1156
rect 2954 1124 2968 1156
rect 3008 1124 3023 1156
rect 3023 1124 3042 1156
rect 3082 1124 3092 1156
rect 3092 1124 3116 1156
rect 3156 1124 3161 1156
rect 3161 1124 3190 1156
rect 3230 1124 3264 1156
rect 2786 1122 2820 1124
rect 2860 1122 2894 1124
rect 2934 1122 2968 1124
rect 3008 1122 3042 1124
rect 3082 1122 3116 1124
rect 3156 1122 3190 1124
rect 3230 1122 3264 1124
rect 3606 1226 3640 1228
rect 3680 1226 3714 1228
rect 3754 1226 3788 1228
rect 3828 1226 3862 1228
rect 3902 1226 3936 1228
rect 3976 1226 4010 1228
rect 4050 1226 4084 1228
rect 3606 1194 3640 1226
rect 3680 1194 3709 1226
rect 3709 1194 3714 1226
rect 3754 1194 3778 1226
rect 3778 1194 3788 1226
rect 3828 1194 3847 1226
rect 3847 1194 3862 1226
rect 3902 1194 3916 1226
rect 3916 1194 3936 1226
rect 3976 1194 3985 1226
rect 3985 1194 4010 1226
rect 4050 1194 4054 1226
rect 4054 1194 4084 1226
rect 4124 1194 4158 1228
rect 4198 1226 4232 1228
rect 4272 1226 4306 1228
rect 4346 1226 4380 1228
rect 4420 1226 4454 1228
rect 4494 1226 4528 1228
rect 4568 1226 4602 1228
rect 4642 1226 4676 1228
rect 4716 1226 4750 1228
rect 4790 1226 4824 1228
rect 4864 1226 4898 1228
rect 4938 1226 4972 1228
rect 5012 1226 5046 1228
rect 5085 1226 5119 1228
rect 5158 1226 5192 1228
rect 5231 1226 5265 1228
rect 5304 1226 5338 1228
rect 5377 1226 5411 1228
rect 5450 1226 5484 1228
rect 5523 1226 5557 1228
rect 5596 1226 5630 1228
rect 5669 1226 5703 1228
rect 5742 1226 5776 1228
rect 5815 1226 5849 1228
rect 5888 1226 5922 1228
rect 5961 1226 5995 1228
rect 6034 1226 6068 1228
rect 6107 1226 6141 1228
rect 6180 1226 6214 1228
rect 6253 1226 6287 1228
rect 6326 1226 6360 1228
rect 6399 1226 6433 1228
rect 6472 1226 6506 1228
rect 4198 1194 4227 1226
rect 4227 1194 4232 1226
rect 4272 1194 4296 1226
rect 4296 1194 4306 1226
rect 4346 1194 4380 1226
rect 4420 1194 4454 1226
rect 4494 1194 4528 1226
rect 4568 1194 4602 1226
rect 4642 1194 4676 1226
rect 4716 1194 4750 1226
rect 4790 1194 4824 1226
rect 4864 1194 4898 1226
rect 4938 1194 4972 1226
rect 5012 1194 5046 1226
rect 5085 1194 5119 1226
rect 5158 1194 5192 1226
rect 5231 1194 5265 1226
rect 5304 1194 5338 1226
rect 5377 1194 5411 1226
rect 5450 1194 5484 1226
rect 5523 1194 5557 1226
rect 5596 1194 5630 1226
rect 5669 1194 5703 1226
rect 5742 1194 5776 1226
rect 5815 1194 5849 1226
rect 5888 1194 5922 1226
rect 5961 1194 5995 1226
rect 6034 1194 6068 1226
rect 6107 1194 6141 1226
rect 6180 1194 6214 1226
rect 6253 1194 6287 1226
rect 6326 1194 6360 1226
rect 6399 1194 6433 1226
rect 6472 1194 6506 1226
rect 3606 1124 3640 1156
rect 3680 1124 3709 1156
rect 3709 1124 3714 1156
rect 3754 1124 3778 1156
rect 3778 1124 3788 1156
rect 3828 1124 3847 1156
rect 3847 1124 3862 1156
rect 3902 1124 3916 1156
rect 3916 1124 3936 1156
rect 3976 1124 3985 1156
rect 3985 1124 4010 1156
rect 4050 1124 4054 1156
rect 4054 1124 4084 1156
rect 3606 1122 3640 1124
rect 3680 1122 3714 1124
rect 3754 1122 3788 1124
rect 3828 1122 3862 1124
rect 3902 1122 3936 1124
rect 3976 1122 4010 1124
rect 4050 1122 4084 1124
rect 4124 1122 4158 1156
rect 4198 1124 4227 1156
rect 4227 1124 4232 1156
rect 4272 1124 4296 1156
rect 4296 1124 4306 1156
rect 4346 1124 4380 1156
rect 4420 1124 4454 1156
rect 4494 1124 4528 1156
rect 4568 1124 4602 1156
rect 4642 1124 4676 1156
rect 4716 1124 4750 1156
rect 4790 1124 4824 1156
rect 4864 1124 4898 1156
rect 4938 1124 4972 1156
rect 5012 1124 5046 1156
rect 5085 1124 5119 1156
rect 5158 1124 5192 1156
rect 5231 1124 5265 1156
rect 5304 1124 5338 1156
rect 5377 1124 5411 1156
rect 5450 1124 5484 1156
rect 5523 1124 5557 1156
rect 5596 1124 5630 1156
rect 5669 1124 5703 1156
rect 5742 1124 5776 1156
rect 5815 1124 5849 1156
rect 5888 1124 5922 1156
rect 5961 1124 5995 1156
rect 6034 1124 6068 1156
rect 6107 1124 6141 1156
rect 6180 1124 6214 1156
rect 6253 1124 6287 1156
rect 6326 1124 6360 1156
rect 6399 1124 6433 1156
rect 6472 1124 6506 1156
rect 4198 1122 4232 1124
rect 4272 1122 4306 1124
rect 4346 1122 4380 1124
rect 4420 1122 4454 1124
rect 4494 1122 4528 1124
rect 4568 1122 4602 1124
rect 4642 1122 4676 1124
rect 4716 1122 4750 1124
rect 4790 1122 4824 1124
rect 4864 1122 4898 1124
rect 4938 1122 4972 1124
rect 5012 1122 5046 1124
rect 5085 1122 5119 1124
rect 5158 1122 5192 1124
rect 5231 1122 5265 1124
rect 5304 1122 5338 1124
rect 5377 1122 5411 1124
rect 5450 1122 5484 1124
rect 5523 1122 5557 1124
rect 5596 1122 5630 1124
rect 5669 1122 5703 1124
rect 5742 1122 5776 1124
rect 5815 1122 5849 1124
rect 5888 1122 5922 1124
rect 5961 1122 5995 1124
rect 6034 1122 6068 1124
rect 6107 1122 6141 1124
rect 6180 1122 6214 1124
rect 6253 1122 6287 1124
rect 6326 1122 6360 1124
rect 6399 1122 6433 1124
rect 6472 1122 6506 1124
rect 6848 1226 6882 1228
rect 6921 1226 6955 1228
rect 6994 1226 7028 1228
rect 7067 1226 7101 1228
rect 7140 1226 7174 1228
rect 7213 1226 7247 1228
rect 7286 1226 7320 1228
rect 7359 1226 7393 1228
rect 7432 1226 7466 1228
rect 7505 1226 7539 1228
rect 7578 1226 7612 1228
rect 7651 1226 7685 1228
rect 7724 1226 7758 1228
rect 7797 1226 7831 1228
rect 7870 1226 7904 1228
rect 7943 1226 7977 1228
rect 8016 1226 8050 1228
rect 8089 1226 8123 1228
rect 8162 1226 8196 1228
rect 8235 1226 8269 1228
rect 8308 1226 8342 1228
rect 8382 1226 8416 1228
rect 8456 1226 8490 1228
rect 8530 1226 8564 1228
rect 8604 1226 8638 1228
rect 8678 1226 8712 1228
rect 8752 1226 8786 1228
rect 8826 1226 8860 1228
rect 8900 1226 8934 1228
rect 8974 1226 9008 1228
rect 9048 1226 9082 1228
rect 9122 1226 9156 1228
rect 6848 1194 6882 1226
rect 6921 1194 6955 1226
rect 6994 1194 7028 1226
rect 7067 1194 7101 1226
rect 7140 1194 7174 1226
rect 7213 1194 7247 1226
rect 7286 1194 7320 1226
rect 7359 1194 7393 1226
rect 7432 1194 7466 1226
rect 7505 1194 7539 1226
rect 7578 1194 7612 1226
rect 7651 1194 7685 1226
rect 7724 1194 7758 1226
rect 7797 1194 7831 1226
rect 7870 1194 7904 1226
rect 7943 1194 7977 1226
rect 8016 1194 8050 1226
rect 8089 1194 8123 1226
rect 8162 1194 8196 1226
rect 8235 1194 8269 1226
rect 8308 1194 8342 1226
rect 8382 1194 8416 1226
rect 8456 1194 8490 1226
rect 8530 1194 8564 1226
rect 8604 1194 8638 1226
rect 8678 1194 8712 1226
rect 8752 1194 8786 1226
rect 8826 1194 8860 1226
rect 8900 1194 8934 1226
rect 8974 1194 9008 1226
rect 9048 1194 9058 1226
rect 9058 1194 9082 1226
rect 9122 1194 9127 1226
rect 9127 1194 9156 1226
rect 9196 1194 9230 1228
rect 9270 1226 9304 1228
rect 9344 1226 9378 1228
rect 9418 1226 9452 1228
rect 9492 1226 9526 1228
rect 9566 1226 9600 1228
rect 9640 1226 9674 1228
rect 9714 1226 9748 1228
rect 9270 1194 9300 1226
rect 9300 1194 9304 1226
rect 9344 1194 9369 1226
rect 9369 1194 9378 1226
rect 9418 1194 9438 1226
rect 9438 1194 9452 1226
rect 9492 1194 9507 1226
rect 9507 1194 9526 1226
rect 9566 1194 9576 1226
rect 9576 1194 9600 1226
rect 9640 1194 9645 1226
rect 9645 1194 9674 1226
rect 9714 1194 9748 1226
rect 6848 1124 6882 1156
rect 6921 1124 6955 1156
rect 6994 1124 7028 1156
rect 7067 1124 7101 1156
rect 7140 1124 7174 1156
rect 7213 1124 7247 1156
rect 7286 1124 7320 1156
rect 7359 1124 7393 1156
rect 7432 1124 7466 1156
rect 7505 1124 7539 1156
rect 7578 1124 7612 1156
rect 7651 1124 7685 1156
rect 7724 1124 7758 1156
rect 7797 1124 7831 1156
rect 7870 1124 7904 1156
rect 7943 1124 7977 1156
rect 8016 1124 8050 1156
rect 8089 1124 8123 1156
rect 8162 1124 8196 1156
rect 8235 1124 8269 1156
rect 8308 1124 8342 1156
rect 8382 1124 8416 1156
rect 8456 1124 8490 1156
rect 8530 1124 8564 1156
rect 8604 1124 8638 1156
rect 8678 1124 8712 1156
rect 8752 1124 8786 1156
rect 8826 1124 8860 1156
rect 8900 1124 8934 1156
rect 8974 1124 9008 1156
rect 9048 1124 9058 1156
rect 9058 1124 9082 1156
rect 9122 1124 9127 1156
rect 9127 1124 9156 1156
rect 6848 1122 6882 1124
rect 6921 1122 6955 1124
rect 6994 1122 7028 1124
rect 7067 1122 7101 1124
rect 7140 1122 7174 1124
rect 7213 1122 7247 1124
rect 7286 1122 7320 1124
rect 7359 1122 7393 1124
rect 7432 1122 7466 1124
rect 7505 1122 7539 1124
rect 7578 1122 7612 1124
rect 7651 1122 7685 1124
rect 7724 1122 7758 1124
rect 7797 1122 7831 1124
rect 7870 1122 7904 1124
rect 7943 1122 7977 1124
rect 8016 1122 8050 1124
rect 8089 1122 8123 1124
rect 8162 1122 8196 1124
rect 8235 1122 8269 1124
rect 8308 1122 8342 1124
rect 8382 1122 8416 1124
rect 8456 1122 8490 1124
rect 8530 1122 8564 1124
rect 8604 1122 8638 1124
rect 8678 1122 8712 1124
rect 8752 1122 8786 1124
rect 8826 1122 8860 1124
rect 8900 1122 8934 1124
rect 8974 1122 9008 1124
rect 9048 1122 9082 1124
rect 9122 1122 9156 1124
rect 9196 1122 9230 1156
rect 9270 1124 9300 1156
rect 9300 1124 9304 1156
rect 9344 1124 9369 1156
rect 9369 1124 9378 1156
rect 9418 1124 9438 1156
rect 9438 1124 9452 1156
rect 9492 1124 9507 1156
rect 9507 1124 9526 1156
rect 9566 1124 9576 1156
rect 9576 1124 9600 1156
rect 9640 1124 9645 1156
rect 9645 1124 9674 1156
rect 9714 1124 9748 1156
rect 9270 1122 9304 1124
rect 9344 1122 9378 1124
rect 9418 1122 9452 1124
rect 9492 1122 9526 1124
rect 9566 1122 9600 1124
rect 9640 1122 9674 1124
rect 9714 1122 9748 1124
rect 10090 1226 10124 1228
rect 10164 1226 10198 1228
rect 10238 1226 10272 1228
rect 10312 1226 10346 1228
rect 10386 1226 10420 1228
rect 10460 1226 10494 1228
rect 10534 1226 10568 1228
rect 10090 1194 10124 1226
rect 10164 1194 10193 1226
rect 10193 1194 10198 1226
rect 10238 1194 10262 1226
rect 10262 1194 10272 1226
rect 10312 1194 10331 1226
rect 10331 1194 10346 1226
rect 10386 1194 10400 1226
rect 10400 1194 10420 1226
rect 10460 1194 10469 1226
rect 10469 1194 10494 1226
rect 10534 1194 10538 1226
rect 10538 1194 10568 1226
rect 10608 1194 10642 1228
rect 10682 1226 10716 1228
rect 10756 1226 10790 1228
rect 10830 1226 10864 1228
rect 10904 1226 10938 1228
rect 10978 1226 11012 1228
rect 11052 1226 11086 1228
rect 11126 1226 11160 1228
rect 11200 1226 11234 1228
rect 11274 1226 11308 1228
rect 11348 1226 11382 1228
rect 11422 1226 11456 1228
rect 11496 1226 11530 1228
rect 11569 1226 11603 1228
rect 11642 1226 11676 1228
rect 11715 1226 11749 1228
rect 11788 1226 11822 1228
rect 11861 1226 11895 1228
rect 11934 1226 11968 1228
rect 12007 1226 12041 1228
rect 12080 1226 12114 1228
rect 12153 1226 12187 1228
rect 12226 1226 12260 1228
rect 12299 1226 12333 1228
rect 12372 1226 12406 1228
rect 12445 1226 12479 1228
rect 12518 1226 12552 1228
rect 12591 1226 12625 1228
rect 12664 1226 12698 1228
rect 12737 1226 12771 1228
rect 12810 1226 12844 1228
rect 12883 1226 12917 1228
rect 12956 1226 12990 1228
rect 10682 1194 10711 1226
rect 10711 1194 10716 1226
rect 10756 1194 10780 1226
rect 10780 1194 10790 1226
rect 10830 1194 10864 1226
rect 10904 1194 10938 1226
rect 10978 1194 11012 1226
rect 11052 1194 11086 1226
rect 11126 1194 11160 1226
rect 11200 1194 11234 1226
rect 11274 1194 11308 1226
rect 11348 1194 11382 1226
rect 11422 1194 11456 1226
rect 11496 1194 11530 1226
rect 11569 1194 11603 1226
rect 11642 1194 11676 1226
rect 11715 1194 11749 1226
rect 11788 1194 11822 1226
rect 11861 1194 11895 1226
rect 11934 1194 11968 1226
rect 12007 1194 12041 1226
rect 12080 1194 12114 1226
rect 12153 1194 12187 1226
rect 12226 1194 12260 1226
rect 12299 1194 12333 1226
rect 12372 1194 12406 1226
rect 12445 1194 12479 1226
rect 12518 1194 12552 1226
rect 12591 1194 12625 1226
rect 12664 1194 12698 1226
rect 12737 1194 12771 1226
rect 12810 1194 12844 1226
rect 12883 1194 12917 1226
rect 12956 1194 12990 1226
rect 10090 1124 10124 1156
rect 10164 1124 10193 1156
rect 10193 1124 10198 1156
rect 10238 1124 10262 1156
rect 10262 1124 10272 1156
rect 10312 1124 10331 1156
rect 10331 1124 10346 1156
rect 10386 1124 10400 1156
rect 10400 1124 10420 1156
rect 10460 1124 10469 1156
rect 10469 1124 10494 1156
rect 10534 1124 10538 1156
rect 10538 1124 10568 1156
rect 10090 1122 10124 1124
rect 10164 1122 10198 1124
rect 10238 1122 10272 1124
rect 10312 1122 10346 1124
rect 10386 1122 10420 1124
rect 10460 1122 10494 1124
rect 10534 1122 10568 1124
rect 10608 1122 10642 1156
rect 10682 1124 10711 1156
rect 10711 1124 10716 1156
rect 10756 1124 10780 1156
rect 10780 1124 10790 1156
rect 10830 1124 10864 1156
rect 10904 1124 10938 1156
rect 10978 1124 11012 1156
rect 11052 1124 11086 1156
rect 11126 1124 11160 1156
rect 11200 1124 11234 1156
rect 11274 1124 11308 1156
rect 11348 1124 11382 1156
rect 11422 1124 11456 1156
rect 11496 1124 11530 1156
rect 11569 1124 11603 1156
rect 11642 1124 11676 1156
rect 11715 1124 11749 1156
rect 11788 1124 11822 1156
rect 11861 1124 11895 1156
rect 11934 1124 11968 1156
rect 12007 1124 12041 1156
rect 12080 1124 12114 1156
rect 12153 1124 12187 1156
rect 12226 1124 12260 1156
rect 12299 1124 12333 1156
rect 12372 1124 12406 1156
rect 12445 1124 12479 1156
rect 12518 1124 12552 1156
rect 12591 1124 12625 1156
rect 12664 1124 12698 1156
rect 12737 1124 12771 1156
rect 12810 1124 12844 1156
rect 12883 1124 12917 1156
rect 12956 1124 12990 1156
rect 10682 1122 10716 1124
rect 10756 1122 10790 1124
rect 10830 1122 10864 1124
rect 10904 1122 10938 1124
rect 10978 1122 11012 1124
rect 11052 1122 11086 1124
rect 11126 1122 11160 1124
rect 11200 1122 11234 1124
rect 11274 1122 11308 1124
rect 11348 1122 11382 1124
rect 11422 1122 11456 1124
rect 11496 1122 11530 1124
rect 11569 1122 11603 1124
rect 11642 1122 11676 1124
rect 11715 1122 11749 1124
rect 11788 1122 11822 1124
rect 11861 1122 11895 1124
rect 11934 1122 11968 1124
rect 12007 1122 12041 1124
rect 12080 1122 12114 1124
rect 12153 1122 12187 1124
rect 12226 1122 12260 1124
rect 12299 1122 12333 1124
rect 12372 1122 12406 1124
rect 12445 1122 12479 1124
rect 12518 1122 12552 1124
rect 12591 1122 12625 1124
rect 12664 1122 12698 1124
rect 12737 1122 12771 1124
rect 12810 1122 12844 1124
rect 12883 1122 12917 1124
rect 12956 1122 12990 1124
rect 13332 1226 13366 1228
rect 13405 1226 13439 1228
rect 13478 1226 13512 1228
rect 13551 1226 13585 1228
rect 13624 1226 13658 1228
rect 13697 1226 13731 1228
rect 13770 1226 13804 1228
rect 13843 1226 13877 1228
rect 13916 1226 13950 1228
rect 13989 1226 14023 1228
rect 14062 1226 14096 1228
rect 14135 1226 14169 1228
rect 14208 1226 14242 1228
rect 14281 1226 14315 1228
rect 14354 1226 14388 1228
rect 14427 1226 14461 1228
rect 14500 1226 14534 1228
rect 14573 1226 14607 1228
rect 14646 1226 14680 1228
rect 14719 1226 14753 1228
rect 14792 1226 14826 1228
rect 14866 1226 14900 1228
rect 14940 1226 14974 1228
rect 15014 1226 15048 1228
rect 15088 1226 15122 1228
rect 15162 1226 15196 1228
rect 15236 1226 15270 1228
rect 15310 1226 15344 1228
rect 15384 1226 15418 1228
rect 15458 1226 15492 1228
rect 15532 1226 15566 1228
rect 15606 1226 15640 1228
rect 13332 1194 13366 1226
rect 13405 1194 13439 1226
rect 13478 1194 13512 1226
rect 13551 1194 13585 1226
rect 13624 1194 13658 1226
rect 13697 1194 13731 1226
rect 13770 1194 13804 1226
rect 13843 1194 13877 1226
rect 13916 1194 13950 1226
rect 13989 1194 14023 1226
rect 14062 1194 14096 1226
rect 14135 1194 14169 1226
rect 14208 1194 14242 1226
rect 14281 1194 14315 1226
rect 14354 1194 14388 1226
rect 14427 1194 14461 1226
rect 14500 1194 14534 1226
rect 14573 1194 14607 1226
rect 14646 1194 14680 1226
rect 14719 1194 14753 1226
rect 14792 1194 14826 1226
rect 14866 1194 14900 1226
rect 14940 1194 14974 1226
rect 15014 1194 15048 1226
rect 15088 1194 15122 1226
rect 15162 1194 15196 1226
rect 15236 1194 15270 1226
rect 15310 1194 15344 1226
rect 15384 1194 15418 1226
rect 15458 1194 15492 1226
rect 15532 1194 15542 1226
rect 15542 1194 15566 1226
rect 15606 1194 15611 1226
rect 15611 1194 15640 1226
rect 15680 1194 15714 1228
rect 15754 1226 15788 1228
rect 15828 1226 15862 1228
rect 15902 1226 15936 1228
rect 15976 1226 16010 1228
rect 16050 1226 16084 1228
rect 16124 1226 16158 1228
rect 16198 1226 16232 1228
rect 15754 1194 15784 1226
rect 15784 1194 15788 1226
rect 15828 1194 15853 1226
rect 15853 1194 15862 1226
rect 15902 1194 15922 1226
rect 15922 1194 15936 1226
rect 15976 1194 15991 1226
rect 15991 1194 16010 1226
rect 16050 1194 16060 1226
rect 16060 1194 16084 1226
rect 16124 1194 16129 1226
rect 16129 1194 16158 1226
rect 16198 1194 16232 1226
rect 13332 1124 13366 1156
rect 13405 1124 13439 1156
rect 13478 1124 13512 1156
rect 13551 1124 13585 1156
rect 13624 1124 13658 1156
rect 13697 1124 13731 1156
rect 13770 1124 13804 1156
rect 13843 1124 13877 1156
rect 13916 1124 13950 1156
rect 13989 1124 14023 1156
rect 14062 1124 14096 1156
rect 14135 1124 14169 1156
rect 14208 1124 14242 1156
rect 14281 1124 14315 1156
rect 14354 1124 14388 1156
rect 14427 1124 14461 1156
rect 14500 1124 14534 1156
rect 14573 1124 14607 1156
rect 14646 1124 14680 1156
rect 14719 1124 14753 1156
rect 14792 1124 14826 1156
rect 14866 1124 14900 1156
rect 14940 1124 14974 1156
rect 15014 1124 15048 1156
rect 15088 1124 15122 1156
rect 15162 1124 15196 1156
rect 15236 1124 15270 1156
rect 15310 1124 15344 1156
rect 15384 1124 15418 1156
rect 15458 1124 15492 1156
rect 15532 1124 15542 1156
rect 15542 1124 15566 1156
rect 15606 1124 15611 1156
rect 15611 1124 15640 1156
rect 13332 1122 13366 1124
rect 13405 1122 13439 1124
rect 13478 1122 13512 1124
rect 13551 1122 13585 1124
rect 13624 1122 13658 1124
rect 13697 1122 13731 1124
rect 13770 1122 13804 1124
rect 13843 1122 13877 1124
rect 13916 1122 13950 1124
rect 13989 1122 14023 1124
rect 14062 1122 14096 1124
rect 14135 1122 14169 1124
rect 14208 1122 14242 1124
rect 14281 1122 14315 1124
rect 14354 1122 14388 1124
rect 14427 1122 14461 1124
rect 14500 1122 14534 1124
rect 14573 1122 14607 1124
rect 14646 1122 14680 1124
rect 14719 1122 14753 1124
rect 14792 1122 14826 1124
rect 14866 1122 14900 1124
rect 14940 1122 14974 1124
rect 15014 1122 15048 1124
rect 15088 1122 15122 1124
rect 15162 1122 15196 1124
rect 15236 1122 15270 1124
rect 15310 1122 15344 1124
rect 15384 1122 15418 1124
rect 15458 1122 15492 1124
rect 15532 1122 15566 1124
rect 15606 1122 15640 1124
rect 15680 1122 15714 1156
rect 15754 1124 15784 1156
rect 15784 1124 15788 1156
rect 15828 1124 15853 1156
rect 15853 1124 15862 1156
rect 15902 1124 15922 1156
rect 15922 1124 15936 1156
rect 15976 1124 15991 1156
rect 15991 1124 16010 1156
rect 16050 1124 16060 1156
rect 16060 1124 16084 1156
rect 16124 1124 16129 1156
rect 16129 1124 16158 1156
rect 16198 1124 16232 1156
rect 15754 1122 15788 1124
rect 15828 1122 15862 1124
rect 15902 1122 15936 1124
rect 15976 1122 16010 1124
rect 16050 1122 16084 1124
rect 16124 1122 16158 1124
rect 16198 1122 16232 1124
rect 16574 1226 16608 1228
rect 16648 1226 16682 1228
rect 16722 1226 16756 1228
rect 16796 1226 16830 1228
rect 16870 1226 16904 1228
rect 16944 1226 16978 1228
rect 17018 1226 17052 1228
rect 16574 1194 16608 1226
rect 16648 1194 16677 1226
rect 16677 1194 16682 1226
rect 16722 1194 16746 1226
rect 16746 1194 16756 1226
rect 16796 1194 16815 1226
rect 16815 1194 16830 1226
rect 16870 1194 16884 1226
rect 16884 1194 16904 1226
rect 16944 1194 16953 1226
rect 16953 1194 16978 1226
rect 17018 1194 17022 1226
rect 17022 1194 17052 1226
rect 17092 1194 17126 1228
rect 17166 1226 17200 1228
rect 17240 1226 17274 1228
rect 17314 1226 17348 1228
rect 17388 1226 17422 1228
rect 17462 1226 17496 1228
rect 17536 1226 17570 1228
rect 17610 1226 17644 1228
rect 17684 1226 17718 1228
rect 17758 1226 17792 1228
rect 17832 1226 17866 1228
rect 17906 1226 17940 1228
rect 17980 1226 18014 1228
rect 18053 1226 18087 1228
rect 18126 1226 18160 1228
rect 18199 1226 18233 1228
rect 18272 1226 18306 1228
rect 18345 1226 18379 1228
rect 18418 1226 18452 1228
rect 18491 1226 18525 1228
rect 18564 1226 18598 1228
rect 18637 1226 18671 1228
rect 18710 1226 18744 1228
rect 18783 1226 18817 1228
rect 18856 1226 18890 1228
rect 18929 1226 18963 1228
rect 19002 1226 19036 1228
rect 19075 1226 19109 1228
rect 19148 1226 19182 1228
rect 19221 1226 19255 1228
rect 19294 1226 19328 1228
rect 19367 1226 19401 1228
rect 19440 1226 19474 1228
rect 17166 1194 17195 1226
rect 17195 1194 17200 1226
rect 17240 1194 17264 1226
rect 17264 1194 17274 1226
rect 17314 1194 17348 1226
rect 17388 1194 17422 1226
rect 17462 1194 17496 1226
rect 17536 1194 17570 1226
rect 17610 1194 17644 1226
rect 17684 1194 17718 1226
rect 17758 1194 17792 1226
rect 17832 1194 17866 1226
rect 17906 1194 17940 1226
rect 17980 1194 18014 1226
rect 18053 1194 18087 1226
rect 18126 1194 18160 1226
rect 18199 1194 18233 1226
rect 18272 1194 18306 1226
rect 18345 1194 18379 1226
rect 18418 1194 18452 1226
rect 18491 1194 18525 1226
rect 18564 1194 18598 1226
rect 18637 1194 18671 1226
rect 18710 1194 18744 1226
rect 18783 1194 18817 1226
rect 18856 1194 18890 1226
rect 18929 1194 18963 1226
rect 19002 1194 19036 1226
rect 19075 1194 19109 1226
rect 19148 1194 19182 1226
rect 19221 1194 19255 1226
rect 19294 1194 19328 1226
rect 19367 1194 19401 1226
rect 19440 1194 19474 1226
rect 16574 1124 16608 1156
rect 16648 1124 16677 1156
rect 16677 1124 16682 1156
rect 16722 1124 16746 1156
rect 16746 1124 16756 1156
rect 16796 1124 16815 1156
rect 16815 1124 16830 1156
rect 16870 1124 16884 1156
rect 16884 1124 16904 1156
rect 16944 1124 16953 1156
rect 16953 1124 16978 1156
rect 17018 1124 17022 1156
rect 17022 1124 17052 1156
rect 16574 1122 16608 1124
rect 16648 1122 16682 1124
rect 16722 1122 16756 1124
rect 16796 1122 16830 1124
rect 16870 1122 16904 1124
rect 16944 1122 16978 1124
rect 17018 1122 17052 1124
rect 17092 1122 17126 1156
rect 17166 1124 17195 1156
rect 17195 1124 17200 1156
rect 17240 1124 17264 1156
rect 17264 1124 17274 1156
rect 17314 1124 17348 1156
rect 17388 1124 17422 1156
rect 17462 1124 17496 1156
rect 17536 1124 17570 1156
rect 17610 1124 17644 1156
rect 17684 1124 17718 1156
rect 17758 1124 17792 1156
rect 17832 1124 17866 1156
rect 17906 1124 17940 1156
rect 17980 1124 18014 1156
rect 18053 1124 18087 1156
rect 18126 1124 18160 1156
rect 18199 1124 18233 1156
rect 18272 1124 18306 1156
rect 18345 1124 18379 1156
rect 18418 1124 18452 1156
rect 18491 1124 18525 1156
rect 18564 1124 18598 1156
rect 18637 1124 18671 1156
rect 18710 1124 18744 1156
rect 18783 1124 18817 1156
rect 18856 1124 18890 1156
rect 18929 1124 18963 1156
rect 19002 1124 19036 1156
rect 19075 1124 19109 1156
rect 19148 1124 19182 1156
rect 19221 1124 19255 1156
rect 19294 1124 19328 1156
rect 19367 1124 19401 1156
rect 19440 1124 19474 1156
rect 17166 1122 17200 1124
rect 17240 1122 17274 1124
rect 17314 1122 17348 1124
rect 17388 1122 17422 1124
rect 17462 1122 17496 1124
rect 17536 1122 17570 1124
rect 17610 1122 17644 1124
rect 17684 1122 17718 1124
rect 17758 1122 17792 1124
rect 17832 1122 17866 1124
rect 17906 1122 17940 1124
rect 17980 1122 18014 1124
rect 18053 1122 18087 1124
rect 18126 1122 18160 1124
rect 18199 1122 18233 1124
rect 18272 1122 18306 1124
rect 18345 1122 18379 1124
rect 18418 1122 18452 1124
rect 18491 1122 18525 1124
rect 18564 1122 18598 1124
rect 18637 1122 18671 1124
rect 18710 1122 18744 1124
rect 18783 1122 18817 1124
rect 18856 1122 18890 1124
rect 18929 1122 18963 1124
rect 19002 1122 19036 1124
rect 19075 1122 19109 1124
rect 19148 1122 19182 1124
rect 19221 1122 19255 1124
rect 19294 1122 19328 1124
rect 19367 1122 19401 1124
rect 19440 1122 19474 1124
rect 19882 1178 19916 1194
rect 19882 1160 19888 1178
rect 19888 1160 19916 1178
rect -46 1075 -12 1109
rect 42 1075 76 1109
rect -46 1001 -12 1035
rect 19882 1109 19916 1121
rect 19882 1087 19888 1109
rect 19888 1087 19916 1109
rect 42 1001 76 1035
rect -46 927 -12 961
rect 42 927 76 961
rect 168 918 182 938
rect 182 918 202 938
rect 168 904 202 918
rect 240 904 274 938
rect 3386 904 3420 938
rect 3458 904 3492 938
rect 6628 904 6662 938
rect 6700 904 6734 938
rect 9870 904 9904 938
rect 9942 904 9976 938
rect 13136 918 13150 938
rect 13150 918 13170 938
rect 13136 904 13170 918
rect 13208 904 13242 938
rect 19588 904 19622 938
rect 19882 1040 19916 1048
rect 19882 1014 19888 1040
rect 19888 1014 19916 1040
rect 19882 971 19916 975
rect 19882 941 19888 971
rect 19888 941 19916 971
rect 19660 904 19694 938
rect -46 853 -12 887
rect 42 853 76 887
rect -46 779 -12 813
rect 19882 868 19888 902
rect 19888 868 19916 902
rect 42 779 76 813
rect -46 705 -12 739
rect 42 705 76 739
rect 364 814 398 816
rect 437 814 471 816
rect 510 814 544 816
rect 583 814 617 816
rect 656 814 690 816
rect 729 814 763 816
rect 802 814 836 816
rect 875 814 909 816
rect 948 814 982 816
rect 1021 814 1055 816
rect 1094 814 1128 816
rect 1167 814 1201 816
rect 1240 814 1274 816
rect 1313 814 1347 816
rect 1386 814 1420 816
rect 1459 814 1493 816
rect 1532 814 1566 816
rect 1605 814 1639 816
rect 1678 814 1712 816
rect 1751 814 1785 816
rect 1824 814 1858 816
rect 1898 814 1932 816
rect 1972 814 2006 816
rect 2046 814 2080 816
rect 2120 814 2154 816
rect 2194 814 2228 816
rect 2268 814 2302 816
rect 2342 814 2376 816
rect 2416 814 2450 816
rect 2490 814 2524 816
rect 2564 814 2598 816
rect 2638 814 2672 816
rect 364 782 398 814
rect 437 782 471 814
rect 510 782 544 814
rect 583 782 617 814
rect 656 782 690 814
rect 729 782 763 814
rect 802 782 836 814
rect 875 782 909 814
rect 948 782 982 814
rect 1021 782 1055 814
rect 1094 782 1128 814
rect 1167 782 1201 814
rect 1240 782 1274 814
rect 1313 782 1347 814
rect 1386 782 1420 814
rect 1459 782 1493 814
rect 1532 782 1566 814
rect 1605 782 1639 814
rect 1678 782 1712 814
rect 1751 782 1785 814
rect 1824 782 1858 814
rect 1898 782 1932 814
rect 1972 782 2006 814
rect 2046 782 2080 814
rect 2120 782 2154 814
rect 2194 782 2228 814
rect 2268 782 2302 814
rect 2342 782 2376 814
rect 2416 782 2450 814
rect 2490 782 2524 814
rect 2564 782 2574 814
rect 2574 782 2598 814
rect 2638 782 2643 814
rect 2643 782 2672 814
rect 2712 782 2746 816
rect 2786 814 2820 816
rect 2860 814 2894 816
rect 2934 814 2968 816
rect 3008 814 3042 816
rect 3082 814 3116 816
rect 3156 814 3190 816
rect 3230 814 3264 816
rect 2786 782 2816 814
rect 2816 782 2820 814
rect 2860 782 2885 814
rect 2885 782 2894 814
rect 2934 782 2954 814
rect 2954 782 2968 814
rect 3008 782 3023 814
rect 3023 782 3042 814
rect 3082 782 3092 814
rect 3092 782 3116 814
rect 3156 782 3161 814
rect 3161 782 3190 814
rect 3230 782 3264 814
rect 364 712 398 744
rect 437 712 471 744
rect 510 712 544 744
rect 583 712 617 744
rect 656 712 690 744
rect 729 712 763 744
rect 802 712 836 744
rect 875 712 909 744
rect 948 712 982 744
rect 1021 712 1055 744
rect 1094 712 1128 744
rect 1167 712 1201 744
rect 1240 712 1274 744
rect 1313 712 1347 744
rect 1386 712 1420 744
rect 1459 712 1493 744
rect 1532 712 1566 744
rect 1605 712 1639 744
rect 1678 712 1712 744
rect 1751 712 1785 744
rect 1824 712 1858 744
rect 1898 712 1932 744
rect 1972 712 2006 744
rect 2046 712 2080 744
rect 2120 712 2154 744
rect 2194 712 2228 744
rect 2268 712 2302 744
rect 2342 712 2376 744
rect 2416 712 2450 744
rect 2490 712 2524 744
rect 2564 712 2574 744
rect 2574 712 2598 744
rect 2638 712 2643 744
rect 2643 712 2672 744
rect 364 710 398 712
rect 437 710 471 712
rect 510 710 544 712
rect 583 710 617 712
rect 656 710 690 712
rect 729 710 763 712
rect 802 710 836 712
rect 875 710 909 712
rect 948 710 982 712
rect 1021 710 1055 712
rect 1094 710 1128 712
rect 1167 710 1201 712
rect 1240 710 1274 712
rect 1313 710 1347 712
rect 1386 710 1420 712
rect 1459 710 1493 712
rect 1532 710 1566 712
rect 1605 710 1639 712
rect 1678 710 1712 712
rect 1751 710 1785 712
rect 1824 710 1858 712
rect 1898 710 1932 712
rect 1972 710 2006 712
rect 2046 710 2080 712
rect 2120 710 2154 712
rect 2194 710 2228 712
rect 2268 710 2302 712
rect 2342 710 2376 712
rect 2416 710 2450 712
rect 2490 710 2524 712
rect 2564 710 2598 712
rect 2638 710 2672 712
rect 2712 710 2746 744
rect 2786 712 2816 744
rect 2816 712 2820 744
rect 2860 712 2885 744
rect 2885 712 2894 744
rect 2934 712 2954 744
rect 2954 712 2968 744
rect 3008 712 3023 744
rect 3023 712 3042 744
rect 3082 712 3092 744
rect 3092 712 3116 744
rect 3156 712 3161 744
rect 3161 712 3190 744
rect 3230 712 3264 744
rect 2786 710 2820 712
rect 2860 710 2894 712
rect 2934 710 2968 712
rect 3008 710 3042 712
rect 3082 710 3116 712
rect 3156 710 3190 712
rect 3230 710 3264 712
rect 3606 814 3640 816
rect 3680 814 3714 816
rect 3754 814 3788 816
rect 3828 814 3862 816
rect 3902 814 3936 816
rect 3976 814 4010 816
rect 4050 814 4084 816
rect 3606 782 3640 814
rect 3680 782 3709 814
rect 3709 782 3714 814
rect 3754 782 3778 814
rect 3778 782 3788 814
rect 3828 782 3847 814
rect 3847 782 3862 814
rect 3902 782 3916 814
rect 3916 782 3936 814
rect 3976 782 3985 814
rect 3985 782 4010 814
rect 4050 782 4054 814
rect 4054 782 4084 814
rect 4124 782 4158 816
rect 4198 814 4232 816
rect 4272 814 4306 816
rect 4346 814 4380 816
rect 4420 814 4454 816
rect 4494 814 4528 816
rect 4568 814 4602 816
rect 4642 814 4676 816
rect 4716 814 4750 816
rect 4790 814 4824 816
rect 4864 814 4898 816
rect 4938 814 4972 816
rect 5012 814 5046 816
rect 5085 814 5119 816
rect 5158 814 5192 816
rect 5231 814 5265 816
rect 5304 814 5338 816
rect 5377 814 5411 816
rect 5450 814 5484 816
rect 5523 814 5557 816
rect 5596 814 5630 816
rect 5669 814 5703 816
rect 5742 814 5776 816
rect 5815 814 5849 816
rect 5888 814 5922 816
rect 5961 814 5995 816
rect 6034 814 6068 816
rect 6107 814 6141 816
rect 6180 814 6214 816
rect 6253 814 6287 816
rect 6326 814 6360 816
rect 6399 814 6433 816
rect 6472 814 6506 816
rect 4198 782 4227 814
rect 4227 782 4232 814
rect 4272 782 4296 814
rect 4296 782 4306 814
rect 4346 782 4380 814
rect 4420 782 4454 814
rect 4494 782 4528 814
rect 4568 782 4602 814
rect 4642 782 4676 814
rect 4716 782 4750 814
rect 4790 782 4824 814
rect 4864 782 4898 814
rect 4938 782 4972 814
rect 5012 782 5046 814
rect 5085 782 5119 814
rect 5158 782 5192 814
rect 5231 782 5265 814
rect 5304 782 5338 814
rect 5377 782 5411 814
rect 5450 782 5484 814
rect 5523 782 5557 814
rect 5596 782 5630 814
rect 5669 782 5703 814
rect 5742 782 5776 814
rect 5815 782 5849 814
rect 5888 782 5922 814
rect 5961 782 5995 814
rect 6034 782 6068 814
rect 6107 782 6141 814
rect 6180 782 6214 814
rect 6253 782 6287 814
rect 6326 782 6360 814
rect 6399 782 6433 814
rect 6472 782 6506 814
rect 3606 712 3640 744
rect 3680 712 3709 744
rect 3709 712 3714 744
rect 3754 712 3778 744
rect 3778 712 3788 744
rect 3828 712 3847 744
rect 3847 712 3862 744
rect 3902 712 3916 744
rect 3916 712 3936 744
rect 3976 712 3985 744
rect 3985 712 4010 744
rect 4050 712 4054 744
rect 4054 712 4084 744
rect 3606 710 3640 712
rect 3680 710 3714 712
rect 3754 710 3788 712
rect 3828 710 3862 712
rect 3902 710 3936 712
rect 3976 710 4010 712
rect 4050 710 4084 712
rect 4124 710 4158 744
rect 4198 712 4227 744
rect 4227 712 4232 744
rect 4272 712 4296 744
rect 4296 712 4306 744
rect 4346 712 4380 744
rect 4420 712 4454 744
rect 4494 712 4528 744
rect 4568 712 4602 744
rect 4642 712 4676 744
rect 4716 712 4750 744
rect 4790 712 4824 744
rect 4864 712 4898 744
rect 4938 712 4972 744
rect 5012 712 5046 744
rect 5085 712 5119 744
rect 5158 712 5192 744
rect 5231 712 5265 744
rect 5304 712 5338 744
rect 5377 712 5411 744
rect 5450 712 5484 744
rect 5523 712 5557 744
rect 5596 712 5630 744
rect 5669 712 5703 744
rect 5742 712 5776 744
rect 5815 712 5849 744
rect 5888 712 5922 744
rect 5961 712 5995 744
rect 6034 712 6068 744
rect 6107 712 6141 744
rect 6180 712 6214 744
rect 6253 712 6287 744
rect 6326 712 6360 744
rect 6399 712 6433 744
rect 6472 712 6506 744
rect 4198 710 4232 712
rect 4272 710 4306 712
rect 4346 710 4380 712
rect 4420 710 4454 712
rect 4494 710 4528 712
rect 4568 710 4602 712
rect 4642 710 4676 712
rect 4716 710 4750 712
rect 4790 710 4824 712
rect 4864 710 4898 712
rect 4938 710 4972 712
rect 5012 710 5046 712
rect 5085 710 5119 712
rect 5158 710 5192 712
rect 5231 710 5265 712
rect 5304 710 5338 712
rect 5377 710 5411 712
rect 5450 710 5484 712
rect 5523 710 5557 712
rect 5596 710 5630 712
rect 5669 710 5703 712
rect 5742 710 5776 712
rect 5815 710 5849 712
rect 5888 710 5922 712
rect 5961 710 5995 712
rect 6034 710 6068 712
rect 6107 710 6141 712
rect 6180 710 6214 712
rect 6253 710 6287 712
rect 6326 710 6360 712
rect 6399 710 6433 712
rect 6472 710 6506 712
rect 6848 814 6882 816
rect 6921 814 6955 816
rect 6994 814 7028 816
rect 7067 814 7101 816
rect 7140 814 7174 816
rect 7213 814 7247 816
rect 7286 814 7320 816
rect 7359 814 7393 816
rect 7432 814 7466 816
rect 7505 814 7539 816
rect 7578 814 7612 816
rect 7651 814 7685 816
rect 7724 814 7758 816
rect 7797 814 7831 816
rect 7870 814 7904 816
rect 7943 814 7977 816
rect 8016 814 8050 816
rect 8089 814 8123 816
rect 8162 814 8196 816
rect 8235 814 8269 816
rect 8308 814 8342 816
rect 8382 814 8416 816
rect 8456 814 8490 816
rect 8530 814 8564 816
rect 8604 814 8638 816
rect 8678 814 8712 816
rect 8752 814 8786 816
rect 8826 814 8860 816
rect 8900 814 8934 816
rect 8974 814 9008 816
rect 9048 814 9082 816
rect 9122 814 9156 816
rect 6848 782 6882 814
rect 6921 782 6955 814
rect 6994 782 7028 814
rect 7067 782 7101 814
rect 7140 782 7174 814
rect 7213 782 7247 814
rect 7286 782 7320 814
rect 7359 782 7393 814
rect 7432 782 7466 814
rect 7505 782 7539 814
rect 7578 782 7612 814
rect 7651 782 7685 814
rect 7724 782 7758 814
rect 7797 782 7831 814
rect 7870 782 7904 814
rect 7943 782 7977 814
rect 8016 782 8050 814
rect 8089 782 8123 814
rect 8162 782 8196 814
rect 8235 782 8269 814
rect 8308 782 8342 814
rect 8382 782 8416 814
rect 8456 782 8490 814
rect 8530 782 8564 814
rect 8604 782 8638 814
rect 8678 782 8712 814
rect 8752 782 8786 814
rect 8826 782 8860 814
rect 8900 782 8934 814
rect 8974 782 9008 814
rect 9048 782 9058 814
rect 9058 782 9082 814
rect 9122 782 9127 814
rect 9127 782 9156 814
rect 9196 782 9230 816
rect 9270 814 9304 816
rect 9344 814 9378 816
rect 9418 814 9452 816
rect 9492 814 9526 816
rect 9566 814 9600 816
rect 9640 814 9674 816
rect 9714 814 9748 816
rect 9270 782 9300 814
rect 9300 782 9304 814
rect 9344 782 9369 814
rect 9369 782 9378 814
rect 9418 782 9438 814
rect 9438 782 9452 814
rect 9492 782 9507 814
rect 9507 782 9526 814
rect 9566 782 9576 814
rect 9576 782 9600 814
rect 9640 782 9645 814
rect 9645 782 9674 814
rect 9714 782 9748 814
rect 6848 712 6882 744
rect 6921 712 6955 744
rect 6994 712 7028 744
rect 7067 712 7101 744
rect 7140 712 7174 744
rect 7213 712 7247 744
rect 7286 712 7320 744
rect 7359 712 7393 744
rect 7432 712 7466 744
rect 7505 712 7539 744
rect 7578 712 7612 744
rect 7651 712 7685 744
rect 7724 712 7758 744
rect 7797 712 7831 744
rect 7870 712 7904 744
rect 7943 712 7977 744
rect 8016 712 8050 744
rect 8089 712 8123 744
rect 8162 712 8196 744
rect 8235 712 8269 744
rect 8308 712 8342 744
rect 8382 712 8416 744
rect 8456 712 8490 744
rect 8530 712 8564 744
rect 8604 712 8638 744
rect 8678 712 8712 744
rect 8752 712 8786 744
rect 8826 712 8860 744
rect 8900 712 8934 744
rect 8974 712 9008 744
rect 9048 712 9058 744
rect 9058 712 9082 744
rect 9122 712 9127 744
rect 9127 712 9156 744
rect 6848 710 6882 712
rect 6921 710 6955 712
rect 6994 710 7028 712
rect 7067 710 7101 712
rect 7140 710 7174 712
rect 7213 710 7247 712
rect 7286 710 7320 712
rect 7359 710 7393 712
rect 7432 710 7466 712
rect 7505 710 7539 712
rect 7578 710 7612 712
rect 7651 710 7685 712
rect 7724 710 7758 712
rect 7797 710 7831 712
rect 7870 710 7904 712
rect 7943 710 7977 712
rect 8016 710 8050 712
rect 8089 710 8123 712
rect 8162 710 8196 712
rect 8235 710 8269 712
rect 8308 710 8342 712
rect 8382 710 8416 712
rect 8456 710 8490 712
rect 8530 710 8564 712
rect 8604 710 8638 712
rect 8678 710 8712 712
rect 8752 710 8786 712
rect 8826 710 8860 712
rect 8900 710 8934 712
rect 8974 710 9008 712
rect 9048 710 9082 712
rect 9122 710 9156 712
rect 9196 710 9230 744
rect 9270 712 9300 744
rect 9300 712 9304 744
rect 9344 712 9369 744
rect 9369 712 9378 744
rect 9418 712 9438 744
rect 9438 712 9452 744
rect 9492 712 9507 744
rect 9507 712 9526 744
rect 9566 712 9576 744
rect 9576 712 9600 744
rect 9640 712 9645 744
rect 9645 712 9674 744
rect 9714 712 9748 744
rect 9270 710 9304 712
rect 9344 710 9378 712
rect 9418 710 9452 712
rect 9492 710 9526 712
rect 9566 710 9600 712
rect 9640 710 9674 712
rect 9714 710 9748 712
rect 10090 814 10124 816
rect 10164 814 10198 816
rect 10238 814 10272 816
rect 10312 814 10346 816
rect 10386 814 10420 816
rect 10460 814 10494 816
rect 10534 814 10568 816
rect 10090 782 10124 814
rect 10164 782 10193 814
rect 10193 782 10198 814
rect 10238 782 10262 814
rect 10262 782 10272 814
rect 10312 782 10331 814
rect 10331 782 10346 814
rect 10386 782 10400 814
rect 10400 782 10420 814
rect 10460 782 10469 814
rect 10469 782 10494 814
rect 10534 782 10538 814
rect 10538 782 10568 814
rect 10608 782 10642 816
rect 10682 814 10716 816
rect 10756 814 10790 816
rect 10830 814 10864 816
rect 10904 814 10938 816
rect 10978 814 11012 816
rect 11052 814 11086 816
rect 11126 814 11160 816
rect 11200 814 11234 816
rect 11274 814 11308 816
rect 11348 814 11382 816
rect 11422 814 11456 816
rect 11496 814 11530 816
rect 11569 814 11603 816
rect 11642 814 11676 816
rect 11715 814 11749 816
rect 11788 814 11822 816
rect 11861 814 11895 816
rect 11934 814 11968 816
rect 12007 814 12041 816
rect 12080 814 12114 816
rect 12153 814 12187 816
rect 12226 814 12260 816
rect 12299 814 12333 816
rect 12372 814 12406 816
rect 12445 814 12479 816
rect 12518 814 12552 816
rect 12591 814 12625 816
rect 12664 814 12698 816
rect 12737 814 12771 816
rect 12810 814 12844 816
rect 12883 814 12917 816
rect 12956 814 12990 816
rect 10682 782 10711 814
rect 10711 782 10716 814
rect 10756 782 10780 814
rect 10780 782 10790 814
rect 10830 782 10864 814
rect 10904 782 10938 814
rect 10978 782 11012 814
rect 11052 782 11086 814
rect 11126 782 11160 814
rect 11200 782 11234 814
rect 11274 782 11308 814
rect 11348 782 11382 814
rect 11422 782 11456 814
rect 11496 782 11530 814
rect 11569 782 11603 814
rect 11642 782 11676 814
rect 11715 782 11749 814
rect 11788 782 11822 814
rect 11861 782 11895 814
rect 11934 782 11968 814
rect 12007 782 12041 814
rect 12080 782 12114 814
rect 12153 782 12187 814
rect 12226 782 12260 814
rect 12299 782 12333 814
rect 12372 782 12406 814
rect 12445 782 12479 814
rect 12518 782 12552 814
rect 12591 782 12625 814
rect 12664 782 12698 814
rect 12737 782 12771 814
rect 12810 782 12844 814
rect 12883 782 12917 814
rect 12956 782 12990 814
rect 10090 712 10124 744
rect 10164 712 10193 744
rect 10193 712 10198 744
rect 10238 712 10262 744
rect 10262 712 10272 744
rect 10312 712 10331 744
rect 10331 712 10346 744
rect 10386 712 10400 744
rect 10400 712 10420 744
rect 10460 712 10469 744
rect 10469 712 10494 744
rect 10534 712 10538 744
rect 10538 712 10568 744
rect 10090 710 10124 712
rect 10164 710 10198 712
rect 10238 710 10272 712
rect 10312 710 10346 712
rect 10386 710 10420 712
rect 10460 710 10494 712
rect 10534 710 10568 712
rect 10608 710 10642 744
rect 10682 712 10711 744
rect 10711 712 10716 744
rect 10756 712 10780 744
rect 10780 712 10790 744
rect 10830 712 10864 744
rect 10904 712 10938 744
rect 10978 712 11012 744
rect 11052 712 11086 744
rect 11126 712 11160 744
rect 11200 712 11234 744
rect 11274 712 11308 744
rect 11348 712 11382 744
rect 11422 712 11456 744
rect 11496 712 11530 744
rect 11569 712 11603 744
rect 11642 712 11676 744
rect 11715 712 11749 744
rect 11788 712 11822 744
rect 11861 712 11895 744
rect 11934 712 11968 744
rect 12007 712 12041 744
rect 12080 712 12114 744
rect 12153 712 12187 744
rect 12226 712 12260 744
rect 12299 712 12333 744
rect 12372 712 12406 744
rect 12445 712 12479 744
rect 12518 712 12552 744
rect 12591 712 12625 744
rect 12664 712 12698 744
rect 12737 712 12771 744
rect 12810 712 12844 744
rect 12883 712 12917 744
rect 12956 712 12990 744
rect 10682 710 10716 712
rect 10756 710 10790 712
rect 10830 710 10864 712
rect 10904 710 10938 712
rect 10978 710 11012 712
rect 11052 710 11086 712
rect 11126 710 11160 712
rect 11200 710 11234 712
rect 11274 710 11308 712
rect 11348 710 11382 712
rect 11422 710 11456 712
rect 11496 710 11530 712
rect 11569 710 11603 712
rect 11642 710 11676 712
rect 11715 710 11749 712
rect 11788 710 11822 712
rect 11861 710 11895 712
rect 11934 710 11968 712
rect 12007 710 12041 712
rect 12080 710 12114 712
rect 12153 710 12187 712
rect 12226 710 12260 712
rect 12299 710 12333 712
rect 12372 710 12406 712
rect 12445 710 12479 712
rect 12518 710 12552 712
rect 12591 710 12625 712
rect 12664 710 12698 712
rect 12737 710 12771 712
rect 12810 710 12844 712
rect 12883 710 12917 712
rect 12956 710 12990 712
rect 13332 814 13366 816
rect 13405 814 13439 816
rect 13478 814 13512 816
rect 13551 814 13585 816
rect 13624 814 13658 816
rect 13697 814 13731 816
rect 13770 814 13804 816
rect 13843 814 13877 816
rect 13916 814 13950 816
rect 13989 814 14023 816
rect 14062 814 14096 816
rect 14135 814 14169 816
rect 14208 814 14242 816
rect 14281 814 14315 816
rect 14354 814 14388 816
rect 14427 814 14461 816
rect 14500 814 14534 816
rect 14573 814 14607 816
rect 14646 814 14680 816
rect 14719 814 14753 816
rect 14792 814 14826 816
rect 14866 814 14900 816
rect 14940 814 14974 816
rect 15014 814 15048 816
rect 15088 814 15122 816
rect 15162 814 15196 816
rect 15236 814 15270 816
rect 15310 814 15344 816
rect 15384 814 15418 816
rect 15458 814 15492 816
rect 15532 814 15566 816
rect 15606 814 15640 816
rect 13332 782 13366 814
rect 13405 782 13439 814
rect 13478 782 13512 814
rect 13551 782 13585 814
rect 13624 782 13658 814
rect 13697 782 13731 814
rect 13770 782 13804 814
rect 13843 782 13877 814
rect 13916 782 13950 814
rect 13989 782 14023 814
rect 14062 782 14096 814
rect 14135 782 14169 814
rect 14208 782 14242 814
rect 14281 782 14315 814
rect 14354 782 14388 814
rect 14427 782 14461 814
rect 14500 782 14534 814
rect 14573 782 14607 814
rect 14646 782 14680 814
rect 14719 782 14753 814
rect 14792 782 14826 814
rect 14866 782 14900 814
rect 14940 782 14974 814
rect 15014 782 15048 814
rect 15088 782 15122 814
rect 15162 782 15196 814
rect 15236 782 15270 814
rect 15310 782 15344 814
rect 15384 782 15418 814
rect 15458 782 15492 814
rect 15532 782 15542 814
rect 15542 782 15566 814
rect 15606 782 15611 814
rect 15611 782 15640 814
rect 15680 782 15714 816
rect 15754 814 15788 816
rect 15828 814 15862 816
rect 15902 814 15936 816
rect 15976 814 16010 816
rect 16050 814 16084 816
rect 16124 814 16158 816
rect 16198 814 16232 816
rect 15754 782 15784 814
rect 15784 782 15788 814
rect 15828 782 15853 814
rect 15853 782 15862 814
rect 15902 782 15922 814
rect 15922 782 15936 814
rect 15976 782 15991 814
rect 15991 782 16010 814
rect 16050 782 16060 814
rect 16060 782 16084 814
rect 16124 782 16129 814
rect 16129 782 16158 814
rect 16198 782 16232 814
rect 13332 712 13366 744
rect 13405 712 13439 744
rect 13478 712 13512 744
rect 13551 712 13585 744
rect 13624 712 13658 744
rect 13697 712 13731 744
rect 13770 712 13804 744
rect 13843 712 13877 744
rect 13916 712 13950 744
rect 13989 712 14023 744
rect 14062 712 14096 744
rect 14135 712 14169 744
rect 14208 712 14242 744
rect 14281 712 14315 744
rect 14354 712 14388 744
rect 14427 712 14461 744
rect 14500 712 14534 744
rect 14573 712 14607 744
rect 14646 712 14680 744
rect 14719 712 14753 744
rect 14792 712 14826 744
rect 14866 712 14900 744
rect 14940 712 14974 744
rect 15014 712 15048 744
rect 15088 712 15122 744
rect 15162 712 15196 744
rect 15236 712 15270 744
rect 15310 712 15344 744
rect 15384 712 15418 744
rect 15458 712 15492 744
rect 15532 712 15542 744
rect 15542 712 15566 744
rect 15606 712 15611 744
rect 15611 712 15640 744
rect 13332 710 13366 712
rect 13405 710 13439 712
rect 13478 710 13512 712
rect 13551 710 13585 712
rect 13624 710 13658 712
rect 13697 710 13731 712
rect 13770 710 13804 712
rect 13843 710 13877 712
rect 13916 710 13950 712
rect 13989 710 14023 712
rect 14062 710 14096 712
rect 14135 710 14169 712
rect 14208 710 14242 712
rect 14281 710 14315 712
rect 14354 710 14388 712
rect 14427 710 14461 712
rect 14500 710 14534 712
rect 14573 710 14607 712
rect 14646 710 14680 712
rect 14719 710 14753 712
rect 14792 710 14826 712
rect 14866 710 14900 712
rect 14940 710 14974 712
rect 15014 710 15048 712
rect 15088 710 15122 712
rect 15162 710 15196 712
rect 15236 710 15270 712
rect 15310 710 15344 712
rect 15384 710 15418 712
rect 15458 710 15492 712
rect 15532 710 15566 712
rect 15606 710 15640 712
rect 15680 710 15714 744
rect 15754 712 15784 744
rect 15784 712 15788 744
rect 15828 712 15853 744
rect 15853 712 15862 744
rect 15902 712 15922 744
rect 15922 712 15936 744
rect 15976 712 15991 744
rect 15991 712 16010 744
rect 16050 712 16060 744
rect 16060 712 16084 744
rect 16124 712 16129 744
rect 16129 712 16158 744
rect 16198 712 16232 744
rect 15754 710 15788 712
rect 15828 710 15862 712
rect 15902 710 15936 712
rect 15976 710 16010 712
rect 16050 710 16084 712
rect 16124 710 16158 712
rect 16198 710 16232 712
rect 16574 814 16608 816
rect 16648 814 16682 816
rect 16722 814 16756 816
rect 16796 814 16830 816
rect 16870 814 16904 816
rect 16944 814 16978 816
rect 17018 814 17052 816
rect 16574 782 16608 814
rect 16648 782 16677 814
rect 16677 782 16682 814
rect 16722 782 16746 814
rect 16746 782 16756 814
rect 16796 782 16815 814
rect 16815 782 16830 814
rect 16870 782 16884 814
rect 16884 782 16904 814
rect 16944 782 16953 814
rect 16953 782 16978 814
rect 17018 782 17022 814
rect 17022 782 17052 814
rect 17092 782 17126 816
rect 17166 814 17200 816
rect 17240 814 17274 816
rect 17314 814 17348 816
rect 17388 814 17422 816
rect 17462 814 17496 816
rect 17536 814 17570 816
rect 17610 814 17644 816
rect 17684 814 17718 816
rect 17758 814 17792 816
rect 17832 814 17866 816
rect 17906 814 17940 816
rect 17980 814 18014 816
rect 18053 814 18087 816
rect 18126 814 18160 816
rect 18199 814 18233 816
rect 18272 814 18306 816
rect 18345 814 18379 816
rect 18418 814 18452 816
rect 18491 814 18525 816
rect 18564 814 18598 816
rect 18637 814 18671 816
rect 18710 814 18744 816
rect 18783 814 18817 816
rect 18856 814 18890 816
rect 18929 814 18963 816
rect 19002 814 19036 816
rect 19075 814 19109 816
rect 19148 814 19182 816
rect 19221 814 19255 816
rect 19294 814 19328 816
rect 19367 814 19401 816
rect 19440 814 19474 816
rect 17166 782 17195 814
rect 17195 782 17200 814
rect 17240 782 17264 814
rect 17264 782 17274 814
rect 17314 782 17348 814
rect 17388 782 17422 814
rect 17462 782 17496 814
rect 17536 782 17570 814
rect 17610 782 17644 814
rect 17684 782 17718 814
rect 17758 782 17792 814
rect 17832 782 17866 814
rect 17906 782 17940 814
rect 17980 782 18014 814
rect 18053 782 18087 814
rect 18126 782 18160 814
rect 18199 782 18233 814
rect 18272 782 18306 814
rect 18345 782 18379 814
rect 18418 782 18452 814
rect 18491 782 18525 814
rect 18564 782 18598 814
rect 18637 782 18671 814
rect 18710 782 18744 814
rect 18783 782 18817 814
rect 18856 782 18890 814
rect 18929 782 18963 814
rect 19002 782 19036 814
rect 19075 782 19109 814
rect 19148 782 19182 814
rect 19221 782 19255 814
rect 19294 782 19328 814
rect 19367 782 19401 814
rect 19440 782 19474 814
rect 16574 712 16608 744
rect 16648 712 16677 744
rect 16677 712 16682 744
rect 16722 712 16746 744
rect 16746 712 16756 744
rect 16796 712 16815 744
rect 16815 712 16830 744
rect 16870 712 16884 744
rect 16884 712 16904 744
rect 16944 712 16953 744
rect 16953 712 16978 744
rect 17018 712 17022 744
rect 17022 712 17052 744
rect 16574 710 16608 712
rect 16648 710 16682 712
rect 16722 710 16756 712
rect 16796 710 16830 712
rect 16870 710 16904 712
rect 16944 710 16978 712
rect 17018 710 17052 712
rect 17092 710 17126 744
rect 17166 712 17195 744
rect 17195 712 17200 744
rect 17240 712 17264 744
rect 17264 712 17274 744
rect 17314 712 17348 744
rect 17388 712 17422 744
rect 17462 712 17496 744
rect 17536 712 17570 744
rect 17610 712 17644 744
rect 17684 712 17718 744
rect 17758 712 17792 744
rect 17832 712 17866 744
rect 17906 712 17940 744
rect 17980 712 18014 744
rect 18053 712 18087 744
rect 18126 712 18160 744
rect 18199 712 18233 744
rect 18272 712 18306 744
rect 18345 712 18379 744
rect 18418 712 18452 744
rect 18491 712 18525 744
rect 18564 712 18598 744
rect 18637 712 18671 744
rect 18710 712 18744 744
rect 18783 712 18817 744
rect 18856 712 18890 744
rect 18929 712 18963 744
rect 19002 712 19036 744
rect 19075 712 19109 744
rect 19148 712 19182 744
rect 19221 712 19255 744
rect 19294 712 19328 744
rect 19367 712 19401 744
rect 19440 712 19474 744
rect 17166 710 17200 712
rect 17240 710 17274 712
rect 17314 710 17348 712
rect 17388 710 17422 712
rect 17462 710 17496 712
rect 17536 710 17570 712
rect 17610 710 17644 712
rect 17684 710 17718 712
rect 17758 710 17792 712
rect 17832 710 17866 712
rect 17906 710 17940 712
rect 17980 710 18014 712
rect 18053 710 18087 712
rect 18126 710 18160 712
rect 18199 710 18233 712
rect 18272 710 18306 712
rect 18345 710 18379 712
rect 18418 710 18452 712
rect 18491 710 18525 712
rect 18564 710 18598 712
rect 18637 710 18671 712
rect 18710 710 18744 712
rect 18783 710 18817 712
rect 18856 710 18890 712
rect 18929 710 18963 712
rect 19002 710 19036 712
rect 19075 710 19109 712
rect 19148 710 19182 712
rect 19221 710 19255 712
rect 19294 710 19328 712
rect 19367 710 19401 712
rect 19440 710 19474 712
rect 19882 799 19888 829
rect 19888 799 19916 829
rect 19882 795 19916 799
rect 19882 729 19888 756
rect 19888 729 19916 756
rect 19882 722 19916 729
rect -46 631 -12 665
rect 42 631 76 665
rect 19882 659 19888 683
rect 19888 659 19916 683
rect 19882 649 19916 659
rect -46 557 -12 591
rect 42 557 76 591
rect 144 588 178 622
rect -46 483 -12 517
rect 42 483 76 517
rect 216 588 250 622
rect 3386 588 3420 622
rect 3458 588 3492 622
rect 6628 588 6662 622
rect 6700 588 6734 622
rect 9870 588 9904 622
rect 9942 588 9976 622
rect 13112 588 13146 622
rect 13184 588 13218 622
rect 16354 588 16388 622
rect 16426 588 16460 622
rect 19564 588 19598 622
rect 19636 608 19670 622
rect 19636 588 19656 608
rect 19656 588 19670 608
rect 19882 589 19888 610
rect 19888 589 19916 610
rect 19882 576 19916 589
rect 19882 519 19888 537
rect 19888 519 19916 537
rect 19882 503 19916 519
rect -46 409 -12 443
rect 42 409 76 443
rect 19882 449 19888 465
rect 19888 449 19916 465
rect 19882 431 19916 449
rect -46 335 -12 369
rect 42 335 76 369
rect 364 402 398 404
rect 437 402 471 404
rect 510 402 544 404
rect 583 402 617 404
rect 656 402 690 404
rect 729 402 763 404
rect 802 402 836 404
rect 875 402 909 404
rect 948 402 982 404
rect 1021 402 1055 404
rect 1094 402 1128 404
rect 1167 402 1201 404
rect 1240 402 1274 404
rect 1313 402 1347 404
rect 1386 402 1420 404
rect 1459 402 1493 404
rect 1532 402 1566 404
rect 1605 402 1639 404
rect 1678 402 1712 404
rect 1751 402 1785 404
rect 1824 402 1858 404
rect 1898 402 1932 404
rect 1972 402 2006 404
rect 2046 402 2080 404
rect 2120 402 2154 404
rect 2194 402 2228 404
rect 2268 402 2302 404
rect 2342 402 2376 404
rect 2416 402 2450 404
rect 2490 402 2524 404
rect 2564 402 2598 404
rect 2638 402 2672 404
rect 364 370 398 402
rect 437 370 471 402
rect 510 370 544 402
rect 583 370 617 402
rect 656 370 690 402
rect 729 370 763 402
rect 802 370 836 402
rect 875 370 909 402
rect 948 370 982 402
rect 1021 370 1055 402
rect 1094 370 1128 402
rect 1167 370 1201 402
rect 1240 370 1274 402
rect 1313 370 1347 402
rect 1386 370 1420 402
rect 1459 370 1493 402
rect 1532 370 1566 402
rect 1605 370 1639 402
rect 1678 370 1712 402
rect 1751 370 1785 402
rect 1824 370 1858 402
rect 1898 370 1932 402
rect 1972 370 2006 402
rect 2046 370 2080 402
rect 2120 370 2154 402
rect 2194 370 2228 402
rect 2268 370 2302 402
rect 2342 370 2376 402
rect 2416 370 2450 402
rect 2490 370 2524 402
rect 2564 370 2574 402
rect 2574 370 2598 402
rect 2638 370 2643 402
rect 2643 370 2672 402
rect 2712 370 2746 404
rect 2786 402 2820 404
rect 2860 402 2894 404
rect 2934 402 2968 404
rect 3008 402 3042 404
rect 3082 402 3116 404
rect 3156 402 3190 404
rect 3230 402 3264 404
rect 2786 370 2816 402
rect 2816 370 2820 402
rect 2860 370 2885 402
rect 2885 370 2894 402
rect 2934 370 2954 402
rect 2954 370 2968 402
rect 3008 370 3023 402
rect 3023 370 3042 402
rect 3082 370 3092 402
rect 3092 370 3116 402
rect 3156 370 3161 402
rect 3161 370 3190 402
rect 3230 370 3264 402
rect 364 300 398 332
rect 437 300 471 332
rect 510 300 544 332
rect 583 300 617 332
rect 656 300 690 332
rect 729 300 763 332
rect 802 300 836 332
rect 875 300 909 332
rect 948 300 982 332
rect 1021 300 1055 332
rect 1094 300 1128 332
rect 1167 300 1201 332
rect 1240 300 1274 332
rect 1313 300 1347 332
rect 1386 300 1420 332
rect 1459 300 1493 332
rect 1532 300 1566 332
rect 1605 300 1639 332
rect 1678 300 1712 332
rect 1751 300 1785 332
rect 1824 300 1858 332
rect 1898 300 1932 332
rect 1972 300 2006 332
rect 2046 300 2080 332
rect 2120 300 2154 332
rect 2194 300 2228 332
rect 2268 300 2302 332
rect 2342 300 2376 332
rect 2416 300 2450 332
rect 2490 300 2524 332
rect 2564 300 2574 332
rect 2574 300 2598 332
rect 2638 300 2643 332
rect 2643 300 2672 332
rect 364 298 398 300
rect 437 298 471 300
rect 510 298 544 300
rect 583 298 617 300
rect 656 298 690 300
rect 729 298 763 300
rect 802 298 836 300
rect 875 298 909 300
rect 948 298 982 300
rect 1021 298 1055 300
rect 1094 298 1128 300
rect 1167 298 1201 300
rect 1240 298 1274 300
rect 1313 298 1347 300
rect 1386 298 1420 300
rect 1459 298 1493 300
rect 1532 298 1566 300
rect 1605 298 1639 300
rect 1678 298 1712 300
rect 1751 298 1785 300
rect 1824 298 1858 300
rect 1898 298 1932 300
rect 1972 298 2006 300
rect 2046 298 2080 300
rect 2120 298 2154 300
rect 2194 298 2228 300
rect 2268 298 2302 300
rect 2342 298 2376 300
rect 2416 298 2450 300
rect 2490 298 2524 300
rect 2564 298 2598 300
rect 2638 298 2672 300
rect 2712 298 2746 332
rect 2786 300 2816 332
rect 2816 300 2820 332
rect 2860 300 2885 332
rect 2885 300 2894 332
rect 2934 300 2954 332
rect 2954 300 2968 332
rect 3008 300 3023 332
rect 3023 300 3042 332
rect 3082 300 3092 332
rect 3092 300 3116 332
rect 3156 300 3161 332
rect 3161 300 3190 332
rect 3230 300 3264 332
rect 2786 298 2820 300
rect 2860 298 2894 300
rect 2934 298 2968 300
rect 3008 298 3042 300
rect 3082 298 3116 300
rect 3156 298 3190 300
rect 3230 298 3264 300
rect 3606 402 3640 404
rect 3680 402 3714 404
rect 3754 402 3788 404
rect 3828 402 3862 404
rect 3902 402 3936 404
rect 3976 402 4010 404
rect 4050 402 4084 404
rect 3606 370 3640 402
rect 3680 370 3709 402
rect 3709 370 3714 402
rect 3754 370 3778 402
rect 3778 370 3788 402
rect 3828 370 3847 402
rect 3847 370 3862 402
rect 3902 370 3916 402
rect 3916 370 3936 402
rect 3976 370 3985 402
rect 3985 370 4010 402
rect 4050 370 4054 402
rect 4054 370 4084 402
rect 4124 370 4158 404
rect 4198 402 4232 404
rect 4272 402 4306 404
rect 4346 402 4380 404
rect 4420 402 4454 404
rect 4494 402 4528 404
rect 4568 402 4602 404
rect 4642 402 4676 404
rect 4716 402 4750 404
rect 4790 402 4824 404
rect 4864 402 4898 404
rect 4938 402 4972 404
rect 5012 402 5046 404
rect 5085 402 5119 404
rect 5158 402 5192 404
rect 5231 402 5265 404
rect 5304 402 5338 404
rect 5377 402 5411 404
rect 5450 402 5484 404
rect 5523 402 5557 404
rect 5596 402 5630 404
rect 5669 402 5703 404
rect 5742 402 5776 404
rect 5815 402 5849 404
rect 5888 402 5922 404
rect 5961 402 5995 404
rect 6034 402 6068 404
rect 6107 402 6141 404
rect 6180 402 6214 404
rect 6253 402 6287 404
rect 6326 402 6360 404
rect 6399 402 6433 404
rect 6472 402 6506 404
rect 4198 370 4227 402
rect 4227 370 4232 402
rect 4272 370 4296 402
rect 4296 370 4306 402
rect 4346 370 4380 402
rect 4420 370 4454 402
rect 4494 370 4528 402
rect 4568 370 4602 402
rect 4642 370 4676 402
rect 4716 370 4750 402
rect 4790 370 4824 402
rect 4864 370 4898 402
rect 4938 370 4972 402
rect 5012 370 5046 402
rect 5085 370 5119 402
rect 5158 370 5192 402
rect 5231 370 5265 402
rect 5304 370 5338 402
rect 5377 370 5411 402
rect 5450 370 5484 402
rect 5523 370 5557 402
rect 5596 370 5630 402
rect 5669 370 5703 402
rect 5742 370 5776 402
rect 5815 370 5849 402
rect 5888 370 5922 402
rect 5961 370 5995 402
rect 6034 370 6068 402
rect 6107 370 6141 402
rect 6180 370 6214 402
rect 6253 370 6287 402
rect 6326 370 6360 402
rect 6399 370 6433 402
rect 6472 370 6506 402
rect 3606 300 3640 332
rect 3680 300 3709 332
rect 3709 300 3714 332
rect 3754 300 3778 332
rect 3778 300 3788 332
rect 3828 300 3847 332
rect 3847 300 3862 332
rect 3902 300 3916 332
rect 3916 300 3936 332
rect 3976 300 3985 332
rect 3985 300 4010 332
rect 4050 300 4054 332
rect 4054 300 4084 332
rect 3606 298 3640 300
rect 3680 298 3714 300
rect 3754 298 3788 300
rect 3828 298 3862 300
rect 3902 298 3936 300
rect 3976 298 4010 300
rect 4050 298 4084 300
rect 4124 298 4158 332
rect 4198 300 4227 332
rect 4227 300 4232 332
rect 4272 300 4296 332
rect 4296 300 4306 332
rect 4346 300 4380 332
rect 4420 300 4454 332
rect 4494 300 4528 332
rect 4568 300 4602 332
rect 4642 300 4676 332
rect 4716 300 4750 332
rect 4790 300 4824 332
rect 4864 300 4898 332
rect 4938 300 4972 332
rect 5012 300 5046 332
rect 5085 300 5119 332
rect 5158 300 5192 332
rect 5231 300 5265 332
rect 5304 300 5338 332
rect 5377 300 5411 332
rect 5450 300 5484 332
rect 5523 300 5557 332
rect 5596 300 5630 332
rect 5669 300 5703 332
rect 5742 300 5776 332
rect 5815 300 5849 332
rect 5888 300 5922 332
rect 5961 300 5995 332
rect 6034 300 6068 332
rect 6107 300 6141 332
rect 6180 300 6214 332
rect 6253 300 6287 332
rect 6326 300 6360 332
rect 6399 300 6433 332
rect 6472 300 6506 332
rect 4198 298 4232 300
rect 4272 298 4306 300
rect 4346 298 4380 300
rect 4420 298 4454 300
rect 4494 298 4528 300
rect 4568 298 4602 300
rect 4642 298 4676 300
rect 4716 298 4750 300
rect 4790 298 4824 300
rect 4864 298 4898 300
rect 4938 298 4972 300
rect 5012 298 5046 300
rect 5085 298 5119 300
rect 5158 298 5192 300
rect 5231 298 5265 300
rect 5304 298 5338 300
rect 5377 298 5411 300
rect 5450 298 5484 300
rect 5523 298 5557 300
rect 5596 298 5630 300
rect 5669 298 5703 300
rect 5742 298 5776 300
rect 5815 298 5849 300
rect 5888 298 5922 300
rect 5961 298 5995 300
rect 6034 298 6068 300
rect 6107 298 6141 300
rect 6180 298 6214 300
rect 6253 298 6287 300
rect 6326 298 6360 300
rect 6399 298 6433 300
rect 6472 298 6506 300
rect 6848 402 6882 404
rect 6921 402 6955 404
rect 6994 402 7028 404
rect 7067 402 7101 404
rect 7140 402 7174 404
rect 7213 402 7247 404
rect 7286 402 7320 404
rect 7359 402 7393 404
rect 7432 402 7466 404
rect 7505 402 7539 404
rect 7578 402 7612 404
rect 7651 402 7685 404
rect 7724 402 7758 404
rect 7797 402 7831 404
rect 7870 402 7904 404
rect 7943 402 7977 404
rect 8016 402 8050 404
rect 8089 402 8123 404
rect 8162 402 8196 404
rect 8235 402 8269 404
rect 8308 402 8342 404
rect 8382 402 8416 404
rect 8456 402 8490 404
rect 8530 402 8564 404
rect 8604 402 8638 404
rect 8678 402 8712 404
rect 8752 402 8786 404
rect 8826 402 8860 404
rect 8900 402 8934 404
rect 8974 402 9008 404
rect 9048 402 9082 404
rect 9122 402 9156 404
rect 6848 370 6882 402
rect 6921 370 6955 402
rect 6994 370 7028 402
rect 7067 370 7101 402
rect 7140 370 7174 402
rect 7213 370 7247 402
rect 7286 370 7320 402
rect 7359 370 7393 402
rect 7432 370 7466 402
rect 7505 370 7539 402
rect 7578 370 7612 402
rect 7651 370 7685 402
rect 7724 370 7758 402
rect 7797 370 7831 402
rect 7870 370 7904 402
rect 7943 370 7977 402
rect 8016 370 8050 402
rect 8089 370 8123 402
rect 8162 370 8196 402
rect 8235 370 8269 402
rect 8308 370 8342 402
rect 8382 370 8416 402
rect 8456 370 8490 402
rect 8530 370 8564 402
rect 8604 370 8638 402
rect 8678 370 8712 402
rect 8752 370 8786 402
rect 8826 370 8860 402
rect 8900 370 8934 402
rect 8974 370 9008 402
rect 9048 370 9058 402
rect 9058 370 9082 402
rect 9122 370 9127 402
rect 9127 370 9156 402
rect 9196 370 9230 404
rect 9270 402 9304 404
rect 9344 402 9378 404
rect 9418 402 9452 404
rect 9492 402 9526 404
rect 9566 402 9600 404
rect 9640 402 9674 404
rect 9714 402 9748 404
rect 9270 370 9300 402
rect 9300 370 9304 402
rect 9344 370 9369 402
rect 9369 370 9378 402
rect 9418 370 9438 402
rect 9438 370 9452 402
rect 9492 370 9507 402
rect 9507 370 9526 402
rect 9566 370 9576 402
rect 9576 370 9600 402
rect 9640 370 9645 402
rect 9645 370 9674 402
rect 9714 370 9748 402
rect 6848 300 6882 332
rect 6921 300 6955 332
rect 6994 300 7028 332
rect 7067 300 7101 332
rect 7140 300 7174 332
rect 7213 300 7247 332
rect 7286 300 7320 332
rect 7359 300 7393 332
rect 7432 300 7466 332
rect 7505 300 7539 332
rect 7578 300 7612 332
rect 7651 300 7685 332
rect 7724 300 7758 332
rect 7797 300 7831 332
rect 7870 300 7904 332
rect 7943 300 7977 332
rect 8016 300 8050 332
rect 8089 300 8123 332
rect 8162 300 8196 332
rect 8235 300 8269 332
rect 8308 300 8342 332
rect 8382 300 8416 332
rect 8456 300 8490 332
rect 8530 300 8564 332
rect 8604 300 8638 332
rect 8678 300 8712 332
rect 8752 300 8786 332
rect 8826 300 8860 332
rect 8900 300 8934 332
rect 8974 300 9008 332
rect 9048 300 9058 332
rect 9058 300 9082 332
rect 9122 300 9127 332
rect 9127 300 9156 332
rect 6848 298 6882 300
rect 6921 298 6955 300
rect 6994 298 7028 300
rect 7067 298 7101 300
rect 7140 298 7174 300
rect 7213 298 7247 300
rect 7286 298 7320 300
rect 7359 298 7393 300
rect 7432 298 7466 300
rect 7505 298 7539 300
rect 7578 298 7612 300
rect 7651 298 7685 300
rect 7724 298 7758 300
rect 7797 298 7831 300
rect 7870 298 7904 300
rect 7943 298 7977 300
rect 8016 298 8050 300
rect 8089 298 8123 300
rect 8162 298 8196 300
rect 8235 298 8269 300
rect 8308 298 8342 300
rect 8382 298 8416 300
rect 8456 298 8490 300
rect 8530 298 8564 300
rect 8604 298 8638 300
rect 8678 298 8712 300
rect 8752 298 8786 300
rect 8826 298 8860 300
rect 8900 298 8934 300
rect 8974 298 9008 300
rect 9048 298 9082 300
rect 9122 298 9156 300
rect 9196 298 9230 332
rect 9270 300 9300 332
rect 9300 300 9304 332
rect 9344 300 9369 332
rect 9369 300 9378 332
rect 9418 300 9438 332
rect 9438 300 9452 332
rect 9492 300 9507 332
rect 9507 300 9526 332
rect 9566 300 9576 332
rect 9576 300 9600 332
rect 9640 300 9645 332
rect 9645 300 9674 332
rect 9714 300 9748 332
rect 9270 298 9304 300
rect 9344 298 9378 300
rect 9418 298 9452 300
rect 9492 298 9526 300
rect 9566 298 9600 300
rect 9640 298 9674 300
rect 9714 298 9748 300
rect 10090 402 10124 404
rect 10164 402 10198 404
rect 10238 402 10272 404
rect 10312 402 10346 404
rect 10386 402 10420 404
rect 10460 402 10494 404
rect 10534 402 10568 404
rect 10090 370 10124 402
rect 10164 370 10193 402
rect 10193 370 10198 402
rect 10238 370 10262 402
rect 10262 370 10272 402
rect 10312 370 10331 402
rect 10331 370 10346 402
rect 10386 370 10400 402
rect 10400 370 10420 402
rect 10460 370 10469 402
rect 10469 370 10494 402
rect 10534 370 10538 402
rect 10538 370 10568 402
rect 10608 370 10642 404
rect 10682 402 10716 404
rect 10756 402 10790 404
rect 10830 402 10864 404
rect 10904 402 10938 404
rect 10978 402 11012 404
rect 11052 402 11086 404
rect 11126 402 11160 404
rect 11200 402 11234 404
rect 11274 402 11308 404
rect 11348 402 11382 404
rect 11422 402 11456 404
rect 11496 402 11530 404
rect 11569 402 11603 404
rect 11642 402 11676 404
rect 11715 402 11749 404
rect 11788 402 11822 404
rect 11861 402 11895 404
rect 11934 402 11968 404
rect 12007 402 12041 404
rect 12080 402 12114 404
rect 12153 402 12187 404
rect 12226 402 12260 404
rect 12299 402 12333 404
rect 12372 402 12406 404
rect 12445 402 12479 404
rect 12518 402 12552 404
rect 12591 402 12625 404
rect 12664 402 12698 404
rect 12737 402 12771 404
rect 12810 402 12844 404
rect 12883 402 12917 404
rect 12956 402 12990 404
rect 10682 370 10711 402
rect 10711 370 10716 402
rect 10756 370 10780 402
rect 10780 370 10790 402
rect 10830 370 10864 402
rect 10904 370 10938 402
rect 10978 370 11012 402
rect 11052 370 11086 402
rect 11126 370 11160 402
rect 11200 370 11234 402
rect 11274 370 11308 402
rect 11348 370 11382 402
rect 11422 370 11456 402
rect 11496 370 11530 402
rect 11569 370 11603 402
rect 11642 370 11676 402
rect 11715 370 11749 402
rect 11788 370 11822 402
rect 11861 370 11895 402
rect 11934 370 11968 402
rect 12007 370 12041 402
rect 12080 370 12114 402
rect 12153 370 12187 402
rect 12226 370 12260 402
rect 12299 370 12333 402
rect 12372 370 12406 402
rect 12445 370 12479 402
rect 12518 370 12552 402
rect 12591 370 12625 402
rect 12664 370 12698 402
rect 12737 370 12771 402
rect 12810 370 12844 402
rect 12883 370 12917 402
rect 12956 370 12990 402
rect 10090 300 10124 332
rect 10164 300 10193 332
rect 10193 300 10198 332
rect 10238 300 10262 332
rect 10262 300 10272 332
rect 10312 300 10331 332
rect 10331 300 10346 332
rect 10386 300 10400 332
rect 10400 300 10420 332
rect 10460 300 10469 332
rect 10469 300 10494 332
rect 10534 300 10538 332
rect 10538 300 10568 332
rect 10090 298 10124 300
rect 10164 298 10198 300
rect 10238 298 10272 300
rect 10312 298 10346 300
rect 10386 298 10420 300
rect 10460 298 10494 300
rect 10534 298 10568 300
rect 10608 298 10642 332
rect 10682 300 10711 332
rect 10711 300 10716 332
rect 10756 300 10780 332
rect 10780 300 10790 332
rect 10830 300 10864 332
rect 10904 300 10938 332
rect 10978 300 11012 332
rect 11052 300 11086 332
rect 11126 300 11160 332
rect 11200 300 11234 332
rect 11274 300 11308 332
rect 11348 300 11382 332
rect 11422 300 11456 332
rect 11496 300 11530 332
rect 11569 300 11603 332
rect 11642 300 11676 332
rect 11715 300 11749 332
rect 11788 300 11822 332
rect 11861 300 11895 332
rect 11934 300 11968 332
rect 12007 300 12041 332
rect 12080 300 12114 332
rect 12153 300 12187 332
rect 12226 300 12260 332
rect 12299 300 12333 332
rect 12372 300 12406 332
rect 12445 300 12479 332
rect 12518 300 12552 332
rect 12591 300 12625 332
rect 12664 300 12698 332
rect 12737 300 12771 332
rect 12810 300 12844 332
rect 12883 300 12917 332
rect 12956 300 12990 332
rect 10682 298 10716 300
rect 10756 298 10790 300
rect 10830 298 10864 300
rect 10904 298 10938 300
rect 10978 298 11012 300
rect 11052 298 11086 300
rect 11126 298 11160 300
rect 11200 298 11234 300
rect 11274 298 11308 300
rect 11348 298 11382 300
rect 11422 298 11456 300
rect 11496 298 11530 300
rect 11569 298 11603 300
rect 11642 298 11676 300
rect 11715 298 11749 300
rect 11788 298 11822 300
rect 11861 298 11895 300
rect 11934 298 11968 300
rect 12007 298 12041 300
rect 12080 298 12114 300
rect 12153 298 12187 300
rect 12226 298 12260 300
rect 12299 298 12333 300
rect 12372 298 12406 300
rect 12445 298 12479 300
rect 12518 298 12552 300
rect 12591 298 12625 300
rect 12664 298 12698 300
rect 12737 298 12771 300
rect 12810 298 12844 300
rect 12883 298 12917 300
rect 12956 298 12990 300
rect 13332 402 13366 404
rect 13405 402 13439 404
rect 13478 402 13512 404
rect 13551 402 13585 404
rect 13624 402 13658 404
rect 13697 402 13731 404
rect 13770 402 13804 404
rect 13843 402 13877 404
rect 13916 402 13950 404
rect 13989 402 14023 404
rect 14062 402 14096 404
rect 14135 402 14169 404
rect 14208 402 14242 404
rect 14281 402 14315 404
rect 14354 402 14388 404
rect 14427 402 14461 404
rect 14500 402 14534 404
rect 14573 402 14607 404
rect 14646 402 14680 404
rect 14719 402 14753 404
rect 14792 402 14826 404
rect 14866 402 14900 404
rect 14940 402 14974 404
rect 15014 402 15048 404
rect 15088 402 15122 404
rect 15162 402 15196 404
rect 15236 402 15270 404
rect 15310 402 15344 404
rect 15384 402 15418 404
rect 15458 402 15492 404
rect 15532 402 15566 404
rect 15606 402 15640 404
rect 13332 370 13366 402
rect 13405 370 13439 402
rect 13478 370 13512 402
rect 13551 370 13585 402
rect 13624 370 13658 402
rect 13697 370 13731 402
rect 13770 370 13804 402
rect 13843 370 13877 402
rect 13916 370 13950 402
rect 13989 370 14023 402
rect 14062 370 14096 402
rect 14135 370 14169 402
rect 14208 370 14242 402
rect 14281 370 14315 402
rect 14354 370 14388 402
rect 14427 370 14461 402
rect 14500 370 14534 402
rect 14573 370 14607 402
rect 14646 370 14680 402
rect 14719 370 14753 402
rect 14792 370 14826 402
rect 14866 370 14900 402
rect 14940 370 14974 402
rect 15014 370 15048 402
rect 15088 370 15122 402
rect 15162 370 15196 402
rect 15236 370 15270 402
rect 15310 370 15344 402
rect 15384 370 15418 402
rect 15458 370 15492 402
rect 15532 370 15542 402
rect 15542 370 15566 402
rect 15606 370 15611 402
rect 15611 370 15640 402
rect 15680 370 15714 404
rect 15754 402 15788 404
rect 15828 402 15862 404
rect 15902 402 15936 404
rect 15976 402 16010 404
rect 16050 402 16084 404
rect 16124 402 16158 404
rect 16198 402 16232 404
rect 15754 370 15784 402
rect 15784 370 15788 402
rect 15828 370 15853 402
rect 15853 370 15862 402
rect 15902 370 15922 402
rect 15922 370 15936 402
rect 15976 370 15991 402
rect 15991 370 16010 402
rect 16050 370 16060 402
rect 16060 370 16084 402
rect 16124 370 16129 402
rect 16129 370 16158 402
rect 16198 370 16232 402
rect 13332 300 13366 332
rect 13405 300 13439 332
rect 13478 300 13512 332
rect 13551 300 13585 332
rect 13624 300 13658 332
rect 13697 300 13731 332
rect 13770 300 13804 332
rect 13843 300 13877 332
rect 13916 300 13950 332
rect 13989 300 14023 332
rect 14062 300 14096 332
rect 14135 300 14169 332
rect 14208 300 14242 332
rect 14281 300 14315 332
rect 14354 300 14388 332
rect 14427 300 14461 332
rect 14500 300 14534 332
rect 14573 300 14607 332
rect 14646 300 14680 332
rect 14719 300 14753 332
rect 14792 300 14826 332
rect 14866 300 14900 332
rect 14940 300 14974 332
rect 15014 300 15048 332
rect 15088 300 15122 332
rect 15162 300 15196 332
rect 15236 300 15270 332
rect 15310 300 15344 332
rect 15384 300 15418 332
rect 15458 300 15492 332
rect 15532 300 15542 332
rect 15542 300 15566 332
rect 15606 300 15611 332
rect 15611 300 15640 332
rect 13332 298 13366 300
rect 13405 298 13439 300
rect 13478 298 13512 300
rect 13551 298 13585 300
rect 13624 298 13658 300
rect 13697 298 13731 300
rect 13770 298 13804 300
rect 13843 298 13877 300
rect 13916 298 13950 300
rect 13989 298 14023 300
rect 14062 298 14096 300
rect 14135 298 14169 300
rect 14208 298 14242 300
rect 14281 298 14315 300
rect 14354 298 14388 300
rect 14427 298 14461 300
rect 14500 298 14534 300
rect 14573 298 14607 300
rect 14646 298 14680 300
rect 14719 298 14753 300
rect 14792 298 14826 300
rect 14866 298 14900 300
rect 14940 298 14974 300
rect 15014 298 15048 300
rect 15088 298 15122 300
rect 15162 298 15196 300
rect 15236 298 15270 300
rect 15310 298 15344 300
rect 15384 298 15418 300
rect 15458 298 15492 300
rect 15532 298 15566 300
rect 15606 298 15640 300
rect 15680 298 15714 332
rect 15754 300 15784 332
rect 15784 300 15788 332
rect 15828 300 15853 332
rect 15853 300 15862 332
rect 15902 300 15922 332
rect 15922 300 15936 332
rect 15976 300 15991 332
rect 15991 300 16010 332
rect 16050 300 16060 332
rect 16060 300 16084 332
rect 16124 300 16129 332
rect 16129 300 16158 332
rect 16198 300 16232 332
rect 15754 298 15788 300
rect 15828 298 15862 300
rect 15902 298 15936 300
rect 15976 298 16010 300
rect 16050 298 16084 300
rect 16124 298 16158 300
rect 16198 298 16232 300
rect 16574 402 16608 404
rect 16648 402 16682 404
rect 16722 402 16756 404
rect 16796 402 16830 404
rect 16870 402 16904 404
rect 16944 402 16978 404
rect 17018 402 17052 404
rect 16574 370 16608 402
rect 16648 370 16677 402
rect 16677 370 16682 402
rect 16722 370 16746 402
rect 16746 370 16756 402
rect 16796 370 16815 402
rect 16815 370 16830 402
rect 16870 370 16884 402
rect 16884 370 16904 402
rect 16944 370 16953 402
rect 16953 370 16978 402
rect 17018 370 17022 402
rect 17022 370 17052 402
rect 17092 370 17126 404
rect 17166 402 17200 404
rect 17240 402 17274 404
rect 17314 402 17348 404
rect 17388 402 17422 404
rect 17462 402 17496 404
rect 17536 402 17570 404
rect 17610 402 17644 404
rect 17684 402 17718 404
rect 17758 402 17792 404
rect 17832 402 17866 404
rect 17906 402 17940 404
rect 17980 402 18014 404
rect 18053 402 18087 404
rect 18126 402 18160 404
rect 18199 402 18233 404
rect 18272 402 18306 404
rect 18345 402 18379 404
rect 18418 402 18452 404
rect 18491 402 18525 404
rect 18564 402 18598 404
rect 18637 402 18671 404
rect 18710 402 18744 404
rect 18783 402 18817 404
rect 18856 402 18890 404
rect 18929 402 18963 404
rect 19002 402 19036 404
rect 19075 402 19109 404
rect 19148 402 19182 404
rect 19221 402 19255 404
rect 19294 402 19328 404
rect 19367 402 19401 404
rect 19440 402 19474 404
rect 17166 370 17195 402
rect 17195 370 17200 402
rect 17240 370 17264 402
rect 17264 370 17274 402
rect 17314 370 17348 402
rect 17388 370 17422 402
rect 17462 370 17496 402
rect 17536 370 17570 402
rect 17610 370 17644 402
rect 17684 370 17718 402
rect 17758 370 17792 402
rect 17832 370 17866 402
rect 17906 370 17940 402
rect 17980 370 18014 402
rect 18053 370 18087 402
rect 18126 370 18160 402
rect 18199 370 18233 402
rect 18272 370 18306 402
rect 18345 370 18379 402
rect 18418 370 18452 402
rect 18491 370 18525 402
rect 18564 370 18598 402
rect 18637 370 18671 402
rect 18710 370 18744 402
rect 18783 370 18817 402
rect 18856 370 18890 402
rect 18929 370 18963 402
rect 19002 370 19036 402
rect 19075 370 19109 402
rect 19148 370 19182 402
rect 19221 370 19255 402
rect 19294 370 19328 402
rect 19367 370 19401 402
rect 19440 370 19474 402
rect 16574 300 16608 332
rect 16648 300 16677 332
rect 16677 300 16682 332
rect 16722 300 16746 332
rect 16746 300 16756 332
rect 16796 300 16815 332
rect 16815 300 16830 332
rect 16870 300 16884 332
rect 16884 300 16904 332
rect 16944 300 16953 332
rect 16953 300 16978 332
rect 17018 300 17022 332
rect 17022 300 17052 332
rect 16574 298 16608 300
rect 16648 298 16682 300
rect 16722 298 16756 300
rect 16796 298 16830 300
rect 16870 298 16904 300
rect 16944 298 16978 300
rect 17018 298 17052 300
rect 17092 298 17126 332
rect 17166 300 17195 332
rect 17195 300 17200 332
rect 17240 300 17264 332
rect 17264 300 17274 332
rect 17314 300 17348 332
rect 17388 300 17422 332
rect 17462 300 17496 332
rect 17536 300 17570 332
rect 17610 300 17644 332
rect 17684 300 17718 332
rect 17758 300 17792 332
rect 17832 300 17866 332
rect 17906 300 17940 332
rect 17980 300 18014 332
rect 18053 300 18087 332
rect 18126 300 18160 332
rect 18199 300 18233 332
rect 18272 300 18306 332
rect 18345 300 18379 332
rect 18418 300 18452 332
rect 18491 300 18525 332
rect 18564 300 18598 332
rect 18637 300 18671 332
rect 18710 300 18744 332
rect 18783 300 18817 332
rect 18856 300 18890 332
rect 18929 300 18963 332
rect 19002 300 19036 332
rect 19075 300 19109 332
rect 19148 300 19182 332
rect 19221 300 19255 332
rect 19294 300 19328 332
rect 19367 300 19401 332
rect 19440 300 19474 332
rect 17166 298 17200 300
rect 17240 298 17274 300
rect 17314 298 17348 300
rect 17388 298 17422 300
rect 17462 298 17496 300
rect 17536 298 17570 300
rect 17610 298 17644 300
rect 17684 298 17718 300
rect 17758 298 17792 300
rect 17832 298 17866 300
rect 17906 298 17940 300
rect 17980 298 18014 300
rect 18053 298 18087 300
rect 18126 298 18160 300
rect 18199 298 18233 300
rect 18272 298 18306 300
rect 18345 298 18379 300
rect 18418 298 18452 300
rect 18491 298 18525 300
rect 18564 298 18598 300
rect 18637 298 18671 300
rect 18710 298 18744 300
rect 18783 298 18817 300
rect 18856 298 18890 300
rect 18929 298 18963 300
rect 19002 298 19036 300
rect 19075 298 19109 300
rect 19148 298 19182 300
rect 19221 298 19255 300
rect 19294 298 19328 300
rect 19367 298 19401 300
rect 19440 298 19474 300
rect 19882 379 19888 393
rect 19888 379 19916 393
rect 19882 359 19916 379
rect -46 261 -12 295
rect 42 261 76 295
rect -46 187 -12 221
rect 42 187 76 221
rect 19882 309 19888 321
rect 19888 309 19916 321
rect 19882 287 19916 309
rect 19882 239 19888 249
rect 19888 239 19916 249
rect 19882 215 19916 239
rect -46 113 -12 147
rect 42 113 76 147
rect 168 94 182 114
rect 182 94 202 114
rect 168 80 202 94
rect 240 80 274 114
rect 3386 80 3420 114
rect 3458 80 3492 114
rect 9870 80 9904 114
rect 9942 80 9976 114
rect 16354 80 16388 114
rect 16426 80 16460 114
rect 19588 80 19622 114
rect 19882 169 19888 177
rect 19888 169 19916 177
rect 19882 143 19916 169
rect 19660 80 19694 114
rect -46 39 -12 73
rect 42 39 76 73
rect -46 -35 -12 -1
rect 42 -35 76 -1
rect 19882 99 19888 105
rect 19888 99 19916 105
rect 19882 71 19916 99
rect 19882 29 19888 33
rect 19888 29 19916 33
rect 19882 -1 19916 29
rect -46 -109 -12 -75
rect 42 -109 76 -75
rect 364 -10 398 -8
rect 437 -10 471 -8
rect 510 -10 544 -8
rect 583 -10 617 -8
rect 656 -10 690 -8
rect 729 -10 763 -8
rect 802 -10 836 -8
rect 875 -10 909 -8
rect 948 -10 982 -8
rect 1021 -10 1055 -8
rect 1094 -10 1128 -8
rect 1167 -10 1201 -8
rect 1240 -10 1274 -8
rect 1313 -10 1347 -8
rect 1386 -10 1420 -8
rect 1459 -10 1493 -8
rect 1532 -10 1566 -8
rect 1605 -10 1639 -8
rect 1678 -10 1712 -8
rect 1751 -10 1785 -8
rect 1824 -10 1858 -8
rect 1898 -10 1932 -8
rect 1972 -10 2006 -8
rect 2046 -10 2080 -8
rect 2120 -10 2154 -8
rect 2194 -10 2228 -8
rect 2268 -10 2302 -8
rect 2342 -10 2376 -8
rect 2416 -10 2450 -8
rect 2490 -10 2524 -8
rect 2564 -10 2598 -8
rect 2638 -10 2672 -8
rect 364 -42 398 -10
rect 437 -42 471 -10
rect 510 -42 544 -10
rect 583 -42 617 -10
rect 656 -42 690 -10
rect 729 -42 763 -10
rect 802 -42 836 -10
rect 875 -42 909 -10
rect 948 -42 982 -10
rect 1021 -42 1055 -10
rect 1094 -42 1128 -10
rect 1167 -42 1201 -10
rect 1240 -42 1274 -10
rect 1313 -42 1347 -10
rect 1386 -42 1420 -10
rect 1459 -42 1493 -10
rect 1532 -42 1566 -10
rect 1605 -42 1639 -10
rect 1678 -42 1712 -10
rect 1751 -42 1785 -10
rect 1824 -42 1858 -10
rect 1898 -42 1932 -10
rect 1972 -42 2006 -10
rect 2046 -42 2080 -10
rect 2120 -42 2154 -10
rect 2194 -42 2228 -10
rect 2268 -42 2302 -10
rect 2342 -42 2376 -10
rect 2416 -42 2450 -10
rect 2490 -42 2524 -10
rect 2564 -42 2574 -10
rect 2574 -42 2598 -10
rect 2638 -42 2643 -10
rect 2643 -42 2672 -10
rect 2712 -42 2746 -8
rect 2786 -10 2820 -8
rect 2860 -10 2894 -8
rect 2934 -10 2968 -8
rect 3008 -10 3042 -8
rect 3082 -10 3116 -8
rect 3156 -10 3190 -8
rect 3230 -10 3264 -8
rect 2786 -42 2816 -10
rect 2816 -42 2820 -10
rect 2860 -42 2885 -10
rect 2885 -42 2894 -10
rect 2934 -42 2954 -10
rect 2954 -42 2968 -10
rect 3008 -42 3023 -10
rect 3023 -42 3042 -10
rect 3082 -42 3092 -10
rect 3092 -42 3116 -10
rect 3156 -42 3161 -10
rect 3161 -42 3190 -10
rect 3230 -42 3264 -10
rect 364 -112 398 -80
rect 437 -112 471 -80
rect 510 -112 544 -80
rect 583 -112 617 -80
rect 656 -112 690 -80
rect 729 -112 763 -80
rect 802 -112 836 -80
rect 875 -112 909 -80
rect 948 -112 982 -80
rect 1021 -112 1055 -80
rect 1094 -112 1128 -80
rect 1167 -112 1201 -80
rect 1240 -112 1274 -80
rect 1313 -112 1347 -80
rect 1386 -112 1420 -80
rect 1459 -112 1493 -80
rect 1532 -112 1566 -80
rect 1605 -112 1639 -80
rect 1678 -112 1712 -80
rect 1751 -112 1785 -80
rect 1824 -112 1858 -80
rect 1898 -112 1932 -80
rect 1972 -112 2006 -80
rect 2046 -112 2080 -80
rect 2120 -112 2154 -80
rect 2194 -112 2228 -80
rect 2268 -112 2302 -80
rect 2342 -112 2376 -80
rect 2416 -112 2450 -80
rect 2490 -112 2524 -80
rect 2564 -112 2574 -80
rect 2574 -112 2598 -80
rect 2638 -112 2643 -80
rect 2643 -112 2672 -80
rect 364 -114 398 -112
rect 437 -114 471 -112
rect 510 -114 544 -112
rect 583 -114 617 -112
rect 656 -114 690 -112
rect 729 -114 763 -112
rect 802 -114 836 -112
rect 875 -114 909 -112
rect 948 -114 982 -112
rect 1021 -114 1055 -112
rect 1094 -114 1128 -112
rect 1167 -114 1201 -112
rect 1240 -114 1274 -112
rect 1313 -114 1347 -112
rect 1386 -114 1420 -112
rect 1459 -114 1493 -112
rect 1532 -114 1566 -112
rect 1605 -114 1639 -112
rect 1678 -114 1712 -112
rect 1751 -114 1785 -112
rect 1824 -114 1858 -112
rect 1898 -114 1932 -112
rect 1972 -114 2006 -112
rect 2046 -114 2080 -112
rect 2120 -114 2154 -112
rect 2194 -114 2228 -112
rect 2268 -114 2302 -112
rect 2342 -114 2376 -112
rect 2416 -114 2450 -112
rect 2490 -114 2524 -112
rect 2564 -114 2598 -112
rect 2638 -114 2672 -112
rect 2712 -114 2746 -80
rect 2786 -112 2816 -80
rect 2816 -112 2820 -80
rect 2860 -112 2885 -80
rect 2885 -112 2894 -80
rect 2934 -112 2954 -80
rect 2954 -112 2968 -80
rect 3008 -112 3023 -80
rect 3023 -112 3042 -80
rect 3082 -112 3092 -80
rect 3092 -112 3116 -80
rect 3156 -112 3161 -80
rect 3161 -112 3190 -80
rect 3230 -112 3264 -80
rect 2786 -114 2820 -112
rect 2860 -114 2894 -112
rect 2934 -114 2968 -112
rect 3008 -114 3042 -112
rect 3082 -114 3116 -112
rect 3156 -114 3190 -112
rect 3230 -114 3264 -112
rect 3606 -10 3640 -8
rect 3680 -10 3714 -8
rect 3754 -10 3788 -8
rect 3828 -10 3862 -8
rect 3902 -10 3936 -8
rect 3976 -10 4010 -8
rect 4050 -10 4084 -8
rect 3606 -42 3640 -10
rect 3680 -42 3709 -10
rect 3709 -42 3714 -10
rect 3754 -42 3778 -10
rect 3778 -42 3788 -10
rect 3828 -42 3847 -10
rect 3847 -42 3862 -10
rect 3902 -42 3916 -10
rect 3916 -42 3936 -10
rect 3976 -42 3985 -10
rect 3985 -42 4010 -10
rect 4050 -42 4054 -10
rect 4054 -42 4084 -10
rect 4124 -42 4158 -8
rect 4198 -10 4232 -8
rect 4272 -10 4306 -8
rect 4346 -10 4380 -8
rect 4420 -10 4454 -8
rect 4494 -10 4528 -8
rect 4568 -10 4602 -8
rect 4642 -10 4676 -8
rect 4716 -10 4750 -8
rect 4790 -10 4824 -8
rect 4864 -10 4898 -8
rect 4938 -10 4972 -8
rect 5012 -10 5046 -8
rect 5085 -10 5119 -8
rect 5158 -10 5192 -8
rect 5231 -10 5265 -8
rect 5304 -10 5338 -8
rect 5377 -10 5411 -8
rect 5450 -10 5484 -8
rect 5523 -10 5557 -8
rect 5596 -10 5630 -8
rect 5669 -10 5703 -8
rect 5742 -10 5776 -8
rect 5815 -10 5849 -8
rect 5888 -10 5922 -8
rect 5961 -10 5995 -8
rect 6034 -10 6068 -8
rect 6107 -10 6141 -8
rect 6180 -10 6214 -8
rect 6253 -10 6287 -8
rect 6326 -10 6360 -8
rect 6399 -10 6433 -8
rect 6472 -10 6506 -8
rect 4198 -42 4227 -10
rect 4227 -42 4232 -10
rect 4272 -42 4296 -10
rect 4296 -42 4306 -10
rect 4346 -42 4380 -10
rect 4420 -42 4454 -10
rect 4494 -42 4528 -10
rect 4568 -42 4602 -10
rect 4642 -42 4676 -10
rect 4716 -42 4750 -10
rect 4790 -42 4824 -10
rect 4864 -42 4898 -10
rect 4938 -42 4972 -10
rect 5012 -42 5046 -10
rect 5085 -42 5119 -10
rect 5158 -42 5192 -10
rect 5231 -42 5265 -10
rect 5304 -42 5338 -10
rect 5377 -42 5411 -10
rect 5450 -42 5484 -10
rect 5523 -42 5557 -10
rect 5596 -42 5630 -10
rect 5669 -42 5703 -10
rect 5742 -42 5776 -10
rect 5815 -42 5849 -10
rect 5888 -42 5922 -10
rect 5961 -42 5995 -10
rect 6034 -42 6068 -10
rect 6107 -42 6141 -10
rect 6180 -42 6214 -10
rect 6253 -42 6287 -10
rect 6326 -42 6360 -10
rect 6399 -42 6433 -10
rect 6472 -42 6506 -10
rect 3606 -112 3640 -80
rect 3680 -112 3709 -80
rect 3709 -112 3714 -80
rect 3754 -112 3778 -80
rect 3778 -112 3788 -80
rect 3828 -112 3847 -80
rect 3847 -112 3862 -80
rect 3902 -112 3916 -80
rect 3916 -112 3936 -80
rect 3976 -112 3985 -80
rect 3985 -112 4010 -80
rect 4050 -112 4054 -80
rect 4054 -112 4084 -80
rect 3606 -114 3640 -112
rect 3680 -114 3714 -112
rect 3754 -114 3788 -112
rect 3828 -114 3862 -112
rect 3902 -114 3936 -112
rect 3976 -114 4010 -112
rect 4050 -114 4084 -112
rect 4124 -114 4158 -80
rect 4198 -112 4227 -80
rect 4227 -112 4232 -80
rect 4272 -112 4296 -80
rect 4296 -112 4306 -80
rect 4346 -112 4380 -80
rect 4420 -112 4454 -80
rect 4494 -112 4528 -80
rect 4568 -112 4602 -80
rect 4642 -112 4676 -80
rect 4716 -112 4750 -80
rect 4790 -112 4824 -80
rect 4864 -112 4898 -80
rect 4938 -112 4972 -80
rect 5012 -112 5046 -80
rect 5085 -112 5119 -80
rect 5158 -112 5192 -80
rect 5231 -112 5265 -80
rect 5304 -112 5338 -80
rect 5377 -112 5411 -80
rect 5450 -112 5484 -80
rect 5523 -112 5557 -80
rect 5596 -112 5630 -80
rect 5669 -112 5703 -80
rect 5742 -112 5776 -80
rect 5815 -112 5849 -80
rect 5888 -112 5922 -80
rect 5961 -112 5995 -80
rect 6034 -112 6068 -80
rect 6107 -112 6141 -80
rect 6180 -112 6214 -80
rect 6253 -112 6287 -80
rect 6326 -112 6360 -80
rect 6399 -112 6433 -80
rect 6472 -112 6506 -80
rect 4198 -114 4232 -112
rect 4272 -114 4306 -112
rect 4346 -114 4380 -112
rect 4420 -114 4454 -112
rect 4494 -114 4528 -112
rect 4568 -114 4602 -112
rect 4642 -114 4676 -112
rect 4716 -114 4750 -112
rect 4790 -114 4824 -112
rect 4864 -114 4898 -112
rect 4938 -114 4972 -112
rect 5012 -114 5046 -112
rect 5085 -114 5119 -112
rect 5158 -114 5192 -112
rect 5231 -114 5265 -112
rect 5304 -114 5338 -112
rect 5377 -114 5411 -112
rect 5450 -114 5484 -112
rect 5523 -114 5557 -112
rect 5596 -114 5630 -112
rect 5669 -114 5703 -112
rect 5742 -114 5776 -112
rect 5815 -114 5849 -112
rect 5888 -114 5922 -112
rect 5961 -114 5995 -112
rect 6034 -114 6068 -112
rect 6107 -114 6141 -112
rect 6180 -114 6214 -112
rect 6253 -114 6287 -112
rect 6326 -114 6360 -112
rect 6399 -114 6433 -112
rect 6472 -114 6506 -112
rect 6848 -10 6882 -8
rect 6921 -10 6955 -8
rect 6994 -10 7028 -8
rect 7067 -10 7101 -8
rect 7140 -10 7174 -8
rect 7213 -10 7247 -8
rect 7286 -10 7320 -8
rect 7359 -10 7393 -8
rect 7432 -10 7466 -8
rect 7505 -10 7539 -8
rect 7578 -10 7612 -8
rect 7651 -10 7685 -8
rect 7724 -10 7758 -8
rect 7797 -10 7831 -8
rect 7870 -10 7904 -8
rect 7943 -10 7977 -8
rect 8016 -10 8050 -8
rect 8089 -10 8123 -8
rect 8162 -10 8196 -8
rect 8235 -10 8269 -8
rect 8308 -10 8342 -8
rect 8382 -10 8416 -8
rect 8456 -10 8490 -8
rect 8530 -10 8564 -8
rect 8604 -10 8638 -8
rect 8678 -10 8712 -8
rect 8752 -10 8786 -8
rect 8826 -10 8860 -8
rect 8900 -10 8934 -8
rect 8974 -10 9008 -8
rect 9048 -10 9082 -8
rect 9122 -10 9156 -8
rect 6848 -42 6882 -10
rect 6921 -42 6955 -10
rect 6994 -42 7028 -10
rect 7067 -42 7101 -10
rect 7140 -42 7174 -10
rect 7213 -42 7247 -10
rect 7286 -42 7320 -10
rect 7359 -42 7393 -10
rect 7432 -42 7466 -10
rect 7505 -42 7539 -10
rect 7578 -42 7612 -10
rect 7651 -42 7685 -10
rect 7724 -42 7758 -10
rect 7797 -42 7831 -10
rect 7870 -42 7904 -10
rect 7943 -42 7977 -10
rect 8016 -42 8050 -10
rect 8089 -42 8123 -10
rect 8162 -42 8196 -10
rect 8235 -42 8269 -10
rect 8308 -42 8342 -10
rect 8382 -42 8416 -10
rect 8456 -42 8490 -10
rect 8530 -42 8564 -10
rect 8604 -42 8638 -10
rect 8678 -42 8712 -10
rect 8752 -42 8786 -10
rect 8826 -42 8860 -10
rect 8900 -42 8934 -10
rect 8974 -42 9008 -10
rect 9048 -42 9058 -10
rect 9058 -42 9082 -10
rect 9122 -42 9127 -10
rect 9127 -42 9156 -10
rect 9196 -42 9230 -8
rect 9270 -10 9304 -8
rect 9344 -10 9378 -8
rect 9418 -10 9452 -8
rect 9492 -10 9526 -8
rect 9566 -10 9600 -8
rect 9640 -10 9674 -8
rect 9714 -10 9748 -8
rect 9270 -42 9300 -10
rect 9300 -42 9304 -10
rect 9344 -42 9369 -10
rect 9369 -42 9378 -10
rect 9418 -42 9438 -10
rect 9438 -42 9452 -10
rect 9492 -42 9507 -10
rect 9507 -42 9526 -10
rect 9566 -42 9576 -10
rect 9576 -42 9600 -10
rect 9640 -42 9645 -10
rect 9645 -42 9674 -10
rect 9714 -42 9748 -10
rect 6848 -112 6882 -80
rect 6921 -112 6955 -80
rect 6994 -112 7028 -80
rect 7067 -112 7101 -80
rect 7140 -112 7174 -80
rect 7213 -112 7247 -80
rect 7286 -112 7320 -80
rect 7359 -112 7393 -80
rect 7432 -112 7466 -80
rect 7505 -112 7539 -80
rect 7578 -112 7612 -80
rect 7651 -112 7685 -80
rect 7724 -112 7758 -80
rect 7797 -112 7831 -80
rect 7870 -112 7904 -80
rect 7943 -112 7977 -80
rect 8016 -112 8050 -80
rect 8089 -112 8123 -80
rect 8162 -112 8196 -80
rect 8235 -112 8269 -80
rect 8308 -112 8342 -80
rect 8382 -112 8416 -80
rect 8456 -112 8490 -80
rect 8530 -112 8564 -80
rect 8604 -112 8638 -80
rect 8678 -112 8712 -80
rect 8752 -112 8786 -80
rect 8826 -112 8860 -80
rect 8900 -112 8934 -80
rect 8974 -112 9008 -80
rect 9048 -112 9058 -80
rect 9058 -112 9082 -80
rect 9122 -112 9127 -80
rect 9127 -112 9156 -80
rect 6848 -114 6882 -112
rect 6921 -114 6955 -112
rect 6994 -114 7028 -112
rect 7067 -114 7101 -112
rect 7140 -114 7174 -112
rect 7213 -114 7247 -112
rect 7286 -114 7320 -112
rect 7359 -114 7393 -112
rect 7432 -114 7466 -112
rect 7505 -114 7539 -112
rect 7578 -114 7612 -112
rect 7651 -114 7685 -112
rect 7724 -114 7758 -112
rect 7797 -114 7831 -112
rect 7870 -114 7904 -112
rect 7943 -114 7977 -112
rect 8016 -114 8050 -112
rect 8089 -114 8123 -112
rect 8162 -114 8196 -112
rect 8235 -114 8269 -112
rect 8308 -114 8342 -112
rect 8382 -114 8416 -112
rect 8456 -114 8490 -112
rect 8530 -114 8564 -112
rect 8604 -114 8638 -112
rect 8678 -114 8712 -112
rect 8752 -114 8786 -112
rect 8826 -114 8860 -112
rect 8900 -114 8934 -112
rect 8974 -114 9008 -112
rect 9048 -114 9082 -112
rect 9122 -114 9156 -112
rect 9196 -114 9230 -80
rect 9270 -112 9300 -80
rect 9300 -112 9304 -80
rect 9344 -112 9369 -80
rect 9369 -112 9378 -80
rect 9418 -112 9438 -80
rect 9438 -112 9452 -80
rect 9492 -112 9507 -80
rect 9507 -112 9526 -80
rect 9566 -112 9576 -80
rect 9576 -112 9600 -80
rect 9640 -112 9645 -80
rect 9645 -112 9674 -80
rect 9714 -112 9748 -80
rect 9270 -114 9304 -112
rect 9344 -114 9378 -112
rect 9418 -114 9452 -112
rect 9492 -114 9526 -112
rect 9566 -114 9600 -112
rect 9640 -114 9674 -112
rect 9714 -114 9748 -112
rect 10090 -10 10124 -8
rect 10164 -10 10198 -8
rect 10238 -10 10272 -8
rect 10312 -10 10346 -8
rect 10386 -10 10420 -8
rect 10460 -10 10494 -8
rect 10534 -10 10568 -8
rect 10090 -42 10124 -10
rect 10164 -42 10193 -10
rect 10193 -42 10198 -10
rect 10238 -42 10262 -10
rect 10262 -42 10272 -10
rect 10312 -42 10331 -10
rect 10331 -42 10346 -10
rect 10386 -42 10400 -10
rect 10400 -42 10420 -10
rect 10460 -42 10469 -10
rect 10469 -42 10494 -10
rect 10534 -42 10538 -10
rect 10538 -42 10568 -10
rect 10608 -42 10642 -8
rect 10682 -10 10716 -8
rect 10756 -10 10790 -8
rect 10830 -10 10864 -8
rect 10904 -10 10938 -8
rect 10978 -10 11012 -8
rect 11052 -10 11086 -8
rect 11126 -10 11160 -8
rect 11200 -10 11234 -8
rect 11274 -10 11308 -8
rect 11348 -10 11382 -8
rect 11422 -10 11456 -8
rect 11496 -10 11530 -8
rect 11569 -10 11603 -8
rect 11642 -10 11676 -8
rect 11715 -10 11749 -8
rect 11788 -10 11822 -8
rect 11861 -10 11895 -8
rect 11934 -10 11968 -8
rect 12007 -10 12041 -8
rect 12080 -10 12114 -8
rect 12153 -10 12187 -8
rect 12226 -10 12260 -8
rect 12299 -10 12333 -8
rect 12372 -10 12406 -8
rect 12445 -10 12479 -8
rect 12518 -10 12552 -8
rect 12591 -10 12625 -8
rect 12664 -10 12698 -8
rect 12737 -10 12771 -8
rect 12810 -10 12844 -8
rect 12883 -10 12917 -8
rect 12956 -10 12990 -8
rect 10682 -42 10711 -10
rect 10711 -42 10716 -10
rect 10756 -42 10780 -10
rect 10780 -42 10790 -10
rect 10830 -42 10864 -10
rect 10904 -42 10938 -10
rect 10978 -42 11012 -10
rect 11052 -42 11086 -10
rect 11126 -42 11160 -10
rect 11200 -42 11234 -10
rect 11274 -42 11308 -10
rect 11348 -42 11382 -10
rect 11422 -42 11456 -10
rect 11496 -42 11530 -10
rect 11569 -42 11603 -10
rect 11642 -42 11676 -10
rect 11715 -42 11749 -10
rect 11788 -42 11822 -10
rect 11861 -42 11895 -10
rect 11934 -42 11968 -10
rect 12007 -42 12041 -10
rect 12080 -42 12114 -10
rect 12153 -42 12187 -10
rect 12226 -42 12260 -10
rect 12299 -42 12333 -10
rect 12372 -42 12406 -10
rect 12445 -42 12479 -10
rect 12518 -42 12552 -10
rect 12591 -42 12625 -10
rect 12664 -42 12698 -10
rect 12737 -42 12771 -10
rect 12810 -42 12844 -10
rect 12883 -42 12917 -10
rect 12956 -42 12990 -10
rect 10090 -112 10124 -80
rect 10164 -112 10193 -80
rect 10193 -112 10198 -80
rect 10238 -112 10262 -80
rect 10262 -112 10272 -80
rect 10312 -112 10331 -80
rect 10331 -112 10346 -80
rect 10386 -112 10400 -80
rect 10400 -112 10420 -80
rect 10460 -112 10469 -80
rect 10469 -112 10494 -80
rect 10534 -112 10538 -80
rect 10538 -112 10568 -80
rect 10090 -114 10124 -112
rect 10164 -114 10198 -112
rect 10238 -114 10272 -112
rect 10312 -114 10346 -112
rect 10386 -114 10420 -112
rect 10460 -114 10494 -112
rect 10534 -114 10568 -112
rect 10608 -114 10642 -80
rect 10682 -112 10711 -80
rect 10711 -112 10716 -80
rect 10756 -112 10780 -80
rect 10780 -112 10790 -80
rect 10830 -112 10864 -80
rect 10904 -112 10938 -80
rect 10978 -112 11012 -80
rect 11052 -112 11086 -80
rect 11126 -112 11160 -80
rect 11200 -112 11234 -80
rect 11274 -112 11308 -80
rect 11348 -112 11382 -80
rect 11422 -112 11456 -80
rect 11496 -112 11530 -80
rect 11569 -112 11603 -80
rect 11642 -112 11676 -80
rect 11715 -112 11749 -80
rect 11788 -112 11822 -80
rect 11861 -112 11895 -80
rect 11934 -112 11968 -80
rect 12007 -112 12041 -80
rect 12080 -112 12114 -80
rect 12153 -112 12187 -80
rect 12226 -112 12260 -80
rect 12299 -112 12333 -80
rect 12372 -112 12406 -80
rect 12445 -112 12479 -80
rect 12518 -112 12552 -80
rect 12591 -112 12625 -80
rect 12664 -112 12698 -80
rect 12737 -112 12771 -80
rect 12810 -112 12844 -80
rect 12883 -112 12917 -80
rect 12956 -112 12990 -80
rect 10682 -114 10716 -112
rect 10756 -114 10790 -112
rect 10830 -114 10864 -112
rect 10904 -114 10938 -112
rect 10978 -114 11012 -112
rect 11052 -114 11086 -112
rect 11126 -114 11160 -112
rect 11200 -114 11234 -112
rect 11274 -114 11308 -112
rect 11348 -114 11382 -112
rect 11422 -114 11456 -112
rect 11496 -114 11530 -112
rect 11569 -114 11603 -112
rect 11642 -114 11676 -112
rect 11715 -114 11749 -112
rect 11788 -114 11822 -112
rect 11861 -114 11895 -112
rect 11934 -114 11968 -112
rect 12007 -114 12041 -112
rect 12080 -114 12114 -112
rect 12153 -114 12187 -112
rect 12226 -114 12260 -112
rect 12299 -114 12333 -112
rect 12372 -114 12406 -112
rect 12445 -114 12479 -112
rect 12518 -114 12552 -112
rect 12591 -114 12625 -112
rect 12664 -114 12698 -112
rect 12737 -114 12771 -112
rect 12810 -114 12844 -112
rect 12883 -114 12917 -112
rect 12956 -114 12990 -112
rect 13332 -10 13366 -8
rect 13405 -10 13439 -8
rect 13478 -10 13512 -8
rect 13551 -10 13585 -8
rect 13624 -10 13658 -8
rect 13697 -10 13731 -8
rect 13770 -10 13804 -8
rect 13843 -10 13877 -8
rect 13916 -10 13950 -8
rect 13989 -10 14023 -8
rect 14062 -10 14096 -8
rect 14135 -10 14169 -8
rect 14208 -10 14242 -8
rect 14281 -10 14315 -8
rect 14354 -10 14388 -8
rect 14427 -10 14461 -8
rect 14500 -10 14534 -8
rect 14573 -10 14607 -8
rect 14646 -10 14680 -8
rect 14719 -10 14753 -8
rect 14792 -10 14826 -8
rect 14866 -10 14900 -8
rect 14940 -10 14974 -8
rect 15014 -10 15048 -8
rect 15088 -10 15122 -8
rect 15162 -10 15196 -8
rect 15236 -10 15270 -8
rect 15310 -10 15344 -8
rect 15384 -10 15418 -8
rect 15458 -10 15492 -8
rect 15532 -10 15566 -8
rect 15606 -10 15640 -8
rect 13332 -42 13366 -10
rect 13405 -42 13439 -10
rect 13478 -42 13512 -10
rect 13551 -42 13585 -10
rect 13624 -42 13658 -10
rect 13697 -42 13731 -10
rect 13770 -42 13804 -10
rect 13843 -42 13877 -10
rect 13916 -42 13950 -10
rect 13989 -42 14023 -10
rect 14062 -42 14096 -10
rect 14135 -42 14169 -10
rect 14208 -42 14242 -10
rect 14281 -42 14315 -10
rect 14354 -42 14388 -10
rect 14427 -42 14461 -10
rect 14500 -42 14534 -10
rect 14573 -42 14607 -10
rect 14646 -42 14680 -10
rect 14719 -42 14753 -10
rect 14792 -42 14826 -10
rect 14866 -42 14900 -10
rect 14940 -42 14974 -10
rect 15014 -42 15048 -10
rect 15088 -42 15122 -10
rect 15162 -42 15196 -10
rect 15236 -42 15270 -10
rect 15310 -42 15344 -10
rect 15384 -42 15418 -10
rect 15458 -42 15492 -10
rect 15532 -42 15542 -10
rect 15542 -42 15566 -10
rect 15606 -42 15611 -10
rect 15611 -42 15640 -10
rect 15680 -42 15714 -8
rect 15754 -10 15788 -8
rect 15828 -10 15862 -8
rect 15902 -10 15936 -8
rect 15976 -10 16010 -8
rect 16050 -10 16084 -8
rect 16124 -10 16158 -8
rect 16198 -10 16232 -8
rect 15754 -42 15784 -10
rect 15784 -42 15788 -10
rect 15828 -42 15853 -10
rect 15853 -42 15862 -10
rect 15902 -42 15922 -10
rect 15922 -42 15936 -10
rect 15976 -42 15991 -10
rect 15991 -42 16010 -10
rect 16050 -42 16060 -10
rect 16060 -42 16084 -10
rect 16124 -42 16129 -10
rect 16129 -42 16158 -10
rect 16198 -42 16232 -10
rect 13332 -112 13366 -80
rect 13405 -112 13439 -80
rect 13478 -112 13512 -80
rect 13551 -112 13585 -80
rect 13624 -112 13658 -80
rect 13697 -112 13731 -80
rect 13770 -112 13804 -80
rect 13843 -112 13877 -80
rect 13916 -112 13950 -80
rect 13989 -112 14023 -80
rect 14062 -112 14096 -80
rect 14135 -112 14169 -80
rect 14208 -112 14242 -80
rect 14281 -112 14315 -80
rect 14354 -112 14388 -80
rect 14427 -112 14461 -80
rect 14500 -112 14534 -80
rect 14573 -112 14607 -80
rect 14646 -112 14680 -80
rect 14719 -112 14753 -80
rect 14792 -112 14826 -80
rect 14866 -112 14900 -80
rect 14940 -112 14974 -80
rect 15014 -112 15048 -80
rect 15088 -112 15122 -80
rect 15162 -112 15196 -80
rect 15236 -112 15270 -80
rect 15310 -112 15344 -80
rect 15384 -112 15418 -80
rect 15458 -112 15492 -80
rect 15532 -112 15542 -80
rect 15542 -112 15566 -80
rect 15606 -112 15611 -80
rect 15611 -112 15640 -80
rect 13332 -114 13366 -112
rect 13405 -114 13439 -112
rect 13478 -114 13512 -112
rect 13551 -114 13585 -112
rect 13624 -114 13658 -112
rect 13697 -114 13731 -112
rect 13770 -114 13804 -112
rect 13843 -114 13877 -112
rect 13916 -114 13950 -112
rect 13989 -114 14023 -112
rect 14062 -114 14096 -112
rect 14135 -114 14169 -112
rect 14208 -114 14242 -112
rect 14281 -114 14315 -112
rect 14354 -114 14388 -112
rect 14427 -114 14461 -112
rect 14500 -114 14534 -112
rect 14573 -114 14607 -112
rect 14646 -114 14680 -112
rect 14719 -114 14753 -112
rect 14792 -114 14826 -112
rect 14866 -114 14900 -112
rect 14940 -114 14974 -112
rect 15014 -114 15048 -112
rect 15088 -114 15122 -112
rect 15162 -114 15196 -112
rect 15236 -114 15270 -112
rect 15310 -114 15344 -112
rect 15384 -114 15418 -112
rect 15458 -114 15492 -112
rect 15532 -114 15566 -112
rect 15606 -114 15640 -112
rect 15680 -114 15714 -80
rect 15754 -112 15784 -80
rect 15784 -112 15788 -80
rect 15828 -112 15853 -80
rect 15853 -112 15862 -80
rect 15902 -112 15922 -80
rect 15922 -112 15936 -80
rect 15976 -112 15991 -80
rect 15991 -112 16010 -80
rect 16050 -112 16060 -80
rect 16060 -112 16084 -80
rect 16124 -112 16129 -80
rect 16129 -112 16158 -80
rect 16198 -112 16232 -80
rect 15754 -114 15788 -112
rect 15828 -114 15862 -112
rect 15902 -114 15936 -112
rect 15976 -114 16010 -112
rect 16050 -114 16084 -112
rect 16124 -114 16158 -112
rect 16198 -114 16232 -112
rect 16574 -10 16608 -8
rect 16648 -10 16682 -8
rect 16722 -10 16756 -8
rect 16796 -10 16830 -8
rect 16870 -10 16904 -8
rect 16944 -10 16978 -8
rect 17018 -10 17052 -8
rect 16574 -42 16608 -10
rect 16648 -42 16677 -10
rect 16677 -42 16682 -10
rect 16722 -42 16746 -10
rect 16746 -42 16756 -10
rect 16796 -42 16815 -10
rect 16815 -42 16830 -10
rect 16870 -42 16884 -10
rect 16884 -42 16904 -10
rect 16944 -42 16953 -10
rect 16953 -42 16978 -10
rect 17018 -42 17022 -10
rect 17022 -42 17052 -10
rect 17092 -42 17126 -8
rect 17166 -10 17200 -8
rect 17240 -10 17274 -8
rect 17314 -10 17348 -8
rect 17388 -10 17422 -8
rect 17462 -10 17496 -8
rect 17536 -10 17570 -8
rect 17610 -10 17644 -8
rect 17684 -10 17718 -8
rect 17758 -10 17792 -8
rect 17832 -10 17866 -8
rect 17906 -10 17940 -8
rect 17980 -10 18014 -8
rect 18053 -10 18087 -8
rect 18126 -10 18160 -8
rect 18199 -10 18233 -8
rect 18272 -10 18306 -8
rect 18345 -10 18379 -8
rect 18418 -10 18452 -8
rect 18491 -10 18525 -8
rect 18564 -10 18598 -8
rect 18637 -10 18671 -8
rect 18710 -10 18744 -8
rect 18783 -10 18817 -8
rect 18856 -10 18890 -8
rect 18929 -10 18963 -8
rect 19002 -10 19036 -8
rect 19075 -10 19109 -8
rect 19148 -10 19182 -8
rect 19221 -10 19255 -8
rect 19294 -10 19328 -8
rect 19367 -10 19401 -8
rect 19440 -10 19474 -8
rect 17166 -42 17195 -10
rect 17195 -42 17200 -10
rect 17240 -42 17264 -10
rect 17264 -42 17274 -10
rect 17314 -42 17348 -10
rect 17388 -42 17422 -10
rect 17462 -42 17496 -10
rect 17536 -42 17570 -10
rect 17610 -42 17644 -10
rect 17684 -42 17718 -10
rect 17758 -42 17792 -10
rect 17832 -42 17866 -10
rect 17906 -42 17940 -10
rect 17980 -42 18014 -10
rect 18053 -42 18087 -10
rect 18126 -42 18160 -10
rect 18199 -42 18233 -10
rect 18272 -42 18306 -10
rect 18345 -42 18379 -10
rect 18418 -42 18452 -10
rect 18491 -42 18525 -10
rect 18564 -42 18598 -10
rect 18637 -42 18671 -10
rect 18710 -42 18744 -10
rect 18783 -42 18817 -10
rect 18856 -42 18890 -10
rect 18929 -42 18963 -10
rect 19002 -42 19036 -10
rect 19075 -42 19109 -10
rect 19148 -42 19182 -10
rect 19221 -42 19255 -10
rect 19294 -42 19328 -10
rect 19367 -42 19401 -10
rect 19440 -42 19474 -10
rect 16574 -112 16608 -80
rect 16648 -112 16677 -80
rect 16677 -112 16682 -80
rect 16722 -112 16746 -80
rect 16746 -112 16756 -80
rect 16796 -112 16815 -80
rect 16815 -112 16830 -80
rect 16870 -112 16884 -80
rect 16884 -112 16904 -80
rect 16944 -112 16953 -80
rect 16953 -112 16978 -80
rect 17018 -112 17022 -80
rect 17022 -112 17052 -80
rect 16574 -114 16608 -112
rect 16648 -114 16682 -112
rect 16722 -114 16756 -112
rect 16796 -114 16830 -112
rect 16870 -114 16904 -112
rect 16944 -114 16978 -112
rect 17018 -114 17052 -112
rect 17092 -114 17126 -80
rect 17166 -112 17195 -80
rect 17195 -112 17200 -80
rect 17240 -112 17264 -80
rect 17264 -112 17274 -80
rect 17314 -112 17348 -80
rect 17388 -112 17422 -80
rect 17462 -112 17496 -80
rect 17536 -112 17570 -80
rect 17610 -112 17644 -80
rect 17684 -112 17718 -80
rect 17758 -112 17792 -80
rect 17832 -112 17866 -80
rect 17906 -112 17940 -80
rect 17980 -112 18014 -80
rect 18053 -112 18087 -80
rect 18126 -112 18160 -80
rect 18199 -112 18233 -80
rect 18272 -112 18306 -80
rect 18345 -112 18379 -80
rect 18418 -112 18452 -80
rect 18491 -112 18525 -80
rect 18564 -112 18598 -80
rect 18637 -112 18671 -80
rect 18710 -112 18744 -80
rect 18783 -112 18817 -80
rect 18856 -112 18890 -80
rect 18929 -112 18963 -80
rect 19002 -112 19036 -80
rect 19075 -112 19109 -80
rect 19148 -112 19182 -80
rect 19221 -112 19255 -80
rect 19294 -112 19328 -80
rect 19367 -112 19401 -80
rect 19440 -112 19474 -80
rect 17166 -114 17200 -112
rect 17240 -114 17274 -112
rect 17314 -114 17348 -112
rect 17388 -114 17422 -112
rect 17462 -114 17496 -112
rect 17536 -114 17570 -112
rect 17610 -114 17644 -112
rect 17684 -114 17718 -112
rect 17758 -114 17792 -112
rect 17832 -114 17866 -112
rect 17906 -114 17940 -112
rect 17980 -114 18014 -112
rect 18053 -114 18087 -112
rect 18126 -114 18160 -112
rect 18199 -114 18233 -112
rect 18272 -114 18306 -112
rect 18345 -114 18379 -112
rect 18418 -114 18452 -112
rect 18491 -114 18525 -112
rect 18564 -114 18598 -112
rect 18637 -114 18671 -112
rect 18710 -114 18744 -112
rect 18783 -114 18817 -112
rect 18856 -114 18890 -112
rect 18929 -114 18963 -112
rect 19002 -114 19036 -112
rect 19075 -114 19109 -112
rect 19148 -114 19182 -112
rect 19221 -114 19255 -112
rect 19294 -114 19328 -112
rect 19367 -114 19401 -112
rect 19440 -114 19474 -112
rect 19882 -41 19888 -39
rect 19888 -41 19916 -39
rect 19882 -73 19916 -41
rect -46 -183 -12 -149
rect 42 -183 76 -149
rect 19882 -145 19916 -111
rect 8 -272 42 -238
rect 80 -272 82 -238
rect 82 -272 114 -238
rect 152 -272 184 -238
rect 184 -272 186 -238
rect 224 -272 252 -238
rect 252 -272 258 -238
rect 296 -272 320 -238
rect 320 -272 330 -238
rect 368 -272 388 -238
rect 388 -272 402 -238
rect 440 -272 456 -238
rect 456 -272 474 -238
rect 512 -272 524 -238
rect 524 -272 546 -238
rect 584 -272 592 -238
rect 592 -272 618 -238
rect 656 -272 660 -238
rect 660 -272 690 -238
rect 728 -272 762 -238
rect 800 -272 830 -238
rect 830 -272 834 -238
rect 872 -272 898 -238
rect 898 -272 906 -238
rect 944 -272 966 -238
rect 966 -272 978 -238
rect 1016 -272 1034 -238
rect 1034 -272 1050 -238
rect 1088 -272 1102 -238
rect 1102 -272 1122 -238
rect 1160 -272 1170 -238
rect 1170 -272 1194 -238
rect 1232 -272 1238 -238
rect 1238 -272 1266 -238
rect 1304 -272 1306 -238
rect 1306 -272 1338 -238
rect 1376 -272 1408 -238
rect 1408 -272 1410 -238
rect 1448 -272 1476 -238
rect 1476 -272 1482 -238
rect 1520 -272 1544 -238
rect 1544 -272 1554 -238
rect 1592 -272 1612 -238
rect 1612 -272 1626 -238
rect 1664 -272 1680 -238
rect 1680 -272 1698 -238
rect 1736 -272 1748 -238
rect 1748 -272 1770 -238
rect 1808 -272 1816 -238
rect 1816 -272 1842 -238
rect 1880 -272 1884 -238
rect 1884 -272 1914 -238
rect 1952 -272 1986 -238
rect 2024 -272 2054 -238
rect 2054 -272 2058 -238
rect 2096 -272 2122 -238
rect 2122 -272 2130 -238
rect 2168 -272 2190 -238
rect 2190 -272 2202 -238
rect 2240 -272 2258 -238
rect 2258 -272 2274 -238
rect 2312 -272 2326 -238
rect 2326 -272 2346 -238
rect 2384 -272 2394 -238
rect 2394 -272 2418 -238
rect 2456 -272 2462 -238
rect 2462 -272 2490 -238
rect 2528 -272 2530 -238
rect 2530 -272 2562 -238
rect 2600 -272 2632 -238
rect 2632 -272 2634 -238
rect 2672 -272 2700 -238
rect 2700 -272 2706 -238
rect 2744 -272 2768 -238
rect 2768 -272 2778 -238
rect 2816 -272 2836 -238
rect 2836 -272 2850 -238
rect 2888 -272 2904 -238
rect 2904 -272 2922 -238
rect 2960 -272 2972 -238
rect 2972 -272 2994 -238
rect 3032 -272 3040 -238
rect 3040 -272 3066 -238
rect 3104 -272 3108 -238
rect 3108 -272 3138 -238
rect 3176 -272 3210 -238
rect 3248 -272 3278 -238
rect 3278 -272 3282 -238
rect 3320 -272 3346 -238
rect 3346 -272 3354 -238
rect 3392 -272 3414 -238
rect 3414 -272 3426 -238
rect 3464 -272 3482 -238
rect 3482 -272 3498 -238
rect 3536 -272 3550 -238
rect 3550 -272 3570 -238
rect 3608 -272 3618 -238
rect 3618 -272 3642 -238
rect 3680 -272 3686 -238
rect 3686 -272 3714 -238
rect 3752 -272 3754 -238
rect 3754 -272 3786 -238
rect 3824 -272 3856 -238
rect 3856 -272 3858 -238
rect 3896 -272 3924 -238
rect 3924 -272 3930 -238
rect 3968 -272 3992 -238
rect 3992 -272 4002 -238
rect 4040 -272 4060 -238
rect 4060 -272 4074 -238
rect 4112 -272 4128 -238
rect 4128 -272 4146 -238
rect 4184 -272 4196 -238
rect 4196 -272 4218 -238
rect 4256 -272 4264 -238
rect 4264 -272 4290 -238
rect 4328 -272 4332 -238
rect 4332 -272 4362 -238
rect 4400 -272 4434 -238
rect 4472 -272 4502 -238
rect 4502 -272 4506 -238
rect 4544 -272 4570 -238
rect 4570 -272 4578 -238
rect 4616 -272 4638 -238
rect 4638 -272 4650 -238
rect 4688 -272 4706 -238
rect 4706 -272 4722 -238
rect 4760 -272 4774 -238
rect 4774 -272 4794 -238
rect 4832 -272 4842 -238
rect 4842 -272 4866 -238
rect 4904 -272 4910 -238
rect 4910 -272 4938 -238
rect 4976 -272 4978 -238
rect 4978 -272 5010 -238
rect 5048 -272 5080 -238
rect 5080 -272 5082 -238
rect 5120 -272 5148 -238
rect 5148 -272 5154 -238
rect 5192 -272 5216 -238
rect 5216 -272 5226 -238
rect 5264 -272 5284 -238
rect 5284 -272 5298 -238
rect 5336 -272 5352 -238
rect 5352 -272 5370 -238
rect 5408 -272 5420 -238
rect 5420 -272 5442 -238
rect 5480 -272 5488 -238
rect 5488 -272 5514 -238
rect 5552 -272 5556 -238
rect 5556 -272 5586 -238
rect 5624 -272 5658 -238
rect 5696 -272 5726 -238
rect 5726 -272 5730 -238
rect 5768 -272 5794 -238
rect 5794 -272 5802 -238
rect 5840 -272 5862 -238
rect 5862 -272 5874 -238
rect 5912 -272 5930 -238
rect 5930 -272 5946 -238
rect 5984 -272 5998 -238
rect 5998 -272 6018 -238
rect 6056 -272 6066 -238
rect 6066 -272 6090 -238
rect 6128 -272 6134 -238
rect 6134 -272 6162 -238
rect 6200 -272 6202 -238
rect 6202 -272 6234 -238
rect 6272 -272 6304 -238
rect 6304 -272 6306 -238
rect 6344 -272 6372 -238
rect 6372 -272 6378 -238
rect 6416 -272 6440 -238
rect 6440 -272 6450 -238
rect 6488 -272 6508 -238
rect 6508 -272 6522 -238
rect 6560 -272 6576 -238
rect 6576 -272 6594 -238
rect 6632 -272 6644 -238
rect 6644 -272 6666 -238
rect 6704 -272 6712 -238
rect 6712 -272 6738 -238
rect 6776 -272 6780 -238
rect 6780 -272 6810 -238
rect 6848 -272 6882 -238
rect 6920 -272 6950 -238
rect 6950 -272 6954 -238
rect 6992 -272 7018 -238
rect 7018 -272 7026 -238
rect 7064 -272 7086 -238
rect 7086 -272 7098 -238
rect 7136 -272 7154 -238
rect 7154 -272 7170 -238
rect 7208 -272 7222 -238
rect 7222 -272 7242 -238
rect 7280 -272 7290 -238
rect 7290 -272 7314 -238
rect 7352 -272 7358 -238
rect 7358 -272 7386 -238
rect 7424 -272 7426 -238
rect 7426 -272 7458 -238
rect 7496 -272 7528 -238
rect 7528 -272 7530 -238
rect 7568 -272 7596 -238
rect 7596 -272 7602 -238
rect 7640 -272 7664 -238
rect 7664 -272 7674 -238
rect 7712 -272 7732 -238
rect 7732 -272 7746 -238
rect 7784 -272 7800 -238
rect 7800 -272 7818 -238
rect 7856 -272 7868 -238
rect 7868 -272 7890 -238
rect 7928 -272 7936 -238
rect 7936 -272 7962 -238
rect 8000 -272 8004 -238
rect 8004 -272 8034 -238
rect 8072 -272 8106 -238
rect 8144 -272 8174 -238
rect 8174 -272 8178 -238
rect 8216 -272 8242 -238
rect 8242 -272 8250 -238
rect 8288 -272 8310 -238
rect 8310 -272 8322 -238
rect 8360 -272 8378 -238
rect 8378 -272 8394 -238
rect 8432 -272 8446 -238
rect 8446 -272 8466 -238
rect 8504 -272 8514 -238
rect 8514 -272 8538 -238
rect 8576 -272 8582 -238
rect 8582 -272 8610 -238
rect 8648 -272 8650 -238
rect 8650 -272 8682 -238
rect 8720 -272 8752 -238
rect 8752 -272 8754 -238
rect 8792 -272 8820 -238
rect 8820 -272 8826 -238
rect 8864 -272 8888 -238
rect 8888 -272 8898 -238
rect 8936 -272 8956 -238
rect 8956 -272 8970 -238
rect 9008 -272 9024 -238
rect 9024 -272 9042 -238
rect 9080 -272 9092 -238
rect 9092 -272 9114 -238
rect 9152 -272 9160 -238
rect 9160 -272 9186 -238
rect 9224 -272 9228 -238
rect 9228 -272 9258 -238
rect 9296 -272 9330 -238
rect 9368 -272 9398 -238
rect 9398 -272 9402 -238
rect 9440 -272 9466 -238
rect 9466 -272 9474 -238
rect 9512 -272 9534 -238
rect 9534 -272 9546 -238
rect 9584 -272 9602 -238
rect 9602 -272 9618 -238
rect 9656 -272 9670 -238
rect 9670 -272 9690 -238
rect 9728 -272 9738 -238
rect 9738 -272 9762 -238
rect 9800 -272 9806 -238
rect 9806 -272 9834 -238
rect 9872 -272 9874 -238
rect 9874 -272 9906 -238
rect 9944 -272 9976 -238
rect 9976 -272 9978 -238
rect 10016 -272 10044 -238
rect 10044 -272 10050 -238
rect 10088 -272 10112 -238
rect 10112 -272 10122 -238
rect 10160 -272 10180 -238
rect 10180 -272 10194 -238
rect 10232 -272 10248 -238
rect 10248 -272 10266 -238
rect 10304 -272 10316 -238
rect 10316 -272 10338 -238
rect 10376 -272 10384 -238
rect 10384 -272 10410 -238
rect 10448 -272 10452 -238
rect 10452 -272 10482 -238
rect 10520 -272 10554 -238
rect 10592 -272 10622 -238
rect 10622 -272 10626 -238
rect 10664 -272 10690 -238
rect 10690 -272 10698 -238
rect 10736 -272 10758 -238
rect 10758 -272 10770 -238
rect 10808 -272 10826 -238
rect 10826 -272 10842 -238
rect 10880 -272 10894 -238
rect 10894 -272 10914 -238
rect 10952 -272 10962 -238
rect 10962 -272 10986 -238
rect 11024 -272 11030 -238
rect 11030 -272 11058 -238
rect 11096 -272 11098 -238
rect 11098 -272 11130 -238
rect 11168 -272 11200 -238
rect 11200 -272 11202 -238
rect 11240 -272 11268 -238
rect 11268 -272 11274 -238
rect 11312 -272 11336 -238
rect 11336 -272 11346 -238
rect 11384 -272 11404 -238
rect 11404 -272 11418 -238
rect 11456 -272 11472 -238
rect 11472 -272 11490 -238
rect 11528 -272 11540 -238
rect 11540 -272 11562 -238
rect 11600 -272 11608 -238
rect 11608 -272 11634 -238
rect 11672 -272 11676 -238
rect 11676 -272 11706 -238
rect 11744 -272 11778 -238
rect 11816 -272 11846 -238
rect 11846 -272 11850 -238
rect 11888 -272 11914 -238
rect 11914 -272 11922 -238
rect 11960 -272 11982 -238
rect 11982 -272 11994 -238
rect 12032 -272 12050 -238
rect 12050 -272 12066 -238
rect 12104 -272 12118 -238
rect 12118 -272 12138 -238
rect 12176 -272 12186 -238
rect 12186 -272 12210 -238
rect 12248 -272 12254 -238
rect 12254 -272 12282 -238
rect 12320 -272 12322 -238
rect 12322 -272 12354 -238
rect 12392 -272 12424 -238
rect 12424 -272 12426 -238
rect 12464 -272 12492 -238
rect 12492 -272 12498 -238
rect 12536 -272 12560 -238
rect 12560 -272 12570 -238
rect 12608 -272 12628 -238
rect 12628 -272 12642 -238
rect 12680 -272 12696 -238
rect 12696 -272 12714 -238
rect 12752 -272 12764 -238
rect 12764 -272 12786 -238
rect 12824 -272 12832 -238
rect 12832 -272 12858 -238
rect 12896 -272 12900 -238
rect 12900 -272 12930 -238
rect 12968 -272 13002 -238
rect 13040 -272 13070 -238
rect 13070 -272 13074 -238
rect 13112 -272 13138 -238
rect 13138 -272 13146 -238
rect 13184 -272 13206 -238
rect 13206 -272 13218 -238
rect 13256 -272 13274 -238
rect 13274 -272 13290 -238
rect 13328 -272 13342 -238
rect 13342 -272 13362 -238
rect 13400 -272 13410 -238
rect 13410 -272 13434 -238
rect 13472 -272 13478 -238
rect 13478 -272 13506 -238
rect 13544 -272 13546 -238
rect 13546 -272 13578 -238
rect 13616 -272 13648 -238
rect 13648 -272 13650 -238
rect 13688 -272 13716 -238
rect 13716 -272 13722 -238
rect 13760 -272 13784 -238
rect 13784 -272 13794 -238
rect 13832 -272 13852 -238
rect 13852 -272 13866 -238
rect 13904 -272 13920 -238
rect 13920 -272 13938 -238
rect 13976 -272 13988 -238
rect 13988 -272 14010 -238
rect 14048 -272 14056 -238
rect 14056 -272 14082 -238
rect 14120 -272 14124 -238
rect 14124 -272 14154 -238
rect 14192 -272 14226 -238
rect 14264 -272 14294 -238
rect 14294 -272 14298 -238
rect 14336 -272 14362 -238
rect 14362 -272 14370 -238
rect 14408 -272 14430 -238
rect 14430 -272 14442 -238
rect 14480 -272 14498 -238
rect 14498 -272 14514 -238
rect 14552 -272 14566 -238
rect 14566 -272 14586 -238
rect 14624 -272 14634 -238
rect 14634 -272 14658 -238
rect 14696 -272 14702 -238
rect 14702 -272 14730 -238
rect 14768 -272 14770 -238
rect 14770 -272 14802 -238
rect 14840 -272 14872 -238
rect 14872 -272 14874 -238
rect 14912 -272 14940 -238
rect 14940 -272 14946 -238
rect 14984 -272 15008 -238
rect 15008 -272 15018 -238
rect 15056 -272 15076 -238
rect 15076 -272 15090 -238
rect 15128 -272 15144 -238
rect 15144 -272 15162 -238
rect 15200 -272 15212 -238
rect 15212 -272 15234 -238
rect 15272 -272 15280 -238
rect 15280 -272 15306 -238
rect 15344 -272 15348 -238
rect 15348 -272 15378 -238
rect 15416 -272 15450 -238
rect 15488 -272 15518 -238
rect 15518 -272 15522 -238
rect 15560 -272 15586 -238
rect 15586 -272 15594 -238
rect 15632 -272 15654 -238
rect 15654 -272 15666 -238
rect 15704 -272 15722 -238
rect 15722 -272 15738 -238
rect 15776 -272 15790 -238
rect 15790 -272 15810 -238
rect 15848 -272 15858 -238
rect 15858 -272 15882 -238
rect 15920 -272 15926 -238
rect 15926 -272 15954 -238
rect 15992 -272 15994 -238
rect 15994 -272 16026 -238
rect 16064 -272 16096 -238
rect 16096 -272 16098 -238
rect 16136 -272 16164 -238
rect 16164 -272 16170 -238
rect 16208 -272 16232 -238
rect 16232 -272 16242 -238
rect 16280 -272 16300 -238
rect 16300 -272 16314 -238
rect 16352 -272 16368 -238
rect 16368 -272 16386 -238
rect 16424 -272 16436 -238
rect 16436 -272 16458 -238
rect 16496 -272 16504 -238
rect 16504 -272 16530 -238
rect 16568 -272 16572 -238
rect 16572 -272 16602 -238
rect 16640 -272 16674 -238
rect 16712 -272 16742 -238
rect 16742 -272 16746 -238
rect 16784 -272 16810 -238
rect 16810 -272 16818 -238
rect 16856 -272 16878 -238
rect 16878 -272 16890 -238
rect 16928 -272 16946 -238
rect 16946 -272 16962 -238
rect 17000 -272 17014 -238
rect 17014 -272 17034 -238
rect 17072 -272 17082 -238
rect 17082 -272 17106 -238
rect 17144 -272 17150 -238
rect 17150 -272 17178 -238
rect 17216 -272 17218 -238
rect 17218 -272 17250 -238
rect 17288 -272 17320 -238
rect 17320 -272 17322 -238
rect 17360 -272 17388 -238
rect 17388 -272 17394 -238
rect 17432 -272 17456 -238
rect 17456 -272 17466 -238
rect 17504 -272 17524 -238
rect 17524 -272 17538 -238
rect 17576 -272 17592 -238
rect 17592 -272 17610 -238
rect 17648 -272 17660 -238
rect 17660 -272 17682 -238
rect 17720 -272 17728 -238
rect 17728 -272 17754 -238
rect 17792 -272 17796 -238
rect 17796 -272 17826 -238
rect 17864 -272 17898 -238
rect 17936 -272 17966 -238
rect 17966 -272 17970 -238
rect 18008 -272 18034 -238
rect 18034 -272 18042 -238
rect 18080 -272 18102 -238
rect 18102 -272 18114 -238
rect 18152 -272 18170 -238
rect 18170 -272 18186 -238
rect 18224 -272 18238 -238
rect 18238 -272 18258 -238
rect 18296 -272 18306 -238
rect 18306 -272 18330 -238
rect 18368 -272 18374 -238
rect 18374 -272 18402 -238
rect 18440 -272 18442 -238
rect 18442 -272 18474 -238
rect 18513 -272 18544 -238
rect 18544 -272 18547 -238
rect 18586 -272 18612 -238
rect 18612 -272 18620 -238
rect 18659 -272 18680 -238
rect 18680 -272 18693 -238
rect 18732 -272 18748 -238
rect 18748 -272 18766 -238
rect 18805 -272 18816 -238
rect 18816 -272 18839 -238
rect 18878 -272 18884 -238
rect 18884 -272 18912 -238
rect 18951 -272 18952 -238
rect 18952 -272 18985 -238
rect 19024 -272 19054 -238
rect 19054 -272 19058 -238
rect 19097 -272 19122 -238
rect 19122 -272 19131 -238
rect 19170 -272 19190 -238
rect 19190 -272 19204 -238
rect 19243 -272 19258 -238
rect 19258 -272 19277 -238
rect 19316 -272 19326 -238
rect 19326 -272 19350 -238
rect 19389 -272 19394 -238
rect 19394 -272 19423 -238
rect 19462 -272 19496 -238
rect 19535 -272 19564 -238
rect 19564 -272 19569 -238
rect 19608 -272 19632 -238
rect 19632 -272 19642 -238
rect 19681 -272 19700 -238
rect 19700 -272 19715 -238
rect 19754 -272 19768 -238
rect 19768 -272 19788 -238
rect 19827 -272 19836 -238
rect 19836 -272 19861 -238
<< metal1 >>
rect -2119 14521 -647 14527
rect -2119 14487 -2040 14521
rect -2006 14487 -1967 14521
rect -1933 14487 -1894 14521
rect -1860 14487 -1821 14521
rect -1787 14487 -1748 14521
rect -1714 14487 -1675 14521
rect -1641 14487 -1601 14521
rect -1567 14487 -1527 14521
rect -1493 14487 -1453 14521
rect -1419 14487 -1379 14521
rect -1345 14487 -1305 14521
rect -1271 14487 -1231 14521
rect -1197 14487 -1157 14521
rect -1123 14487 -1083 14521
rect -1049 14487 -1009 14521
rect -975 14487 -935 14521
rect -901 14487 -861 14521
rect -827 14487 -787 14521
rect -753 14487 -713 14521
rect -679 14487 -647 14521
rect -2119 14449 -647 14487
rect -2119 14415 -2113 14449
rect -2079 14415 -2041 14449
rect -2007 14415 -1967 14449
rect -1933 14415 -1894 14449
rect -1860 14415 -1821 14449
rect -1787 14415 -1748 14449
rect -1714 14415 -1675 14449
rect -1641 14415 -1601 14449
rect -1567 14415 -1527 14449
rect -1493 14415 -1453 14449
rect -1419 14415 -1379 14449
rect -1345 14415 -1305 14449
rect -1271 14415 -1231 14449
rect -1197 14415 -1157 14449
rect -1123 14415 -1083 14449
rect -1049 14415 -1009 14449
rect -975 14415 -935 14449
rect -901 14415 -861 14449
rect -827 14415 -787 14449
rect -753 14415 -713 14449
rect -679 14415 -647 14449
rect -2119 14377 -647 14415
rect -2119 14376 -1969 14377
rect -2119 14342 -2113 14376
rect -2079 14342 -2041 14376
rect -2007 14343 -1969 14376
rect -1935 14343 -1896 14377
rect -1862 14343 -1823 14377
rect -1789 14343 -1749 14377
rect -1715 14343 -1675 14377
rect -1641 14343 -1601 14377
rect -1567 14343 -1527 14377
rect -1493 14343 -1453 14377
rect -1419 14343 -1379 14377
rect -1345 14343 -1305 14377
rect -1271 14343 -1231 14377
rect -1197 14343 -1157 14377
rect -1123 14343 -1083 14377
rect -1049 14343 -1009 14377
rect -975 14343 -935 14377
rect -901 14343 -861 14377
rect -827 14343 -787 14377
rect -753 14343 -713 14377
rect -679 14343 -647 14377
rect -2007 14342 -647 14343
rect -2119 14337 -647 14342
rect -2119 14304 -1929 14337
rect -2119 14303 -1969 14304
rect -2119 14269 -2113 14303
rect -2079 14269 -2041 14303
rect -2007 14270 -1969 14303
rect -1935 14270 -1929 14304
rect -2007 14269 -1929 14270
rect -2119 14231 -1929 14269
rect -2119 14230 -1969 14231
rect -2119 14196 -2113 14230
rect -2079 14196 -2041 14230
rect -2007 14197 -1969 14230
rect -1935 14197 -1929 14231
rect -2007 14196 -1929 14197
rect -2119 14158 -1929 14196
rect -2119 14157 -1969 14158
rect -2119 14123 -2113 14157
rect -2079 14123 -2041 14157
rect -2007 14124 -1969 14157
rect -1935 14124 -1929 14158
rect -2007 14123 -1929 14124
rect -2119 14085 -1929 14123
rect -2119 14084 -1969 14085
rect -2119 14050 -2113 14084
rect -2079 14050 -2041 14084
rect -2007 14051 -1969 14084
rect -1935 14051 -1929 14085
rect -2007 14050 -1929 14051
rect -2119 14012 -1929 14050
rect -2119 14011 -1969 14012
rect -2119 13977 -2113 14011
rect -2079 13977 -2041 14011
rect -2007 13978 -1969 14011
rect -1935 13978 -1929 14012
rect -2007 13977 -1929 13978
rect -2119 13939 -1929 13977
rect -2119 13938 -1969 13939
rect -2119 13904 -2113 13938
rect -2079 13904 -2041 13938
rect -2007 13905 -1969 13938
rect -1935 13905 -1929 13939
rect -2007 13904 -1929 13905
rect -2119 13866 -1929 13904
rect -2119 13865 -1969 13866
rect -2119 13831 -2113 13865
rect -2079 13831 -2041 13865
rect -2007 13832 -1969 13865
rect -1935 13832 -1929 13866
rect -2007 13831 -1929 13832
rect -2119 13793 -1929 13831
rect -2119 13792 -1969 13793
rect -2119 13758 -2113 13792
rect -2079 13758 -2041 13792
rect -2007 13759 -1969 13792
rect -1935 13759 -1929 13793
rect -2007 13758 -1929 13759
rect -2119 13720 -1929 13758
rect -2119 13719 -1969 13720
rect -2119 13685 -2113 13719
rect -2079 13685 -2041 13719
rect -2007 13686 -1969 13719
rect -1935 13686 -1929 13720
rect -2007 13685 -1929 13686
rect -2119 13647 -1929 13685
rect -2119 13646 -1969 13647
rect -2119 13612 -2113 13646
rect -2079 13612 -2041 13646
rect -2007 13613 -1969 13646
rect -1935 13613 -1929 13647
rect -2007 13612 -1929 13613
rect -2119 13574 -1929 13612
rect -2119 13573 -1969 13574
rect -2119 13539 -2113 13573
rect -2079 13539 -2041 13573
rect -2007 13540 -1969 13573
rect -1935 13540 -1929 13574
rect -2007 13539 -1929 13540
rect -2119 13501 -1929 13539
rect -2119 13500 -1969 13501
rect -2119 13466 -2113 13500
rect -2079 13466 -2041 13500
rect -2007 13467 -1969 13500
rect -1935 13467 -1929 13501
rect -2007 13466 -1929 13467
rect -2119 13428 -1929 13466
rect -2119 13427 -1969 13428
rect -2119 13393 -2113 13427
rect -2079 13393 -2041 13427
rect -2007 13394 -1969 13427
rect -1935 13394 -1929 13428
rect -2007 13393 -1929 13394
rect -2119 13355 -1929 13393
rect -2119 13354 -1969 13355
rect -2119 13320 -2113 13354
rect -2079 13320 -2041 13354
rect -2007 13321 -1969 13354
rect -1935 13321 -1929 13355
rect -2007 13320 -1929 13321
rect -2119 13282 -1929 13320
rect -2119 13281 -1969 13282
rect -2119 13247 -2113 13281
rect -2079 13247 -2041 13281
rect -2007 13248 -1969 13281
rect -1935 13248 -1929 13282
rect -2007 13247 -1929 13248
rect -2119 13209 -1929 13247
rect -2119 13208 -1969 13209
rect -2119 13174 -2113 13208
rect -2079 13174 -2041 13208
rect -2007 13175 -1969 13208
rect -1935 13175 -1929 13209
rect -2007 13174 -1929 13175
rect -2119 13136 -1929 13174
rect -2119 13135 -1969 13136
rect -2119 13101 -2113 13135
rect -2079 13101 -2041 13135
rect -2007 13102 -1969 13135
rect -1935 13102 -1929 13136
rect -2007 13101 -1929 13102
rect -2119 13063 -1929 13101
rect -2119 13062 -1969 13063
rect -2119 13028 -2113 13062
rect -2079 13028 -2041 13062
rect -2007 13029 -1969 13062
rect -1935 13029 -1929 13063
rect -2007 13028 -1929 13029
rect -2119 12990 -1929 13028
rect -2119 12989 -1969 12990
rect -2119 12955 -2113 12989
rect -2079 12955 -2041 12989
rect -2007 12956 -1969 12989
rect -1935 12956 -1929 12990
rect -2007 12955 -1929 12956
rect -2119 12917 -1929 12955
rect -2119 12916 -1969 12917
rect -2119 12882 -2113 12916
rect -2079 12882 -2041 12916
rect -2007 12883 -1969 12916
rect -1935 12883 -1929 12917
rect -2007 12882 -1929 12883
rect -2119 12844 -1929 12882
rect -2119 12843 -1969 12844
rect -2119 12809 -2113 12843
rect -2079 12809 -2041 12843
rect -2007 12810 -1969 12843
rect -1935 12810 -1929 12844
rect -2007 12809 -1929 12810
rect -2119 12771 -1929 12809
rect -2119 12770 -1969 12771
rect -2119 12736 -2113 12770
rect -2079 12736 -2041 12770
rect -2007 12737 -1969 12770
rect -1935 12737 -1929 12771
rect -2007 12736 -1929 12737
rect -2119 12698 -1929 12736
rect -2119 12697 -1969 12698
rect -2119 12663 -2113 12697
rect -2079 12663 -2041 12697
rect -2007 12664 -1969 12697
rect -1935 12664 -1929 12698
rect -2007 12663 -1929 12664
rect -2119 12625 -1929 12663
rect -2119 12624 -1969 12625
rect -2119 12590 -2113 12624
rect -2079 12590 -2041 12624
rect -2007 12591 -1969 12624
rect -1935 12591 -1929 12625
rect -2007 12590 -1929 12591
rect -2119 12552 -1929 12590
rect -2119 12551 -1969 12552
rect -2119 12517 -2113 12551
rect -2079 12517 -2041 12551
rect -2007 12518 -1969 12551
rect -1935 12518 -1929 12552
rect -2007 12517 -1929 12518
rect -2119 12479 -1929 12517
rect -2119 12478 -1969 12479
rect -2119 12444 -2113 12478
rect -2079 12444 -2041 12478
rect -2007 12445 -1969 12478
rect -1935 12445 -1929 12479
rect -2007 12444 -1929 12445
rect -2119 12406 -1929 12444
rect -2119 12405 -1969 12406
rect -2119 12371 -2113 12405
rect -2079 12371 -2041 12405
rect -2007 12372 -1969 12405
rect -1935 12372 -1929 12406
rect -2007 12371 -1929 12372
rect -2119 12333 -1929 12371
rect -2119 12332 -1969 12333
rect -2119 12298 -2113 12332
rect -2079 12298 -2041 12332
rect -2007 12299 -1969 12332
rect -1935 12299 -1929 12333
rect -2007 12298 -1929 12299
rect -2119 12260 -1929 12298
rect -2119 12259 -1969 12260
rect -2119 12225 -2113 12259
rect -2079 12225 -2041 12259
rect -2007 12226 -1969 12259
rect -1935 12226 -1929 12260
rect -2007 12225 -1929 12226
rect -2119 12187 -1929 12225
rect -2119 12186 -1969 12187
rect -2119 7616 -2113 12186
rect -2007 12153 -1969 12186
rect -1935 12153 -1929 12187
rect -2007 12114 -1929 12153
rect -1935 7728 -1929 12114
rect -1795 14197 -1053 14203
rect -1795 14163 -1711 14197
rect -1677 14163 -1633 14197
rect -1599 14169 -1555 14197
rect -1521 14169 -1477 14197
rect -1443 14169 -1399 14197
rect -1521 14163 -1511 14169
rect -1443 14163 -1418 14169
rect -1365 14163 -1321 14197
rect -1287 14163 -1243 14197
rect -1209 14163 -1165 14197
rect -1131 14163 -1053 14197
rect -1795 14125 -1604 14163
rect -1552 14125 -1511 14163
rect -1459 14125 -1418 14163
rect -1366 14125 -1053 14163
rect -1795 14091 -1789 14125
rect -1755 14091 -1717 14125
rect -1683 14091 -1633 14125
rect -1521 14117 -1511 14125
rect -1443 14117 -1418 14125
rect -1599 14091 -1555 14117
rect -1521 14091 -1477 14117
rect -1443 14091 -1399 14117
rect -1365 14091 -1321 14125
rect -1287 14091 -1243 14125
rect -1209 14091 -1165 14125
rect -1795 14085 -1165 14091
rect -1795 14052 -1677 14085
rect -1795 14018 -1789 14052
rect -1755 14018 -1717 14052
rect -1683 14018 -1677 14052
rect -1795 13979 -1677 14018
rect -1171 14019 -1165 14085
rect -1059 14019 -1053 14125
rect -1795 13945 -1789 13979
rect -1755 13945 -1717 13979
rect -1683 13945 -1677 13979
rect -1795 13906 -1677 13945
rect -1795 13872 -1789 13906
rect -1755 13872 -1717 13906
rect -1683 13872 -1677 13906
rect -1795 13833 -1677 13872
rect -1795 13799 -1789 13833
rect -1755 13799 -1717 13833
rect -1683 13799 -1677 13833
rect -1795 13760 -1677 13799
rect -1795 13726 -1789 13760
rect -1755 13726 -1717 13760
rect -1683 13726 -1677 13760
rect -1795 13687 -1677 13726
rect -1795 13653 -1789 13687
rect -1755 13653 -1717 13687
rect -1683 13653 -1677 13687
rect -1795 13614 -1677 13653
rect -1795 13580 -1789 13614
rect -1755 13580 -1717 13614
rect -1683 13580 -1677 13614
rect -1795 13541 -1677 13580
rect -1795 13507 -1789 13541
rect -1755 13507 -1717 13541
rect -1683 13507 -1677 13541
rect -1795 13468 -1677 13507
rect -1795 7962 -1789 13468
rect -1683 8035 -1677 13468
rect -1525 12506 -1479 13982
rect -1525 12472 -1519 12506
rect -1485 12472 -1479 12506
rect -1525 12434 -1479 12472
rect -1525 12400 -1519 12434
rect -1485 12400 -1479 12434
rect -1603 12321 -1557 12333
rect -1603 12287 -1597 12321
rect -1563 12287 -1557 12321
rect -1603 12249 -1557 12287
rect -1603 12215 -1597 12249
rect -1563 12215 -1557 12249
rect -1603 12177 -1557 12215
rect -1603 12143 -1597 12177
rect -1563 12143 -1557 12177
rect -1603 12105 -1557 12143
rect -1603 12071 -1597 12105
rect -1563 12071 -1557 12105
rect -1603 12033 -1557 12071
rect -1603 11999 -1597 12033
rect -1563 11999 -1557 12033
tri -1606 11979 -1603 11982 se
rect -1603 11979 -1557 11999
tri -1557 11979 -1554 11982 sw
rect -1606 11973 -1554 11979
rect -1606 11909 -1554 11921
rect -1606 11855 -1597 11857
rect -1563 11855 -1554 11857
rect -1606 11845 -1554 11855
rect -1525 11853 -1479 12400
rect -1369 12506 -1323 13982
rect -1369 12472 -1363 12506
rect -1329 12472 -1323 12506
rect -1369 12434 -1323 12472
rect -1369 12400 -1363 12434
rect -1329 12400 -1323 12434
rect -1450 12321 -1398 12333
rect -1450 12311 -1441 12321
rect -1407 12311 -1398 12321
rect -1450 12249 -1398 12259
rect -1450 12247 -1441 12249
rect -1407 12247 -1398 12249
rect -1450 12183 -1398 12195
rect -1450 12125 -1398 12131
tri -1450 12122 -1447 12125 ne
rect -1447 12105 -1401 12125
tri -1401 12122 -1398 12125 nw
rect -1447 12071 -1441 12105
rect -1407 12071 -1401 12105
rect -1447 12033 -1401 12071
rect -1447 11999 -1441 12033
rect -1407 11999 -1401 12033
rect -1447 11961 -1401 11999
rect -1447 11927 -1441 11961
rect -1407 11927 -1401 11961
rect -1447 11889 -1401 11927
rect -1447 11855 -1441 11889
rect -1407 11855 -1401 11889
rect -1447 11817 -1401 11855
rect -1369 11853 -1323 12400
rect -1171 13980 -1053 14019
rect -1171 13946 -1165 13980
rect -1131 13946 -1093 13980
rect -1059 13946 -1053 13980
rect -1171 13907 -1053 13946
rect -1171 13873 -1165 13907
rect -1131 13873 -1093 13907
rect -1059 13873 -1053 13907
rect -1171 13834 -1053 13873
rect -1171 13800 -1165 13834
rect -1131 13800 -1093 13834
rect -1059 13800 -1053 13834
rect -1171 13761 -1053 13800
rect -1171 13727 -1165 13761
rect -1131 13727 -1093 13761
rect -1059 13727 -1053 13761
rect -1171 13688 -1053 13727
rect -1171 13654 -1165 13688
rect -1131 13654 -1093 13688
rect -1059 13654 -1053 13688
rect -1171 13615 -1053 13654
rect -1171 13581 -1165 13615
rect -1131 13581 -1093 13615
rect -1059 13581 -1053 13615
rect -1171 13542 -1053 13581
rect -1171 13508 -1165 13542
rect -1131 13508 -1093 13542
rect -1059 13508 -1053 13542
rect -1171 13469 -1053 13508
rect -1171 13435 -1165 13469
rect -1131 13435 -1093 13469
rect -1059 13435 -1053 13469
rect -1171 13396 -1053 13435
rect -1171 13362 -1165 13396
rect -1131 13362 -1093 13396
rect -1059 13362 -1053 13396
rect -1171 13323 -1053 13362
rect -1171 13289 -1165 13323
rect -1131 13289 -1093 13323
rect -1059 13289 -1053 13323
rect -1171 13250 -1053 13289
rect -1171 13216 -1165 13250
rect -1131 13216 -1093 13250
rect -1059 13216 -1053 13250
rect -1171 13177 -1053 13216
rect -1171 13143 -1165 13177
rect -1131 13143 -1093 13177
rect -1059 13143 -1053 13177
rect -1171 13104 -1053 13143
rect -1171 13070 -1165 13104
rect -1131 13070 -1093 13104
rect -1059 13070 -1053 13104
rect -1171 13031 -1053 13070
rect -1171 12997 -1165 13031
rect -1131 12997 -1093 13031
rect -1059 12997 -1053 13031
rect -1171 12958 -1053 12997
rect -1171 12924 -1165 12958
rect -1131 12924 -1093 12958
rect -1059 12924 -1053 12958
rect -1171 12885 -1053 12924
rect -1171 12851 -1165 12885
rect -1131 12851 -1093 12885
rect -1059 12851 -1053 12885
rect -1171 12812 -1053 12851
rect -1171 12778 -1165 12812
rect -1131 12778 -1093 12812
rect -1059 12778 -1053 12812
rect -1171 12739 -1053 12778
rect -1171 12705 -1165 12739
rect -1131 12705 -1093 12739
rect -1059 12705 -1053 12739
rect -1171 12666 -1053 12705
rect -1171 12632 -1165 12666
rect -1131 12632 -1093 12666
rect -1059 12632 -1053 12666
rect -1171 12568 -1053 12632
rect -1171 12534 -1165 12568
rect -1131 12534 -1093 12568
rect -1059 12534 -1053 12568
rect -1171 12495 -1053 12534
rect -1171 12461 -1165 12495
rect -1131 12461 -1093 12495
rect -1059 12461 -1053 12495
rect -1171 12422 -1053 12461
rect -1171 12388 -1165 12422
rect -1131 12388 -1093 12422
rect -1059 12388 -1053 12422
rect -1171 12349 -1053 12388
rect -1291 12321 -1245 12333
rect -1291 12287 -1285 12321
rect -1251 12287 -1245 12321
rect -1291 12249 -1245 12287
rect -1291 12215 -1285 12249
rect -1251 12215 -1245 12249
rect -1291 12177 -1245 12215
rect -1291 12143 -1285 12177
rect -1251 12143 -1245 12177
rect -1291 12105 -1245 12143
rect -1291 12071 -1285 12105
rect -1251 12071 -1245 12105
rect -1291 12033 -1245 12071
rect -1291 11999 -1285 12033
rect -1251 11999 -1245 12033
tri -1294 11979 -1291 11982 se
rect -1291 11979 -1245 11999
rect -1171 12315 -1165 12349
rect -1131 12315 -1093 12349
rect -1059 12315 -1053 12349
rect -1171 12276 -1053 12315
rect -1171 12242 -1165 12276
rect -1131 12242 -1093 12276
rect -1059 12242 -1053 12276
rect -1171 12203 -1053 12242
rect -1171 12169 -1165 12203
rect -1131 12169 -1093 12203
rect -1059 12169 -1053 12203
rect -1171 12130 -1053 12169
rect -1171 12096 -1165 12130
rect -1131 12096 -1093 12130
rect -1059 12096 -1053 12130
rect -1171 12057 -1053 12096
rect -1171 12023 -1165 12057
rect -1131 12023 -1093 12057
rect -1059 12023 -1053 12057
rect -1171 11984 -1053 12023
tri -1245 11979 -1242 11982 sw
rect -1294 11973 -1242 11979
rect -1294 11909 -1242 11921
rect -1294 11855 -1285 11857
rect -1251 11855 -1242 11857
rect -1606 11783 -1597 11793
rect -1563 11783 -1554 11793
rect -1606 11771 -1554 11783
rect -1525 11774 -1479 11797
rect -1525 11740 -1519 11774
rect -1485 11740 -1479 11774
rect -1447 11783 -1441 11817
rect -1407 11783 -1401 11817
rect -1294 11845 -1242 11855
rect -1447 11771 -1401 11783
rect -1369 11774 -1323 11797
rect -1525 11702 -1479 11740
rect -1606 11659 -1554 11671
rect -1606 11649 -1597 11659
rect -1563 11649 -1554 11659
rect -1606 11587 -1554 11597
rect -1606 11585 -1597 11587
rect -1563 11585 -1554 11587
rect -1606 11521 -1554 11533
rect -1606 11463 -1554 11469
tri -1606 11460 -1603 11463 ne
rect -1603 11443 -1557 11463
tri -1557 11460 -1554 11463 nw
rect -1525 11668 -1519 11702
rect -1485 11668 -1479 11702
rect -1369 11740 -1363 11774
rect -1329 11740 -1323 11774
rect -1294 11783 -1285 11793
rect -1251 11783 -1242 11793
rect -1294 11771 -1242 11783
rect -1171 11950 -1165 11984
rect -1131 11950 -1093 11984
rect -1059 11950 -1053 11984
rect -1171 11911 -1053 11950
rect -1171 11877 -1165 11911
rect -1131 11877 -1093 11911
rect -1059 11877 -1053 11911
rect -1171 11838 -1053 11877
rect -1171 11804 -1165 11838
rect -1131 11804 -1093 11838
rect -1059 11804 -1053 11838
rect -1369 11702 -1323 11740
rect -1603 11409 -1597 11443
rect -1563 11409 -1557 11443
rect -1603 11371 -1557 11409
rect -1603 11337 -1597 11371
rect -1563 11337 -1557 11371
rect -1603 11299 -1557 11337
rect -1603 11265 -1597 11299
rect -1563 11265 -1557 11299
rect -1603 11227 -1557 11265
rect -1603 11193 -1597 11227
rect -1563 11193 -1557 11227
rect -1603 11155 -1557 11193
rect -1603 11121 -1597 11155
rect -1563 11121 -1557 11155
rect -1603 11109 -1557 11121
rect -1525 11108 -1479 11668
rect -1447 11659 -1401 11671
rect -1447 11625 -1441 11659
rect -1407 11625 -1401 11659
rect -1447 11587 -1401 11625
rect -1447 11553 -1441 11587
rect -1407 11553 -1401 11587
rect -1447 11515 -1401 11553
rect -1447 11481 -1441 11515
rect -1407 11481 -1401 11515
rect -1447 11443 -1401 11481
rect -1447 11409 -1441 11443
rect -1407 11409 -1401 11443
rect -1447 11371 -1401 11409
rect -1447 11337 -1441 11371
rect -1407 11337 -1401 11371
rect -1447 11317 -1401 11337
rect -1369 11668 -1363 11702
rect -1329 11668 -1323 11702
rect -1171 11765 -1053 11804
rect -1171 11731 -1165 11765
rect -1131 11731 -1093 11765
rect -1059 11731 -1053 11765
rect -1171 11692 -1053 11731
rect -1450 11311 -1398 11317
rect -1450 11247 -1398 11259
rect -1450 11193 -1441 11195
rect -1407 11193 -1398 11195
rect -1450 11183 -1398 11193
rect -1450 11125 -1441 11131
rect -1447 11121 -1441 11125
rect -1407 11125 -1398 11131
rect -1407 11121 -1401 11125
rect -1447 11109 -1401 11121
rect -1369 11108 -1323 11668
rect -1294 11659 -1242 11671
rect -1294 11649 -1285 11659
rect -1251 11649 -1242 11659
rect -1294 11587 -1242 11597
rect -1294 11585 -1285 11587
rect -1251 11585 -1242 11587
rect -1294 11521 -1242 11533
rect -1294 11463 -1242 11469
tri -1294 11460 -1291 11463 ne
rect -1291 11443 -1245 11463
tri -1245 11460 -1242 11463 nw
rect -1171 11658 -1165 11692
rect -1131 11658 -1093 11692
rect -1059 11658 -1053 11692
rect -1171 11619 -1053 11658
rect -1171 11585 -1165 11619
rect -1131 11585 -1093 11619
rect -1059 11585 -1053 11619
rect -1171 11546 -1053 11585
rect -1171 11512 -1165 11546
rect -1131 11512 -1093 11546
rect -1059 11512 -1053 11546
rect -1171 11473 -1053 11512
rect -1291 11409 -1285 11443
rect -1251 11409 -1245 11443
rect -1291 11371 -1245 11409
rect -1291 11337 -1285 11371
rect -1251 11337 -1245 11371
rect -1291 11299 -1245 11337
rect -1291 11265 -1285 11299
rect -1251 11265 -1245 11299
rect -1291 11227 -1245 11265
rect -1291 11193 -1285 11227
rect -1251 11193 -1245 11227
rect -1291 11155 -1245 11193
rect -1291 11121 -1285 11155
rect -1251 11121 -1245 11155
rect -1291 11109 -1245 11121
rect -1171 11439 -1165 11473
rect -1131 11439 -1093 11473
rect -1059 11439 -1053 11473
rect -1171 11400 -1053 11439
rect -1171 11366 -1165 11400
rect -1131 11366 -1093 11400
rect -1059 11366 -1053 11400
rect -1171 11327 -1053 11366
rect -1171 11293 -1165 11327
rect -1131 11293 -1093 11327
rect -1059 11293 -1053 11327
rect -1171 11254 -1053 11293
rect -1171 11220 -1165 11254
rect -1131 11220 -1093 11254
rect -1059 11220 -1053 11254
rect -1171 11181 -1053 11220
rect -1171 11147 -1165 11181
rect -1131 11147 -1093 11181
rect -1059 11147 -1053 11181
rect -1171 11108 -1053 11147
rect -1171 11074 -1165 11108
rect -1131 11074 -1093 11108
rect -1059 11074 -1053 11108
rect -1525 11042 -1479 11065
rect -1525 11008 -1519 11042
rect -1485 11008 -1479 11042
rect -1525 10970 -1479 11008
rect -1525 10936 -1519 10970
rect -1485 10936 -1479 10970
rect -1603 10857 -1557 10869
rect -1603 10823 -1597 10857
rect -1563 10823 -1557 10857
rect -1603 10785 -1557 10823
rect -1603 10751 -1597 10785
rect -1563 10751 -1557 10785
rect -1603 10713 -1557 10751
rect -1603 10679 -1597 10713
rect -1563 10679 -1557 10713
rect -1603 10641 -1557 10679
rect -1603 10607 -1597 10641
rect -1563 10607 -1557 10641
rect -1603 10569 -1557 10607
rect -1603 10535 -1597 10569
rect -1563 10535 -1557 10569
rect -1603 10515 -1557 10535
rect -1606 10509 -1554 10515
rect -1606 10445 -1554 10457
rect -1606 10391 -1597 10393
rect -1563 10391 -1554 10393
rect -1606 10381 -1554 10391
rect -1606 10323 -1597 10329
rect -1603 10319 -1597 10323
rect -1563 10323 -1554 10329
rect -1563 10319 -1557 10323
rect -1603 10307 -1557 10319
rect -1525 9590 -1479 10936
rect -1369 11042 -1323 11065
rect -1369 11008 -1363 11042
rect -1329 11008 -1323 11042
rect -1369 10970 -1323 11008
rect -1369 10936 -1363 10970
rect -1329 10936 -1323 10970
rect -1450 10857 -1398 10869
rect -1450 10847 -1441 10857
rect -1407 10847 -1398 10857
rect -1450 10785 -1398 10795
rect -1450 10783 -1441 10785
rect -1407 10783 -1398 10785
rect -1450 10719 -1398 10731
rect -1450 10661 -1398 10667
tri -1450 10658 -1447 10661 ne
rect -1447 10641 -1401 10661
tri -1401 10658 -1398 10661 nw
rect -1447 10607 -1441 10641
rect -1407 10607 -1401 10641
rect -1447 10569 -1401 10607
rect -1447 10535 -1441 10569
rect -1407 10535 -1401 10569
rect -1447 10497 -1401 10535
rect -1447 10463 -1441 10497
rect -1407 10463 -1401 10497
rect -1447 10425 -1401 10463
rect -1447 10391 -1441 10425
rect -1407 10391 -1401 10425
rect -1447 10353 -1401 10391
rect -1447 10319 -1441 10353
rect -1407 10319 -1401 10353
rect -1447 10307 -1401 10319
rect -1369 9590 -1323 10936
rect -1171 11035 -1053 11074
rect -1171 11001 -1165 11035
rect -1131 11001 -1093 11035
rect -1059 11001 -1053 11035
rect -1171 10962 -1053 11001
rect -1171 10928 -1165 10962
rect -1131 10928 -1093 10962
rect -1059 10928 -1053 10962
rect -1171 10889 -1053 10928
rect -1291 10857 -1245 10869
rect -1291 10823 -1285 10857
rect -1251 10823 -1245 10857
rect -1291 10785 -1245 10823
rect -1291 10751 -1285 10785
rect -1251 10751 -1245 10785
rect -1291 10713 -1245 10751
rect -1291 10679 -1285 10713
rect -1251 10679 -1245 10713
rect -1291 10641 -1245 10679
rect -1291 10607 -1285 10641
rect -1251 10607 -1245 10641
rect -1291 10569 -1245 10607
rect -1291 10535 -1285 10569
rect -1251 10535 -1245 10569
rect -1291 10515 -1245 10535
rect -1171 10855 -1165 10889
rect -1131 10855 -1093 10889
rect -1059 10855 -1053 10889
rect -1171 10816 -1053 10855
rect -1171 10782 -1165 10816
rect -1131 10782 -1093 10816
rect -1059 10782 -1053 10816
rect -1171 10743 -1053 10782
rect -1171 10709 -1165 10743
rect -1131 10709 -1093 10743
rect -1059 10709 -1053 10743
rect -1171 10670 -1053 10709
rect -1171 10636 -1165 10670
rect -1131 10636 -1093 10670
rect -1059 10636 -1053 10670
rect -1171 10597 -1053 10636
rect -1171 10563 -1165 10597
rect -1131 10563 -1093 10597
rect -1059 10563 -1053 10597
rect -1171 10524 -1053 10563
rect -1294 10509 -1242 10515
rect -1294 10445 -1242 10457
rect -1294 10391 -1285 10393
rect -1251 10391 -1242 10393
rect -1294 10381 -1242 10391
rect -1294 10323 -1285 10329
rect -1291 10319 -1285 10323
rect -1251 10323 -1242 10329
rect -1171 10490 -1165 10524
rect -1131 10490 -1093 10524
rect -1059 10490 -1053 10524
rect -1171 10451 -1053 10490
rect -1171 10417 -1165 10451
rect -1131 10417 -1093 10451
rect -1059 10417 -1053 10451
rect -1171 10378 -1053 10417
rect -1171 10344 -1165 10378
rect -1131 10344 -1093 10378
rect -1059 10344 -1053 10378
rect -1251 10319 -1245 10323
rect -1291 10307 -1245 10319
rect -1171 10305 -1053 10344
rect -1171 10271 -1165 10305
rect -1131 10271 -1093 10305
rect -1059 10271 -1053 10305
rect -1171 10232 -1053 10271
rect -1171 10198 -1165 10232
rect -1131 10198 -1093 10232
rect -1059 10198 -1053 10232
rect -1171 10159 -1053 10198
rect -1171 10125 -1165 10159
rect -1131 10125 -1093 10159
rect -1059 10125 -1053 10159
rect -1171 10086 -1053 10125
rect -1171 10052 -1165 10086
rect -1131 10052 -1093 10086
rect -1059 10052 -1053 10086
rect -1171 10013 -1053 10052
tri -1677 8035 -1640 8072 sw
tri -1208 8035 -1171 8072 se
rect -1171 8035 -1165 10013
rect -1059 8035 -1053 10013
rect -1683 8002 -1640 8035
tri -1640 8002 -1607 8035 sw
tri -1241 8002 -1208 8035 se
rect -1208 8002 -1053 8035
rect -1683 7996 -1053 8002
rect -1683 7962 -1641 7996
rect -1607 7962 -1565 7996
rect -1531 7962 -1490 7996
rect -1456 7962 -1415 7996
rect -1381 7962 -1340 7996
rect -1306 7962 -1265 7996
rect -1231 7962 -1190 7996
rect -1156 7962 -1053 7996
rect -1795 7947 -1053 7962
rect -1795 7924 -1093 7947
rect -1795 7890 -1717 7924
rect -1683 7890 -1639 7924
rect -1605 7890 -1561 7924
rect -1527 7890 -1483 7924
rect -1449 7890 -1405 7924
rect -1371 7890 -1327 7924
rect -1293 7890 -1249 7924
rect -1215 7890 -1171 7924
rect -1137 7913 -1093 7924
rect -1059 7913 -1053 7947
rect -1137 7890 -1053 7913
rect -1795 7884 -1053 7890
rect -1935 7722 -647 7728
rect -1935 7688 -1895 7722
rect -1861 7688 -1821 7722
rect -1787 7688 -1747 7722
rect -1713 7688 -1673 7722
rect -1639 7688 -1599 7722
rect -1565 7688 -1525 7722
rect -1491 7688 -1451 7722
rect -1417 7688 -1377 7722
rect -1343 7688 -1303 7722
rect -1269 7688 -1229 7722
rect -1195 7688 -1155 7722
rect -1121 7688 -1081 7722
rect -1047 7688 -1007 7722
rect -973 7688 -933 7722
rect -899 7688 -859 7722
rect -825 7688 -786 7722
rect -752 7688 -713 7722
rect -679 7688 -647 7722
rect -2007 7650 -647 7688
rect -2007 7616 -1967 7650
rect -1933 7616 -1893 7650
rect -1859 7616 -1819 7650
rect -1785 7616 -1745 7650
rect -1711 7616 -1671 7650
rect -1637 7616 -1597 7650
rect -1563 7616 -1523 7650
rect -1489 7616 -1449 7650
rect -1415 7616 -1375 7650
rect -1341 7616 -1301 7650
rect -1267 7616 -1227 7650
rect -1193 7616 -1153 7650
rect -1119 7616 -1079 7650
rect -1045 7616 -1005 7650
rect -971 7616 -932 7650
rect -898 7616 -859 7650
rect -825 7616 -786 7650
rect -752 7616 -713 7650
rect -679 7616 -647 7650
rect -2119 7578 -647 7616
rect -2119 7544 -2041 7578
rect -2007 7544 -1967 7578
rect -1933 7544 -1893 7578
rect -1859 7544 -1819 7578
rect -1785 7544 -1745 7578
rect -1711 7544 -1671 7578
rect -1637 7544 -1597 7578
rect -1563 7544 -1523 7578
rect -1489 7544 -1449 7578
rect -1415 7544 -1375 7578
rect -1341 7544 -1301 7578
rect -1267 7544 -1227 7578
rect -1193 7544 -1153 7578
rect -1119 7544 -1079 7578
rect -1045 7544 -1005 7578
rect -971 7544 -932 7578
rect -898 7544 -859 7578
rect -825 7544 -786 7578
rect -752 7544 -713 7578
rect -679 7544 -647 7578
rect -2119 7538 -647 7544
rect -957 6223 -905 6229
tri -991 6117 -957 6151 se
rect -957 6148 -905 6171
tri -996 6112 -991 6117 se
rect -991 6112 -957 6117
tri -1586 6090 -1564 6112 se
rect -1564 6096 -957 6112
rect 21783 6171 21901 6177
rect 21835 6165 21847 6171
rect 19684 6123 19690 6126
rect -1564 6090 -905 6096
tri -1593 6083 -1586 6090 se
rect -1586 6083 -913 6090
tri -913 6083 -906 6090 nw
tri -1617 6059 -1593 6083 se
rect -1593 6060 -936 6083
tri -936 6060 -913 6083 nw
rect 19681 6077 19690 6123
rect 19684 6074 19690 6077
rect 19742 6074 19757 6126
rect 19809 6074 19824 6126
rect 19876 6074 19882 6126
rect 21899 6119 21901 6171
rect 21783 6104 21789 6119
rect 21895 6104 21901 6119
rect -1593 6059 -1534 6060
tri -1534 6059 -1533 6060 nw
tri -1636 6040 -1617 6059 se
rect -1617 6040 -1553 6059
tri -1553 6040 -1534 6059 nw
rect 21835 6052 21847 6059
rect 21899 6052 21901 6104
rect 21783 6047 21901 6052
rect 21783 6046 21899 6047
rect -1636 5832 -1584 6040
tri -1584 6009 -1553 6040 nw
rect -1636 5757 -1584 5780
rect -1636 5699 -1584 5705
rect 20005 5526 21890 5532
rect 19684 5496 19690 5499
rect 19681 5450 19690 5496
rect 19684 5447 19690 5450
rect 19742 5447 19754 5499
rect 19806 5447 19812 5499
rect 20005 5420 21772 5526
rect 21878 5420 21890 5526
rect 20005 5414 21890 5420
rect 3023 5079 3029 5131
rect 3081 5079 3095 5131
rect 3147 5079 3161 5131
rect 3213 5079 3227 5131
rect 3279 5079 3293 5131
rect 3345 5079 3358 5131
rect 3410 5079 3423 5131
rect 3475 5079 3488 5131
rect 3540 5079 3553 5131
rect 3605 5079 3618 5131
rect 3670 5079 3683 5131
rect 3735 5079 3748 5131
rect 3800 5079 3813 5131
rect 3865 5079 3878 5131
rect 3930 5079 3943 5131
rect 3995 5079 4008 5131
rect 4060 5079 4073 5131
rect 4125 5079 4138 5131
rect 4190 5079 4203 5131
rect 4255 5079 4268 5131
rect 4320 5079 4326 5131
rect 3023 5015 4326 5079
rect 3023 4963 3029 5015
rect 3081 4963 3095 5015
rect 3147 4963 3161 5015
rect 3213 4963 3227 5015
rect 3279 4963 3293 5015
rect 3345 4963 3358 5015
rect 3410 4963 3423 5015
rect 3475 4963 3488 5015
rect 3540 4963 3553 5015
rect 3605 4963 3618 5015
rect 3670 4963 3683 5015
rect 3735 4963 3748 5015
rect 3800 4963 3813 5015
rect 3865 4963 3878 5015
rect 3930 4963 3943 5015
rect 3995 4963 4008 5015
rect 4060 4963 4073 5015
rect 4125 4963 4138 5015
rect 4190 4963 4203 5015
rect 4255 4963 4268 5015
rect 4320 4963 4326 5015
rect 8554 5079 8560 5131
rect 8612 5079 8627 5131
rect 8679 5079 8694 5131
rect 8746 5079 8761 5131
rect 8813 5079 8828 5131
rect 8880 5079 8895 5131
rect 8947 5079 8962 5131
rect 9014 5079 9028 5131
rect 9080 5079 9094 5131
rect 9146 5079 9160 5131
rect 9212 5079 9226 5131
rect 9278 5079 9292 5131
rect 9344 5079 9358 5131
rect 9410 5079 9424 5131
rect 9476 5079 9490 5131
rect 9542 5079 9556 5131
rect 9608 5079 9614 5131
rect 8554 5015 9614 5079
rect 8554 4963 8560 5015
rect 8612 4963 8627 5015
rect 8679 4963 8694 5015
rect 8746 4963 8761 5015
rect 8813 4963 8828 5015
rect 8880 4963 8895 5015
rect 8947 4963 8962 5015
rect 9014 4963 9028 5015
rect 9080 4963 9094 5015
rect 9146 4963 9160 5015
rect 9212 4963 9226 5015
rect 9278 4963 9292 5015
rect 9344 4963 9358 5015
rect 9410 4963 9424 5015
rect 9476 4963 9490 5015
rect 9542 4963 9556 5015
rect 9608 4963 9614 5015
rect 11008 5079 11014 5131
rect 11066 5079 11082 5131
rect 11134 5079 11150 5131
rect 11202 5079 11217 5131
rect 11269 5079 11275 5131
rect 11008 5015 11275 5079
rect 11008 4963 11014 5015
rect 11066 4963 11082 5015
rect 11134 4963 11150 5015
rect 11202 4963 11217 5015
rect 11269 4963 11275 5015
rect 15043 5079 15049 5131
rect 15101 5079 15118 5131
rect 15170 5079 15187 5131
rect 15239 5079 15255 5131
rect 15307 5079 15323 5131
rect 15375 5079 15391 5131
rect 15443 5079 15459 5131
rect 15511 5079 15527 5131
rect 15579 5079 15595 5131
rect 15647 5079 15663 5131
rect 15715 5079 15731 5131
rect 15783 5079 15799 5131
rect 15851 5079 15867 5131
rect 15919 5079 15925 5131
rect 15043 5015 15925 5079
rect 15043 4963 15049 5015
rect 15101 4963 15118 5015
rect 15170 4963 15187 5015
rect 15239 4963 15255 5015
rect 15307 4963 15323 5015
rect 15375 4963 15391 5015
rect 15443 4963 15459 5015
rect 15511 4963 15527 5015
rect 15579 4963 15595 5015
rect 15647 4963 15663 5015
rect 15715 4963 15731 5015
rect 15783 4963 15799 5015
rect 15851 4963 15867 5015
rect 15919 4963 15925 5015
rect 16882 5079 16888 5131
rect 16940 5079 16957 5131
rect 17009 5079 17026 5131
rect 17078 5079 17094 5131
rect 17146 5079 17162 5131
rect 17214 5079 17230 5131
rect 17282 5079 17298 5131
rect 17350 5079 17366 5131
rect 17418 5079 17434 5131
rect 17486 5079 17502 5131
rect 17554 5079 17570 5131
rect 17622 5079 17638 5131
rect 17690 5079 17706 5131
rect 17758 5079 17764 5131
rect 16882 5015 17764 5079
rect 16882 4963 16888 5015
rect 16940 4963 16957 5015
rect 17009 4963 17026 5015
rect 17078 4963 17094 5015
rect 17146 4963 17162 5015
rect 17214 4963 17230 5015
rect 17282 4963 17298 5015
rect 17350 4963 17366 5015
rect 17418 4963 17434 5015
rect 17486 4963 17502 5015
rect 17554 4963 17570 5015
rect 17622 4963 17638 5015
rect 17690 4963 17706 5015
rect 17758 4963 17764 5015
rect 19665 5079 19671 5131
rect 19723 5079 19762 5131
rect 19814 5079 19820 5131
rect 19665 5015 19820 5079
rect 19665 4963 19671 5015
rect 19723 4963 19762 5015
rect 19814 4963 19820 5015
rect 3625 4706 3631 4758
rect 3683 4706 3698 4758
rect 3750 4706 3765 4758
rect 3817 4706 3832 4758
rect 3884 4706 3899 4758
rect 3951 4706 3966 4758
rect 4018 4706 4033 4758
rect 4085 4706 4099 4758
rect 4151 4706 4165 4758
rect 4217 4706 4223 4758
rect 3625 4694 4223 4706
rect 3625 4642 3631 4694
rect 3683 4642 3698 4694
rect 3750 4642 3765 4694
rect 3817 4642 3832 4694
rect 3884 4642 3899 4694
rect 3951 4642 3966 4694
rect 4018 4642 4033 4694
rect 4085 4642 4099 4694
rect 4151 4642 4165 4694
rect 4217 4642 4223 4694
rect 3625 4630 4223 4642
rect 3625 4578 3631 4630
rect 3683 4578 3698 4630
rect 3750 4578 3765 4630
rect 3817 4578 3832 4630
rect 3884 4578 3899 4630
rect 3951 4578 3966 4630
rect 4018 4578 4033 4630
rect 4085 4578 4099 4630
rect 4151 4578 4165 4630
rect 4217 4578 4223 4630
rect -1176 4526 -1124 4532
rect -1176 4462 -1124 4474
rect -1176 4404 -1124 4410
rect -1084 4406 -1078 4458
rect -1026 4406 -1014 4458
rect -962 4406 -956 4458
tri 19842 4376 19844 4378 se
rect 19844 4372 19960 4378
tri 19960 4376 19962 4378 sw
rect 643 4295 649 4347
rect 701 4295 725 4347
rect 777 4295 800 4347
rect 852 4295 858 4347
rect 643 4267 858 4295
rect 643 4215 649 4267
rect 701 4215 725 4267
rect 777 4215 800 4267
rect 852 4215 858 4267
rect 6012 4295 6018 4347
rect 6070 4295 6085 4347
rect 6137 4295 6152 4347
rect 6204 4295 6219 4347
rect 6271 4295 6286 4347
rect 6338 4295 6353 4347
rect 6405 4295 6411 4347
rect 6012 4267 6411 4295
rect 6012 4215 6018 4267
rect 6070 4215 6085 4267
rect 6137 4215 6152 4267
rect 6204 4215 6219 4267
rect 6271 4215 6286 4267
rect 6338 4215 6353 4267
rect 6405 4215 6411 4267
rect 6943 4295 6949 4347
rect 7001 4295 7016 4347
rect 7068 4295 7083 4347
rect 7135 4295 7150 4347
rect 7202 4295 7217 4347
rect 7269 4295 7284 4347
rect 7336 4295 7342 4347
rect 6943 4267 7342 4295
rect 6943 4215 6949 4267
rect 7001 4215 7016 4267
rect 7068 4215 7083 4267
rect 7135 4215 7150 4267
rect 7202 4215 7217 4267
rect 7269 4215 7284 4267
rect 7336 4215 7342 4267
rect 12496 4295 12502 4347
rect 12554 4295 12569 4347
rect 12621 4295 12636 4347
rect 12688 4295 12703 4347
rect 12755 4295 12770 4347
rect 12822 4295 12837 4347
rect 12889 4295 12895 4347
rect 12496 4267 12895 4295
rect 12496 4215 12502 4267
rect 12554 4215 12569 4267
rect 12621 4215 12636 4267
rect 12688 4215 12703 4267
rect 12755 4215 12770 4267
rect 12822 4215 12837 4267
rect 12889 4215 12895 4267
rect 13427 4295 13433 4347
rect 13485 4295 13500 4347
rect 13552 4295 13567 4347
rect 13619 4295 13634 4347
rect 13686 4295 13701 4347
rect 13753 4295 13768 4347
rect 13820 4295 13826 4347
rect 13427 4267 13826 4295
rect 13427 4215 13433 4267
rect 13485 4215 13500 4267
rect 13552 4215 13567 4267
rect 13619 4215 13634 4267
rect 13686 4215 13701 4267
rect 13753 4215 13768 4267
rect 13820 4215 13826 4267
rect 19061 4295 19067 4347
rect 19119 4295 19152 4347
rect 19204 4295 19237 4347
rect 19289 4295 19321 4347
rect 19373 4295 19379 4347
rect 19061 4267 19379 4295
rect 19061 4215 19067 4267
rect 19119 4215 19152 4267
rect 19204 4215 19237 4267
rect 19289 4215 19321 4267
rect 19373 4215 19379 4267
rect 19844 4186 19960 4192
rect -630 3333 -624 3385
rect -572 3333 -560 3385
rect -508 3380 -502 3385
rect -508 3334 -12 3380
rect -508 3333 -502 3334
rect -310 3017 20058 3023
rect -258 2991 20058 3017
rect -310 2953 -258 2965
rect -897 2895 -799 2926
tri -799 2895 -768 2926 sw
rect -310 2895 -258 2901
rect -52 2928 644 2959
rect 696 2928 728 2959
rect 780 2928 812 2959
rect 864 2928 895 2959
rect 947 2928 6018 2959
rect 6070 2928 6085 2959
rect 6137 2928 6152 2959
rect -897 2894 -768 2895
tri -768 2894 -767 2895 sw
rect -52 2894 -20 2928
rect 14 2894 53 2928
rect 87 2894 126 2928
rect 160 2894 199 2928
rect 233 2894 272 2928
rect 306 2894 345 2928
rect 379 2894 418 2928
rect 452 2894 491 2928
rect 525 2894 564 2928
rect 598 2894 637 2928
rect 696 2907 710 2928
rect 780 2907 783 2928
rect 890 2907 895 2928
rect 671 2894 710 2907
rect 744 2894 783 2907
rect 817 2894 856 2907
rect 890 2894 929 2907
rect 963 2894 1002 2928
rect 1036 2894 1075 2928
rect 1109 2894 1148 2928
rect 1182 2894 1221 2928
rect 1255 2894 1294 2928
rect 1328 2894 1367 2928
rect 1401 2894 1440 2928
rect 1474 2894 1513 2928
rect 1547 2894 1586 2928
rect 1620 2894 1659 2928
rect 1693 2894 1732 2928
rect 1766 2894 1805 2928
rect 1839 2894 1878 2928
rect 1912 2894 1951 2928
rect 1985 2894 2024 2928
rect 2058 2894 2097 2928
rect 2131 2894 2170 2928
rect 2204 2894 2243 2928
rect 2277 2894 2316 2928
rect 2350 2894 2389 2928
rect 2423 2894 2462 2928
rect 2496 2894 2535 2928
rect 2569 2894 2608 2928
rect 2642 2894 2681 2928
rect 2715 2894 2754 2928
rect 2788 2894 2827 2928
rect 2861 2894 2900 2928
rect 2934 2894 2973 2928
rect 3007 2894 3046 2928
rect 3080 2894 3119 2928
rect 3153 2894 3192 2928
rect 3226 2894 3265 2928
rect 3299 2894 3338 2928
rect 3372 2894 3411 2928
rect 3445 2894 3483 2928
rect 3517 2894 3555 2928
rect 3589 2894 3627 2928
rect 3661 2894 3699 2928
rect 3733 2894 3771 2928
rect 3805 2894 3843 2928
rect 3877 2894 3915 2928
rect 3949 2894 3987 2928
rect 4021 2894 4059 2928
rect 4093 2894 4131 2928
rect 4165 2894 4203 2928
rect 4237 2894 4275 2928
rect 4309 2894 4347 2928
rect 4381 2894 4419 2928
rect 4453 2894 4491 2928
rect 4525 2894 4563 2928
rect 4597 2894 4635 2928
rect 4669 2894 4707 2928
rect 4741 2894 4779 2928
rect 4813 2894 4851 2928
rect 4885 2894 4923 2928
rect 4957 2894 4995 2928
rect 5029 2894 5067 2928
rect 5101 2894 5139 2928
rect 5173 2894 5211 2928
rect 5245 2894 5283 2928
rect 5317 2894 5355 2928
rect 5389 2894 5427 2928
rect 5461 2894 5499 2928
rect 5533 2894 5571 2928
rect 5605 2894 5643 2928
rect 5677 2894 5715 2928
rect 5749 2894 5787 2928
rect 5821 2894 5859 2928
rect 5893 2894 5931 2928
rect 5965 2894 6003 2928
rect 6070 2907 6075 2928
rect 6137 2907 6147 2928
rect 6204 2907 6219 2959
rect 6271 2907 6286 2959
rect 6338 2907 6353 2959
rect 6405 2928 6949 2959
rect 7001 2928 7016 2959
rect 6405 2907 6435 2928
rect 6037 2894 6075 2907
rect 6109 2894 6147 2907
rect 6181 2894 6219 2907
rect 6253 2894 6291 2907
rect 6325 2894 6363 2907
rect 6397 2894 6435 2907
rect 6469 2894 6507 2928
rect 6541 2894 6579 2928
rect 6613 2894 6651 2928
rect 6685 2894 6723 2928
rect 6757 2894 6795 2928
rect 6829 2894 6867 2928
rect 6901 2894 6939 2928
rect 7001 2907 7011 2928
rect 7068 2907 7083 2959
rect 7135 2907 7150 2959
rect 7202 2907 7217 2959
rect 7269 2907 7284 2959
rect 7336 2928 12502 2959
rect 12554 2928 12569 2959
rect 12621 2928 12636 2959
rect 12688 2928 12703 2959
rect 7336 2907 7371 2928
rect 6973 2894 7011 2907
rect 7045 2894 7083 2907
rect 7117 2894 7155 2907
rect 7189 2894 7227 2907
rect 7261 2894 7299 2907
rect 7333 2894 7371 2907
rect 7405 2894 7443 2928
rect 7477 2894 7515 2928
rect 7549 2894 7587 2928
rect 7621 2894 7659 2928
rect 7693 2894 7731 2928
rect 7765 2894 7803 2928
rect 7837 2894 7875 2928
rect 7909 2894 7947 2928
rect 7981 2894 8019 2928
rect 8053 2894 8091 2928
rect 8125 2894 8163 2928
rect 8197 2894 8235 2928
rect 8269 2894 8307 2928
rect 8341 2894 8379 2928
rect 8413 2894 8451 2928
rect 8485 2894 8523 2928
rect 8557 2894 8595 2928
rect 8629 2894 8667 2928
rect 8701 2894 8739 2928
rect 8773 2894 8811 2928
rect 8845 2894 8883 2928
rect 8917 2894 8955 2928
rect 8989 2894 9027 2928
rect 9061 2894 9099 2928
rect 9133 2894 9171 2928
rect 9205 2894 9243 2928
rect 9277 2894 9315 2928
rect 9349 2894 9387 2928
rect 9421 2894 9459 2928
rect 9493 2894 9531 2928
rect 9565 2894 9603 2928
rect 9637 2894 9675 2928
rect 9709 2894 9747 2928
rect 9781 2894 9819 2928
rect 9853 2894 9891 2928
rect 9925 2894 9963 2928
rect 9997 2894 10035 2928
rect 10069 2894 10107 2928
rect 10141 2894 10179 2928
rect 10213 2894 10251 2928
rect 10285 2894 10323 2928
rect 10357 2894 10395 2928
rect 10429 2894 10467 2928
rect 10501 2894 10539 2928
rect 10573 2894 10611 2928
rect 10645 2894 10683 2928
rect 10717 2894 10755 2928
rect 10789 2894 10827 2928
rect 10861 2894 10899 2928
rect 10933 2894 10971 2928
rect 11005 2894 11043 2928
rect 11077 2894 11115 2928
rect 11149 2894 11187 2928
rect 11221 2894 11259 2928
rect 11293 2894 11331 2928
rect 11365 2894 11403 2928
rect 11437 2894 11475 2928
rect 11509 2894 11547 2928
rect 11581 2894 11619 2928
rect 11653 2894 11691 2928
rect 11725 2894 11763 2928
rect 11797 2894 11835 2928
rect 11869 2894 11907 2928
rect 11941 2894 11979 2928
rect 12013 2894 12051 2928
rect 12085 2894 12123 2928
rect 12157 2894 12195 2928
rect 12229 2894 12267 2928
rect 12301 2894 12339 2928
rect 12373 2894 12411 2928
rect 12445 2894 12483 2928
rect 12554 2907 12555 2928
rect 12621 2907 12627 2928
rect 12688 2907 12699 2928
rect 12755 2907 12770 2959
rect 12822 2907 12837 2959
rect 12889 2928 13433 2959
rect 13485 2928 13500 2959
rect 13552 2928 13567 2959
rect 12889 2907 12915 2928
rect 12517 2894 12555 2907
rect 12589 2894 12627 2907
rect 12661 2894 12699 2907
rect 12733 2894 12771 2907
rect 12805 2894 12843 2907
rect 12877 2894 12915 2907
rect 12949 2894 12987 2928
rect 13021 2894 13059 2928
rect 13093 2894 13131 2928
rect 13165 2894 13203 2928
rect 13237 2894 13275 2928
rect 13309 2894 13347 2928
rect 13381 2894 13419 2928
rect 13485 2907 13491 2928
rect 13552 2907 13563 2928
rect 13619 2907 13634 2959
rect 13686 2907 13701 2959
rect 13753 2907 13768 2959
rect 13820 2928 19071 2959
rect 19123 2928 19155 2959
rect 19207 2928 19238 2959
rect 13820 2907 13851 2928
rect 13453 2894 13491 2907
rect 13525 2894 13563 2907
rect 13597 2894 13635 2907
rect 13669 2894 13707 2907
rect 13741 2894 13779 2907
rect 13813 2894 13851 2907
rect 13885 2894 13923 2928
rect 13957 2894 13995 2928
rect 14029 2894 14067 2928
rect 14101 2894 14139 2928
rect 14173 2894 14211 2928
rect 14245 2894 14283 2928
rect 14317 2894 14355 2928
rect 14389 2894 14427 2928
rect 14461 2894 14499 2928
rect 14533 2894 14571 2928
rect 14605 2894 14643 2928
rect 14677 2894 14715 2928
rect 14749 2894 14787 2928
rect 14821 2894 14859 2928
rect 14893 2894 14931 2928
rect 14965 2894 15003 2928
rect 15037 2894 15075 2928
rect 15109 2894 15147 2928
rect 15181 2894 15219 2928
rect 15253 2894 15291 2928
rect 15325 2894 15363 2928
rect 15397 2894 15435 2928
rect 15469 2894 15507 2928
rect 15541 2894 15579 2928
rect 15613 2894 15651 2928
rect 15685 2894 15723 2928
rect 15757 2894 15795 2928
rect 15829 2894 15867 2928
rect 15901 2894 15939 2928
rect 15973 2894 16011 2928
rect 16045 2894 16083 2928
rect 16117 2894 16155 2928
rect 16189 2894 16227 2928
rect 16261 2894 16299 2928
rect 16333 2894 16371 2928
rect 16405 2894 16443 2928
rect 16477 2894 16515 2928
rect 16549 2894 16587 2928
rect 16621 2894 16659 2928
rect 16693 2894 16731 2928
rect 16765 2894 16803 2928
rect 16837 2894 16875 2928
rect 16909 2894 16947 2928
rect 16981 2894 17019 2928
rect 17053 2894 17091 2928
rect 17125 2894 17163 2928
rect 17197 2894 17235 2928
rect 17269 2894 17307 2928
rect 17341 2894 17379 2928
rect 17413 2894 17451 2928
rect 17485 2894 17523 2928
rect 17557 2894 17595 2928
rect 17629 2894 17667 2928
rect 17701 2894 17739 2928
rect 17773 2894 17811 2928
rect 17845 2894 17883 2928
rect 17917 2894 17955 2928
rect 17989 2894 18027 2928
rect 18061 2894 18099 2928
rect 18133 2894 18171 2928
rect 18205 2894 18243 2928
rect 18277 2894 18315 2928
rect 18349 2894 18387 2928
rect 18421 2894 18459 2928
rect 18493 2894 18531 2928
rect 18565 2894 18603 2928
rect 18637 2894 18675 2928
rect 18709 2894 18747 2928
rect 18781 2894 18819 2928
rect 18853 2894 18891 2928
rect 18925 2894 18963 2928
rect 18997 2894 19035 2928
rect 19069 2907 19071 2928
rect 19141 2907 19155 2928
rect 19213 2907 19238 2928
rect 19290 2907 19321 2959
rect 19373 2951 19939 2959
tri 19939 2951 19947 2959 sw
rect 19373 2928 19947 2951
rect 19373 2907 19395 2928
rect 19069 2894 19107 2907
rect 19141 2894 19179 2907
rect 19213 2894 19251 2907
rect 19285 2894 19323 2907
rect 19357 2894 19395 2907
rect 19429 2894 19467 2928
rect 19501 2894 19539 2928
rect 19573 2894 19611 2928
rect 19645 2894 19683 2928
rect 19717 2894 19755 2928
rect 19789 2927 19947 2928
tri 19947 2927 19971 2951 sw
rect 19789 2894 19971 2927
rect -897 2883 -767 2894
tri -767 2883 -756 2894 sw
rect -897 2880 -414 2883
tri -835 2873 -828 2880 ne
rect -828 2877 -414 2880
rect -828 2873 -466 2877
tri -828 2845 -800 2873 ne
rect -800 2845 -466 2873
rect -1647 2829 -1289 2835
rect -1647 2823 -1360 2829
rect -1308 2823 -1289 2829
rect -1647 2789 -1641 2823
rect -1607 2789 -1360 2823
rect -1295 2789 -1289 2823
rect -1647 2777 -1360 2789
rect -1308 2777 -1289 2789
rect -1647 2759 -1289 2777
rect -1647 2750 -1360 2759
rect -1308 2750 -1289 2759
rect -1647 2716 -1641 2750
rect -1607 2716 -1360 2750
rect -1295 2716 -1289 2750
rect -1647 2707 -1360 2716
rect -1308 2707 -1289 2716
rect -1647 2688 -1289 2707
rect -1647 2676 -1360 2688
rect -1308 2676 -1289 2688
rect -1737 2645 -1685 2651
rect -1647 2642 -1641 2676
rect -1607 2642 -1360 2676
rect -1295 2642 -1289 2676
rect -1647 2636 -1360 2642
rect -1308 2636 -1289 2642
rect -1647 2630 -1289 2636
rect -1204 2829 -846 2835
rect -1204 2823 -1084 2829
rect -1204 2789 -1198 2823
rect -1164 2789 -1084 2823
rect -1204 2777 -1084 2789
rect -1032 2823 -846 2829
rect -1032 2789 -886 2823
rect -852 2789 -846 2823
rect -1032 2777 -846 2789
rect -1204 2759 -846 2777
rect -1204 2750 -1084 2759
rect -1204 2716 -1198 2750
rect -1164 2716 -1084 2750
rect -1204 2707 -1084 2716
rect -1032 2750 -846 2759
rect -466 2813 -414 2825
rect -466 2755 -414 2761
rect -52 2879 19971 2894
rect -52 2827 644 2879
rect 696 2827 728 2879
rect 780 2827 812 2879
rect 864 2827 895 2879
rect 947 2827 6018 2879
rect 6070 2827 6085 2879
rect 6137 2827 6152 2879
rect 6204 2827 6219 2879
rect 6271 2827 6286 2879
rect 6338 2827 6353 2879
rect 6405 2827 6949 2879
rect 7001 2827 7016 2879
rect 7068 2827 7083 2879
rect 7135 2827 7150 2879
rect 7202 2827 7217 2879
rect 7269 2827 7284 2879
rect 7336 2827 12502 2879
rect 12554 2827 12569 2879
rect 12621 2827 12636 2879
rect 12688 2827 12703 2879
rect 12755 2827 12770 2879
rect 12822 2827 12837 2879
rect 12889 2827 13433 2879
rect 13485 2827 13500 2879
rect 13552 2827 13567 2879
rect 13619 2827 13634 2879
rect 13686 2827 13701 2879
rect 13753 2827 13768 2879
rect 13820 2827 19071 2879
rect 19123 2827 19155 2879
rect 19207 2827 19238 2879
rect 19290 2827 19321 2879
rect 19373 2873 19971 2879
rect 19373 2839 19882 2873
rect 19916 2839 19971 2873
rect 19373 2827 19971 2839
rect -52 2818 187 2827
tri 187 2818 196 2827 nw
tri 19729 2818 19738 2827 ne
rect 19738 2818 19971 2827
rect -52 2800 169 2818
tri 169 2800 187 2818 nw
tri 19738 2800 19756 2818 ne
rect 19756 2800 19971 2818
rect -52 2794 135 2800
rect -52 2760 -46 2794
rect -12 2760 42 2794
rect 76 2766 135 2794
tri 135 2766 169 2800 nw
tri 19756 2766 19790 2800 ne
rect 19790 2766 19882 2800
rect 19916 2766 19971 2800
rect 76 2760 107 2766
rect -1032 2716 -886 2750
rect -852 2716 -846 2750
rect -1032 2707 -846 2716
rect -1204 2688 -846 2707
rect -1204 2676 -1084 2688
rect -1204 2642 -1198 2676
rect -1164 2642 -1084 2676
rect -1204 2636 -1084 2642
rect -1032 2676 -846 2688
rect -1032 2642 -886 2676
rect -852 2642 -846 2676
rect -1032 2636 -846 2642
rect -1204 2630 -846 2636
rect -52 2738 107 2760
tri 107 2738 135 2766 nw
tri 19790 2738 19818 2766 ne
rect 19818 2738 19971 2766
rect -52 2727 96 2738
tri 96 2727 107 2738 nw
rect -52 2721 82 2727
rect -52 2687 -46 2721
rect -12 2687 42 2721
rect 76 2687 82 2721
tri 82 2713 96 2727 nw
rect -52 2648 82 2687
rect -1737 2581 -1685 2593
rect -52 2614 -46 2648
rect -12 2614 42 2648
rect 76 2614 82 2648
rect -52 2575 82 2614
rect -1685 2567 -170 2573
rect -1685 2561 -222 2567
rect -1685 2529 -1485 2561
rect -1737 2527 -1485 2529
rect -1451 2527 -222 2561
rect -1737 2523 -222 2527
rect -1491 2489 -1445 2523
tri -253 2508 -238 2523 ne
rect -238 2515 -222 2523
rect -238 2508 -170 2515
tri -238 2502 -232 2508 ne
rect -232 2503 -170 2508
rect -232 2502 -222 2503
tri -232 2492 -222 2502 ne
rect -1491 2455 -1485 2489
rect -1451 2455 -1445 2489
rect -1491 2443 -1445 2455
rect -1048 2475 -1002 2487
rect -1048 2441 -1042 2475
rect -1008 2441 -1002 2475
rect -1048 2406 -1002 2441
rect -310 2461 -258 2467
rect -222 2444 -170 2451
rect -52 2541 -46 2575
rect -12 2541 42 2575
rect 76 2541 82 2575
rect 638 2686 644 2738
rect 696 2686 728 2738
rect 780 2686 812 2738
rect 864 2686 895 2738
rect 947 2686 953 2738
rect 638 2674 953 2686
rect 638 2622 644 2674
rect 696 2622 728 2674
rect 780 2622 812 2674
rect 864 2622 895 2674
rect 947 2622 953 2674
rect 638 2610 953 2622
rect 638 2558 644 2610
rect 696 2558 728 2610
rect 780 2558 812 2610
rect 864 2558 895 2610
rect 947 2558 953 2610
rect 6012 2686 6018 2738
rect 6070 2686 6085 2738
rect 6137 2686 6152 2738
rect 6204 2686 6219 2738
rect 6271 2686 6286 2738
rect 6338 2686 6353 2738
rect 6405 2686 6411 2738
rect 6012 2674 6411 2686
rect 6012 2622 6018 2674
rect 6070 2622 6085 2674
rect 6137 2622 6152 2674
rect 6204 2622 6219 2674
rect 6271 2622 6286 2674
rect 6338 2622 6353 2674
rect 6405 2622 6411 2674
rect 6012 2610 6411 2622
rect 6012 2558 6018 2610
rect 6070 2558 6085 2610
rect 6137 2558 6152 2610
rect 6204 2558 6219 2610
rect 6271 2558 6286 2610
rect 6338 2558 6353 2610
rect 6405 2558 6411 2610
rect 6943 2686 6949 2738
rect 7001 2686 7016 2738
rect 7068 2686 7083 2738
rect 7135 2686 7150 2738
rect 7202 2686 7217 2738
rect 7269 2686 7284 2738
rect 7336 2686 7342 2738
rect 6943 2674 7342 2686
rect 6943 2622 6949 2674
rect 7001 2622 7016 2674
rect 7068 2622 7083 2674
rect 7135 2622 7150 2674
rect 7202 2622 7217 2674
rect 7269 2622 7284 2674
rect 7336 2622 7342 2674
rect 6943 2610 7342 2622
rect 6943 2558 6949 2610
rect 7001 2558 7016 2610
rect 7068 2558 7083 2610
rect 7135 2558 7150 2610
rect 7202 2558 7217 2610
rect 7269 2558 7284 2610
rect 7336 2558 7342 2610
rect 12496 2686 12502 2738
rect 12554 2686 12569 2738
rect 12621 2686 12636 2738
rect 12688 2686 12703 2738
rect 12755 2686 12770 2738
rect 12822 2686 12837 2738
rect 12889 2686 12895 2738
rect 12496 2674 12895 2686
rect 12496 2622 12502 2674
rect 12554 2622 12569 2674
rect 12621 2622 12636 2674
rect 12688 2622 12703 2674
rect 12755 2622 12770 2674
rect 12822 2622 12837 2674
rect 12889 2622 12895 2674
rect 12496 2610 12895 2622
rect 12496 2558 12502 2610
rect 12554 2558 12569 2610
rect 12621 2558 12636 2610
rect 12688 2558 12703 2610
rect 12755 2558 12770 2610
rect 12822 2558 12837 2610
rect 12889 2558 12895 2610
rect 13427 2686 13433 2738
rect 13485 2686 13500 2738
rect 13552 2686 13567 2738
rect 13619 2686 13634 2738
rect 13686 2686 13701 2738
rect 13753 2686 13768 2738
rect 13820 2686 13826 2738
rect 13427 2674 13826 2686
rect 13427 2622 13433 2674
rect 13485 2622 13500 2674
rect 13552 2622 13567 2674
rect 13619 2622 13634 2674
rect 13686 2622 13701 2674
rect 13753 2622 13768 2674
rect 13820 2622 13826 2674
rect 13427 2610 13826 2622
rect 13427 2558 13433 2610
rect 13485 2558 13500 2610
rect 13552 2558 13567 2610
rect 13619 2558 13634 2610
rect 13686 2558 13701 2610
rect 13753 2558 13768 2610
rect 13820 2558 13826 2610
rect 19065 2686 19071 2738
rect 19123 2686 19154 2738
rect 19206 2686 19237 2738
rect 19289 2686 19321 2738
rect 19373 2686 19379 2738
tri 19818 2727 19829 2738 ne
rect 19829 2727 19971 2738
tri 19829 2715 19841 2727 ne
rect 19065 2674 19379 2686
rect 19065 2622 19071 2674
rect 19123 2622 19154 2674
rect 19206 2622 19237 2674
rect 19289 2622 19321 2674
rect 19373 2622 19379 2674
rect 19065 2610 19379 2622
rect 19065 2558 19071 2610
rect 19123 2558 19154 2610
rect 19206 2558 19237 2610
rect 19289 2558 19321 2610
rect 19373 2558 19379 2610
rect 19841 2693 19882 2727
rect 19916 2693 19971 2727
rect 19841 2654 19971 2693
rect 19841 2620 19882 2654
rect 19916 2620 19971 2654
rect 19841 2581 19971 2620
rect -52 2502 82 2541
rect -52 2468 -46 2502
rect -12 2468 42 2502
rect 76 2468 82 2502
rect -310 2406 -258 2409
rect -1722 2403 -258 2406
rect -1722 2400 -1042 2403
rect -1670 2369 -1042 2400
rect -1008 2397 -258 2403
rect -1008 2369 -310 2397
rect -1670 2356 -310 2369
rect -1722 2336 -1670 2348
rect -310 2339 -258 2345
rect -52 2429 82 2468
rect 19841 2547 19882 2581
rect 19916 2547 19971 2581
rect 19841 2508 19971 2547
rect 19841 2474 19882 2508
rect 19916 2474 19971 2508
rect -52 2395 -46 2429
rect -12 2395 42 2429
rect 76 2395 82 2429
rect -52 2356 82 2395
rect -1722 2278 -1670 2284
rect -52 2322 -46 2356
rect -12 2322 42 2356
rect 76 2322 82 2356
rect -52 2283 82 2322
rect -52 2249 -46 2283
rect -12 2249 42 2283
rect 76 2249 82 2283
rect -52 2210 82 2249
rect -52 2176 -46 2210
rect -12 2176 42 2210
rect 76 2176 82 2210
rect -52 2137 82 2176
rect -1596 2114 -799 2120
rect -1596 2080 -1584 2114
rect -1550 2080 -1503 2114
rect -1469 2080 -1423 2114
rect -1389 2080 -1343 2114
rect -1309 2080 -1263 2114
rect -1229 2080 -1183 2114
rect -1149 2080 -1103 2114
rect -1069 2080 -1023 2114
rect -989 2080 -943 2114
rect -909 2103 -799 2114
tri -799 2103 -782 2120 sw
rect -52 2103 -46 2137
rect -12 2103 42 2137
rect 76 2103 82 2137
rect -909 2080 -782 2103
rect -1596 2077 -782 2080
tri -782 2077 -756 2103 sw
rect -1596 2074 -414 2077
tri -835 2070 -831 2074 ne
rect -831 2071 -414 2074
rect -831 2070 -466 2071
tri -831 2064 -825 2070 ne
rect -825 2064 -466 2070
tri -825 2041 -802 2064 ne
rect -802 2041 -466 2064
rect -1647 2035 -1289 2041
tri -802 2039 -800 2041 ne
rect -800 2039 -466 2041
rect -1647 2029 -1636 2035
rect -1584 2029 -1289 2035
rect -1647 1995 -1641 2029
rect -1584 1995 -1329 2029
rect -1295 1995 -1289 2029
rect -1647 1983 -1636 1995
rect -1584 1983 -1289 1995
rect -1647 1965 -1289 1983
rect -1647 1956 -1636 1965
rect -1584 1956 -1289 1965
rect -1647 1922 -1641 1956
rect -1584 1922 -1329 1956
rect -1295 1922 -1289 1956
rect -466 2007 -414 2019
rect -466 1949 -414 1955
rect -52 2064 82 2103
rect -52 2030 -46 2064
rect -12 2030 42 2064
rect 76 2030 82 2064
rect 1021 2437 1920 2441
rect 1021 2385 1027 2437
rect 1079 2385 1092 2437
rect 1144 2385 1157 2437
rect 1209 2385 1222 2437
rect 1274 2385 1286 2437
rect 1338 2385 1350 2437
rect 1402 2385 1414 2437
rect 1466 2385 1478 2437
rect 1530 2385 1542 2437
rect 1594 2385 1606 2437
rect 1658 2385 1670 2437
rect 1722 2385 1734 2437
rect 1786 2385 1798 2437
rect 1850 2385 1862 2437
rect 1914 2385 1920 2437
rect 1021 2369 1920 2385
rect 1021 2317 1027 2369
rect 1079 2317 1092 2369
rect 1144 2317 1157 2369
rect 1209 2317 1222 2369
rect 1274 2317 1286 2369
rect 1338 2317 1350 2369
rect 1402 2317 1414 2369
rect 1466 2317 1478 2369
rect 1530 2317 1542 2369
rect 1594 2317 1606 2369
rect 1658 2317 1670 2369
rect 1722 2317 1734 2369
rect 1786 2317 1798 2369
rect 1850 2317 1862 2369
rect 1914 2317 1920 2369
rect 1021 2301 1920 2317
rect 1021 2249 1027 2301
rect 1079 2249 1092 2301
rect 1144 2249 1157 2301
rect 1209 2249 1222 2301
rect 1274 2249 1286 2301
rect 1338 2249 1350 2301
rect 1402 2249 1414 2301
rect 1466 2249 1478 2301
rect 1530 2249 1542 2301
rect 1594 2249 1606 2301
rect 1658 2249 1670 2301
rect 1722 2249 1734 2301
rect 1786 2249 1798 2301
rect 1850 2249 1862 2301
rect 1914 2249 1920 2301
rect 1021 2233 1920 2249
rect 1021 2181 1027 2233
rect 1079 2181 1092 2233
rect 1144 2181 1157 2233
rect 1209 2181 1222 2233
rect 1274 2181 1286 2233
rect 1338 2181 1350 2233
rect 1402 2181 1414 2233
rect 1466 2181 1478 2233
rect 1530 2181 1542 2233
rect 1594 2181 1606 2233
rect 1658 2181 1670 2233
rect 1722 2181 1734 2233
rect 1786 2181 1798 2233
rect 1850 2181 1862 2233
rect 1914 2181 1920 2233
rect 1021 2165 1920 2181
rect 1021 2113 1027 2165
rect 1079 2113 1092 2165
rect 1144 2113 1157 2165
rect 1209 2113 1222 2165
rect 1274 2113 1286 2165
rect 1338 2113 1350 2165
rect 1402 2113 1414 2165
rect 1466 2113 1478 2165
rect 1530 2113 1542 2165
rect 1594 2113 1606 2165
rect 1658 2113 1670 2165
rect 1722 2113 1734 2165
rect 1786 2113 1798 2165
rect 1850 2113 1862 2165
rect 1914 2113 1920 2165
rect 1021 2097 1920 2113
rect 1021 2045 1027 2097
rect 1079 2045 1092 2097
rect 1144 2045 1157 2097
rect 1209 2045 1222 2097
rect 1274 2045 1286 2097
rect 1338 2045 1350 2097
rect 1402 2045 1414 2097
rect 1466 2045 1478 2097
rect 1530 2045 1542 2097
rect 1594 2045 1606 2097
rect 1658 2045 1670 2097
rect 1722 2045 1734 2097
rect 1786 2045 1798 2097
rect 1850 2045 1862 2097
rect 1914 2045 1920 2097
rect 1021 2041 1920 2045
rect 7505 2437 8404 2441
rect 7505 2385 7511 2437
rect 7563 2385 7576 2437
rect 7628 2385 7641 2437
rect 7693 2385 7706 2437
rect 7758 2385 7770 2437
rect 7822 2385 7834 2437
rect 7886 2385 7898 2437
rect 7950 2385 7962 2437
rect 8014 2385 8026 2437
rect 8078 2385 8090 2437
rect 8142 2385 8154 2437
rect 8206 2385 8218 2437
rect 8270 2385 8282 2437
rect 8334 2385 8346 2437
rect 8398 2385 8404 2437
rect 7505 2369 8404 2385
rect 7505 2317 7511 2369
rect 7563 2317 7576 2369
rect 7628 2317 7641 2369
rect 7693 2317 7706 2369
rect 7758 2317 7770 2369
rect 7822 2317 7834 2369
rect 7886 2317 7898 2369
rect 7950 2317 7962 2369
rect 8014 2317 8026 2369
rect 8078 2317 8090 2369
rect 8142 2317 8154 2369
rect 8206 2317 8218 2369
rect 8270 2317 8282 2369
rect 8334 2317 8346 2369
rect 8398 2317 8404 2369
rect 7505 2301 8404 2317
rect 7505 2249 7511 2301
rect 7563 2249 7576 2301
rect 7628 2249 7641 2301
rect 7693 2249 7706 2301
rect 7758 2249 7770 2301
rect 7822 2249 7834 2301
rect 7886 2249 7898 2301
rect 7950 2249 7962 2301
rect 8014 2249 8026 2301
rect 8078 2249 8090 2301
rect 8142 2249 8154 2301
rect 8206 2249 8218 2301
rect 8270 2249 8282 2301
rect 8334 2249 8346 2301
rect 8398 2249 8404 2301
rect 7505 2233 8404 2249
rect 7505 2181 7511 2233
rect 7563 2181 7576 2233
rect 7628 2181 7641 2233
rect 7693 2181 7706 2233
rect 7758 2181 7770 2233
rect 7822 2181 7834 2233
rect 7886 2181 7898 2233
rect 7950 2181 7962 2233
rect 8014 2181 8026 2233
rect 8078 2181 8090 2233
rect 8142 2181 8154 2233
rect 8206 2181 8218 2233
rect 8270 2181 8282 2233
rect 8334 2181 8346 2233
rect 8398 2181 8404 2233
rect 7505 2165 8404 2181
rect 7505 2113 7511 2165
rect 7563 2113 7576 2165
rect 7628 2113 7641 2165
rect 7693 2113 7706 2165
rect 7758 2113 7770 2165
rect 7822 2113 7834 2165
rect 7886 2113 7898 2165
rect 7950 2113 7962 2165
rect 8014 2113 8026 2165
rect 8078 2113 8090 2165
rect 8142 2113 8154 2165
rect 8206 2113 8218 2165
rect 8270 2113 8282 2165
rect 8334 2113 8346 2165
rect 8398 2113 8404 2165
rect 7505 2097 8404 2113
rect 7505 2045 7511 2097
rect 7563 2045 7576 2097
rect 7628 2045 7641 2097
rect 7693 2045 7706 2097
rect 7758 2045 7770 2097
rect 7822 2045 7834 2097
rect 7886 2045 7898 2097
rect 7950 2045 7962 2097
rect 8014 2045 8026 2097
rect 8078 2045 8090 2097
rect 8142 2045 8154 2097
rect 8206 2045 8218 2097
rect 8270 2045 8282 2097
rect 8334 2045 8346 2097
rect 8398 2045 8404 2097
rect 7505 2041 8404 2045
rect 11434 2437 12333 2441
rect 11434 2385 11440 2437
rect 11492 2385 11504 2437
rect 11556 2385 11568 2437
rect 11620 2385 11632 2437
rect 11684 2385 11696 2437
rect 11748 2385 11760 2437
rect 11812 2385 11824 2437
rect 11876 2385 11888 2437
rect 11940 2385 11952 2437
rect 12004 2385 12016 2437
rect 12068 2385 12080 2437
rect 12132 2385 12145 2437
rect 12197 2385 12210 2437
rect 12262 2385 12275 2437
rect 12327 2385 12333 2437
rect 11434 2369 12333 2385
rect 11434 2317 11440 2369
rect 11492 2317 11504 2369
rect 11556 2317 11568 2369
rect 11620 2317 11632 2369
rect 11684 2317 11696 2369
rect 11748 2317 11760 2369
rect 11812 2317 11824 2369
rect 11876 2317 11888 2369
rect 11940 2317 11952 2369
rect 12004 2317 12016 2369
rect 12068 2317 12080 2369
rect 12132 2317 12145 2369
rect 12197 2317 12210 2369
rect 12262 2317 12275 2369
rect 12327 2317 12333 2369
rect 11434 2301 12333 2317
rect 11434 2249 11440 2301
rect 11492 2249 11504 2301
rect 11556 2249 11568 2301
rect 11620 2249 11632 2301
rect 11684 2249 11696 2301
rect 11748 2249 11760 2301
rect 11812 2249 11824 2301
rect 11876 2249 11888 2301
rect 11940 2249 11952 2301
rect 12004 2249 12016 2301
rect 12068 2249 12080 2301
rect 12132 2249 12145 2301
rect 12197 2249 12210 2301
rect 12262 2249 12275 2301
rect 12327 2249 12333 2301
rect 11434 2233 12333 2249
rect 11434 2181 11440 2233
rect 11492 2181 11504 2233
rect 11556 2181 11568 2233
rect 11620 2181 11632 2233
rect 11684 2181 11696 2233
rect 11748 2181 11760 2233
rect 11812 2181 11824 2233
rect 11876 2181 11888 2233
rect 11940 2181 11952 2233
rect 12004 2181 12016 2233
rect 12068 2181 12080 2233
rect 12132 2181 12145 2233
rect 12197 2181 12210 2233
rect 12262 2181 12275 2233
rect 12327 2181 12333 2233
rect 11434 2165 12333 2181
rect 11434 2113 11440 2165
rect 11492 2113 11504 2165
rect 11556 2113 11568 2165
rect 11620 2113 11632 2165
rect 11684 2113 11696 2165
rect 11748 2113 11760 2165
rect 11812 2113 11824 2165
rect 11876 2113 11888 2165
rect 11940 2113 11952 2165
rect 12004 2113 12016 2165
rect 12068 2113 12080 2165
rect 12132 2113 12145 2165
rect 12197 2113 12210 2165
rect 12262 2113 12275 2165
rect 12327 2113 12333 2165
rect 11434 2097 12333 2113
rect 11434 2045 11440 2097
rect 11492 2045 11504 2097
rect 11556 2045 11568 2097
rect 11620 2045 11632 2097
rect 11684 2045 11696 2097
rect 11748 2045 11760 2097
rect 11812 2045 11824 2097
rect 11876 2045 11888 2097
rect 11940 2045 11952 2097
rect 12004 2045 12016 2097
rect 12068 2045 12080 2097
rect 12132 2045 12145 2097
rect 12197 2045 12210 2097
rect 12262 2045 12275 2097
rect 12327 2045 12333 2097
rect 11434 2041 12333 2045
rect 13989 2437 14888 2441
rect 13989 2385 13995 2437
rect 14047 2385 14060 2437
rect 14112 2385 14125 2437
rect 14177 2385 14190 2437
rect 14242 2385 14254 2437
rect 14306 2385 14318 2437
rect 14370 2385 14382 2437
rect 14434 2385 14446 2437
rect 14498 2385 14510 2437
rect 14562 2385 14574 2437
rect 14626 2385 14638 2437
rect 14690 2385 14702 2437
rect 14754 2385 14766 2437
rect 14818 2385 14830 2437
rect 14882 2385 14888 2437
rect 13989 2369 14888 2385
rect 13989 2317 13995 2369
rect 14047 2317 14060 2369
rect 14112 2317 14125 2369
rect 14177 2317 14190 2369
rect 14242 2317 14254 2369
rect 14306 2317 14318 2369
rect 14370 2317 14382 2369
rect 14434 2317 14446 2369
rect 14498 2317 14510 2369
rect 14562 2317 14574 2369
rect 14626 2317 14638 2369
rect 14690 2317 14702 2369
rect 14754 2317 14766 2369
rect 14818 2317 14830 2369
rect 14882 2317 14888 2369
rect 13989 2301 14888 2317
rect 13989 2249 13995 2301
rect 14047 2249 14060 2301
rect 14112 2249 14125 2301
rect 14177 2249 14190 2301
rect 14242 2249 14254 2301
rect 14306 2249 14318 2301
rect 14370 2249 14382 2301
rect 14434 2249 14446 2301
rect 14498 2249 14510 2301
rect 14562 2249 14574 2301
rect 14626 2249 14638 2301
rect 14690 2249 14702 2301
rect 14754 2249 14766 2301
rect 14818 2249 14830 2301
rect 14882 2249 14888 2301
rect 13989 2233 14888 2249
rect 13989 2181 13995 2233
rect 14047 2181 14060 2233
rect 14112 2181 14125 2233
rect 14177 2181 14190 2233
rect 14242 2181 14254 2233
rect 14306 2181 14318 2233
rect 14370 2181 14382 2233
rect 14434 2181 14446 2233
rect 14498 2181 14510 2233
rect 14562 2181 14574 2233
rect 14626 2181 14638 2233
rect 14690 2181 14702 2233
rect 14754 2181 14766 2233
rect 14818 2181 14830 2233
rect 14882 2181 14888 2233
rect 13989 2165 14888 2181
rect 13989 2113 13995 2165
rect 14047 2113 14060 2165
rect 14112 2113 14125 2165
rect 14177 2113 14190 2165
rect 14242 2113 14254 2165
rect 14306 2113 14318 2165
rect 14370 2113 14382 2165
rect 14434 2113 14446 2165
rect 14498 2113 14510 2165
rect 14562 2113 14574 2165
rect 14626 2113 14638 2165
rect 14690 2113 14702 2165
rect 14754 2113 14766 2165
rect 14818 2113 14830 2165
rect 14882 2113 14888 2165
rect 13989 2097 14888 2113
rect 13989 2045 13995 2097
rect 14047 2045 14060 2097
rect 14112 2045 14125 2097
rect 14177 2045 14190 2097
rect 14242 2045 14254 2097
rect 14306 2045 14318 2097
rect 14370 2045 14382 2097
rect 14434 2045 14446 2097
rect 14498 2045 14510 2097
rect 14562 2045 14574 2097
rect 14626 2045 14638 2097
rect 14690 2045 14702 2097
rect 14754 2045 14766 2097
rect 14818 2045 14830 2097
rect 14882 2045 14888 2097
rect 13989 2041 14888 2045
rect 17918 2437 18817 2441
rect 17918 2385 17924 2437
rect 17976 2385 17988 2437
rect 18040 2385 18052 2437
rect 18104 2385 18116 2437
rect 18168 2385 18180 2437
rect 18232 2385 18244 2437
rect 18296 2385 18308 2437
rect 18360 2385 18372 2437
rect 18424 2385 18436 2437
rect 18488 2385 18500 2437
rect 18552 2385 18564 2437
rect 18616 2385 18629 2437
rect 18681 2385 18694 2437
rect 18746 2385 18759 2437
rect 18811 2385 18817 2437
rect 17918 2369 18817 2385
rect 17918 2317 17924 2369
rect 17976 2317 17988 2369
rect 18040 2317 18052 2369
rect 18104 2317 18116 2369
rect 18168 2317 18180 2369
rect 18232 2317 18244 2369
rect 18296 2317 18308 2369
rect 18360 2317 18372 2369
rect 18424 2317 18436 2369
rect 18488 2317 18500 2369
rect 18552 2317 18564 2369
rect 18616 2317 18629 2369
rect 18681 2317 18694 2369
rect 18746 2317 18759 2369
rect 18811 2317 18817 2369
rect 17918 2301 18817 2317
rect 17918 2249 17924 2301
rect 17976 2249 17988 2301
rect 18040 2249 18052 2301
rect 18104 2249 18116 2301
rect 18168 2249 18180 2301
rect 18232 2249 18244 2301
rect 18296 2249 18308 2301
rect 18360 2249 18372 2301
rect 18424 2249 18436 2301
rect 18488 2249 18500 2301
rect 18552 2249 18564 2301
rect 18616 2249 18629 2301
rect 18681 2249 18694 2301
rect 18746 2249 18759 2301
rect 18811 2249 18817 2301
rect 17918 2233 18817 2249
rect 17918 2181 17924 2233
rect 17976 2181 17988 2233
rect 18040 2181 18052 2233
rect 18104 2181 18116 2233
rect 18168 2181 18180 2233
rect 18232 2181 18244 2233
rect 18296 2181 18308 2233
rect 18360 2181 18372 2233
rect 18424 2181 18436 2233
rect 18488 2181 18500 2233
rect 18552 2181 18564 2233
rect 18616 2181 18629 2233
rect 18681 2181 18694 2233
rect 18746 2181 18759 2233
rect 18811 2181 18817 2233
rect 17918 2165 18817 2181
rect 17918 2113 17924 2165
rect 17976 2113 17988 2165
rect 18040 2113 18052 2165
rect 18104 2113 18116 2165
rect 18168 2113 18180 2165
rect 18232 2113 18244 2165
rect 18296 2113 18308 2165
rect 18360 2113 18372 2165
rect 18424 2113 18436 2165
rect 18488 2113 18500 2165
rect 18552 2113 18564 2165
rect 18616 2113 18629 2165
rect 18681 2113 18694 2165
rect 18746 2113 18759 2165
rect 18811 2113 18817 2165
rect 17918 2097 18817 2113
rect 17918 2045 17924 2097
rect 17976 2045 17988 2097
rect 18040 2045 18052 2097
rect 18104 2045 18116 2097
rect 18168 2045 18180 2097
rect 18232 2045 18244 2097
rect 18296 2045 18308 2097
rect 18360 2045 18372 2097
rect 18424 2045 18436 2097
rect 18488 2045 18500 2097
rect 18552 2045 18564 2097
rect 18616 2045 18629 2097
rect 18681 2045 18694 2097
rect 18746 2045 18759 2097
rect 18811 2045 18817 2097
rect 17918 2041 18817 2045
rect 19841 2435 19971 2474
rect 19841 2401 19882 2435
rect 19916 2401 19971 2435
rect 19841 2362 19971 2401
rect 19841 2328 19882 2362
rect 19916 2328 19971 2362
rect 19841 2289 19971 2328
rect 19841 2255 19882 2289
rect 19916 2255 19971 2289
rect 19841 2216 19971 2255
rect 19841 2182 19882 2216
rect 19916 2182 19971 2216
rect 19841 2143 19971 2182
rect 19841 2109 19882 2143
rect 19916 2109 19971 2143
rect 19841 2070 19971 2109
rect -52 1991 82 2030
rect -52 1957 -46 1991
rect -12 1957 42 1991
rect 76 1957 82 1991
rect -1647 1913 -1636 1922
rect -1584 1913 -1289 1922
rect -1647 1894 -1289 1913
rect -1647 1882 -1636 1894
rect -1584 1882 -1289 1894
rect -1736 1849 -1684 1855
rect -1647 1848 -1641 1882
rect -1584 1848 -1329 1882
rect -1295 1848 -1289 1882
rect -1647 1842 -1636 1848
rect -1584 1842 -1289 1848
rect -1647 1836 -1289 1842
rect -52 1918 82 1957
rect 19841 2036 19882 2070
rect 19916 2036 19971 2070
rect 19841 1997 19971 2036
rect 19841 1963 19882 1997
rect 19916 1963 19971 1997
tri 306 1924 311 1929 se
rect 311 1924 3317 1929
tri 3317 1924 3322 1929 sw
tri 3548 1924 3553 1929 se
rect 3553 1924 6559 1929
tri 6559 1924 6564 1929 sw
tri 6790 1924 6795 1929 se
rect 6795 1924 9801 1929
tri 9801 1924 9806 1929 sw
rect 19841 1924 19971 1963
rect -52 1884 -46 1918
rect -12 1884 42 1918
rect 76 1884 82 1918
tri 272 1890 306 1924 se
rect 306 1919 3322 1924
rect 306 1890 644 1919
rect -52 1845 82 1884
rect -1736 1785 -1684 1797
rect -630 1807 -578 1813
rect -1684 1765 -630 1777
rect -1684 1733 -1485 1765
rect -1736 1731 -1485 1733
rect -1451 1755 -630 1765
rect -1451 1743 -578 1755
rect -1451 1731 -630 1743
rect -1736 1727 -630 1731
rect -1491 1693 -1445 1727
rect -1491 1659 -1485 1693
rect -1451 1659 -1445 1693
rect -630 1685 -578 1691
rect -52 1811 -46 1845
rect -12 1811 42 1845
rect 76 1811 82 1845
rect -52 1772 82 1811
rect -52 1738 -46 1772
rect -12 1738 42 1772
rect 76 1738 82 1772
tri 264 1882 272 1890 se
rect 272 1882 644 1890
rect 264 1867 644 1882
rect 696 1867 728 1919
rect 780 1867 812 1919
rect 864 1867 895 1919
rect 947 1890 3322 1919
tri 3322 1890 3356 1924 sw
tri 3514 1890 3548 1924 se
rect 3548 1919 6564 1924
rect 3548 1890 6018 1919
rect 947 1882 3356 1890
tri 3356 1882 3364 1890 sw
tri 3506 1882 3514 1890 se
rect 3514 1882 6018 1890
rect 947 1867 6018 1882
rect 6070 1867 6085 1919
rect 6137 1867 6152 1919
rect 6204 1867 6219 1919
rect 6271 1867 6286 1919
rect 6338 1867 6353 1919
rect 6405 1890 6564 1919
tri 6564 1890 6598 1924 sw
tri 6756 1890 6790 1924 se
rect 6790 1919 9806 1924
rect 6790 1890 6949 1919
rect 6405 1882 6598 1890
tri 6598 1882 6606 1890 sw
tri 6748 1882 6756 1890 se
rect 6756 1882 6949 1890
rect 6405 1867 6949 1882
rect 7001 1867 7016 1919
rect 7068 1867 7083 1919
rect 7135 1867 7150 1919
rect 7202 1867 7217 1919
rect 7269 1867 7284 1919
rect 7336 1890 9806 1919
tri 9806 1890 9840 1924 sw
rect 7336 1882 9840 1890
tri 9840 1882 9848 1890 sw
rect 12496 1882 12502 1919
rect 7336 1867 12502 1882
rect 12554 1867 12569 1919
rect 12621 1867 12636 1919
rect 12688 1867 12703 1919
rect 12755 1867 12770 1919
rect 12822 1867 12837 1919
rect 12889 1882 12895 1919
rect 12889 1867 13043 1882
rect 264 1855 13043 1867
rect 264 1803 644 1855
rect 696 1803 728 1855
rect 780 1803 812 1855
rect 864 1803 895 1855
rect 947 1803 6018 1855
rect 6070 1803 6085 1855
rect 6137 1803 6152 1855
rect 6204 1803 6219 1855
rect 6271 1803 6286 1855
rect 6338 1803 6353 1855
rect 6405 1803 6949 1855
rect 7001 1803 7016 1855
rect 7068 1803 7083 1855
rect 7135 1803 7150 1855
rect 7202 1803 7217 1855
rect 7269 1803 7284 1855
rect 7336 1803 12502 1855
rect 12554 1803 12569 1855
rect 12621 1803 12636 1855
rect 12688 1803 12703 1855
rect 12755 1803 12770 1855
rect 12822 1803 12837 1855
rect 12889 1803 13043 1855
rect 264 1791 13043 1803
rect 264 1776 644 1791
tri 264 1744 296 1776 ne
rect 296 1744 644 1776
rect -52 1699 82 1738
tri 296 1729 311 1744 ne
rect 311 1739 644 1744
rect 696 1739 728 1791
rect 780 1739 812 1791
rect 864 1739 895 1791
rect 947 1776 6018 1791
rect 947 1744 3332 1776
tri 3332 1744 3364 1776 nw
tri 3506 1744 3538 1776 ne
rect 3538 1744 6018 1776
rect 947 1739 3317 1744
rect 311 1729 3317 1739
tri 3317 1729 3332 1744 nw
tri 3538 1729 3553 1744 ne
rect 3553 1739 6018 1744
rect 6070 1739 6085 1791
rect 6137 1739 6152 1791
rect 6204 1739 6219 1791
rect 6271 1739 6286 1791
rect 6338 1739 6353 1791
rect 6405 1776 6949 1791
rect 6405 1744 6574 1776
tri 6574 1744 6606 1776 nw
tri 6748 1744 6780 1776 ne
rect 6780 1744 6949 1776
rect 6405 1739 6559 1744
rect 3553 1729 6559 1739
tri 6559 1729 6574 1744 nw
tri 6780 1729 6795 1744 ne
rect 6795 1739 6949 1744
rect 7001 1739 7016 1791
rect 7068 1739 7083 1791
rect 7135 1739 7150 1791
rect 7202 1739 7217 1791
rect 7269 1739 7284 1791
rect 7336 1776 12502 1791
rect 7336 1744 9816 1776
tri 9816 1744 9848 1776 nw
rect 7336 1739 9801 1744
rect 6795 1729 9801 1739
tri 9801 1729 9816 1744 nw
rect 12496 1739 12502 1776
rect 12554 1739 12569 1791
rect 12621 1739 12636 1791
rect 12688 1739 12703 1791
rect 12755 1739 12770 1791
rect 12822 1739 12837 1791
rect 12889 1776 13043 1791
rect 13427 1867 13433 1919
rect 13485 1867 13500 1919
rect 13552 1867 13567 1919
rect 13619 1867 13634 1919
rect 13686 1867 13701 1919
rect 13753 1867 13768 1919
rect 13820 1867 13826 1919
rect 13427 1855 13826 1867
rect 13427 1803 13433 1855
rect 13485 1803 13500 1855
rect 13552 1803 13567 1855
rect 13619 1803 13634 1855
rect 13686 1803 13701 1855
rect 13753 1803 13768 1855
rect 13820 1803 13826 1855
rect 13427 1791 13826 1803
rect 12889 1739 12895 1776
rect 13427 1739 13433 1791
rect 13485 1739 13500 1791
rect 13552 1739 13567 1791
rect 13619 1739 13634 1791
rect 13686 1739 13701 1791
rect 13753 1739 13768 1791
rect 13820 1739 13826 1791
rect 19065 1867 19071 1919
rect 19123 1867 19154 1919
rect 19206 1867 19237 1919
rect 19289 1867 19321 1919
rect 19373 1867 19379 1919
rect 19065 1855 19379 1867
rect 19065 1803 19071 1855
rect 19123 1803 19154 1855
rect 19206 1803 19237 1855
rect 19289 1803 19321 1855
rect 19373 1803 19379 1855
rect 19065 1791 19379 1803
rect 19065 1739 19071 1791
rect 19123 1739 19154 1791
rect 19206 1739 19237 1791
rect 19289 1739 19321 1791
rect 19373 1739 19379 1791
rect 19841 1890 19882 1924
rect 19916 1890 19971 1924
rect 19841 1851 19971 1890
rect 19841 1817 19882 1851
rect 19916 1817 19971 1851
rect 19841 1778 19971 1817
rect 19841 1744 19882 1778
rect 19916 1744 19971 1778
rect -1491 1647 -1445 1659
rect -52 1665 -46 1699
rect -12 1665 42 1699
rect 76 1665 82 1699
rect 19841 1705 19971 1744
tri 310 1686 311 1687 se
rect 311 1686 3317 1687
tri 3317 1686 3318 1687 sw
tri 3552 1686 3553 1687 se
rect 3553 1686 6559 1687
tri 6559 1686 6560 1687 sw
tri 6794 1686 6795 1687 se
rect 6795 1686 9801 1687
tri 9801 1686 9802 1687 sw
tri 10036 1686 10037 1687 se
rect 10037 1686 13043 1687
tri 13043 1686 13044 1687 sw
tri 13278 1686 13279 1687 se
rect 13279 1686 16285 1687
tri 16285 1686 16286 1687 sw
tri 16520 1686 16521 1687 se
rect 16521 1686 19527 1687
tri 19527 1686 19528 1687 sw
tri 295 1671 310 1686 se
rect 310 1685 9802 1686
rect 310 1671 2677 1685
rect -52 1626 82 1665
tri 271 1647 295 1671 se
rect 295 1647 2677 1671
rect -52 1592 -46 1626
rect -12 1592 42 1626
rect 76 1592 82 1626
rect -52 1553 82 1592
tri -151 1519 -132 1538 se
rect -132 1532 -80 1538
tri -161 1509 -151 1519 se
rect -151 1509 -132 1519
rect -630 1503 -132 1509
rect -578 1480 -132 1503
rect -578 1468 -80 1480
rect -578 1451 -132 1468
rect -630 1440 -132 1451
rect -630 1439 -515 1440
rect -578 1412 -515 1439
tri -515 1412 -487 1440 nw
rect -578 1410 -517 1412
tri -517 1410 -515 1412 nw
rect -132 1410 -80 1416
rect -52 1519 -46 1553
rect -12 1519 42 1553
rect 76 1519 82 1553
tri 264 1640 271 1647 se
rect 271 1640 2677 1647
rect 2729 1640 2744 1685
rect 2796 1640 2811 1685
rect 2863 1640 2878 1685
rect 2930 1640 2945 1685
rect 2997 1640 3012 1685
rect 264 1606 364 1640
rect 398 1606 437 1640
rect 471 1606 510 1640
rect 544 1606 583 1640
rect 617 1606 656 1640
rect 690 1606 729 1640
rect 763 1606 802 1640
rect 836 1606 875 1640
rect 909 1606 948 1640
rect 982 1606 1021 1640
rect 1055 1606 1094 1640
rect 1128 1606 1167 1640
rect 1201 1606 1240 1640
rect 1274 1606 1313 1640
rect 1347 1606 1386 1640
rect 1420 1606 1459 1640
rect 1493 1606 1532 1640
rect 1566 1606 1605 1640
rect 1639 1606 1678 1640
rect 1712 1606 1751 1640
rect 1785 1606 1824 1640
rect 1858 1606 1898 1640
rect 1932 1606 1972 1640
rect 2006 1606 2046 1640
rect 2080 1606 2120 1640
rect 2154 1606 2194 1640
rect 2228 1606 2268 1640
rect 2302 1606 2342 1640
rect 2376 1606 2416 1640
rect 2450 1606 2490 1640
rect 2524 1606 2564 1640
rect 2598 1606 2638 1640
rect 2672 1633 2677 1640
rect 2930 1633 2934 1640
rect 2997 1633 3008 1640
rect 3064 1633 3079 1685
rect 3131 1633 3146 1685
rect 3198 1633 3213 1685
rect 3265 1633 3279 1685
rect 3331 1633 3345 1685
rect 3397 1633 3411 1685
rect 3463 1633 3477 1685
rect 3529 1633 3543 1685
rect 3595 1640 4882 1685
rect 4934 1640 4971 1685
rect 5023 1640 5059 1685
rect 5111 1640 5720 1685
rect 5772 1640 5799 1685
rect 3595 1633 3606 1640
rect 2672 1613 2712 1633
rect 2746 1613 2786 1633
rect 2820 1613 2860 1633
rect 2894 1613 2934 1633
rect 2968 1613 3008 1633
rect 3042 1613 3082 1633
rect 3116 1613 3156 1633
rect 3190 1613 3230 1633
rect 3264 1613 3606 1633
rect 2672 1606 2677 1613
rect 2930 1606 2934 1613
rect 2997 1606 3008 1613
rect 264 1568 2677 1606
rect 2729 1568 2744 1606
rect 2796 1568 2811 1606
rect 2863 1568 2878 1606
rect 2930 1568 2945 1606
rect 2997 1568 3012 1606
rect 264 1534 364 1568
rect 398 1534 437 1568
rect 471 1534 510 1568
rect 544 1534 583 1568
rect 617 1534 656 1568
rect 690 1534 729 1568
rect 763 1534 802 1568
rect 836 1534 875 1568
rect 909 1534 948 1568
rect 982 1534 1021 1568
rect 1055 1534 1094 1568
rect 1128 1534 1167 1568
rect 1201 1534 1240 1568
rect 1274 1534 1313 1568
rect 1347 1534 1386 1568
rect 1420 1534 1459 1568
rect 1493 1534 1532 1568
rect 1566 1534 1605 1568
rect 1639 1534 1678 1568
rect 1712 1534 1751 1568
rect 1785 1534 1824 1568
rect 1858 1534 1898 1568
rect 1932 1534 1972 1568
rect 2006 1534 2046 1568
rect 2080 1534 2120 1568
rect 2154 1534 2194 1568
rect 2228 1534 2268 1568
rect 2302 1534 2342 1568
rect 2376 1534 2416 1568
rect 2450 1534 2490 1568
rect 2524 1534 2564 1568
rect 2598 1534 2638 1568
rect 2672 1561 2677 1568
rect 2930 1561 2934 1568
rect 2997 1561 3008 1568
rect 3064 1561 3079 1613
rect 3131 1561 3146 1613
rect 3198 1561 3213 1613
rect 3265 1561 3279 1613
rect 3331 1561 3345 1613
rect 3397 1561 3411 1613
rect 3463 1561 3477 1613
rect 3529 1561 3543 1613
rect 3595 1606 3606 1613
rect 3640 1606 3680 1640
rect 3714 1606 3754 1640
rect 3788 1606 3828 1640
rect 3862 1606 3902 1640
rect 3936 1606 3976 1640
rect 4010 1606 4050 1640
rect 4084 1606 4124 1640
rect 4158 1606 4198 1640
rect 4232 1606 4272 1640
rect 4306 1606 4346 1640
rect 4380 1606 4420 1640
rect 4454 1606 4494 1640
rect 4528 1606 4568 1640
rect 4602 1606 4642 1640
rect 4676 1606 4716 1640
rect 4750 1606 4790 1640
rect 4824 1606 4864 1640
rect 4934 1633 4938 1640
rect 5046 1633 5059 1640
rect 4898 1613 4938 1633
rect 4972 1613 5012 1633
rect 5046 1613 5085 1633
rect 4934 1606 4938 1613
rect 5046 1606 5059 1613
rect 5119 1606 5158 1640
rect 5192 1606 5231 1640
rect 5265 1606 5304 1640
rect 5338 1606 5377 1640
rect 5411 1606 5450 1640
rect 5484 1606 5523 1640
rect 5557 1606 5596 1640
rect 5630 1606 5669 1640
rect 5703 1633 5720 1640
rect 5776 1633 5799 1640
rect 5851 1633 5878 1685
rect 5930 1640 6497 1685
rect 5930 1633 5961 1640
rect 5703 1613 5742 1633
rect 5776 1613 5815 1633
rect 5849 1613 5888 1633
rect 5922 1613 5961 1633
rect 5703 1606 5720 1613
rect 5776 1606 5799 1613
rect 3595 1568 4882 1606
rect 4934 1568 4971 1606
rect 5023 1568 5059 1606
rect 5111 1568 5720 1606
rect 5772 1568 5799 1606
rect 3595 1561 3606 1568
rect 2672 1541 2712 1561
rect 2746 1541 2786 1561
rect 2820 1541 2860 1561
rect 2894 1541 2934 1561
rect 2968 1541 3008 1561
rect 3042 1541 3082 1561
rect 3116 1541 3156 1561
rect 3190 1541 3230 1561
rect 3264 1541 3606 1561
rect 2672 1534 2677 1541
rect 2930 1534 2934 1541
rect 2997 1534 3008 1541
tri 264 1525 273 1534 ne
rect 273 1525 2677 1534
rect -52 1479 82 1519
tri 273 1488 310 1525 ne
rect 310 1489 2677 1525
rect 2729 1489 2744 1534
rect 2796 1489 2811 1534
rect 2863 1489 2878 1534
rect 2930 1489 2945 1534
rect 2997 1489 3012 1534
rect 3064 1489 3079 1541
rect 3131 1489 3146 1541
rect 3198 1489 3213 1541
rect 3265 1489 3279 1541
rect 3331 1489 3345 1541
rect 3397 1489 3411 1541
rect 3463 1489 3477 1541
rect 3529 1489 3543 1541
rect 3595 1534 3606 1541
rect 3640 1534 3680 1568
rect 3714 1534 3754 1568
rect 3788 1534 3828 1568
rect 3862 1534 3902 1568
rect 3936 1534 3976 1568
rect 4010 1534 4050 1568
rect 4084 1534 4124 1568
rect 4158 1534 4198 1568
rect 4232 1534 4272 1568
rect 4306 1534 4346 1568
rect 4380 1534 4420 1568
rect 4454 1534 4494 1568
rect 4528 1534 4568 1568
rect 4602 1534 4642 1568
rect 4676 1534 4716 1568
rect 4750 1534 4790 1568
rect 4824 1534 4864 1568
rect 4934 1561 4938 1568
rect 5046 1561 5059 1568
rect 4898 1541 4938 1561
rect 4972 1541 5012 1561
rect 5046 1541 5085 1561
rect 4934 1534 4938 1541
rect 5046 1534 5059 1541
rect 5119 1534 5158 1568
rect 5192 1534 5231 1568
rect 5265 1534 5304 1568
rect 5338 1534 5377 1568
rect 5411 1534 5450 1568
rect 5484 1534 5523 1568
rect 5557 1534 5596 1568
rect 5630 1534 5669 1568
rect 5703 1561 5720 1568
rect 5776 1561 5799 1568
rect 5851 1561 5878 1613
rect 5930 1606 5961 1613
rect 5995 1606 6034 1640
rect 6068 1606 6107 1640
rect 6141 1606 6180 1640
rect 6214 1606 6253 1640
rect 6287 1606 6326 1640
rect 6360 1606 6399 1640
rect 6433 1606 6472 1640
rect 6549 1633 6574 1685
rect 6626 1633 6651 1685
rect 6703 1633 6728 1685
rect 6780 1633 6805 1685
rect 6857 1640 9525 1685
rect 9577 1640 9592 1685
rect 9644 1640 9659 1685
rect 9711 1640 9726 1685
rect 9778 1671 9802 1685
tri 9802 1671 9817 1686 sw
tri 10021 1671 10036 1686 se
rect 10036 1671 13044 1686
tri 13044 1671 13059 1686 sw
tri 13263 1671 13278 1686 se
rect 13278 1671 16286 1686
tri 16286 1671 16301 1686 sw
rect 16397 1685 19528 1686
rect 9778 1640 9817 1671
tri 9817 1640 9848 1671 sw
tri 9990 1640 10021 1671 se
rect 10021 1640 13059 1671
tri 13059 1640 13090 1671 sw
tri 13232 1640 13263 1671 se
rect 13263 1640 16301 1671
tri 16301 1640 16332 1671 sw
rect 16397 1640 16403 1685
rect 6506 1613 6848 1633
rect 5930 1568 6497 1606
rect 5930 1561 5961 1568
rect 5703 1541 5742 1561
rect 5776 1541 5815 1561
rect 5849 1541 5888 1561
rect 5922 1541 5961 1561
rect 5703 1534 5720 1541
rect 5776 1534 5799 1541
rect 3595 1489 4882 1534
rect 4934 1489 4971 1534
rect 5023 1489 5059 1534
rect 5111 1489 5720 1534
rect 5772 1489 5799 1534
rect 5851 1489 5878 1541
rect 5930 1534 5961 1541
rect 5995 1534 6034 1568
rect 6068 1534 6107 1568
rect 6141 1534 6180 1568
rect 6214 1534 6253 1568
rect 6287 1534 6326 1568
rect 6360 1534 6399 1568
rect 6433 1534 6472 1568
rect 6549 1561 6574 1613
rect 6626 1561 6651 1613
rect 6703 1561 6728 1613
rect 6780 1561 6805 1613
rect 6882 1606 6921 1640
rect 6955 1606 6994 1640
rect 7028 1606 7067 1640
rect 7101 1606 7140 1640
rect 7174 1606 7213 1640
rect 7247 1606 7286 1640
rect 7320 1606 7359 1640
rect 7393 1606 7432 1640
rect 7466 1606 7505 1640
rect 7539 1606 7578 1640
rect 7612 1606 7651 1640
rect 7685 1606 7724 1640
rect 7758 1606 7797 1640
rect 7831 1606 7870 1640
rect 7904 1606 7943 1640
rect 7977 1606 8016 1640
rect 8050 1606 8089 1640
rect 8123 1606 8162 1640
rect 8196 1606 8235 1640
rect 8269 1606 8308 1640
rect 8342 1606 8382 1640
rect 8416 1606 8456 1640
rect 8490 1606 8530 1640
rect 8564 1606 8604 1640
rect 8638 1606 8678 1640
rect 8712 1606 8752 1640
rect 8786 1606 8826 1640
rect 8860 1606 8900 1640
rect 8934 1606 8974 1640
rect 9008 1606 9048 1640
rect 9082 1606 9122 1640
rect 9156 1606 9196 1640
rect 9230 1606 9270 1640
rect 9304 1606 9344 1640
rect 9378 1606 9418 1640
rect 9452 1606 9492 1640
rect 9711 1633 9714 1640
rect 9778 1633 10090 1640
rect 9526 1613 9566 1633
rect 9600 1613 9640 1633
rect 9674 1613 9714 1633
rect 9748 1613 10090 1633
rect 9711 1606 9714 1613
rect 9778 1606 10090 1613
rect 10124 1606 10164 1640
rect 10198 1606 10238 1640
rect 10272 1606 10312 1640
rect 10346 1606 10386 1640
rect 10420 1606 10460 1640
rect 10494 1606 10534 1640
rect 10568 1606 10608 1640
rect 10642 1606 10682 1640
rect 10716 1606 10756 1640
rect 10790 1606 10830 1640
rect 10864 1606 10904 1640
rect 10938 1606 10978 1640
rect 11012 1606 11052 1640
rect 11086 1606 11126 1640
rect 11160 1606 11200 1640
rect 11234 1606 11274 1640
rect 11308 1606 11348 1640
rect 11382 1606 11422 1640
rect 11456 1606 11496 1640
rect 11530 1606 11569 1640
rect 11603 1606 11642 1640
rect 11676 1606 11715 1640
rect 11749 1606 11788 1640
rect 11822 1606 11861 1640
rect 11895 1606 11934 1640
rect 11968 1606 12007 1640
rect 12041 1606 12080 1640
rect 12114 1606 12153 1640
rect 12187 1606 12226 1640
rect 12260 1606 12299 1640
rect 12333 1606 12372 1640
rect 12406 1606 12445 1640
rect 12479 1606 12518 1640
rect 12552 1606 12591 1640
rect 12625 1606 12664 1640
rect 12698 1606 12737 1640
rect 12771 1606 12810 1640
rect 12844 1606 12883 1640
rect 12917 1606 12956 1640
rect 12990 1606 13332 1640
rect 13366 1606 13405 1640
rect 13439 1606 13478 1640
rect 13512 1606 13551 1640
rect 13585 1606 13624 1640
rect 13658 1606 13697 1640
rect 13731 1606 13770 1640
rect 13804 1606 13843 1640
rect 13877 1606 13916 1640
rect 13950 1606 13989 1640
rect 14023 1606 14062 1640
rect 14096 1606 14135 1640
rect 14169 1606 14208 1640
rect 14242 1606 14281 1640
rect 14315 1606 14354 1640
rect 14388 1606 14427 1640
rect 14461 1606 14500 1640
rect 14534 1606 14573 1640
rect 14607 1606 14646 1640
rect 14680 1606 14719 1640
rect 14753 1606 14792 1640
rect 14826 1606 14866 1640
rect 14900 1606 14940 1640
rect 14974 1606 15014 1640
rect 15048 1606 15088 1640
rect 15122 1606 15162 1640
rect 15196 1606 15236 1640
rect 15270 1606 15310 1640
rect 15344 1606 15384 1640
rect 15418 1606 15458 1640
rect 15492 1606 15532 1640
rect 15566 1606 15606 1640
rect 15640 1606 15680 1640
rect 15714 1606 15754 1640
rect 15788 1606 15828 1640
rect 15862 1606 15902 1640
rect 15936 1606 15976 1640
rect 16010 1606 16050 1640
rect 16084 1606 16124 1640
rect 16158 1606 16198 1640
rect 16232 1633 16403 1640
rect 16455 1633 16471 1685
rect 16523 1633 16539 1685
rect 16591 1640 16607 1685
rect 16659 1640 16674 1685
rect 16726 1640 16741 1685
rect 16793 1671 19528 1685
tri 19528 1671 19543 1686 sw
rect 19841 1671 19882 1705
rect 19916 1671 19971 1705
rect 16793 1640 19543 1671
tri 19543 1640 19574 1671 sw
rect 16793 1633 16796 1640
rect 16232 1613 16574 1633
rect 16608 1613 16648 1633
rect 16682 1613 16722 1633
rect 16756 1613 16796 1633
rect 16232 1606 16403 1613
rect 6857 1568 9525 1606
rect 9577 1568 9592 1606
rect 9644 1568 9659 1606
rect 9711 1568 9726 1606
rect 9778 1568 16403 1606
rect 6506 1541 6848 1561
rect 5930 1489 6497 1534
rect 6549 1489 6574 1541
rect 6626 1489 6651 1541
rect 6703 1489 6728 1541
rect 6780 1489 6805 1541
rect 6882 1534 6921 1568
rect 6955 1534 6994 1568
rect 7028 1534 7067 1568
rect 7101 1534 7140 1568
rect 7174 1534 7213 1568
rect 7247 1534 7286 1568
rect 7320 1534 7359 1568
rect 7393 1534 7432 1568
rect 7466 1534 7505 1568
rect 7539 1534 7578 1568
rect 7612 1534 7651 1568
rect 7685 1534 7724 1568
rect 7758 1534 7797 1568
rect 7831 1534 7870 1568
rect 7904 1534 7943 1568
rect 7977 1534 8016 1568
rect 8050 1534 8089 1568
rect 8123 1534 8162 1568
rect 8196 1534 8235 1568
rect 8269 1534 8308 1568
rect 8342 1534 8382 1568
rect 8416 1534 8456 1568
rect 8490 1534 8530 1568
rect 8564 1534 8604 1568
rect 8638 1534 8678 1568
rect 8712 1534 8752 1568
rect 8786 1534 8826 1568
rect 8860 1534 8900 1568
rect 8934 1534 8974 1568
rect 9008 1534 9048 1568
rect 9082 1534 9122 1568
rect 9156 1534 9196 1568
rect 9230 1534 9270 1568
rect 9304 1534 9344 1568
rect 9378 1534 9418 1568
rect 9452 1534 9492 1568
rect 9711 1561 9714 1568
rect 9778 1561 10090 1568
rect 9526 1541 9566 1561
rect 9600 1541 9640 1561
rect 9674 1541 9714 1561
rect 9748 1541 10090 1561
rect 9711 1534 9714 1541
rect 9778 1534 10090 1541
rect 10124 1534 10164 1568
rect 10198 1534 10238 1568
rect 10272 1534 10312 1568
rect 10346 1534 10386 1568
rect 10420 1534 10460 1568
rect 10494 1534 10534 1568
rect 10568 1534 10608 1568
rect 10642 1534 10682 1568
rect 10716 1534 10756 1568
rect 10790 1534 10830 1568
rect 10864 1534 10904 1568
rect 10938 1534 10978 1568
rect 11012 1534 11052 1568
rect 11086 1534 11126 1568
rect 11160 1534 11200 1568
rect 11234 1534 11274 1568
rect 11308 1534 11348 1568
rect 11382 1534 11422 1568
rect 11456 1534 11496 1568
rect 11530 1534 11569 1568
rect 11603 1534 11642 1568
rect 11676 1534 11715 1568
rect 11749 1534 11788 1568
rect 11822 1534 11861 1568
rect 11895 1534 11934 1568
rect 11968 1534 12007 1568
rect 12041 1534 12080 1568
rect 12114 1534 12153 1568
rect 12187 1534 12226 1568
rect 12260 1534 12299 1568
rect 12333 1534 12372 1568
rect 12406 1534 12445 1568
rect 12479 1534 12518 1568
rect 12552 1534 12591 1568
rect 12625 1534 12664 1568
rect 12698 1534 12737 1568
rect 12771 1534 12810 1568
rect 12844 1534 12883 1568
rect 12917 1534 12956 1568
rect 12990 1534 13332 1568
rect 13366 1534 13405 1568
rect 13439 1534 13478 1568
rect 13512 1534 13551 1568
rect 13585 1534 13624 1568
rect 13658 1534 13697 1568
rect 13731 1534 13770 1568
rect 13804 1534 13843 1568
rect 13877 1534 13916 1568
rect 13950 1534 13989 1568
rect 14023 1534 14062 1568
rect 14096 1534 14135 1568
rect 14169 1534 14208 1568
rect 14242 1534 14281 1568
rect 14315 1534 14354 1568
rect 14388 1534 14427 1568
rect 14461 1534 14500 1568
rect 14534 1534 14573 1568
rect 14607 1534 14646 1568
rect 14680 1534 14719 1568
rect 14753 1534 14792 1568
rect 14826 1534 14866 1568
rect 14900 1534 14940 1568
rect 14974 1534 15014 1568
rect 15048 1534 15088 1568
rect 15122 1534 15162 1568
rect 15196 1534 15236 1568
rect 15270 1534 15310 1568
rect 15344 1534 15384 1568
rect 15418 1534 15458 1568
rect 15492 1534 15532 1568
rect 15566 1534 15606 1568
rect 15640 1534 15680 1568
rect 15714 1534 15754 1568
rect 15788 1534 15828 1568
rect 15862 1534 15902 1568
rect 15936 1534 15976 1568
rect 16010 1534 16050 1568
rect 16084 1534 16124 1568
rect 16158 1534 16198 1568
rect 16232 1561 16403 1568
rect 16455 1561 16471 1613
rect 16523 1561 16539 1613
rect 16793 1606 16796 1613
rect 16830 1606 16870 1640
rect 16904 1606 16944 1640
rect 16978 1606 17018 1640
rect 17052 1606 17092 1640
rect 17126 1606 17166 1640
rect 17200 1606 17240 1640
rect 17274 1606 17314 1640
rect 17348 1606 17388 1640
rect 17422 1606 17462 1640
rect 17496 1606 17536 1640
rect 17570 1606 17610 1640
rect 17644 1606 17684 1640
rect 17718 1606 17758 1640
rect 17792 1606 17832 1640
rect 17866 1606 17906 1640
rect 17940 1606 17980 1640
rect 18014 1606 18053 1640
rect 18087 1606 18126 1640
rect 18160 1606 18199 1640
rect 18233 1606 18272 1640
rect 18306 1606 18345 1640
rect 18379 1606 18418 1640
rect 18452 1606 18491 1640
rect 18525 1606 18564 1640
rect 18598 1606 18637 1640
rect 18671 1606 18710 1640
rect 18744 1606 18783 1640
rect 18817 1606 18856 1640
rect 18890 1606 18929 1640
rect 18963 1606 19002 1640
rect 19036 1606 19075 1640
rect 19109 1606 19148 1640
rect 19182 1606 19221 1640
rect 19255 1606 19294 1640
rect 19328 1606 19367 1640
rect 19401 1606 19440 1640
rect 19474 1606 19574 1640
rect 16591 1568 16607 1606
rect 16659 1568 16674 1606
rect 16726 1568 16741 1606
rect 16793 1568 19574 1606
rect 16793 1561 16796 1568
rect 16232 1541 16574 1561
rect 16608 1541 16648 1561
rect 16682 1541 16722 1561
rect 16756 1541 16796 1561
rect 16232 1534 16403 1541
rect 6857 1489 9525 1534
rect 9577 1489 9592 1534
rect 9644 1489 9659 1534
rect 9711 1489 9726 1534
rect 9778 1525 9839 1534
tri 9839 1525 9848 1534 nw
tri 9990 1525 9999 1534 ne
rect 9999 1525 13081 1534
tri 13081 1525 13090 1534 nw
tri 13232 1525 13241 1534 ne
rect 13241 1525 16323 1534
tri 16323 1525 16332 1534 nw
rect 9778 1489 9802 1525
rect 310 1488 9802 1489
tri 9802 1488 9839 1525 nw
tri 9999 1496 10028 1525 ne
rect 10028 1496 13044 1525
rect 9897 1490 9949 1496
tri 310 1487 311 1488 ne
rect 311 1487 3317 1488
tri 3317 1487 3318 1488 nw
tri 3552 1487 3553 1488 ne
rect 3553 1487 6559 1488
tri 6559 1487 6560 1488 nw
tri 6794 1487 6795 1488 ne
rect 6795 1487 9801 1488
tri 9801 1487 9802 1488 nw
rect -52 1445 -46 1479
rect -12 1445 42 1479
rect 76 1445 82 1479
rect 3370 1452 3376 1455
rect -578 1405 -522 1410
tri -522 1405 -517 1410 nw
rect -52 1405 82 1445
rect 156 1446 3376 1452
rect 156 1412 168 1446
rect 202 1439 240 1446
rect 228 1412 240 1439
rect 274 1412 3376 1446
rect 156 1406 176 1412
rect -578 1387 -546 1405
rect -630 1381 -546 1387
tri -546 1381 -522 1405 nw
rect -52 1371 -46 1405
rect -12 1371 42 1405
rect 76 1371 82 1405
rect -52 1331 82 1371
rect -52 1297 -46 1331
rect -12 1297 42 1331
rect 76 1297 82 1331
rect 228 1406 3376 1412
rect 3370 1403 3376 1406
rect 3428 1403 3440 1455
rect 3492 1452 3498 1455
rect 3492 1406 6648 1452
rect 6649 1407 6650 1451
rect 6710 1407 6711 1451
rect 6712 1446 9897 1452
tri 10028 1488 10036 1496 ne
rect 10036 1488 13044 1496
tri 13044 1488 13081 1525 nw
tri 13241 1488 13278 1525 ne
rect 13278 1488 16286 1525
tri 16286 1488 16323 1525 nw
rect 16397 1489 16403 1534
rect 16455 1489 16471 1541
rect 16523 1489 16539 1541
rect 16793 1534 16796 1541
rect 16830 1534 16870 1568
rect 16904 1534 16944 1568
rect 16978 1534 17018 1568
rect 17052 1534 17092 1568
rect 17126 1534 17166 1568
rect 17200 1534 17240 1568
rect 17274 1534 17314 1568
rect 17348 1534 17388 1568
rect 17422 1534 17462 1568
rect 17496 1534 17536 1568
rect 17570 1534 17610 1568
rect 17644 1534 17684 1568
rect 17718 1534 17758 1568
rect 17792 1534 17832 1568
rect 17866 1534 17906 1568
rect 17940 1534 17980 1568
rect 18014 1534 18053 1568
rect 18087 1534 18126 1568
rect 18160 1534 18199 1568
rect 18233 1534 18272 1568
rect 18306 1534 18345 1568
rect 18379 1534 18418 1568
rect 18452 1534 18491 1568
rect 18525 1534 18564 1568
rect 18598 1534 18637 1568
rect 18671 1534 18710 1568
rect 18744 1534 18783 1568
rect 18817 1534 18856 1568
rect 18890 1534 18929 1568
rect 18963 1534 19002 1568
rect 19036 1534 19075 1568
rect 19109 1534 19148 1568
rect 19182 1534 19221 1568
rect 19255 1534 19294 1568
rect 19328 1534 19367 1568
rect 19401 1534 19440 1568
rect 19474 1534 19574 1568
rect 16591 1489 16607 1534
rect 16659 1489 16674 1534
rect 16726 1489 16741 1534
rect 16793 1525 19565 1534
tri 19565 1525 19574 1534 nw
rect 19841 1632 19971 1671
rect 19841 1598 19882 1632
rect 19916 1598 19971 1632
rect 19841 1559 19971 1598
rect 19841 1525 19882 1559
rect 19916 1525 19971 1559
rect 16793 1489 19528 1525
rect 16397 1488 19528 1489
tri 19528 1488 19565 1525 nw
tri 10036 1487 10037 1488 ne
rect 10037 1487 13043 1488
tri 13043 1487 13044 1488 nw
tri 13278 1487 13279 1488 ne
rect 13279 1487 16285 1488
tri 16285 1487 16286 1488 nw
tri 16520 1487 16521 1488 ne
rect 16521 1487 19527 1488
tri 19527 1487 19528 1488 nw
rect 19841 1486 19971 1525
rect 19841 1452 19882 1486
rect 19916 1452 19971 1486
rect 9949 1446 13113 1452
rect 6712 1412 9870 1446
rect 9904 1426 9942 1438
rect 9976 1412 13113 1446
rect 6712 1406 9897 1412
rect 3492 1403 3498 1406
rect 176 1375 228 1387
tri 276 1340 311 1375 se
rect 311 1371 3317 1375
rect 311 1340 1027 1371
rect 176 1317 228 1323
tri 264 1328 276 1340 se
rect 276 1328 1027 1340
rect 264 1319 1027 1328
rect 1079 1319 1092 1371
rect 1144 1319 1157 1371
rect 1209 1319 1222 1371
rect 1274 1319 1286 1371
rect 1338 1319 1350 1371
rect 1402 1319 1414 1371
rect 1466 1319 1478 1371
rect 1530 1319 1542 1371
rect 1594 1319 1606 1371
rect 1658 1319 1670 1371
rect 1722 1319 1734 1371
rect 1786 1319 1798 1371
rect 1850 1319 1862 1371
rect 1914 1340 3317 1371
tri 3317 1340 3352 1375 sw
tri 3518 1340 3553 1375 se
rect 3553 1371 6559 1375
rect 3553 1340 5199 1371
rect 1914 1328 3352 1340
tri 3352 1328 3364 1340 sw
tri 3506 1328 3518 1340 se
rect 3518 1328 5199 1340
rect 1914 1319 5199 1328
rect 5251 1319 5263 1371
rect 5315 1319 5327 1371
rect 5379 1319 5392 1371
rect 5444 1319 5457 1371
rect 5509 1319 5522 1371
rect 5574 1319 5587 1371
rect 5639 1340 6559 1371
tri 6559 1340 6594 1375 sw
tri 6760 1340 6795 1375 se
rect 6795 1371 9801 1375
rect 6795 1340 7511 1371
rect 5639 1328 6594 1340
tri 6594 1328 6606 1340 sw
tri 6748 1328 6760 1340 se
rect 6760 1328 7511 1340
rect 5639 1319 7511 1328
rect 7563 1319 7576 1371
rect 7628 1319 7641 1371
rect 7693 1319 7706 1371
rect 7758 1319 7770 1371
rect 7822 1319 7834 1371
rect 7886 1319 7898 1371
rect 7950 1319 7962 1371
rect 8014 1319 8026 1371
rect 8078 1319 8090 1371
rect 8142 1319 8154 1371
rect 8206 1319 8218 1371
rect 8270 1319 8282 1371
rect 8334 1319 8346 1371
rect 8398 1340 9801 1371
tri 9801 1340 9836 1375 sw
rect 9949 1406 13113 1412
rect 13209 1446 19706 1452
rect 13209 1412 16354 1446
rect 16388 1412 16426 1446
rect 16460 1412 19564 1446
rect 19598 1412 19636 1446
rect 19670 1412 19706 1446
rect 13209 1406 19706 1412
rect 19610 1396 19706 1406
rect 9897 1368 9949 1374
tri 10030 1368 10037 1375 se
rect 10037 1371 13043 1375
rect 10037 1368 11440 1371
tri 10002 1340 10030 1368 se
rect 10030 1340 11440 1368
rect 8398 1328 9836 1340
tri 9836 1328 9848 1340 sw
tri 9990 1328 10002 1340 se
rect 10002 1328 11440 1340
rect 8398 1319 11440 1328
rect 11492 1319 11504 1371
rect 11556 1319 11568 1371
rect 11620 1319 11632 1371
rect 11684 1319 11696 1371
rect 11748 1319 11760 1371
rect 11812 1319 11824 1371
rect 11876 1319 11888 1371
rect 11940 1319 11952 1371
rect 12004 1319 12016 1371
rect 12068 1319 12080 1371
rect 12132 1319 12145 1371
rect 12197 1319 12210 1371
rect 12262 1319 12275 1371
rect 12327 1340 13043 1371
tri 13043 1340 13078 1375 sw
tri 13244 1340 13279 1375 se
rect 13279 1371 16285 1375
rect 13279 1340 13995 1371
rect 12327 1328 13078 1340
tri 13078 1328 13090 1340 sw
tri 13232 1328 13244 1340 se
rect 13244 1328 13995 1340
rect 12327 1319 13995 1328
rect 14047 1319 14060 1371
rect 14112 1319 14125 1371
rect 14177 1319 14190 1371
rect 14242 1319 14254 1371
rect 14306 1319 14318 1371
rect 14370 1319 14382 1371
rect 14434 1319 14446 1371
rect 14498 1319 14510 1371
rect 14562 1319 14574 1371
rect 14626 1319 14638 1371
rect 14690 1319 14702 1371
rect 14754 1319 14766 1371
rect 14818 1319 14830 1371
rect 14882 1340 16285 1371
tri 16285 1340 16320 1375 sw
tri 16486 1340 16521 1375 se
rect 16521 1371 19527 1375
rect 16521 1340 17924 1371
rect 14882 1328 16320 1340
tri 16320 1328 16332 1340 sw
tri 16474 1328 16486 1340 se
rect 16486 1328 17924 1340
rect 14882 1319 17924 1328
rect 17976 1319 17988 1371
rect 18040 1319 18052 1371
rect 18104 1319 18116 1371
rect 18168 1319 18180 1371
rect 18232 1319 18244 1371
rect 18296 1319 18308 1371
rect 18360 1319 18372 1371
rect 18424 1319 18436 1371
rect 18488 1319 18500 1371
rect 18552 1319 18564 1371
rect 18616 1319 18629 1371
rect 18681 1319 18694 1371
rect 18746 1319 18759 1371
rect 18811 1340 19527 1371
tri 19527 1340 19562 1375 sw
rect 19662 1344 19706 1396
rect 18811 1328 19562 1340
tri 19562 1328 19574 1340 sw
rect 18811 1319 19574 1328
rect -52 1257 82 1297
rect -52 1223 -46 1257
rect -12 1223 42 1257
rect 76 1223 82 1257
rect -52 1183 82 1223
rect -52 1149 -46 1183
rect -12 1149 42 1183
rect 76 1149 82 1183
rect -52 1109 82 1149
rect -52 1075 -46 1109
rect -12 1075 42 1109
rect 76 1075 82 1109
rect -52 1035 82 1075
rect -52 1001 -46 1035
rect -12 1001 42 1035
rect 76 1001 82 1035
rect 264 1303 19574 1319
rect 264 1251 1027 1303
rect 1079 1251 1092 1303
rect 1144 1251 1157 1303
rect 1209 1251 1222 1303
rect 1274 1251 1286 1303
rect 1338 1251 1350 1303
rect 1402 1251 1414 1303
rect 1466 1251 1478 1303
rect 1530 1251 1542 1303
rect 1594 1251 1606 1303
rect 1658 1251 1670 1303
rect 1722 1251 1734 1303
rect 1786 1251 1798 1303
rect 1850 1251 1862 1303
rect 1914 1251 5199 1303
rect 5251 1251 5263 1303
rect 5315 1251 5327 1303
rect 5379 1251 5392 1303
rect 5444 1251 5457 1303
rect 5509 1251 5522 1303
rect 5574 1251 5587 1303
rect 5639 1251 7511 1303
rect 7563 1251 7576 1303
rect 7628 1251 7641 1303
rect 7693 1251 7706 1303
rect 7758 1251 7770 1303
rect 7822 1251 7834 1303
rect 7886 1251 7898 1303
rect 7950 1251 7962 1303
rect 8014 1251 8026 1303
rect 8078 1251 8090 1303
rect 8142 1251 8154 1303
rect 8206 1251 8218 1303
rect 8270 1251 8282 1303
rect 8334 1251 8346 1303
rect 8398 1251 11440 1303
rect 11492 1251 11504 1303
rect 11556 1251 11568 1303
rect 11620 1251 11632 1303
rect 11684 1251 11696 1303
rect 11748 1251 11760 1303
rect 11812 1251 11824 1303
rect 11876 1251 11888 1303
rect 11940 1251 11952 1303
rect 12004 1251 12016 1303
rect 12068 1251 12080 1303
rect 12132 1251 12145 1303
rect 12197 1251 12210 1303
rect 12262 1251 12275 1303
rect 12327 1251 13995 1303
rect 14047 1251 14060 1303
rect 14112 1251 14125 1303
rect 14177 1251 14190 1303
rect 14242 1251 14254 1303
rect 14306 1251 14318 1303
rect 14370 1251 14382 1303
rect 14434 1251 14446 1303
rect 14498 1251 14510 1303
rect 14562 1251 14574 1303
rect 14626 1251 14638 1303
rect 14690 1251 14702 1303
rect 14754 1251 14766 1303
rect 14818 1251 14830 1303
rect 14882 1251 17924 1303
rect 17976 1251 17988 1303
rect 18040 1251 18052 1303
rect 18104 1251 18116 1303
rect 18168 1251 18180 1303
rect 18232 1251 18244 1303
rect 18296 1251 18308 1303
rect 18360 1251 18372 1303
rect 18424 1251 18436 1303
rect 18488 1251 18500 1303
rect 18552 1251 18564 1303
rect 18616 1251 18629 1303
rect 18681 1251 18694 1303
rect 18746 1251 18759 1303
rect 18811 1251 19574 1303
rect 19610 1332 19706 1344
rect 19662 1280 19706 1332
rect 19610 1274 19706 1280
rect 19841 1413 19971 1452
rect 19841 1379 19882 1413
rect 19916 1379 19971 1413
rect 19841 1340 19971 1379
rect 19841 1306 19882 1340
rect 19916 1306 19971 1340
rect 264 1235 19574 1251
rect 264 1228 1027 1235
rect 264 1194 364 1228
rect 398 1194 437 1228
rect 471 1194 510 1228
rect 544 1194 583 1228
rect 617 1194 656 1228
rect 690 1194 729 1228
rect 763 1194 802 1228
rect 836 1194 875 1228
rect 909 1194 948 1228
rect 982 1194 1021 1228
rect 264 1183 1027 1194
rect 1079 1183 1092 1235
rect 1144 1183 1157 1235
rect 1209 1183 1222 1235
rect 1274 1183 1286 1235
rect 1338 1228 1350 1235
rect 1402 1228 1414 1235
rect 1466 1228 1478 1235
rect 1530 1228 1542 1235
rect 1594 1228 1606 1235
rect 1347 1194 1350 1228
rect 1530 1194 1532 1228
rect 1594 1194 1605 1228
rect 1338 1183 1350 1194
rect 1402 1183 1414 1194
rect 1466 1183 1478 1194
rect 1530 1183 1542 1194
rect 1594 1183 1606 1194
rect 1658 1183 1670 1235
rect 1722 1183 1734 1235
rect 1786 1183 1798 1235
rect 1850 1228 1862 1235
rect 1914 1228 5199 1235
rect 5251 1228 5263 1235
rect 5315 1228 5327 1235
rect 5379 1228 5392 1235
rect 5444 1228 5457 1235
rect 1858 1194 1862 1228
rect 1932 1194 1972 1228
rect 2006 1194 2046 1228
rect 2080 1194 2120 1228
rect 2154 1194 2194 1228
rect 2228 1194 2268 1228
rect 2302 1194 2342 1228
rect 2376 1194 2416 1228
rect 2450 1194 2490 1228
rect 2524 1194 2564 1228
rect 2598 1194 2638 1228
rect 2672 1194 2712 1228
rect 2746 1194 2786 1228
rect 2820 1194 2860 1228
rect 2894 1194 2934 1228
rect 2968 1194 3008 1228
rect 3042 1194 3082 1228
rect 3116 1194 3156 1228
rect 3190 1194 3230 1228
rect 3264 1194 3606 1228
rect 3640 1194 3680 1228
rect 3714 1194 3754 1228
rect 3788 1194 3828 1228
rect 3862 1194 3902 1228
rect 3936 1194 3976 1228
rect 4010 1194 4050 1228
rect 4084 1194 4124 1228
rect 4158 1194 4198 1228
rect 4232 1194 4272 1228
rect 4306 1194 4346 1228
rect 4380 1194 4420 1228
rect 4454 1194 4494 1228
rect 4528 1194 4568 1228
rect 4602 1194 4642 1228
rect 4676 1194 4716 1228
rect 4750 1194 4790 1228
rect 4824 1194 4864 1228
rect 4898 1194 4938 1228
rect 4972 1194 5012 1228
rect 5046 1194 5085 1228
rect 5119 1194 5158 1228
rect 5192 1194 5199 1228
rect 5444 1194 5450 1228
rect 1850 1183 1862 1194
rect 1914 1183 5199 1194
rect 5251 1183 5263 1194
rect 5315 1183 5327 1194
rect 5379 1183 5392 1194
rect 5444 1183 5457 1194
rect 5509 1183 5522 1235
rect 5574 1183 5587 1235
rect 5639 1228 7511 1235
rect 5639 1194 5669 1228
rect 5703 1194 5742 1228
rect 5776 1194 5815 1228
rect 5849 1194 5888 1228
rect 5922 1194 5961 1228
rect 5995 1194 6034 1228
rect 6068 1194 6107 1228
rect 6141 1194 6180 1228
rect 6214 1194 6253 1228
rect 6287 1194 6326 1228
rect 6360 1194 6399 1228
rect 6433 1194 6472 1228
rect 6506 1194 6848 1228
rect 6882 1194 6921 1228
rect 6955 1194 6994 1228
rect 7028 1194 7067 1228
rect 7101 1194 7140 1228
rect 7174 1194 7213 1228
rect 7247 1194 7286 1228
rect 7320 1194 7359 1228
rect 7393 1194 7432 1228
rect 7466 1194 7505 1228
rect 5639 1183 7511 1194
rect 7563 1183 7576 1235
rect 7628 1183 7641 1235
rect 7693 1183 7706 1235
rect 7758 1183 7770 1235
rect 7822 1228 7834 1235
rect 7886 1228 7898 1235
rect 7950 1228 7962 1235
rect 8014 1228 8026 1235
rect 8078 1228 8090 1235
rect 7831 1194 7834 1228
rect 8014 1194 8016 1228
rect 8078 1194 8089 1228
rect 7822 1183 7834 1194
rect 7886 1183 7898 1194
rect 7950 1183 7962 1194
rect 8014 1183 8026 1194
rect 8078 1183 8090 1194
rect 8142 1183 8154 1235
rect 8206 1183 8218 1235
rect 8270 1183 8282 1235
rect 8334 1228 8346 1235
rect 8398 1228 11440 1235
rect 11492 1228 11504 1235
rect 8342 1194 8346 1228
rect 8416 1194 8456 1228
rect 8490 1194 8530 1228
rect 8564 1194 8604 1228
rect 8638 1194 8678 1228
rect 8712 1194 8752 1228
rect 8786 1194 8826 1228
rect 8860 1194 8900 1228
rect 8934 1194 8974 1228
rect 9008 1194 9048 1228
rect 9082 1194 9122 1228
rect 9156 1194 9196 1228
rect 9230 1194 9270 1228
rect 9304 1194 9344 1228
rect 9378 1194 9418 1228
rect 9452 1194 9492 1228
rect 9526 1194 9566 1228
rect 9600 1194 9640 1228
rect 9674 1194 9714 1228
rect 9748 1194 10090 1228
rect 10124 1194 10164 1228
rect 10198 1194 10238 1228
rect 10272 1194 10312 1228
rect 10346 1194 10386 1228
rect 10420 1194 10460 1228
rect 10494 1194 10534 1228
rect 10568 1194 10608 1228
rect 10642 1194 10682 1228
rect 10716 1194 10756 1228
rect 10790 1194 10830 1228
rect 10864 1194 10904 1228
rect 10938 1194 10978 1228
rect 11012 1194 11052 1228
rect 11086 1194 11126 1228
rect 11160 1194 11200 1228
rect 11234 1194 11274 1228
rect 11308 1194 11348 1228
rect 11382 1194 11422 1228
rect 11492 1194 11496 1228
rect 8334 1183 8346 1194
rect 8398 1183 11440 1194
rect 11492 1183 11504 1194
rect 11556 1183 11568 1235
rect 11620 1183 11632 1235
rect 11684 1183 11696 1235
rect 11748 1228 11760 1235
rect 11812 1228 11824 1235
rect 11876 1228 11888 1235
rect 11940 1228 11952 1235
rect 12004 1228 12016 1235
rect 11749 1194 11760 1228
rect 11822 1194 11824 1228
rect 12004 1194 12007 1228
rect 11748 1183 11760 1194
rect 11812 1183 11824 1194
rect 11876 1183 11888 1194
rect 11940 1183 11952 1194
rect 12004 1183 12016 1194
rect 12068 1183 12080 1235
rect 12132 1183 12145 1235
rect 12197 1183 12210 1235
rect 12262 1183 12275 1235
rect 12327 1228 13995 1235
rect 12333 1194 12372 1228
rect 12406 1194 12445 1228
rect 12479 1194 12518 1228
rect 12552 1194 12591 1228
rect 12625 1194 12664 1228
rect 12698 1194 12737 1228
rect 12771 1194 12810 1228
rect 12844 1194 12883 1228
rect 12917 1194 12956 1228
rect 12990 1194 13332 1228
rect 13366 1194 13405 1228
rect 13439 1194 13478 1228
rect 13512 1194 13551 1228
rect 13585 1194 13624 1228
rect 13658 1194 13697 1228
rect 13731 1194 13770 1228
rect 13804 1194 13843 1228
rect 13877 1194 13916 1228
rect 13950 1194 13989 1228
rect 12327 1183 13995 1194
rect 14047 1183 14060 1235
rect 14112 1183 14125 1235
rect 14177 1183 14190 1235
rect 14242 1183 14254 1235
rect 14306 1228 14318 1235
rect 14370 1228 14382 1235
rect 14434 1228 14446 1235
rect 14498 1228 14510 1235
rect 14562 1228 14574 1235
rect 14315 1194 14318 1228
rect 14498 1194 14500 1228
rect 14562 1194 14573 1228
rect 14306 1183 14318 1194
rect 14370 1183 14382 1194
rect 14434 1183 14446 1194
rect 14498 1183 14510 1194
rect 14562 1183 14574 1194
rect 14626 1183 14638 1235
rect 14690 1183 14702 1235
rect 14754 1183 14766 1235
rect 14818 1228 14830 1235
rect 14882 1228 17924 1235
rect 17976 1228 17988 1235
rect 14826 1194 14830 1228
rect 14900 1194 14940 1228
rect 14974 1194 15014 1228
rect 15048 1194 15088 1228
rect 15122 1194 15162 1228
rect 15196 1194 15236 1228
rect 15270 1194 15310 1228
rect 15344 1194 15384 1228
rect 15418 1194 15458 1228
rect 15492 1194 15532 1228
rect 15566 1194 15606 1228
rect 15640 1194 15680 1228
rect 15714 1194 15754 1228
rect 15788 1194 15828 1228
rect 15862 1194 15902 1228
rect 15936 1194 15976 1228
rect 16010 1194 16050 1228
rect 16084 1194 16124 1228
rect 16158 1194 16198 1228
rect 16232 1194 16574 1228
rect 16608 1194 16648 1228
rect 16682 1194 16722 1228
rect 16756 1194 16796 1228
rect 16830 1194 16870 1228
rect 16904 1194 16944 1228
rect 16978 1194 17018 1228
rect 17052 1194 17092 1228
rect 17126 1194 17166 1228
rect 17200 1194 17240 1228
rect 17274 1194 17314 1228
rect 17348 1194 17388 1228
rect 17422 1194 17462 1228
rect 17496 1194 17536 1228
rect 17570 1194 17610 1228
rect 17644 1194 17684 1228
rect 17718 1194 17758 1228
rect 17792 1194 17832 1228
rect 17866 1194 17906 1228
rect 17976 1194 17980 1228
rect 14818 1183 14830 1194
rect 14882 1183 17924 1194
rect 17976 1183 17988 1194
rect 18040 1183 18052 1235
rect 18104 1183 18116 1235
rect 18168 1183 18180 1235
rect 18232 1228 18244 1235
rect 18296 1228 18308 1235
rect 18360 1228 18372 1235
rect 18424 1228 18436 1235
rect 18488 1228 18500 1235
rect 18233 1194 18244 1228
rect 18306 1194 18308 1228
rect 18488 1194 18491 1228
rect 18232 1183 18244 1194
rect 18296 1183 18308 1194
rect 18360 1183 18372 1194
rect 18424 1183 18436 1194
rect 18488 1183 18500 1194
rect 18552 1183 18564 1235
rect 18616 1183 18629 1235
rect 18681 1183 18694 1235
rect 18746 1183 18759 1235
rect 18811 1228 19574 1235
rect 18817 1194 18856 1228
rect 18890 1194 18929 1228
rect 18963 1194 19002 1228
rect 19036 1194 19075 1228
rect 19109 1194 19148 1228
rect 19182 1194 19221 1228
rect 19255 1194 19294 1228
rect 19328 1194 19367 1228
rect 19401 1194 19440 1228
rect 19474 1194 19574 1228
rect 19841 1267 19971 1306
rect 19841 1233 19882 1267
rect 19916 1233 19971 1267
rect 18811 1183 19574 1194
rect 264 1167 19574 1183
rect 264 1156 1027 1167
rect 264 1122 364 1156
rect 398 1122 437 1156
rect 471 1122 510 1156
rect 544 1122 583 1156
rect 617 1122 656 1156
rect 690 1122 729 1156
rect 763 1122 802 1156
rect 836 1122 875 1156
rect 909 1122 948 1156
rect 982 1122 1021 1156
rect 264 1115 1027 1122
rect 1079 1115 1092 1167
rect 1144 1115 1157 1167
rect 1209 1115 1222 1167
rect 1274 1115 1286 1167
rect 1338 1156 1350 1167
rect 1402 1156 1414 1167
rect 1466 1156 1478 1167
rect 1530 1156 1542 1167
rect 1594 1156 1606 1167
rect 1347 1122 1350 1156
rect 1530 1122 1532 1156
rect 1594 1122 1605 1156
rect 1338 1115 1350 1122
rect 1402 1115 1414 1122
rect 1466 1115 1478 1122
rect 1530 1115 1542 1122
rect 1594 1115 1606 1122
rect 1658 1115 1670 1167
rect 1722 1115 1734 1167
rect 1786 1115 1798 1167
rect 1850 1156 1862 1167
rect 1914 1156 5199 1167
rect 5251 1156 5263 1167
rect 5315 1156 5327 1167
rect 5379 1156 5392 1167
rect 5444 1156 5457 1167
rect 1858 1122 1862 1156
rect 1932 1122 1972 1156
rect 2006 1122 2046 1156
rect 2080 1122 2120 1156
rect 2154 1122 2194 1156
rect 2228 1122 2268 1156
rect 2302 1122 2342 1156
rect 2376 1122 2416 1156
rect 2450 1122 2490 1156
rect 2524 1122 2564 1156
rect 2598 1122 2638 1156
rect 2672 1122 2712 1156
rect 2746 1122 2786 1156
rect 2820 1122 2860 1156
rect 2894 1122 2934 1156
rect 2968 1122 3008 1156
rect 3042 1122 3082 1156
rect 3116 1122 3156 1156
rect 3190 1122 3230 1156
rect 3264 1122 3606 1156
rect 3640 1122 3680 1156
rect 3714 1122 3754 1156
rect 3788 1122 3828 1156
rect 3862 1122 3902 1156
rect 3936 1122 3976 1156
rect 4010 1122 4050 1156
rect 4084 1122 4124 1156
rect 4158 1122 4198 1156
rect 4232 1122 4272 1156
rect 4306 1122 4346 1156
rect 4380 1122 4420 1156
rect 4454 1122 4494 1156
rect 4528 1122 4568 1156
rect 4602 1122 4642 1156
rect 4676 1122 4716 1156
rect 4750 1122 4790 1156
rect 4824 1122 4864 1156
rect 4898 1122 4938 1156
rect 4972 1122 5012 1156
rect 5046 1122 5085 1156
rect 5119 1122 5158 1156
rect 5192 1122 5199 1156
rect 5444 1122 5450 1156
rect 1850 1115 1862 1122
rect 1914 1115 5199 1122
rect 5251 1115 5263 1122
rect 5315 1115 5327 1122
rect 5379 1115 5392 1122
rect 5444 1115 5457 1122
rect 5509 1115 5522 1167
rect 5574 1115 5587 1167
rect 5639 1156 7511 1167
rect 5639 1122 5669 1156
rect 5703 1122 5742 1156
rect 5776 1122 5815 1156
rect 5849 1122 5888 1156
rect 5922 1122 5961 1156
rect 5995 1122 6034 1156
rect 6068 1122 6107 1156
rect 6141 1122 6180 1156
rect 6214 1122 6253 1156
rect 6287 1122 6326 1156
rect 6360 1122 6399 1156
rect 6433 1122 6472 1156
rect 6506 1122 6848 1156
rect 6882 1122 6921 1156
rect 6955 1122 6994 1156
rect 7028 1122 7067 1156
rect 7101 1122 7140 1156
rect 7174 1122 7213 1156
rect 7247 1122 7286 1156
rect 7320 1122 7359 1156
rect 7393 1122 7432 1156
rect 7466 1122 7505 1156
rect 5639 1115 7511 1122
rect 7563 1115 7576 1167
rect 7628 1115 7641 1167
rect 7693 1115 7706 1167
rect 7758 1115 7770 1167
rect 7822 1156 7834 1167
rect 7886 1156 7898 1167
rect 7950 1156 7962 1167
rect 8014 1156 8026 1167
rect 8078 1156 8090 1167
rect 7831 1122 7834 1156
rect 8014 1122 8016 1156
rect 8078 1122 8089 1156
rect 7822 1115 7834 1122
rect 7886 1115 7898 1122
rect 7950 1115 7962 1122
rect 8014 1115 8026 1122
rect 8078 1115 8090 1122
rect 8142 1115 8154 1167
rect 8206 1115 8218 1167
rect 8270 1115 8282 1167
rect 8334 1156 8346 1167
rect 8398 1156 11440 1167
rect 11492 1156 11504 1167
rect 8342 1122 8346 1156
rect 8416 1122 8456 1156
rect 8490 1122 8530 1156
rect 8564 1122 8604 1156
rect 8638 1122 8678 1156
rect 8712 1122 8752 1156
rect 8786 1122 8826 1156
rect 8860 1122 8900 1156
rect 8934 1122 8974 1156
rect 9008 1122 9048 1156
rect 9082 1122 9122 1156
rect 9156 1122 9196 1156
rect 9230 1122 9270 1156
rect 9304 1122 9344 1156
rect 9378 1122 9418 1156
rect 9452 1122 9492 1156
rect 9526 1122 9566 1156
rect 9600 1122 9640 1156
rect 9674 1122 9714 1156
rect 9748 1122 10090 1156
rect 10124 1122 10164 1156
rect 10198 1122 10238 1156
rect 10272 1122 10312 1156
rect 10346 1122 10386 1156
rect 10420 1122 10460 1156
rect 10494 1122 10534 1156
rect 10568 1122 10608 1156
rect 10642 1122 10682 1156
rect 10716 1122 10756 1156
rect 10790 1122 10830 1156
rect 10864 1122 10904 1156
rect 10938 1122 10978 1156
rect 11012 1122 11052 1156
rect 11086 1122 11126 1156
rect 11160 1122 11200 1156
rect 11234 1122 11274 1156
rect 11308 1122 11348 1156
rect 11382 1122 11422 1156
rect 11492 1122 11496 1156
rect 8334 1115 8346 1122
rect 8398 1115 11440 1122
rect 11492 1115 11504 1122
rect 11556 1115 11568 1167
rect 11620 1115 11632 1167
rect 11684 1115 11696 1167
rect 11748 1156 11760 1167
rect 11812 1156 11824 1167
rect 11876 1156 11888 1167
rect 11940 1156 11952 1167
rect 12004 1156 12016 1167
rect 11749 1122 11760 1156
rect 11822 1122 11824 1156
rect 12004 1122 12007 1156
rect 11748 1115 11760 1122
rect 11812 1115 11824 1122
rect 11876 1115 11888 1122
rect 11940 1115 11952 1122
rect 12004 1115 12016 1122
rect 12068 1115 12080 1167
rect 12132 1115 12145 1167
rect 12197 1115 12210 1167
rect 12262 1115 12275 1167
rect 12327 1156 13995 1167
rect 12333 1122 12372 1156
rect 12406 1122 12445 1156
rect 12479 1122 12518 1156
rect 12552 1122 12591 1156
rect 12625 1122 12664 1156
rect 12698 1122 12737 1156
rect 12771 1122 12810 1156
rect 12844 1122 12883 1156
rect 12917 1122 12956 1156
rect 12990 1122 13332 1156
rect 13366 1122 13405 1156
rect 13439 1122 13478 1156
rect 13512 1122 13551 1156
rect 13585 1122 13624 1156
rect 13658 1122 13697 1156
rect 13731 1122 13770 1156
rect 13804 1122 13843 1156
rect 13877 1122 13916 1156
rect 13950 1122 13989 1156
rect 12327 1115 13995 1122
rect 14047 1115 14060 1167
rect 14112 1115 14125 1167
rect 14177 1115 14190 1167
rect 14242 1115 14254 1167
rect 14306 1156 14318 1167
rect 14370 1156 14382 1167
rect 14434 1156 14446 1167
rect 14498 1156 14510 1167
rect 14562 1156 14574 1167
rect 14315 1122 14318 1156
rect 14498 1122 14500 1156
rect 14562 1122 14573 1156
rect 14306 1115 14318 1122
rect 14370 1115 14382 1122
rect 14434 1115 14446 1122
rect 14498 1115 14510 1122
rect 14562 1115 14574 1122
rect 14626 1115 14638 1167
rect 14690 1115 14702 1167
rect 14754 1115 14766 1167
rect 14818 1156 14830 1167
rect 14882 1156 17924 1167
rect 17976 1156 17988 1167
rect 14826 1122 14830 1156
rect 14900 1122 14940 1156
rect 14974 1122 15014 1156
rect 15048 1122 15088 1156
rect 15122 1122 15162 1156
rect 15196 1122 15236 1156
rect 15270 1122 15310 1156
rect 15344 1122 15384 1156
rect 15418 1122 15458 1156
rect 15492 1122 15532 1156
rect 15566 1122 15606 1156
rect 15640 1122 15680 1156
rect 15714 1122 15754 1156
rect 15788 1122 15828 1156
rect 15862 1122 15902 1156
rect 15936 1122 15976 1156
rect 16010 1122 16050 1156
rect 16084 1122 16124 1156
rect 16158 1122 16198 1156
rect 16232 1122 16574 1156
rect 16608 1122 16648 1156
rect 16682 1122 16722 1156
rect 16756 1122 16796 1156
rect 16830 1122 16870 1156
rect 16904 1122 16944 1156
rect 16978 1122 17018 1156
rect 17052 1122 17092 1156
rect 17126 1122 17166 1156
rect 17200 1122 17240 1156
rect 17274 1122 17314 1156
rect 17348 1122 17388 1156
rect 17422 1122 17462 1156
rect 17496 1122 17536 1156
rect 17570 1122 17610 1156
rect 17644 1122 17684 1156
rect 17718 1122 17758 1156
rect 17792 1122 17832 1156
rect 17866 1122 17906 1156
rect 17976 1122 17980 1156
rect 14818 1115 14830 1122
rect 14882 1115 17924 1122
rect 17976 1115 17988 1122
rect 18040 1115 18052 1167
rect 18104 1115 18116 1167
rect 18168 1115 18180 1167
rect 18232 1156 18244 1167
rect 18296 1156 18308 1167
rect 18360 1156 18372 1167
rect 18424 1156 18436 1167
rect 18488 1156 18500 1167
rect 18233 1122 18244 1156
rect 18306 1122 18308 1156
rect 18488 1122 18491 1156
rect 18232 1115 18244 1122
rect 18296 1115 18308 1122
rect 18360 1115 18372 1122
rect 18424 1115 18436 1122
rect 18488 1115 18500 1122
rect 18552 1115 18564 1167
rect 18616 1115 18629 1167
rect 18681 1115 18694 1167
rect 18746 1115 18759 1167
rect 18811 1156 19574 1167
rect 18817 1122 18856 1156
rect 18890 1122 18929 1156
rect 18963 1122 19002 1156
rect 19036 1122 19075 1156
rect 19109 1122 19148 1156
rect 19182 1122 19221 1156
rect 19255 1122 19294 1156
rect 19328 1122 19367 1156
rect 19401 1122 19440 1156
rect 19474 1122 19574 1156
rect 18811 1115 19574 1122
rect 264 1099 19574 1115
rect 264 1047 1027 1099
rect 1079 1047 1092 1099
rect 1144 1047 1157 1099
rect 1209 1047 1222 1099
rect 1274 1047 1286 1099
rect 1338 1047 1350 1099
rect 1402 1047 1414 1099
rect 1466 1047 1478 1099
rect 1530 1047 1542 1099
rect 1594 1047 1606 1099
rect 1658 1047 1670 1099
rect 1722 1047 1734 1099
rect 1786 1047 1798 1099
rect 1850 1047 1862 1099
rect 1914 1047 5199 1099
rect 5251 1047 5263 1099
rect 5315 1047 5327 1099
rect 5379 1047 5392 1099
rect 5444 1047 5457 1099
rect 5509 1047 5522 1099
rect 5574 1047 5587 1099
rect 5639 1047 7511 1099
rect 7563 1047 7576 1099
rect 7628 1047 7641 1099
rect 7693 1047 7706 1099
rect 7758 1047 7770 1099
rect 7822 1047 7834 1099
rect 7886 1047 7898 1099
rect 7950 1047 7962 1099
rect 8014 1047 8026 1099
rect 8078 1047 8090 1099
rect 8142 1047 8154 1099
rect 8206 1047 8218 1099
rect 8270 1047 8282 1099
rect 8334 1047 8346 1099
rect 8398 1047 11440 1099
rect 11492 1047 11504 1099
rect 11556 1047 11568 1099
rect 11620 1047 11632 1099
rect 11684 1047 11696 1099
rect 11748 1047 11760 1099
rect 11812 1047 11824 1099
rect 11876 1047 11888 1099
rect 11940 1047 11952 1099
rect 12004 1047 12016 1099
rect 12068 1047 12080 1099
rect 12132 1047 12145 1099
rect 12197 1047 12210 1099
rect 12262 1047 12275 1099
rect 12327 1047 13995 1099
rect 14047 1047 14060 1099
rect 14112 1047 14125 1099
rect 14177 1047 14190 1099
rect 14242 1047 14254 1099
rect 14306 1047 14318 1099
rect 14370 1047 14382 1099
rect 14434 1047 14446 1099
rect 14498 1047 14510 1099
rect 14562 1047 14574 1099
rect 14626 1047 14638 1099
rect 14690 1047 14702 1099
rect 14754 1047 14766 1099
rect 14818 1047 14830 1099
rect 14882 1047 17924 1099
rect 17976 1047 17988 1099
rect 18040 1047 18052 1099
rect 18104 1047 18116 1099
rect 18168 1047 18180 1099
rect 18232 1047 18244 1099
rect 18296 1047 18308 1099
rect 18360 1047 18372 1099
rect 18424 1047 18436 1099
rect 18488 1047 18500 1099
rect 18552 1047 18564 1099
rect 18616 1047 18629 1099
rect 18681 1047 18694 1099
rect 18746 1047 18759 1099
rect 18811 1047 19574 1099
rect 264 1031 19574 1047
rect 19759 1203 19811 1211
rect 19759 1139 19811 1151
rect -52 961 82 1001
rect -52 927 -46 961
rect -12 927 42 961
rect 76 927 82 961
rect 176 1020 228 1026
rect 264 1022 1027 1031
tri 264 1014 272 1022 ne
rect 272 1014 1027 1022
tri 272 975 311 1014 ne
rect 311 979 1027 1014
rect 1079 979 1092 1031
rect 1144 979 1157 1031
rect 1209 979 1222 1031
rect 1274 979 1286 1031
rect 1338 979 1350 1031
rect 1402 979 1414 1031
rect 1466 979 1478 1031
rect 1530 979 1542 1031
rect 1594 979 1606 1031
rect 1658 979 1670 1031
rect 1722 979 1734 1031
rect 1786 979 1798 1031
rect 1850 979 1862 1031
rect 1914 1022 5199 1031
rect 1914 1014 3356 1022
tri 3356 1014 3364 1022 nw
tri 3506 1014 3514 1022 ne
rect 3514 1014 5199 1022
rect 1914 979 3317 1014
rect 311 975 3317 979
tri 3317 975 3356 1014 nw
tri 3514 975 3553 1014 ne
rect 3553 979 5199 1014
rect 5251 979 5263 1031
rect 5315 979 5327 1031
rect 5379 979 5392 1031
rect 5444 979 5457 1031
rect 5509 979 5522 1031
rect 5574 979 5587 1031
rect 5639 1022 7511 1031
rect 5639 1014 6598 1022
tri 6598 1014 6606 1022 nw
tri 6748 1014 6756 1022 ne
rect 6756 1014 7511 1022
rect 5639 979 6559 1014
rect 3553 975 6559 979
tri 6559 975 6598 1014 nw
tri 6756 975 6795 1014 ne
rect 6795 979 7511 1014
rect 7563 979 7576 1031
rect 7628 979 7641 1031
rect 7693 979 7706 1031
rect 7758 979 7770 1031
rect 7822 979 7834 1031
rect 7886 979 7898 1031
rect 7950 979 7962 1031
rect 8014 979 8026 1031
rect 8078 979 8090 1031
rect 8142 979 8154 1031
rect 8206 979 8218 1031
rect 8270 979 8282 1031
rect 8334 979 8346 1031
rect 8398 1022 11440 1031
rect 8398 1014 9840 1022
tri 9840 1014 9848 1022 nw
tri 9990 1014 9998 1022 ne
rect 9998 1014 11440 1022
rect 8398 979 9801 1014
rect 6795 975 9801 979
tri 9801 975 9840 1014 nw
tri 9998 975 10037 1014 ne
rect 10037 979 11440 1014
rect 11492 979 11504 1031
rect 11556 979 11568 1031
rect 11620 979 11632 1031
rect 11684 979 11696 1031
rect 11748 979 11760 1031
rect 11812 979 11824 1031
rect 11876 979 11888 1031
rect 11940 979 11952 1031
rect 12004 979 12016 1031
rect 12068 979 12080 1031
rect 12132 979 12145 1031
rect 12197 979 12210 1031
rect 12262 979 12275 1031
rect 12327 1022 13995 1031
rect 12327 1014 13082 1022
tri 13082 1014 13090 1022 nw
tri 13232 1014 13240 1022 ne
rect 13240 1014 13995 1022
rect 12327 979 13043 1014
rect 10037 975 13043 979
tri 13043 975 13082 1014 nw
tri 13240 975 13279 1014 ne
rect 13279 979 13995 1014
rect 14047 979 14060 1031
rect 14112 979 14125 1031
rect 14177 979 14190 1031
rect 14242 979 14254 1031
rect 14306 979 14318 1031
rect 14370 979 14382 1031
rect 14434 979 14446 1031
rect 14498 979 14510 1031
rect 14562 979 14574 1031
rect 14626 979 14638 1031
rect 14690 979 14702 1031
rect 14754 979 14766 1031
rect 14818 979 14830 1031
rect 14882 1022 17924 1031
rect 14882 1014 16324 1022
tri 16324 1014 16332 1022 nw
tri 16474 1014 16482 1022 ne
rect 16482 1014 17924 1022
rect 14882 979 16285 1014
rect 13279 975 16285 979
tri 16285 975 16324 1014 nw
tri 16482 975 16521 1014 ne
rect 16521 979 17924 1014
rect 17976 979 17988 1031
rect 18040 979 18052 1031
rect 18104 979 18116 1031
rect 18168 979 18180 1031
rect 18232 979 18244 1031
rect 18296 979 18308 1031
rect 18360 979 18372 1031
rect 18424 979 18436 1031
rect 18488 979 18500 1031
rect 18552 979 18564 1031
rect 18616 979 18629 1031
rect 18681 979 18694 1031
rect 18746 979 18759 1031
rect 18811 1022 19574 1031
rect 18811 1014 19566 1022
tri 19566 1014 19574 1022 nw
rect 19610 1027 19662 1033
rect 18811 979 19527 1014
rect 16521 975 19527 979
tri 19527 975 19566 1014 nw
rect 19662 975 19706 994
rect 176 956 228 968
rect -52 887 82 927
rect 156 938 176 944
rect 19610 963 19706 975
rect 228 938 16332 944
rect 156 904 168 938
rect 228 904 240 938
rect 274 904 3386 938
rect 3420 904 3458 938
rect 3492 904 6628 938
rect 6662 904 6700 938
rect 6734 904 9870 938
rect 9904 904 9942 938
rect 9976 904 13136 938
rect 13170 904 13208 938
rect 13242 904 16332 938
rect 156 898 16332 904
rect 16474 938 19610 944
rect 19662 938 19706 963
rect 16474 904 19588 938
rect 19622 904 19660 911
rect 19694 904 19706 938
rect 16474 898 19706 904
rect -630 870 -306 876
rect -578 818 -306 870
rect -630 806 -306 818
rect -578 754 -306 806
rect -630 748 -306 754
rect -52 853 -46 887
rect -12 853 42 887
rect 76 853 82 887
tri 19638 875 19661 898 ne
rect -52 813 82 853
tri 277 829 311 863 se
rect 311 829 3317 863
tri 3317 829 3351 863 sw
tri 3519 829 3553 863 se
rect 3553 861 6559 863
rect 3553 829 3913 861
rect -52 779 -46 813
rect -12 779 42 813
rect 76 779 82 813
rect -52 739 82 779
rect -222 727 -170 735
rect -222 663 -170 675
rect -222 605 -170 611
rect -52 705 -46 739
rect -12 705 42 739
rect 76 705 82 739
rect -52 665 82 705
tri 264 816 277 829 se
rect 277 816 3351 829
tri 3351 816 3364 829 sw
tri 3506 816 3519 829 se
rect 3519 816 3913 829
rect 3965 816 3977 861
rect 264 782 364 816
rect 398 782 437 816
rect 471 782 510 816
rect 544 782 583 816
rect 617 782 656 816
rect 690 782 729 816
rect 763 782 802 816
rect 836 782 875 816
rect 909 782 948 816
rect 982 782 1021 816
rect 1055 782 1094 816
rect 1128 782 1167 816
rect 1201 782 1240 816
rect 1274 782 1313 816
rect 1347 782 1386 816
rect 1420 782 1459 816
rect 1493 782 1532 816
rect 1566 782 1605 816
rect 1639 782 1678 816
rect 1712 782 1751 816
rect 1785 782 1824 816
rect 1858 782 1898 816
rect 1932 782 1972 816
rect 2006 782 2046 816
rect 2080 782 2120 816
rect 2154 782 2194 816
rect 2228 782 2268 816
rect 2302 782 2342 816
rect 2376 782 2416 816
rect 2450 782 2490 816
rect 2524 782 2564 816
rect 2598 782 2638 816
rect 2672 782 2712 816
rect 2746 782 2786 816
rect 2820 782 2860 816
rect 2894 782 2934 816
rect 2968 782 3008 816
rect 3042 782 3082 816
rect 3116 782 3156 816
rect 3190 782 3230 816
rect 3264 782 3606 816
rect 3640 782 3680 816
rect 3714 782 3754 816
rect 3788 782 3828 816
rect 3862 782 3902 816
rect 3965 809 3976 816
rect 4029 809 4041 861
rect 4093 809 4105 861
rect 4157 816 4169 861
rect 4221 816 4233 861
rect 4285 816 4297 861
rect 4349 816 4361 861
rect 4413 816 4425 861
rect 4158 809 4169 816
rect 4232 809 4233 816
rect 4413 809 4420 816
rect 4477 809 4489 861
rect 4541 809 4553 861
rect 4605 809 4617 861
rect 4669 816 4681 861
rect 4733 816 4746 861
rect 4798 829 6559 861
tri 6559 829 6593 863 sw
tri 6761 829 6795 863 se
rect 6795 861 9801 863
rect 6795 829 8556 861
rect 4798 816 6593 829
tri 6593 816 6606 829 sw
tri 6748 816 6761 829 se
rect 6761 816 8556 829
rect 8608 816 8621 861
rect 8673 816 8685 861
rect 4676 809 4681 816
rect 3936 789 3976 809
rect 4010 789 4050 809
rect 4084 789 4124 809
rect 4158 789 4198 809
rect 4232 789 4272 809
rect 4306 789 4346 809
rect 4380 789 4420 809
rect 4454 789 4494 809
rect 4528 789 4568 809
rect 4602 789 4642 809
rect 4676 789 4716 809
rect 4750 789 4790 809
rect 3965 782 3976 789
rect 264 744 3913 782
rect 3965 744 3977 782
rect 264 710 364 744
rect 398 710 437 744
rect 471 710 510 744
rect 544 710 583 744
rect 617 710 656 744
rect 690 710 729 744
rect 763 710 802 744
rect 836 710 875 744
rect 909 710 948 744
rect 982 710 1021 744
rect 1055 710 1094 744
rect 1128 710 1167 744
rect 1201 710 1240 744
rect 1274 710 1313 744
rect 1347 710 1386 744
rect 1420 710 1459 744
rect 1493 710 1532 744
rect 1566 710 1605 744
rect 1639 710 1678 744
rect 1712 710 1751 744
rect 1785 710 1824 744
rect 1858 710 1898 744
rect 1932 710 1972 744
rect 2006 710 2046 744
rect 2080 710 2120 744
rect 2154 710 2194 744
rect 2228 710 2268 744
rect 2302 710 2342 744
rect 2376 710 2416 744
rect 2450 710 2490 744
rect 2524 710 2564 744
rect 2598 710 2638 744
rect 2672 710 2712 744
rect 2746 710 2786 744
rect 2820 710 2860 744
rect 2894 710 2934 744
rect 2968 710 3008 744
rect 3042 710 3082 744
rect 3116 710 3156 744
rect 3190 710 3230 744
rect 3264 710 3606 744
rect 3640 710 3680 744
rect 3714 710 3754 744
rect 3788 710 3828 744
rect 3862 710 3902 744
rect 3965 737 3976 744
rect 4029 737 4041 789
rect 4093 737 4105 789
rect 4158 782 4169 789
rect 4232 782 4233 789
rect 4413 782 4420 789
rect 4157 744 4169 782
rect 4221 744 4233 782
rect 4285 744 4297 782
rect 4349 744 4361 782
rect 4413 744 4425 782
rect 4158 737 4169 744
rect 4232 737 4233 744
rect 4413 737 4420 744
rect 4477 737 4489 789
rect 4541 737 4553 789
rect 4605 737 4617 789
rect 4676 782 4681 789
rect 4824 782 4864 816
rect 4898 782 4938 816
rect 4972 782 5012 816
rect 5046 782 5085 816
rect 5119 782 5158 816
rect 5192 782 5231 816
rect 5265 782 5304 816
rect 5338 782 5377 816
rect 5411 782 5450 816
rect 5484 782 5523 816
rect 5557 782 5596 816
rect 5630 782 5669 816
rect 5703 782 5742 816
rect 5776 782 5815 816
rect 5849 782 5888 816
rect 5922 782 5961 816
rect 5995 782 6034 816
rect 6068 782 6107 816
rect 6141 782 6180 816
rect 6214 782 6253 816
rect 6287 782 6326 816
rect 6360 782 6399 816
rect 6433 782 6472 816
rect 6506 782 6848 816
rect 6882 782 6921 816
rect 6955 782 6994 816
rect 7028 782 7067 816
rect 7101 782 7140 816
rect 7174 782 7213 816
rect 7247 782 7286 816
rect 7320 782 7359 816
rect 7393 782 7432 816
rect 7466 782 7505 816
rect 7539 782 7578 816
rect 7612 782 7651 816
rect 7685 782 7724 816
rect 7758 782 7797 816
rect 7831 782 7870 816
rect 7904 782 7943 816
rect 7977 782 8016 816
rect 8050 782 8089 816
rect 8123 782 8162 816
rect 8196 782 8235 816
rect 8269 782 8308 816
rect 8342 782 8382 816
rect 8416 782 8456 816
rect 8490 782 8530 816
rect 8673 809 8678 816
rect 8737 809 8749 861
rect 8801 809 8813 861
rect 8865 809 8877 861
rect 8929 816 8941 861
rect 8993 816 9005 861
rect 9057 816 9069 861
rect 9121 816 9133 861
rect 9185 816 9197 861
rect 8934 809 8941 816
rect 9121 809 9122 816
rect 9185 809 9196 816
rect 9249 809 9261 861
rect 9313 809 9325 861
rect 9377 816 9389 861
rect 9441 829 9801 861
tri 9801 829 9835 863 sw
tri 10003 829 10037 863 se
rect 10037 861 13043 863
rect 10037 829 10397 861
rect 9441 816 9835 829
tri 9835 816 9848 829 sw
tri 9990 816 10003 829 se
rect 10003 816 10397 829
rect 10449 816 10461 861
rect 9378 809 9389 816
rect 8564 789 8604 809
rect 8638 789 8678 809
rect 8712 789 8752 809
rect 8786 789 8826 809
rect 8860 789 8900 809
rect 8934 789 8974 809
rect 9008 789 9048 809
rect 9082 789 9122 809
rect 9156 789 9196 809
rect 9230 789 9270 809
rect 9304 789 9344 809
rect 9378 789 9418 809
rect 8673 782 8678 789
rect 4669 744 4681 782
rect 4733 744 4746 782
rect 4798 744 8556 782
rect 8608 744 8621 782
rect 8673 744 8685 782
rect 4676 737 4681 744
rect 3936 717 3976 737
rect 4010 717 4050 737
rect 4084 717 4124 737
rect 4158 717 4198 737
rect 4232 717 4272 737
rect 4306 717 4346 737
rect 4380 717 4420 737
rect 4454 717 4494 737
rect 4528 717 4568 737
rect 4602 717 4642 737
rect 4676 717 4716 737
rect 4750 717 4790 737
rect 3965 710 3976 717
tri 264 683 291 710 ne
rect 291 683 3337 710
tri 3337 683 3364 710 nw
tri 3506 683 3533 710 ne
rect 3533 683 3913 710
rect -52 631 -46 665
rect -12 631 42 665
rect 76 631 82 665
tri 291 663 311 683 ne
rect 311 663 3317 683
tri 3317 663 3337 683 nw
tri 3533 663 3553 683 ne
rect 3553 665 3913 683
rect 3965 665 3977 710
rect 4029 665 4041 717
rect 4093 665 4105 717
rect 4158 710 4169 717
rect 4232 710 4233 717
rect 4413 710 4420 717
rect 4157 665 4169 710
rect 4221 665 4233 710
rect 4285 665 4297 710
rect 4349 665 4361 710
rect 4413 665 4425 710
rect 4477 665 4489 717
rect 4541 665 4553 717
rect 4605 665 4617 717
rect 4676 710 4681 717
rect 4824 710 4864 744
rect 4898 710 4938 744
rect 4972 710 5012 744
rect 5046 710 5085 744
rect 5119 710 5158 744
rect 5192 710 5231 744
rect 5265 710 5304 744
rect 5338 710 5377 744
rect 5411 710 5450 744
rect 5484 710 5523 744
rect 5557 710 5596 744
rect 5630 710 5669 744
rect 5703 710 5742 744
rect 5776 710 5815 744
rect 5849 710 5888 744
rect 5922 710 5961 744
rect 5995 710 6034 744
rect 6068 710 6107 744
rect 6141 710 6180 744
rect 6214 710 6253 744
rect 6287 710 6326 744
rect 6360 710 6399 744
rect 6433 710 6472 744
rect 6506 710 6848 744
rect 6882 710 6921 744
rect 6955 710 6994 744
rect 7028 710 7067 744
rect 7101 710 7140 744
rect 7174 710 7213 744
rect 7247 710 7286 744
rect 7320 710 7359 744
rect 7393 710 7432 744
rect 7466 710 7505 744
rect 7539 710 7578 744
rect 7612 710 7651 744
rect 7685 710 7724 744
rect 7758 710 7797 744
rect 7831 710 7870 744
rect 7904 710 7943 744
rect 7977 710 8016 744
rect 8050 710 8089 744
rect 8123 710 8162 744
rect 8196 710 8235 744
rect 8269 710 8308 744
rect 8342 710 8382 744
rect 8416 710 8456 744
rect 8490 710 8530 744
rect 8673 737 8678 744
rect 8737 737 8749 789
rect 8801 737 8813 789
rect 8865 737 8877 789
rect 8934 782 8941 789
rect 9121 782 9122 789
rect 9185 782 9196 789
rect 8929 744 8941 782
rect 8993 744 9005 782
rect 9057 744 9069 782
rect 9121 744 9133 782
rect 9185 744 9197 782
rect 8934 737 8941 744
rect 9121 737 9122 744
rect 9185 737 9196 744
rect 9249 737 9261 789
rect 9313 737 9325 789
rect 9378 782 9389 789
rect 9452 782 9492 816
rect 9526 782 9566 816
rect 9600 782 9640 816
rect 9674 782 9714 816
rect 9748 782 10090 816
rect 10124 782 10164 816
rect 10198 782 10238 816
rect 10272 782 10312 816
rect 10346 782 10386 816
rect 10449 809 10460 816
rect 10513 809 10525 861
rect 10577 809 10589 861
rect 10641 816 10653 861
rect 10705 816 10717 861
rect 10769 816 10781 861
rect 10833 816 10845 861
rect 10897 816 10909 861
rect 10642 809 10653 816
rect 10716 809 10717 816
rect 10897 809 10904 816
rect 10961 809 10973 861
rect 11025 809 11037 861
rect 11089 809 11101 861
rect 11153 816 11165 861
rect 11217 816 11230 861
rect 11282 829 13043 861
tri 13043 829 13077 863 sw
tri 13245 829 13279 863 se
rect 13279 861 16285 863
rect 13279 829 15040 861
rect 11282 816 13077 829
tri 13077 816 13090 829 sw
tri 13232 816 13245 829 se
rect 13245 816 15040 829
rect 15092 816 15105 861
rect 15157 816 15169 861
rect 11160 809 11165 816
rect 10420 789 10460 809
rect 10494 789 10534 809
rect 10568 789 10608 809
rect 10642 789 10682 809
rect 10716 789 10756 809
rect 10790 789 10830 809
rect 10864 789 10904 809
rect 10938 789 10978 809
rect 11012 789 11052 809
rect 11086 789 11126 809
rect 11160 789 11200 809
rect 11234 789 11274 809
rect 10449 782 10460 789
rect 9377 744 9389 782
rect 9441 744 10397 782
rect 10449 744 10461 782
rect 9378 737 9389 744
rect 8564 717 8604 737
rect 8638 717 8678 737
rect 8712 717 8752 737
rect 8786 717 8826 737
rect 8860 717 8900 737
rect 8934 717 8974 737
rect 9008 717 9048 737
rect 9082 717 9122 737
rect 9156 717 9196 737
rect 9230 717 9270 737
rect 9304 717 9344 737
rect 9378 717 9418 737
rect 8673 710 8678 717
rect 4669 665 4681 710
rect 4733 665 4746 710
rect 4798 683 6579 710
tri 6579 683 6606 710 nw
tri 6748 683 6775 710 ne
rect 6775 683 8556 710
rect 4798 665 6559 683
rect 3553 663 6559 665
tri 6559 663 6579 683 nw
tri 6775 663 6795 683 ne
rect 6795 665 8556 683
rect 8608 665 8621 710
rect 8673 665 8685 710
rect 8737 665 8749 717
rect 8801 665 8813 717
rect 8865 665 8877 717
rect 8934 710 8941 717
rect 9121 710 9122 717
rect 9185 710 9196 717
rect 8929 665 8941 710
rect 8993 665 9005 710
rect 9057 665 9069 710
rect 9121 665 9133 710
rect 9185 665 9197 710
rect 9249 665 9261 717
rect 9313 665 9325 717
rect 9378 710 9389 717
rect 9452 710 9492 744
rect 9526 710 9566 744
rect 9600 710 9640 744
rect 9674 710 9714 744
rect 9748 710 10090 744
rect 10124 710 10164 744
rect 10198 710 10238 744
rect 10272 710 10312 744
rect 10346 710 10386 744
rect 10449 737 10460 744
rect 10513 737 10525 789
rect 10577 737 10589 789
rect 10642 782 10653 789
rect 10716 782 10717 789
rect 10897 782 10904 789
rect 10641 744 10653 782
rect 10705 744 10717 782
rect 10769 744 10781 782
rect 10833 744 10845 782
rect 10897 744 10909 782
rect 10642 737 10653 744
rect 10716 737 10717 744
rect 10897 737 10904 744
rect 10961 737 10973 789
rect 11025 737 11037 789
rect 11089 737 11101 789
rect 11160 782 11165 789
rect 11308 782 11348 816
rect 11382 782 11422 816
rect 11456 782 11496 816
rect 11530 782 11569 816
rect 11603 782 11642 816
rect 11676 782 11715 816
rect 11749 782 11788 816
rect 11822 782 11861 816
rect 11895 782 11934 816
rect 11968 782 12007 816
rect 12041 782 12080 816
rect 12114 782 12153 816
rect 12187 782 12226 816
rect 12260 782 12299 816
rect 12333 782 12372 816
rect 12406 782 12445 816
rect 12479 782 12518 816
rect 12552 782 12591 816
rect 12625 782 12664 816
rect 12698 782 12737 816
rect 12771 782 12810 816
rect 12844 782 12883 816
rect 12917 782 12956 816
rect 12990 782 13332 816
rect 13366 782 13405 816
rect 13439 782 13478 816
rect 13512 782 13551 816
rect 13585 782 13624 816
rect 13658 782 13697 816
rect 13731 782 13770 816
rect 13804 782 13843 816
rect 13877 782 13916 816
rect 13950 782 13989 816
rect 14023 782 14062 816
rect 14096 782 14135 816
rect 14169 782 14208 816
rect 14242 782 14281 816
rect 14315 782 14354 816
rect 14388 782 14427 816
rect 14461 782 14500 816
rect 14534 782 14573 816
rect 14607 782 14646 816
rect 14680 782 14719 816
rect 14753 782 14792 816
rect 14826 782 14866 816
rect 14900 782 14940 816
rect 14974 782 15014 816
rect 15157 809 15162 816
rect 15221 809 15233 861
rect 15285 809 15297 861
rect 15349 809 15361 861
rect 15413 816 15425 861
rect 15477 816 15489 861
rect 15541 816 15553 861
rect 15605 816 15617 861
rect 15669 816 15681 861
rect 15418 809 15425 816
rect 15605 809 15606 816
rect 15669 809 15680 816
rect 15733 809 15745 861
rect 15797 809 15809 861
rect 15861 816 15873 861
rect 15925 829 16285 861
tri 16285 829 16319 863 sw
tri 16487 829 16521 863 se
rect 16521 861 19527 863
rect 16521 829 16881 861
rect 15925 816 16319 829
tri 16319 816 16332 829 sw
tri 16474 816 16487 829 se
rect 16487 816 16881 829
rect 16933 816 16945 861
rect 15862 809 15873 816
rect 15048 789 15088 809
rect 15122 789 15162 809
rect 15196 789 15236 809
rect 15270 789 15310 809
rect 15344 789 15384 809
rect 15418 789 15458 809
rect 15492 789 15532 809
rect 15566 789 15606 809
rect 15640 789 15680 809
rect 15714 789 15754 809
rect 15788 789 15828 809
rect 15862 789 15902 809
rect 15157 782 15162 789
rect 11153 744 11165 782
rect 11217 744 11230 782
rect 11282 744 15040 782
rect 15092 744 15105 782
rect 15157 744 15169 782
rect 11160 737 11165 744
rect 10420 717 10460 737
rect 10494 717 10534 737
rect 10568 717 10608 737
rect 10642 717 10682 737
rect 10716 717 10756 737
rect 10790 717 10830 737
rect 10864 717 10904 737
rect 10938 717 10978 737
rect 11012 717 11052 737
rect 11086 717 11126 737
rect 11160 717 11200 737
rect 11234 717 11274 737
rect 10449 710 10460 717
rect 9377 665 9389 710
rect 9441 683 9821 710
tri 9821 683 9848 710 nw
tri 9990 683 10017 710 ne
rect 10017 683 10397 710
rect 9441 665 9801 683
rect 6795 663 9801 665
tri 9801 663 9821 683 nw
tri 10017 663 10037 683 ne
rect 10037 665 10397 683
rect 10449 665 10461 710
rect 10513 665 10525 717
rect 10577 665 10589 717
rect 10642 710 10653 717
rect 10716 710 10717 717
rect 10897 710 10904 717
rect 10641 665 10653 710
rect 10705 665 10717 710
rect 10769 665 10781 710
rect 10833 665 10845 710
rect 10897 665 10909 710
rect 10961 665 10973 717
rect 11025 665 11037 717
rect 11089 665 11101 717
rect 11160 710 11165 717
rect 11308 710 11348 744
rect 11382 710 11422 744
rect 11456 710 11496 744
rect 11530 710 11569 744
rect 11603 710 11642 744
rect 11676 710 11715 744
rect 11749 710 11788 744
rect 11822 710 11861 744
rect 11895 710 11934 744
rect 11968 710 12007 744
rect 12041 710 12080 744
rect 12114 710 12153 744
rect 12187 710 12226 744
rect 12260 710 12299 744
rect 12333 710 12372 744
rect 12406 710 12445 744
rect 12479 710 12518 744
rect 12552 710 12591 744
rect 12625 710 12664 744
rect 12698 710 12737 744
rect 12771 710 12810 744
rect 12844 710 12883 744
rect 12917 710 12956 744
rect 12990 710 13332 744
rect 13366 710 13405 744
rect 13439 710 13478 744
rect 13512 710 13551 744
rect 13585 710 13624 744
rect 13658 710 13697 744
rect 13731 710 13770 744
rect 13804 710 13843 744
rect 13877 710 13916 744
rect 13950 710 13989 744
rect 14023 710 14062 744
rect 14096 710 14135 744
rect 14169 710 14208 744
rect 14242 710 14281 744
rect 14315 710 14354 744
rect 14388 710 14427 744
rect 14461 710 14500 744
rect 14534 710 14573 744
rect 14607 710 14646 744
rect 14680 710 14719 744
rect 14753 710 14792 744
rect 14826 710 14866 744
rect 14900 710 14940 744
rect 14974 710 15014 744
rect 15157 737 15162 744
rect 15221 737 15233 789
rect 15285 737 15297 789
rect 15349 737 15361 789
rect 15418 782 15425 789
rect 15605 782 15606 789
rect 15669 782 15680 789
rect 15413 744 15425 782
rect 15477 744 15489 782
rect 15541 744 15553 782
rect 15605 744 15617 782
rect 15669 744 15681 782
rect 15418 737 15425 744
rect 15605 737 15606 744
rect 15669 737 15680 744
rect 15733 737 15745 789
rect 15797 737 15809 789
rect 15862 782 15873 789
rect 15936 782 15976 816
rect 16010 782 16050 816
rect 16084 782 16124 816
rect 16158 782 16198 816
rect 16232 782 16574 816
rect 16608 782 16648 816
rect 16682 782 16722 816
rect 16756 782 16796 816
rect 16830 782 16870 816
rect 16933 809 16944 816
rect 16997 809 17009 861
rect 17061 809 17073 861
rect 17125 816 17137 861
rect 17189 816 17201 861
rect 17253 816 17265 861
rect 17317 816 17329 861
rect 17381 816 17393 861
rect 17126 809 17137 816
rect 17200 809 17201 816
rect 17381 809 17388 816
rect 17445 809 17457 861
rect 17509 809 17521 861
rect 17573 809 17585 861
rect 17637 816 17649 861
rect 17701 816 17714 861
rect 17766 829 19527 861
tri 19527 829 19561 863 sw
rect 17766 816 19561 829
tri 19561 816 19574 829 sw
rect 17644 809 17649 816
rect 16904 789 16944 809
rect 16978 789 17018 809
rect 17052 789 17092 809
rect 17126 789 17166 809
rect 17200 789 17240 809
rect 17274 789 17314 809
rect 17348 789 17388 809
rect 17422 789 17462 809
rect 17496 789 17536 809
rect 17570 789 17610 809
rect 17644 789 17684 809
rect 17718 789 17758 809
rect 16933 782 16944 789
rect 15861 744 15873 782
rect 15925 744 16881 782
rect 16933 744 16945 782
rect 15862 737 15873 744
rect 15048 717 15088 737
rect 15122 717 15162 737
rect 15196 717 15236 737
rect 15270 717 15310 737
rect 15344 717 15384 737
rect 15418 717 15458 737
rect 15492 717 15532 737
rect 15566 717 15606 737
rect 15640 717 15680 737
rect 15714 717 15754 737
rect 15788 717 15828 737
rect 15862 717 15902 737
rect 15157 710 15162 717
rect 11153 665 11165 710
rect 11217 665 11230 710
rect 11282 683 13063 710
tri 13063 683 13090 710 nw
tri 13232 683 13259 710 ne
rect 13259 683 15040 710
rect 11282 665 13043 683
rect 10037 663 13043 665
tri 13043 663 13063 683 nw
tri 13259 663 13279 683 ne
rect 13279 665 15040 683
rect 15092 665 15105 710
rect 15157 665 15169 710
rect 15221 665 15233 717
rect 15285 665 15297 717
rect 15349 665 15361 717
rect 15418 710 15425 717
rect 15605 710 15606 717
rect 15669 710 15680 717
rect 15413 665 15425 710
rect 15477 665 15489 710
rect 15541 665 15553 710
rect 15605 665 15617 710
rect 15669 665 15681 710
rect 15733 665 15745 717
rect 15797 665 15809 717
rect 15862 710 15873 717
rect 15936 710 15976 744
rect 16010 710 16050 744
rect 16084 710 16124 744
rect 16158 710 16198 744
rect 16232 710 16574 744
rect 16608 710 16648 744
rect 16682 710 16722 744
rect 16756 710 16796 744
rect 16830 710 16870 744
rect 16933 737 16944 744
rect 16997 737 17009 789
rect 17061 737 17073 789
rect 17126 782 17137 789
rect 17200 782 17201 789
rect 17381 782 17388 789
rect 17125 744 17137 782
rect 17189 744 17201 782
rect 17253 744 17265 782
rect 17317 744 17329 782
rect 17381 744 17393 782
rect 17126 737 17137 744
rect 17200 737 17201 744
rect 17381 737 17388 744
rect 17445 737 17457 789
rect 17509 737 17521 789
rect 17573 737 17585 789
rect 17644 782 17649 789
rect 17792 782 17832 816
rect 17866 782 17906 816
rect 17940 782 17980 816
rect 18014 782 18053 816
rect 18087 782 18126 816
rect 18160 782 18199 816
rect 18233 782 18272 816
rect 18306 782 18345 816
rect 18379 782 18418 816
rect 18452 782 18491 816
rect 18525 782 18564 816
rect 18598 782 18637 816
rect 18671 782 18710 816
rect 18744 782 18783 816
rect 18817 782 18856 816
rect 18890 782 18929 816
rect 18963 782 19002 816
rect 19036 782 19075 816
rect 19109 782 19148 816
rect 19182 782 19221 816
rect 19255 782 19294 816
rect 19328 782 19367 816
rect 19401 782 19440 816
rect 19474 782 19574 816
rect 17637 744 17649 782
rect 17701 744 17714 782
rect 17766 744 19574 782
rect 17644 737 17649 744
rect 16904 717 16944 737
rect 16978 717 17018 737
rect 17052 717 17092 737
rect 17126 717 17166 737
rect 17200 717 17240 737
rect 17274 717 17314 737
rect 17348 717 17388 737
rect 17422 717 17462 737
rect 17496 717 17536 737
rect 17570 717 17610 737
rect 17644 717 17684 737
rect 17718 717 17758 737
rect 16933 710 16944 717
rect 15861 665 15873 710
rect 15925 683 16305 710
tri 16305 683 16332 710 nw
tri 16474 683 16501 710 ne
rect 16501 683 16881 710
rect 15925 665 16285 683
rect 13279 663 16285 665
tri 16285 663 16305 683 nw
tri 16501 663 16521 683 ne
rect 16521 665 16881 683
rect 16933 665 16945 710
rect 16997 665 17009 717
rect 17061 665 17073 717
rect 17126 710 17137 717
rect 17200 710 17201 717
rect 17381 710 17388 717
rect 17125 665 17137 710
rect 17189 665 17201 710
rect 17253 665 17265 710
rect 17317 665 17329 710
rect 17381 665 17393 710
rect 17445 665 17457 717
rect 17509 665 17521 717
rect 17573 665 17585 717
rect 17644 710 17649 717
rect 17792 710 17832 744
rect 17866 710 17906 744
rect 17940 710 17980 744
rect 18014 710 18053 744
rect 18087 710 18126 744
rect 18160 710 18199 744
rect 18233 710 18272 744
rect 18306 710 18345 744
rect 18379 710 18418 744
rect 18452 710 18491 744
rect 18525 710 18564 744
rect 18598 710 18637 744
rect 18671 710 18710 744
rect 18744 710 18783 744
rect 18817 710 18856 744
rect 18890 710 18929 744
rect 18963 710 19002 744
rect 19036 710 19075 744
rect 19109 710 19148 744
rect 19182 710 19221 744
rect 19255 710 19294 744
rect 19328 710 19367 744
rect 19401 710 19440 744
rect 19474 710 19574 744
rect 17637 665 17649 710
rect 17701 665 17714 710
rect 17766 683 19547 710
tri 19547 683 19574 710 nw
rect 17766 665 19527 683
rect 16521 663 19527 665
tri 19527 663 19547 683 nw
rect -52 591 82 631
tri 19642 628 19661 647 se
rect 19661 628 19706 898
rect -52 557 -46 591
rect -12 557 42 591
rect 76 557 82 591
rect 132 622 19706 628
rect 132 588 144 622
rect 178 588 216 622
rect 250 588 3386 622
rect 3420 588 3458 622
rect 3492 588 6628 622
rect 6662 588 6700 622
rect 6734 588 9870 622
rect 9904 588 9942 622
rect 9976 588 13112 622
rect 13146 588 13184 622
rect 13218 588 16354 622
rect 16388 588 16426 622
rect 16460 588 19564 622
rect 19598 615 19636 622
rect 19598 588 19610 615
rect 19670 588 19706 622
rect 132 582 19610 588
rect -52 517 82 557
rect 19662 563 19706 588
rect 19610 551 19706 563
tri 297 537 311 551 se
rect 311 547 3317 551
rect 311 537 1027 547
rect -52 483 -46 517
rect -12 483 42 517
rect 76 483 82 517
rect -52 443 82 483
rect -52 409 -46 443
rect -12 409 42 443
rect 76 409 82 443
rect -52 369 82 409
rect -52 335 -46 369
rect -12 335 42 369
rect 76 335 82 369
rect -52 295 82 335
rect -52 261 -46 295
rect -12 261 42 295
rect 76 261 82 295
rect -52 221 82 261
rect -52 187 -46 221
rect -12 187 42 221
rect 76 187 82 221
tri 264 504 297 537 se
rect 297 504 1027 537
rect 264 495 1027 504
rect 1079 495 1092 547
rect 1144 495 1157 547
rect 1209 495 1222 547
rect 1274 495 1286 547
rect 1338 495 1350 547
rect 1402 495 1414 547
rect 1466 495 1478 547
rect 1530 495 1542 547
rect 1594 495 1606 547
rect 1658 495 1670 547
rect 1722 495 1734 547
rect 1786 495 1798 547
rect 1850 495 1862 547
rect 1914 537 3317 547
tri 3317 537 3331 551 sw
tri 3539 537 3553 551 se
rect 3553 547 6559 551
rect 3553 537 5199 547
rect 1914 504 3331 537
tri 3331 504 3364 537 sw
tri 3506 504 3539 537 se
rect 3539 504 5199 537
rect 1914 495 5199 504
rect 5251 495 5263 547
rect 5315 495 5327 547
rect 5379 495 5392 547
rect 5444 495 5457 547
rect 5509 495 5522 547
rect 5574 495 5587 547
rect 5639 537 6559 547
tri 6559 537 6573 551 sw
tri 6781 537 6795 551 se
rect 6795 547 9801 551
rect 6795 537 7511 547
rect 5639 504 6573 537
tri 6573 504 6606 537 sw
tri 6748 504 6781 537 se
rect 6781 504 7511 537
rect 5639 495 7511 504
rect 7563 495 7576 547
rect 7628 495 7641 547
rect 7693 495 7706 547
rect 7758 495 7770 547
rect 7822 495 7834 547
rect 7886 495 7898 547
rect 7950 495 7962 547
rect 8014 495 8026 547
rect 8078 495 8090 547
rect 8142 495 8154 547
rect 8206 495 8218 547
rect 8270 495 8282 547
rect 8334 495 8346 547
rect 8398 537 9801 547
tri 9801 537 9815 551 sw
tri 10023 537 10037 551 se
rect 10037 547 13043 551
rect 10037 537 11440 547
rect 8398 504 9815 537
tri 9815 504 9848 537 sw
tri 9990 504 10023 537 se
rect 10023 504 11440 537
rect 8398 495 11440 504
rect 11492 495 11504 547
rect 11556 495 11568 547
rect 11620 495 11632 547
rect 11684 495 11696 547
rect 11748 495 11760 547
rect 11812 495 11824 547
rect 11876 495 11888 547
rect 11940 495 11952 547
rect 12004 495 12016 547
rect 12068 495 12080 547
rect 12132 495 12145 547
rect 12197 495 12210 547
rect 12262 495 12275 547
rect 12327 537 13043 547
tri 13043 537 13057 551 sw
tri 13265 537 13279 551 se
rect 13279 547 16285 551
rect 13279 537 13995 547
rect 12327 504 13057 537
tri 13057 504 13090 537 sw
tri 13232 504 13265 537 se
rect 13265 504 13995 537
rect 12327 495 13995 504
rect 14047 495 14060 547
rect 14112 495 14125 547
rect 14177 495 14190 547
rect 14242 495 14254 547
rect 14306 495 14318 547
rect 14370 495 14382 547
rect 14434 495 14446 547
rect 14498 495 14510 547
rect 14562 495 14574 547
rect 14626 495 14638 547
rect 14690 495 14702 547
rect 14754 495 14766 547
rect 14818 495 14830 547
rect 14882 537 16285 547
tri 16285 537 16299 551 sw
tri 16507 537 16521 551 se
rect 16521 547 19527 551
rect 16521 537 17924 547
rect 14882 504 16299 537
tri 16299 504 16332 537 sw
tri 16474 504 16507 537 se
rect 16507 504 17924 537
rect 14882 495 17924 504
rect 17976 495 17988 547
rect 18040 495 18052 547
rect 18104 495 18116 547
rect 18168 495 18180 547
rect 18232 495 18244 547
rect 18296 495 18308 547
rect 18360 495 18372 547
rect 18424 495 18436 547
rect 18488 495 18500 547
rect 18552 495 18564 547
rect 18616 495 18629 547
rect 18681 495 18694 547
rect 18746 495 18759 547
rect 18811 537 19527 547
tri 19527 537 19541 551 sw
rect 18811 504 19541 537
tri 19541 504 19574 537 sw
rect 18811 495 19574 504
rect 264 479 19574 495
rect 19662 499 19706 551
rect 19610 493 19706 499
rect 264 427 1027 479
rect 1079 427 1092 479
rect 1144 427 1157 479
rect 1209 427 1222 479
rect 1274 427 1286 479
rect 1338 427 1350 479
rect 1402 427 1414 479
rect 1466 427 1478 479
rect 1530 427 1542 479
rect 1594 427 1606 479
rect 1658 427 1670 479
rect 1722 427 1734 479
rect 1786 427 1798 479
rect 1850 427 1862 479
rect 1914 427 5199 479
rect 5251 427 5263 479
rect 5315 427 5327 479
rect 5379 427 5392 479
rect 5444 427 5457 479
rect 5509 427 5522 479
rect 5574 427 5587 479
rect 5639 427 7511 479
rect 7563 427 7576 479
rect 7628 427 7641 479
rect 7693 427 7706 479
rect 7758 427 7770 479
rect 7822 427 7834 479
rect 7886 427 7898 479
rect 7950 427 7962 479
rect 8014 427 8026 479
rect 8078 427 8090 479
rect 8142 427 8154 479
rect 8206 427 8218 479
rect 8270 427 8282 479
rect 8334 427 8346 479
rect 8398 427 11440 479
rect 11492 427 11504 479
rect 11556 427 11568 479
rect 11620 427 11632 479
rect 11684 427 11696 479
rect 11748 427 11760 479
rect 11812 427 11824 479
rect 11876 427 11888 479
rect 11940 427 11952 479
rect 12004 427 12016 479
rect 12068 427 12080 479
rect 12132 427 12145 479
rect 12197 427 12210 479
rect 12262 427 12275 479
rect 12327 427 13995 479
rect 14047 427 14060 479
rect 14112 427 14125 479
rect 14177 427 14190 479
rect 14242 427 14254 479
rect 14306 427 14318 479
rect 14370 427 14382 479
rect 14434 427 14446 479
rect 14498 427 14510 479
rect 14562 427 14574 479
rect 14626 427 14638 479
rect 14690 427 14702 479
rect 14754 427 14766 479
rect 14818 427 14830 479
rect 14882 427 17924 479
rect 17976 427 17988 479
rect 18040 427 18052 479
rect 18104 427 18116 479
rect 18168 427 18180 479
rect 18232 427 18244 479
rect 18296 427 18308 479
rect 18360 427 18372 479
rect 18424 427 18436 479
rect 18488 427 18500 479
rect 18552 427 18564 479
rect 18616 427 18629 479
rect 18681 427 18694 479
rect 18746 427 18759 479
rect 18811 427 19574 479
tri 19629 465 19657 493 ne
rect 19657 465 19706 493
tri 19657 463 19659 465 ne
rect 19659 463 19706 465
rect 264 411 19574 427
rect 264 404 1027 411
rect 264 370 364 404
rect 398 370 437 404
rect 471 370 510 404
rect 544 370 583 404
rect 617 370 656 404
rect 690 370 729 404
rect 763 370 802 404
rect 836 370 875 404
rect 909 370 948 404
rect 982 370 1021 404
rect 264 359 1027 370
rect 1079 359 1092 411
rect 1144 359 1157 411
rect 1209 359 1222 411
rect 1274 359 1286 411
rect 1338 404 1350 411
rect 1402 404 1414 411
rect 1466 404 1478 411
rect 1530 404 1542 411
rect 1594 404 1606 411
rect 1347 370 1350 404
rect 1530 370 1532 404
rect 1594 370 1605 404
rect 1338 359 1350 370
rect 1402 359 1414 370
rect 1466 359 1478 370
rect 1530 359 1542 370
rect 1594 359 1606 370
rect 1658 359 1670 411
rect 1722 359 1734 411
rect 1786 359 1798 411
rect 1850 404 1862 411
rect 1914 404 5199 411
rect 5251 404 5263 411
rect 5315 404 5327 411
rect 5379 404 5392 411
rect 5444 404 5457 411
rect 1858 370 1862 404
rect 1932 370 1972 404
rect 2006 370 2046 404
rect 2080 370 2120 404
rect 2154 370 2194 404
rect 2228 370 2268 404
rect 2302 370 2342 404
rect 2376 370 2416 404
rect 2450 370 2490 404
rect 2524 370 2564 404
rect 2598 370 2638 404
rect 2672 370 2712 404
rect 2746 370 2786 404
rect 2820 370 2860 404
rect 2894 370 2934 404
rect 2968 370 3008 404
rect 3042 370 3082 404
rect 3116 370 3156 404
rect 3190 370 3230 404
rect 3264 370 3606 404
rect 3640 370 3680 404
rect 3714 370 3754 404
rect 3788 370 3828 404
rect 3862 370 3902 404
rect 3936 370 3976 404
rect 4010 370 4050 404
rect 4084 370 4124 404
rect 4158 370 4198 404
rect 4232 370 4272 404
rect 4306 370 4346 404
rect 4380 370 4420 404
rect 4454 370 4494 404
rect 4528 370 4568 404
rect 4602 370 4642 404
rect 4676 370 4716 404
rect 4750 370 4790 404
rect 4824 370 4864 404
rect 4898 370 4938 404
rect 4972 370 5012 404
rect 5046 370 5085 404
rect 5119 370 5158 404
rect 5192 370 5199 404
rect 5444 370 5450 404
rect 1850 359 1862 370
rect 1914 359 5199 370
rect 5251 359 5263 370
rect 5315 359 5327 370
rect 5379 359 5392 370
rect 5444 359 5457 370
rect 5509 359 5522 411
rect 5574 359 5587 411
rect 5639 404 7511 411
rect 5639 370 5669 404
rect 5703 370 5742 404
rect 5776 370 5815 404
rect 5849 370 5888 404
rect 5922 370 5961 404
rect 5995 370 6034 404
rect 6068 370 6107 404
rect 6141 370 6180 404
rect 6214 370 6253 404
rect 6287 370 6326 404
rect 6360 370 6399 404
rect 6433 370 6472 404
rect 6506 370 6848 404
rect 6882 370 6921 404
rect 6955 370 6994 404
rect 7028 370 7067 404
rect 7101 370 7140 404
rect 7174 370 7213 404
rect 7247 370 7286 404
rect 7320 370 7359 404
rect 7393 370 7432 404
rect 7466 370 7505 404
rect 5639 359 7511 370
rect 7563 359 7576 411
rect 7628 359 7641 411
rect 7693 359 7706 411
rect 7758 359 7770 411
rect 7822 404 7834 411
rect 7886 404 7898 411
rect 7950 404 7962 411
rect 8014 404 8026 411
rect 8078 404 8090 411
rect 7831 370 7834 404
rect 8014 370 8016 404
rect 8078 370 8089 404
rect 7822 359 7834 370
rect 7886 359 7898 370
rect 7950 359 7962 370
rect 8014 359 8026 370
rect 8078 359 8090 370
rect 8142 359 8154 411
rect 8206 359 8218 411
rect 8270 359 8282 411
rect 8334 404 8346 411
rect 8398 404 11440 411
rect 11492 404 11504 411
rect 8342 370 8346 404
rect 8416 370 8456 404
rect 8490 370 8530 404
rect 8564 370 8604 404
rect 8638 370 8678 404
rect 8712 370 8752 404
rect 8786 370 8826 404
rect 8860 370 8900 404
rect 8934 370 8974 404
rect 9008 370 9048 404
rect 9082 370 9122 404
rect 9156 370 9196 404
rect 9230 370 9270 404
rect 9304 370 9344 404
rect 9378 370 9418 404
rect 9452 370 9492 404
rect 9526 370 9566 404
rect 9600 370 9640 404
rect 9674 370 9714 404
rect 9748 370 10090 404
rect 10124 370 10164 404
rect 10198 370 10238 404
rect 10272 370 10312 404
rect 10346 370 10386 404
rect 10420 370 10460 404
rect 10494 370 10534 404
rect 10568 370 10608 404
rect 10642 370 10682 404
rect 10716 370 10756 404
rect 10790 370 10830 404
rect 10864 370 10904 404
rect 10938 370 10978 404
rect 11012 370 11052 404
rect 11086 370 11126 404
rect 11160 370 11200 404
rect 11234 370 11274 404
rect 11308 370 11348 404
rect 11382 370 11422 404
rect 11492 370 11496 404
rect 8334 359 8346 370
rect 8398 359 11440 370
rect 11492 359 11504 370
rect 11556 359 11568 411
rect 11620 359 11632 411
rect 11684 359 11696 411
rect 11748 404 11760 411
rect 11812 404 11824 411
rect 11876 404 11888 411
rect 11940 404 11952 411
rect 12004 404 12016 411
rect 11749 370 11760 404
rect 11822 370 11824 404
rect 12004 370 12007 404
rect 11748 359 11760 370
rect 11812 359 11824 370
rect 11876 359 11888 370
rect 11940 359 11952 370
rect 12004 359 12016 370
rect 12068 359 12080 411
rect 12132 359 12145 411
rect 12197 359 12210 411
rect 12262 359 12275 411
rect 12327 404 13995 411
rect 12333 370 12372 404
rect 12406 370 12445 404
rect 12479 370 12518 404
rect 12552 370 12591 404
rect 12625 370 12664 404
rect 12698 370 12737 404
rect 12771 370 12810 404
rect 12844 370 12883 404
rect 12917 370 12956 404
rect 12990 370 13332 404
rect 13366 370 13405 404
rect 13439 370 13478 404
rect 13512 370 13551 404
rect 13585 370 13624 404
rect 13658 370 13697 404
rect 13731 370 13770 404
rect 13804 370 13843 404
rect 13877 370 13916 404
rect 13950 370 13989 404
rect 12327 359 13995 370
rect 14047 359 14060 411
rect 14112 359 14125 411
rect 14177 359 14190 411
rect 14242 359 14254 411
rect 14306 404 14318 411
rect 14370 404 14382 411
rect 14434 404 14446 411
rect 14498 404 14510 411
rect 14562 404 14574 411
rect 14315 370 14318 404
rect 14498 370 14500 404
rect 14562 370 14573 404
rect 14306 359 14318 370
rect 14370 359 14382 370
rect 14434 359 14446 370
rect 14498 359 14510 370
rect 14562 359 14574 370
rect 14626 359 14638 411
rect 14690 359 14702 411
rect 14754 359 14766 411
rect 14818 404 14830 411
rect 14882 404 17924 411
rect 17976 404 17988 411
rect 14826 370 14830 404
rect 14900 370 14940 404
rect 14974 370 15014 404
rect 15048 370 15088 404
rect 15122 370 15162 404
rect 15196 370 15236 404
rect 15270 370 15310 404
rect 15344 370 15384 404
rect 15418 370 15458 404
rect 15492 370 15532 404
rect 15566 370 15606 404
rect 15640 370 15680 404
rect 15714 370 15754 404
rect 15788 370 15828 404
rect 15862 370 15902 404
rect 15936 370 15976 404
rect 16010 370 16050 404
rect 16084 370 16124 404
rect 16158 370 16198 404
rect 16232 370 16574 404
rect 16608 370 16648 404
rect 16682 370 16722 404
rect 16756 370 16796 404
rect 16830 370 16870 404
rect 16904 370 16944 404
rect 16978 370 17018 404
rect 17052 370 17092 404
rect 17126 370 17166 404
rect 17200 370 17240 404
rect 17274 370 17314 404
rect 17348 370 17388 404
rect 17422 370 17462 404
rect 17496 370 17536 404
rect 17570 370 17610 404
rect 17644 370 17684 404
rect 17718 370 17758 404
rect 17792 370 17832 404
rect 17866 370 17906 404
rect 17976 370 17980 404
rect 14818 359 14830 370
rect 14882 359 17924 370
rect 17976 359 17988 370
rect 18040 359 18052 411
rect 18104 359 18116 411
rect 18168 359 18180 411
rect 18232 404 18244 411
rect 18296 404 18308 411
rect 18360 404 18372 411
rect 18424 404 18436 411
rect 18488 404 18500 411
rect 18233 370 18244 404
rect 18306 370 18308 404
rect 18488 370 18491 404
rect 18232 359 18244 370
rect 18296 359 18308 370
rect 18360 359 18372 370
rect 18424 359 18436 370
rect 18488 359 18500 370
rect 18552 359 18564 411
rect 18616 359 18629 411
rect 18681 359 18694 411
rect 18746 359 18759 411
rect 18811 404 19574 411
rect 18817 370 18856 404
rect 18890 370 18929 404
rect 18963 370 19002 404
rect 19036 370 19075 404
rect 19109 370 19148 404
rect 19182 370 19221 404
rect 19255 370 19294 404
rect 19328 370 19367 404
rect 19401 370 19440 404
rect 19474 370 19574 404
rect 18811 359 19574 370
rect 264 343 19574 359
rect 264 332 1027 343
rect 264 298 364 332
rect 398 298 437 332
rect 471 298 510 332
rect 544 298 583 332
rect 617 298 656 332
rect 690 298 729 332
rect 763 298 802 332
rect 836 298 875 332
rect 909 298 948 332
rect 982 298 1021 332
rect 264 291 1027 298
rect 1079 291 1092 343
rect 1144 291 1157 343
rect 1209 291 1222 343
rect 1274 291 1286 343
rect 1338 332 1350 343
rect 1402 332 1414 343
rect 1466 332 1478 343
rect 1530 332 1542 343
rect 1594 332 1606 343
rect 1347 298 1350 332
rect 1530 298 1532 332
rect 1594 298 1605 332
rect 1338 291 1350 298
rect 1402 291 1414 298
rect 1466 291 1478 298
rect 1530 291 1542 298
rect 1594 291 1606 298
rect 1658 291 1670 343
rect 1722 291 1734 343
rect 1786 291 1798 343
rect 1850 332 1862 343
rect 1914 332 5199 343
rect 5251 332 5263 343
rect 5315 332 5327 343
rect 5379 332 5392 343
rect 5444 332 5457 343
rect 1858 298 1862 332
rect 1932 298 1972 332
rect 2006 298 2046 332
rect 2080 298 2120 332
rect 2154 298 2194 332
rect 2228 298 2268 332
rect 2302 298 2342 332
rect 2376 298 2416 332
rect 2450 298 2490 332
rect 2524 298 2564 332
rect 2598 298 2638 332
rect 2672 298 2712 332
rect 2746 298 2786 332
rect 2820 298 2860 332
rect 2894 298 2934 332
rect 2968 298 3008 332
rect 3042 298 3082 332
rect 3116 298 3156 332
rect 3190 298 3230 332
rect 3264 298 3606 332
rect 3640 298 3680 332
rect 3714 298 3754 332
rect 3788 298 3828 332
rect 3862 298 3902 332
rect 3936 298 3976 332
rect 4010 298 4050 332
rect 4084 298 4124 332
rect 4158 298 4198 332
rect 4232 298 4272 332
rect 4306 298 4346 332
rect 4380 298 4420 332
rect 4454 298 4494 332
rect 4528 298 4568 332
rect 4602 298 4642 332
rect 4676 298 4716 332
rect 4750 298 4790 332
rect 4824 298 4864 332
rect 4898 298 4938 332
rect 4972 298 5012 332
rect 5046 298 5085 332
rect 5119 298 5158 332
rect 5192 298 5199 332
rect 5444 298 5450 332
rect 1850 291 1862 298
rect 1914 291 5199 298
rect 5251 291 5263 298
rect 5315 291 5327 298
rect 5379 291 5392 298
rect 5444 291 5457 298
rect 5509 291 5522 343
rect 5574 291 5587 343
rect 5639 332 7511 343
rect 5639 298 5669 332
rect 5703 298 5742 332
rect 5776 298 5815 332
rect 5849 298 5888 332
rect 5922 298 5961 332
rect 5995 298 6034 332
rect 6068 298 6107 332
rect 6141 298 6180 332
rect 6214 298 6253 332
rect 6287 298 6326 332
rect 6360 298 6399 332
rect 6433 298 6472 332
rect 6506 298 6848 332
rect 6882 298 6921 332
rect 6955 298 6994 332
rect 7028 298 7067 332
rect 7101 298 7140 332
rect 7174 298 7213 332
rect 7247 298 7286 332
rect 7320 298 7359 332
rect 7393 298 7432 332
rect 7466 298 7505 332
rect 5639 291 7511 298
rect 7563 291 7576 343
rect 7628 291 7641 343
rect 7693 291 7706 343
rect 7758 291 7770 343
rect 7822 332 7834 343
rect 7886 332 7898 343
rect 7950 332 7962 343
rect 8014 332 8026 343
rect 8078 332 8090 343
rect 7831 298 7834 332
rect 8014 298 8016 332
rect 8078 298 8089 332
rect 7822 291 7834 298
rect 7886 291 7898 298
rect 7950 291 7962 298
rect 8014 291 8026 298
rect 8078 291 8090 298
rect 8142 291 8154 343
rect 8206 291 8218 343
rect 8270 291 8282 343
rect 8334 332 8346 343
rect 8398 332 11440 343
rect 11492 332 11504 343
rect 8342 298 8346 332
rect 8416 298 8456 332
rect 8490 298 8530 332
rect 8564 298 8604 332
rect 8638 298 8678 332
rect 8712 298 8752 332
rect 8786 298 8826 332
rect 8860 298 8900 332
rect 8934 298 8974 332
rect 9008 298 9048 332
rect 9082 298 9122 332
rect 9156 298 9196 332
rect 9230 298 9270 332
rect 9304 298 9344 332
rect 9378 298 9418 332
rect 9452 298 9492 332
rect 9526 298 9566 332
rect 9600 298 9640 332
rect 9674 298 9714 332
rect 9748 298 10090 332
rect 10124 298 10164 332
rect 10198 298 10238 332
rect 10272 298 10312 332
rect 10346 298 10386 332
rect 10420 298 10460 332
rect 10494 298 10534 332
rect 10568 298 10608 332
rect 10642 298 10682 332
rect 10716 298 10756 332
rect 10790 298 10830 332
rect 10864 298 10904 332
rect 10938 298 10978 332
rect 11012 298 11052 332
rect 11086 298 11126 332
rect 11160 298 11200 332
rect 11234 298 11274 332
rect 11308 298 11348 332
rect 11382 298 11422 332
rect 11492 298 11496 332
rect 8334 291 8346 298
rect 8398 291 11440 298
rect 11492 291 11504 298
rect 11556 291 11568 343
rect 11620 291 11632 343
rect 11684 291 11696 343
rect 11748 332 11760 343
rect 11812 332 11824 343
rect 11876 332 11888 343
rect 11940 332 11952 343
rect 12004 332 12016 343
rect 11749 298 11760 332
rect 11822 298 11824 332
rect 12004 298 12007 332
rect 11748 291 11760 298
rect 11812 291 11824 298
rect 11876 291 11888 298
rect 11940 291 11952 298
rect 12004 291 12016 298
rect 12068 291 12080 343
rect 12132 291 12145 343
rect 12197 291 12210 343
rect 12262 291 12275 343
rect 12327 332 13995 343
rect 12333 298 12372 332
rect 12406 298 12445 332
rect 12479 298 12518 332
rect 12552 298 12591 332
rect 12625 298 12664 332
rect 12698 298 12737 332
rect 12771 298 12810 332
rect 12844 298 12883 332
rect 12917 298 12956 332
rect 12990 298 13332 332
rect 13366 298 13405 332
rect 13439 298 13478 332
rect 13512 298 13551 332
rect 13585 298 13624 332
rect 13658 298 13697 332
rect 13731 298 13770 332
rect 13804 298 13843 332
rect 13877 298 13916 332
rect 13950 298 13989 332
rect 12327 291 13995 298
rect 14047 291 14060 343
rect 14112 291 14125 343
rect 14177 291 14190 343
rect 14242 291 14254 343
rect 14306 332 14318 343
rect 14370 332 14382 343
rect 14434 332 14446 343
rect 14498 332 14510 343
rect 14562 332 14574 343
rect 14315 298 14318 332
rect 14498 298 14500 332
rect 14562 298 14573 332
rect 14306 291 14318 298
rect 14370 291 14382 298
rect 14434 291 14446 298
rect 14498 291 14510 298
rect 14562 291 14574 298
rect 14626 291 14638 343
rect 14690 291 14702 343
rect 14754 291 14766 343
rect 14818 332 14830 343
rect 14882 332 17924 343
rect 17976 332 17988 343
rect 14826 298 14830 332
rect 14900 298 14940 332
rect 14974 298 15014 332
rect 15048 298 15088 332
rect 15122 298 15162 332
rect 15196 298 15236 332
rect 15270 298 15310 332
rect 15344 298 15384 332
rect 15418 298 15458 332
rect 15492 298 15532 332
rect 15566 298 15606 332
rect 15640 298 15680 332
rect 15714 298 15754 332
rect 15788 298 15828 332
rect 15862 298 15902 332
rect 15936 298 15976 332
rect 16010 298 16050 332
rect 16084 298 16124 332
rect 16158 298 16198 332
rect 16232 298 16574 332
rect 16608 298 16648 332
rect 16682 298 16722 332
rect 16756 298 16796 332
rect 16830 298 16870 332
rect 16904 298 16944 332
rect 16978 298 17018 332
rect 17052 298 17092 332
rect 17126 298 17166 332
rect 17200 298 17240 332
rect 17274 298 17314 332
rect 17348 298 17388 332
rect 17422 298 17462 332
rect 17496 298 17536 332
rect 17570 298 17610 332
rect 17644 298 17684 332
rect 17718 298 17758 332
rect 17792 298 17832 332
rect 17866 298 17906 332
rect 17976 298 17980 332
rect 14818 291 14830 298
rect 14882 291 17924 298
rect 17976 291 17988 298
rect 18040 291 18052 343
rect 18104 291 18116 343
rect 18168 291 18180 343
rect 18232 332 18244 343
rect 18296 332 18308 343
rect 18360 332 18372 343
rect 18424 332 18436 343
rect 18488 332 18500 343
rect 18233 298 18244 332
rect 18306 298 18308 332
rect 18488 298 18491 332
rect 18232 291 18244 298
rect 18296 291 18308 298
rect 18360 291 18372 298
rect 18424 291 18436 298
rect 18488 291 18500 298
rect 18552 291 18564 343
rect 18616 291 18629 343
rect 18681 291 18694 343
rect 18746 291 18759 343
rect 18811 332 19574 343
rect 18817 298 18856 332
rect 18890 298 18929 332
rect 18963 298 19002 332
rect 19036 298 19075 332
rect 19109 298 19148 332
rect 19182 298 19221 332
rect 19255 298 19294 332
rect 19328 298 19367 332
rect 19401 298 19440 332
rect 19474 298 19574 332
rect 18811 291 19574 298
rect 264 275 19574 291
rect 264 223 1027 275
rect 1079 223 1092 275
rect 1144 223 1157 275
rect 1209 223 1222 275
rect 1274 223 1286 275
rect 1338 223 1350 275
rect 1402 223 1414 275
rect 1466 223 1478 275
rect 1530 223 1542 275
rect 1594 223 1606 275
rect 1658 223 1670 275
rect 1722 223 1734 275
rect 1786 223 1798 275
rect 1850 223 1862 275
rect 1914 223 5199 275
rect 5251 223 5263 275
rect 5315 223 5327 275
rect 5379 223 5392 275
rect 5444 223 5457 275
rect 5509 223 5522 275
rect 5574 223 5587 275
rect 5639 223 7511 275
rect 7563 223 7576 275
rect 7628 223 7641 275
rect 7693 223 7706 275
rect 7758 223 7770 275
rect 7822 223 7834 275
rect 7886 223 7898 275
rect 7950 223 7962 275
rect 8014 223 8026 275
rect 8078 223 8090 275
rect 8142 223 8154 275
rect 8206 223 8218 275
rect 8270 223 8282 275
rect 8334 223 8346 275
rect 8398 223 11440 275
rect 11492 223 11504 275
rect 11556 223 11568 275
rect 11620 223 11632 275
rect 11684 223 11696 275
rect 11748 223 11760 275
rect 11812 223 11824 275
rect 11876 223 11888 275
rect 11940 223 11952 275
rect 12004 223 12016 275
rect 12068 223 12080 275
rect 12132 223 12145 275
rect 12197 223 12210 275
rect 12262 223 12275 275
rect 12327 223 13995 275
rect 14047 223 14060 275
rect 14112 223 14125 275
rect 14177 223 14190 275
rect 14242 223 14254 275
rect 14306 223 14318 275
rect 14370 223 14382 275
rect 14434 223 14446 275
rect 14498 223 14510 275
rect 14562 223 14574 275
rect 14626 223 14638 275
rect 14690 223 14702 275
rect 14754 223 14766 275
rect 14818 223 14830 275
rect 14882 223 17924 275
rect 17976 223 17988 275
rect 18040 223 18052 275
rect 18104 223 18116 275
rect 18168 223 18180 275
rect 18232 223 18244 275
rect 18296 223 18308 275
rect 18360 223 18372 275
rect 18424 223 18436 275
rect 18488 223 18500 275
rect 18552 223 18564 275
rect 18616 223 18629 275
rect 18681 223 18694 275
rect 18746 223 18759 275
rect 18811 223 19574 275
rect -138 152 -86 160
rect -138 88 -86 100
rect -138 -146 -86 36
rect -138 -210 -86 -198
rect -138 -268 -86 -262
rect -52 147 82 187
rect -52 113 -46 147
rect -12 113 42 147
rect 76 113 82 147
rect 176 203 228 209
rect 264 207 19574 223
tri 19637 215 19659 237 se
rect 19659 215 19706 237
tri 19631 209 19637 215 se
rect 19637 209 19706 215
rect 264 198 1027 207
tri 264 177 285 198 ne
rect 285 177 1027 198
tri 285 151 311 177 ne
rect 311 155 1027 177
rect 1079 155 1092 207
rect 1144 155 1157 207
rect 1209 155 1222 207
rect 1274 155 1286 207
rect 1338 155 1350 207
rect 1402 155 1414 207
rect 1466 155 1478 207
rect 1530 155 1542 207
rect 1594 155 1606 207
rect 1658 155 1670 207
rect 1722 155 1734 207
rect 1786 155 1798 207
rect 1850 155 1862 207
rect 1914 198 5199 207
rect 1914 177 3343 198
tri 3343 177 3364 198 nw
tri 3506 177 3527 198 ne
rect 3527 177 5199 198
rect 1914 155 3317 177
rect 311 151 3317 155
tri 3317 151 3343 177 nw
tri 3527 151 3553 177 ne
rect 3553 155 5199 177
rect 5251 155 5263 207
rect 5315 155 5327 207
rect 5379 155 5392 207
rect 5444 155 5457 207
rect 5509 155 5522 207
rect 5574 155 5587 207
rect 5639 198 7511 207
rect 5639 177 6585 198
tri 6585 177 6606 198 nw
tri 6748 177 6769 198 ne
rect 6769 177 7511 198
rect 5639 155 6559 177
rect 3553 151 6559 155
tri 6559 151 6585 177 nw
tri 6769 151 6795 177 ne
rect 6795 155 7511 177
rect 7563 155 7576 207
rect 7628 155 7641 207
rect 7693 155 7706 207
rect 7758 155 7770 207
rect 7822 155 7834 207
rect 7886 155 7898 207
rect 7950 155 7962 207
rect 8014 155 8026 207
rect 8078 155 8090 207
rect 8142 155 8154 207
rect 8206 155 8218 207
rect 8270 155 8282 207
rect 8334 155 8346 207
rect 8398 198 11440 207
rect 8398 177 9827 198
tri 9827 177 9848 198 nw
tri 9990 177 10011 198 ne
rect 10011 177 11440 198
rect 8398 155 9801 177
rect 6795 151 9801 155
tri 9801 151 9827 177 nw
tri 10011 151 10037 177 ne
rect 10037 155 11440 177
rect 11492 155 11504 207
rect 11556 155 11568 207
rect 11620 155 11632 207
rect 11684 155 11696 207
rect 11748 155 11760 207
rect 11812 155 11824 207
rect 11876 155 11888 207
rect 11940 155 11952 207
rect 12004 155 12016 207
rect 12068 155 12080 207
rect 12132 155 12145 207
rect 12197 155 12210 207
rect 12262 155 12275 207
rect 12327 198 13995 207
rect 12327 177 13069 198
tri 13069 177 13090 198 nw
tri 13232 177 13253 198 ne
rect 13253 177 13995 198
rect 12327 155 13043 177
rect 10037 151 13043 155
tri 13043 151 13069 177 nw
tri 13253 151 13279 177 ne
rect 13279 155 13995 177
rect 14047 155 14060 207
rect 14112 155 14125 207
rect 14177 155 14190 207
rect 14242 155 14254 207
rect 14306 155 14318 207
rect 14370 155 14382 207
rect 14434 155 14446 207
rect 14498 155 14510 207
rect 14562 155 14574 207
rect 14626 155 14638 207
rect 14690 155 14702 207
rect 14754 155 14766 207
rect 14818 155 14830 207
rect 14882 198 17924 207
rect 14882 177 16311 198
tri 16311 177 16332 198 nw
tri 16474 177 16495 198 ne
rect 16495 177 17924 198
rect 14882 155 16285 177
rect 13279 151 16285 155
tri 16285 151 16311 177 nw
tri 16495 151 16521 177 ne
rect 16521 155 17924 177
rect 17976 155 17988 207
rect 18040 155 18052 207
rect 18104 155 18116 207
rect 18168 155 18180 207
rect 18232 155 18244 207
rect 18296 155 18308 207
rect 18360 155 18372 207
rect 18424 155 18436 207
rect 18488 155 18500 207
rect 18552 155 18564 207
rect 18616 155 18629 207
rect 18681 155 18694 207
rect 18746 155 18759 207
rect 18811 198 19574 207
rect 18811 177 19553 198
tri 19553 177 19574 198 nw
rect 19610 203 19706 209
rect 18811 155 19527 177
rect 16521 151 19527 155
tri 19527 151 19553 177 nw
rect 19662 151 19706 203
rect 176 139 228 151
rect -52 73 82 113
rect 156 114 176 120
rect 19610 139 19706 151
rect 228 114 13090 120
rect 156 80 168 114
rect 228 87 240 114
rect 202 80 240 87
rect 274 80 3386 114
rect 3420 80 3458 114
rect 3492 80 9870 114
rect 9904 80 9942 114
rect 9976 80 13090 114
rect 156 74 13090 80
rect 13233 114 19610 120
rect 19662 114 19706 139
rect 13233 80 16354 114
rect 16388 80 16426 114
rect 16460 80 19588 114
rect 19622 80 19660 87
rect 19694 80 19706 114
rect 13233 74 19706 80
rect -52 39 -46 73
rect -12 39 42 73
rect 76 39 82 73
rect -52 -1 82 39
tri 305 33 311 39 se
rect 311 33 3317 39
tri 3317 33 3323 39 sw
tri 3547 33 3553 39 se
rect 3553 38 6559 39
rect 3553 33 3913 38
tri 271 -1 305 33 se
rect 305 -1 3323 33
tri 3323 -1 3357 33 sw
tri 3513 -1 3547 33 se
rect 3547 -1 3913 33
rect -52 -35 -46 -1
rect -12 -35 42 -1
rect 76 -35 82 -1
rect -52 -75 82 -35
rect -52 -109 -46 -75
rect -12 -109 42 -75
rect 76 -109 82 -75
rect -52 -149 82 -109
tri 264 -8 271 -1 se
rect 271 -8 3357 -1
tri 3357 -8 3364 -1 sw
tri 3506 -8 3513 -1 se
rect 3513 -8 3913 -1
rect 3965 -8 3978 38
rect 264 -42 364 -8
rect 398 -42 437 -8
rect 471 -42 510 -8
rect 544 -42 583 -8
rect 617 -42 656 -8
rect 690 -42 729 -8
rect 763 -42 802 -8
rect 836 -42 875 -8
rect 909 -42 948 -8
rect 982 -42 1021 -8
rect 1055 -42 1094 -8
rect 1128 -42 1167 -8
rect 1201 -42 1240 -8
rect 1274 -42 1313 -8
rect 1347 -42 1386 -8
rect 1420 -42 1459 -8
rect 1493 -42 1532 -8
rect 1566 -42 1605 -8
rect 1639 -42 1678 -8
rect 1712 -42 1751 -8
rect 1785 -42 1824 -8
rect 1858 -42 1898 -8
rect 1932 -42 1972 -8
rect 2006 -42 2046 -8
rect 2080 -42 2120 -8
rect 2154 -42 2194 -8
rect 2228 -42 2268 -8
rect 2302 -42 2342 -8
rect 2376 -42 2416 -8
rect 2450 -42 2490 -8
rect 2524 -42 2564 -8
rect 2598 -42 2638 -8
rect 2672 -42 2712 -8
rect 2746 -42 2786 -8
rect 2820 -42 2860 -8
rect 2894 -42 2934 -8
rect 2968 -42 3008 -8
rect 3042 -42 3082 -8
rect 3116 -42 3156 -8
rect 3190 -42 3230 -8
rect 3264 -42 3606 -8
rect 3640 -42 3680 -8
rect 3714 -42 3754 -8
rect 3788 -42 3828 -8
rect 3862 -42 3902 -8
rect 3965 -14 3976 -8
rect 4030 -14 4042 38
rect 4094 -14 4106 38
rect 4158 -14 4170 38
rect 4222 -8 4234 38
rect 4286 -8 4298 38
rect 4350 -8 4362 38
rect 4414 -8 4426 38
rect 4232 -14 4234 -8
rect 4414 -14 4420 -8
rect 4478 -14 4490 38
rect 4542 -14 4554 38
rect 4606 -14 4618 38
rect 4670 -8 4682 38
rect 4734 -8 4746 38
rect 4798 33 6559 38
tri 6559 33 6565 39 sw
tri 6789 33 6795 39 se
rect 6795 38 9801 39
rect 6795 33 8556 38
rect 4798 -1 6565 33
tri 6565 -1 6599 33 sw
tri 6755 -1 6789 33 se
rect 6789 -1 8556 33
rect 4798 -8 6599 -1
tri 6599 -8 6606 -1 sw
tri 6748 -8 6755 -1 se
rect 6755 -8 8556 -1
rect 8608 -8 8621 38
rect 8673 -8 8685 38
rect 4676 -14 4682 -8
rect 3936 -34 3976 -14
rect 4010 -34 4050 -14
rect 4084 -34 4124 -14
rect 4158 -34 4198 -14
rect 4232 -34 4272 -14
rect 4306 -34 4346 -14
rect 4380 -34 4420 -14
rect 4454 -34 4494 -14
rect 4528 -34 4568 -14
rect 4602 -34 4642 -14
rect 4676 -34 4716 -14
rect 4750 -34 4790 -14
rect 3965 -42 3976 -34
rect 264 -80 3913 -42
rect 3965 -80 3978 -42
rect 264 -114 364 -80
rect 398 -114 437 -80
rect 471 -114 510 -80
rect 544 -114 583 -80
rect 617 -114 656 -80
rect 690 -114 729 -80
rect 763 -114 802 -80
rect 836 -114 875 -80
rect 909 -114 948 -80
rect 982 -114 1021 -80
rect 1055 -114 1094 -80
rect 1128 -114 1167 -80
rect 1201 -114 1240 -80
rect 1274 -114 1313 -80
rect 1347 -114 1386 -80
rect 1420 -114 1459 -80
rect 1493 -114 1532 -80
rect 1566 -114 1605 -80
rect 1639 -114 1678 -80
rect 1712 -114 1751 -80
rect 1785 -114 1824 -80
rect 1858 -114 1898 -80
rect 1932 -114 1972 -80
rect 2006 -114 2046 -80
rect 2080 -114 2120 -80
rect 2154 -114 2194 -80
rect 2228 -114 2268 -80
rect 2302 -114 2342 -80
rect 2376 -114 2416 -80
rect 2450 -114 2490 -80
rect 2524 -114 2564 -80
rect 2598 -114 2638 -80
rect 2672 -114 2712 -80
rect 2746 -114 2786 -80
rect 2820 -114 2860 -80
rect 2894 -114 2934 -80
rect 2968 -114 3008 -80
rect 3042 -114 3082 -80
rect 3116 -114 3156 -80
rect 3190 -114 3230 -80
rect 3264 -114 3606 -80
rect 3640 -114 3680 -80
rect 3714 -114 3754 -80
rect 3788 -114 3828 -80
rect 3862 -114 3902 -80
rect 3965 -86 3976 -80
rect 4030 -86 4042 -34
rect 4094 -86 4106 -34
rect 4158 -86 4170 -34
rect 4232 -42 4234 -34
rect 4414 -42 4420 -34
rect 4222 -80 4234 -42
rect 4286 -80 4298 -42
rect 4350 -80 4362 -42
rect 4414 -80 4426 -42
rect 4232 -86 4234 -80
rect 4414 -86 4420 -80
rect 4478 -86 4490 -34
rect 4542 -86 4554 -34
rect 4606 -86 4618 -34
rect 4676 -42 4682 -34
rect 4824 -42 4864 -8
rect 4898 -42 4938 -8
rect 4972 -42 5012 -8
rect 5046 -42 5085 -8
rect 5119 -42 5158 -8
rect 5192 -42 5231 -8
rect 5265 -42 5304 -8
rect 5338 -42 5377 -8
rect 5411 -42 5450 -8
rect 5484 -42 5523 -8
rect 5557 -42 5596 -8
rect 5630 -42 5669 -8
rect 5703 -42 5742 -8
rect 5776 -42 5815 -8
rect 5849 -42 5888 -8
rect 5922 -42 5961 -8
rect 5995 -42 6034 -8
rect 6068 -42 6107 -8
rect 6141 -42 6180 -8
rect 6214 -42 6253 -8
rect 6287 -42 6326 -8
rect 6360 -42 6399 -8
rect 6433 -42 6472 -8
rect 6506 -42 6848 -8
rect 6882 -42 6921 -8
rect 6955 -42 6994 -8
rect 7028 -42 7067 -8
rect 7101 -42 7140 -8
rect 7174 -42 7213 -8
rect 7247 -42 7286 -8
rect 7320 -42 7359 -8
rect 7393 -42 7432 -8
rect 7466 -42 7505 -8
rect 7539 -42 7578 -8
rect 7612 -42 7651 -8
rect 7685 -42 7724 -8
rect 7758 -42 7797 -8
rect 7831 -42 7870 -8
rect 7904 -42 7943 -8
rect 7977 -42 8016 -8
rect 8050 -42 8089 -8
rect 8123 -42 8162 -8
rect 8196 -42 8235 -8
rect 8269 -42 8308 -8
rect 8342 -42 8382 -8
rect 8416 -42 8456 -8
rect 8490 -42 8530 -8
rect 8673 -14 8678 -8
rect 8737 -14 8749 38
rect 8801 -14 8813 38
rect 8865 -14 8877 38
rect 8929 -8 8941 38
rect 8993 -8 9005 38
rect 9057 -8 9069 38
rect 9121 -8 9133 38
rect 9185 -8 9197 38
rect 8934 -14 8941 -8
rect 9121 -14 9122 -8
rect 9185 -14 9196 -8
rect 9249 -14 9261 38
rect 9313 -14 9325 38
rect 9377 -8 9389 38
rect 9441 33 9801 38
tri 9801 33 9807 39 sw
tri 10031 33 10037 39 se
rect 10037 38 13043 39
rect 10037 33 10397 38
rect 9441 -1 9807 33
tri 9807 -1 9841 33 sw
tri 9997 -1 10031 33 se
rect 10031 -1 10397 33
rect 9441 -8 9841 -1
tri 9841 -8 9848 -1 sw
tri 9990 -8 9997 -1 se
rect 9997 -8 10397 -1
rect 10449 -8 10462 38
rect 9378 -14 9389 -8
rect 8564 -34 8604 -14
rect 8638 -34 8678 -14
rect 8712 -34 8752 -14
rect 8786 -34 8826 -14
rect 8860 -34 8900 -14
rect 8934 -34 8974 -14
rect 9008 -34 9048 -14
rect 9082 -34 9122 -14
rect 9156 -34 9196 -14
rect 9230 -34 9270 -14
rect 9304 -34 9344 -14
rect 9378 -34 9418 -14
rect 8673 -42 8678 -34
rect 4670 -80 4682 -42
rect 4734 -80 4746 -42
rect 4798 -80 8556 -42
rect 8608 -80 8621 -42
rect 8673 -80 8685 -42
rect 4676 -86 4682 -80
rect 3936 -106 3976 -86
rect 4010 -106 4050 -86
rect 4084 -106 4124 -86
rect 4158 -106 4198 -86
rect 4232 -106 4272 -86
rect 4306 -106 4346 -86
rect 4380 -106 4420 -86
rect 4454 -106 4494 -86
rect 4528 -106 4568 -86
rect 4602 -106 4642 -86
rect 4676 -106 4716 -86
rect 4750 -106 4790 -86
rect 3965 -114 3976 -106
tri 264 -145 295 -114 ne
rect 295 -145 3333 -114
tri 3333 -145 3364 -114 nw
tri 3506 -145 3537 -114 ne
rect 3537 -145 3913 -114
rect -52 -183 -46 -149
rect -12 -183 42 -149
rect 76 -183 82 -149
tri 295 -161 311 -145 ne
rect 311 -161 3317 -145
tri 3317 -161 3333 -145 nw
tri 3537 -161 3553 -145 ne
rect 3553 -158 3913 -145
rect 3965 -158 3978 -114
rect 4030 -158 4042 -106
rect 4094 -158 4106 -106
rect 4158 -158 4170 -106
rect 4232 -114 4234 -106
rect 4414 -114 4420 -106
rect 4222 -158 4234 -114
rect 4286 -158 4298 -114
rect 4350 -158 4362 -114
rect 4414 -158 4426 -114
rect 4478 -158 4490 -106
rect 4542 -158 4554 -106
rect 4606 -158 4618 -106
rect 4676 -114 4682 -106
rect 4824 -114 4864 -80
rect 4898 -114 4938 -80
rect 4972 -114 5012 -80
rect 5046 -114 5085 -80
rect 5119 -114 5158 -80
rect 5192 -114 5231 -80
rect 5265 -114 5304 -80
rect 5338 -114 5377 -80
rect 5411 -114 5450 -80
rect 5484 -114 5523 -80
rect 5557 -114 5596 -80
rect 5630 -114 5669 -80
rect 5703 -114 5742 -80
rect 5776 -114 5815 -80
rect 5849 -114 5888 -80
rect 5922 -114 5961 -80
rect 5995 -114 6034 -80
rect 6068 -114 6107 -80
rect 6141 -114 6180 -80
rect 6214 -114 6253 -80
rect 6287 -114 6326 -80
rect 6360 -114 6399 -80
rect 6433 -114 6472 -80
rect 6506 -114 6848 -80
rect 6882 -114 6921 -80
rect 6955 -114 6994 -80
rect 7028 -114 7067 -80
rect 7101 -114 7140 -80
rect 7174 -114 7213 -80
rect 7247 -114 7286 -80
rect 7320 -114 7359 -80
rect 7393 -114 7432 -80
rect 7466 -114 7505 -80
rect 7539 -114 7578 -80
rect 7612 -114 7651 -80
rect 7685 -114 7724 -80
rect 7758 -114 7797 -80
rect 7831 -114 7870 -80
rect 7904 -114 7943 -80
rect 7977 -114 8016 -80
rect 8050 -114 8089 -80
rect 8123 -114 8162 -80
rect 8196 -114 8235 -80
rect 8269 -114 8308 -80
rect 8342 -114 8382 -80
rect 8416 -114 8456 -80
rect 8490 -114 8530 -80
rect 8673 -86 8678 -80
rect 8737 -86 8749 -34
rect 8801 -86 8813 -34
rect 8865 -86 8877 -34
rect 8934 -42 8941 -34
rect 9121 -42 9122 -34
rect 9185 -42 9196 -34
rect 8929 -80 8941 -42
rect 8993 -80 9005 -42
rect 9057 -80 9069 -42
rect 9121 -80 9133 -42
rect 9185 -80 9197 -42
rect 8934 -86 8941 -80
rect 9121 -86 9122 -80
rect 9185 -86 9196 -80
rect 9249 -86 9261 -34
rect 9313 -86 9325 -34
rect 9378 -42 9389 -34
rect 9452 -42 9492 -8
rect 9526 -42 9566 -8
rect 9600 -42 9640 -8
rect 9674 -42 9714 -8
rect 9748 -42 10090 -8
rect 10124 -42 10164 -8
rect 10198 -42 10238 -8
rect 10272 -42 10312 -8
rect 10346 -42 10386 -8
rect 10449 -14 10460 -8
rect 10514 -14 10526 38
rect 10578 -14 10590 38
rect 10642 -14 10654 38
rect 10706 -8 10718 38
rect 10770 -8 10782 38
rect 10834 -8 10846 38
rect 10898 -8 10910 38
rect 10716 -14 10718 -8
rect 10898 -14 10904 -8
rect 10962 -14 10974 38
rect 11026 -14 11038 38
rect 11090 -14 11102 38
rect 11154 -8 11166 38
rect 11218 -8 11230 38
rect 11282 33 13043 38
tri 13043 33 13049 39 sw
tri 13273 33 13279 39 se
rect 13279 37 16285 39
rect 13279 33 15040 37
rect 11282 -1 13049 33
tri 13049 -1 13083 33 sw
tri 13239 -1 13273 33 se
rect 13273 -1 15040 33
rect 11282 -8 13083 -1
tri 13083 -8 13090 -1 sw
tri 13232 -8 13239 -1 se
rect 13239 -8 15040 -1
rect 15092 -8 15105 37
rect 15157 -8 15169 37
rect 11160 -14 11166 -8
rect 10420 -34 10460 -14
rect 10494 -34 10534 -14
rect 10568 -34 10608 -14
rect 10642 -34 10682 -14
rect 10716 -34 10756 -14
rect 10790 -34 10830 -14
rect 10864 -34 10904 -14
rect 10938 -34 10978 -14
rect 11012 -34 11052 -14
rect 11086 -34 11126 -14
rect 11160 -34 11200 -14
rect 11234 -34 11274 -14
rect 10449 -42 10460 -34
rect 9377 -80 9389 -42
rect 9441 -80 10397 -42
rect 10449 -80 10462 -42
rect 9378 -86 9389 -80
rect 8564 -106 8604 -86
rect 8638 -106 8678 -86
rect 8712 -106 8752 -86
rect 8786 -106 8826 -86
rect 8860 -106 8900 -86
rect 8934 -106 8974 -86
rect 9008 -106 9048 -86
rect 9082 -106 9122 -86
rect 9156 -106 9196 -86
rect 9230 -106 9270 -86
rect 9304 -106 9344 -86
rect 9378 -106 9418 -86
rect 8673 -114 8678 -106
rect 4670 -158 4682 -114
rect 4734 -158 4746 -114
rect 4798 -145 6575 -114
tri 6575 -145 6606 -114 nw
tri 6748 -145 6779 -114 ne
rect 6779 -145 8556 -114
rect 4798 -158 6559 -145
rect 3553 -161 6559 -158
tri 6559 -161 6575 -145 nw
tri 6779 -161 6795 -145 ne
rect 6795 -158 8556 -145
rect 8608 -158 8621 -114
rect 8673 -158 8685 -114
rect 8737 -158 8749 -106
rect 8801 -158 8813 -106
rect 8865 -158 8877 -106
rect 8934 -114 8941 -106
rect 9121 -114 9122 -106
rect 9185 -114 9196 -106
rect 8929 -158 8941 -114
rect 8993 -158 9005 -114
rect 9057 -158 9069 -114
rect 9121 -158 9133 -114
rect 9185 -158 9197 -114
rect 9249 -158 9261 -106
rect 9313 -158 9325 -106
rect 9378 -114 9389 -106
rect 9452 -114 9492 -80
rect 9526 -114 9566 -80
rect 9600 -114 9640 -80
rect 9674 -114 9714 -80
rect 9748 -114 10090 -80
rect 10124 -114 10164 -80
rect 10198 -114 10238 -80
rect 10272 -114 10312 -80
rect 10346 -114 10386 -80
rect 10449 -86 10460 -80
rect 10514 -86 10526 -34
rect 10578 -86 10590 -34
rect 10642 -86 10654 -34
rect 10716 -42 10718 -34
rect 10898 -42 10904 -34
rect 10706 -80 10718 -42
rect 10770 -80 10782 -42
rect 10834 -80 10846 -42
rect 10898 -80 10910 -42
rect 10716 -86 10718 -80
rect 10898 -86 10904 -80
rect 10962 -86 10974 -34
rect 11026 -86 11038 -34
rect 11090 -86 11102 -34
rect 11160 -42 11166 -34
rect 11308 -42 11348 -8
rect 11382 -42 11422 -8
rect 11456 -42 11496 -8
rect 11530 -42 11569 -8
rect 11603 -42 11642 -8
rect 11676 -42 11715 -8
rect 11749 -42 11788 -8
rect 11822 -42 11861 -8
rect 11895 -42 11934 -8
rect 11968 -42 12007 -8
rect 12041 -42 12080 -8
rect 12114 -42 12153 -8
rect 12187 -42 12226 -8
rect 12260 -42 12299 -8
rect 12333 -42 12372 -8
rect 12406 -42 12445 -8
rect 12479 -42 12518 -8
rect 12552 -42 12591 -8
rect 12625 -42 12664 -8
rect 12698 -42 12737 -8
rect 12771 -42 12810 -8
rect 12844 -42 12883 -8
rect 12917 -42 12956 -8
rect 12990 -42 13332 -8
rect 13366 -42 13405 -8
rect 13439 -42 13478 -8
rect 13512 -42 13551 -8
rect 13585 -42 13624 -8
rect 13658 -42 13697 -8
rect 13731 -42 13770 -8
rect 13804 -42 13843 -8
rect 13877 -42 13916 -8
rect 13950 -42 13989 -8
rect 14023 -42 14062 -8
rect 14096 -42 14135 -8
rect 14169 -42 14208 -8
rect 14242 -42 14281 -8
rect 14315 -42 14354 -8
rect 14388 -42 14427 -8
rect 14461 -42 14500 -8
rect 14534 -42 14573 -8
rect 14607 -42 14646 -8
rect 14680 -42 14719 -8
rect 14753 -42 14792 -8
rect 14826 -42 14866 -8
rect 14900 -42 14940 -8
rect 14974 -42 15014 -8
rect 15157 -15 15162 -8
rect 15221 -15 15233 37
rect 15285 -15 15297 37
rect 15349 -15 15361 37
rect 15413 -8 15425 37
rect 15477 -8 15489 37
rect 15541 -8 15553 37
rect 15605 -8 15617 37
rect 15669 -8 15681 37
rect 15418 -15 15425 -8
rect 15605 -15 15606 -8
rect 15669 -15 15680 -8
rect 15733 -15 15745 37
rect 15797 -15 15809 37
rect 15861 -8 15873 37
rect 15925 33 16285 37
tri 16285 33 16291 39 sw
tri 16515 33 16521 39 se
rect 16521 37 19527 39
rect 16521 33 16881 37
rect 15925 -1 16291 33
tri 16291 -1 16325 33 sw
tri 16481 -1 16515 33 se
rect 16515 -1 16881 33
rect 15925 -8 16325 -1
tri 16325 -8 16332 -1 sw
tri 16474 -8 16481 -1 se
rect 16481 -8 16881 -1
rect 16933 -8 16946 37
rect 15862 -15 15873 -8
rect 15048 -35 15088 -15
rect 15122 -35 15162 -15
rect 15196 -35 15236 -15
rect 15270 -35 15310 -15
rect 15344 -35 15384 -15
rect 15418 -35 15458 -15
rect 15492 -35 15532 -15
rect 15566 -35 15606 -15
rect 15640 -35 15680 -15
rect 15714 -35 15754 -15
rect 15788 -35 15828 -15
rect 15862 -35 15902 -15
rect 15157 -42 15162 -35
rect 11154 -80 11166 -42
rect 11218 -80 11230 -42
rect 11282 -80 15040 -42
rect 15092 -80 15105 -42
rect 15157 -80 15169 -42
rect 11160 -86 11166 -80
rect 10420 -106 10460 -86
rect 10494 -106 10534 -86
rect 10568 -106 10608 -86
rect 10642 -106 10682 -86
rect 10716 -106 10756 -86
rect 10790 -106 10830 -86
rect 10864 -106 10904 -86
rect 10938 -106 10978 -86
rect 11012 -106 11052 -86
rect 11086 -106 11126 -86
rect 11160 -106 11200 -86
rect 11234 -106 11274 -86
rect 10449 -114 10460 -106
rect 9377 -158 9389 -114
rect 9441 -145 9817 -114
tri 9817 -145 9848 -114 nw
tri 9990 -145 10021 -114 ne
rect 10021 -145 10397 -114
rect 9441 -158 9801 -145
rect 6795 -161 9801 -158
tri 9801 -161 9817 -145 nw
tri 10021 -161 10037 -145 ne
rect 10037 -158 10397 -145
rect 10449 -158 10462 -114
rect 10514 -158 10526 -106
rect 10578 -158 10590 -106
rect 10642 -158 10654 -106
rect 10716 -114 10718 -106
rect 10898 -114 10904 -106
rect 10706 -158 10718 -114
rect 10770 -158 10782 -114
rect 10834 -158 10846 -114
rect 10898 -158 10910 -114
rect 10962 -158 10974 -106
rect 11026 -158 11038 -106
rect 11090 -158 11102 -106
rect 11160 -114 11166 -106
rect 11308 -114 11348 -80
rect 11382 -114 11422 -80
rect 11456 -114 11496 -80
rect 11530 -114 11569 -80
rect 11603 -114 11642 -80
rect 11676 -114 11715 -80
rect 11749 -114 11788 -80
rect 11822 -114 11861 -80
rect 11895 -114 11934 -80
rect 11968 -114 12007 -80
rect 12041 -114 12080 -80
rect 12114 -114 12153 -80
rect 12187 -114 12226 -80
rect 12260 -114 12299 -80
rect 12333 -114 12372 -80
rect 12406 -114 12445 -80
rect 12479 -114 12518 -80
rect 12552 -114 12591 -80
rect 12625 -114 12664 -80
rect 12698 -114 12737 -80
rect 12771 -114 12810 -80
rect 12844 -114 12883 -80
rect 12917 -114 12956 -80
rect 12990 -114 13332 -80
rect 13366 -114 13405 -80
rect 13439 -114 13478 -80
rect 13512 -114 13551 -80
rect 13585 -114 13624 -80
rect 13658 -114 13697 -80
rect 13731 -114 13770 -80
rect 13804 -114 13843 -80
rect 13877 -114 13916 -80
rect 13950 -114 13989 -80
rect 14023 -114 14062 -80
rect 14096 -114 14135 -80
rect 14169 -114 14208 -80
rect 14242 -114 14281 -80
rect 14315 -114 14354 -80
rect 14388 -114 14427 -80
rect 14461 -114 14500 -80
rect 14534 -114 14573 -80
rect 14607 -114 14646 -80
rect 14680 -114 14719 -80
rect 14753 -114 14792 -80
rect 14826 -114 14866 -80
rect 14900 -114 14940 -80
rect 14974 -114 15014 -80
rect 15157 -87 15162 -80
rect 15221 -87 15233 -35
rect 15285 -87 15297 -35
rect 15349 -87 15361 -35
rect 15418 -42 15425 -35
rect 15605 -42 15606 -35
rect 15669 -42 15680 -35
rect 15413 -80 15425 -42
rect 15477 -80 15489 -42
rect 15541 -80 15553 -42
rect 15605 -80 15617 -42
rect 15669 -80 15681 -42
rect 15418 -87 15425 -80
rect 15605 -87 15606 -80
rect 15669 -87 15680 -80
rect 15733 -87 15745 -35
rect 15797 -87 15809 -35
rect 15862 -42 15873 -35
rect 15936 -42 15976 -8
rect 16010 -42 16050 -8
rect 16084 -42 16124 -8
rect 16158 -42 16198 -8
rect 16232 -42 16574 -8
rect 16608 -42 16648 -8
rect 16682 -42 16722 -8
rect 16756 -42 16796 -8
rect 16830 -42 16870 -8
rect 16933 -15 16944 -8
rect 16998 -15 17010 37
rect 17062 -15 17074 37
rect 17126 -15 17138 37
rect 17190 -8 17202 37
rect 17254 -8 17266 37
rect 17318 -8 17330 37
rect 17382 -8 17394 37
rect 17200 -15 17202 -8
rect 17382 -15 17388 -8
rect 17446 -15 17458 37
rect 17510 -15 17522 37
rect 17574 -15 17586 37
rect 17638 -8 17650 37
rect 17702 -8 17714 37
rect 17766 33 19527 37
tri 19527 33 19533 39 sw
rect 17766 -1 19533 33
tri 19533 -1 19567 33 sw
rect 17766 -8 19567 -1
tri 19567 -8 19574 -1 sw
rect 17644 -15 17650 -8
rect 16904 -35 16944 -15
rect 16978 -35 17018 -15
rect 17052 -35 17092 -15
rect 17126 -35 17166 -15
rect 17200 -35 17240 -15
rect 17274 -35 17314 -15
rect 17348 -35 17388 -15
rect 17422 -35 17462 -15
rect 17496 -35 17536 -15
rect 17570 -35 17610 -15
rect 17644 -35 17684 -15
rect 17718 -35 17758 -15
rect 16933 -42 16944 -35
rect 15861 -80 15873 -42
rect 15925 -80 16881 -42
rect 16933 -80 16946 -42
rect 15862 -87 15873 -80
rect 15048 -107 15088 -87
rect 15122 -107 15162 -87
rect 15196 -107 15236 -87
rect 15270 -107 15310 -87
rect 15344 -107 15384 -87
rect 15418 -107 15458 -87
rect 15492 -107 15532 -87
rect 15566 -107 15606 -87
rect 15640 -107 15680 -87
rect 15714 -107 15754 -87
rect 15788 -107 15828 -87
rect 15862 -107 15902 -87
rect 15157 -114 15162 -107
rect 11154 -158 11166 -114
rect 11218 -158 11230 -114
rect 11282 -145 13059 -114
tri 13059 -145 13090 -114 nw
tri 13232 -145 13263 -114 ne
rect 13263 -145 15040 -114
rect 11282 -158 13043 -145
rect 10037 -161 13043 -158
tri 13043 -161 13059 -145 nw
tri 13263 -161 13279 -145 ne
rect 13279 -159 15040 -145
rect 15092 -159 15105 -114
rect 15157 -159 15169 -114
rect 15221 -159 15233 -107
rect 15285 -159 15297 -107
rect 15349 -159 15361 -107
rect 15418 -114 15425 -107
rect 15605 -114 15606 -107
rect 15669 -114 15680 -107
rect 15413 -159 15425 -114
rect 15477 -159 15489 -114
rect 15541 -159 15553 -114
rect 15605 -159 15617 -114
rect 15669 -159 15681 -114
rect 15733 -159 15745 -107
rect 15797 -159 15809 -107
rect 15862 -114 15873 -107
rect 15936 -114 15976 -80
rect 16010 -114 16050 -80
rect 16084 -114 16124 -80
rect 16158 -114 16198 -80
rect 16232 -114 16574 -80
rect 16608 -114 16648 -80
rect 16682 -114 16722 -80
rect 16756 -114 16796 -80
rect 16830 -114 16870 -80
rect 16933 -87 16944 -80
rect 16998 -87 17010 -35
rect 17062 -87 17074 -35
rect 17126 -87 17138 -35
rect 17200 -42 17202 -35
rect 17382 -42 17388 -35
rect 17190 -80 17202 -42
rect 17254 -80 17266 -42
rect 17318 -80 17330 -42
rect 17382 -80 17394 -42
rect 17200 -87 17202 -80
rect 17382 -87 17388 -80
rect 17446 -87 17458 -35
rect 17510 -87 17522 -35
rect 17574 -87 17586 -35
rect 17644 -42 17650 -35
rect 17792 -42 17832 -8
rect 17866 -42 17906 -8
rect 17940 -42 17980 -8
rect 18014 -42 18053 -8
rect 18087 -42 18126 -8
rect 18160 -42 18199 -8
rect 18233 -42 18272 -8
rect 18306 -42 18345 -8
rect 18379 -42 18418 -8
rect 18452 -42 18491 -8
rect 18525 -42 18564 -8
rect 18598 -42 18637 -8
rect 18671 -42 18710 -8
rect 18744 -42 18783 -8
rect 18817 -42 18856 -8
rect 18890 -42 18929 -8
rect 18963 -42 19002 -8
rect 19036 -42 19075 -8
rect 19109 -42 19148 -8
rect 19182 -42 19221 -8
rect 19255 -42 19294 -8
rect 19328 -42 19367 -8
rect 19401 -42 19440 -8
rect 19474 -42 19574 -8
rect 17638 -80 17650 -42
rect 17702 -80 17714 -42
rect 17766 -80 19574 -42
rect 17644 -87 17650 -80
rect 16904 -107 16944 -87
rect 16978 -107 17018 -87
rect 17052 -107 17092 -87
rect 17126 -107 17166 -87
rect 17200 -107 17240 -87
rect 17274 -107 17314 -87
rect 17348 -107 17388 -87
rect 17422 -107 17462 -87
rect 17496 -107 17536 -87
rect 17570 -107 17610 -87
rect 17644 -107 17684 -87
rect 17718 -107 17758 -87
rect 16933 -114 16944 -107
rect 15861 -159 15873 -114
rect 15925 -145 16301 -114
tri 16301 -145 16332 -114 nw
tri 16474 -145 16505 -114 ne
rect 16505 -145 16881 -114
rect 15925 -159 16285 -145
rect 13279 -161 16285 -159
tri 16285 -161 16301 -145 nw
tri 16505 -161 16521 -145 ne
rect 16521 -159 16881 -145
rect 16933 -159 16946 -114
rect 16998 -159 17010 -107
rect 17062 -159 17074 -107
rect 17126 -159 17138 -107
rect 17200 -114 17202 -107
rect 17382 -114 17388 -107
rect 17190 -159 17202 -114
rect 17254 -159 17266 -114
rect 17318 -159 17330 -114
rect 17382 -159 17394 -114
rect 17446 -159 17458 -107
rect 17510 -159 17522 -107
rect 17574 -159 17586 -107
rect 17644 -114 17650 -107
rect 17792 -114 17832 -80
rect 17866 -114 17906 -80
rect 17940 -114 17980 -80
rect 18014 -114 18053 -80
rect 18087 -114 18126 -80
rect 18160 -114 18199 -80
rect 18233 -114 18272 -80
rect 18306 -114 18345 -80
rect 18379 -114 18418 -80
rect 18452 -114 18491 -80
rect 18525 -114 18564 -80
rect 18598 -114 18637 -80
rect 18671 -114 18710 -80
rect 18744 -114 18783 -80
rect 18817 -114 18856 -80
rect 18890 -114 18929 -80
rect 18963 -114 19002 -80
rect 19036 -114 19075 -80
rect 19109 -114 19148 -80
rect 19182 -114 19221 -80
rect 19255 -114 19294 -80
rect 19328 -114 19367 -80
rect 19401 -114 19440 -80
rect 19474 -114 19574 -80
rect 17638 -159 17650 -114
rect 17702 -159 17714 -114
rect 17766 -145 19543 -114
tri 19543 -145 19574 -114 nw
rect 19759 -18 19811 1087
rect 19759 -82 19811 -70
rect 19759 -140 19811 -134
rect 19841 1194 19971 1233
rect 19841 1160 19882 1194
rect 19916 1160 19971 1194
rect 19841 1121 19971 1160
rect 19841 1087 19882 1121
rect 19916 1087 19971 1121
rect 19841 1048 19971 1087
rect 19841 1014 19882 1048
rect 19916 1014 19971 1048
rect 19841 975 19971 1014
rect 19841 941 19882 975
rect 19916 941 19971 975
rect 19841 902 19971 941
rect 19841 868 19882 902
rect 19916 868 19971 902
rect 19841 829 19971 868
rect 19841 795 19882 829
rect 19916 795 19971 829
rect 19841 756 19971 795
rect 19841 722 19882 756
rect 19916 722 19971 756
rect 19841 683 19971 722
rect 19841 649 19882 683
rect 19916 649 19971 683
rect 19841 610 19971 649
rect 19841 576 19882 610
rect 19916 576 19971 610
rect 19841 537 19971 576
rect 19841 503 19882 537
rect 19916 503 19971 537
rect 19841 465 19971 503
rect 19841 431 19882 465
rect 19916 431 19971 465
rect 19841 393 19971 431
rect 19841 359 19882 393
rect 19916 359 19971 393
rect 19841 321 19971 359
rect 19841 287 19882 321
rect 19916 287 19971 321
rect 19841 249 19971 287
rect 19841 215 19882 249
rect 19916 215 19971 249
rect 19841 177 19971 215
rect 19841 143 19882 177
rect 19916 143 19971 177
rect 19841 105 19971 143
rect 20006 1027 20058 2991
rect 20006 963 20058 975
rect 20006 615 20058 911
rect 20006 551 20058 563
rect 20006 234 20058 499
rect 20006 170 20058 182
rect 20006 112 20058 118
rect 20198 1027 20250 1035
rect 20198 963 20250 975
rect 19841 71 19882 105
rect 19916 71 19971 105
rect 19841 33 19971 71
rect 19841 -1 19882 33
rect 19916 -1 19971 33
rect 19841 -39 19971 -1
rect 19841 -73 19882 -39
rect 19916 -73 19971 -39
rect 20006 63 20058 71
rect 20006 -1 20058 11
rect 20006 -59 20058 -53
rect 19841 -111 19971 -73
rect 19841 -145 19882 -111
rect 19916 -145 19971 -111
rect 17766 -159 19527 -145
rect 16521 -161 19527 -159
tri 19527 -161 19543 -145 nw
rect -52 -215 82 -183
tri 82 -215 135 -162 sw
tri 19788 -215 19841 -162 se
rect 19841 -215 19971 -145
rect -52 -228 19971 -215
rect -52 -229 12502 -228
rect -52 -238 673 -229
rect 725 -238 747 -229
rect 799 -238 821 -229
rect 873 -238 895 -229
rect 947 -238 6018 -229
rect 6070 -238 6085 -229
rect 6137 -238 6152 -229
rect 6204 -238 6219 -229
rect 6271 -238 6286 -229
rect 6338 -238 6353 -229
rect 6405 -238 6949 -229
rect 7001 -238 7016 -229
rect 7068 -238 7083 -229
rect 7135 -238 7150 -229
rect 7202 -238 7217 -229
rect 7269 -238 7284 -229
rect 7336 -238 12502 -229
rect 12554 -238 12569 -228
rect 12621 -238 12636 -228
rect 12688 -238 12703 -228
rect 12755 -238 12770 -228
rect 12822 -238 12837 -228
rect 12889 -229 19971 -228
rect 12889 -238 13433 -229
rect 13485 -238 13500 -229
rect 13552 -238 13567 -229
rect 13619 -238 13634 -229
rect 13686 -238 13701 -229
rect 13753 -238 13768 -229
rect 13820 -238 19071 -229
rect 19123 -238 19155 -229
rect -52 -267 8 -238
tri -52 -268 -51 -267 ne
rect -51 -268 8 -267
tri -51 -272 -47 -268 ne
rect -47 -272 8 -268
rect 42 -272 80 -238
rect 114 -272 152 -238
rect 186 -272 224 -238
rect 258 -272 296 -238
rect 330 -272 368 -238
rect 402 -272 440 -238
rect 474 -272 512 -238
rect 546 -272 584 -238
rect 618 -272 656 -238
rect 725 -272 728 -238
rect 799 -272 800 -238
rect 978 -272 1016 -238
rect 1050 -272 1088 -238
rect 1122 -272 1160 -238
rect 1194 -272 1232 -238
rect 1266 -272 1304 -238
rect 1338 -272 1376 -238
rect 1410 -272 1448 -238
rect 1482 -272 1520 -238
rect 1554 -272 1592 -238
rect 1626 -272 1664 -238
rect 1698 -272 1736 -238
rect 1770 -272 1808 -238
rect 1842 -272 1880 -238
rect 1914 -272 1952 -238
rect 1986 -272 2024 -238
rect 2058 -272 2096 -238
rect 2130 -272 2168 -238
rect 2202 -272 2240 -238
rect 2274 -272 2312 -238
rect 2346 -272 2384 -238
rect 2418 -272 2456 -238
rect 2490 -272 2528 -238
rect 2562 -272 2600 -238
rect 2634 -272 2672 -238
rect 2706 -272 2744 -238
rect 2778 -272 2816 -238
rect 2850 -272 2888 -238
rect 2922 -272 2960 -238
rect 2994 -272 3032 -238
rect 3066 -272 3104 -238
rect 3138 -272 3176 -238
rect 3210 -272 3248 -238
rect 3282 -272 3320 -238
rect 3354 -272 3392 -238
rect 3426 -272 3464 -238
rect 3498 -272 3536 -238
rect 3570 -272 3608 -238
rect 3642 -272 3680 -238
rect 3714 -272 3752 -238
rect 3786 -272 3824 -238
rect 3858 -272 3896 -238
rect 3930 -272 3968 -238
rect 4002 -272 4040 -238
rect 4074 -272 4112 -238
rect 4146 -272 4184 -238
rect 4218 -272 4256 -238
rect 4290 -272 4328 -238
rect 4362 -272 4400 -238
rect 4434 -272 4472 -238
rect 4506 -272 4544 -238
rect 4578 -272 4616 -238
rect 4650 -272 4688 -238
rect 4722 -272 4760 -238
rect 4794 -272 4832 -238
rect 4866 -272 4904 -238
rect 4938 -272 4976 -238
rect 5010 -272 5048 -238
rect 5082 -272 5120 -238
rect 5154 -272 5192 -238
rect 5226 -272 5264 -238
rect 5298 -272 5336 -238
rect 5370 -272 5408 -238
rect 5442 -272 5480 -238
rect 5514 -272 5552 -238
rect 5586 -272 5624 -238
rect 5658 -272 5696 -238
rect 5730 -272 5768 -238
rect 5802 -272 5840 -238
rect 5874 -272 5912 -238
rect 5946 -272 5984 -238
rect 6271 -272 6272 -238
rect 6338 -272 6344 -238
rect 6405 -272 6416 -238
rect 6450 -272 6488 -238
rect 6522 -272 6560 -238
rect 6594 -272 6632 -238
rect 6666 -272 6704 -238
rect 6738 -272 6776 -238
rect 6810 -272 6848 -238
rect 6882 -272 6920 -238
rect 7135 -272 7136 -238
rect 7202 -272 7208 -238
rect 7269 -272 7280 -238
rect 7336 -272 7352 -238
rect 7386 -272 7424 -238
rect 7458 -272 7496 -238
rect 7530 -272 7568 -238
rect 7602 -272 7640 -238
rect 7674 -272 7712 -238
rect 7746 -272 7784 -238
rect 7818 -272 7856 -238
rect 7890 -272 7928 -238
rect 7962 -272 8000 -238
rect 8034 -272 8072 -238
rect 8106 -272 8144 -238
rect 8178 -272 8216 -238
rect 8250 -272 8288 -238
rect 8322 -272 8360 -238
rect 8394 -272 8432 -238
rect 8466 -272 8504 -238
rect 8538 -272 8576 -238
rect 8610 -272 8648 -238
rect 8682 -272 8720 -238
rect 8754 -272 8792 -238
rect 8826 -272 8864 -238
rect 8898 -272 8936 -238
rect 8970 -272 9008 -238
rect 9042 -272 9080 -238
rect 9114 -272 9152 -238
rect 9186 -272 9224 -238
rect 9258 -272 9296 -238
rect 9330 -272 9368 -238
rect 9402 -272 9440 -238
rect 9474 -272 9512 -238
rect 9546 -272 9584 -238
rect 9618 -272 9656 -238
rect 9690 -272 9728 -238
rect 9762 -272 9800 -238
rect 9834 -272 9872 -238
rect 9906 -272 9944 -238
rect 9978 -272 10016 -238
rect 10050 -272 10088 -238
rect 10122 -272 10160 -238
rect 10194 -272 10232 -238
rect 10266 -272 10304 -238
rect 10338 -272 10376 -238
rect 10410 -272 10448 -238
rect 10482 -272 10520 -238
rect 10554 -272 10592 -238
rect 10626 -272 10664 -238
rect 10698 -272 10736 -238
rect 10770 -272 10808 -238
rect 10842 -272 10880 -238
rect 10914 -272 10952 -238
rect 10986 -272 11024 -238
rect 11058 -272 11096 -238
rect 11130 -272 11168 -238
rect 11202 -272 11240 -238
rect 11274 -272 11312 -238
rect 11346 -272 11384 -238
rect 11418 -272 11456 -238
rect 11490 -272 11528 -238
rect 11562 -272 11600 -238
rect 11634 -272 11672 -238
rect 11706 -272 11744 -238
rect 11778 -272 11816 -238
rect 11850 -272 11888 -238
rect 11922 -272 11960 -238
rect 11994 -272 12032 -238
rect 12066 -272 12104 -238
rect 12138 -272 12176 -238
rect 12210 -272 12248 -238
rect 12282 -272 12320 -238
rect 12354 -272 12392 -238
rect 12426 -272 12464 -238
rect 12498 -272 12502 -238
rect 12822 -272 12824 -238
rect 12889 -272 12896 -238
rect 12930 -272 12968 -238
rect 13002 -272 13040 -238
rect 13074 -272 13112 -238
rect 13146 -272 13184 -238
rect 13218 -272 13256 -238
rect 13290 -272 13328 -238
rect 13362 -272 13400 -238
rect 13686 -272 13688 -238
rect 13753 -272 13760 -238
rect 13820 -272 13832 -238
rect 13866 -272 13904 -238
rect 13938 -272 13976 -238
rect 14010 -272 14048 -238
rect 14082 -272 14120 -238
rect 14154 -272 14192 -238
rect 14226 -272 14264 -238
rect 14298 -272 14336 -238
rect 14370 -272 14408 -238
rect 14442 -272 14480 -238
rect 14514 -272 14552 -238
rect 14586 -272 14624 -238
rect 14658 -272 14696 -238
rect 14730 -272 14768 -238
rect 14802 -272 14840 -238
rect 14874 -272 14912 -238
rect 14946 -272 14984 -238
rect 15018 -272 15056 -238
rect 15090 -272 15128 -238
rect 15162 -272 15200 -238
rect 15234 -272 15272 -238
rect 15306 -272 15344 -238
rect 15378 -272 15416 -238
rect 15450 -272 15488 -238
rect 15522 -272 15560 -238
rect 15594 -272 15632 -238
rect 15666 -272 15704 -238
rect 15738 -272 15776 -238
rect 15810 -272 15848 -238
rect 15882 -272 15920 -238
rect 15954 -272 15992 -238
rect 16026 -272 16064 -238
rect 16098 -272 16136 -238
rect 16170 -272 16208 -238
rect 16242 -272 16280 -238
rect 16314 -272 16352 -238
rect 16386 -272 16424 -238
rect 16458 -272 16496 -238
rect 16530 -272 16568 -238
rect 16602 -272 16640 -238
rect 16674 -272 16712 -238
rect 16746 -272 16784 -238
rect 16818 -272 16856 -238
rect 16890 -272 16928 -238
rect 16962 -272 17000 -238
rect 17034 -272 17072 -238
rect 17106 -272 17144 -238
rect 17178 -272 17216 -238
rect 17250 -272 17288 -238
rect 17322 -272 17360 -238
rect 17394 -272 17432 -238
rect 17466 -272 17504 -238
rect 17538 -272 17576 -238
rect 17610 -272 17648 -238
rect 17682 -272 17720 -238
rect 17754 -272 17792 -238
rect 17826 -272 17864 -238
rect 17898 -272 17936 -238
rect 17970 -272 18008 -238
rect 18042 -272 18080 -238
rect 18114 -272 18152 -238
rect 18186 -272 18224 -238
rect 18258 -272 18296 -238
rect 18330 -272 18368 -238
rect 18402 -272 18440 -238
rect 18474 -272 18513 -238
rect 18547 -272 18586 -238
rect 18620 -272 18659 -238
rect 18693 -272 18732 -238
rect 18766 -272 18805 -238
rect 18839 -272 18878 -238
rect 18912 -272 18951 -238
rect 18985 -272 19024 -238
rect 19058 -272 19071 -238
rect 19131 -272 19155 -238
tri -47 -295 -24 -272 ne
rect -24 -281 673 -272
rect 725 -281 747 -272
rect 799 -281 821 -272
rect 873 -281 895 -272
rect 947 -281 6018 -272
rect 6070 -281 6085 -272
rect 6137 -281 6152 -272
rect 6204 -281 6219 -272
rect 6271 -281 6286 -272
rect 6338 -281 6353 -272
rect 6405 -281 6949 -272
rect 7001 -281 7016 -272
rect 7068 -281 7083 -272
rect 7135 -281 7150 -272
rect 7202 -281 7217 -272
rect 7269 -281 7284 -272
rect 7336 -280 12502 -272
rect 12554 -280 12569 -272
rect 12621 -280 12636 -272
rect 12688 -280 12703 -272
rect 12755 -280 12770 -272
rect 12822 -280 12837 -272
rect 12889 -280 13433 -272
rect 7336 -281 13433 -280
rect 13485 -281 13500 -272
rect 13552 -281 13567 -272
rect 13619 -281 13634 -272
rect 13686 -281 13701 -272
rect 13753 -281 13768 -272
rect 13820 -281 19071 -272
rect 19123 -281 19155 -272
rect 19207 -281 19238 -229
rect 19290 -238 19321 -229
rect 19373 -238 19971 -229
rect 19290 -272 19316 -238
rect 19373 -272 19389 -238
rect 19423 -272 19462 -238
rect 19496 -272 19535 -238
rect 19569 -272 19608 -238
rect 19642 -272 19681 -238
rect 19715 -272 19754 -238
rect 19788 -272 19827 -238
rect 19861 -272 19971 -238
rect 19290 -281 19321 -272
rect 19373 -281 19971 -272
rect -24 -295 19971 -281
tri -24 -345 26 -295 ne
rect 26 -345 19971 -295
rect 3708 -469 3714 -417
rect 3766 -469 3778 -417
rect 3830 -469 3836 -417
tri 3742 -503 3776 -469 ne
rect 3776 -838 3836 -469
tri 20191 -808 20198 -801 se
rect 20198 -808 20250 911
rect 20430 222 20482 228
rect 20430 158 20482 170
rect 20430 63 20482 106
tri 20482 63 20504 85 sw
rect 20430 58 20504 63
tri 20504 58 20509 63 sw
rect 22755 58 22871 63
rect 20430 57 22871 58
rect 20430 -22 22755 57
rect 22755 -65 22871 -59
tri 3836 -838 3866 -808 sw
tri 20161 -838 20191 -808 se
rect 20191 -838 20250 -808
rect 3776 -842 20250 -838
tri 3776 -874 3808 -842 ne
rect 3808 -872 20250 -842
rect 3808 -874 5849 -872
tri 5849 -874 5851 -872 nw
rect -2190 -2789 -2049 -2651
rect 15039 -2923 15045 -2871
rect 15097 -2923 15113 -2871
rect 15165 -2923 15181 -2871
rect 15233 -2923 15249 -2871
rect 15301 -2923 15317 -2871
rect 15369 -2923 15385 -2871
rect 15437 -2923 15453 -2871
rect 15505 -2923 15521 -2871
rect 15573 -2923 15589 -2871
rect 15641 -2923 15657 -2871
rect 15709 -2923 15725 -2871
rect 15777 -2923 15793 -2871
rect 15845 -2923 15861 -2871
rect 15913 -2923 15919 -2871
rect 16880 -2923 16886 -2871
rect 16938 -2923 16954 -2871
rect 17006 -2923 17022 -2871
rect 17074 -2923 17090 -2871
rect 17142 -2923 17158 -2871
rect 17210 -2923 17226 -2871
rect 17278 -2923 17294 -2871
rect 17346 -2923 17362 -2871
rect 17414 -2923 17430 -2871
rect 17482 -2923 17498 -2871
rect 17550 -2923 17566 -2871
rect 17618 -2923 17634 -2871
rect 17686 -2923 17702 -2871
rect 17754 -2923 17760 -2871
tri 14953 -3009 15039 -2923 se
rect 15039 -3009 15919 -2923
tri 15919 -3009 16005 -2923 sw
tri 16794 -3009 16880 -2923 se
rect 16880 -3009 17760 -2923
tri 17760 -3009 17846 -2923 sw
rect -2635 -3184 -2456 -3020
<< rmetal1 >>
rect 6648 1451 6650 1452
rect 6648 1407 6649 1451
rect 6648 1406 6650 1407
rect 6710 1451 6712 1452
rect 6711 1407 6712 1451
rect 6710 1406 6712 1407
<< via1 >>
rect -1604 14163 -1599 14169
rect -1599 14163 -1555 14169
rect -1555 14163 -1552 14169
rect -1511 14163 -1477 14169
rect -1477 14163 -1459 14169
rect -1418 14163 -1399 14169
rect -1399 14163 -1366 14169
rect -1604 14125 -1552 14163
rect -1511 14125 -1459 14163
rect -1418 14125 -1366 14163
rect -1604 14117 -1599 14125
rect -1599 14117 -1555 14125
rect -1555 14117 -1552 14125
rect -1511 14117 -1477 14125
rect -1477 14117 -1459 14125
rect -1418 14117 -1399 14125
rect -1399 14117 -1366 14125
rect -1606 11961 -1554 11973
rect -1606 11927 -1597 11961
rect -1597 11927 -1563 11961
rect -1563 11927 -1554 11961
rect -1606 11921 -1554 11927
rect -1606 11889 -1554 11909
rect -1606 11857 -1597 11889
rect -1597 11857 -1563 11889
rect -1563 11857 -1554 11889
rect -1450 12287 -1441 12311
rect -1441 12287 -1407 12311
rect -1407 12287 -1398 12311
rect -1450 12259 -1398 12287
rect -1450 12215 -1441 12247
rect -1441 12215 -1407 12247
rect -1407 12215 -1398 12247
rect -1450 12195 -1398 12215
rect -1450 12177 -1398 12183
rect -1450 12143 -1441 12177
rect -1441 12143 -1407 12177
rect -1407 12143 -1398 12177
rect -1450 12131 -1398 12143
rect -1606 11817 -1554 11845
rect -1606 11793 -1597 11817
rect -1597 11793 -1563 11817
rect -1563 11793 -1554 11817
rect -1294 11961 -1242 11973
rect -1294 11927 -1285 11961
rect -1285 11927 -1251 11961
rect -1251 11927 -1242 11961
rect -1294 11921 -1242 11927
rect -1294 11889 -1242 11909
rect -1294 11857 -1285 11889
rect -1285 11857 -1251 11889
rect -1251 11857 -1242 11889
rect -1294 11817 -1242 11845
rect -1606 11625 -1597 11649
rect -1597 11625 -1563 11649
rect -1563 11625 -1554 11649
rect -1606 11597 -1554 11625
rect -1606 11553 -1597 11585
rect -1597 11553 -1563 11585
rect -1563 11553 -1554 11585
rect -1606 11533 -1554 11553
rect -1606 11515 -1554 11521
rect -1606 11481 -1597 11515
rect -1597 11481 -1563 11515
rect -1563 11481 -1554 11515
rect -1606 11469 -1554 11481
rect -1294 11793 -1285 11817
rect -1285 11793 -1251 11817
rect -1251 11793 -1242 11817
rect -1450 11299 -1398 11311
rect -1450 11265 -1441 11299
rect -1441 11265 -1407 11299
rect -1407 11265 -1398 11299
rect -1450 11259 -1398 11265
rect -1450 11227 -1398 11247
rect -1450 11195 -1441 11227
rect -1441 11195 -1407 11227
rect -1407 11195 -1398 11227
rect -1450 11155 -1398 11183
rect -1450 11131 -1441 11155
rect -1441 11131 -1407 11155
rect -1407 11131 -1398 11155
rect -1294 11625 -1285 11649
rect -1285 11625 -1251 11649
rect -1251 11625 -1242 11649
rect -1294 11597 -1242 11625
rect -1294 11553 -1285 11585
rect -1285 11553 -1251 11585
rect -1251 11553 -1242 11585
rect -1294 11533 -1242 11553
rect -1294 11515 -1242 11521
rect -1294 11481 -1285 11515
rect -1285 11481 -1251 11515
rect -1251 11481 -1242 11515
rect -1294 11469 -1242 11481
rect -1606 10497 -1554 10509
rect -1606 10463 -1597 10497
rect -1597 10463 -1563 10497
rect -1563 10463 -1554 10497
rect -1606 10457 -1554 10463
rect -1606 10425 -1554 10445
rect -1606 10393 -1597 10425
rect -1597 10393 -1563 10425
rect -1563 10393 -1554 10425
rect -1606 10353 -1554 10381
rect -1606 10329 -1597 10353
rect -1597 10329 -1563 10353
rect -1563 10329 -1554 10353
rect -1450 10823 -1441 10847
rect -1441 10823 -1407 10847
rect -1407 10823 -1398 10847
rect -1450 10795 -1398 10823
rect -1450 10751 -1441 10783
rect -1441 10751 -1407 10783
rect -1407 10751 -1398 10783
rect -1450 10731 -1398 10751
rect -1450 10713 -1398 10719
rect -1450 10679 -1441 10713
rect -1441 10679 -1407 10713
rect -1407 10679 -1398 10713
rect -1450 10667 -1398 10679
rect -1294 10497 -1242 10509
rect -1294 10463 -1285 10497
rect -1285 10463 -1251 10497
rect -1251 10463 -1242 10497
rect -1294 10457 -1242 10463
rect -1294 10425 -1242 10445
rect -1294 10393 -1285 10425
rect -1285 10393 -1251 10425
rect -1251 10393 -1242 10425
rect -1294 10353 -1242 10381
rect -1294 10329 -1285 10353
rect -1285 10329 -1251 10353
rect -1251 10329 -1242 10353
rect -957 6171 -905 6223
rect -957 6096 -905 6148
rect 21783 6165 21835 6171
rect 21847 6165 21899 6171
rect 19690 6117 19742 6126
rect 19690 6083 19693 6117
rect 19693 6083 19727 6117
rect 19727 6083 19742 6117
rect 19690 6074 19742 6083
rect 19757 6117 19809 6126
rect 19757 6083 19765 6117
rect 19765 6083 19799 6117
rect 19799 6083 19809 6117
rect 19757 6074 19809 6083
rect 19824 6074 19876 6126
rect 21783 6119 21789 6165
rect 21789 6119 21835 6165
rect 21847 6119 21895 6165
rect 21895 6119 21899 6165
rect 21783 6059 21789 6104
rect 21789 6059 21835 6104
rect 21847 6059 21895 6104
rect 21895 6059 21899 6104
rect 21783 6052 21835 6059
rect 21847 6052 21899 6059
rect -1636 5780 -1584 5832
rect -1636 5705 -1584 5757
rect 19690 5490 19742 5499
rect 19690 5456 19693 5490
rect 19693 5456 19727 5490
rect 19727 5456 19742 5490
rect 19690 5447 19742 5456
rect 19754 5490 19806 5499
rect 19754 5456 19765 5490
rect 19765 5456 19799 5490
rect 19799 5456 19806 5490
rect 19754 5447 19806 5456
rect 3029 5079 3081 5131
rect 3095 5079 3147 5131
rect 3161 5079 3213 5131
rect 3227 5079 3279 5131
rect 3293 5079 3345 5131
rect 3358 5079 3410 5131
rect 3423 5079 3475 5131
rect 3488 5079 3540 5131
rect 3553 5079 3605 5131
rect 3618 5079 3670 5131
rect 3683 5079 3735 5131
rect 3748 5079 3800 5131
rect 3813 5079 3865 5131
rect 3878 5079 3930 5131
rect 3943 5079 3995 5131
rect 4008 5079 4060 5131
rect 4073 5079 4125 5131
rect 4138 5079 4190 5131
rect 4203 5079 4255 5131
rect 4268 5079 4320 5131
rect 3029 4963 3081 5015
rect 3095 4963 3147 5015
rect 3161 4963 3213 5015
rect 3227 4963 3279 5015
rect 3293 4963 3345 5015
rect 3358 4963 3410 5015
rect 3423 4963 3475 5015
rect 3488 4963 3540 5015
rect 3553 4963 3605 5015
rect 3618 4963 3670 5015
rect 3683 4963 3735 5015
rect 3748 4963 3800 5015
rect 3813 4963 3865 5015
rect 3878 4963 3930 5015
rect 3943 4963 3995 5015
rect 4008 4963 4060 5015
rect 4073 4963 4125 5015
rect 4138 4963 4190 5015
rect 4203 4963 4255 5015
rect 4268 4963 4320 5015
rect 8560 5079 8612 5131
rect 8627 5079 8679 5131
rect 8694 5079 8746 5131
rect 8761 5079 8813 5131
rect 8828 5079 8880 5131
rect 8895 5079 8947 5131
rect 8962 5079 9014 5131
rect 9028 5079 9080 5131
rect 9094 5079 9146 5131
rect 9160 5079 9212 5131
rect 9226 5079 9278 5131
rect 9292 5079 9344 5131
rect 9358 5079 9410 5131
rect 9424 5079 9476 5131
rect 9490 5079 9542 5131
rect 9556 5079 9608 5131
rect 8560 4963 8612 5015
rect 8627 4963 8679 5015
rect 8694 4963 8746 5015
rect 8761 4963 8813 5015
rect 8828 4963 8880 5015
rect 8895 4963 8947 5015
rect 8962 4963 9014 5015
rect 9028 4963 9080 5015
rect 9094 4963 9146 5015
rect 9160 4963 9212 5015
rect 9226 4963 9278 5015
rect 9292 4963 9344 5015
rect 9358 4963 9410 5015
rect 9424 4963 9476 5015
rect 9490 4963 9542 5015
rect 9556 4963 9608 5015
rect 11014 5079 11066 5131
rect 11082 5079 11134 5131
rect 11150 5079 11202 5131
rect 11217 5079 11269 5131
rect 11014 4963 11066 5015
rect 11082 4963 11134 5015
rect 11150 4963 11202 5015
rect 11217 4963 11269 5015
rect 15049 5079 15101 5131
rect 15118 5079 15170 5131
rect 15187 5079 15239 5131
rect 15255 5079 15307 5131
rect 15323 5079 15375 5131
rect 15391 5079 15443 5131
rect 15459 5079 15511 5131
rect 15527 5079 15579 5131
rect 15595 5079 15647 5131
rect 15663 5079 15715 5131
rect 15731 5079 15783 5131
rect 15799 5079 15851 5131
rect 15867 5079 15919 5131
rect 15049 4963 15101 5015
rect 15118 4963 15170 5015
rect 15187 4963 15239 5015
rect 15255 4963 15307 5015
rect 15323 4963 15375 5015
rect 15391 4963 15443 5015
rect 15459 4963 15511 5015
rect 15527 4963 15579 5015
rect 15595 4963 15647 5015
rect 15663 4963 15715 5015
rect 15731 4963 15783 5015
rect 15799 4963 15851 5015
rect 15867 4963 15919 5015
rect 16888 5079 16940 5131
rect 16957 5079 17009 5131
rect 17026 5079 17078 5131
rect 17094 5079 17146 5131
rect 17162 5079 17214 5131
rect 17230 5079 17282 5131
rect 17298 5079 17350 5131
rect 17366 5079 17418 5131
rect 17434 5079 17486 5131
rect 17502 5079 17554 5131
rect 17570 5079 17622 5131
rect 17638 5079 17690 5131
rect 17706 5079 17758 5131
rect 16888 4963 16940 5015
rect 16957 4963 17009 5015
rect 17026 4963 17078 5015
rect 17094 4963 17146 5015
rect 17162 4963 17214 5015
rect 17230 4963 17282 5015
rect 17298 4963 17350 5015
rect 17366 4963 17418 5015
rect 17434 4963 17486 5015
rect 17502 4963 17554 5015
rect 17570 4963 17622 5015
rect 17638 4963 17690 5015
rect 17706 4963 17758 5015
rect 19671 5079 19723 5131
rect 19762 5079 19814 5131
rect 19671 4963 19723 5015
rect 19762 4963 19814 5015
rect 3631 4706 3683 4758
rect 3698 4706 3750 4758
rect 3765 4706 3817 4758
rect 3832 4706 3884 4758
rect 3899 4706 3951 4758
rect 3966 4706 4018 4758
rect 4033 4706 4085 4758
rect 4099 4706 4151 4758
rect 4165 4706 4217 4758
rect 3631 4642 3683 4694
rect 3698 4642 3750 4694
rect 3765 4642 3817 4694
rect 3832 4642 3884 4694
rect 3899 4642 3951 4694
rect 3966 4642 4018 4694
rect 4033 4642 4085 4694
rect 4099 4642 4151 4694
rect 4165 4642 4217 4694
rect 3631 4578 3683 4630
rect 3698 4578 3750 4630
rect 3765 4578 3817 4630
rect 3832 4578 3884 4630
rect 3899 4578 3951 4630
rect 3966 4578 4018 4630
rect 4033 4578 4085 4630
rect 4099 4578 4151 4630
rect 4165 4578 4217 4630
rect -1176 4474 -1124 4526
rect -1176 4410 -1124 4462
rect -1078 4406 -1026 4458
rect -1014 4406 -962 4458
rect 649 4295 701 4347
rect 725 4295 777 4347
rect 800 4295 852 4347
rect 649 4215 701 4267
rect 725 4215 777 4267
rect 800 4215 852 4267
rect 6018 4295 6070 4347
rect 6085 4295 6137 4347
rect 6152 4295 6204 4347
rect 6219 4295 6271 4347
rect 6286 4295 6338 4347
rect 6353 4295 6405 4347
rect 6018 4215 6070 4267
rect 6085 4215 6137 4267
rect 6152 4215 6204 4267
rect 6219 4215 6271 4267
rect 6286 4215 6338 4267
rect 6353 4215 6405 4267
rect 6949 4295 7001 4347
rect 7016 4295 7068 4347
rect 7083 4295 7135 4347
rect 7150 4295 7202 4347
rect 7217 4295 7269 4347
rect 7284 4295 7336 4347
rect 6949 4215 7001 4267
rect 7016 4215 7068 4267
rect 7083 4215 7135 4267
rect 7150 4215 7202 4267
rect 7217 4215 7269 4267
rect 7284 4215 7336 4267
rect 12502 4295 12554 4347
rect 12569 4295 12621 4347
rect 12636 4295 12688 4347
rect 12703 4295 12755 4347
rect 12770 4295 12822 4347
rect 12837 4295 12889 4347
rect 12502 4215 12554 4267
rect 12569 4215 12621 4267
rect 12636 4215 12688 4267
rect 12703 4215 12755 4267
rect 12770 4215 12822 4267
rect 12837 4215 12889 4267
rect 13433 4295 13485 4347
rect 13500 4295 13552 4347
rect 13567 4295 13619 4347
rect 13634 4295 13686 4347
rect 13701 4295 13753 4347
rect 13768 4295 13820 4347
rect 13433 4215 13485 4267
rect 13500 4215 13552 4267
rect 13567 4215 13619 4267
rect 13634 4215 13686 4267
rect 13701 4215 13753 4267
rect 13768 4215 13820 4267
rect 19067 4295 19119 4347
rect 19152 4295 19204 4347
rect 19237 4295 19289 4347
rect 19321 4295 19373 4347
rect 19067 4215 19119 4267
rect 19152 4215 19204 4267
rect 19237 4215 19289 4267
rect 19321 4215 19373 4267
rect 19844 4192 19960 4372
rect -624 3333 -572 3385
rect -560 3333 -508 3385
rect -310 2965 -258 3017
rect -310 2901 -258 2953
rect 644 2928 696 2959
rect 728 2928 780 2959
rect 812 2928 864 2959
rect 895 2928 947 2959
rect 6018 2928 6070 2959
rect 6085 2928 6137 2959
rect 6152 2928 6204 2959
rect 644 2907 671 2928
rect 671 2907 696 2928
rect 728 2907 744 2928
rect 744 2907 780 2928
rect 812 2907 817 2928
rect 817 2907 856 2928
rect 856 2907 864 2928
rect 895 2907 929 2928
rect 929 2907 947 2928
rect 6018 2907 6037 2928
rect 6037 2907 6070 2928
rect 6085 2907 6109 2928
rect 6109 2907 6137 2928
rect 6152 2907 6181 2928
rect 6181 2907 6204 2928
rect 6219 2928 6271 2959
rect 6219 2907 6253 2928
rect 6253 2907 6271 2928
rect 6286 2928 6338 2959
rect 6286 2907 6291 2928
rect 6291 2907 6325 2928
rect 6325 2907 6338 2928
rect 6353 2928 6405 2959
rect 6949 2928 7001 2959
rect 7016 2928 7068 2959
rect 6353 2907 6363 2928
rect 6363 2907 6397 2928
rect 6397 2907 6405 2928
rect 6949 2907 6973 2928
rect 6973 2907 7001 2928
rect 7016 2907 7045 2928
rect 7045 2907 7068 2928
rect 7083 2928 7135 2959
rect 7083 2907 7117 2928
rect 7117 2907 7135 2928
rect 7150 2928 7202 2959
rect 7150 2907 7155 2928
rect 7155 2907 7189 2928
rect 7189 2907 7202 2928
rect 7217 2928 7269 2959
rect 7217 2907 7227 2928
rect 7227 2907 7261 2928
rect 7261 2907 7269 2928
rect 7284 2928 7336 2959
rect 12502 2928 12554 2959
rect 12569 2928 12621 2959
rect 12636 2928 12688 2959
rect 12703 2928 12755 2959
rect 7284 2907 7299 2928
rect 7299 2907 7333 2928
rect 7333 2907 7336 2928
rect 12502 2907 12517 2928
rect 12517 2907 12554 2928
rect 12569 2907 12589 2928
rect 12589 2907 12621 2928
rect 12636 2907 12661 2928
rect 12661 2907 12688 2928
rect 12703 2907 12733 2928
rect 12733 2907 12755 2928
rect 12770 2928 12822 2959
rect 12770 2907 12771 2928
rect 12771 2907 12805 2928
rect 12805 2907 12822 2928
rect 12837 2928 12889 2959
rect 13433 2928 13485 2959
rect 13500 2928 13552 2959
rect 13567 2928 13619 2959
rect 12837 2907 12843 2928
rect 12843 2907 12877 2928
rect 12877 2907 12889 2928
rect 13433 2907 13453 2928
rect 13453 2907 13485 2928
rect 13500 2907 13525 2928
rect 13525 2907 13552 2928
rect 13567 2907 13597 2928
rect 13597 2907 13619 2928
rect 13634 2928 13686 2959
rect 13634 2907 13635 2928
rect 13635 2907 13669 2928
rect 13669 2907 13686 2928
rect 13701 2928 13753 2959
rect 13701 2907 13707 2928
rect 13707 2907 13741 2928
rect 13741 2907 13753 2928
rect 13768 2928 13820 2959
rect 19071 2928 19123 2959
rect 19155 2928 19207 2959
rect 19238 2928 19290 2959
rect 13768 2907 13779 2928
rect 13779 2907 13813 2928
rect 13813 2907 13820 2928
rect 19071 2907 19107 2928
rect 19107 2907 19123 2928
rect 19155 2907 19179 2928
rect 19179 2907 19207 2928
rect 19238 2907 19251 2928
rect 19251 2907 19285 2928
rect 19285 2907 19290 2928
rect 19321 2928 19373 2959
rect 19321 2907 19323 2928
rect 19323 2907 19357 2928
rect 19357 2907 19373 2928
rect -1360 2823 -1308 2829
rect -1360 2789 -1329 2823
rect -1329 2789 -1308 2823
rect -1360 2777 -1308 2789
rect -1360 2750 -1308 2759
rect -1360 2716 -1329 2750
rect -1329 2716 -1308 2750
rect -1360 2707 -1308 2716
rect -1360 2676 -1308 2688
rect -1737 2593 -1685 2645
rect -1360 2642 -1329 2676
rect -1329 2642 -1308 2676
rect -1360 2636 -1308 2642
rect -1084 2777 -1032 2829
rect -1084 2707 -1032 2759
rect -466 2825 -414 2877
rect -466 2761 -414 2813
rect 644 2827 696 2879
rect 728 2827 780 2879
rect 812 2827 864 2879
rect 895 2827 947 2879
rect 6018 2827 6070 2879
rect 6085 2827 6137 2879
rect 6152 2827 6204 2879
rect 6219 2827 6271 2879
rect 6286 2827 6338 2879
rect 6353 2827 6405 2879
rect 6949 2827 7001 2879
rect 7016 2827 7068 2879
rect 7083 2827 7135 2879
rect 7150 2827 7202 2879
rect 7217 2827 7269 2879
rect 7284 2827 7336 2879
rect 12502 2827 12554 2879
rect 12569 2827 12621 2879
rect 12636 2827 12688 2879
rect 12703 2827 12755 2879
rect 12770 2827 12822 2879
rect 12837 2827 12889 2879
rect 13433 2827 13485 2879
rect 13500 2827 13552 2879
rect 13567 2827 13619 2879
rect 13634 2827 13686 2879
rect 13701 2827 13753 2879
rect 13768 2827 13820 2879
rect 19071 2827 19123 2879
rect 19155 2827 19207 2879
rect 19238 2827 19290 2879
rect 19321 2827 19373 2879
rect -1084 2636 -1032 2688
rect -1737 2529 -1685 2581
rect -222 2515 -170 2567
rect -310 2409 -258 2461
rect -222 2451 -170 2503
rect 644 2686 696 2738
rect 728 2686 780 2738
rect 812 2686 864 2738
rect 895 2686 947 2738
rect 644 2622 696 2674
rect 728 2622 780 2674
rect 812 2622 864 2674
rect 895 2622 947 2674
rect 644 2558 696 2610
rect 728 2558 780 2610
rect 812 2558 864 2610
rect 895 2558 947 2610
rect 6018 2686 6070 2738
rect 6085 2686 6137 2738
rect 6152 2686 6204 2738
rect 6219 2686 6271 2738
rect 6286 2686 6338 2738
rect 6353 2686 6405 2738
rect 6018 2622 6070 2674
rect 6085 2622 6137 2674
rect 6152 2622 6204 2674
rect 6219 2622 6271 2674
rect 6286 2622 6338 2674
rect 6353 2622 6405 2674
rect 6018 2558 6070 2610
rect 6085 2558 6137 2610
rect 6152 2558 6204 2610
rect 6219 2558 6271 2610
rect 6286 2558 6338 2610
rect 6353 2558 6405 2610
rect 6949 2686 7001 2738
rect 7016 2686 7068 2738
rect 7083 2686 7135 2738
rect 7150 2686 7202 2738
rect 7217 2686 7269 2738
rect 7284 2686 7336 2738
rect 6949 2622 7001 2674
rect 7016 2622 7068 2674
rect 7083 2622 7135 2674
rect 7150 2622 7202 2674
rect 7217 2622 7269 2674
rect 7284 2622 7336 2674
rect 6949 2558 7001 2610
rect 7016 2558 7068 2610
rect 7083 2558 7135 2610
rect 7150 2558 7202 2610
rect 7217 2558 7269 2610
rect 7284 2558 7336 2610
rect 12502 2686 12554 2738
rect 12569 2686 12621 2738
rect 12636 2686 12688 2738
rect 12703 2686 12755 2738
rect 12770 2686 12822 2738
rect 12837 2686 12889 2738
rect 12502 2622 12554 2674
rect 12569 2622 12621 2674
rect 12636 2622 12688 2674
rect 12703 2622 12755 2674
rect 12770 2622 12822 2674
rect 12837 2622 12889 2674
rect 12502 2558 12554 2610
rect 12569 2558 12621 2610
rect 12636 2558 12688 2610
rect 12703 2558 12755 2610
rect 12770 2558 12822 2610
rect 12837 2558 12889 2610
rect 13433 2686 13485 2738
rect 13500 2686 13552 2738
rect 13567 2686 13619 2738
rect 13634 2686 13686 2738
rect 13701 2686 13753 2738
rect 13768 2686 13820 2738
rect 13433 2622 13485 2674
rect 13500 2622 13552 2674
rect 13567 2622 13619 2674
rect 13634 2622 13686 2674
rect 13701 2622 13753 2674
rect 13768 2622 13820 2674
rect 13433 2558 13485 2610
rect 13500 2558 13552 2610
rect 13567 2558 13619 2610
rect 13634 2558 13686 2610
rect 13701 2558 13753 2610
rect 13768 2558 13820 2610
rect 19071 2686 19123 2738
rect 19154 2686 19206 2738
rect 19237 2686 19289 2738
rect 19321 2686 19373 2738
rect 19071 2622 19123 2674
rect 19154 2622 19206 2674
rect 19237 2622 19289 2674
rect 19321 2622 19373 2674
rect 19071 2558 19123 2610
rect 19154 2558 19206 2610
rect 19237 2558 19289 2610
rect 19321 2558 19373 2610
rect -1722 2348 -1670 2400
rect -310 2345 -258 2397
rect -1722 2284 -1670 2336
rect -1636 2029 -1584 2035
rect -1636 1995 -1607 2029
rect -1607 1995 -1584 2029
rect -1636 1983 -1584 1995
rect -1636 1956 -1584 1965
rect -1636 1922 -1607 1956
rect -1607 1922 -1584 1956
rect -466 2019 -414 2071
rect -466 1955 -414 2007
rect 1027 2385 1079 2437
rect 1092 2385 1144 2437
rect 1157 2385 1209 2437
rect 1222 2385 1274 2437
rect 1286 2385 1338 2437
rect 1350 2385 1402 2437
rect 1414 2385 1466 2437
rect 1478 2385 1530 2437
rect 1542 2385 1594 2437
rect 1606 2385 1658 2437
rect 1670 2385 1722 2437
rect 1734 2385 1786 2437
rect 1798 2385 1850 2437
rect 1862 2385 1914 2437
rect 1027 2317 1079 2369
rect 1092 2317 1144 2369
rect 1157 2317 1209 2369
rect 1222 2317 1274 2369
rect 1286 2317 1338 2369
rect 1350 2317 1402 2369
rect 1414 2317 1466 2369
rect 1478 2317 1530 2369
rect 1542 2317 1594 2369
rect 1606 2317 1658 2369
rect 1670 2317 1722 2369
rect 1734 2317 1786 2369
rect 1798 2317 1850 2369
rect 1862 2317 1914 2369
rect 1027 2249 1079 2301
rect 1092 2249 1144 2301
rect 1157 2249 1209 2301
rect 1222 2249 1274 2301
rect 1286 2249 1338 2301
rect 1350 2249 1402 2301
rect 1414 2249 1466 2301
rect 1478 2249 1530 2301
rect 1542 2249 1594 2301
rect 1606 2249 1658 2301
rect 1670 2249 1722 2301
rect 1734 2249 1786 2301
rect 1798 2249 1850 2301
rect 1862 2249 1914 2301
rect 1027 2181 1079 2233
rect 1092 2181 1144 2233
rect 1157 2181 1209 2233
rect 1222 2181 1274 2233
rect 1286 2181 1338 2233
rect 1350 2181 1402 2233
rect 1414 2181 1466 2233
rect 1478 2181 1530 2233
rect 1542 2181 1594 2233
rect 1606 2181 1658 2233
rect 1670 2181 1722 2233
rect 1734 2181 1786 2233
rect 1798 2181 1850 2233
rect 1862 2181 1914 2233
rect 1027 2113 1079 2165
rect 1092 2113 1144 2165
rect 1157 2113 1209 2165
rect 1222 2113 1274 2165
rect 1286 2113 1338 2165
rect 1350 2113 1402 2165
rect 1414 2113 1466 2165
rect 1478 2113 1530 2165
rect 1542 2113 1594 2165
rect 1606 2113 1658 2165
rect 1670 2113 1722 2165
rect 1734 2113 1786 2165
rect 1798 2113 1850 2165
rect 1862 2113 1914 2165
rect 1027 2045 1079 2097
rect 1092 2045 1144 2097
rect 1157 2045 1209 2097
rect 1222 2045 1274 2097
rect 1286 2045 1338 2097
rect 1350 2045 1402 2097
rect 1414 2045 1466 2097
rect 1478 2045 1530 2097
rect 1542 2045 1594 2097
rect 1606 2045 1658 2097
rect 1670 2045 1722 2097
rect 1734 2045 1786 2097
rect 1798 2045 1850 2097
rect 1862 2045 1914 2097
rect 7511 2385 7563 2437
rect 7576 2385 7628 2437
rect 7641 2385 7693 2437
rect 7706 2385 7758 2437
rect 7770 2385 7822 2437
rect 7834 2385 7886 2437
rect 7898 2385 7950 2437
rect 7962 2385 8014 2437
rect 8026 2385 8078 2437
rect 8090 2385 8142 2437
rect 8154 2385 8206 2437
rect 8218 2385 8270 2437
rect 8282 2385 8334 2437
rect 8346 2385 8398 2437
rect 7511 2317 7563 2369
rect 7576 2317 7628 2369
rect 7641 2317 7693 2369
rect 7706 2317 7758 2369
rect 7770 2317 7822 2369
rect 7834 2317 7886 2369
rect 7898 2317 7950 2369
rect 7962 2317 8014 2369
rect 8026 2317 8078 2369
rect 8090 2317 8142 2369
rect 8154 2317 8206 2369
rect 8218 2317 8270 2369
rect 8282 2317 8334 2369
rect 8346 2317 8398 2369
rect 7511 2249 7563 2301
rect 7576 2249 7628 2301
rect 7641 2249 7693 2301
rect 7706 2249 7758 2301
rect 7770 2249 7822 2301
rect 7834 2249 7886 2301
rect 7898 2249 7950 2301
rect 7962 2249 8014 2301
rect 8026 2249 8078 2301
rect 8090 2249 8142 2301
rect 8154 2249 8206 2301
rect 8218 2249 8270 2301
rect 8282 2249 8334 2301
rect 8346 2249 8398 2301
rect 7511 2181 7563 2233
rect 7576 2181 7628 2233
rect 7641 2181 7693 2233
rect 7706 2181 7758 2233
rect 7770 2181 7822 2233
rect 7834 2181 7886 2233
rect 7898 2181 7950 2233
rect 7962 2181 8014 2233
rect 8026 2181 8078 2233
rect 8090 2181 8142 2233
rect 8154 2181 8206 2233
rect 8218 2181 8270 2233
rect 8282 2181 8334 2233
rect 8346 2181 8398 2233
rect 7511 2113 7563 2165
rect 7576 2113 7628 2165
rect 7641 2113 7693 2165
rect 7706 2113 7758 2165
rect 7770 2113 7822 2165
rect 7834 2113 7886 2165
rect 7898 2113 7950 2165
rect 7962 2113 8014 2165
rect 8026 2113 8078 2165
rect 8090 2113 8142 2165
rect 8154 2113 8206 2165
rect 8218 2113 8270 2165
rect 8282 2113 8334 2165
rect 8346 2113 8398 2165
rect 7511 2045 7563 2097
rect 7576 2045 7628 2097
rect 7641 2045 7693 2097
rect 7706 2045 7758 2097
rect 7770 2045 7822 2097
rect 7834 2045 7886 2097
rect 7898 2045 7950 2097
rect 7962 2045 8014 2097
rect 8026 2045 8078 2097
rect 8090 2045 8142 2097
rect 8154 2045 8206 2097
rect 8218 2045 8270 2097
rect 8282 2045 8334 2097
rect 8346 2045 8398 2097
rect 11440 2385 11492 2437
rect 11504 2385 11556 2437
rect 11568 2385 11620 2437
rect 11632 2385 11684 2437
rect 11696 2385 11748 2437
rect 11760 2385 11812 2437
rect 11824 2385 11876 2437
rect 11888 2385 11940 2437
rect 11952 2385 12004 2437
rect 12016 2385 12068 2437
rect 12080 2385 12132 2437
rect 12145 2385 12197 2437
rect 12210 2385 12262 2437
rect 12275 2385 12327 2437
rect 11440 2317 11492 2369
rect 11504 2317 11556 2369
rect 11568 2317 11620 2369
rect 11632 2317 11684 2369
rect 11696 2317 11748 2369
rect 11760 2317 11812 2369
rect 11824 2317 11876 2369
rect 11888 2317 11940 2369
rect 11952 2317 12004 2369
rect 12016 2317 12068 2369
rect 12080 2317 12132 2369
rect 12145 2317 12197 2369
rect 12210 2317 12262 2369
rect 12275 2317 12327 2369
rect 11440 2249 11492 2301
rect 11504 2249 11556 2301
rect 11568 2249 11620 2301
rect 11632 2249 11684 2301
rect 11696 2249 11748 2301
rect 11760 2249 11812 2301
rect 11824 2249 11876 2301
rect 11888 2249 11940 2301
rect 11952 2249 12004 2301
rect 12016 2249 12068 2301
rect 12080 2249 12132 2301
rect 12145 2249 12197 2301
rect 12210 2249 12262 2301
rect 12275 2249 12327 2301
rect 11440 2181 11492 2233
rect 11504 2181 11556 2233
rect 11568 2181 11620 2233
rect 11632 2181 11684 2233
rect 11696 2181 11748 2233
rect 11760 2181 11812 2233
rect 11824 2181 11876 2233
rect 11888 2181 11940 2233
rect 11952 2181 12004 2233
rect 12016 2181 12068 2233
rect 12080 2181 12132 2233
rect 12145 2181 12197 2233
rect 12210 2181 12262 2233
rect 12275 2181 12327 2233
rect 11440 2113 11492 2165
rect 11504 2113 11556 2165
rect 11568 2113 11620 2165
rect 11632 2113 11684 2165
rect 11696 2113 11748 2165
rect 11760 2113 11812 2165
rect 11824 2113 11876 2165
rect 11888 2113 11940 2165
rect 11952 2113 12004 2165
rect 12016 2113 12068 2165
rect 12080 2113 12132 2165
rect 12145 2113 12197 2165
rect 12210 2113 12262 2165
rect 12275 2113 12327 2165
rect 11440 2045 11492 2097
rect 11504 2045 11556 2097
rect 11568 2045 11620 2097
rect 11632 2045 11684 2097
rect 11696 2045 11748 2097
rect 11760 2045 11812 2097
rect 11824 2045 11876 2097
rect 11888 2045 11940 2097
rect 11952 2045 12004 2097
rect 12016 2045 12068 2097
rect 12080 2045 12132 2097
rect 12145 2045 12197 2097
rect 12210 2045 12262 2097
rect 12275 2045 12327 2097
rect 13995 2385 14047 2437
rect 14060 2385 14112 2437
rect 14125 2385 14177 2437
rect 14190 2385 14242 2437
rect 14254 2385 14306 2437
rect 14318 2385 14370 2437
rect 14382 2385 14434 2437
rect 14446 2385 14498 2437
rect 14510 2385 14562 2437
rect 14574 2385 14626 2437
rect 14638 2385 14690 2437
rect 14702 2385 14754 2437
rect 14766 2385 14818 2437
rect 14830 2385 14882 2437
rect 13995 2317 14047 2369
rect 14060 2317 14112 2369
rect 14125 2317 14177 2369
rect 14190 2317 14242 2369
rect 14254 2317 14306 2369
rect 14318 2317 14370 2369
rect 14382 2317 14434 2369
rect 14446 2317 14498 2369
rect 14510 2317 14562 2369
rect 14574 2317 14626 2369
rect 14638 2317 14690 2369
rect 14702 2317 14754 2369
rect 14766 2317 14818 2369
rect 14830 2317 14882 2369
rect 13995 2249 14047 2301
rect 14060 2249 14112 2301
rect 14125 2249 14177 2301
rect 14190 2249 14242 2301
rect 14254 2249 14306 2301
rect 14318 2249 14370 2301
rect 14382 2249 14434 2301
rect 14446 2249 14498 2301
rect 14510 2249 14562 2301
rect 14574 2249 14626 2301
rect 14638 2249 14690 2301
rect 14702 2249 14754 2301
rect 14766 2249 14818 2301
rect 14830 2249 14882 2301
rect 13995 2181 14047 2233
rect 14060 2181 14112 2233
rect 14125 2181 14177 2233
rect 14190 2181 14242 2233
rect 14254 2181 14306 2233
rect 14318 2181 14370 2233
rect 14382 2181 14434 2233
rect 14446 2181 14498 2233
rect 14510 2181 14562 2233
rect 14574 2181 14626 2233
rect 14638 2181 14690 2233
rect 14702 2181 14754 2233
rect 14766 2181 14818 2233
rect 14830 2181 14882 2233
rect 13995 2113 14047 2165
rect 14060 2113 14112 2165
rect 14125 2113 14177 2165
rect 14190 2113 14242 2165
rect 14254 2113 14306 2165
rect 14318 2113 14370 2165
rect 14382 2113 14434 2165
rect 14446 2113 14498 2165
rect 14510 2113 14562 2165
rect 14574 2113 14626 2165
rect 14638 2113 14690 2165
rect 14702 2113 14754 2165
rect 14766 2113 14818 2165
rect 14830 2113 14882 2165
rect 13995 2045 14047 2097
rect 14060 2045 14112 2097
rect 14125 2045 14177 2097
rect 14190 2045 14242 2097
rect 14254 2045 14306 2097
rect 14318 2045 14370 2097
rect 14382 2045 14434 2097
rect 14446 2045 14498 2097
rect 14510 2045 14562 2097
rect 14574 2045 14626 2097
rect 14638 2045 14690 2097
rect 14702 2045 14754 2097
rect 14766 2045 14818 2097
rect 14830 2045 14882 2097
rect 17924 2385 17976 2437
rect 17988 2385 18040 2437
rect 18052 2385 18104 2437
rect 18116 2385 18168 2437
rect 18180 2385 18232 2437
rect 18244 2385 18296 2437
rect 18308 2385 18360 2437
rect 18372 2385 18424 2437
rect 18436 2385 18488 2437
rect 18500 2385 18552 2437
rect 18564 2385 18616 2437
rect 18629 2385 18681 2437
rect 18694 2385 18746 2437
rect 18759 2385 18811 2437
rect 17924 2317 17976 2369
rect 17988 2317 18040 2369
rect 18052 2317 18104 2369
rect 18116 2317 18168 2369
rect 18180 2317 18232 2369
rect 18244 2317 18296 2369
rect 18308 2317 18360 2369
rect 18372 2317 18424 2369
rect 18436 2317 18488 2369
rect 18500 2317 18552 2369
rect 18564 2317 18616 2369
rect 18629 2317 18681 2369
rect 18694 2317 18746 2369
rect 18759 2317 18811 2369
rect 17924 2249 17976 2301
rect 17988 2249 18040 2301
rect 18052 2249 18104 2301
rect 18116 2249 18168 2301
rect 18180 2249 18232 2301
rect 18244 2249 18296 2301
rect 18308 2249 18360 2301
rect 18372 2249 18424 2301
rect 18436 2249 18488 2301
rect 18500 2249 18552 2301
rect 18564 2249 18616 2301
rect 18629 2249 18681 2301
rect 18694 2249 18746 2301
rect 18759 2249 18811 2301
rect 17924 2181 17976 2233
rect 17988 2181 18040 2233
rect 18052 2181 18104 2233
rect 18116 2181 18168 2233
rect 18180 2181 18232 2233
rect 18244 2181 18296 2233
rect 18308 2181 18360 2233
rect 18372 2181 18424 2233
rect 18436 2181 18488 2233
rect 18500 2181 18552 2233
rect 18564 2181 18616 2233
rect 18629 2181 18681 2233
rect 18694 2181 18746 2233
rect 18759 2181 18811 2233
rect 17924 2113 17976 2165
rect 17988 2113 18040 2165
rect 18052 2113 18104 2165
rect 18116 2113 18168 2165
rect 18180 2113 18232 2165
rect 18244 2113 18296 2165
rect 18308 2113 18360 2165
rect 18372 2113 18424 2165
rect 18436 2113 18488 2165
rect 18500 2113 18552 2165
rect 18564 2113 18616 2165
rect 18629 2113 18681 2165
rect 18694 2113 18746 2165
rect 18759 2113 18811 2165
rect 17924 2045 17976 2097
rect 17988 2045 18040 2097
rect 18052 2045 18104 2097
rect 18116 2045 18168 2097
rect 18180 2045 18232 2097
rect 18244 2045 18296 2097
rect 18308 2045 18360 2097
rect 18372 2045 18424 2097
rect 18436 2045 18488 2097
rect 18500 2045 18552 2097
rect 18564 2045 18616 2097
rect 18629 2045 18681 2097
rect 18694 2045 18746 2097
rect 18759 2045 18811 2097
rect -1636 1913 -1584 1922
rect -1636 1882 -1584 1894
rect -1736 1797 -1684 1849
rect -1636 1848 -1607 1882
rect -1607 1848 -1584 1882
rect -1636 1842 -1584 1848
rect -1736 1733 -1684 1785
rect -630 1755 -578 1807
rect -630 1691 -578 1743
rect 644 1867 696 1919
rect 728 1867 780 1919
rect 812 1867 864 1919
rect 895 1867 947 1919
rect 6018 1867 6070 1919
rect 6085 1867 6137 1919
rect 6152 1867 6204 1919
rect 6219 1867 6271 1919
rect 6286 1867 6338 1919
rect 6353 1867 6405 1919
rect 6949 1867 7001 1919
rect 7016 1867 7068 1919
rect 7083 1867 7135 1919
rect 7150 1867 7202 1919
rect 7217 1867 7269 1919
rect 7284 1867 7336 1919
rect 12502 1867 12554 1919
rect 12569 1867 12621 1919
rect 12636 1867 12688 1919
rect 12703 1867 12755 1919
rect 12770 1867 12822 1919
rect 12837 1867 12889 1919
rect 644 1803 696 1855
rect 728 1803 780 1855
rect 812 1803 864 1855
rect 895 1803 947 1855
rect 6018 1803 6070 1855
rect 6085 1803 6137 1855
rect 6152 1803 6204 1855
rect 6219 1803 6271 1855
rect 6286 1803 6338 1855
rect 6353 1803 6405 1855
rect 6949 1803 7001 1855
rect 7016 1803 7068 1855
rect 7083 1803 7135 1855
rect 7150 1803 7202 1855
rect 7217 1803 7269 1855
rect 7284 1803 7336 1855
rect 12502 1803 12554 1855
rect 12569 1803 12621 1855
rect 12636 1803 12688 1855
rect 12703 1803 12755 1855
rect 12770 1803 12822 1855
rect 12837 1803 12889 1855
rect 644 1739 696 1791
rect 728 1739 780 1791
rect 812 1739 864 1791
rect 895 1739 947 1791
rect 6018 1739 6070 1791
rect 6085 1739 6137 1791
rect 6152 1739 6204 1791
rect 6219 1739 6271 1791
rect 6286 1739 6338 1791
rect 6353 1739 6405 1791
rect 6949 1739 7001 1791
rect 7016 1739 7068 1791
rect 7083 1739 7135 1791
rect 7150 1739 7202 1791
rect 7217 1739 7269 1791
rect 7284 1739 7336 1791
rect 12502 1739 12554 1791
rect 12569 1739 12621 1791
rect 12636 1739 12688 1791
rect 12703 1739 12755 1791
rect 12770 1739 12822 1791
rect 12837 1739 12889 1791
rect 13433 1867 13485 1919
rect 13500 1867 13552 1919
rect 13567 1867 13619 1919
rect 13634 1867 13686 1919
rect 13701 1867 13753 1919
rect 13768 1867 13820 1919
rect 13433 1803 13485 1855
rect 13500 1803 13552 1855
rect 13567 1803 13619 1855
rect 13634 1803 13686 1855
rect 13701 1803 13753 1855
rect 13768 1803 13820 1855
rect 13433 1739 13485 1791
rect 13500 1739 13552 1791
rect 13567 1739 13619 1791
rect 13634 1739 13686 1791
rect 13701 1739 13753 1791
rect 13768 1739 13820 1791
rect 19071 1867 19123 1919
rect 19154 1867 19206 1919
rect 19237 1867 19289 1919
rect 19321 1867 19373 1919
rect 19071 1803 19123 1855
rect 19154 1803 19206 1855
rect 19237 1803 19289 1855
rect 19321 1803 19373 1855
rect 19071 1739 19123 1791
rect 19154 1739 19206 1791
rect 19237 1739 19289 1791
rect 19321 1739 19373 1791
rect -630 1451 -578 1503
rect -132 1480 -80 1532
rect -630 1387 -578 1439
rect -132 1416 -80 1468
rect 2677 1640 2729 1685
rect 2744 1640 2796 1685
rect 2811 1640 2863 1685
rect 2878 1640 2930 1685
rect 2945 1640 2997 1685
rect 3012 1640 3064 1685
rect 2677 1633 2712 1640
rect 2712 1633 2729 1640
rect 2744 1633 2746 1640
rect 2746 1633 2786 1640
rect 2786 1633 2796 1640
rect 2811 1633 2820 1640
rect 2820 1633 2860 1640
rect 2860 1633 2863 1640
rect 2878 1633 2894 1640
rect 2894 1633 2930 1640
rect 2945 1633 2968 1640
rect 2968 1633 2997 1640
rect 3012 1633 3042 1640
rect 3042 1633 3064 1640
rect 3079 1640 3131 1685
rect 3079 1633 3082 1640
rect 3082 1633 3116 1640
rect 3116 1633 3131 1640
rect 3146 1640 3198 1685
rect 3146 1633 3156 1640
rect 3156 1633 3190 1640
rect 3190 1633 3198 1640
rect 3213 1640 3265 1685
rect 3213 1633 3230 1640
rect 3230 1633 3264 1640
rect 3264 1633 3265 1640
rect 3279 1633 3331 1685
rect 3345 1633 3397 1685
rect 3411 1633 3463 1685
rect 3477 1633 3529 1685
rect 3543 1633 3595 1685
rect 4882 1640 4934 1685
rect 4971 1640 5023 1685
rect 5059 1640 5111 1685
rect 5720 1640 5772 1685
rect 5799 1640 5851 1685
rect 2677 1606 2712 1613
rect 2712 1606 2729 1613
rect 2744 1606 2746 1613
rect 2746 1606 2786 1613
rect 2786 1606 2796 1613
rect 2811 1606 2820 1613
rect 2820 1606 2860 1613
rect 2860 1606 2863 1613
rect 2878 1606 2894 1613
rect 2894 1606 2930 1613
rect 2945 1606 2968 1613
rect 2968 1606 2997 1613
rect 3012 1606 3042 1613
rect 3042 1606 3064 1613
rect 2677 1568 2729 1606
rect 2744 1568 2796 1606
rect 2811 1568 2863 1606
rect 2878 1568 2930 1606
rect 2945 1568 2997 1606
rect 3012 1568 3064 1606
rect 2677 1561 2712 1568
rect 2712 1561 2729 1568
rect 2744 1561 2746 1568
rect 2746 1561 2786 1568
rect 2786 1561 2796 1568
rect 2811 1561 2820 1568
rect 2820 1561 2860 1568
rect 2860 1561 2863 1568
rect 2878 1561 2894 1568
rect 2894 1561 2930 1568
rect 2945 1561 2968 1568
rect 2968 1561 2997 1568
rect 3012 1561 3042 1568
rect 3042 1561 3064 1568
rect 3079 1606 3082 1613
rect 3082 1606 3116 1613
rect 3116 1606 3131 1613
rect 3079 1568 3131 1606
rect 3079 1561 3082 1568
rect 3082 1561 3116 1568
rect 3116 1561 3131 1568
rect 3146 1606 3156 1613
rect 3156 1606 3190 1613
rect 3190 1606 3198 1613
rect 3146 1568 3198 1606
rect 3146 1561 3156 1568
rect 3156 1561 3190 1568
rect 3190 1561 3198 1568
rect 3213 1606 3230 1613
rect 3230 1606 3264 1613
rect 3264 1606 3265 1613
rect 3213 1568 3265 1606
rect 3213 1561 3230 1568
rect 3230 1561 3264 1568
rect 3264 1561 3265 1568
rect 3279 1561 3331 1613
rect 3345 1561 3397 1613
rect 3411 1561 3463 1613
rect 3477 1561 3529 1613
rect 3543 1561 3595 1613
rect 4882 1633 4898 1640
rect 4898 1633 4934 1640
rect 4971 1633 4972 1640
rect 4972 1633 5012 1640
rect 5012 1633 5023 1640
rect 5059 1633 5085 1640
rect 5085 1633 5111 1640
rect 4882 1606 4898 1613
rect 4898 1606 4934 1613
rect 4971 1606 4972 1613
rect 4972 1606 5012 1613
rect 5012 1606 5023 1613
rect 5059 1606 5085 1613
rect 5085 1606 5111 1613
rect 5720 1633 5742 1640
rect 5742 1633 5772 1640
rect 5799 1633 5815 1640
rect 5815 1633 5849 1640
rect 5849 1633 5851 1640
rect 5878 1640 5930 1685
rect 6497 1640 6549 1685
rect 5878 1633 5888 1640
rect 5888 1633 5922 1640
rect 5922 1633 5930 1640
rect 5720 1606 5742 1613
rect 5742 1606 5772 1613
rect 5799 1606 5815 1613
rect 5815 1606 5849 1613
rect 5849 1606 5851 1613
rect 4882 1568 4934 1606
rect 4971 1568 5023 1606
rect 5059 1568 5111 1606
rect 5720 1568 5772 1606
rect 5799 1568 5851 1606
rect 2677 1534 2712 1541
rect 2712 1534 2729 1541
rect 2744 1534 2746 1541
rect 2746 1534 2786 1541
rect 2786 1534 2796 1541
rect 2811 1534 2820 1541
rect 2820 1534 2860 1541
rect 2860 1534 2863 1541
rect 2878 1534 2894 1541
rect 2894 1534 2930 1541
rect 2945 1534 2968 1541
rect 2968 1534 2997 1541
rect 3012 1534 3042 1541
rect 3042 1534 3064 1541
rect 2677 1489 2729 1534
rect 2744 1489 2796 1534
rect 2811 1489 2863 1534
rect 2878 1489 2930 1534
rect 2945 1489 2997 1534
rect 3012 1489 3064 1534
rect 3079 1534 3082 1541
rect 3082 1534 3116 1541
rect 3116 1534 3131 1541
rect 3079 1489 3131 1534
rect 3146 1534 3156 1541
rect 3156 1534 3190 1541
rect 3190 1534 3198 1541
rect 3146 1489 3198 1534
rect 3213 1534 3230 1541
rect 3230 1534 3264 1541
rect 3264 1534 3265 1541
rect 3213 1489 3265 1534
rect 3279 1489 3331 1541
rect 3345 1489 3397 1541
rect 3411 1489 3463 1541
rect 3477 1489 3529 1541
rect 3543 1489 3595 1541
rect 4882 1561 4898 1568
rect 4898 1561 4934 1568
rect 4971 1561 4972 1568
rect 4972 1561 5012 1568
rect 5012 1561 5023 1568
rect 5059 1561 5085 1568
rect 5085 1561 5111 1568
rect 4882 1534 4898 1541
rect 4898 1534 4934 1541
rect 4971 1534 4972 1541
rect 4972 1534 5012 1541
rect 5012 1534 5023 1541
rect 5059 1534 5085 1541
rect 5085 1534 5111 1541
rect 5720 1561 5742 1568
rect 5742 1561 5772 1568
rect 5799 1561 5815 1568
rect 5815 1561 5849 1568
rect 5849 1561 5851 1568
rect 5878 1606 5888 1613
rect 5888 1606 5922 1613
rect 5922 1606 5930 1613
rect 6497 1633 6506 1640
rect 6506 1633 6549 1640
rect 6574 1633 6626 1685
rect 6651 1633 6703 1685
rect 6728 1633 6780 1685
rect 6805 1640 6857 1685
rect 9525 1640 9577 1685
rect 9592 1640 9644 1685
rect 9659 1640 9711 1685
rect 9726 1640 9778 1685
rect 6805 1633 6848 1640
rect 6848 1633 6857 1640
rect 6497 1606 6506 1613
rect 6506 1606 6549 1613
rect 5878 1568 5930 1606
rect 6497 1568 6549 1606
rect 5878 1561 5888 1568
rect 5888 1561 5922 1568
rect 5922 1561 5930 1568
rect 5720 1534 5742 1541
rect 5742 1534 5772 1541
rect 5799 1534 5815 1541
rect 5815 1534 5849 1541
rect 5849 1534 5851 1541
rect 4882 1489 4934 1534
rect 4971 1489 5023 1534
rect 5059 1489 5111 1534
rect 5720 1489 5772 1534
rect 5799 1489 5851 1534
rect 5878 1534 5888 1541
rect 5888 1534 5922 1541
rect 5922 1534 5930 1541
rect 6497 1561 6506 1568
rect 6506 1561 6549 1568
rect 6574 1561 6626 1613
rect 6651 1561 6703 1613
rect 6728 1561 6780 1613
rect 6805 1606 6848 1613
rect 6848 1606 6857 1613
rect 9525 1633 9526 1640
rect 9526 1633 9566 1640
rect 9566 1633 9577 1640
rect 9592 1633 9600 1640
rect 9600 1633 9640 1640
rect 9640 1633 9644 1640
rect 9659 1633 9674 1640
rect 9674 1633 9711 1640
rect 9726 1633 9748 1640
rect 9748 1633 9778 1640
rect 9525 1606 9526 1613
rect 9526 1606 9566 1613
rect 9566 1606 9577 1613
rect 9592 1606 9600 1613
rect 9600 1606 9640 1613
rect 9640 1606 9644 1613
rect 9659 1606 9674 1613
rect 9674 1606 9711 1613
rect 9726 1606 9748 1613
rect 9748 1606 9778 1613
rect 16403 1633 16455 1685
rect 16471 1633 16523 1685
rect 16539 1640 16591 1685
rect 16607 1640 16659 1685
rect 16674 1640 16726 1685
rect 16741 1640 16793 1685
rect 16539 1633 16574 1640
rect 16574 1633 16591 1640
rect 16607 1633 16608 1640
rect 16608 1633 16648 1640
rect 16648 1633 16659 1640
rect 16674 1633 16682 1640
rect 16682 1633 16722 1640
rect 16722 1633 16726 1640
rect 16741 1633 16756 1640
rect 16756 1633 16793 1640
rect 6805 1568 6857 1606
rect 9525 1568 9577 1606
rect 9592 1568 9644 1606
rect 9659 1568 9711 1606
rect 9726 1568 9778 1606
rect 6805 1561 6848 1568
rect 6848 1561 6857 1568
rect 6497 1534 6506 1541
rect 6506 1534 6549 1541
rect 5878 1489 5930 1534
rect 6497 1489 6549 1534
rect 6574 1489 6626 1541
rect 6651 1489 6703 1541
rect 6728 1489 6780 1541
rect 6805 1534 6848 1541
rect 6848 1534 6857 1541
rect 9525 1561 9526 1568
rect 9526 1561 9566 1568
rect 9566 1561 9577 1568
rect 9592 1561 9600 1568
rect 9600 1561 9640 1568
rect 9640 1561 9644 1568
rect 9659 1561 9674 1568
rect 9674 1561 9711 1568
rect 9726 1561 9748 1568
rect 9748 1561 9778 1568
rect 9525 1534 9526 1541
rect 9526 1534 9566 1541
rect 9566 1534 9577 1541
rect 9592 1534 9600 1541
rect 9600 1534 9640 1541
rect 9640 1534 9644 1541
rect 9659 1534 9674 1541
rect 9674 1534 9711 1541
rect 9726 1534 9748 1541
rect 9748 1534 9778 1541
rect 16403 1561 16455 1613
rect 16471 1561 16523 1613
rect 16539 1606 16574 1613
rect 16574 1606 16591 1613
rect 16607 1606 16608 1613
rect 16608 1606 16648 1613
rect 16648 1606 16659 1613
rect 16674 1606 16682 1613
rect 16682 1606 16722 1613
rect 16722 1606 16726 1613
rect 16741 1606 16756 1613
rect 16756 1606 16793 1613
rect 16539 1568 16591 1606
rect 16607 1568 16659 1606
rect 16674 1568 16726 1606
rect 16741 1568 16793 1606
rect 16539 1561 16574 1568
rect 16574 1561 16591 1568
rect 16607 1561 16608 1568
rect 16608 1561 16648 1568
rect 16648 1561 16659 1568
rect 16674 1561 16682 1568
rect 16682 1561 16722 1568
rect 16722 1561 16726 1568
rect 16741 1561 16756 1568
rect 16756 1561 16793 1568
rect 6805 1489 6857 1534
rect 9525 1489 9577 1534
rect 9592 1489 9644 1534
rect 9659 1489 9711 1534
rect 9726 1489 9778 1534
rect 3376 1446 3428 1455
rect 176 1412 202 1439
rect 202 1412 228 1439
rect 3376 1412 3386 1446
rect 3386 1412 3420 1446
rect 3420 1412 3428 1446
rect 176 1387 228 1412
rect 3376 1403 3428 1412
rect 3440 1446 3492 1455
rect 3440 1412 3458 1446
rect 3458 1412 3492 1446
rect 3440 1403 3492 1412
rect 9897 1446 9949 1490
rect 16403 1489 16455 1541
rect 16471 1489 16523 1541
rect 16539 1534 16574 1541
rect 16574 1534 16591 1541
rect 16607 1534 16608 1541
rect 16608 1534 16648 1541
rect 16648 1534 16659 1541
rect 16674 1534 16682 1541
rect 16682 1534 16722 1541
rect 16722 1534 16726 1541
rect 16741 1534 16756 1541
rect 16756 1534 16793 1541
rect 16539 1489 16591 1534
rect 16607 1489 16659 1534
rect 16674 1489 16726 1534
rect 16741 1489 16793 1534
rect 9897 1438 9904 1446
rect 9904 1438 9942 1446
rect 9942 1438 9949 1446
rect 9897 1412 9904 1426
rect 9904 1412 9942 1426
rect 9942 1412 9949 1426
rect 176 1323 228 1375
rect 1027 1319 1079 1371
rect 1092 1319 1144 1371
rect 1157 1319 1209 1371
rect 1222 1319 1274 1371
rect 1286 1319 1338 1371
rect 1350 1319 1402 1371
rect 1414 1319 1466 1371
rect 1478 1319 1530 1371
rect 1542 1319 1594 1371
rect 1606 1319 1658 1371
rect 1670 1319 1722 1371
rect 1734 1319 1786 1371
rect 1798 1319 1850 1371
rect 1862 1319 1914 1371
rect 5199 1319 5251 1371
rect 5263 1319 5315 1371
rect 5327 1319 5379 1371
rect 5392 1319 5444 1371
rect 5457 1319 5509 1371
rect 5522 1319 5574 1371
rect 5587 1319 5639 1371
rect 7511 1319 7563 1371
rect 7576 1319 7628 1371
rect 7641 1319 7693 1371
rect 7706 1319 7758 1371
rect 7770 1319 7822 1371
rect 7834 1319 7886 1371
rect 7898 1319 7950 1371
rect 7962 1319 8014 1371
rect 8026 1319 8078 1371
rect 8090 1319 8142 1371
rect 8154 1319 8206 1371
rect 8218 1319 8270 1371
rect 8282 1319 8334 1371
rect 8346 1319 8398 1371
rect 9897 1374 9949 1412
rect 11440 1319 11492 1371
rect 11504 1319 11556 1371
rect 11568 1319 11620 1371
rect 11632 1319 11684 1371
rect 11696 1319 11748 1371
rect 11760 1319 11812 1371
rect 11824 1319 11876 1371
rect 11888 1319 11940 1371
rect 11952 1319 12004 1371
rect 12016 1319 12068 1371
rect 12080 1319 12132 1371
rect 12145 1319 12197 1371
rect 12210 1319 12262 1371
rect 12275 1319 12327 1371
rect 13995 1319 14047 1371
rect 14060 1319 14112 1371
rect 14125 1319 14177 1371
rect 14190 1319 14242 1371
rect 14254 1319 14306 1371
rect 14318 1319 14370 1371
rect 14382 1319 14434 1371
rect 14446 1319 14498 1371
rect 14510 1319 14562 1371
rect 14574 1319 14626 1371
rect 14638 1319 14690 1371
rect 14702 1319 14754 1371
rect 14766 1319 14818 1371
rect 14830 1319 14882 1371
rect 17924 1319 17976 1371
rect 17988 1319 18040 1371
rect 18052 1319 18104 1371
rect 18116 1319 18168 1371
rect 18180 1319 18232 1371
rect 18244 1319 18296 1371
rect 18308 1319 18360 1371
rect 18372 1319 18424 1371
rect 18436 1319 18488 1371
rect 18500 1319 18552 1371
rect 18564 1319 18616 1371
rect 18629 1319 18681 1371
rect 18694 1319 18746 1371
rect 18759 1319 18811 1371
rect 19610 1344 19662 1396
rect 1027 1251 1079 1303
rect 1092 1251 1144 1303
rect 1157 1251 1209 1303
rect 1222 1251 1274 1303
rect 1286 1251 1338 1303
rect 1350 1251 1402 1303
rect 1414 1251 1466 1303
rect 1478 1251 1530 1303
rect 1542 1251 1594 1303
rect 1606 1251 1658 1303
rect 1670 1251 1722 1303
rect 1734 1251 1786 1303
rect 1798 1251 1850 1303
rect 1862 1251 1914 1303
rect 5199 1251 5251 1303
rect 5263 1251 5315 1303
rect 5327 1251 5379 1303
rect 5392 1251 5444 1303
rect 5457 1251 5509 1303
rect 5522 1251 5574 1303
rect 5587 1251 5639 1303
rect 7511 1251 7563 1303
rect 7576 1251 7628 1303
rect 7641 1251 7693 1303
rect 7706 1251 7758 1303
rect 7770 1251 7822 1303
rect 7834 1251 7886 1303
rect 7898 1251 7950 1303
rect 7962 1251 8014 1303
rect 8026 1251 8078 1303
rect 8090 1251 8142 1303
rect 8154 1251 8206 1303
rect 8218 1251 8270 1303
rect 8282 1251 8334 1303
rect 8346 1251 8398 1303
rect 11440 1251 11492 1303
rect 11504 1251 11556 1303
rect 11568 1251 11620 1303
rect 11632 1251 11684 1303
rect 11696 1251 11748 1303
rect 11760 1251 11812 1303
rect 11824 1251 11876 1303
rect 11888 1251 11940 1303
rect 11952 1251 12004 1303
rect 12016 1251 12068 1303
rect 12080 1251 12132 1303
rect 12145 1251 12197 1303
rect 12210 1251 12262 1303
rect 12275 1251 12327 1303
rect 13995 1251 14047 1303
rect 14060 1251 14112 1303
rect 14125 1251 14177 1303
rect 14190 1251 14242 1303
rect 14254 1251 14306 1303
rect 14318 1251 14370 1303
rect 14382 1251 14434 1303
rect 14446 1251 14498 1303
rect 14510 1251 14562 1303
rect 14574 1251 14626 1303
rect 14638 1251 14690 1303
rect 14702 1251 14754 1303
rect 14766 1251 14818 1303
rect 14830 1251 14882 1303
rect 17924 1251 17976 1303
rect 17988 1251 18040 1303
rect 18052 1251 18104 1303
rect 18116 1251 18168 1303
rect 18180 1251 18232 1303
rect 18244 1251 18296 1303
rect 18308 1251 18360 1303
rect 18372 1251 18424 1303
rect 18436 1251 18488 1303
rect 18500 1251 18552 1303
rect 18564 1251 18616 1303
rect 18629 1251 18681 1303
rect 18694 1251 18746 1303
rect 18759 1251 18811 1303
rect 19610 1280 19662 1332
rect 1027 1228 1079 1235
rect 1027 1194 1055 1228
rect 1055 1194 1079 1228
rect 1027 1183 1079 1194
rect 1092 1228 1144 1235
rect 1092 1194 1094 1228
rect 1094 1194 1128 1228
rect 1128 1194 1144 1228
rect 1092 1183 1144 1194
rect 1157 1228 1209 1235
rect 1157 1194 1167 1228
rect 1167 1194 1201 1228
rect 1201 1194 1209 1228
rect 1157 1183 1209 1194
rect 1222 1228 1274 1235
rect 1222 1194 1240 1228
rect 1240 1194 1274 1228
rect 1222 1183 1274 1194
rect 1286 1228 1338 1235
rect 1350 1228 1402 1235
rect 1414 1228 1466 1235
rect 1478 1228 1530 1235
rect 1542 1228 1594 1235
rect 1606 1228 1658 1235
rect 1286 1194 1313 1228
rect 1313 1194 1338 1228
rect 1350 1194 1386 1228
rect 1386 1194 1402 1228
rect 1414 1194 1420 1228
rect 1420 1194 1459 1228
rect 1459 1194 1466 1228
rect 1478 1194 1493 1228
rect 1493 1194 1530 1228
rect 1542 1194 1566 1228
rect 1566 1194 1594 1228
rect 1606 1194 1639 1228
rect 1639 1194 1658 1228
rect 1286 1183 1338 1194
rect 1350 1183 1402 1194
rect 1414 1183 1466 1194
rect 1478 1183 1530 1194
rect 1542 1183 1594 1194
rect 1606 1183 1658 1194
rect 1670 1228 1722 1235
rect 1670 1194 1678 1228
rect 1678 1194 1712 1228
rect 1712 1194 1722 1228
rect 1670 1183 1722 1194
rect 1734 1228 1786 1235
rect 1734 1194 1751 1228
rect 1751 1194 1785 1228
rect 1785 1194 1786 1228
rect 1734 1183 1786 1194
rect 1798 1228 1850 1235
rect 1862 1228 1914 1235
rect 5199 1228 5251 1235
rect 5263 1228 5315 1235
rect 5327 1228 5379 1235
rect 5392 1228 5444 1235
rect 5457 1228 5509 1235
rect 1798 1194 1824 1228
rect 1824 1194 1850 1228
rect 1862 1194 1898 1228
rect 1898 1194 1914 1228
rect 5199 1194 5231 1228
rect 5231 1194 5251 1228
rect 5263 1194 5265 1228
rect 5265 1194 5304 1228
rect 5304 1194 5315 1228
rect 5327 1194 5338 1228
rect 5338 1194 5377 1228
rect 5377 1194 5379 1228
rect 5392 1194 5411 1228
rect 5411 1194 5444 1228
rect 5457 1194 5484 1228
rect 5484 1194 5509 1228
rect 1798 1183 1850 1194
rect 1862 1183 1914 1194
rect 5199 1183 5251 1194
rect 5263 1183 5315 1194
rect 5327 1183 5379 1194
rect 5392 1183 5444 1194
rect 5457 1183 5509 1194
rect 5522 1228 5574 1235
rect 5522 1194 5523 1228
rect 5523 1194 5557 1228
rect 5557 1194 5574 1228
rect 5522 1183 5574 1194
rect 5587 1228 5639 1235
rect 7511 1228 7563 1235
rect 5587 1194 5596 1228
rect 5596 1194 5630 1228
rect 5630 1194 5639 1228
rect 7511 1194 7539 1228
rect 7539 1194 7563 1228
rect 5587 1183 5639 1194
rect 7511 1183 7563 1194
rect 7576 1228 7628 1235
rect 7576 1194 7578 1228
rect 7578 1194 7612 1228
rect 7612 1194 7628 1228
rect 7576 1183 7628 1194
rect 7641 1228 7693 1235
rect 7641 1194 7651 1228
rect 7651 1194 7685 1228
rect 7685 1194 7693 1228
rect 7641 1183 7693 1194
rect 7706 1228 7758 1235
rect 7706 1194 7724 1228
rect 7724 1194 7758 1228
rect 7706 1183 7758 1194
rect 7770 1228 7822 1235
rect 7834 1228 7886 1235
rect 7898 1228 7950 1235
rect 7962 1228 8014 1235
rect 8026 1228 8078 1235
rect 8090 1228 8142 1235
rect 7770 1194 7797 1228
rect 7797 1194 7822 1228
rect 7834 1194 7870 1228
rect 7870 1194 7886 1228
rect 7898 1194 7904 1228
rect 7904 1194 7943 1228
rect 7943 1194 7950 1228
rect 7962 1194 7977 1228
rect 7977 1194 8014 1228
rect 8026 1194 8050 1228
rect 8050 1194 8078 1228
rect 8090 1194 8123 1228
rect 8123 1194 8142 1228
rect 7770 1183 7822 1194
rect 7834 1183 7886 1194
rect 7898 1183 7950 1194
rect 7962 1183 8014 1194
rect 8026 1183 8078 1194
rect 8090 1183 8142 1194
rect 8154 1228 8206 1235
rect 8154 1194 8162 1228
rect 8162 1194 8196 1228
rect 8196 1194 8206 1228
rect 8154 1183 8206 1194
rect 8218 1228 8270 1235
rect 8218 1194 8235 1228
rect 8235 1194 8269 1228
rect 8269 1194 8270 1228
rect 8218 1183 8270 1194
rect 8282 1228 8334 1235
rect 8346 1228 8398 1235
rect 11440 1228 11492 1235
rect 11504 1228 11556 1235
rect 8282 1194 8308 1228
rect 8308 1194 8334 1228
rect 8346 1194 8382 1228
rect 8382 1194 8398 1228
rect 11440 1194 11456 1228
rect 11456 1194 11492 1228
rect 11504 1194 11530 1228
rect 11530 1194 11556 1228
rect 8282 1183 8334 1194
rect 8346 1183 8398 1194
rect 11440 1183 11492 1194
rect 11504 1183 11556 1194
rect 11568 1228 11620 1235
rect 11568 1194 11569 1228
rect 11569 1194 11603 1228
rect 11603 1194 11620 1228
rect 11568 1183 11620 1194
rect 11632 1228 11684 1235
rect 11632 1194 11642 1228
rect 11642 1194 11676 1228
rect 11676 1194 11684 1228
rect 11632 1183 11684 1194
rect 11696 1228 11748 1235
rect 11760 1228 11812 1235
rect 11824 1228 11876 1235
rect 11888 1228 11940 1235
rect 11952 1228 12004 1235
rect 12016 1228 12068 1235
rect 11696 1194 11715 1228
rect 11715 1194 11748 1228
rect 11760 1194 11788 1228
rect 11788 1194 11812 1228
rect 11824 1194 11861 1228
rect 11861 1194 11876 1228
rect 11888 1194 11895 1228
rect 11895 1194 11934 1228
rect 11934 1194 11940 1228
rect 11952 1194 11968 1228
rect 11968 1194 12004 1228
rect 12016 1194 12041 1228
rect 12041 1194 12068 1228
rect 11696 1183 11748 1194
rect 11760 1183 11812 1194
rect 11824 1183 11876 1194
rect 11888 1183 11940 1194
rect 11952 1183 12004 1194
rect 12016 1183 12068 1194
rect 12080 1228 12132 1235
rect 12080 1194 12114 1228
rect 12114 1194 12132 1228
rect 12080 1183 12132 1194
rect 12145 1228 12197 1235
rect 12145 1194 12153 1228
rect 12153 1194 12187 1228
rect 12187 1194 12197 1228
rect 12145 1183 12197 1194
rect 12210 1228 12262 1235
rect 12210 1194 12226 1228
rect 12226 1194 12260 1228
rect 12260 1194 12262 1228
rect 12210 1183 12262 1194
rect 12275 1228 12327 1235
rect 13995 1228 14047 1235
rect 12275 1194 12299 1228
rect 12299 1194 12327 1228
rect 13995 1194 14023 1228
rect 14023 1194 14047 1228
rect 12275 1183 12327 1194
rect 13995 1183 14047 1194
rect 14060 1228 14112 1235
rect 14060 1194 14062 1228
rect 14062 1194 14096 1228
rect 14096 1194 14112 1228
rect 14060 1183 14112 1194
rect 14125 1228 14177 1235
rect 14125 1194 14135 1228
rect 14135 1194 14169 1228
rect 14169 1194 14177 1228
rect 14125 1183 14177 1194
rect 14190 1228 14242 1235
rect 14190 1194 14208 1228
rect 14208 1194 14242 1228
rect 14190 1183 14242 1194
rect 14254 1228 14306 1235
rect 14318 1228 14370 1235
rect 14382 1228 14434 1235
rect 14446 1228 14498 1235
rect 14510 1228 14562 1235
rect 14574 1228 14626 1235
rect 14254 1194 14281 1228
rect 14281 1194 14306 1228
rect 14318 1194 14354 1228
rect 14354 1194 14370 1228
rect 14382 1194 14388 1228
rect 14388 1194 14427 1228
rect 14427 1194 14434 1228
rect 14446 1194 14461 1228
rect 14461 1194 14498 1228
rect 14510 1194 14534 1228
rect 14534 1194 14562 1228
rect 14574 1194 14607 1228
rect 14607 1194 14626 1228
rect 14254 1183 14306 1194
rect 14318 1183 14370 1194
rect 14382 1183 14434 1194
rect 14446 1183 14498 1194
rect 14510 1183 14562 1194
rect 14574 1183 14626 1194
rect 14638 1228 14690 1235
rect 14638 1194 14646 1228
rect 14646 1194 14680 1228
rect 14680 1194 14690 1228
rect 14638 1183 14690 1194
rect 14702 1228 14754 1235
rect 14702 1194 14719 1228
rect 14719 1194 14753 1228
rect 14753 1194 14754 1228
rect 14702 1183 14754 1194
rect 14766 1228 14818 1235
rect 14830 1228 14882 1235
rect 17924 1228 17976 1235
rect 17988 1228 18040 1235
rect 14766 1194 14792 1228
rect 14792 1194 14818 1228
rect 14830 1194 14866 1228
rect 14866 1194 14882 1228
rect 17924 1194 17940 1228
rect 17940 1194 17976 1228
rect 17988 1194 18014 1228
rect 18014 1194 18040 1228
rect 14766 1183 14818 1194
rect 14830 1183 14882 1194
rect 17924 1183 17976 1194
rect 17988 1183 18040 1194
rect 18052 1228 18104 1235
rect 18052 1194 18053 1228
rect 18053 1194 18087 1228
rect 18087 1194 18104 1228
rect 18052 1183 18104 1194
rect 18116 1228 18168 1235
rect 18116 1194 18126 1228
rect 18126 1194 18160 1228
rect 18160 1194 18168 1228
rect 18116 1183 18168 1194
rect 18180 1228 18232 1235
rect 18244 1228 18296 1235
rect 18308 1228 18360 1235
rect 18372 1228 18424 1235
rect 18436 1228 18488 1235
rect 18500 1228 18552 1235
rect 18180 1194 18199 1228
rect 18199 1194 18232 1228
rect 18244 1194 18272 1228
rect 18272 1194 18296 1228
rect 18308 1194 18345 1228
rect 18345 1194 18360 1228
rect 18372 1194 18379 1228
rect 18379 1194 18418 1228
rect 18418 1194 18424 1228
rect 18436 1194 18452 1228
rect 18452 1194 18488 1228
rect 18500 1194 18525 1228
rect 18525 1194 18552 1228
rect 18180 1183 18232 1194
rect 18244 1183 18296 1194
rect 18308 1183 18360 1194
rect 18372 1183 18424 1194
rect 18436 1183 18488 1194
rect 18500 1183 18552 1194
rect 18564 1228 18616 1235
rect 18564 1194 18598 1228
rect 18598 1194 18616 1228
rect 18564 1183 18616 1194
rect 18629 1228 18681 1235
rect 18629 1194 18637 1228
rect 18637 1194 18671 1228
rect 18671 1194 18681 1228
rect 18629 1183 18681 1194
rect 18694 1228 18746 1235
rect 18694 1194 18710 1228
rect 18710 1194 18744 1228
rect 18744 1194 18746 1228
rect 18694 1183 18746 1194
rect 18759 1228 18811 1235
rect 18759 1194 18783 1228
rect 18783 1194 18811 1228
rect 18759 1183 18811 1194
rect 1027 1156 1079 1167
rect 1027 1122 1055 1156
rect 1055 1122 1079 1156
rect 1027 1115 1079 1122
rect 1092 1156 1144 1167
rect 1092 1122 1094 1156
rect 1094 1122 1128 1156
rect 1128 1122 1144 1156
rect 1092 1115 1144 1122
rect 1157 1156 1209 1167
rect 1157 1122 1167 1156
rect 1167 1122 1201 1156
rect 1201 1122 1209 1156
rect 1157 1115 1209 1122
rect 1222 1156 1274 1167
rect 1222 1122 1240 1156
rect 1240 1122 1274 1156
rect 1222 1115 1274 1122
rect 1286 1156 1338 1167
rect 1350 1156 1402 1167
rect 1414 1156 1466 1167
rect 1478 1156 1530 1167
rect 1542 1156 1594 1167
rect 1606 1156 1658 1167
rect 1286 1122 1313 1156
rect 1313 1122 1338 1156
rect 1350 1122 1386 1156
rect 1386 1122 1402 1156
rect 1414 1122 1420 1156
rect 1420 1122 1459 1156
rect 1459 1122 1466 1156
rect 1478 1122 1493 1156
rect 1493 1122 1530 1156
rect 1542 1122 1566 1156
rect 1566 1122 1594 1156
rect 1606 1122 1639 1156
rect 1639 1122 1658 1156
rect 1286 1115 1338 1122
rect 1350 1115 1402 1122
rect 1414 1115 1466 1122
rect 1478 1115 1530 1122
rect 1542 1115 1594 1122
rect 1606 1115 1658 1122
rect 1670 1156 1722 1167
rect 1670 1122 1678 1156
rect 1678 1122 1712 1156
rect 1712 1122 1722 1156
rect 1670 1115 1722 1122
rect 1734 1156 1786 1167
rect 1734 1122 1751 1156
rect 1751 1122 1785 1156
rect 1785 1122 1786 1156
rect 1734 1115 1786 1122
rect 1798 1156 1850 1167
rect 1862 1156 1914 1167
rect 5199 1156 5251 1167
rect 5263 1156 5315 1167
rect 5327 1156 5379 1167
rect 5392 1156 5444 1167
rect 5457 1156 5509 1167
rect 1798 1122 1824 1156
rect 1824 1122 1850 1156
rect 1862 1122 1898 1156
rect 1898 1122 1914 1156
rect 5199 1122 5231 1156
rect 5231 1122 5251 1156
rect 5263 1122 5265 1156
rect 5265 1122 5304 1156
rect 5304 1122 5315 1156
rect 5327 1122 5338 1156
rect 5338 1122 5377 1156
rect 5377 1122 5379 1156
rect 5392 1122 5411 1156
rect 5411 1122 5444 1156
rect 5457 1122 5484 1156
rect 5484 1122 5509 1156
rect 1798 1115 1850 1122
rect 1862 1115 1914 1122
rect 5199 1115 5251 1122
rect 5263 1115 5315 1122
rect 5327 1115 5379 1122
rect 5392 1115 5444 1122
rect 5457 1115 5509 1122
rect 5522 1156 5574 1167
rect 5522 1122 5523 1156
rect 5523 1122 5557 1156
rect 5557 1122 5574 1156
rect 5522 1115 5574 1122
rect 5587 1156 5639 1167
rect 7511 1156 7563 1167
rect 5587 1122 5596 1156
rect 5596 1122 5630 1156
rect 5630 1122 5639 1156
rect 7511 1122 7539 1156
rect 7539 1122 7563 1156
rect 5587 1115 5639 1122
rect 7511 1115 7563 1122
rect 7576 1156 7628 1167
rect 7576 1122 7578 1156
rect 7578 1122 7612 1156
rect 7612 1122 7628 1156
rect 7576 1115 7628 1122
rect 7641 1156 7693 1167
rect 7641 1122 7651 1156
rect 7651 1122 7685 1156
rect 7685 1122 7693 1156
rect 7641 1115 7693 1122
rect 7706 1156 7758 1167
rect 7706 1122 7724 1156
rect 7724 1122 7758 1156
rect 7706 1115 7758 1122
rect 7770 1156 7822 1167
rect 7834 1156 7886 1167
rect 7898 1156 7950 1167
rect 7962 1156 8014 1167
rect 8026 1156 8078 1167
rect 8090 1156 8142 1167
rect 7770 1122 7797 1156
rect 7797 1122 7822 1156
rect 7834 1122 7870 1156
rect 7870 1122 7886 1156
rect 7898 1122 7904 1156
rect 7904 1122 7943 1156
rect 7943 1122 7950 1156
rect 7962 1122 7977 1156
rect 7977 1122 8014 1156
rect 8026 1122 8050 1156
rect 8050 1122 8078 1156
rect 8090 1122 8123 1156
rect 8123 1122 8142 1156
rect 7770 1115 7822 1122
rect 7834 1115 7886 1122
rect 7898 1115 7950 1122
rect 7962 1115 8014 1122
rect 8026 1115 8078 1122
rect 8090 1115 8142 1122
rect 8154 1156 8206 1167
rect 8154 1122 8162 1156
rect 8162 1122 8196 1156
rect 8196 1122 8206 1156
rect 8154 1115 8206 1122
rect 8218 1156 8270 1167
rect 8218 1122 8235 1156
rect 8235 1122 8269 1156
rect 8269 1122 8270 1156
rect 8218 1115 8270 1122
rect 8282 1156 8334 1167
rect 8346 1156 8398 1167
rect 11440 1156 11492 1167
rect 11504 1156 11556 1167
rect 8282 1122 8308 1156
rect 8308 1122 8334 1156
rect 8346 1122 8382 1156
rect 8382 1122 8398 1156
rect 11440 1122 11456 1156
rect 11456 1122 11492 1156
rect 11504 1122 11530 1156
rect 11530 1122 11556 1156
rect 8282 1115 8334 1122
rect 8346 1115 8398 1122
rect 11440 1115 11492 1122
rect 11504 1115 11556 1122
rect 11568 1156 11620 1167
rect 11568 1122 11569 1156
rect 11569 1122 11603 1156
rect 11603 1122 11620 1156
rect 11568 1115 11620 1122
rect 11632 1156 11684 1167
rect 11632 1122 11642 1156
rect 11642 1122 11676 1156
rect 11676 1122 11684 1156
rect 11632 1115 11684 1122
rect 11696 1156 11748 1167
rect 11760 1156 11812 1167
rect 11824 1156 11876 1167
rect 11888 1156 11940 1167
rect 11952 1156 12004 1167
rect 12016 1156 12068 1167
rect 11696 1122 11715 1156
rect 11715 1122 11748 1156
rect 11760 1122 11788 1156
rect 11788 1122 11812 1156
rect 11824 1122 11861 1156
rect 11861 1122 11876 1156
rect 11888 1122 11895 1156
rect 11895 1122 11934 1156
rect 11934 1122 11940 1156
rect 11952 1122 11968 1156
rect 11968 1122 12004 1156
rect 12016 1122 12041 1156
rect 12041 1122 12068 1156
rect 11696 1115 11748 1122
rect 11760 1115 11812 1122
rect 11824 1115 11876 1122
rect 11888 1115 11940 1122
rect 11952 1115 12004 1122
rect 12016 1115 12068 1122
rect 12080 1156 12132 1167
rect 12080 1122 12114 1156
rect 12114 1122 12132 1156
rect 12080 1115 12132 1122
rect 12145 1156 12197 1167
rect 12145 1122 12153 1156
rect 12153 1122 12187 1156
rect 12187 1122 12197 1156
rect 12145 1115 12197 1122
rect 12210 1156 12262 1167
rect 12210 1122 12226 1156
rect 12226 1122 12260 1156
rect 12260 1122 12262 1156
rect 12210 1115 12262 1122
rect 12275 1156 12327 1167
rect 13995 1156 14047 1167
rect 12275 1122 12299 1156
rect 12299 1122 12327 1156
rect 13995 1122 14023 1156
rect 14023 1122 14047 1156
rect 12275 1115 12327 1122
rect 13995 1115 14047 1122
rect 14060 1156 14112 1167
rect 14060 1122 14062 1156
rect 14062 1122 14096 1156
rect 14096 1122 14112 1156
rect 14060 1115 14112 1122
rect 14125 1156 14177 1167
rect 14125 1122 14135 1156
rect 14135 1122 14169 1156
rect 14169 1122 14177 1156
rect 14125 1115 14177 1122
rect 14190 1156 14242 1167
rect 14190 1122 14208 1156
rect 14208 1122 14242 1156
rect 14190 1115 14242 1122
rect 14254 1156 14306 1167
rect 14318 1156 14370 1167
rect 14382 1156 14434 1167
rect 14446 1156 14498 1167
rect 14510 1156 14562 1167
rect 14574 1156 14626 1167
rect 14254 1122 14281 1156
rect 14281 1122 14306 1156
rect 14318 1122 14354 1156
rect 14354 1122 14370 1156
rect 14382 1122 14388 1156
rect 14388 1122 14427 1156
rect 14427 1122 14434 1156
rect 14446 1122 14461 1156
rect 14461 1122 14498 1156
rect 14510 1122 14534 1156
rect 14534 1122 14562 1156
rect 14574 1122 14607 1156
rect 14607 1122 14626 1156
rect 14254 1115 14306 1122
rect 14318 1115 14370 1122
rect 14382 1115 14434 1122
rect 14446 1115 14498 1122
rect 14510 1115 14562 1122
rect 14574 1115 14626 1122
rect 14638 1156 14690 1167
rect 14638 1122 14646 1156
rect 14646 1122 14680 1156
rect 14680 1122 14690 1156
rect 14638 1115 14690 1122
rect 14702 1156 14754 1167
rect 14702 1122 14719 1156
rect 14719 1122 14753 1156
rect 14753 1122 14754 1156
rect 14702 1115 14754 1122
rect 14766 1156 14818 1167
rect 14830 1156 14882 1167
rect 17924 1156 17976 1167
rect 17988 1156 18040 1167
rect 14766 1122 14792 1156
rect 14792 1122 14818 1156
rect 14830 1122 14866 1156
rect 14866 1122 14882 1156
rect 17924 1122 17940 1156
rect 17940 1122 17976 1156
rect 17988 1122 18014 1156
rect 18014 1122 18040 1156
rect 14766 1115 14818 1122
rect 14830 1115 14882 1122
rect 17924 1115 17976 1122
rect 17988 1115 18040 1122
rect 18052 1156 18104 1167
rect 18052 1122 18053 1156
rect 18053 1122 18087 1156
rect 18087 1122 18104 1156
rect 18052 1115 18104 1122
rect 18116 1156 18168 1167
rect 18116 1122 18126 1156
rect 18126 1122 18160 1156
rect 18160 1122 18168 1156
rect 18116 1115 18168 1122
rect 18180 1156 18232 1167
rect 18244 1156 18296 1167
rect 18308 1156 18360 1167
rect 18372 1156 18424 1167
rect 18436 1156 18488 1167
rect 18500 1156 18552 1167
rect 18180 1122 18199 1156
rect 18199 1122 18232 1156
rect 18244 1122 18272 1156
rect 18272 1122 18296 1156
rect 18308 1122 18345 1156
rect 18345 1122 18360 1156
rect 18372 1122 18379 1156
rect 18379 1122 18418 1156
rect 18418 1122 18424 1156
rect 18436 1122 18452 1156
rect 18452 1122 18488 1156
rect 18500 1122 18525 1156
rect 18525 1122 18552 1156
rect 18180 1115 18232 1122
rect 18244 1115 18296 1122
rect 18308 1115 18360 1122
rect 18372 1115 18424 1122
rect 18436 1115 18488 1122
rect 18500 1115 18552 1122
rect 18564 1156 18616 1167
rect 18564 1122 18598 1156
rect 18598 1122 18616 1156
rect 18564 1115 18616 1122
rect 18629 1156 18681 1167
rect 18629 1122 18637 1156
rect 18637 1122 18671 1156
rect 18671 1122 18681 1156
rect 18629 1115 18681 1122
rect 18694 1156 18746 1167
rect 18694 1122 18710 1156
rect 18710 1122 18744 1156
rect 18744 1122 18746 1156
rect 18694 1115 18746 1122
rect 18759 1156 18811 1167
rect 18759 1122 18783 1156
rect 18783 1122 18811 1156
rect 18759 1115 18811 1122
rect 1027 1047 1079 1099
rect 1092 1047 1144 1099
rect 1157 1047 1209 1099
rect 1222 1047 1274 1099
rect 1286 1047 1338 1099
rect 1350 1047 1402 1099
rect 1414 1047 1466 1099
rect 1478 1047 1530 1099
rect 1542 1047 1594 1099
rect 1606 1047 1658 1099
rect 1670 1047 1722 1099
rect 1734 1047 1786 1099
rect 1798 1047 1850 1099
rect 1862 1047 1914 1099
rect 5199 1047 5251 1099
rect 5263 1047 5315 1099
rect 5327 1047 5379 1099
rect 5392 1047 5444 1099
rect 5457 1047 5509 1099
rect 5522 1047 5574 1099
rect 5587 1047 5639 1099
rect 7511 1047 7563 1099
rect 7576 1047 7628 1099
rect 7641 1047 7693 1099
rect 7706 1047 7758 1099
rect 7770 1047 7822 1099
rect 7834 1047 7886 1099
rect 7898 1047 7950 1099
rect 7962 1047 8014 1099
rect 8026 1047 8078 1099
rect 8090 1047 8142 1099
rect 8154 1047 8206 1099
rect 8218 1047 8270 1099
rect 8282 1047 8334 1099
rect 8346 1047 8398 1099
rect 11440 1047 11492 1099
rect 11504 1047 11556 1099
rect 11568 1047 11620 1099
rect 11632 1047 11684 1099
rect 11696 1047 11748 1099
rect 11760 1047 11812 1099
rect 11824 1047 11876 1099
rect 11888 1047 11940 1099
rect 11952 1047 12004 1099
rect 12016 1047 12068 1099
rect 12080 1047 12132 1099
rect 12145 1047 12197 1099
rect 12210 1047 12262 1099
rect 12275 1047 12327 1099
rect 13995 1047 14047 1099
rect 14060 1047 14112 1099
rect 14125 1047 14177 1099
rect 14190 1047 14242 1099
rect 14254 1047 14306 1099
rect 14318 1047 14370 1099
rect 14382 1047 14434 1099
rect 14446 1047 14498 1099
rect 14510 1047 14562 1099
rect 14574 1047 14626 1099
rect 14638 1047 14690 1099
rect 14702 1047 14754 1099
rect 14766 1047 14818 1099
rect 14830 1047 14882 1099
rect 17924 1047 17976 1099
rect 17988 1047 18040 1099
rect 18052 1047 18104 1099
rect 18116 1047 18168 1099
rect 18180 1047 18232 1099
rect 18244 1047 18296 1099
rect 18308 1047 18360 1099
rect 18372 1047 18424 1099
rect 18436 1047 18488 1099
rect 18500 1047 18552 1099
rect 18564 1047 18616 1099
rect 18629 1047 18681 1099
rect 18694 1047 18746 1099
rect 18759 1047 18811 1099
rect 19759 1151 19811 1203
rect 19759 1087 19811 1139
rect 176 968 228 1020
rect 1027 979 1079 1031
rect 1092 979 1144 1031
rect 1157 979 1209 1031
rect 1222 979 1274 1031
rect 1286 979 1338 1031
rect 1350 979 1402 1031
rect 1414 979 1466 1031
rect 1478 979 1530 1031
rect 1542 979 1594 1031
rect 1606 979 1658 1031
rect 1670 979 1722 1031
rect 1734 979 1786 1031
rect 1798 979 1850 1031
rect 1862 979 1914 1031
rect 5199 979 5251 1031
rect 5263 979 5315 1031
rect 5327 979 5379 1031
rect 5392 979 5444 1031
rect 5457 979 5509 1031
rect 5522 979 5574 1031
rect 5587 979 5639 1031
rect 7511 979 7563 1031
rect 7576 979 7628 1031
rect 7641 979 7693 1031
rect 7706 979 7758 1031
rect 7770 979 7822 1031
rect 7834 979 7886 1031
rect 7898 979 7950 1031
rect 7962 979 8014 1031
rect 8026 979 8078 1031
rect 8090 979 8142 1031
rect 8154 979 8206 1031
rect 8218 979 8270 1031
rect 8282 979 8334 1031
rect 8346 979 8398 1031
rect 11440 979 11492 1031
rect 11504 979 11556 1031
rect 11568 979 11620 1031
rect 11632 979 11684 1031
rect 11696 979 11748 1031
rect 11760 979 11812 1031
rect 11824 979 11876 1031
rect 11888 979 11940 1031
rect 11952 979 12004 1031
rect 12016 979 12068 1031
rect 12080 979 12132 1031
rect 12145 979 12197 1031
rect 12210 979 12262 1031
rect 12275 979 12327 1031
rect 13995 979 14047 1031
rect 14060 979 14112 1031
rect 14125 979 14177 1031
rect 14190 979 14242 1031
rect 14254 979 14306 1031
rect 14318 979 14370 1031
rect 14382 979 14434 1031
rect 14446 979 14498 1031
rect 14510 979 14562 1031
rect 14574 979 14626 1031
rect 14638 979 14690 1031
rect 14702 979 14754 1031
rect 14766 979 14818 1031
rect 14830 979 14882 1031
rect 17924 979 17976 1031
rect 17988 979 18040 1031
rect 18052 979 18104 1031
rect 18116 979 18168 1031
rect 18180 979 18232 1031
rect 18244 979 18296 1031
rect 18308 979 18360 1031
rect 18372 979 18424 1031
rect 18436 979 18488 1031
rect 18500 979 18552 1031
rect 18564 979 18616 1031
rect 18629 979 18681 1031
rect 18694 979 18746 1031
rect 18759 979 18811 1031
rect 19610 975 19662 1027
rect 176 938 228 956
rect 176 904 202 938
rect 202 904 228 938
rect 19610 938 19662 963
rect 19610 911 19622 938
rect 19622 911 19660 938
rect 19660 911 19662 938
rect -630 818 -578 870
rect -630 754 -578 806
rect -222 675 -170 727
rect -222 611 -170 663
rect 3913 816 3965 861
rect 3977 816 4029 861
rect 3913 809 3936 816
rect 3936 809 3965 816
rect 3977 809 4010 816
rect 4010 809 4029 816
rect 4041 816 4093 861
rect 4041 809 4050 816
rect 4050 809 4084 816
rect 4084 809 4093 816
rect 4105 816 4157 861
rect 4169 816 4221 861
rect 4233 816 4285 861
rect 4297 816 4349 861
rect 4361 816 4413 861
rect 4425 816 4477 861
rect 4105 809 4124 816
rect 4124 809 4157 816
rect 4169 809 4198 816
rect 4198 809 4221 816
rect 4233 809 4272 816
rect 4272 809 4285 816
rect 4297 809 4306 816
rect 4306 809 4346 816
rect 4346 809 4349 816
rect 4361 809 4380 816
rect 4380 809 4413 816
rect 4425 809 4454 816
rect 4454 809 4477 816
rect 4489 816 4541 861
rect 4489 809 4494 816
rect 4494 809 4528 816
rect 4528 809 4541 816
rect 4553 816 4605 861
rect 4553 809 4568 816
rect 4568 809 4602 816
rect 4602 809 4605 816
rect 4617 816 4669 861
rect 4681 816 4733 861
rect 4746 816 4798 861
rect 8556 816 8608 861
rect 8621 816 8673 861
rect 8685 816 8737 861
rect 4617 809 4642 816
rect 4642 809 4669 816
rect 4681 809 4716 816
rect 4716 809 4733 816
rect 4746 809 4750 816
rect 4750 809 4790 816
rect 4790 809 4798 816
rect 3913 782 3936 789
rect 3936 782 3965 789
rect 3977 782 4010 789
rect 4010 782 4029 789
rect 3913 744 3965 782
rect 3977 744 4029 782
rect 3913 737 3936 744
rect 3936 737 3965 744
rect 3977 737 4010 744
rect 4010 737 4029 744
rect 4041 782 4050 789
rect 4050 782 4084 789
rect 4084 782 4093 789
rect 4041 744 4093 782
rect 4041 737 4050 744
rect 4050 737 4084 744
rect 4084 737 4093 744
rect 4105 782 4124 789
rect 4124 782 4157 789
rect 4169 782 4198 789
rect 4198 782 4221 789
rect 4233 782 4272 789
rect 4272 782 4285 789
rect 4297 782 4306 789
rect 4306 782 4346 789
rect 4346 782 4349 789
rect 4361 782 4380 789
rect 4380 782 4413 789
rect 4425 782 4454 789
rect 4454 782 4477 789
rect 4105 744 4157 782
rect 4169 744 4221 782
rect 4233 744 4285 782
rect 4297 744 4349 782
rect 4361 744 4413 782
rect 4425 744 4477 782
rect 4105 737 4124 744
rect 4124 737 4157 744
rect 4169 737 4198 744
rect 4198 737 4221 744
rect 4233 737 4272 744
rect 4272 737 4285 744
rect 4297 737 4306 744
rect 4306 737 4346 744
rect 4346 737 4349 744
rect 4361 737 4380 744
rect 4380 737 4413 744
rect 4425 737 4454 744
rect 4454 737 4477 744
rect 4489 782 4494 789
rect 4494 782 4528 789
rect 4528 782 4541 789
rect 4489 744 4541 782
rect 4489 737 4494 744
rect 4494 737 4528 744
rect 4528 737 4541 744
rect 4553 782 4568 789
rect 4568 782 4602 789
rect 4602 782 4605 789
rect 4553 744 4605 782
rect 4553 737 4568 744
rect 4568 737 4602 744
rect 4602 737 4605 744
rect 4617 782 4642 789
rect 4642 782 4669 789
rect 4681 782 4716 789
rect 4716 782 4733 789
rect 4746 782 4750 789
rect 4750 782 4790 789
rect 4790 782 4798 789
rect 8556 809 8564 816
rect 8564 809 8604 816
rect 8604 809 8608 816
rect 8621 809 8638 816
rect 8638 809 8673 816
rect 8685 809 8712 816
rect 8712 809 8737 816
rect 8749 816 8801 861
rect 8749 809 8752 816
rect 8752 809 8786 816
rect 8786 809 8801 816
rect 8813 816 8865 861
rect 8813 809 8826 816
rect 8826 809 8860 816
rect 8860 809 8865 816
rect 8877 816 8929 861
rect 8941 816 8993 861
rect 9005 816 9057 861
rect 9069 816 9121 861
rect 9133 816 9185 861
rect 9197 816 9249 861
rect 8877 809 8900 816
rect 8900 809 8929 816
rect 8941 809 8974 816
rect 8974 809 8993 816
rect 9005 809 9008 816
rect 9008 809 9048 816
rect 9048 809 9057 816
rect 9069 809 9082 816
rect 9082 809 9121 816
rect 9133 809 9156 816
rect 9156 809 9185 816
rect 9197 809 9230 816
rect 9230 809 9249 816
rect 9261 816 9313 861
rect 9261 809 9270 816
rect 9270 809 9304 816
rect 9304 809 9313 816
rect 9325 816 9377 861
rect 9389 816 9441 861
rect 10397 816 10449 861
rect 10461 816 10513 861
rect 9325 809 9344 816
rect 9344 809 9377 816
rect 9389 809 9418 816
rect 9418 809 9441 816
rect 8556 782 8564 789
rect 8564 782 8604 789
rect 8604 782 8608 789
rect 8621 782 8638 789
rect 8638 782 8673 789
rect 8685 782 8712 789
rect 8712 782 8737 789
rect 4617 744 4669 782
rect 4681 744 4733 782
rect 4746 744 4798 782
rect 8556 744 8608 782
rect 8621 744 8673 782
rect 8685 744 8737 782
rect 4617 737 4642 744
rect 4642 737 4669 744
rect 4681 737 4716 744
rect 4716 737 4733 744
rect 4746 737 4750 744
rect 4750 737 4790 744
rect 4790 737 4798 744
rect 3913 710 3936 717
rect 3936 710 3965 717
rect 3977 710 4010 717
rect 4010 710 4029 717
rect 3913 665 3965 710
rect 3977 665 4029 710
rect 4041 710 4050 717
rect 4050 710 4084 717
rect 4084 710 4093 717
rect 4041 665 4093 710
rect 4105 710 4124 717
rect 4124 710 4157 717
rect 4169 710 4198 717
rect 4198 710 4221 717
rect 4233 710 4272 717
rect 4272 710 4285 717
rect 4297 710 4306 717
rect 4306 710 4346 717
rect 4346 710 4349 717
rect 4361 710 4380 717
rect 4380 710 4413 717
rect 4425 710 4454 717
rect 4454 710 4477 717
rect 4105 665 4157 710
rect 4169 665 4221 710
rect 4233 665 4285 710
rect 4297 665 4349 710
rect 4361 665 4413 710
rect 4425 665 4477 710
rect 4489 710 4494 717
rect 4494 710 4528 717
rect 4528 710 4541 717
rect 4489 665 4541 710
rect 4553 710 4568 717
rect 4568 710 4602 717
rect 4602 710 4605 717
rect 4553 665 4605 710
rect 4617 710 4642 717
rect 4642 710 4669 717
rect 4681 710 4716 717
rect 4716 710 4733 717
rect 4746 710 4750 717
rect 4750 710 4790 717
rect 4790 710 4798 717
rect 8556 737 8564 744
rect 8564 737 8604 744
rect 8604 737 8608 744
rect 8621 737 8638 744
rect 8638 737 8673 744
rect 8685 737 8712 744
rect 8712 737 8737 744
rect 8749 782 8752 789
rect 8752 782 8786 789
rect 8786 782 8801 789
rect 8749 744 8801 782
rect 8749 737 8752 744
rect 8752 737 8786 744
rect 8786 737 8801 744
rect 8813 782 8826 789
rect 8826 782 8860 789
rect 8860 782 8865 789
rect 8813 744 8865 782
rect 8813 737 8826 744
rect 8826 737 8860 744
rect 8860 737 8865 744
rect 8877 782 8900 789
rect 8900 782 8929 789
rect 8941 782 8974 789
rect 8974 782 8993 789
rect 9005 782 9008 789
rect 9008 782 9048 789
rect 9048 782 9057 789
rect 9069 782 9082 789
rect 9082 782 9121 789
rect 9133 782 9156 789
rect 9156 782 9185 789
rect 9197 782 9230 789
rect 9230 782 9249 789
rect 8877 744 8929 782
rect 8941 744 8993 782
rect 9005 744 9057 782
rect 9069 744 9121 782
rect 9133 744 9185 782
rect 9197 744 9249 782
rect 8877 737 8900 744
rect 8900 737 8929 744
rect 8941 737 8974 744
rect 8974 737 8993 744
rect 9005 737 9008 744
rect 9008 737 9048 744
rect 9048 737 9057 744
rect 9069 737 9082 744
rect 9082 737 9121 744
rect 9133 737 9156 744
rect 9156 737 9185 744
rect 9197 737 9230 744
rect 9230 737 9249 744
rect 9261 782 9270 789
rect 9270 782 9304 789
rect 9304 782 9313 789
rect 9261 744 9313 782
rect 9261 737 9270 744
rect 9270 737 9304 744
rect 9304 737 9313 744
rect 9325 782 9344 789
rect 9344 782 9377 789
rect 9389 782 9418 789
rect 9418 782 9441 789
rect 10397 809 10420 816
rect 10420 809 10449 816
rect 10461 809 10494 816
rect 10494 809 10513 816
rect 10525 816 10577 861
rect 10525 809 10534 816
rect 10534 809 10568 816
rect 10568 809 10577 816
rect 10589 816 10641 861
rect 10653 816 10705 861
rect 10717 816 10769 861
rect 10781 816 10833 861
rect 10845 816 10897 861
rect 10909 816 10961 861
rect 10589 809 10608 816
rect 10608 809 10641 816
rect 10653 809 10682 816
rect 10682 809 10705 816
rect 10717 809 10756 816
rect 10756 809 10769 816
rect 10781 809 10790 816
rect 10790 809 10830 816
rect 10830 809 10833 816
rect 10845 809 10864 816
rect 10864 809 10897 816
rect 10909 809 10938 816
rect 10938 809 10961 816
rect 10973 816 11025 861
rect 10973 809 10978 816
rect 10978 809 11012 816
rect 11012 809 11025 816
rect 11037 816 11089 861
rect 11037 809 11052 816
rect 11052 809 11086 816
rect 11086 809 11089 816
rect 11101 816 11153 861
rect 11165 816 11217 861
rect 11230 816 11282 861
rect 15040 816 15092 861
rect 15105 816 15157 861
rect 15169 816 15221 861
rect 11101 809 11126 816
rect 11126 809 11153 816
rect 11165 809 11200 816
rect 11200 809 11217 816
rect 11230 809 11234 816
rect 11234 809 11274 816
rect 11274 809 11282 816
rect 10397 782 10420 789
rect 10420 782 10449 789
rect 10461 782 10494 789
rect 10494 782 10513 789
rect 9325 744 9377 782
rect 9389 744 9441 782
rect 10397 744 10449 782
rect 10461 744 10513 782
rect 9325 737 9344 744
rect 9344 737 9377 744
rect 9389 737 9418 744
rect 9418 737 9441 744
rect 8556 710 8564 717
rect 8564 710 8604 717
rect 8604 710 8608 717
rect 8621 710 8638 717
rect 8638 710 8673 717
rect 8685 710 8712 717
rect 8712 710 8737 717
rect 4617 665 4669 710
rect 4681 665 4733 710
rect 4746 665 4798 710
rect 8556 665 8608 710
rect 8621 665 8673 710
rect 8685 665 8737 710
rect 8749 710 8752 717
rect 8752 710 8786 717
rect 8786 710 8801 717
rect 8749 665 8801 710
rect 8813 710 8826 717
rect 8826 710 8860 717
rect 8860 710 8865 717
rect 8813 665 8865 710
rect 8877 710 8900 717
rect 8900 710 8929 717
rect 8941 710 8974 717
rect 8974 710 8993 717
rect 9005 710 9008 717
rect 9008 710 9048 717
rect 9048 710 9057 717
rect 9069 710 9082 717
rect 9082 710 9121 717
rect 9133 710 9156 717
rect 9156 710 9185 717
rect 9197 710 9230 717
rect 9230 710 9249 717
rect 8877 665 8929 710
rect 8941 665 8993 710
rect 9005 665 9057 710
rect 9069 665 9121 710
rect 9133 665 9185 710
rect 9197 665 9249 710
rect 9261 710 9270 717
rect 9270 710 9304 717
rect 9304 710 9313 717
rect 9261 665 9313 710
rect 9325 710 9344 717
rect 9344 710 9377 717
rect 9389 710 9418 717
rect 9418 710 9441 717
rect 10397 737 10420 744
rect 10420 737 10449 744
rect 10461 737 10494 744
rect 10494 737 10513 744
rect 10525 782 10534 789
rect 10534 782 10568 789
rect 10568 782 10577 789
rect 10525 744 10577 782
rect 10525 737 10534 744
rect 10534 737 10568 744
rect 10568 737 10577 744
rect 10589 782 10608 789
rect 10608 782 10641 789
rect 10653 782 10682 789
rect 10682 782 10705 789
rect 10717 782 10756 789
rect 10756 782 10769 789
rect 10781 782 10790 789
rect 10790 782 10830 789
rect 10830 782 10833 789
rect 10845 782 10864 789
rect 10864 782 10897 789
rect 10909 782 10938 789
rect 10938 782 10961 789
rect 10589 744 10641 782
rect 10653 744 10705 782
rect 10717 744 10769 782
rect 10781 744 10833 782
rect 10845 744 10897 782
rect 10909 744 10961 782
rect 10589 737 10608 744
rect 10608 737 10641 744
rect 10653 737 10682 744
rect 10682 737 10705 744
rect 10717 737 10756 744
rect 10756 737 10769 744
rect 10781 737 10790 744
rect 10790 737 10830 744
rect 10830 737 10833 744
rect 10845 737 10864 744
rect 10864 737 10897 744
rect 10909 737 10938 744
rect 10938 737 10961 744
rect 10973 782 10978 789
rect 10978 782 11012 789
rect 11012 782 11025 789
rect 10973 744 11025 782
rect 10973 737 10978 744
rect 10978 737 11012 744
rect 11012 737 11025 744
rect 11037 782 11052 789
rect 11052 782 11086 789
rect 11086 782 11089 789
rect 11037 744 11089 782
rect 11037 737 11052 744
rect 11052 737 11086 744
rect 11086 737 11089 744
rect 11101 782 11126 789
rect 11126 782 11153 789
rect 11165 782 11200 789
rect 11200 782 11217 789
rect 11230 782 11234 789
rect 11234 782 11274 789
rect 11274 782 11282 789
rect 15040 809 15048 816
rect 15048 809 15088 816
rect 15088 809 15092 816
rect 15105 809 15122 816
rect 15122 809 15157 816
rect 15169 809 15196 816
rect 15196 809 15221 816
rect 15233 816 15285 861
rect 15233 809 15236 816
rect 15236 809 15270 816
rect 15270 809 15285 816
rect 15297 816 15349 861
rect 15297 809 15310 816
rect 15310 809 15344 816
rect 15344 809 15349 816
rect 15361 816 15413 861
rect 15425 816 15477 861
rect 15489 816 15541 861
rect 15553 816 15605 861
rect 15617 816 15669 861
rect 15681 816 15733 861
rect 15361 809 15384 816
rect 15384 809 15413 816
rect 15425 809 15458 816
rect 15458 809 15477 816
rect 15489 809 15492 816
rect 15492 809 15532 816
rect 15532 809 15541 816
rect 15553 809 15566 816
rect 15566 809 15605 816
rect 15617 809 15640 816
rect 15640 809 15669 816
rect 15681 809 15714 816
rect 15714 809 15733 816
rect 15745 816 15797 861
rect 15745 809 15754 816
rect 15754 809 15788 816
rect 15788 809 15797 816
rect 15809 816 15861 861
rect 15873 816 15925 861
rect 16881 816 16933 861
rect 16945 816 16997 861
rect 15809 809 15828 816
rect 15828 809 15861 816
rect 15873 809 15902 816
rect 15902 809 15925 816
rect 15040 782 15048 789
rect 15048 782 15088 789
rect 15088 782 15092 789
rect 15105 782 15122 789
rect 15122 782 15157 789
rect 15169 782 15196 789
rect 15196 782 15221 789
rect 11101 744 11153 782
rect 11165 744 11217 782
rect 11230 744 11282 782
rect 15040 744 15092 782
rect 15105 744 15157 782
rect 15169 744 15221 782
rect 11101 737 11126 744
rect 11126 737 11153 744
rect 11165 737 11200 744
rect 11200 737 11217 744
rect 11230 737 11234 744
rect 11234 737 11274 744
rect 11274 737 11282 744
rect 10397 710 10420 717
rect 10420 710 10449 717
rect 10461 710 10494 717
rect 10494 710 10513 717
rect 9325 665 9377 710
rect 9389 665 9441 710
rect 10397 665 10449 710
rect 10461 665 10513 710
rect 10525 710 10534 717
rect 10534 710 10568 717
rect 10568 710 10577 717
rect 10525 665 10577 710
rect 10589 710 10608 717
rect 10608 710 10641 717
rect 10653 710 10682 717
rect 10682 710 10705 717
rect 10717 710 10756 717
rect 10756 710 10769 717
rect 10781 710 10790 717
rect 10790 710 10830 717
rect 10830 710 10833 717
rect 10845 710 10864 717
rect 10864 710 10897 717
rect 10909 710 10938 717
rect 10938 710 10961 717
rect 10589 665 10641 710
rect 10653 665 10705 710
rect 10717 665 10769 710
rect 10781 665 10833 710
rect 10845 665 10897 710
rect 10909 665 10961 710
rect 10973 710 10978 717
rect 10978 710 11012 717
rect 11012 710 11025 717
rect 10973 665 11025 710
rect 11037 710 11052 717
rect 11052 710 11086 717
rect 11086 710 11089 717
rect 11037 665 11089 710
rect 11101 710 11126 717
rect 11126 710 11153 717
rect 11165 710 11200 717
rect 11200 710 11217 717
rect 11230 710 11234 717
rect 11234 710 11274 717
rect 11274 710 11282 717
rect 15040 737 15048 744
rect 15048 737 15088 744
rect 15088 737 15092 744
rect 15105 737 15122 744
rect 15122 737 15157 744
rect 15169 737 15196 744
rect 15196 737 15221 744
rect 15233 782 15236 789
rect 15236 782 15270 789
rect 15270 782 15285 789
rect 15233 744 15285 782
rect 15233 737 15236 744
rect 15236 737 15270 744
rect 15270 737 15285 744
rect 15297 782 15310 789
rect 15310 782 15344 789
rect 15344 782 15349 789
rect 15297 744 15349 782
rect 15297 737 15310 744
rect 15310 737 15344 744
rect 15344 737 15349 744
rect 15361 782 15384 789
rect 15384 782 15413 789
rect 15425 782 15458 789
rect 15458 782 15477 789
rect 15489 782 15492 789
rect 15492 782 15532 789
rect 15532 782 15541 789
rect 15553 782 15566 789
rect 15566 782 15605 789
rect 15617 782 15640 789
rect 15640 782 15669 789
rect 15681 782 15714 789
rect 15714 782 15733 789
rect 15361 744 15413 782
rect 15425 744 15477 782
rect 15489 744 15541 782
rect 15553 744 15605 782
rect 15617 744 15669 782
rect 15681 744 15733 782
rect 15361 737 15384 744
rect 15384 737 15413 744
rect 15425 737 15458 744
rect 15458 737 15477 744
rect 15489 737 15492 744
rect 15492 737 15532 744
rect 15532 737 15541 744
rect 15553 737 15566 744
rect 15566 737 15605 744
rect 15617 737 15640 744
rect 15640 737 15669 744
rect 15681 737 15714 744
rect 15714 737 15733 744
rect 15745 782 15754 789
rect 15754 782 15788 789
rect 15788 782 15797 789
rect 15745 744 15797 782
rect 15745 737 15754 744
rect 15754 737 15788 744
rect 15788 737 15797 744
rect 15809 782 15828 789
rect 15828 782 15861 789
rect 15873 782 15902 789
rect 15902 782 15925 789
rect 16881 809 16904 816
rect 16904 809 16933 816
rect 16945 809 16978 816
rect 16978 809 16997 816
rect 17009 816 17061 861
rect 17009 809 17018 816
rect 17018 809 17052 816
rect 17052 809 17061 816
rect 17073 816 17125 861
rect 17137 816 17189 861
rect 17201 816 17253 861
rect 17265 816 17317 861
rect 17329 816 17381 861
rect 17393 816 17445 861
rect 17073 809 17092 816
rect 17092 809 17125 816
rect 17137 809 17166 816
rect 17166 809 17189 816
rect 17201 809 17240 816
rect 17240 809 17253 816
rect 17265 809 17274 816
rect 17274 809 17314 816
rect 17314 809 17317 816
rect 17329 809 17348 816
rect 17348 809 17381 816
rect 17393 809 17422 816
rect 17422 809 17445 816
rect 17457 816 17509 861
rect 17457 809 17462 816
rect 17462 809 17496 816
rect 17496 809 17509 816
rect 17521 816 17573 861
rect 17521 809 17536 816
rect 17536 809 17570 816
rect 17570 809 17573 816
rect 17585 816 17637 861
rect 17649 816 17701 861
rect 17714 816 17766 861
rect 17585 809 17610 816
rect 17610 809 17637 816
rect 17649 809 17684 816
rect 17684 809 17701 816
rect 17714 809 17718 816
rect 17718 809 17758 816
rect 17758 809 17766 816
rect 16881 782 16904 789
rect 16904 782 16933 789
rect 16945 782 16978 789
rect 16978 782 16997 789
rect 15809 744 15861 782
rect 15873 744 15925 782
rect 16881 744 16933 782
rect 16945 744 16997 782
rect 15809 737 15828 744
rect 15828 737 15861 744
rect 15873 737 15902 744
rect 15902 737 15925 744
rect 15040 710 15048 717
rect 15048 710 15088 717
rect 15088 710 15092 717
rect 15105 710 15122 717
rect 15122 710 15157 717
rect 15169 710 15196 717
rect 15196 710 15221 717
rect 11101 665 11153 710
rect 11165 665 11217 710
rect 11230 665 11282 710
rect 15040 665 15092 710
rect 15105 665 15157 710
rect 15169 665 15221 710
rect 15233 710 15236 717
rect 15236 710 15270 717
rect 15270 710 15285 717
rect 15233 665 15285 710
rect 15297 710 15310 717
rect 15310 710 15344 717
rect 15344 710 15349 717
rect 15297 665 15349 710
rect 15361 710 15384 717
rect 15384 710 15413 717
rect 15425 710 15458 717
rect 15458 710 15477 717
rect 15489 710 15492 717
rect 15492 710 15532 717
rect 15532 710 15541 717
rect 15553 710 15566 717
rect 15566 710 15605 717
rect 15617 710 15640 717
rect 15640 710 15669 717
rect 15681 710 15714 717
rect 15714 710 15733 717
rect 15361 665 15413 710
rect 15425 665 15477 710
rect 15489 665 15541 710
rect 15553 665 15605 710
rect 15617 665 15669 710
rect 15681 665 15733 710
rect 15745 710 15754 717
rect 15754 710 15788 717
rect 15788 710 15797 717
rect 15745 665 15797 710
rect 15809 710 15828 717
rect 15828 710 15861 717
rect 15873 710 15902 717
rect 15902 710 15925 717
rect 16881 737 16904 744
rect 16904 737 16933 744
rect 16945 737 16978 744
rect 16978 737 16997 744
rect 17009 782 17018 789
rect 17018 782 17052 789
rect 17052 782 17061 789
rect 17009 744 17061 782
rect 17009 737 17018 744
rect 17018 737 17052 744
rect 17052 737 17061 744
rect 17073 782 17092 789
rect 17092 782 17125 789
rect 17137 782 17166 789
rect 17166 782 17189 789
rect 17201 782 17240 789
rect 17240 782 17253 789
rect 17265 782 17274 789
rect 17274 782 17314 789
rect 17314 782 17317 789
rect 17329 782 17348 789
rect 17348 782 17381 789
rect 17393 782 17422 789
rect 17422 782 17445 789
rect 17073 744 17125 782
rect 17137 744 17189 782
rect 17201 744 17253 782
rect 17265 744 17317 782
rect 17329 744 17381 782
rect 17393 744 17445 782
rect 17073 737 17092 744
rect 17092 737 17125 744
rect 17137 737 17166 744
rect 17166 737 17189 744
rect 17201 737 17240 744
rect 17240 737 17253 744
rect 17265 737 17274 744
rect 17274 737 17314 744
rect 17314 737 17317 744
rect 17329 737 17348 744
rect 17348 737 17381 744
rect 17393 737 17422 744
rect 17422 737 17445 744
rect 17457 782 17462 789
rect 17462 782 17496 789
rect 17496 782 17509 789
rect 17457 744 17509 782
rect 17457 737 17462 744
rect 17462 737 17496 744
rect 17496 737 17509 744
rect 17521 782 17536 789
rect 17536 782 17570 789
rect 17570 782 17573 789
rect 17521 744 17573 782
rect 17521 737 17536 744
rect 17536 737 17570 744
rect 17570 737 17573 744
rect 17585 782 17610 789
rect 17610 782 17637 789
rect 17649 782 17684 789
rect 17684 782 17701 789
rect 17714 782 17718 789
rect 17718 782 17758 789
rect 17758 782 17766 789
rect 17585 744 17637 782
rect 17649 744 17701 782
rect 17714 744 17766 782
rect 17585 737 17610 744
rect 17610 737 17637 744
rect 17649 737 17684 744
rect 17684 737 17701 744
rect 17714 737 17718 744
rect 17718 737 17758 744
rect 17758 737 17766 744
rect 16881 710 16904 717
rect 16904 710 16933 717
rect 16945 710 16978 717
rect 16978 710 16997 717
rect 15809 665 15861 710
rect 15873 665 15925 710
rect 16881 665 16933 710
rect 16945 665 16997 710
rect 17009 710 17018 717
rect 17018 710 17052 717
rect 17052 710 17061 717
rect 17009 665 17061 710
rect 17073 710 17092 717
rect 17092 710 17125 717
rect 17137 710 17166 717
rect 17166 710 17189 717
rect 17201 710 17240 717
rect 17240 710 17253 717
rect 17265 710 17274 717
rect 17274 710 17314 717
rect 17314 710 17317 717
rect 17329 710 17348 717
rect 17348 710 17381 717
rect 17393 710 17422 717
rect 17422 710 17445 717
rect 17073 665 17125 710
rect 17137 665 17189 710
rect 17201 665 17253 710
rect 17265 665 17317 710
rect 17329 665 17381 710
rect 17393 665 17445 710
rect 17457 710 17462 717
rect 17462 710 17496 717
rect 17496 710 17509 717
rect 17457 665 17509 710
rect 17521 710 17536 717
rect 17536 710 17570 717
rect 17570 710 17573 717
rect 17521 665 17573 710
rect 17585 710 17610 717
rect 17610 710 17637 717
rect 17649 710 17684 717
rect 17684 710 17701 717
rect 17714 710 17718 717
rect 17718 710 17758 717
rect 17758 710 17766 717
rect 17585 665 17637 710
rect 17649 665 17701 710
rect 17714 665 17766 710
rect 19610 588 19636 615
rect 19636 588 19662 615
rect 19610 563 19662 588
rect 1027 495 1079 547
rect 1092 495 1144 547
rect 1157 495 1209 547
rect 1222 495 1274 547
rect 1286 495 1338 547
rect 1350 495 1402 547
rect 1414 495 1466 547
rect 1478 495 1530 547
rect 1542 495 1594 547
rect 1606 495 1658 547
rect 1670 495 1722 547
rect 1734 495 1786 547
rect 1798 495 1850 547
rect 1862 495 1914 547
rect 5199 495 5251 547
rect 5263 495 5315 547
rect 5327 495 5379 547
rect 5392 495 5444 547
rect 5457 495 5509 547
rect 5522 495 5574 547
rect 5587 495 5639 547
rect 7511 495 7563 547
rect 7576 495 7628 547
rect 7641 495 7693 547
rect 7706 495 7758 547
rect 7770 495 7822 547
rect 7834 495 7886 547
rect 7898 495 7950 547
rect 7962 495 8014 547
rect 8026 495 8078 547
rect 8090 495 8142 547
rect 8154 495 8206 547
rect 8218 495 8270 547
rect 8282 495 8334 547
rect 8346 495 8398 547
rect 11440 495 11492 547
rect 11504 495 11556 547
rect 11568 495 11620 547
rect 11632 495 11684 547
rect 11696 495 11748 547
rect 11760 495 11812 547
rect 11824 495 11876 547
rect 11888 495 11940 547
rect 11952 495 12004 547
rect 12016 495 12068 547
rect 12080 495 12132 547
rect 12145 495 12197 547
rect 12210 495 12262 547
rect 12275 495 12327 547
rect 13995 495 14047 547
rect 14060 495 14112 547
rect 14125 495 14177 547
rect 14190 495 14242 547
rect 14254 495 14306 547
rect 14318 495 14370 547
rect 14382 495 14434 547
rect 14446 495 14498 547
rect 14510 495 14562 547
rect 14574 495 14626 547
rect 14638 495 14690 547
rect 14702 495 14754 547
rect 14766 495 14818 547
rect 14830 495 14882 547
rect 17924 495 17976 547
rect 17988 495 18040 547
rect 18052 495 18104 547
rect 18116 495 18168 547
rect 18180 495 18232 547
rect 18244 495 18296 547
rect 18308 495 18360 547
rect 18372 495 18424 547
rect 18436 495 18488 547
rect 18500 495 18552 547
rect 18564 495 18616 547
rect 18629 495 18681 547
rect 18694 495 18746 547
rect 18759 495 18811 547
rect 19610 499 19662 551
rect 1027 427 1079 479
rect 1092 427 1144 479
rect 1157 427 1209 479
rect 1222 427 1274 479
rect 1286 427 1338 479
rect 1350 427 1402 479
rect 1414 427 1466 479
rect 1478 427 1530 479
rect 1542 427 1594 479
rect 1606 427 1658 479
rect 1670 427 1722 479
rect 1734 427 1786 479
rect 1798 427 1850 479
rect 1862 427 1914 479
rect 5199 427 5251 479
rect 5263 427 5315 479
rect 5327 427 5379 479
rect 5392 427 5444 479
rect 5457 427 5509 479
rect 5522 427 5574 479
rect 5587 427 5639 479
rect 7511 427 7563 479
rect 7576 427 7628 479
rect 7641 427 7693 479
rect 7706 427 7758 479
rect 7770 427 7822 479
rect 7834 427 7886 479
rect 7898 427 7950 479
rect 7962 427 8014 479
rect 8026 427 8078 479
rect 8090 427 8142 479
rect 8154 427 8206 479
rect 8218 427 8270 479
rect 8282 427 8334 479
rect 8346 427 8398 479
rect 11440 427 11492 479
rect 11504 427 11556 479
rect 11568 427 11620 479
rect 11632 427 11684 479
rect 11696 427 11748 479
rect 11760 427 11812 479
rect 11824 427 11876 479
rect 11888 427 11940 479
rect 11952 427 12004 479
rect 12016 427 12068 479
rect 12080 427 12132 479
rect 12145 427 12197 479
rect 12210 427 12262 479
rect 12275 427 12327 479
rect 13995 427 14047 479
rect 14060 427 14112 479
rect 14125 427 14177 479
rect 14190 427 14242 479
rect 14254 427 14306 479
rect 14318 427 14370 479
rect 14382 427 14434 479
rect 14446 427 14498 479
rect 14510 427 14562 479
rect 14574 427 14626 479
rect 14638 427 14690 479
rect 14702 427 14754 479
rect 14766 427 14818 479
rect 14830 427 14882 479
rect 17924 427 17976 479
rect 17988 427 18040 479
rect 18052 427 18104 479
rect 18116 427 18168 479
rect 18180 427 18232 479
rect 18244 427 18296 479
rect 18308 427 18360 479
rect 18372 427 18424 479
rect 18436 427 18488 479
rect 18500 427 18552 479
rect 18564 427 18616 479
rect 18629 427 18681 479
rect 18694 427 18746 479
rect 18759 427 18811 479
rect 1027 404 1079 411
rect 1027 370 1055 404
rect 1055 370 1079 404
rect 1027 359 1079 370
rect 1092 404 1144 411
rect 1092 370 1094 404
rect 1094 370 1128 404
rect 1128 370 1144 404
rect 1092 359 1144 370
rect 1157 404 1209 411
rect 1157 370 1167 404
rect 1167 370 1201 404
rect 1201 370 1209 404
rect 1157 359 1209 370
rect 1222 404 1274 411
rect 1222 370 1240 404
rect 1240 370 1274 404
rect 1222 359 1274 370
rect 1286 404 1338 411
rect 1350 404 1402 411
rect 1414 404 1466 411
rect 1478 404 1530 411
rect 1542 404 1594 411
rect 1606 404 1658 411
rect 1286 370 1313 404
rect 1313 370 1338 404
rect 1350 370 1386 404
rect 1386 370 1402 404
rect 1414 370 1420 404
rect 1420 370 1459 404
rect 1459 370 1466 404
rect 1478 370 1493 404
rect 1493 370 1530 404
rect 1542 370 1566 404
rect 1566 370 1594 404
rect 1606 370 1639 404
rect 1639 370 1658 404
rect 1286 359 1338 370
rect 1350 359 1402 370
rect 1414 359 1466 370
rect 1478 359 1530 370
rect 1542 359 1594 370
rect 1606 359 1658 370
rect 1670 404 1722 411
rect 1670 370 1678 404
rect 1678 370 1712 404
rect 1712 370 1722 404
rect 1670 359 1722 370
rect 1734 404 1786 411
rect 1734 370 1751 404
rect 1751 370 1785 404
rect 1785 370 1786 404
rect 1734 359 1786 370
rect 1798 404 1850 411
rect 1862 404 1914 411
rect 5199 404 5251 411
rect 5263 404 5315 411
rect 5327 404 5379 411
rect 5392 404 5444 411
rect 5457 404 5509 411
rect 1798 370 1824 404
rect 1824 370 1850 404
rect 1862 370 1898 404
rect 1898 370 1914 404
rect 5199 370 5231 404
rect 5231 370 5251 404
rect 5263 370 5265 404
rect 5265 370 5304 404
rect 5304 370 5315 404
rect 5327 370 5338 404
rect 5338 370 5377 404
rect 5377 370 5379 404
rect 5392 370 5411 404
rect 5411 370 5444 404
rect 5457 370 5484 404
rect 5484 370 5509 404
rect 1798 359 1850 370
rect 1862 359 1914 370
rect 5199 359 5251 370
rect 5263 359 5315 370
rect 5327 359 5379 370
rect 5392 359 5444 370
rect 5457 359 5509 370
rect 5522 404 5574 411
rect 5522 370 5523 404
rect 5523 370 5557 404
rect 5557 370 5574 404
rect 5522 359 5574 370
rect 5587 404 5639 411
rect 7511 404 7563 411
rect 5587 370 5596 404
rect 5596 370 5630 404
rect 5630 370 5639 404
rect 7511 370 7539 404
rect 7539 370 7563 404
rect 5587 359 5639 370
rect 7511 359 7563 370
rect 7576 404 7628 411
rect 7576 370 7578 404
rect 7578 370 7612 404
rect 7612 370 7628 404
rect 7576 359 7628 370
rect 7641 404 7693 411
rect 7641 370 7651 404
rect 7651 370 7685 404
rect 7685 370 7693 404
rect 7641 359 7693 370
rect 7706 404 7758 411
rect 7706 370 7724 404
rect 7724 370 7758 404
rect 7706 359 7758 370
rect 7770 404 7822 411
rect 7834 404 7886 411
rect 7898 404 7950 411
rect 7962 404 8014 411
rect 8026 404 8078 411
rect 8090 404 8142 411
rect 7770 370 7797 404
rect 7797 370 7822 404
rect 7834 370 7870 404
rect 7870 370 7886 404
rect 7898 370 7904 404
rect 7904 370 7943 404
rect 7943 370 7950 404
rect 7962 370 7977 404
rect 7977 370 8014 404
rect 8026 370 8050 404
rect 8050 370 8078 404
rect 8090 370 8123 404
rect 8123 370 8142 404
rect 7770 359 7822 370
rect 7834 359 7886 370
rect 7898 359 7950 370
rect 7962 359 8014 370
rect 8026 359 8078 370
rect 8090 359 8142 370
rect 8154 404 8206 411
rect 8154 370 8162 404
rect 8162 370 8196 404
rect 8196 370 8206 404
rect 8154 359 8206 370
rect 8218 404 8270 411
rect 8218 370 8235 404
rect 8235 370 8269 404
rect 8269 370 8270 404
rect 8218 359 8270 370
rect 8282 404 8334 411
rect 8346 404 8398 411
rect 11440 404 11492 411
rect 11504 404 11556 411
rect 8282 370 8308 404
rect 8308 370 8334 404
rect 8346 370 8382 404
rect 8382 370 8398 404
rect 11440 370 11456 404
rect 11456 370 11492 404
rect 11504 370 11530 404
rect 11530 370 11556 404
rect 8282 359 8334 370
rect 8346 359 8398 370
rect 11440 359 11492 370
rect 11504 359 11556 370
rect 11568 404 11620 411
rect 11568 370 11569 404
rect 11569 370 11603 404
rect 11603 370 11620 404
rect 11568 359 11620 370
rect 11632 404 11684 411
rect 11632 370 11642 404
rect 11642 370 11676 404
rect 11676 370 11684 404
rect 11632 359 11684 370
rect 11696 404 11748 411
rect 11760 404 11812 411
rect 11824 404 11876 411
rect 11888 404 11940 411
rect 11952 404 12004 411
rect 12016 404 12068 411
rect 11696 370 11715 404
rect 11715 370 11748 404
rect 11760 370 11788 404
rect 11788 370 11812 404
rect 11824 370 11861 404
rect 11861 370 11876 404
rect 11888 370 11895 404
rect 11895 370 11934 404
rect 11934 370 11940 404
rect 11952 370 11968 404
rect 11968 370 12004 404
rect 12016 370 12041 404
rect 12041 370 12068 404
rect 11696 359 11748 370
rect 11760 359 11812 370
rect 11824 359 11876 370
rect 11888 359 11940 370
rect 11952 359 12004 370
rect 12016 359 12068 370
rect 12080 404 12132 411
rect 12080 370 12114 404
rect 12114 370 12132 404
rect 12080 359 12132 370
rect 12145 404 12197 411
rect 12145 370 12153 404
rect 12153 370 12187 404
rect 12187 370 12197 404
rect 12145 359 12197 370
rect 12210 404 12262 411
rect 12210 370 12226 404
rect 12226 370 12260 404
rect 12260 370 12262 404
rect 12210 359 12262 370
rect 12275 404 12327 411
rect 13995 404 14047 411
rect 12275 370 12299 404
rect 12299 370 12327 404
rect 13995 370 14023 404
rect 14023 370 14047 404
rect 12275 359 12327 370
rect 13995 359 14047 370
rect 14060 404 14112 411
rect 14060 370 14062 404
rect 14062 370 14096 404
rect 14096 370 14112 404
rect 14060 359 14112 370
rect 14125 404 14177 411
rect 14125 370 14135 404
rect 14135 370 14169 404
rect 14169 370 14177 404
rect 14125 359 14177 370
rect 14190 404 14242 411
rect 14190 370 14208 404
rect 14208 370 14242 404
rect 14190 359 14242 370
rect 14254 404 14306 411
rect 14318 404 14370 411
rect 14382 404 14434 411
rect 14446 404 14498 411
rect 14510 404 14562 411
rect 14574 404 14626 411
rect 14254 370 14281 404
rect 14281 370 14306 404
rect 14318 370 14354 404
rect 14354 370 14370 404
rect 14382 370 14388 404
rect 14388 370 14427 404
rect 14427 370 14434 404
rect 14446 370 14461 404
rect 14461 370 14498 404
rect 14510 370 14534 404
rect 14534 370 14562 404
rect 14574 370 14607 404
rect 14607 370 14626 404
rect 14254 359 14306 370
rect 14318 359 14370 370
rect 14382 359 14434 370
rect 14446 359 14498 370
rect 14510 359 14562 370
rect 14574 359 14626 370
rect 14638 404 14690 411
rect 14638 370 14646 404
rect 14646 370 14680 404
rect 14680 370 14690 404
rect 14638 359 14690 370
rect 14702 404 14754 411
rect 14702 370 14719 404
rect 14719 370 14753 404
rect 14753 370 14754 404
rect 14702 359 14754 370
rect 14766 404 14818 411
rect 14830 404 14882 411
rect 17924 404 17976 411
rect 17988 404 18040 411
rect 14766 370 14792 404
rect 14792 370 14818 404
rect 14830 370 14866 404
rect 14866 370 14882 404
rect 17924 370 17940 404
rect 17940 370 17976 404
rect 17988 370 18014 404
rect 18014 370 18040 404
rect 14766 359 14818 370
rect 14830 359 14882 370
rect 17924 359 17976 370
rect 17988 359 18040 370
rect 18052 404 18104 411
rect 18052 370 18053 404
rect 18053 370 18087 404
rect 18087 370 18104 404
rect 18052 359 18104 370
rect 18116 404 18168 411
rect 18116 370 18126 404
rect 18126 370 18160 404
rect 18160 370 18168 404
rect 18116 359 18168 370
rect 18180 404 18232 411
rect 18244 404 18296 411
rect 18308 404 18360 411
rect 18372 404 18424 411
rect 18436 404 18488 411
rect 18500 404 18552 411
rect 18180 370 18199 404
rect 18199 370 18232 404
rect 18244 370 18272 404
rect 18272 370 18296 404
rect 18308 370 18345 404
rect 18345 370 18360 404
rect 18372 370 18379 404
rect 18379 370 18418 404
rect 18418 370 18424 404
rect 18436 370 18452 404
rect 18452 370 18488 404
rect 18500 370 18525 404
rect 18525 370 18552 404
rect 18180 359 18232 370
rect 18244 359 18296 370
rect 18308 359 18360 370
rect 18372 359 18424 370
rect 18436 359 18488 370
rect 18500 359 18552 370
rect 18564 404 18616 411
rect 18564 370 18598 404
rect 18598 370 18616 404
rect 18564 359 18616 370
rect 18629 404 18681 411
rect 18629 370 18637 404
rect 18637 370 18671 404
rect 18671 370 18681 404
rect 18629 359 18681 370
rect 18694 404 18746 411
rect 18694 370 18710 404
rect 18710 370 18744 404
rect 18744 370 18746 404
rect 18694 359 18746 370
rect 18759 404 18811 411
rect 18759 370 18783 404
rect 18783 370 18811 404
rect 18759 359 18811 370
rect 1027 332 1079 343
rect 1027 298 1055 332
rect 1055 298 1079 332
rect 1027 291 1079 298
rect 1092 332 1144 343
rect 1092 298 1094 332
rect 1094 298 1128 332
rect 1128 298 1144 332
rect 1092 291 1144 298
rect 1157 332 1209 343
rect 1157 298 1167 332
rect 1167 298 1201 332
rect 1201 298 1209 332
rect 1157 291 1209 298
rect 1222 332 1274 343
rect 1222 298 1240 332
rect 1240 298 1274 332
rect 1222 291 1274 298
rect 1286 332 1338 343
rect 1350 332 1402 343
rect 1414 332 1466 343
rect 1478 332 1530 343
rect 1542 332 1594 343
rect 1606 332 1658 343
rect 1286 298 1313 332
rect 1313 298 1338 332
rect 1350 298 1386 332
rect 1386 298 1402 332
rect 1414 298 1420 332
rect 1420 298 1459 332
rect 1459 298 1466 332
rect 1478 298 1493 332
rect 1493 298 1530 332
rect 1542 298 1566 332
rect 1566 298 1594 332
rect 1606 298 1639 332
rect 1639 298 1658 332
rect 1286 291 1338 298
rect 1350 291 1402 298
rect 1414 291 1466 298
rect 1478 291 1530 298
rect 1542 291 1594 298
rect 1606 291 1658 298
rect 1670 332 1722 343
rect 1670 298 1678 332
rect 1678 298 1712 332
rect 1712 298 1722 332
rect 1670 291 1722 298
rect 1734 332 1786 343
rect 1734 298 1751 332
rect 1751 298 1785 332
rect 1785 298 1786 332
rect 1734 291 1786 298
rect 1798 332 1850 343
rect 1862 332 1914 343
rect 5199 332 5251 343
rect 5263 332 5315 343
rect 5327 332 5379 343
rect 5392 332 5444 343
rect 5457 332 5509 343
rect 1798 298 1824 332
rect 1824 298 1850 332
rect 1862 298 1898 332
rect 1898 298 1914 332
rect 5199 298 5231 332
rect 5231 298 5251 332
rect 5263 298 5265 332
rect 5265 298 5304 332
rect 5304 298 5315 332
rect 5327 298 5338 332
rect 5338 298 5377 332
rect 5377 298 5379 332
rect 5392 298 5411 332
rect 5411 298 5444 332
rect 5457 298 5484 332
rect 5484 298 5509 332
rect 1798 291 1850 298
rect 1862 291 1914 298
rect 5199 291 5251 298
rect 5263 291 5315 298
rect 5327 291 5379 298
rect 5392 291 5444 298
rect 5457 291 5509 298
rect 5522 332 5574 343
rect 5522 298 5523 332
rect 5523 298 5557 332
rect 5557 298 5574 332
rect 5522 291 5574 298
rect 5587 332 5639 343
rect 7511 332 7563 343
rect 5587 298 5596 332
rect 5596 298 5630 332
rect 5630 298 5639 332
rect 7511 298 7539 332
rect 7539 298 7563 332
rect 5587 291 5639 298
rect 7511 291 7563 298
rect 7576 332 7628 343
rect 7576 298 7578 332
rect 7578 298 7612 332
rect 7612 298 7628 332
rect 7576 291 7628 298
rect 7641 332 7693 343
rect 7641 298 7651 332
rect 7651 298 7685 332
rect 7685 298 7693 332
rect 7641 291 7693 298
rect 7706 332 7758 343
rect 7706 298 7724 332
rect 7724 298 7758 332
rect 7706 291 7758 298
rect 7770 332 7822 343
rect 7834 332 7886 343
rect 7898 332 7950 343
rect 7962 332 8014 343
rect 8026 332 8078 343
rect 8090 332 8142 343
rect 7770 298 7797 332
rect 7797 298 7822 332
rect 7834 298 7870 332
rect 7870 298 7886 332
rect 7898 298 7904 332
rect 7904 298 7943 332
rect 7943 298 7950 332
rect 7962 298 7977 332
rect 7977 298 8014 332
rect 8026 298 8050 332
rect 8050 298 8078 332
rect 8090 298 8123 332
rect 8123 298 8142 332
rect 7770 291 7822 298
rect 7834 291 7886 298
rect 7898 291 7950 298
rect 7962 291 8014 298
rect 8026 291 8078 298
rect 8090 291 8142 298
rect 8154 332 8206 343
rect 8154 298 8162 332
rect 8162 298 8196 332
rect 8196 298 8206 332
rect 8154 291 8206 298
rect 8218 332 8270 343
rect 8218 298 8235 332
rect 8235 298 8269 332
rect 8269 298 8270 332
rect 8218 291 8270 298
rect 8282 332 8334 343
rect 8346 332 8398 343
rect 11440 332 11492 343
rect 11504 332 11556 343
rect 8282 298 8308 332
rect 8308 298 8334 332
rect 8346 298 8382 332
rect 8382 298 8398 332
rect 11440 298 11456 332
rect 11456 298 11492 332
rect 11504 298 11530 332
rect 11530 298 11556 332
rect 8282 291 8334 298
rect 8346 291 8398 298
rect 11440 291 11492 298
rect 11504 291 11556 298
rect 11568 332 11620 343
rect 11568 298 11569 332
rect 11569 298 11603 332
rect 11603 298 11620 332
rect 11568 291 11620 298
rect 11632 332 11684 343
rect 11632 298 11642 332
rect 11642 298 11676 332
rect 11676 298 11684 332
rect 11632 291 11684 298
rect 11696 332 11748 343
rect 11760 332 11812 343
rect 11824 332 11876 343
rect 11888 332 11940 343
rect 11952 332 12004 343
rect 12016 332 12068 343
rect 11696 298 11715 332
rect 11715 298 11748 332
rect 11760 298 11788 332
rect 11788 298 11812 332
rect 11824 298 11861 332
rect 11861 298 11876 332
rect 11888 298 11895 332
rect 11895 298 11934 332
rect 11934 298 11940 332
rect 11952 298 11968 332
rect 11968 298 12004 332
rect 12016 298 12041 332
rect 12041 298 12068 332
rect 11696 291 11748 298
rect 11760 291 11812 298
rect 11824 291 11876 298
rect 11888 291 11940 298
rect 11952 291 12004 298
rect 12016 291 12068 298
rect 12080 332 12132 343
rect 12080 298 12114 332
rect 12114 298 12132 332
rect 12080 291 12132 298
rect 12145 332 12197 343
rect 12145 298 12153 332
rect 12153 298 12187 332
rect 12187 298 12197 332
rect 12145 291 12197 298
rect 12210 332 12262 343
rect 12210 298 12226 332
rect 12226 298 12260 332
rect 12260 298 12262 332
rect 12210 291 12262 298
rect 12275 332 12327 343
rect 13995 332 14047 343
rect 12275 298 12299 332
rect 12299 298 12327 332
rect 13995 298 14023 332
rect 14023 298 14047 332
rect 12275 291 12327 298
rect 13995 291 14047 298
rect 14060 332 14112 343
rect 14060 298 14062 332
rect 14062 298 14096 332
rect 14096 298 14112 332
rect 14060 291 14112 298
rect 14125 332 14177 343
rect 14125 298 14135 332
rect 14135 298 14169 332
rect 14169 298 14177 332
rect 14125 291 14177 298
rect 14190 332 14242 343
rect 14190 298 14208 332
rect 14208 298 14242 332
rect 14190 291 14242 298
rect 14254 332 14306 343
rect 14318 332 14370 343
rect 14382 332 14434 343
rect 14446 332 14498 343
rect 14510 332 14562 343
rect 14574 332 14626 343
rect 14254 298 14281 332
rect 14281 298 14306 332
rect 14318 298 14354 332
rect 14354 298 14370 332
rect 14382 298 14388 332
rect 14388 298 14427 332
rect 14427 298 14434 332
rect 14446 298 14461 332
rect 14461 298 14498 332
rect 14510 298 14534 332
rect 14534 298 14562 332
rect 14574 298 14607 332
rect 14607 298 14626 332
rect 14254 291 14306 298
rect 14318 291 14370 298
rect 14382 291 14434 298
rect 14446 291 14498 298
rect 14510 291 14562 298
rect 14574 291 14626 298
rect 14638 332 14690 343
rect 14638 298 14646 332
rect 14646 298 14680 332
rect 14680 298 14690 332
rect 14638 291 14690 298
rect 14702 332 14754 343
rect 14702 298 14719 332
rect 14719 298 14753 332
rect 14753 298 14754 332
rect 14702 291 14754 298
rect 14766 332 14818 343
rect 14830 332 14882 343
rect 17924 332 17976 343
rect 17988 332 18040 343
rect 14766 298 14792 332
rect 14792 298 14818 332
rect 14830 298 14866 332
rect 14866 298 14882 332
rect 17924 298 17940 332
rect 17940 298 17976 332
rect 17988 298 18014 332
rect 18014 298 18040 332
rect 14766 291 14818 298
rect 14830 291 14882 298
rect 17924 291 17976 298
rect 17988 291 18040 298
rect 18052 332 18104 343
rect 18052 298 18053 332
rect 18053 298 18087 332
rect 18087 298 18104 332
rect 18052 291 18104 298
rect 18116 332 18168 343
rect 18116 298 18126 332
rect 18126 298 18160 332
rect 18160 298 18168 332
rect 18116 291 18168 298
rect 18180 332 18232 343
rect 18244 332 18296 343
rect 18308 332 18360 343
rect 18372 332 18424 343
rect 18436 332 18488 343
rect 18500 332 18552 343
rect 18180 298 18199 332
rect 18199 298 18232 332
rect 18244 298 18272 332
rect 18272 298 18296 332
rect 18308 298 18345 332
rect 18345 298 18360 332
rect 18372 298 18379 332
rect 18379 298 18418 332
rect 18418 298 18424 332
rect 18436 298 18452 332
rect 18452 298 18488 332
rect 18500 298 18525 332
rect 18525 298 18552 332
rect 18180 291 18232 298
rect 18244 291 18296 298
rect 18308 291 18360 298
rect 18372 291 18424 298
rect 18436 291 18488 298
rect 18500 291 18552 298
rect 18564 332 18616 343
rect 18564 298 18598 332
rect 18598 298 18616 332
rect 18564 291 18616 298
rect 18629 332 18681 343
rect 18629 298 18637 332
rect 18637 298 18671 332
rect 18671 298 18681 332
rect 18629 291 18681 298
rect 18694 332 18746 343
rect 18694 298 18710 332
rect 18710 298 18744 332
rect 18744 298 18746 332
rect 18694 291 18746 298
rect 18759 332 18811 343
rect 18759 298 18783 332
rect 18783 298 18811 332
rect 18759 291 18811 298
rect 1027 223 1079 275
rect 1092 223 1144 275
rect 1157 223 1209 275
rect 1222 223 1274 275
rect 1286 223 1338 275
rect 1350 223 1402 275
rect 1414 223 1466 275
rect 1478 223 1530 275
rect 1542 223 1594 275
rect 1606 223 1658 275
rect 1670 223 1722 275
rect 1734 223 1786 275
rect 1798 223 1850 275
rect 1862 223 1914 275
rect 5199 223 5251 275
rect 5263 223 5315 275
rect 5327 223 5379 275
rect 5392 223 5444 275
rect 5457 223 5509 275
rect 5522 223 5574 275
rect 5587 223 5639 275
rect 7511 223 7563 275
rect 7576 223 7628 275
rect 7641 223 7693 275
rect 7706 223 7758 275
rect 7770 223 7822 275
rect 7834 223 7886 275
rect 7898 223 7950 275
rect 7962 223 8014 275
rect 8026 223 8078 275
rect 8090 223 8142 275
rect 8154 223 8206 275
rect 8218 223 8270 275
rect 8282 223 8334 275
rect 8346 223 8398 275
rect 11440 223 11492 275
rect 11504 223 11556 275
rect 11568 223 11620 275
rect 11632 223 11684 275
rect 11696 223 11748 275
rect 11760 223 11812 275
rect 11824 223 11876 275
rect 11888 223 11940 275
rect 11952 223 12004 275
rect 12016 223 12068 275
rect 12080 223 12132 275
rect 12145 223 12197 275
rect 12210 223 12262 275
rect 12275 223 12327 275
rect 13995 223 14047 275
rect 14060 223 14112 275
rect 14125 223 14177 275
rect 14190 223 14242 275
rect 14254 223 14306 275
rect 14318 223 14370 275
rect 14382 223 14434 275
rect 14446 223 14498 275
rect 14510 223 14562 275
rect 14574 223 14626 275
rect 14638 223 14690 275
rect 14702 223 14754 275
rect 14766 223 14818 275
rect 14830 223 14882 275
rect 17924 223 17976 275
rect 17988 223 18040 275
rect 18052 223 18104 275
rect 18116 223 18168 275
rect 18180 223 18232 275
rect 18244 223 18296 275
rect 18308 223 18360 275
rect 18372 223 18424 275
rect 18436 223 18488 275
rect 18500 223 18552 275
rect 18564 223 18616 275
rect 18629 223 18681 275
rect 18694 223 18746 275
rect 18759 223 18811 275
rect -138 100 -86 152
rect -138 36 -86 88
rect -138 -198 -86 -146
rect -138 -262 -86 -210
rect 176 151 228 203
rect 1027 155 1079 207
rect 1092 155 1144 207
rect 1157 155 1209 207
rect 1222 155 1274 207
rect 1286 155 1338 207
rect 1350 155 1402 207
rect 1414 155 1466 207
rect 1478 155 1530 207
rect 1542 155 1594 207
rect 1606 155 1658 207
rect 1670 155 1722 207
rect 1734 155 1786 207
rect 1798 155 1850 207
rect 1862 155 1914 207
rect 5199 155 5251 207
rect 5263 155 5315 207
rect 5327 155 5379 207
rect 5392 155 5444 207
rect 5457 155 5509 207
rect 5522 155 5574 207
rect 5587 155 5639 207
rect 7511 155 7563 207
rect 7576 155 7628 207
rect 7641 155 7693 207
rect 7706 155 7758 207
rect 7770 155 7822 207
rect 7834 155 7886 207
rect 7898 155 7950 207
rect 7962 155 8014 207
rect 8026 155 8078 207
rect 8090 155 8142 207
rect 8154 155 8206 207
rect 8218 155 8270 207
rect 8282 155 8334 207
rect 8346 155 8398 207
rect 11440 155 11492 207
rect 11504 155 11556 207
rect 11568 155 11620 207
rect 11632 155 11684 207
rect 11696 155 11748 207
rect 11760 155 11812 207
rect 11824 155 11876 207
rect 11888 155 11940 207
rect 11952 155 12004 207
rect 12016 155 12068 207
rect 12080 155 12132 207
rect 12145 155 12197 207
rect 12210 155 12262 207
rect 12275 155 12327 207
rect 13995 155 14047 207
rect 14060 155 14112 207
rect 14125 155 14177 207
rect 14190 155 14242 207
rect 14254 155 14306 207
rect 14318 155 14370 207
rect 14382 155 14434 207
rect 14446 155 14498 207
rect 14510 155 14562 207
rect 14574 155 14626 207
rect 14638 155 14690 207
rect 14702 155 14754 207
rect 14766 155 14818 207
rect 14830 155 14882 207
rect 17924 155 17976 207
rect 17988 155 18040 207
rect 18052 155 18104 207
rect 18116 155 18168 207
rect 18180 155 18232 207
rect 18244 155 18296 207
rect 18308 155 18360 207
rect 18372 155 18424 207
rect 18436 155 18488 207
rect 18500 155 18552 207
rect 18564 155 18616 207
rect 18629 155 18681 207
rect 18694 155 18746 207
rect 18759 155 18811 207
rect 19610 151 19662 203
rect 176 114 228 139
rect 176 87 202 114
rect 202 87 228 114
rect 19610 114 19662 139
rect 19610 87 19622 114
rect 19622 87 19660 114
rect 19660 87 19662 114
rect 3913 -8 3965 38
rect 3978 -8 4030 38
rect 3913 -14 3936 -8
rect 3936 -14 3965 -8
rect 3978 -14 4010 -8
rect 4010 -14 4030 -8
rect 4042 -8 4094 38
rect 4042 -14 4050 -8
rect 4050 -14 4084 -8
rect 4084 -14 4094 -8
rect 4106 -8 4158 38
rect 4106 -14 4124 -8
rect 4124 -14 4158 -8
rect 4170 -8 4222 38
rect 4234 -8 4286 38
rect 4298 -8 4350 38
rect 4362 -8 4414 38
rect 4426 -8 4478 38
rect 4170 -14 4198 -8
rect 4198 -14 4222 -8
rect 4234 -14 4272 -8
rect 4272 -14 4286 -8
rect 4298 -14 4306 -8
rect 4306 -14 4346 -8
rect 4346 -14 4350 -8
rect 4362 -14 4380 -8
rect 4380 -14 4414 -8
rect 4426 -14 4454 -8
rect 4454 -14 4478 -8
rect 4490 -8 4542 38
rect 4490 -14 4494 -8
rect 4494 -14 4528 -8
rect 4528 -14 4542 -8
rect 4554 -8 4606 38
rect 4554 -14 4568 -8
rect 4568 -14 4602 -8
rect 4602 -14 4606 -8
rect 4618 -8 4670 38
rect 4682 -8 4734 38
rect 4746 -8 4798 38
rect 8556 -8 8608 38
rect 8621 -8 8673 38
rect 8685 -8 8737 38
rect 4618 -14 4642 -8
rect 4642 -14 4670 -8
rect 4682 -14 4716 -8
rect 4716 -14 4734 -8
rect 4746 -14 4750 -8
rect 4750 -14 4790 -8
rect 4790 -14 4798 -8
rect 3913 -42 3936 -34
rect 3936 -42 3965 -34
rect 3978 -42 4010 -34
rect 4010 -42 4030 -34
rect 3913 -80 3965 -42
rect 3978 -80 4030 -42
rect 3913 -86 3936 -80
rect 3936 -86 3965 -80
rect 3978 -86 4010 -80
rect 4010 -86 4030 -80
rect 4042 -42 4050 -34
rect 4050 -42 4084 -34
rect 4084 -42 4094 -34
rect 4042 -80 4094 -42
rect 4042 -86 4050 -80
rect 4050 -86 4084 -80
rect 4084 -86 4094 -80
rect 4106 -42 4124 -34
rect 4124 -42 4158 -34
rect 4106 -80 4158 -42
rect 4106 -86 4124 -80
rect 4124 -86 4158 -80
rect 4170 -42 4198 -34
rect 4198 -42 4222 -34
rect 4234 -42 4272 -34
rect 4272 -42 4286 -34
rect 4298 -42 4306 -34
rect 4306 -42 4346 -34
rect 4346 -42 4350 -34
rect 4362 -42 4380 -34
rect 4380 -42 4414 -34
rect 4426 -42 4454 -34
rect 4454 -42 4478 -34
rect 4170 -80 4222 -42
rect 4234 -80 4286 -42
rect 4298 -80 4350 -42
rect 4362 -80 4414 -42
rect 4426 -80 4478 -42
rect 4170 -86 4198 -80
rect 4198 -86 4222 -80
rect 4234 -86 4272 -80
rect 4272 -86 4286 -80
rect 4298 -86 4306 -80
rect 4306 -86 4346 -80
rect 4346 -86 4350 -80
rect 4362 -86 4380 -80
rect 4380 -86 4414 -80
rect 4426 -86 4454 -80
rect 4454 -86 4478 -80
rect 4490 -42 4494 -34
rect 4494 -42 4528 -34
rect 4528 -42 4542 -34
rect 4490 -80 4542 -42
rect 4490 -86 4494 -80
rect 4494 -86 4528 -80
rect 4528 -86 4542 -80
rect 4554 -42 4568 -34
rect 4568 -42 4602 -34
rect 4602 -42 4606 -34
rect 4554 -80 4606 -42
rect 4554 -86 4568 -80
rect 4568 -86 4602 -80
rect 4602 -86 4606 -80
rect 4618 -42 4642 -34
rect 4642 -42 4670 -34
rect 4682 -42 4716 -34
rect 4716 -42 4734 -34
rect 4746 -42 4750 -34
rect 4750 -42 4790 -34
rect 4790 -42 4798 -34
rect 8556 -14 8564 -8
rect 8564 -14 8604 -8
rect 8604 -14 8608 -8
rect 8621 -14 8638 -8
rect 8638 -14 8673 -8
rect 8685 -14 8712 -8
rect 8712 -14 8737 -8
rect 8749 -8 8801 38
rect 8749 -14 8752 -8
rect 8752 -14 8786 -8
rect 8786 -14 8801 -8
rect 8813 -8 8865 38
rect 8813 -14 8826 -8
rect 8826 -14 8860 -8
rect 8860 -14 8865 -8
rect 8877 -8 8929 38
rect 8941 -8 8993 38
rect 9005 -8 9057 38
rect 9069 -8 9121 38
rect 9133 -8 9185 38
rect 9197 -8 9249 38
rect 8877 -14 8900 -8
rect 8900 -14 8929 -8
rect 8941 -14 8974 -8
rect 8974 -14 8993 -8
rect 9005 -14 9008 -8
rect 9008 -14 9048 -8
rect 9048 -14 9057 -8
rect 9069 -14 9082 -8
rect 9082 -14 9121 -8
rect 9133 -14 9156 -8
rect 9156 -14 9185 -8
rect 9197 -14 9230 -8
rect 9230 -14 9249 -8
rect 9261 -8 9313 38
rect 9261 -14 9270 -8
rect 9270 -14 9304 -8
rect 9304 -14 9313 -8
rect 9325 -8 9377 38
rect 9389 -8 9441 38
rect 10397 -8 10449 38
rect 10462 -8 10514 38
rect 9325 -14 9344 -8
rect 9344 -14 9377 -8
rect 9389 -14 9418 -8
rect 9418 -14 9441 -8
rect 8556 -42 8564 -34
rect 8564 -42 8604 -34
rect 8604 -42 8608 -34
rect 8621 -42 8638 -34
rect 8638 -42 8673 -34
rect 8685 -42 8712 -34
rect 8712 -42 8737 -34
rect 4618 -80 4670 -42
rect 4682 -80 4734 -42
rect 4746 -80 4798 -42
rect 8556 -80 8608 -42
rect 8621 -80 8673 -42
rect 8685 -80 8737 -42
rect 4618 -86 4642 -80
rect 4642 -86 4670 -80
rect 4682 -86 4716 -80
rect 4716 -86 4734 -80
rect 4746 -86 4750 -80
rect 4750 -86 4790 -80
rect 4790 -86 4798 -80
rect 3913 -114 3936 -106
rect 3936 -114 3965 -106
rect 3978 -114 4010 -106
rect 4010 -114 4030 -106
rect 3913 -158 3965 -114
rect 3978 -158 4030 -114
rect 4042 -114 4050 -106
rect 4050 -114 4084 -106
rect 4084 -114 4094 -106
rect 4042 -158 4094 -114
rect 4106 -114 4124 -106
rect 4124 -114 4158 -106
rect 4106 -158 4158 -114
rect 4170 -114 4198 -106
rect 4198 -114 4222 -106
rect 4234 -114 4272 -106
rect 4272 -114 4286 -106
rect 4298 -114 4306 -106
rect 4306 -114 4346 -106
rect 4346 -114 4350 -106
rect 4362 -114 4380 -106
rect 4380 -114 4414 -106
rect 4426 -114 4454 -106
rect 4454 -114 4478 -106
rect 4170 -158 4222 -114
rect 4234 -158 4286 -114
rect 4298 -158 4350 -114
rect 4362 -158 4414 -114
rect 4426 -158 4478 -114
rect 4490 -114 4494 -106
rect 4494 -114 4528 -106
rect 4528 -114 4542 -106
rect 4490 -158 4542 -114
rect 4554 -114 4568 -106
rect 4568 -114 4602 -106
rect 4602 -114 4606 -106
rect 4554 -158 4606 -114
rect 4618 -114 4642 -106
rect 4642 -114 4670 -106
rect 4682 -114 4716 -106
rect 4716 -114 4734 -106
rect 4746 -114 4750 -106
rect 4750 -114 4790 -106
rect 4790 -114 4798 -106
rect 8556 -86 8564 -80
rect 8564 -86 8604 -80
rect 8604 -86 8608 -80
rect 8621 -86 8638 -80
rect 8638 -86 8673 -80
rect 8685 -86 8712 -80
rect 8712 -86 8737 -80
rect 8749 -42 8752 -34
rect 8752 -42 8786 -34
rect 8786 -42 8801 -34
rect 8749 -80 8801 -42
rect 8749 -86 8752 -80
rect 8752 -86 8786 -80
rect 8786 -86 8801 -80
rect 8813 -42 8826 -34
rect 8826 -42 8860 -34
rect 8860 -42 8865 -34
rect 8813 -80 8865 -42
rect 8813 -86 8826 -80
rect 8826 -86 8860 -80
rect 8860 -86 8865 -80
rect 8877 -42 8900 -34
rect 8900 -42 8929 -34
rect 8941 -42 8974 -34
rect 8974 -42 8993 -34
rect 9005 -42 9008 -34
rect 9008 -42 9048 -34
rect 9048 -42 9057 -34
rect 9069 -42 9082 -34
rect 9082 -42 9121 -34
rect 9133 -42 9156 -34
rect 9156 -42 9185 -34
rect 9197 -42 9230 -34
rect 9230 -42 9249 -34
rect 8877 -80 8929 -42
rect 8941 -80 8993 -42
rect 9005 -80 9057 -42
rect 9069 -80 9121 -42
rect 9133 -80 9185 -42
rect 9197 -80 9249 -42
rect 8877 -86 8900 -80
rect 8900 -86 8929 -80
rect 8941 -86 8974 -80
rect 8974 -86 8993 -80
rect 9005 -86 9008 -80
rect 9008 -86 9048 -80
rect 9048 -86 9057 -80
rect 9069 -86 9082 -80
rect 9082 -86 9121 -80
rect 9133 -86 9156 -80
rect 9156 -86 9185 -80
rect 9197 -86 9230 -80
rect 9230 -86 9249 -80
rect 9261 -42 9270 -34
rect 9270 -42 9304 -34
rect 9304 -42 9313 -34
rect 9261 -80 9313 -42
rect 9261 -86 9270 -80
rect 9270 -86 9304 -80
rect 9304 -86 9313 -80
rect 9325 -42 9344 -34
rect 9344 -42 9377 -34
rect 9389 -42 9418 -34
rect 9418 -42 9441 -34
rect 10397 -14 10420 -8
rect 10420 -14 10449 -8
rect 10462 -14 10494 -8
rect 10494 -14 10514 -8
rect 10526 -8 10578 38
rect 10526 -14 10534 -8
rect 10534 -14 10568 -8
rect 10568 -14 10578 -8
rect 10590 -8 10642 38
rect 10590 -14 10608 -8
rect 10608 -14 10642 -8
rect 10654 -8 10706 38
rect 10718 -8 10770 38
rect 10782 -8 10834 38
rect 10846 -8 10898 38
rect 10910 -8 10962 38
rect 10654 -14 10682 -8
rect 10682 -14 10706 -8
rect 10718 -14 10756 -8
rect 10756 -14 10770 -8
rect 10782 -14 10790 -8
rect 10790 -14 10830 -8
rect 10830 -14 10834 -8
rect 10846 -14 10864 -8
rect 10864 -14 10898 -8
rect 10910 -14 10938 -8
rect 10938 -14 10962 -8
rect 10974 -8 11026 38
rect 10974 -14 10978 -8
rect 10978 -14 11012 -8
rect 11012 -14 11026 -8
rect 11038 -8 11090 38
rect 11038 -14 11052 -8
rect 11052 -14 11086 -8
rect 11086 -14 11090 -8
rect 11102 -8 11154 38
rect 11166 -8 11218 38
rect 11230 -8 11282 38
rect 15040 -8 15092 37
rect 15105 -8 15157 37
rect 15169 -8 15221 37
rect 11102 -14 11126 -8
rect 11126 -14 11154 -8
rect 11166 -14 11200 -8
rect 11200 -14 11218 -8
rect 11230 -14 11234 -8
rect 11234 -14 11274 -8
rect 11274 -14 11282 -8
rect 10397 -42 10420 -34
rect 10420 -42 10449 -34
rect 10462 -42 10494 -34
rect 10494 -42 10514 -34
rect 9325 -80 9377 -42
rect 9389 -80 9441 -42
rect 10397 -80 10449 -42
rect 10462 -80 10514 -42
rect 9325 -86 9344 -80
rect 9344 -86 9377 -80
rect 9389 -86 9418 -80
rect 9418 -86 9441 -80
rect 8556 -114 8564 -106
rect 8564 -114 8604 -106
rect 8604 -114 8608 -106
rect 8621 -114 8638 -106
rect 8638 -114 8673 -106
rect 8685 -114 8712 -106
rect 8712 -114 8737 -106
rect 4618 -158 4670 -114
rect 4682 -158 4734 -114
rect 4746 -158 4798 -114
rect 8556 -158 8608 -114
rect 8621 -158 8673 -114
rect 8685 -158 8737 -114
rect 8749 -114 8752 -106
rect 8752 -114 8786 -106
rect 8786 -114 8801 -106
rect 8749 -158 8801 -114
rect 8813 -114 8826 -106
rect 8826 -114 8860 -106
rect 8860 -114 8865 -106
rect 8813 -158 8865 -114
rect 8877 -114 8900 -106
rect 8900 -114 8929 -106
rect 8941 -114 8974 -106
rect 8974 -114 8993 -106
rect 9005 -114 9008 -106
rect 9008 -114 9048 -106
rect 9048 -114 9057 -106
rect 9069 -114 9082 -106
rect 9082 -114 9121 -106
rect 9133 -114 9156 -106
rect 9156 -114 9185 -106
rect 9197 -114 9230 -106
rect 9230 -114 9249 -106
rect 8877 -158 8929 -114
rect 8941 -158 8993 -114
rect 9005 -158 9057 -114
rect 9069 -158 9121 -114
rect 9133 -158 9185 -114
rect 9197 -158 9249 -114
rect 9261 -114 9270 -106
rect 9270 -114 9304 -106
rect 9304 -114 9313 -106
rect 9261 -158 9313 -114
rect 9325 -114 9344 -106
rect 9344 -114 9377 -106
rect 9389 -114 9418 -106
rect 9418 -114 9441 -106
rect 10397 -86 10420 -80
rect 10420 -86 10449 -80
rect 10462 -86 10494 -80
rect 10494 -86 10514 -80
rect 10526 -42 10534 -34
rect 10534 -42 10568 -34
rect 10568 -42 10578 -34
rect 10526 -80 10578 -42
rect 10526 -86 10534 -80
rect 10534 -86 10568 -80
rect 10568 -86 10578 -80
rect 10590 -42 10608 -34
rect 10608 -42 10642 -34
rect 10590 -80 10642 -42
rect 10590 -86 10608 -80
rect 10608 -86 10642 -80
rect 10654 -42 10682 -34
rect 10682 -42 10706 -34
rect 10718 -42 10756 -34
rect 10756 -42 10770 -34
rect 10782 -42 10790 -34
rect 10790 -42 10830 -34
rect 10830 -42 10834 -34
rect 10846 -42 10864 -34
rect 10864 -42 10898 -34
rect 10910 -42 10938 -34
rect 10938 -42 10962 -34
rect 10654 -80 10706 -42
rect 10718 -80 10770 -42
rect 10782 -80 10834 -42
rect 10846 -80 10898 -42
rect 10910 -80 10962 -42
rect 10654 -86 10682 -80
rect 10682 -86 10706 -80
rect 10718 -86 10756 -80
rect 10756 -86 10770 -80
rect 10782 -86 10790 -80
rect 10790 -86 10830 -80
rect 10830 -86 10834 -80
rect 10846 -86 10864 -80
rect 10864 -86 10898 -80
rect 10910 -86 10938 -80
rect 10938 -86 10962 -80
rect 10974 -42 10978 -34
rect 10978 -42 11012 -34
rect 11012 -42 11026 -34
rect 10974 -80 11026 -42
rect 10974 -86 10978 -80
rect 10978 -86 11012 -80
rect 11012 -86 11026 -80
rect 11038 -42 11052 -34
rect 11052 -42 11086 -34
rect 11086 -42 11090 -34
rect 11038 -80 11090 -42
rect 11038 -86 11052 -80
rect 11052 -86 11086 -80
rect 11086 -86 11090 -80
rect 11102 -42 11126 -34
rect 11126 -42 11154 -34
rect 11166 -42 11200 -34
rect 11200 -42 11218 -34
rect 11230 -42 11234 -34
rect 11234 -42 11274 -34
rect 11274 -42 11282 -34
rect 15040 -15 15048 -8
rect 15048 -15 15088 -8
rect 15088 -15 15092 -8
rect 15105 -15 15122 -8
rect 15122 -15 15157 -8
rect 15169 -15 15196 -8
rect 15196 -15 15221 -8
rect 15233 -8 15285 37
rect 15233 -15 15236 -8
rect 15236 -15 15270 -8
rect 15270 -15 15285 -8
rect 15297 -8 15349 37
rect 15297 -15 15310 -8
rect 15310 -15 15344 -8
rect 15344 -15 15349 -8
rect 15361 -8 15413 37
rect 15425 -8 15477 37
rect 15489 -8 15541 37
rect 15553 -8 15605 37
rect 15617 -8 15669 37
rect 15681 -8 15733 37
rect 15361 -15 15384 -8
rect 15384 -15 15413 -8
rect 15425 -15 15458 -8
rect 15458 -15 15477 -8
rect 15489 -15 15492 -8
rect 15492 -15 15532 -8
rect 15532 -15 15541 -8
rect 15553 -15 15566 -8
rect 15566 -15 15605 -8
rect 15617 -15 15640 -8
rect 15640 -15 15669 -8
rect 15681 -15 15714 -8
rect 15714 -15 15733 -8
rect 15745 -8 15797 37
rect 15745 -15 15754 -8
rect 15754 -15 15788 -8
rect 15788 -15 15797 -8
rect 15809 -8 15861 37
rect 15873 -8 15925 37
rect 16881 -8 16933 37
rect 16946 -8 16998 37
rect 15809 -15 15828 -8
rect 15828 -15 15861 -8
rect 15873 -15 15902 -8
rect 15902 -15 15925 -8
rect 15040 -42 15048 -35
rect 15048 -42 15088 -35
rect 15088 -42 15092 -35
rect 15105 -42 15122 -35
rect 15122 -42 15157 -35
rect 15169 -42 15196 -35
rect 15196 -42 15221 -35
rect 11102 -80 11154 -42
rect 11166 -80 11218 -42
rect 11230 -80 11282 -42
rect 15040 -80 15092 -42
rect 15105 -80 15157 -42
rect 15169 -80 15221 -42
rect 11102 -86 11126 -80
rect 11126 -86 11154 -80
rect 11166 -86 11200 -80
rect 11200 -86 11218 -80
rect 11230 -86 11234 -80
rect 11234 -86 11274 -80
rect 11274 -86 11282 -80
rect 10397 -114 10420 -106
rect 10420 -114 10449 -106
rect 10462 -114 10494 -106
rect 10494 -114 10514 -106
rect 9325 -158 9377 -114
rect 9389 -158 9441 -114
rect 10397 -158 10449 -114
rect 10462 -158 10514 -114
rect 10526 -114 10534 -106
rect 10534 -114 10568 -106
rect 10568 -114 10578 -106
rect 10526 -158 10578 -114
rect 10590 -114 10608 -106
rect 10608 -114 10642 -106
rect 10590 -158 10642 -114
rect 10654 -114 10682 -106
rect 10682 -114 10706 -106
rect 10718 -114 10756 -106
rect 10756 -114 10770 -106
rect 10782 -114 10790 -106
rect 10790 -114 10830 -106
rect 10830 -114 10834 -106
rect 10846 -114 10864 -106
rect 10864 -114 10898 -106
rect 10910 -114 10938 -106
rect 10938 -114 10962 -106
rect 10654 -158 10706 -114
rect 10718 -158 10770 -114
rect 10782 -158 10834 -114
rect 10846 -158 10898 -114
rect 10910 -158 10962 -114
rect 10974 -114 10978 -106
rect 10978 -114 11012 -106
rect 11012 -114 11026 -106
rect 10974 -158 11026 -114
rect 11038 -114 11052 -106
rect 11052 -114 11086 -106
rect 11086 -114 11090 -106
rect 11038 -158 11090 -114
rect 11102 -114 11126 -106
rect 11126 -114 11154 -106
rect 11166 -114 11200 -106
rect 11200 -114 11218 -106
rect 11230 -114 11234 -106
rect 11234 -114 11274 -106
rect 11274 -114 11282 -106
rect 15040 -87 15048 -80
rect 15048 -87 15088 -80
rect 15088 -87 15092 -80
rect 15105 -87 15122 -80
rect 15122 -87 15157 -80
rect 15169 -87 15196 -80
rect 15196 -87 15221 -80
rect 15233 -42 15236 -35
rect 15236 -42 15270 -35
rect 15270 -42 15285 -35
rect 15233 -80 15285 -42
rect 15233 -87 15236 -80
rect 15236 -87 15270 -80
rect 15270 -87 15285 -80
rect 15297 -42 15310 -35
rect 15310 -42 15344 -35
rect 15344 -42 15349 -35
rect 15297 -80 15349 -42
rect 15297 -87 15310 -80
rect 15310 -87 15344 -80
rect 15344 -87 15349 -80
rect 15361 -42 15384 -35
rect 15384 -42 15413 -35
rect 15425 -42 15458 -35
rect 15458 -42 15477 -35
rect 15489 -42 15492 -35
rect 15492 -42 15532 -35
rect 15532 -42 15541 -35
rect 15553 -42 15566 -35
rect 15566 -42 15605 -35
rect 15617 -42 15640 -35
rect 15640 -42 15669 -35
rect 15681 -42 15714 -35
rect 15714 -42 15733 -35
rect 15361 -80 15413 -42
rect 15425 -80 15477 -42
rect 15489 -80 15541 -42
rect 15553 -80 15605 -42
rect 15617 -80 15669 -42
rect 15681 -80 15733 -42
rect 15361 -87 15384 -80
rect 15384 -87 15413 -80
rect 15425 -87 15458 -80
rect 15458 -87 15477 -80
rect 15489 -87 15492 -80
rect 15492 -87 15532 -80
rect 15532 -87 15541 -80
rect 15553 -87 15566 -80
rect 15566 -87 15605 -80
rect 15617 -87 15640 -80
rect 15640 -87 15669 -80
rect 15681 -87 15714 -80
rect 15714 -87 15733 -80
rect 15745 -42 15754 -35
rect 15754 -42 15788 -35
rect 15788 -42 15797 -35
rect 15745 -80 15797 -42
rect 15745 -87 15754 -80
rect 15754 -87 15788 -80
rect 15788 -87 15797 -80
rect 15809 -42 15828 -35
rect 15828 -42 15861 -35
rect 15873 -42 15902 -35
rect 15902 -42 15925 -35
rect 16881 -15 16904 -8
rect 16904 -15 16933 -8
rect 16946 -15 16978 -8
rect 16978 -15 16998 -8
rect 17010 -8 17062 37
rect 17010 -15 17018 -8
rect 17018 -15 17052 -8
rect 17052 -15 17062 -8
rect 17074 -8 17126 37
rect 17074 -15 17092 -8
rect 17092 -15 17126 -8
rect 17138 -8 17190 37
rect 17202 -8 17254 37
rect 17266 -8 17318 37
rect 17330 -8 17382 37
rect 17394 -8 17446 37
rect 17138 -15 17166 -8
rect 17166 -15 17190 -8
rect 17202 -15 17240 -8
rect 17240 -15 17254 -8
rect 17266 -15 17274 -8
rect 17274 -15 17314 -8
rect 17314 -15 17318 -8
rect 17330 -15 17348 -8
rect 17348 -15 17382 -8
rect 17394 -15 17422 -8
rect 17422 -15 17446 -8
rect 17458 -8 17510 37
rect 17458 -15 17462 -8
rect 17462 -15 17496 -8
rect 17496 -15 17510 -8
rect 17522 -8 17574 37
rect 17522 -15 17536 -8
rect 17536 -15 17570 -8
rect 17570 -15 17574 -8
rect 17586 -8 17638 37
rect 17650 -8 17702 37
rect 17714 -8 17766 37
rect 17586 -15 17610 -8
rect 17610 -15 17638 -8
rect 17650 -15 17684 -8
rect 17684 -15 17702 -8
rect 17714 -15 17718 -8
rect 17718 -15 17758 -8
rect 17758 -15 17766 -8
rect 16881 -42 16904 -35
rect 16904 -42 16933 -35
rect 16946 -42 16978 -35
rect 16978 -42 16998 -35
rect 15809 -80 15861 -42
rect 15873 -80 15925 -42
rect 16881 -80 16933 -42
rect 16946 -80 16998 -42
rect 15809 -87 15828 -80
rect 15828 -87 15861 -80
rect 15873 -87 15902 -80
rect 15902 -87 15925 -80
rect 15040 -114 15048 -107
rect 15048 -114 15088 -107
rect 15088 -114 15092 -107
rect 15105 -114 15122 -107
rect 15122 -114 15157 -107
rect 15169 -114 15196 -107
rect 15196 -114 15221 -107
rect 11102 -158 11154 -114
rect 11166 -158 11218 -114
rect 11230 -158 11282 -114
rect 15040 -159 15092 -114
rect 15105 -159 15157 -114
rect 15169 -159 15221 -114
rect 15233 -114 15236 -107
rect 15236 -114 15270 -107
rect 15270 -114 15285 -107
rect 15233 -159 15285 -114
rect 15297 -114 15310 -107
rect 15310 -114 15344 -107
rect 15344 -114 15349 -107
rect 15297 -159 15349 -114
rect 15361 -114 15384 -107
rect 15384 -114 15413 -107
rect 15425 -114 15458 -107
rect 15458 -114 15477 -107
rect 15489 -114 15492 -107
rect 15492 -114 15532 -107
rect 15532 -114 15541 -107
rect 15553 -114 15566 -107
rect 15566 -114 15605 -107
rect 15617 -114 15640 -107
rect 15640 -114 15669 -107
rect 15681 -114 15714 -107
rect 15714 -114 15733 -107
rect 15361 -159 15413 -114
rect 15425 -159 15477 -114
rect 15489 -159 15541 -114
rect 15553 -159 15605 -114
rect 15617 -159 15669 -114
rect 15681 -159 15733 -114
rect 15745 -114 15754 -107
rect 15754 -114 15788 -107
rect 15788 -114 15797 -107
rect 15745 -159 15797 -114
rect 15809 -114 15828 -107
rect 15828 -114 15861 -107
rect 15873 -114 15902 -107
rect 15902 -114 15925 -107
rect 16881 -87 16904 -80
rect 16904 -87 16933 -80
rect 16946 -87 16978 -80
rect 16978 -87 16998 -80
rect 17010 -42 17018 -35
rect 17018 -42 17052 -35
rect 17052 -42 17062 -35
rect 17010 -80 17062 -42
rect 17010 -87 17018 -80
rect 17018 -87 17052 -80
rect 17052 -87 17062 -80
rect 17074 -42 17092 -35
rect 17092 -42 17126 -35
rect 17074 -80 17126 -42
rect 17074 -87 17092 -80
rect 17092 -87 17126 -80
rect 17138 -42 17166 -35
rect 17166 -42 17190 -35
rect 17202 -42 17240 -35
rect 17240 -42 17254 -35
rect 17266 -42 17274 -35
rect 17274 -42 17314 -35
rect 17314 -42 17318 -35
rect 17330 -42 17348 -35
rect 17348 -42 17382 -35
rect 17394 -42 17422 -35
rect 17422 -42 17446 -35
rect 17138 -80 17190 -42
rect 17202 -80 17254 -42
rect 17266 -80 17318 -42
rect 17330 -80 17382 -42
rect 17394 -80 17446 -42
rect 17138 -87 17166 -80
rect 17166 -87 17190 -80
rect 17202 -87 17240 -80
rect 17240 -87 17254 -80
rect 17266 -87 17274 -80
rect 17274 -87 17314 -80
rect 17314 -87 17318 -80
rect 17330 -87 17348 -80
rect 17348 -87 17382 -80
rect 17394 -87 17422 -80
rect 17422 -87 17446 -80
rect 17458 -42 17462 -35
rect 17462 -42 17496 -35
rect 17496 -42 17510 -35
rect 17458 -80 17510 -42
rect 17458 -87 17462 -80
rect 17462 -87 17496 -80
rect 17496 -87 17510 -80
rect 17522 -42 17536 -35
rect 17536 -42 17570 -35
rect 17570 -42 17574 -35
rect 17522 -80 17574 -42
rect 17522 -87 17536 -80
rect 17536 -87 17570 -80
rect 17570 -87 17574 -80
rect 17586 -42 17610 -35
rect 17610 -42 17638 -35
rect 17650 -42 17684 -35
rect 17684 -42 17702 -35
rect 17714 -42 17718 -35
rect 17718 -42 17758 -35
rect 17758 -42 17766 -35
rect 17586 -80 17638 -42
rect 17650 -80 17702 -42
rect 17714 -80 17766 -42
rect 17586 -87 17610 -80
rect 17610 -87 17638 -80
rect 17650 -87 17684 -80
rect 17684 -87 17702 -80
rect 17714 -87 17718 -80
rect 17718 -87 17758 -80
rect 17758 -87 17766 -80
rect 16881 -114 16904 -107
rect 16904 -114 16933 -107
rect 16946 -114 16978 -107
rect 16978 -114 16998 -107
rect 15809 -159 15861 -114
rect 15873 -159 15925 -114
rect 16881 -159 16933 -114
rect 16946 -159 16998 -114
rect 17010 -114 17018 -107
rect 17018 -114 17052 -107
rect 17052 -114 17062 -107
rect 17010 -159 17062 -114
rect 17074 -114 17092 -107
rect 17092 -114 17126 -107
rect 17074 -159 17126 -114
rect 17138 -114 17166 -107
rect 17166 -114 17190 -107
rect 17202 -114 17240 -107
rect 17240 -114 17254 -107
rect 17266 -114 17274 -107
rect 17274 -114 17314 -107
rect 17314 -114 17318 -107
rect 17330 -114 17348 -107
rect 17348 -114 17382 -107
rect 17394 -114 17422 -107
rect 17422 -114 17446 -107
rect 17138 -159 17190 -114
rect 17202 -159 17254 -114
rect 17266 -159 17318 -114
rect 17330 -159 17382 -114
rect 17394 -159 17446 -114
rect 17458 -114 17462 -107
rect 17462 -114 17496 -107
rect 17496 -114 17510 -107
rect 17458 -159 17510 -114
rect 17522 -114 17536 -107
rect 17536 -114 17570 -107
rect 17570 -114 17574 -107
rect 17522 -159 17574 -114
rect 17586 -114 17610 -107
rect 17610 -114 17638 -107
rect 17650 -114 17684 -107
rect 17684 -114 17702 -107
rect 17714 -114 17718 -107
rect 17718 -114 17758 -107
rect 17758 -114 17766 -107
rect 17586 -159 17638 -114
rect 17650 -159 17702 -114
rect 17714 -159 17766 -114
rect 19759 -70 19811 -18
rect 19759 -134 19811 -82
rect 20006 975 20058 1027
rect 20006 911 20058 963
rect 20006 563 20058 615
rect 20006 499 20058 551
rect 20006 182 20058 234
rect 20006 118 20058 170
rect 20198 975 20250 1027
rect 20198 911 20250 963
rect 20006 11 20058 63
rect 20006 -53 20058 -1
rect 673 -238 725 -229
rect 747 -238 799 -229
rect 821 -238 873 -229
rect 895 -238 947 -229
rect 6018 -238 6070 -229
rect 6085 -238 6137 -229
rect 6152 -238 6204 -229
rect 6219 -238 6271 -229
rect 6286 -238 6338 -229
rect 6353 -238 6405 -229
rect 6949 -238 7001 -229
rect 7016 -238 7068 -229
rect 7083 -238 7135 -229
rect 7150 -238 7202 -229
rect 7217 -238 7269 -229
rect 7284 -238 7336 -229
rect 12502 -238 12554 -228
rect 12569 -238 12621 -228
rect 12636 -238 12688 -228
rect 12703 -238 12755 -228
rect 12770 -238 12822 -228
rect 12837 -238 12889 -228
rect 13433 -238 13485 -229
rect 13500 -238 13552 -229
rect 13567 -238 13619 -229
rect 13634 -238 13686 -229
rect 13701 -238 13753 -229
rect 13768 -238 13820 -229
rect 19071 -238 19123 -229
rect 19155 -238 19207 -229
rect 673 -272 690 -238
rect 690 -272 725 -238
rect 747 -272 762 -238
rect 762 -272 799 -238
rect 821 -272 834 -238
rect 834 -272 872 -238
rect 872 -272 873 -238
rect 895 -272 906 -238
rect 906 -272 944 -238
rect 944 -272 947 -238
rect 6018 -272 6056 -238
rect 6056 -272 6070 -238
rect 6085 -272 6090 -238
rect 6090 -272 6128 -238
rect 6128 -272 6137 -238
rect 6152 -272 6162 -238
rect 6162 -272 6200 -238
rect 6200 -272 6204 -238
rect 6219 -272 6234 -238
rect 6234 -272 6271 -238
rect 6286 -272 6306 -238
rect 6306 -272 6338 -238
rect 6353 -272 6378 -238
rect 6378 -272 6405 -238
rect 6949 -272 6954 -238
rect 6954 -272 6992 -238
rect 6992 -272 7001 -238
rect 7016 -272 7026 -238
rect 7026 -272 7064 -238
rect 7064 -272 7068 -238
rect 7083 -272 7098 -238
rect 7098 -272 7135 -238
rect 7150 -272 7170 -238
rect 7170 -272 7202 -238
rect 7217 -272 7242 -238
rect 7242 -272 7269 -238
rect 7284 -272 7314 -238
rect 7314 -272 7336 -238
rect 12502 -272 12536 -238
rect 12536 -272 12554 -238
rect 12569 -272 12570 -238
rect 12570 -272 12608 -238
rect 12608 -272 12621 -238
rect 12636 -272 12642 -238
rect 12642 -272 12680 -238
rect 12680 -272 12688 -238
rect 12703 -272 12714 -238
rect 12714 -272 12752 -238
rect 12752 -272 12755 -238
rect 12770 -272 12786 -238
rect 12786 -272 12822 -238
rect 12837 -272 12858 -238
rect 12858 -272 12889 -238
rect 13433 -272 13434 -238
rect 13434 -272 13472 -238
rect 13472 -272 13485 -238
rect 13500 -272 13506 -238
rect 13506 -272 13544 -238
rect 13544 -272 13552 -238
rect 13567 -272 13578 -238
rect 13578 -272 13616 -238
rect 13616 -272 13619 -238
rect 13634 -272 13650 -238
rect 13650 -272 13686 -238
rect 13701 -272 13722 -238
rect 13722 -272 13753 -238
rect 13768 -272 13794 -238
rect 13794 -272 13820 -238
rect 19071 -272 19097 -238
rect 19097 -272 19123 -238
rect 19155 -272 19170 -238
rect 19170 -272 19204 -238
rect 19204 -272 19207 -238
rect 673 -281 725 -272
rect 747 -281 799 -272
rect 821 -281 873 -272
rect 895 -281 947 -272
rect 6018 -281 6070 -272
rect 6085 -281 6137 -272
rect 6152 -281 6204 -272
rect 6219 -281 6271 -272
rect 6286 -281 6338 -272
rect 6353 -281 6405 -272
rect 6949 -281 7001 -272
rect 7016 -281 7068 -272
rect 7083 -281 7135 -272
rect 7150 -281 7202 -272
rect 7217 -281 7269 -272
rect 7284 -281 7336 -272
rect 12502 -280 12554 -272
rect 12569 -280 12621 -272
rect 12636 -280 12688 -272
rect 12703 -280 12755 -272
rect 12770 -280 12822 -272
rect 12837 -280 12889 -272
rect 13433 -281 13485 -272
rect 13500 -281 13552 -272
rect 13567 -281 13619 -272
rect 13634 -281 13686 -272
rect 13701 -281 13753 -272
rect 13768 -281 13820 -272
rect 19071 -281 19123 -272
rect 19155 -281 19207 -272
rect 19238 -238 19290 -229
rect 19321 -238 19373 -229
rect 19238 -272 19243 -238
rect 19243 -272 19277 -238
rect 19277 -272 19290 -238
rect 19321 -272 19350 -238
rect 19350 -272 19373 -238
rect 19238 -281 19290 -272
rect 19321 -281 19373 -272
rect 3714 -469 3766 -417
rect 3778 -469 3830 -417
rect 20430 170 20482 222
rect 20430 106 20482 158
rect 22755 -59 22871 57
rect 15045 -2923 15097 -2871
rect 15113 -2923 15165 -2871
rect 15181 -2923 15233 -2871
rect 15249 -2923 15301 -2871
rect 15317 -2923 15369 -2871
rect 15385 -2923 15437 -2871
rect 15453 -2923 15505 -2871
rect 15521 -2923 15573 -2871
rect 15589 -2923 15641 -2871
rect 15657 -2923 15709 -2871
rect 15725 -2923 15777 -2871
rect 15793 -2923 15845 -2871
rect 15861 -2923 15913 -2871
rect 16886 -2923 16938 -2871
rect 16954 -2923 17006 -2871
rect 17022 -2923 17074 -2871
rect 17090 -2923 17142 -2871
rect 17158 -2923 17210 -2871
rect 17226 -2923 17278 -2871
rect 17294 -2923 17346 -2871
rect 17362 -2923 17414 -2871
rect 17430 -2923 17482 -2871
rect 17498 -2923 17550 -2871
rect 17566 -2923 17618 -2871
rect 17634 -2923 17686 -2871
rect 17702 -2923 17754 -2871
<< metal2 >>
rect -1610 14169 -1360 14199
rect -1610 14117 -1604 14169
rect -1552 14117 -1511 14169
rect -1459 14117 -1418 14169
rect -1366 14117 -1360 14169
rect -1610 14087 -1360 14117
rect -1450 12311 -1398 12317
tri -1481 12272 -1450 12303 se
rect -2262 12259 -1450 12272
rect -2262 12247 -1398 12259
rect -2262 12220 -1450 12247
rect -2262 12195 -2203 12220
tri -2203 12195 -2178 12220 nw
tri -1480 12195 -1455 12220 ne
rect -1455 12195 -1450 12220
rect -2262 7178 -2210 12195
tri -2210 12188 -2203 12195 nw
tri -1455 12190 -1450 12195 ne
rect -1450 12183 -1398 12195
rect -1450 12125 -1398 12131
rect -1606 11973 -905 11979
rect -1554 11921 -1294 11973
rect -1242 11921 -905 11973
rect -1606 11909 -905 11921
rect -1554 11857 -1294 11909
rect -1242 11857 -905 11909
rect -1606 11845 -905 11857
rect -1554 11793 -1294 11845
rect -1242 11793 -905 11845
rect -1606 11787 -905 11793
tri -1000 11744 -957 11787 ne
rect -1606 11649 -1032 11655
rect -1554 11597 -1294 11649
rect -1242 11597 -1032 11649
rect -1606 11585 -1032 11597
rect -1554 11533 -1294 11585
rect -1242 11533 -1032 11585
rect -1606 11521 -1032 11533
rect -1554 11469 -1294 11521
rect -1242 11469 -1032 11521
rect -1606 11463 -1032 11469
tri -1107 11440 -1084 11463 ne
rect -1450 11311 -1398 11317
tri -1455 11247 -1450 11252 se
rect -1450 11247 -1398 11259
tri -1480 11222 -1455 11247 se
rect -1455 11222 -1450 11247
rect -2422 7126 -2210 7178
rect -2174 11195 -1450 11222
rect -2174 11183 -1398 11195
rect -2174 11170 -1450 11183
rect -2422 1782 -2370 7126
rect -2174 2406 -2122 11170
tri -2122 11138 -2090 11170 nw
tri -1481 11139 -1450 11170 ne
rect -1450 11125 -1398 11131
rect -1450 10847 -1398 10853
tri -1481 10808 -1450 10839 se
rect -2090 10795 -1450 10808
rect -2090 10783 -1398 10795
rect -2090 10756 -1450 10783
rect -2090 10731 -2031 10756
tri -2031 10731 -2006 10756 nw
tri -1480 10731 -1455 10756 ne
rect -1455 10731 -1450 10756
rect -2090 2651 -2038 10731
tri -2038 10724 -2031 10731 nw
tri -1455 10726 -1450 10731 ne
rect -1450 10719 -1398 10731
rect -1450 10661 -1398 10667
rect -1606 10509 -1124 10515
rect -1554 10457 -1294 10509
rect -1242 10457 -1124 10509
rect -1606 10445 -1124 10457
rect -1554 10393 -1294 10445
rect -1242 10393 -1124 10445
rect -1606 10381 -1124 10393
rect -1554 10329 -1294 10381
rect -1242 10329 -1124 10381
rect -1606 10323 -1124 10329
rect -1636 5832 -1584 5838
rect -1636 5757 -1584 5780
rect -1636 4307 -1584 5705
rect -1176 5015 -1124 10323
rect -1084 5061 -1032 11463
rect -957 6223 -905 11787
rect -957 6148 -905 6171
rect 21783 6171 23006 6177
rect -957 6090 -905 6096
rect 19684 6074 19690 6126
rect 19742 6074 19757 6126
rect 19809 6074 19824 6126
rect 19876 6074 19960 6126
tri 19820 6052 19842 6074 ne
rect 19842 6052 19960 6074
tri 19842 6046 19848 6052 ne
rect 19848 6046 19960 6052
rect 21835 6119 21847 6171
rect 21899 6137 23006 6171
tri 23006 6137 23046 6177 sw
rect 21899 6119 23046 6137
rect 21783 6104 23046 6119
rect 21835 6052 21847 6104
rect 21899 6052 23046 6104
rect 21783 6046 23046 6052
tri 19848 6044 19850 6046 ne
tri 19820 5928 19850 5958 se
rect 19850 5928 19960 6046
tri 22906 6016 22936 6046 ne
rect 19820 5876 19960 5928
tri 19820 5846 19850 5876 ne
rect 19666 5445 19675 5501
rect 19731 5499 19755 5501
rect 19742 5447 19754 5499
rect 19731 5445 19755 5447
rect 19811 5445 19820 5501
rect 3023 5079 3029 5131
rect 3081 5128 3095 5131
rect 3147 5128 3161 5131
rect 3213 5128 3227 5131
rect 3279 5128 3293 5131
rect 3089 5079 3095 5128
rect 3345 5079 3358 5131
rect 3410 5128 3423 5131
rect 3475 5128 3488 5131
rect 3540 5128 3553 5131
rect 3605 5128 3618 5131
rect 3417 5079 3423 5128
rect 3605 5079 3607 5128
rect 3670 5079 3683 5131
rect 3735 5128 3748 5131
rect 3800 5128 3813 5131
rect 3865 5128 3878 5131
rect 3930 5128 3943 5131
rect 3745 5079 3748 5128
rect 3930 5079 3935 5128
rect 3995 5079 4008 5131
rect 4060 5128 4073 5131
rect 4125 5128 4138 5131
rect 4190 5128 4203 5131
rect 4255 5128 4268 5131
rect 4072 5079 4073 5128
rect 4255 5079 4259 5128
rect 4320 5079 4326 5131
tri -1084 5021 -1044 5061 ne
rect -1044 5021 -1032 5061
tri -1032 5021 -975 5078 sw
rect 3023 5072 3033 5079
rect 3089 5072 3115 5079
rect 3171 5072 3197 5079
rect 3253 5072 3279 5079
rect 3335 5072 3361 5079
rect 3417 5072 3443 5079
rect 3499 5072 3525 5079
rect 3581 5072 3607 5079
rect 3663 5072 3689 5079
rect 3745 5072 3771 5079
rect 3827 5072 3853 5079
rect 3909 5072 3935 5079
rect 3991 5072 4016 5079
rect 4072 5072 4097 5079
rect 4153 5072 4178 5079
rect 4234 5072 4259 5079
rect 4315 5072 4326 5079
tri -1124 5015 -1118 5021 sw
tri -1044 5015 -1038 5021 ne
rect -1038 5015 -975 5021
tri -975 5015 -969 5021 sw
rect -1176 5009 -1118 5015
tri -1118 5009 -1112 5015 sw
tri -1038 5009 -1032 5015 ne
rect -1032 5009 -969 5015
rect -1176 5004 -1112 5009
tri -1176 4963 -1135 5004 ne
rect -1135 4963 -1112 5004
tri -1112 4963 -1066 5009 sw
tri -1032 4991 -1014 5009 ne
tri -1135 4961 -1133 4963 ne
rect -1133 4961 -1066 4963
tri -1066 4961 -1064 4963 sw
tri -1133 4952 -1124 4961 ne
rect -1124 4952 -1064 4961
tri -1124 4937 -1109 4952 ne
tri -1156 4706 -1109 4753 se
rect -1109 4726 -1064 4952
rect -1109 4713 -1077 4726
tri -1077 4713 -1064 4726 nw
rect -1109 4706 -1084 4713
tri -1084 4706 -1077 4713 nw
tri -1021 4706 -1014 4713 se
rect -1014 4706 -969 5009
rect 3023 5020 4326 5072
rect 3023 5015 3033 5020
rect 3089 5015 3115 5020
rect 3171 5015 3197 5020
rect 3253 5015 3279 5020
rect 3335 5015 3361 5020
rect 3417 5015 3443 5020
rect 3499 5015 3525 5020
rect 3581 5015 3607 5020
rect 3663 5015 3689 5020
rect 3745 5015 3771 5020
rect 3827 5015 3853 5020
rect 3909 5015 3935 5020
rect 3991 5015 4016 5020
rect 4072 5015 4097 5020
rect 4153 5015 4178 5020
rect 4234 5015 4259 5020
rect 4315 5015 4326 5020
rect 3023 4963 3029 5015
rect 3089 4964 3095 5015
rect 3081 4963 3095 4964
rect 3147 4963 3161 4964
rect 3213 4963 3227 4964
rect 3279 4963 3293 4964
rect 3345 4963 3358 5015
rect 3417 4964 3423 5015
rect 3605 4964 3607 5015
rect 3410 4963 3423 4964
rect 3475 4963 3488 4964
rect 3540 4963 3553 4964
rect 3605 4963 3618 4964
rect 3670 4963 3683 5015
rect 3745 4964 3748 5015
rect 3930 4964 3935 5015
rect 3735 4963 3748 4964
rect 3800 4963 3813 4964
rect 3865 4963 3878 4964
rect 3930 4963 3943 4964
rect 3995 4963 4008 5015
rect 4072 4964 4073 5015
rect 4255 4964 4259 5015
rect 4060 4963 4073 4964
rect 4125 4963 4138 4964
rect 4190 4963 4203 4964
rect 4255 4963 4268 4964
rect 4320 4963 4326 5015
rect 8554 5079 8560 5131
rect 8612 5079 8627 5131
rect 8679 5079 8694 5131
rect 8746 5079 8761 5131
rect 8813 5079 8828 5131
rect 8880 5079 8895 5131
rect 8947 5079 8962 5131
rect 9014 5079 9028 5131
rect 9080 5079 9094 5131
rect 9146 5079 9160 5131
rect 9212 5128 9226 5131
rect 9278 5079 9292 5131
rect 9344 5128 9358 5131
rect 9410 5128 9424 5131
rect 9476 5128 9490 5131
rect 9542 5128 9556 5131
rect 9608 5128 9614 5131
rect 9352 5079 9358 5128
rect 9542 5079 9550 5128
rect 9608 5079 9634 5128
rect 8554 5072 9211 5079
rect 9267 5072 9296 5079
rect 9352 5072 9381 5079
rect 9437 5072 9466 5079
rect 9522 5072 9550 5079
rect 9606 5072 9634 5079
rect 9690 5072 9718 5128
rect 9774 5072 9783 5128
rect 8554 5020 9783 5072
rect 8554 5015 9211 5020
rect 9267 5015 9296 5020
rect 9352 5015 9381 5020
rect 9437 5015 9466 5020
rect 9522 5015 9550 5020
rect 9606 5015 9634 5020
rect 8554 4963 8560 5015
rect 8612 4963 8627 5015
rect 8679 4963 8694 5015
rect 8746 4963 8761 5015
rect 8813 4963 8828 5015
rect 8880 4963 8895 5015
rect 8947 4963 8962 5015
rect 9014 4963 9028 5015
rect 9080 4963 9094 5015
rect 9146 4963 9160 5015
rect 9212 4963 9226 4964
rect 9278 4963 9292 5015
rect 9352 4964 9358 5015
rect 9542 4964 9550 5015
rect 9608 4964 9634 5015
rect 9690 4964 9718 5020
rect 9774 4964 9783 5020
rect 11008 5079 11014 5131
rect 11066 5128 11082 5131
rect 11134 5128 11150 5131
rect 11202 5128 11217 5131
rect 11074 5079 11082 5128
rect 11202 5079 11209 5128
rect 11269 5079 11275 5131
rect 11008 5072 11018 5079
rect 11074 5072 11114 5079
rect 11170 5072 11209 5079
rect 11265 5072 11275 5079
rect 11008 5020 11275 5072
rect 11008 5015 11018 5020
rect 11074 5015 11114 5020
rect 11170 5015 11209 5020
rect 11265 5015 11275 5020
rect 9344 4963 9358 4964
rect 9410 4963 9424 4964
rect 9476 4963 9490 4964
rect 9542 4963 9556 4964
rect 9608 4963 9614 4964
rect 11008 4963 11014 5015
rect 11074 4964 11082 5015
rect 11202 4964 11209 5015
rect 11066 4963 11082 4964
rect 11134 4963 11150 4964
rect 11202 4963 11217 4964
rect 11269 4963 11275 5015
rect 15043 5079 15049 5131
rect 15101 5128 15118 5131
rect 15170 5128 15187 5131
rect 15239 5128 15255 5131
rect 15307 5128 15323 5131
rect 15375 5128 15391 5131
rect 15443 5128 15459 5131
rect 15511 5128 15527 5131
rect 15579 5128 15595 5131
rect 15647 5128 15663 5131
rect 15715 5128 15731 5131
rect 15783 5128 15799 5131
rect 15851 5128 15867 5131
rect 15109 5079 15118 5128
rect 15375 5079 15377 5128
rect 15443 5079 15458 5128
rect 15514 5079 15527 5128
rect 15851 5079 15859 5128
rect 15919 5079 15925 5131
rect 15043 5072 15053 5079
rect 15109 5072 15134 5079
rect 15190 5072 15215 5079
rect 15271 5072 15296 5079
rect 15352 5072 15377 5079
rect 15433 5072 15458 5079
rect 15514 5072 15539 5079
rect 15595 5072 15619 5079
rect 15675 5072 15699 5079
rect 15755 5072 15779 5079
rect 15835 5072 15859 5079
rect 15915 5072 15925 5079
rect 15043 5020 15925 5072
rect 15043 5015 15053 5020
rect 15109 5015 15134 5020
rect 15190 5015 15215 5020
rect 15271 5015 15296 5020
rect 15352 5015 15377 5020
rect 15433 5015 15458 5020
rect 15514 5015 15539 5020
rect 15595 5015 15619 5020
rect 15675 5015 15699 5020
rect 15755 5015 15779 5020
rect 15835 5015 15859 5020
rect 15915 5015 15925 5020
rect 15043 4963 15049 5015
rect 15109 4964 15118 5015
rect 15375 4964 15377 5015
rect 15443 4964 15458 5015
rect 15514 4964 15527 5015
rect 15851 4964 15859 5015
rect 15101 4963 15118 4964
rect 15170 4963 15187 4964
rect 15239 4963 15255 4964
rect 15307 4963 15323 4964
rect 15375 4963 15391 4964
rect 15443 4963 15459 4964
rect 15511 4963 15527 4964
rect 15579 4963 15595 4964
rect 15647 4963 15663 4964
rect 15715 4963 15731 4964
rect 15783 4963 15799 4964
rect 15851 4963 15867 4964
rect 15919 4963 15925 5015
rect 16882 5079 16888 5131
rect 16940 5128 16957 5131
rect 17009 5128 17026 5131
rect 17078 5128 17094 5131
rect 17146 5128 17162 5131
rect 17214 5128 17230 5131
rect 17282 5128 17298 5131
rect 17350 5128 17366 5131
rect 17418 5128 17434 5131
rect 17486 5128 17502 5131
rect 17554 5128 17570 5131
rect 17622 5128 17638 5131
rect 17690 5128 17706 5131
rect 16948 5079 16957 5128
rect 17214 5079 17216 5128
rect 17282 5079 17297 5128
rect 17353 5079 17366 5128
rect 17690 5079 17698 5128
rect 17758 5079 17764 5131
rect 16882 5072 16892 5079
rect 16948 5072 16973 5079
rect 17029 5072 17054 5079
rect 17110 5072 17135 5079
rect 17191 5072 17216 5079
rect 17272 5072 17297 5079
rect 17353 5072 17378 5079
rect 17434 5072 17458 5079
rect 17514 5072 17538 5079
rect 17594 5072 17618 5079
rect 17674 5072 17698 5079
rect 17754 5072 17764 5079
rect 16882 5020 17764 5072
rect 16882 5015 16892 5020
rect 16948 5015 16973 5020
rect 17029 5015 17054 5020
rect 17110 5015 17135 5020
rect 17191 5015 17216 5020
rect 17272 5015 17297 5020
rect 17353 5015 17378 5020
rect 17434 5015 17458 5020
rect 17514 5015 17538 5020
rect 17594 5015 17618 5020
rect 17674 5015 17698 5020
rect 17754 5015 17764 5020
rect 16882 4963 16888 5015
rect 16948 4964 16957 5015
rect 17214 4964 17216 5015
rect 17282 4964 17297 5015
rect 17353 4964 17366 5015
rect 17690 4964 17698 5015
rect 16940 4963 16957 4964
rect 17009 4963 17026 4964
rect 17078 4963 17094 4964
rect 17146 4963 17162 4964
rect 17214 4963 17230 4964
rect 17282 4963 17298 4964
rect 17350 4963 17366 4964
rect 17418 4963 17434 4964
rect 17486 4963 17502 4964
rect 17554 4963 17570 4964
rect 17622 4963 17638 4964
rect 17690 4963 17706 4964
rect 17758 4963 17764 5015
rect 19665 5079 19671 5131
rect 19723 5128 19762 5131
rect 19665 5072 19675 5079
rect 19731 5072 19755 5128
rect 19814 5079 19820 5131
rect 19811 5072 19820 5079
rect 19665 5020 19820 5072
rect 19665 5015 19675 5020
rect 19665 4963 19671 5015
rect 19731 4964 19755 5020
rect 19811 5015 19820 5020
rect 19723 4963 19762 4964
rect 19814 4963 19820 5015
tri -1168 4694 -1156 4706 se
rect -1156 4694 -1096 4706
tri -1096 4694 -1084 4706 nw
tri -1033 4694 -1021 4706 se
rect -1021 4694 -969 4706
tri -1176 4686 -1168 4694 se
rect -1168 4686 -1104 4694
tri -1104 4686 -1096 4694 nw
tri -1041 4686 -1033 4694 se
rect -1033 4686 -969 4694
rect -1176 4526 -1124 4686
tri -1124 4666 -1104 4686 nw
tri -1061 4666 -1041 4686 se
rect -1041 4666 -1012 4686
rect -1176 4462 -1124 4474
tri -1584 4307 -1572 4319 sw
rect -1636 4275 -1572 4307
tri -1636 4267 -1628 4275 ne
rect -1628 4267 -1572 4275
tri -1628 4263 -1624 4267 ne
tri -1636 3962 -1624 3974 se
rect -1624 3962 -1572 4267
rect -1636 3930 -1572 3962
rect -2090 2645 -1685 2651
rect -2090 2599 -1737 2645
rect -1737 2581 -1685 2593
rect -1737 2523 -1685 2529
rect -2174 2400 -1670 2406
rect -2174 2354 -1722 2400
rect -1722 2336 -1670 2348
rect -1722 2278 -1670 2284
rect -1636 2035 -1584 3930
tri -1584 3918 -1572 3930 nw
tri -1259 3082 -1176 3165 se
rect -1176 3134 -1124 4410
tri -1084 4643 -1061 4666 se
rect -1061 4643 -1012 4666
tri -1012 4643 -969 4686 nw
rect 3625 4706 3631 4758
rect 3683 4706 3698 4758
rect 3750 4706 3765 4758
rect 3817 4706 3832 4758
rect 3884 4706 3899 4758
rect 3951 4706 3966 4758
rect 4018 4706 4033 4758
rect 4085 4706 4099 4758
rect 4151 4706 4165 4758
rect 4217 4706 4223 4758
rect 3625 4694 4223 4706
rect -1084 4642 -1013 4643
tri -1013 4642 -1012 4643 nw
rect 3625 4642 3631 4694
rect 3683 4642 3698 4694
rect 3750 4642 3765 4694
rect 3817 4642 3832 4694
rect 3884 4642 3899 4694
rect 3951 4642 3966 4694
rect 4018 4642 4033 4694
rect 4085 4642 4099 4694
rect 4151 4642 4165 4694
rect 4217 4642 4223 4694
rect -1084 4630 -1025 4642
tri -1025 4630 -1013 4642 nw
rect 3625 4630 4223 4642
rect -1084 4458 -1032 4630
tri -1032 4623 -1025 4630 nw
rect 3625 4578 3631 4630
rect 3683 4578 3698 4630
rect 3750 4578 3765 4630
rect 3817 4578 3832 4630
rect 3884 4578 3899 4630
rect 3951 4578 3966 4630
rect 4018 4578 4033 4630
rect 4085 4578 4099 4630
rect 4151 4578 4165 4630
rect 4217 4578 4223 4630
rect -1084 4406 -1078 4458
rect -1026 4406 -1014 4458
rect -962 4406 -956 4458
rect -1084 3779 -1032 4406
tri 19844 4378 19850 4384 se
rect 19850 4378 19960 5876
tri 22934 4623 22936 4625 se
rect 22936 4623 23046 6046
rect 19844 4372 19960 4378
rect 638 4295 647 4351
rect 703 4347 729 4351
rect 785 4347 811 4351
rect 703 4295 725 4347
rect 785 4295 800 4347
rect 867 4295 892 4351
rect 948 4295 957 4351
rect 638 4267 957 4295
rect 638 4211 647 4267
rect 703 4215 725 4267
rect 785 4215 800 4267
rect 703 4211 729 4215
rect 785 4211 811 4215
rect 867 4211 892 4267
rect 948 4211 957 4267
rect 6012 4347 6021 4351
rect 6077 4347 6103 4351
rect 6159 4347 6184 4351
rect 6240 4347 6265 4351
rect 6321 4347 6346 4351
rect 6402 4347 6411 4351
rect 6012 4295 6018 4347
rect 6077 4295 6085 4347
rect 6338 4295 6346 4347
rect 6405 4295 6411 4347
rect 6012 4267 6411 4295
rect 6012 4215 6018 4267
rect 6077 4215 6085 4267
rect 6338 4215 6346 4267
rect 6405 4215 6411 4267
rect 6012 4211 6021 4215
rect 6077 4211 6103 4215
rect 6159 4211 6184 4215
rect 6240 4211 6265 4215
rect 6321 4211 6346 4215
rect 6402 4211 6411 4215
rect 6943 4347 6952 4351
rect 7008 4347 7034 4351
rect 7090 4347 7115 4351
rect 7171 4347 7196 4351
rect 7252 4347 7277 4351
rect 7333 4347 7342 4351
rect 6943 4295 6949 4347
rect 7008 4295 7016 4347
rect 7269 4295 7277 4347
rect 7336 4295 7342 4347
rect 6943 4267 7342 4295
rect 6943 4215 6949 4267
rect 7008 4215 7016 4267
rect 7269 4215 7277 4267
rect 7336 4215 7342 4267
rect 6943 4211 6952 4215
rect 7008 4211 7034 4215
rect 7090 4211 7115 4215
rect 7171 4211 7196 4215
rect 7252 4211 7277 4215
rect 7333 4211 7342 4215
rect 12496 4347 12505 4351
rect 12561 4347 12587 4351
rect 12643 4347 12668 4351
rect 12724 4347 12749 4351
rect 12805 4347 12830 4351
rect 12886 4347 12895 4351
rect 12496 4295 12502 4347
rect 12561 4295 12569 4347
rect 12822 4295 12830 4347
rect 12889 4295 12895 4347
rect 12496 4267 12895 4295
rect 12496 4215 12502 4267
rect 12561 4215 12569 4267
rect 12822 4215 12830 4267
rect 12889 4215 12895 4267
rect 12496 4211 12505 4215
rect 12561 4211 12587 4215
rect 12643 4211 12668 4215
rect 12724 4211 12749 4215
rect 12805 4211 12830 4215
rect 12886 4211 12895 4215
rect 13427 4347 13436 4351
rect 13492 4347 13518 4351
rect 13574 4347 13599 4351
rect 13655 4347 13680 4351
rect 13736 4347 13761 4351
rect 13817 4347 13826 4351
rect 13427 4295 13433 4347
rect 13492 4295 13500 4347
rect 13753 4295 13761 4347
rect 13820 4295 13826 4347
rect 13427 4267 13826 4295
rect 13427 4215 13433 4267
rect 13492 4215 13500 4267
rect 13753 4215 13761 4267
rect 13820 4215 13826 4267
rect 13427 4211 13436 4215
rect 13492 4211 13518 4215
rect 13574 4211 13599 4215
rect 13655 4211 13680 4215
rect 13736 4211 13761 4215
rect 13817 4211 13826 4215
rect 19061 4347 19070 4351
rect 19061 4295 19067 4347
rect 19126 4295 19152 4351
rect 19208 4295 19233 4351
rect 19289 4295 19314 4351
rect 19370 4347 19379 4351
rect 19373 4295 19379 4347
rect 19061 4267 19379 4295
rect 19061 4215 19067 4267
rect 19061 4211 19070 4215
rect 19126 4211 19152 4267
rect 19208 4211 19233 4267
rect 19289 4211 19314 4267
rect 19373 4215 19379 4267
rect 19370 4211 19379 4215
rect 19844 4186 19960 4192
tri 22930 4619 22934 4623 se
rect 22934 4619 23046 4623
rect -1095 3727 -1032 3779
rect -1095 3454 -1049 3727
rect -1095 3402 -1032 3454
tri -1176 3082 -1124 3134 nw
tri -1318 3023 -1259 3082 se
rect -1259 3023 -1235 3082
tri -1235 3023 -1176 3082 nw
tri -1324 3017 -1318 3023 se
rect -1318 3017 -1241 3023
tri -1241 3017 -1235 3023 nw
tri -1342 2999 -1324 3017 se
rect -1324 2999 -1259 3017
tri -1259 2999 -1241 3017 nw
tri -1360 2981 -1342 2999 se
rect -1342 2981 -1277 2999
tri -1277 2981 -1259 2999 nw
rect -1360 2965 -1293 2981
tri -1293 2965 -1277 2981 nw
rect -1360 2959 -1299 2965
tri -1299 2959 -1293 2965 nw
rect -1360 2953 -1305 2959
tri -1305 2953 -1299 2959 nw
rect -1360 2829 -1308 2953
tri -1308 2950 -1305 2953 nw
rect -1360 2759 -1308 2777
rect -1360 2688 -1308 2707
rect -1360 2630 -1308 2636
rect -1084 2829 -1032 3402
rect -1084 2759 -1032 2777
rect -1084 2688 -1032 2707
rect -1084 2630 -1032 2636
rect -630 3333 -624 3385
rect -572 3333 -560 3385
rect -508 3333 -502 3385
rect -1636 1965 -1584 1983
rect -1636 1894 -1584 1913
rect -1736 1849 -1684 1855
rect -1736 1785 -1684 1797
rect -2422 1733 -1736 1782
rect -2422 1730 -1684 1733
rect -1736 1727 -1684 1730
rect -1636 788 -1584 1842
rect -630 1807 -578 3333
rect -310 3017 -258 3023
rect -310 2953 -258 2965
rect -310 2895 -258 2901
rect 638 2959 647 2963
rect 638 2907 644 2959
rect 703 2907 728 2963
rect 784 2907 808 2963
rect 864 2907 888 2963
rect 944 2959 953 2963
rect 947 2907 953 2959
rect -466 2877 -414 2883
rect -466 2813 -414 2825
rect -466 2755 -414 2761
rect -310 2467 -270 2895
rect 638 2879 953 2907
rect 638 2827 644 2879
rect 638 2823 647 2827
rect 703 2823 728 2879
rect 784 2823 808 2879
rect 864 2823 888 2879
rect 947 2827 953 2879
rect 944 2823 953 2827
rect 6012 2959 6021 2963
rect 6077 2959 6103 2963
rect 6159 2959 6184 2963
rect 6240 2959 6265 2963
rect 6321 2959 6346 2963
rect 6402 2959 6411 2963
rect 6012 2907 6018 2959
rect 6077 2907 6085 2959
rect 6338 2907 6346 2959
rect 6405 2907 6411 2959
rect 6012 2879 6411 2907
rect 6012 2827 6018 2879
rect 6077 2827 6085 2879
rect 6338 2827 6346 2879
rect 6405 2827 6411 2879
rect 6012 2823 6021 2827
rect 6077 2823 6103 2827
rect 6159 2823 6184 2827
rect 6240 2823 6265 2827
rect 6321 2823 6346 2827
rect 6402 2823 6411 2827
rect 6943 2959 6952 2963
rect 7008 2959 7034 2963
rect 7090 2959 7115 2963
rect 7171 2959 7196 2963
rect 7252 2959 7277 2963
rect 7333 2959 7342 2963
rect 6943 2907 6949 2959
rect 7008 2907 7016 2959
rect 7269 2907 7277 2959
rect 7336 2907 7342 2959
rect 6943 2879 7342 2907
rect 6943 2827 6949 2879
rect 7008 2827 7016 2879
rect 7269 2827 7277 2879
rect 7336 2827 7342 2879
rect 6943 2823 6952 2827
rect 7008 2823 7034 2827
rect 7090 2823 7115 2827
rect 7171 2823 7196 2827
rect 7252 2823 7277 2827
rect 7333 2823 7342 2827
rect 12496 2959 12505 2963
rect 12561 2959 12587 2963
rect 12643 2959 12668 2963
rect 12724 2959 12749 2963
rect 12805 2959 12830 2963
rect 12886 2959 12895 2963
rect 12496 2907 12502 2959
rect 12561 2907 12569 2959
rect 12822 2907 12830 2959
rect 12889 2907 12895 2959
rect 12496 2879 12895 2907
rect 12496 2827 12502 2879
rect 12561 2827 12569 2879
rect 12822 2827 12830 2879
rect 12889 2827 12895 2879
rect 12496 2823 12505 2827
rect 12561 2823 12587 2827
rect 12643 2823 12668 2827
rect 12724 2823 12749 2827
rect 12805 2823 12830 2827
rect 12886 2823 12895 2827
rect 13427 2959 13436 2963
rect 13492 2959 13518 2963
rect 13574 2959 13599 2963
rect 13655 2959 13680 2963
rect 13736 2959 13761 2963
rect 13817 2959 13826 2963
rect 13427 2907 13433 2959
rect 13492 2907 13500 2959
rect 13753 2907 13761 2959
rect 13820 2907 13826 2959
rect 13427 2879 13826 2907
rect 13427 2827 13433 2879
rect 13492 2827 13500 2879
rect 13753 2827 13761 2879
rect 13820 2827 13826 2879
rect 13427 2823 13436 2827
rect 13492 2823 13518 2827
rect 13574 2823 13599 2827
rect 13655 2823 13680 2827
rect 13736 2823 13761 2827
rect 13817 2823 13826 2827
rect 19065 2959 19074 2963
rect 19065 2907 19071 2959
rect 19130 2907 19154 2963
rect 19210 2907 19234 2963
rect 19290 2907 19314 2963
rect 19370 2959 19379 2963
rect 19373 2907 19379 2959
rect 19065 2879 19379 2907
rect 19065 2827 19071 2879
rect 19065 2823 19074 2827
rect 19130 2823 19154 2879
rect 19210 2823 19234 2879
rect 19290 2823 19314 2879
rect 19373 2827 19379 2879
rect 19370 2823 19379 2827
rect 638 2686 644 2738
rect 638 2682 647 2686
rect 703 2682 728 2738
rect 784 2682 808 2738
rect 864 2682 888 2738
rect 947 2686 953 2738
rect 944 2682 953 2686
rect 638 2674 953 2682
rect 638 2622 644 2674
rect 696 2622 728 2674
rect 780 2622 812 2674
rect 864 2622 895 2674
rect 947 2622 953 2674
rect 638 2614 953 2622
rect 638 2610 647 2614
rect -222 2567 -170 2573
rect 638 2558 644 2610
rect 703 2558 728 2614
rect 784 2558 808 2614
rect 864 2558 888 2614
rect 944 2610 953 2614
rect 947 2558 953 2610
rect 6012 2686 6018 2738
rect 6077 2686 6085 2738
rect 6338 2686 6346 2738
rect 6405 2686 6411 2738
rect 6012 2682 6021 2686
rect 6077 2682 6102 2686
rect 6158 2682 6183 2686
rect 6239 2682 6264 2686
rect 6320 2682 6346 2686
rect 6402 2682 6411 2686
rect 6012 2674 6411 2682
rect 6012 2622 6018 2674
rect 6070 2622 6085 2674
rect 6137 2622 6152 2674
rect 6204 2622 6219 2674
rect 6271 2622 6286 2674
rect 6338 2622 6353 2674
rect 6405 2622 6411 2674
rect 6012 2614 6411 2622
rect 6012 2610 6021 2614
rect 6077 2610 6102 2614
rect 6158 2610 6183 2614
rect 6239 2610 6264 2614
rect 6320 2610 6346 2614
rect 6402 2610 6411 2614
rect 6012 2558 6018 2610
rect 6077 2558 6085 2610
rect 6338 2558 6346 2610
rect 6405 2558 6411 2610
rect 6943 2686 6949 2738
rect 7008 2686 7016 2738
rect 7269 2686 7277 2738
rect 7336 2686 7342 2738
rect 6943 2682 6952 2686
rect 7008 2682 7034 2686
rect 7090 2682 7115 2686
rect 7171 2682 7196 2686
rect 7252 2682 7277 2686
rect 7333 2682 7342 2686
rect 6943 2674 7342 2682
rect 6943 2622 6949 2674
rect 7001 2622 7016 2674
rect 7068 2622 7083 2674
rect 7135 2622 7150 2674
rect 7202 2622 7217 2674
rect 7269 2622 7284 2674
rect 7336 2622 7342 2674
rect 6943 2614 7342 2622
rect 6943 2610 6952 2614
rect 7008 2610 7034 2614
rect 7090 2610 7115 2614
rect 7171 2610 7196 2614
rect 7252 2610 7277 2614
rect 7333 2610 7342 2614
rect 6943 2558 6949 2610
rect 7008 2558 7016 2610
rect 7269 2558 7277 2610
rect 7336 2558 7342 2610
rect 12496 2686 12502 2738
rect 12561 2686 12569 2738
rect 12822 2686 12830 2738
rect 12889 2686 12895 2738
rect 12496 2682 12505 2686
rect 12561 2682 12586 2686
rect 12642 2682 12667 2686
rect 12723 2682 12748 2686
rect 12804 2682 12830 2686
rect 12886 2682 12895 2686
rect 12496 2674 12895 2682
rect 12496 2622 12502 2674
rect 12554 2622 12569 2674
rect 12621 2622 12636 2674
rect 12688 2622 12703 2674
rect 12755 2622 12770 2674
rect 12822 2622 12837 2674
rect 12889 2622 12895 2674
rect 12496 2614 12895 2622
rect 12496 2610 12505 2614
rect 12561 2610 12586 2614
rect 12642 2610 12667 2614
rect 12723 2610 12748 2614
rect 12804 2610 12830 2614
rect 12886 2610 12895 2614
rect 12496 2558 12502 2610
rect 12561 2558 12569 2610
rect 12822 2558 12830 2610
rect 12889 2558 12895 2610
rect 13427 2686 13433 2738
rect 13492 2686 13500 2738
rect 13753 2686 13761 2738
rect 13820 2686 13826 2738
rect 13427 2682 13436 2686
rect 13492 2682 13518 2686
rect 13574 2682 13599 2686
rect 13655 2682 13680 2686
rect 13736 2682 13761 2686
rect 13817 2682 13826 2686
rect 13427 2674 13826 2682
rect 13427 2622 13433 2674
rect 13485 2622 13500 2674
rect 13552 2622 13567 2674
rect 13619 2622 13634 2674
rect 13686 2622 13701 2674
rect 13753 2622 13768 2674
rect 13820 2622 13826 2674
rect 13427 2614 13826 2622
rect 13427 2610 13436 2614
rect 13492 2610 13518 2614
rect 13574 2610 13599 2614
rect 13655 2610 13680 2614
rect 13736 2610 13761 2614
rect 13817 2610 13826 2614
rect 13427 2558 13433 2610
rect 13492 2558 13500 2610
rect 13753 2558 13761 2610
rect 13820 2558 13826 2610
rect 19065 2686 19071 2738
rect 19065 2682 19074 2686
rect 19130 2682 19154 2738
rect 19210 2682 19234 2738
rect 19290 2682 19314 2738
rect 19373 2686 19379 2738
rect 19370 2682 19379 2686
rect 19065 2674 19379 2682
rect 19065 2622 19071 2674
rect 19123 2622 19154 2674
rect 19206 2622 19237 2674
rect 19289 2622 19321 2674
rect 19373 2622 19379 2674
rect 19065 2614 19379 2622
rect 19065 2610 19074 2614
rect 19065 2558 19071 2610
rect 19130 2558 19154 2614
rect 19210 2558 19234 2614
rect 19290 2558 19314 2614
rect 19370 2610 19379 2614
rect 19373 2558 19379 2610
rect 19065 2553 19379 2558
rect 19065 2538 19364 2553
tri 19364 2538 19379 2553 nw
rect -222 2503 -170 2515
rect -310 2461 -258 2467
rect -310 2397 -258 2409
rect -310 2339 -258 2345
rect -466 2071 -414 2077
rect -466 2007 -414 2019
rect -466 1949 -414 1955
rect -630 1743 -578 1755
rect -630 1503 -578 1691
rect -630 1439 -578 1451
rect -630 870 -578 1387
rect -630 806 -578 818
tri -1636 758 -1606 788 ne
rect -1606 758 -1584 788
tri -1584 758 -1538 804 sw
tri -1606 754 -1602 758 ne
rect -1602 754 -1538 758
tri -1538 754 -1534 758 sw
tri -1602 737 -1585 754 ne
rect -1585 737 -1534 754
tri -1534 737 -1517 754 sw
rect -630 748 -578 754
rect -222 1047 -170 2451
rect 1021 2437 1920 2441
rect 1021 2385 1027 2437
rect 1274 2385 1284 2437
rect 1340 2385 1350 2437
rect 1594 2385 1606 2437
rect 1667 2385 1670 2437
rect 1850 2385 1854 2437
rect 1914 2385 1920 2437
rect 1021 2381 1038 2385
rect 1094 2381 1120 2385
rect 1176 2381 1202 2385
rect 1258 2381 1284 2385
rect 1340 2381 1366 2385
rect 1422 2381 1448 2385
rect 1504 2381 1530 2385
rect 1586 2381 1611 2385
rect 1667 2381 1692 2385
rect 1748 2381 1773 2385
rect 1829 2381 1854 2385
rect 1910 2381 1920 2385
rect 1021 2369 1920 2381
rect 1021 2317 1027 2369
rect 1079 2353 1092 2369
rect 1144 2353 1157 2369
rect 1209 2353 1222 2369
rect 1274 2353 1286 2369
rect 1338 2353 1350 2369
rect 1402 2353 1414 2369
rect 1466 2353 1478 2369
rect 1530 2353 1542 2369
rect 1274 2317 1284 2353
rect 1340 2317 1350 2353
rect 1594 2317 1606 2369
rect 1658 2353 1670 2369
rect 1722 2353 1734 2369
rect 1786 2353 1798 2369
rect 1850 2353 1862 2369
rect 1667 2317 1670 2353
rect 1850 2317 1854 2353
rect 1914 2317 1920 2369
rect 1021 2301 1038 2317
rect 1094 2301 1120 2317
rect 1176 2301 1202 2317
rect 1258 2301 1284 2317
rect 1340 2301 1366 2317
rect 1422 2301 1448 2317
rect 1504 2301 1530 2317
rect 1586 2301 1611 2317
rect 1667 2301 1692 2317
rect 1748 2301 1773 2317
rect 1829 2301 1854 2317
rect 1910 2301 1920 2317
rect 1021 2249 1027 2301
rect 1274 2297 1284 2301
rect 1340 2297 1350 2301
rect 1079 2269 1092 2297
rect 1144 2269 1157 2297
rect 1209 2269 1222 2297
rect 1274 2269 1286 2297
rect 1338 2269 1350 2297
rect 1402 2269 1414 2297
rect 1466 2269 1478 2297
rect 1530 2269 1542 2297
rect 1274 2249 1284 2269
rect 1340 2249 1350 2269
rect 1594 2249 1606 2301
rect 1667 2297 1670 2301
rect 1850 2297 1854 2301
rect 1658 2269 1670 2297
rect 1722 2269 1734 2297
rect 1786 2269 1798 2297
rect 1850 2269 1862 2297
rect 1667 2249 1670 2269
rect 1850 2249 1854 2269
rect 1914 2249 1920 2301
rect 1021 2233 1038 2249
rect 1094 2233 1120 2249
rect 1176 2233 1202 2249
rect 1258 2233 1284 2249
rect 1340 2233 1366 2249
rect 1422 2233 1448 2249
rect 1504 2233 1530 2249
rect 1586 2233 1611 2249
rect 1667 2233 1692 2249
rect 1748 2233 1773 2249
rect 1829 2233 1854 2249
rect 1910 2233 1920 2249
rect 1021 2181 1027 2233
rect 1274 2213 1284 2233
rect 1340 2213 1350 2233
rect 1079 2185 1092 2213
rect 1144 2185 1157 2213
rect 1209 2185 1222 2213
rect 1274 2185 1286 2213
rect 1338 2185 1350 2213
rect 1402 2185 1414 2213
rect 1466 2185 1478 2213
rect 1530 2185 1542 2213
rect 1274 2181 1284 2185
rect 1340 2181 1350 2185
rect 1594 2181 1606 2233
rect 1667 2213 1670 2233
rect 1850 2213 1854 2233
rect 1658 2185 1670 2213
rect 1722 2185 1734 2213
rect 1786 2185 1798 2213
rect 1850 2185 1862 2213
rect 1667 2181 1670 2185
rect 1850 2181 1854 2185
rect 1914 2181 1920 2233
rect 1021 2165 1038 2181
rect 1094 2165 1120 2181
rect 1176 2165 1202 2181
rect 1258 2165 1284 2181
rect 1340 2165 1366 2181
rect 1422 2165 1448 2181
rect 1504 2165 1530 2181
rect 1586 2165 1611 2181
rect 1667 2165 1692 2181
rect 1748 2165 1773 2181
rect 1829 2165 1854 2181
rect 1910 2165 1920 2181
rect 1021 2113 1027 2165
rect 1274 2129 1284 2165
rect 1340 2129 1350 2165
rect 1079 2113 1092 2129
rect 1144 2113 1157 2129
rect 1209 2113 1222 2129
rect 1274 2113 1286 2129
rect 1338 2113 1350 2129
rect 1402 2113 1414 2129
rect 1466 2113 1478 2129
rect 1530 2113 1542 2129
rect 1594 2113 1606 2165
rect 1667 2129 1670 2165
rect 1850 2129 1854 2165
rect 1658 2113 1670 2129
rect 1722 2113 1734 2129
rect 1786 2113 1798 2129
rect 1850 2113 1862 2129
rect 1914 2113 1920 2165
rect 1021 2101 1920 2113
rect 1021 2097 1038 2101
rect 1094 2097 1120 2101
rect 1176 2097 1202 2101
rect 1258 2097 1284 2101
rect 1340 2097 1366 2101
rect 1422 2097 1448 2101
rect 1504 2097 1530 2101
rect 1586 2097 1611 2101
rect 1667 2097 1692 2101
rect 1748 2097 1773 2101
rect 1829 2097 1854 2101
rect 1910 2097 1920 2101
rect 1021 2045 1027 2097
rect 1274 2045 1284 2097
rect 1340 2045 1350 2097
rect 1594 2045 1606 2097
rect 1667 2045 1670 2097
rect 1850 2045 1854 2097
rect 1914 2045 1920 2097
rect 1021 2041 1920 2045
rect 5194 2437 5841 2439
rect 5194 2381 5203 2437
rect 5259 2381 5284 2437
rect 5340 2381 5366 2437
rect 5422 2381 5448 2437
rect 5504 2381 5530 2437
rect 5586 2381 5612 2437
rect 5668 2381 5694 2437
rect 5750 2381 5776 2437
rect 5832 2381 5841 2437
rect 5194 2353 5841 2381
rect 5194 2297 5203 2353
rect 5259 2297 5284 2353
rect 5340 2297 5366 2353
rect 5422 2297 5448 2353
rect 5504 2297 5530 2353
rect 5586 2297 5612 2353
rect 5668 2297 5694 2353
rect 5750 2297 5776 2353
rect 5832 2297 5841 2353
rect 5194 2269 5841 2297
rect 5194 2213 5203 2269
rect 5259 2213 5284 2269
rect 5340 2213 5366 2269
rect 5422 2213 5448 2269
rect 5504 2213 5530 2269
rect 5586 2213 5612 2269
rect 5668 2213 5694 2269
rect 5750 2213 5776 2269
rect 5832 2213 5841 2269
rect 5194 2185 5841 2213
rect 5194 2129 5203 2185
rect 5259 2129 5284 2185
rect 5340 2129 5366 2185
rect 5422 2129 5448 2185
rect 5504 2129 5530 2185
rect 5586 2129 5612 2185
rect 5668 2129 5694 2185
rect 5750 2129 5776 2185
rect 5832 2129 5841 2185
rect 5194 2101 5841 2129
rect 5194 2045 5203 2101
rect 5259 2045 5284 2101
rect 5340 2045 5366 2101
rect 5422 2045 5448 2101
rect 5504 2045 5530 2101
rect 5586 2045 5612 2101
rect 5668 2045 5694 2101
rect 5750 2045 5776 2101
rect 5832 2045 5841 2101
rect 5194 2043 5841 2045
rect 7505 2437 8404 2441
rect 7505 2385 7511 2437
rect 7758 2385 7768 2437
rect 7824 2385 7834 2437
rect 8078 2385 8090 2437
rect 8151 2385 8154 2437
rect 8334 2385 8338 2437
rect 8398 2385 8404 2437
rect 7505 2381 7522 2385
rect 7578 2381 7604 2385
rect 7660 2381 7686 2385
rect 7742 2381 7768 2385
rect 7824 2381 7850 2385
rect 7906 2381 7932 2385
rect 7988 2381 8014 2385
rect 8070 2381 8095 2385
rect 8151 2381 8176 2385
rect 8232 2381 8257 2385
rect 8313 2381 8338 2385
rect 8394 2381 8404 2385
rect 7505 2369 8404 2381
rect 7505 2317 7511 2369
rect 7563 2353 7576 2369
rect 7628 2353 7641 2369
rect 7693 2353 7706 2369
rect 7758 2353 7770 2369
rect 7822 2353 7834 2369
rect 7886 2353 7898 2369
rect 7950 2353 7962 2369
rect 8014 2353 8026 2369
rect 7758 2317 7768 2353
rect 7824 2317 7834 2353
rect 8078 2317 8090 2369
rect 8142 2353 8154 2369
rect 8206 2353 8218 2369
rect 8270 2353 8282 2369
rect 8334 2353 8346 2369
rect 8151 2317 8154 2353
rect 8334 2317 8338 2353
rect 8398 2317 8404 2369
rect 7505 2301 7522 2317
rect 7578 2301 7604 2317
rect 7660 2301 7686 2317
rect 7742 2301 7768 2317
rect 7824 2301 7850 2317
rect 7906 2301 7932 2317
rect 7988 2301 8014 2317
rect 8070 2301 8095 2317
rect 8151 2301 8176 2317
rect 8232 2301 8257 2317
rect 8313 2301 8338 2317
rect 8394 2301 8404 2317
rect 7505 2249 7511 2301
rect 7758 2297 7768 2301
rect 7824 2297 7834 2301
rect 7563 2269 7576 2297
rect 7628 2269 7641 2297
rect 7693 2269 7706 2297
rect 7758 2269 7770 2297
rect 7822 2269 7834 2297
rect 7886 2269 7898 2297
rect 7950 2269 7962 2297
rect 8014 2269 8026 2297
rect 7758 2249 7768 2269
rect 7824 2249 7834 2269
rect 8078 2249 8090 2301
rect 8151 2297 8154 2301
rect 8334 2297 8338 2301
rect 8142 2269 8154 2297
rect 8206 2269 8218 2297
rect 8270 2269 8282 2297
rect 8334 2269 8346 2297
rect 8151 2249 8154 2269
rect 8334 2249 8338 2269
rect 8398 2249 8404 2301
rect 7505 2233 7522 2249
rect 7578 2233 7604 2249
rect 7660 2233 7686 2249
rect 7742 2233 7768 2249
rect 7824 2233 7850 2249
rect 7906 2233 7932 2249
rect 7988 2233 8014 2249
rect 8070 2233 8095 2249
rect 8151 2233 8176 2249
rect 8232 2233 8257 2249
rect 8313 2233 8338 2249
rect 8394 2233 8404 2249
rect 7505 2181 7511 2233
rect 7758 2213 7768 2233
rect 7824 2213 7834 2233
rect 7563 2185 7576 2213
rect 7628 2185 7641 2213
rect 7693 2185 7706 2213
rect 7758 2185 7770 2213
rect 7822 2185 7834 2213
rect 7886 2185 7898 2213
rect 7950 2185 7962 2213
rect 8014 2185 8026 2213
rect 7758 2181 7768 2185
rect 7824 2181 7834 2185
rect 8078 2181 8090 2233
rect 8151 2213 8154 2233
rect 8334 2213 8338 2233
rect 8142 2185 8154 2213
rect 8206 2185 8218 2213
rect 8270 2185 8282 2213
rect 8334 2185 8346 2213
rect 8151 2181 8154 2185
rect 8334 2181 8338 2185
rect 8398 2181 8404 2233
rect 7505 2165 7522 2181
rect 7578 2165 7604 2181
rect 7660 2165 7686 2181
rect 7742 2165 7768 2181
rect 7824 2165 7850 2181
rect 7906 2165 7932 2181
rect 7988 2165 8014 2181
rect 8070 2165 8095 2181
rect 8151 2165 8176 2181
rect 8232 2165 8257 2181
rect 8313 2165 8338 2181
rect 8394 2165 8404 2181
rect 7505 2113 7511 2165
rect 7758 2129 7768 2165
rect 7824 2129 7834 2165
rect 7563 2113 7576 2129
rect 7628 2113 7641 2129
rect 7693 2113 7706 2129
rect 7758 2113 7770 2129
rect 7822 2113 7834 2129
rect 7886 2113 7898 2129
rect 7950 2113 7962 2129
rect 8014 2113 8026 2129
rect 8078 2113 8090 2165
rect 8151 2129 8154 2165
rect 8334 2129 8338 2165
rect 8142 2113 8154 2129
rect 8206 2113 8218 2129
rect 8270 2113 8282 2129
rect 8334 2113 8346 2129
rect 8398 2113 8404 2165
rect 7505 2101 8404 2113
rect 7505 2097 7522 2101
rect 7578 2097 7604 2101
rect 7660 2097 7686 2101
rect 7742 2097 7768 2101
rect 7824 2097 7850 2101
rect 7906 2097 7932 2101
rect 7988 2097 8014 2101
rect 8070 2097 8095 2101
rect 8151 2097 8176 2101
rect 8232 2097 8257 2101
rect 8313 2097 8338 2101
rect 8394 2097 8404 2101
rect 7505 2045 7511 2097
rect 7758 2045 7768 2097
rect 7824 2045 7834 2097
rect 8078 2045 8090 2097
rect 8151 2045 8154 2097
rect 8334 2045 8338 2097
rect 8398 2045 8404 2097
rect 7505 2041 8404 2045
rect 11434 2437 12333 2441
rect 11434 2385 11440 2437
rect 11500 2385 11504 2437
rect 11684 2385 11687 2437
rect 11748 2385 11760 2437
rect 12004 2385 12014 2437
rect 12070 2385 12080 2437
rect 12327 2385 12333 2437
rect 11434 2381 11444 2385
rect 11500 2381 11525 2385
rect 11581 2381 11606 2385
rect 11662 2381 11687 2385
rect 11743 2381 11768 2385
rect 11824 2381 11850 2385
rect 11906 2381 11932 2385
rect 11988 2381 12014 2385
rect 12070 2381 12096 2385
rect 12152 2381 12178 2385
rect 12234 2381 12260 2385
rect 12316 2381 12333 2385
rect 11434 2369 12333 2381
rect 11434 2317 11440 2369
rect 11492 2353 11504 2369
rect 11556 2353 11568 2369
rect 11620 2353 11632 2369
rect 11684 2353 11696 2369
rect 11500 2317 11504 2353
rect 11684 2317 11687 2353
rect 11748 2317 11760 2369
rect 11812 2353 11824 2369
rect 11876 2353 11888 2369
rect 11940 2353 11952 2369
rect 12004 2353 12016 2369
rect 12068 2353 12080 2369
rect 12132 2353 12145 2369
rect 12197 2353 12210 2369
rect 12262 2353 12275 2369
rect 12004 2317 12014 2353
rect 12070 2317 12080 2353
rect 12327 2317 12333 2369
rect 11434 2301 11444 2317
rect 11500 2301 11525 2317
rect 11581 2301 11606 2317
rect 11662 2301 11687 2317
rect 11743 2301 11768 2317
rect 11824 2301 11850 2317
rect 11906 2301 11932 2317
rect 11988 2301 12014 2317
rect 12070 2301 12096 2317
rect 12152 2301 12178 2317
rect 12234 2301 12260 2317
rect 12316 2301 12333 2317
rect 11434 2249 11440 2301
rect 11500 2297 11504 2301
rect 11684 2297 11687 2301
rect 11492 2269 11504 2297
rect 11556 2269 11568 2297
rect 11620 2269 11632 2297
rect 11684 2269 11696 2297
rect 11500 2249 11504 2269
rect 11684 2249 11687 2269
rect 11748 2249 11760 2301
rect 12004 2297 12014 2301
rect 12070 2297 12080 2301
rect 11812 2269 11824 2297
rect 11876 2269 11888 2297
rect 11940 2269 11952 2297
rect 12004 2269 12016 2297
rect 12068 2269 12080 2297
rect 12132 2269 12145 2297
rect 12197 2269 12210 2297
rect 12262 2269 12275 2297
rect 12004 2249 12014 2269
rect 12070 2249 12080 2269
rect 12327 2249 12333 2301
rect 11434 2233 11444 2249
rect 11500 2233 11525 2249
rect 11581 2233 11606 2249
rect 11662 2233 11687 2249
rect 11743 2233 11768 2249
rect 11824 2233 11850 2249
rect 11906 2233 11932 2249
rect 11988 2233 12014 2249
rect 12070 2233 12096 2249
rect 12152 2233 12178 2249
rect 12234 2233 12260 2249
rect 12316 2233 12333 2249
rect 11434 2181 11440 2233
rect 11500 2213 11504 2233
rect 11684 2213 11687 2233
rect 11492 2185 11504 2213
rect 11556 2185 11568 2213
rect 11620 2185 11632 2213
rect 11684 2185 11696 2213
rect 11500 2181 11504 2185
rect 11684 2181 11687 2185
rect 11748 2181 11760 2233
rect 12004 2213 12014 2233
rect 12070 2213 12080 2233
rect 11812 2185 11824 2213
rect 11876 2185 11888 2213
rect 11940 2185 11952 2213
rect 12004 2185 12016 2213
rect 12068 2185 12080 2213
rect 12132 2185 12145 2213
rect 12197 2185 12210 2213
rect 12262 2185 12275 2213
rect 12004 2181 12014 2185
rect 12070 2181 12080 2185
rect 12327 2181 12333 2233
rect 11434 2165 11444 2181
rect 11500 2165 11525 2181
rect 11581 2165 11606 2181
rect 11662 2165 11687 2181
rect 11743 2165 11768 2181
rect 11824 2165 11850 2181
rect 11906 2165 11932 2181
rect 11988 2165 12014 2181
rect 12070 2165 12096 2181
rect 12152 2165 12178 2181
rect 12234 2165 12260 2181
rect 12316 2165 12333 2181
rect 11434 2113 11440 2165
rect 11500 2129 11504 2165
rect 11684 2129 11687 2165
rect 11492 2113 11504 2129
rect 11556 2113 11568 2129
rect 11620 2113 11632 2129
rect 11684 2113 11696 2129
rect 11748 2113 11760 2165
rect 12004 2129 12014 2165
rect 12070 2129 12080 2165
rect 11812 2113 11824 2129
rect 11876 2113 11888 2129
rect 11940 2113 11952 2129
rect 12004 2113 12016 2129
rect 12068 2113 12080 2129
rect 12132 2113 12145 2129
rect 12197 2113 12210 2129
rect 12262 2113 12275 2129
rect 12327 2113 12333 2165
rect 11434 2101 12333 2113
rect 11434 2097 11444 2101
rect 11500 2097 11525 2101
rect 11581 2097 11606 2101
rect 11662 2097 11687 2101
rect 11743 2097 11768 2101
rect 11824 2097 11850 2101
rect 11906 2097 11932 2101
rect 11988 2097 12014 2101
rect 12070 2097 12096 2101
rect 12152 2097 12178 2101
rect 12234 2097 12260 2101
rect 12316 2097 12333 2101
rect 11434 2045 11440 2097
rect 11500 2045 11504 2097
rect 11684 2045 11687 2097
rect 11748 2045 11760 2097
rect 12004 2045 12014 2097
rect 12070 2045 12080 2097
rect 12327 2045 12333 2097
rect 11434 2041 12333 2045
rect 13989 2437 14888 2441
rect 13989 2385 13995 2437
rect 14242 2385 14252 2437
rect 14308 2385 14318 2437
rect 14562 2385 14574 2437
rect 14635 2385 14638 2437
rect 14818 2385 14822 2437
rect 14882 2385 14888 2437
rect 13989 2381 14006 2385
rect 14062 2381 14088 2385
rect 14144 2381 14170 2385
rect 14226 2381 14252 2385
rect 14308 2381 14334 2385
rect 14390 2381 14416 2385
rect 14472 2381 14498 2385
rect 14554 2381 14579 2385
rect 14635 2381 14660 2385
rect 14716 2381 14741 2385
rect 14797 2381 14822 2385
rect 14878 2381 14888 2385
rect 13989 2369 14888 2381
rect 13989 2317 13995 2369
rect 14047 2353 14060 2369
rect 14112 2353 14125 2369
rect 14177 2353 14190 2369
rect 14242 2353 14254 2369
rect 14306 2353 14318 2369
rect 14370 2353 14382 2369
rect 14434 2353 14446 2369
rect 14498 2353 14510 2369
rect 14242 2317 14252 2353
rect 14308 2317 14318 2353
rect 14562 2317 14574 2369
rect 14626 2353 14638 2369
rect 14690 2353 14702 2369
rect 14754 2353 14766 2369
rect 14818 2353 14830 2369
rect 14635 2317 14638 2353
rect 14818 2317 14822 2353
rect 14882 2317 14888 2369
rect 13989 2301 14006 2317
rect 14062 2301 14088 2317
rect 14144 2301 14170 2317
rect 14226 2301 14252 2317
rect 14308 2301 14334 2317
rect 14390 2301 14416 2317
rect 14472 2301 14498 2317
rect 14554 2301 14579 2317
rect 14635 2301 14660 2317
rect 14716 2301 14741 2317
rect 14797 2301 14822 2317
rect 14878 2301 14888 2317
rect 13989 2249 13995 2301
rect 14242 2297 14252 2301
rect 14308 2297 14318 2301
rect 14047 2269 14060 2297
rect 14112 2269 14125 2297
rect 14177 2269 14190 2297
rect 14242 2269 14254 2297
rect 14306 2269 14318 2297
rect 14370 2269 14382 2297
rect 14434 2269 14446 2297
rect 14498 2269 14510 2297
rect 14242 2249 14252 2269
rect 14308 2249 14318 2269
rect 14562 2249 14574 2301
rect 14635 2297 14638 2301
rect 14818 2297 14822 2301
rect 14626 2269 14638 2297
rect 14690 2269 14702 2297
rect 14754 2269 14766 2297
rect 14818 2269 14830 2297
rect 14635 2249 14638 2269
rect 14818 2249 14822 2269
rect 14882 2249 14888 2301
rect 13989 2233 14006 2249
rect 14062 2233 14088 2249
rect 14144 2233 14170 2249
rect 14226 2233 14252 2249
rect 14308 2233 14334 2249
rect 14390 2233 14416 2249
rect 14472 2233 14498 2249
rect 14554 2233 14579 2249
rect 14635 2233 14660 2249
rect 14716 2233 14741 2249
rect 14797 2233 14822 2249
rect 14878 2233 14888 2249
rect 13989 2181 13995 2233
rect 14242 2213 14252 2233
rect 14308 2213 14318 2233
rect 14047 2185 14060 2213
rect 14112 2185 14125 2213
rect 14177 2185 14190 2213
rect 14242 2185 14254 2213
rect 14306 2185 14318 2213
rect 14370 2185 14382 2213
rect 14434 2185 14446 2213
rect 14498 2185 14510 2213
rect 14242 2181 14252 2185
rect 14308 2181 14318 2185
rect 14562 2181 14574 2233
rect 14635 2213 14638 2233
rect 14818 2213 14822 2233
rect 14626 2185 14638 2213
rect 14690 2185 14702 2213
rect 14754 2185 14766 2213
rect 14818 2185 14830 2213
rect 14635 2181 14638 2185
rect 14818 2181 14822 2185
rect 14882 2181 14888 2233
rect 13989 2165 14006 2181
rect 14062 2165 14088 2181
rect 14144 2165 14170 2181
rect 14226 2165 14252 2181
rect 14308 2165 14334 2181
rect 14390 2165 14416 2181
rect 14472 2165 14498 2181
rect 14554 2165 14579 2181
rect 14635 2165 14660 2181
rect 14716 2165 14741 2181
rect 14797 2165 14822 2181
rect 14878 2165 14888 2181
rect 13989 2113 13995 2165
rect 14242 2129 14252 2165
rect 14308 2129 14318 2165
rect 14047 2113 14060 2129
rect 14112 2113 14125 2129
rect 14177 2113 14190 2129
rect 14242 2113 14254 2129
rect 14306 2113 14318 2129
rect 14370 2113 14382 2129
rect 14434 2113 14446 2129
rect 14498 2113 14510 2129
rect 14562 2113 14574 2165
rect 14635 2129 14638 2165
rect 14818 2129 14822 2165
rect 14626 2113 14638 2129
rect 14690 2113 14702 2129
rect 14754 2113 14766 2129
rect 14818 2113 14830 2129
rect 14882 2113 14888 2165
rect 13989 2101 14888 2113
rect 13989 2097 14006 2101
rect 14062 2097 14088 2101
rect 14144 2097 14170 2101
rect 14226 2097 14252 2101
rect 14308 2097 14334 2101
rect 14390 2097 14416 2101
rect 14472 2097 14498 2101
rect 14554 2097 14579 2101
rect 14635 2097 14660 2101
rect 14716 2097 14741 2101
rect 14797 2097 14822 2101
rect 14878 2097 14888 2101
rect 13989 2045 13995 2097
rect 14242 2045 14252 2097
rect 14308 2045 14318 2097
rect 14562 2045 14574 2097
rect 14635 2045 14638 2097
rect 14818 2045 14822 2097
rect 14882 2045 14888 2097
rect 13989 2041 14888 2045
rect 17918 2437 18817 2441
rect 17918 2385 17924 2437
rect 17984 2385 17988 2437
rect 18168 2385 18171 2437
rect 18232 2385 18244 2437
rect 18488 2385 18498 2437
rect 18554 2385 18564 2437
rect 18811 2385 18817 2437
rect 17918 2381 17928 2385
rect 17984 2381 18009 2385
rect 18065 2381 18090 2385
rect 18146 2381 18171 2385
rect 18227 2381 18252 2385
rect 18308 2381 18334 2385
rect 18390 2381 18416 2385
rect 18472 2381 18498 2385
rect 18554 2381 18580 2385
rect 18636 2381 18662 2385
rect 18718 2381 18744 2385
rect 18800 2381 18817 2385
rect 17918 2369 18817 2381
rect 17918 2317 17924 2369
rect 17976 2353 17988 2369
rect 18040 2353 18052 2369
rect 18104 2353 18116 2369
rect 18168 2353 18180 2369
rect 17984 2317 17988 2353
rect 18168 2317 18171 2353
rect 18232 2317 18244 2369
rect 18296 2353 18308 2369
rect 18360 2353 18372 2369
rect 18424 2353 18436 2369
rect 18488 2353 18500 2369
rect 18552 2353 18564 2369
rect 18616 2353 18629 2369
rect 18681 2353 18694 2369
rect 18746 2353 18759 2369
rect 18488 2317 18498 2353
rect 18554 2317 18564 2353
rect 18811 2317 18817 2369
rect 17918 2301 17928 2317
rect 17984 2301 18009 2317
rect 18065 2301 18090 2317
rect 18146 2301 18171 2317
rect 18227 2301 18252 2317
rect 18308 2301 18334 2317
rect 18390 2301 18416 2317
rect 18472 2301 18498 2317
rect 18554 2301 18580 2317
rect 18636 2301 18662 2317
rect 18718 2301 18744 2317
rect 18800 2301 18817 2317
rect 17918 2249 17924 2301
rect 17984 2297 17988 2301
rect 18168 2297 18171 2301
rect 17976 2269 17988 2297
rect 18040 2269 18052 2297
rect 18104 2269 18116 2297
rect 18168 2269 18180 2297
rect 17984 2249 17988 2269
rect 18168 2249 18171 2269
rect 18232 2249 18244 2301
rect 18488 2297 18498 2301
rect 18554 2297 18564 2301
rect 18296 2269 18308 2297
rect 18360 2269 18372 2297
rect 18424 2269 18436 2297
rect 18488 2269 18500 2297
rect 18552 2269 18564 2297
rect 18616 2269 18629 2297
rect 18681 2269 18694 2297
rect 18746 2269 18759 2297
rect 18488 2249 18498 2269
rect 18554 2249 18564 2269
rect 18811 2249 18817 2301
rect 17918 2233 17928 2249
rect 17984 2233 18009 2249
rect 18065 2233 18090 2249
rect 18146 2233 18171 2249
rect 18227 2233 18252 2249
rect 18308 2233 18334 2249
rect 18390 2233 18416 2249
rect 18472 2233 18498 2249
rect 18554 2233 18580 2249
rect 18636 2233 18662 2249
rect 18718 2233 18744 2249
rect 18800 2233 18817 2249
rect 17918 2181 17924 2233
rect 17984 2213 17988 2233
rect 18168 2213 18171 2233
rect 17976 2185 17988 2213
rect 18040 2185 18052 2213
rect 18104 2185 18116 2213
rect 18168 2185 18180 2213
rect 17984 2181 17988 2185
rect 18168 2181 18171 2185
rect 18232 2181 18244 2233
rect 18488 2213 18498 2233
rect 18554 2213 18564 2233
rect 18296 2185 18308 2213
rect 18360 2185 18372 2213
rect 18424 2185 18436 2213
rect 18488 2185 18500 2213
rect 18552 2185 18564 2213
rect 18616 2185 18629 2213
rect 18681 2185 18694 2213
rect 18746 2185 18759 2213
rect 18488 2181 18498 2185
rect 18554 2181 18564 2185
rect 18811 2181 18817 2233
rect 17918 2165 17928 2181
rect 17984 2165 18009 2181
rect 18065 2165 18090 2181
rect 18146 2165 18171 2181
rect 18227 2165 18252 2181
rect 18308 2165 18334 2181
rect 18390 2165 18416 2181
rect 18472 2165 18498 2181
rect 18554 2165 18580 2181
rect 18636 2165 18662 2181
rect 18718 2165 18744 2181
rect 18800 2165 18817 2181
rect 17918 2113 17924 2165
rect 17984 2129 17988 2165
rect 18168 2129 18171 2165
rect 17976 2113 17988 2129
rect 18040 2113 18052 2129
rect 18104 2113 18116 2129
rect 18168 2113 18180 2129
rect 18232 2113 18244 2165
rect 18488 2129 18498 2165
rect 18554 2129 18564 2165
rect 18296 2113 18308 2129
rect 18360 2113 18372 2129
rect 18424 2113 18436 2129
rect 18488 2113 18500 2129
rect 18552 2113 18564 2129
rect 18616 2113 18629 2129
rect 18681 2113 18694 2129
rect 18746 2113 18759 2129
rect 18811 2113 18817 2165
rect 17918 2101 18817 2113
rect 17918 2097 17928 2101
rect 17984 2097 18009 2101
rect 18065 2097 18090 2101
rect 18146 2097 18171 2101
rect 18227 2097 18252 2101
rect 18308 2097 18334 2101
rect 18390 2097 18416 2101
rect 18472 2097 18498 2101
rect 18554 2097 18580 2101
rect 18636 2097 18662 2101
rect 18718 2097 18744 2101
rect 18800 2097 18817 2101
rect 17918 2045 17924 2097
rect 17984 2045 17988 2097
rect 18168 2045 18171 2097
rect 18232 2045 18244 2097
rect 18488 2045 18498 2097
rect 18554 2045 18564 2097
rect 18811 2045 18817 2097
rect 17918 2041 18817 2045
rect 638 1867 644 1919
rect 638 1863 647 1867
rect 703 1863 728 1919
rect 784 1863 808 1919
rect 864 1863 888 1919
rect 947 1867 953 1919
rect 944 1863 953 1867
rect 638 1855 953 1863
rect 638 1803 644 1855
rect 696 1803 728 1855
rect 780 1803 812 1855
rect 864 1803 895 1855
rect 947 1803 953 1855
rect 638 1795 953 1803
rect 638 1791 647 1795
rect 638 1739 644 1791
rect 703 1739 728 1795
rect 784 1739 808 1795
rect 864 1739 888 1795
rect 944 1791 953 1795
rect 947 1739 953 1791
rect 6012 1867 6018 1919
rect 6077 1867 6085 1919
rect 6338 1867 6346 1919
rect 6405 1867 6411 1919
rect 6012 1863 6021 1867
rect 6077 1863 6102 1867
rect 6158 1863 6183 1867
rect 6239 1863 6264 1867
rect 6320 1863 6346 1867
rect 6402 1863 6411 1867
rect 6012 1855 6411 1863
rect 6012 1803 6018 1855
rect 6070 1803 6085 1855
rect 6137 1803 6152 1855
rect 6204 1803 6219 1855
rect 6271 1803 6286 1855
rect 6338 1803 6353 1855
rect 6405 1803 6411 1855
rect 6012 1795 6411 1803
rect 6012 1791 6021 1795
rect 6077 1791 6102 1795
rect 6158 1791 6183 1795
rect 6239 1791 6264 1795
rect 6320 1791 6346 1795
rect 6402 1791 6411 1795
rect 6012 1739 6018 1791
rect 6077 1739 6085 1791
rect 6338 1739 6346 1791
rect 6405 1739 6411 1791
rect 6943 1867 6949 1919
rect 7008 1867 7016 1919
rect 7269 1867 7277 1919
rect 7336 1867 7342 1919
rect 6943 1863 6952 1867
rect 7008 1863 7034 1867
rect 7090 1863 7115 1867
rect 7171 1863 7196 1867
rect 7252 1863 7277 1867
rect 7333 1863 7342 1867
rect 6943 1855 7342 1863
rect 6943 1803 6949 1855
rect 7001 1803 7016 1855
rect 7068 1803 7083 1855
rect 7135 1803 7150 1855
rect 7202 1803 7217 1855
rect 7269 1803 7284 1855
rect 7336 1803 7342 1855
rect 6943 1795 7342 1803
rect 6943 1791 6952 1795
rect 7008 1791 7034 1795
rect 7090 1791 7115 1795
rect 7171 1791 7196 1795
rect 7252 1791 7277 1795
rect 7333 1791 7342 1795
rect 6943 1739 6949 1791
rect 7008 1739 7016 1791
rect 7269 1739 7277 1791
rect 7336 1739 7342 1791
rect 12496 1867 12502 1919
rect 12561 1867 12569 1919
rect 12822 1867 12830 1919
rect 12889 1867 12895 1919
rect 12496 1863 12505 1867
rect 12561 1863 12586 1867
rect 12642 1863 12667 1867
rect 12723 1863 12748 1867
rect 12804 1863 12830 1867
rect 12886 1863 12895 1867
rect 12496 1855 12895 1863
rect 12496 1803 12502 1855
rect 12554 1803 12569 1855
rect 12621 1803 12636 1855
rect 12688 1803 12703 1855
rect 12755 1803 12770 1855
rect 12822 1803 12837 1855
rect 12889 1803 12895 1855
rect 12496 1795 12895 1803
rect 12496 1791 12505 1795
rect 12561 1791 12586 1795
rect 12642 1791 12667 1795
rect 12723 1791 12748 1795
rect 12804 1791 12830 1795
rect 12886 1791 12895 1795
rect 12496 1739 12502 1791
rect 12561 1739 12569 1791
rect 12822 1739 12830 1791
rect 12889 1739 12895 1791
rect 13427 1867 13433 1919
rect 13492 1867 13500 1919
rect 13753 1867 13761 1919
rect 13820 1867 13826 1919
rect 13427 1863 13436 1867
rect 13492 1863 13518 1867
rect 13574 1863 13599 1867
rect 13655 1863 13680 1867
rect 13736 1863 13761 1867
rect 13817 1863 13826 1867
rect 13427 1855 13826 1863
rect 13427 1803 13433 1855
rect 13485 1803 13500 1855
rect 13552 1803 13567 1855
rect 13619 1803 13634 1855
rect 13686 1803 13701 1855
rect 13753 1803 13768 1855
rect 13820 1803 13826 1855
rect 13427 1795 13826 1803
rect 13427 1791 13436 1795
rect 13492 1791 13518 1795
rect 13574 1791 13599 1795
rect 13655 1791 13680 1795
rect 13736 1791 13761 1795
rect 13817 1791 13826 1795
rect 13427 1739 13433 1791
rect 13492 1739 13500 1791
rect 13753 1739 13761 1791
rect 13820 1739 13826 1791
rect 19065 1867 19071 1919
rect 19065 1863 19074 1867
rect 19130 1863 19154 1919
rect 19210 1863 19234 1919
rect 19290 1863 19314 1919
rect 19373 1867 19379 1919
rect 19370 1863 19379 1867
rect 19065 1855 19379 1863
rect 19065 1803 19071 1855
rect 19123 1803 19154 1855
rect 19206 1803 19237 1855
rect 19289 1803 19321 1855
rect 19373 1803 19379 1855
rect 19065 1795 19379 1803
rect 19065 1791 19074 1795
rect 19065 1739 19071 1791
rect 19130 1739 19154 1795
rect 19210 1739 19234 1795
rect 19290 1739 19314 1795
rect 19370 1791 19379 1795
rect 19373 1739 19379 1791
rect 2671 1685 3601 1686
rect 2671 1633 2677 1685
rect 2729 1682 2744 1685
rect 2796 1682 2811 1685
rect 2863 1682 2878 1685
rect 2930 1682 2945 1685
rect 2736 1633 2744 1682
rect 2930 1633 2938 1682
rect 2997 1633 3012 1685
rect 3064 1682 3079 1685
rect 3131 1682 3146 1685
rect 3198 1682 3213 1685
rect 3265 1633 3279 1685
rect 3331 1682 3345 1685
rect 3397 1682 3411 1685
rect 3463 1682 3477 1685
rect 3529 1682 3543 1685
rect 3337 1633 3345 1682
rect 3529 1633 3536 1682
rect 3595 1633 3601 1685
rect 2671 1626 2680 1633
rect 2736 1626 2766 1633
rect 2822 1626 2852 1633
rect 2908 1626 2938 1633
rect 2994 1626 3024 1633
rect 3080 1626 3110 1633
rect 3166 1626 3196 1633
rect 3252 1626 3281 1633
rect 3337 1626 3366 1633
rect 3422 1626 3451 1633
rect 3507 1626 3536 1633
rect 3592 1626 3601 1633
rect 2671 1613 3601 1626
rect 2671 1561 2677 1613
rect 2729 1561 2744 1613
rect 2796 1561 2811 1613
rect 2863 1561 2878 1613
rect 2930 1561 2945 1613
rect 2997 1561 3012 1613
rect 3064 1561 3079 1613
rect 3131 1561 3146 1613
rect 3198 1561 3213 1613
rect 3265 1561 3279 1613
rect 3331 1561 3345 1613
rect 3397 1561 3411 1613
rect 3463 1561 3477 1613
rect 3529 1561 3543 1613
rect 3595 1561 3601 1613
rect 2671 1548 3601 1561
rect 2671 1541 2680 1548
rect 2736 1541 2766 1548
rect 2822 1541 2852 1548
rect 2908 1541 2938 1548
rect 2994 1541 3024 1548
rect 3080 1541 3110 1548
rect 3166 1541 3196 1548
rect 3252 1541 3281 1548
rect 3337 1541 3366 1548
rect 3422 1541 3451 1548
rect 3507 1541 3536 1548
rect 3592 1541 3601 1548
rect -132 1532 228 1538
rect -80 1480 228 1532
rect 2671 1489 2677 1541
rect 2736 1492 2744 1541
rect 2930 1492 2938 1541
rect 2729 1489 2744 1492
rect 2796 1489 2811 1492
rect 2863 1489 2878 1492
rect 2930 1489 2945 1492
rect 2997 1489 3012 1541
rect 3064 1489 3079 1492
rect 3131 1489 3146 1492
rect 3198 1489 3213 1492
rect 3265 1489 3279 1541
rect 3337 1492 3345 1541
rect 3529 1492 3536 1541
rect 3331 1489 3345 1492
rect 3397 1489 3411 1492
rect 3463 1489 3477 1492
rect 3529 1489 3543 1492
rect 3595 1489 3601 1541
rect 2671 1488 3601 1489
rect 4876 1685 5117 1686
rect 4876 1633 4882 1685
rect 4934 1682 4971 1685
rect 5023 1682 5059 1685
rect 4876 1626 4885 1633
rect 4941 1626 4969 1682
rect 5025 1626 5052 1682
rect 5111 1633 5117 1685
rect 5714 1685 5936 1686
rect 5714 1682 5720 1685
rect 5772 1682 5799 1685
rect 5108 1626 5117 1633
rect 4876 1613 5117 1626
rect 4876 1561 4882 1613
rect 4934 1561 4971 1613
rect 5023 1561 5059 1613
rect 5111 1561 5117 1613
rect 4876 1548 5117 1561
rect 4876 1541 4885 1548
rect 4876 1489 4882 1541
rect 4941 1492 4969 1548
rect 5025 1492 5052 1548
rect 5108 1541 5117 1548
rect 4934 1489 4971 1492
rect 5023 1489 5059 1492
rect 5111 1489 5117 1541
rect 5713 1633 5720 1682
rect 5778 1633 5799 1682
rect 5851 1682 5878 1685
rect 5851 1633 5871 1682
rect 5930 1633 5936 1685
rect 5713 1626 5722 1633
rect 5778 1626 5871 1633
rect 5927 1626 5936 1633
rect 5713 1613 5936 1626
rect 5713 1561 5720 1613
rect 5772 1561 5799 1613
rect 5851 1561 5878 1613
rect 5930 1561 5936 1613
rect 5713 1548 5936 1561
rect 5713 1541 5722 1548
rect 5778 1541 5871 1548
rect 5927 1541 5936 1548
rect 5713 1492 5720 1541
rect 5778 1492 5799 1541
rect 4876 1488 5117 1489
rect 5714 1489 5720 1492
rect 5772 1489 5799 1492
rect 5851 1492 5871 1541
rect 5851 1489 5878 1492
rect 5930 1489 5936 1541
rect 6487 1630 6496 1686
rect 6552 1685 6598 1686
rect 6654 1685 6700 1686
rect 6756 1685 6802 1686
rect 6552 1633 6574 1685
rect 6780 1633 6802 1685
rect 6552 1630 6598 1633
rect 6654 1630 6700 1633
rect 6756 1630 6802 1633
rect 6858 1630 6867 1686
rect 6487 1613 6867 1630
rect 6487 1561 6497 1613
rect 6549 1561 6574 1613
rect 6626 1561 6651 1613
rect 6703 1561 6728 1613
rect 6780 1561 6805 1613
rect 6857 1561 6867 1613
rect 6487 1552 6867 1561
rect 6487 1496 6496 1552
rect 6552 1541 6598 1552
rect 6654 1541 6700 1552
rect 6756 1541 6802 1552
rect 6552 1496 6574 1541
rect 6780 1496 6802 1541
rect 6858 1496 6867 1552
rect 9519 1685 9784 1686
rect 9519 1633 9525 1685
rect 9577 1682 9592 1685
rect 9644 1682 9659 1685
rect 9711 1682 9726 1685
rect 9584 1633 9592 1682
rect 9711 1633 9719 1682
rect 9778 1633 9784 1685
rect 9519 1626 9528 1633
rect 9584 1626 9624 1633
rect 9680 1626 9719 1633
rect 9775 1626 9784 1633
rect 9519 1613 9784 1626
rect 9519 1561 9525 1613
rect 9577 1561 9592 1613
rect 9644 1561 9659 1613
rect 9711 1561 9726 1613
rect 9778 1561 9784 1613
rect 9519 1548 9784 1561
rect 9519 1541 9528 1548
rect 9584 1541 9624 1548
rect 9680 1541 9719 1548
rect 9775 1541 9784 1548
rect 5714 1488 5936 1489
rect 6491 1489 6497 1496
rect 6549 1489 6574 1496
rect 6626 1489 6651 1496
rect 6703 1489 6728 1496
rect 6780 1489 6805 1496
rect 6857 1489 6863 1496
rect 6491 1488 6863 1489
rect 9519 1489 9525 1541
rect 9584 1492 9592 1541
rect 9711 1492 9719 1541
rect 9577 1489 9592 1492
rect 9644 1489 9659 1492
rect 9711 1489 9726 1492
rect 9778 1489 9784 1541
rect 16397 1685 16799 1686
rect 16397 1633 16403 1685
rect 16455 1682 16471 1685
rect 16523 1682 16539 1685
rect 16591 1682 16607 1685
rect 16659 1682 16674 1685
rect 16726 1682 16741 1685
rect 16462 1633 16471 1682
rect 16726 1633 16734 1682
rect 16793 1633 16799 1685
rect 16397 1626 16406 1633
rect 16462 1626 16488 1633
rect 16544 1626 16570 1633
rect 16626 1626 16652 1633
rect 16708 1626 16734 1633
rect 16790 1626 16799 1633
rect 16397 1613 16799 1626
rect 16397 1561 16403 1613
rect 16455 1561 16471 1613
rect 16523 1561 16539 1613
rect 16591 1561 16607 1613
rect 16659 1561 16674 1613
rect 16726 1561 16741 1613
rect 16793 1561 16799 1613
rect 16397 1548 16799 1561
rect 16397 1541 16406 1548
rect 16462 1541 16488 1548
rect 16544 1541 16570 1548
rect 16626 1541 16652 1548
rect 16708 1541 16734 1548
rect 16790 1541 16799 1548
rect 9519 1488 9784 1489
rect 9897 1490 9949 1496
rect -132 1468 228 1480
rect -80 1439 228 1468
rect -80 1416 176 1439
rect -132 1410 176 1416
tri 119 1387 142 1410 ne
rect 142 1387 176 1410
rect 3370 1403 3376 1455
rect 3428 1403 3440 1455
rect 3492 1438 3808 1455
tri 3808 1438 3825 1455 sw
rect 16397 1489 16403 1541
rect 16462 1492 16471 1541
rect 16726 1492 16734 1541
rect 16455 1489 16471 1492
rect 16523 1489 16539 1492
rect 16591 1489 16607 1492
rect 16659 1489 16674 1492
rect 16726 1489 16741 1492
rect 16793 1489 16799 1541
rect 16397 1488 16799 1489
rect 3492 1427 3825 1438
tri 3825 1427 3836 1438 sw
rect 3492 1403 3836 1427
tri 142 1375 154 1387 ne
rect 154 1375 228 1387
tri 3745 1375 3773 1403 ne
rect 3773 1375 3836 1403
rect 9897 1426 9949 1438
tri 154 1353 176 1375 ne
rect 176 1317 228 1323
rect 1021 1371 1920 1375
tri 3773 1374 3774 1375 ne
rect 3774 1374 3836 1375
tri 3774 1371 3777 1374 ne
rect 3777 1371 3836 1374
rect 1021 1319 1027 1371
rect 1274 1319 1284 1371
rect 1340 1319 1350 1371
rect 1594 1319 1606 1371
rect 1667 1319 1670 1371
rect 1850 1319 1854 1371
rect 1914 1319 1920 1371
tri 3777 1355 3793 1371 ne
rect 1021 1315 1038 1319
rect 1094 1315 1120 1319
rect 1176 1315 1202 1319
rect 1258 1315 1284 1319
rect 1340 1315 1366 1319
rect 1422 1315 1448 1319
rect 1504 1315 1530 1319
rect 1586 1315 1611 1319
rect 1667 1315 1692 1319
rect 1748 1315 1773 1319
rect 1829 1315 1854 1319
rect 1910 1315 1920 1319
rect 1021 1303 1920 1315
rect 1021 1251 1027 1303
rect 1079 1287 1092 1303
rect 1144 1287 1157 1303
rect 1209 1287 1222 1303
rect 1274 1287 1286 1303
rect 1338 1287 1350 1303
rect 1402 1287 1414 1303
rect 1466 1287 1478 1303
rect 1530 1287 1542 1303
rect 1274 1251 1284 1287
rect 1340 1251 1350 1287
rect 1594 1251 1606 1303
rect 1658 1287 1670 1303
rect 1722 1287 1734 1303
rect 1786 1287 1798 1303
rect 1850 1287 1862 1303
rect 1667 1251 1670 1287
rect 1850 1251 1854 1287
rect 1914 1251 1920 1303
rect 1021 1235 1038 1251
rect 1094 1235 1120 1251
rect 1176 1235 1202 1251
rect 1258 1235 1284 1251
rect 1340 1235 1366 1251
rect 1422 1235 1448 1251
rect 1504 1235 1530 1251
rect 1586 1235 1611 1251
rect 1667 1235 1692 1251
rect 1748 1235 1773 1251
rect 1829 1235 1854 1251
rect 1910 1235 1920 1251
rect 1021 1183 1027 1235
rect 1274 1231 1284 1235
rect 1340 1231 1350 1235
rect 1079 1203 1092 1231
rect 1144 1203 1157 1231
rect 1209 1203 1222 1231
rect 1274 1203 1286 1231
rect 1338 1203 1350 1231
rect 1402 1203 1414 1231
rect 1466 1203 1478 1231
rect 1530 1203 1542 1231
rect 1274 1183 1284 1203
rect 1340 1183 1350 1203
rect 1594 1183 1606 1235
rect 1667 1231 1670 1235
rect 1850 1231 1854 1235
rect 1658 1203 1670 1231
rect 1722 1203 1734 1231
rect 1786 1203 1798 1231
rect 1850 1203 1862 1231
rect 1667 1183 1670 1203
rect 1850 1183 1854 1203
rect 1914 1183 1920 1235
rect 1021 1167 1038 1183
rect 1094 1167 1120 1183
rect 1176 1167 1202 1183
rect 1258 1167 1284 1183
rect 1340 1167 1366 1183
rect 1422 1167 1448 1183
rect 1504 1167 1530 1183
rect 1586 1167 1611 1183
rect 1667 1167 1692 1183
rect 1748 1167 1773 1183
rect 1829 1167 1854 1183
rect 1910 1167 1920 1183
rect 1021 1115 1027 1167
rect 1274 1147 1284 1167
rect 1340 1147 1350 1167
rect 1079 1119 1092 1147
rect 1144 1119 1157 1147
rect 1209 1119 1222 1147
rect 1274 1119 1286 1147
rect 1338 1119 1350 1147
rect 1402 1119 1414 1147
rect 1466 1119 1478 1147
rect 1530 1119 1542 1147
rect 1274 1115 1284 1119
rect 1340 1115 1350 1119
rect 1594 1115 1606 1167
rect 1667 1147 1670 1167
rect 1850 1147 1854 1167
rect 1658 1119 1670 1147
rect 1722 1119 1734 1147
rect 1786 1119 1798 1147
rect 1850 1119 1862 1147
rect 1667 1115 1670 1119
rect 1850 1115 1854 1119
rect 1914 1115 1920 1167
rect 1021 1099 1038 1115
rect 1094 1099 1120 1115
rect 1176 1099 1202 1115
rect 1258 1099 1284 1115
rect 1340 1099 1366 1115
rect 1422 1099 1448 1115
rect 1504 1099 1530 1115
rect 1586 1099 1611 1115
rect 1667 1099 1692 1115
rect 1748 1099 1773 1115
rect 1829 1099 1854 1115
rect 1910 1099 1920 1115
tri -170 1047 -157 1060 sw
rect 1021 1047 1027 1099
rect 1274 1063 1284 1099
rect 1340 1063 1350 1099
rect 1079 1047 1092 1063
rect 1144 1047 1157 1063
rect 1209 1047 1222 1063
rect 1274 1047 1286 1063
rect 1338 1047 1350 1063
rect 1402 1047 1414 1063
rect 1466 1047 1478 1063
rect 1530 1047 1542 1063
rect 1594 1047 1606 1099
rect 1667 1063 1670 1099
rect 1850 1063 1854 1099
rect 1658 1047 1670 1063
rect 1722 1047 1734 1063
rect 1786 1047 1798 1063
rect 1850 1047 1862 1063
rect 1914 1047 1920 1099
rect -222 1031 -157 1047
tri -157 1031 -141 1047 sw
rect 1021 1035 1920 1047
rect 1021 1031 1038 1035
rect 1094 1031 1120 1035
rect 1176 1031 1202 1035
rect 1258 1031 1284 1035
rect 1340 1031 1366 1035
rect 1422 1031 1448 1035
rect 1504 1031 1530 1035
rect 1586 1031 1611 1035
rect 1667 1031 1692 1035
rect 1748 1031 1773 1035
rect 1829 1031 1854 1035
rect 1910 1031 1920 1035
rect -222 1026 -141 1031
tri -141 1026 -136 1031 sw
rect -222 1020 228 1026
rect -222 977 176 1020
rect -222 968 -148 977
tri -148 968 -139 977 nw
tri 135 968 144 977 ne
rect 144 968 176 977
rect 1021 979 1027 1031
rect 1274 979 1284 1031
rect 1340 979 1350 1031
rect 1594 979 1606 1031
rect 1667 979 1670 1031
rect 1850 979 1854 1031
rect 1914 979 1920 1031
rect 1021 975 1920 979
rect -222 963 -153 968
tri -153 963 -148 968 nw
tri 144 963 149 968 ne
rect 149 963 228 968
rect -222 956 -160 963
tri -160 956 -153 963 nw
tri 149 956 156 963 ne
rect 156 956 228 963
tri -1585 736 -1584 737 ne
rect -1584 736 -1517 737
tri -1584 727 -1575 736 ne
rect -1575 727 -1517 736
tri -1517 727 -1507 737 sw
rect -222 735 -170 956
tri -170 946 -160 956 nw
tri 156 946 166 956 ne
rect 166 946 176 956
tri 166 936 176 946 ne
rect 176 898 228 904
rect -222 727 -86 735
tri -1575 690 -1538 727 ne
rect -1538 690 -1507 727
tri -1507 690 -1470 727 sw
tri -1538 675 -1523 690 ne
rect -1523 675 -1470 690
tri -1470 675 -1455 690 sw
rect -170 675 -86 727
tri -1523 665 -1513 675 ne
rect -1513 665 -1455 675
tri -1455 665 -1445 675 sw
tri -1513 663 -1511 665 ne
rect -1511 663 -1445 665
tri -1445 663 -1443 665 sw
rect -222 663 -86 675
tri -1511 622 -1470 663 ne
rect -1470 622 -1443 663
tri -1443 622 -1402 663 sw
tri -1470 611 -1459 622 ne
rect -1459 611 -1402 622
tri -1402 611 -1391 622 sw
rect -170 611 -86 663
tri -1459 563 -1411 611 ne
rect -1411 605 -1391 611
tri -1391 605 -1385 611 sw
rect -222 605 -86 611
rect -1411 585 -1385 605
tri -1385 585 -1365 605 sw
tri -158 585 -138 605 ne
rect -1411 563 -1365 585
tri -1365 563 -1343 585 sw
tri -1411 554 -1402 563 ne
rect -1402 554 -1343 563
tri -1343 554 -1334 563 sw
tri -1402 551 -1399 554 ne
rect -1399 551 -1334 554
tri -1334 551 -1331 554 sw
tri -1399 547 -1395 551 ne
rect -1395 547 -1331 551
tri -1331 547 -1327 551 sw
tri -1395 495 -1343 547 ne
rect -1343 495 -1327 547
tri -1327 495 -1275 547 sw
tri -1343 486 -1334 495 ne
rect -1334 486 -1275 495
tri -1275 486 -1266 495 sw
tri -1334 479 -1327 486 ne
rect -1327 479 -861 486
tri -861 479 -854 486 sw
tri -1327 472 -1320 479 ne
rect -1320 472 -854 479
tri -854 472 -847 479 sw
tri -1320 432 -1280 472 ne
rect -1280 432 -847 472
tri -933 427 -928 432 ne
rect -928 427 -847 432
tri -928 411 -912 427 ne
rect -912 411 -847 427
tri -912 398 -899 411 ne
tri -967 -1926 -899 -1858 se
rect -899 -1874 -847 411
rect -138 275 -86 605
rect 1021 547 1920 551
rect 1021 495 1027 547
rect 1274 495 1284 547
rect 1340 495 1350 547
rect 1594 495 1606 547
rect 1667 495 1670 547
rect 1850 495 1854 547
rect 1914 495 1920 547
rect 1021 491 1038 495
rect 1094 491 1120 495
rect 1176 491 1202 495
rect 1258 491 1284 495
rect 1340 491 1366 495
rect 1422 491 1448 495
rect 1504 491 1530 495
rect 1586 491 1611 495
rect 1667 491 1692 495
rect 1748 491 1773 495
rect 1829 491 1854 495
rect 1910 491 1920 495
rect 1021 479 1920 491
rect 1021 427 1027 479
rect 1079 463 1092 479
rect 1144 463 1157 479
rect 1209 463 1222 479
rect 1274 463 1286 479
rect 1338 463 1350 479
rect 1402 463 1414 479
rect 1466 463 1478 479
rect 1530 463 1542 479
rect 1274 427 1284 463
rect 1340 427 1350 463
rect 1594 427 1606 479
rect 1658 463 1670 479
rect 1722 463 1734 479
rect 1786 463 1798 479
rect 1850 463 1862 479
rect 1667 427 1670 463
rect 1850 427 1854 463
rect 1914 427 1920 479
rect 1021 411 1038 427
rect 1094 411 1120 427
rect 1176 411 1202 427
rect 1258 411 1284 427
rect 1340 411 1366 427
rect 1422 411 1448 427
rect 1504 411 1530 427
rect 1586 411 1611 427
rect 1667 411 1692 427
rect 1748 411 1773 427
rect 1829 411 1854 427
rect 1910 411 1920 427
rect 1021 359 1027 411
rect 1274 407 1284 411
rect 1340 407 1350 411
rect 1079 379 1092 407
rect 1144 379 1157 407
rect 1209 379 1222 407
rect 1274 379 1286 407
rect 1338 379 1350 407
rect 1402 379 1414 407
rect 1466 379 1478 407
rect 1530 379 1542 407
rect 1274 359 1284 379
rect 1340 359 1350 379
rect 1594 359 1606 411
rect 1667 407 1670 411
rect 1850 407 1854 411
rect 1658 379 1670 407
rect 1722 379 1734 407
rect 1786 379 1798 407
rect 1850 379 1862 407
rect 1667 359 1670 379
rect 1850 359 1854 379
rect 1914 359 1920 411
rect 1021 343 1038 359
rect 1094 343 1120 359
rect 1176 343 1202 359
rect 1258 343 1284 359
rect 1340 343 1366 359
rect 1422 343 1448 359
rect 1504 343 1530 359
rect 1586 343 1611 359
rect 1667 343 1692 359
rect 1748 343 1773 359
rect 1829 343 1854 359
rect 1910 343 1920 359
rect 1021 291 1027 343
rect 1274 323 1284 343
rect 1340 323 1350 343
rect 1079 295 1092 323
rect 1144 295 1157 323
rect 1209 295 1222 323
rect 1274 295 1286 323
rect 1338 295 1350 323
rect 1402 295 1414 323
rect 1466 295 1478 323
rect 1530 295 1542 323
rect 1274 291 1284 295
rect 1340 291 1350 295
rect 1594 291 1606 343
rect 1667 323 1670 343
rect 1850 323 1854 343
rect 1658 295 1670 323
rect 1722 295 1734 323
rect 1786 295 1798 323
rect 1850 295 1862 323
rect 1667 291 1670 295
rect 1850 291 1854 295
rect 1914 291 1920 343
tri -86 275 -84 277 sw
rect 1021 275 1038 291
rect 1094 275 1120 291
rect 1176 275 1202 291
rect 1258 275 1284 291
rect 1340 275 1366 291
rect 1422 275 1448 291
rect 1504 275 1530 291
rect 1586 275 1611 291
rect 1667 275 1692 291
rect 1748 275 1773 291
rect 1829 275 1854 291
rect 1910 275 1920 291
rect -138 241 -84 275
tri -84 241 -50 275 sw
rect -138 201 50 241
rect 51 202 52 240
rect 112 202 113 240
rect 114 203 228 241
rect 114 201 176 203
tri 120 185 136 201 ne
rect -138 152 -86 160
tri -86 151 -83 154 sw
rect 136 151 176 201
rect 1021 223 1027 275
rect 1274 239 1284 275
rect 1340 239 1350 275
rect 1079 223 1092 239
rect 1144 223 1157 239
rect 1209 223 1222 239
rect 1274 223 1286 239
rect 1338 223 1350 239
rect 1402 223 1414 239
rect 1466 223 1478 239
rect 1530 223 1542 239
rect 1594 223 1606 275
rect 1667 239 1670 275
rect 1850 239 1854 275
rect 1658 223 1670 239
rect 1722 223 1734 239
rect 1786 223 1798 239
rect 1850 223 1862 239
rect 1914 223 1920 275
rect 1021 211 1920 223
rect 1021 207 1038 211
rect 1094 207 1120 211
rect 1176 207 1202 211
rect 1258 207 1284 211
rect 1340 207 1366 211
rect 1422 207 1448 211
rect 1504 207 1530 211
rect 1586 207 1611 211
rect 1667 207 1692 211
rect 1748 207 1773 211
rect 1829 207 1854 211
rect 1910 207 1920 211
rect 1021 155 1027 207
rect 1274 155 1284 207
rect 1340 155 1350 207
rect 1594 155 1606 207
rect 1667 155 1670 207
rect 1850 155 1854 207
rect 1914 155 1920 207
rect 1021 151 1920 155
rect -86 139 -83 151
tri -83 139 -71 151 sw
rect 136 139 228 151
rect -86 137 -71 139
tri -71 137 -69 139 sw
rect -86 121 -69 137
tri -69 121 -53 137 sw
tri 120 121 136 137 se
rect 136 121 176 139
rect -86 100 -1 121
rect 1 120 61 121
rect -138 88 -1 100
rect -86 81 -1 88
rect 0 82 62 120
rect 63 87 176 121
rect 1 81 61 82
rect 63 81 228 87
rect -86 63 -71 81
tri -71 63 -53 81 nw
tri -86 48 -71 63 nw
rect -138 30 -86 36
rect -138 -146 -86 -138
rect -138 -210 -86 -198
rect -138 -325 -86 -262
rect 642 -211 651 -155
rect 707 -211 770 -155
rect 826 -211 888 -155
rect 944 -211 953 -155
rect 642 -229 953 -211
rect 642 -239 673 -229
tri -86 -325 -54 -293 sw
rect 642 -295 651 -239
rect 725 -281 747 -229
rect 799 -239 821 -229
rect 873 -239 895 -229
rect 873 -281 888 -239
rect 947 -281 953 -229
rect 707 -295 770 -281
rect 826 -295 888 -281
rect 944 -295 953 -281
rect -138 -377 3486 -325
tri 3464 -388 3475 -377 ne
rect 3475 -388 3486 -377
tri 3486 -388 3549 -325 sw
tri 3475 -399 3486 -388 ne
rect 3486 -399 3549 -388
tri 3486 -410 3497 -399 ne
rect 3497 -495 3549 -399
tri 3764 -417 3793 -388 se
rect 3793 -417 3836 1371
rect 5193 1371 5645 1375
rect 5193 1319 5199 1371
rect 5259 1319 5263 1371
rect 5379 1319 5387 1371
rect 5444 1319 5457 1371
rect 5639 1319 5645 1371
rect 5193 1315 5203 1319
rect 5259 1315 5295 1319
rect 5351 1315 5387 1319
rect 5443 1315 5479 1319
rect 5535 1315 5572 1319
rect 5628 1315 5645 1319
rect 5193 1303 5645 1315
rect 5193 1251 5199 1303
rect 5251 1287 5263 1303
rect 5315 1287 5327 1303
rect 5379 1287 5392 1303
rect 5259 1251 5263 1287
rect 5379 1251 5387 1287
rect 5444 1251 5457 1303
rect 5509 1287 5522 1303
rect 5574 1287 5587 1303
rect 5639 1251 5645 1303
rect 5193 1235 5203 1251
rect 5259 1235 5295 1251
rect 5351 1235 5387 1251
rect 5443 1235 5479 1251
rect 5535 1235 5572 1251
rect 5628 1235 5645 1251
rect 5193 1183 5199 1235
rect 5259 1231 5263 1235
rect 5379 1231 5387 1235
rect 5251 1203 5263 1231
rect 5315 1203 5327 1231
rect 5379 1203 5392 1231
rect 5259 1183 5263 1203
rect 5379 1183 5387 1203
rect 5444 1183 5457 1235
rect 5509 1203 5522 1231
rect 5574 1203 5587 1231
rect 5639 1183 5645 1235
rect 5193 1167 5203 1183
rect 5259 1167 5295 1183
rect 5351 1167 5387 1183
rect 5443 1167 5479 1183
rect 5535 1167 5572 1183
rect 5628 1167 5645 1183
rect 5193 1115 5199 1167
rect 5259 1147 5263 1167
rect 5379 1147 5387 1167
rect 5251 1119 5263 1147
rect 5315 1119 5327 1147
rect 5379 1119 5392 1147
rect 5259 1115 5263 1119
rect 5379 1115 5387 1119
rect 5444 1115 5457 1167
rect 5509 1119 5522 1147
rect 5574 1119 5587 1147
rect 5639 1115 5645 1167
rect 5193 1099 5203 1115
rect 5259 1099 5295 1115
rect 5351 1099 5387 1115
rect 5443 1099 5479 1115
rect 5535 1099 5572 1115
rect 5628 1099 5645 1115
rect 5193 1047 5199 1099
rect 5259 1063 5263 1099
rect 5379 1063 5387 1099
rect 5251 1047 5263 1063
rect 5315 1047 5327 1063
rect 5379 1047 5392 1063
rect 5444 1047 5457 1099
rect 5509 1047 5522 1063
rect 5574 1047 5587 1063
rect 5639 1047 5645 1099
rect 5193 1035 5645 1047
rect 5193 1031 5203 1035
rect 5259 1031 5295 1035
rect 5351 1031 5387 1035
rect 5443 1031 5479 1035
rect 5535 1031 5572 1035
rect 5628 1031 5645 1035
rect 5193 979 5199 1031
rect 5259 979 5263 1031
rect 5379 979 5387 1031
rect 5444 979 5457 1031
rect 5639 979 5645 1031
rect 5193 975 5645 979
rect 7505 1371 8404 1375
rect 7505 1319 7511 1371
rect 7758 1319 7768 1371
rect 7824 1319 7834 1371
rect 8078 1319 8090 1371
rect 8151 1319 8154 1371
rect 8334 1319 8338 1371
rect 8398 1319 8404 1371
rect 7505 1315 7522 1319
rect 7578 1315 7604 1319
rect 7660 1315 7686 1319
rect 7742 1315 7768 1319
rect 7824 1315 7850 1319
rect 7906 1315 7932 1319
rect 7988 1315 8014 1319
rect 8070 1315 8095 1319
rect 8151 1315 8176 1319
rect 8232 1315 8257 1319
rect 8313 1315 8338 1319
rect 8394 1315 8404 1319
rect 7505 1303 8404 1315
rect 7505 1251 7511 1303
rect 7563 1287 7576 1303
rect 7628 1287 7641 1303
rect 7693 1287 7706 1303
rect 7758 1287 7770 1303
rect 7822 1287 7834 1303
rect 7886 1287 7898 1303
rect 7950 1287 7962 1303
rect 8014 1287 8026 1303
rect 7758 1251 7768 1287
rect 7824 1251 7834 1287
rect 8078 1251 8090 1303
rect 8142 1287 8154 1303
rect 8206 1287 8218 1303
rect 8270 1287 8282 1303
rect 8334 1287 8346 1303
rect 8151 1251 8154 1287
rect 8334 1251 8338 1287
rect 8398 1251 8404 1303
rect 7505 1235 7522 1251
rect 7578 1235 7604 1251
rect 7660 1235 7686 1251
rect 7742 1235 7768 1251
rect 7824 1235 7850 1251
rect 7906 1235 7932 1251
rect 7988 1235 8014 1251
rect 8070 1235 8095 1251
rect 8151 1235 8176 1251
rect 8232 1235 8257 1251
rect 8313 1235 8338 1251
rect 8394 1235 8404 1251
rect 7505 1183 7511 1235
rect 7758 1231 7768 1235
rect 7824 1231 7834 1235
rect 7563 1203 7576 1231
rect 7628 1203 7641 1231
rect 7693 1203 7706 1231
rect 7758 1203 7770 1231
rect 7822 1203 7834 1231
rect 7886 1203 7898 1231
rect 7950 1203 7962 1231
rect 8014 1203 8026 1231
rect 7758 1183 7768 1203
rect 7824 1183 7834 1203
rect 8078 1183 8090 1235
rect 8151 1231 8154 1235
rect 8334 1231 8338 1235
rect 8142 1203 8154 1231
rect 8206 1203 8218 1231
rect 8270 1203 8282 1231
rect 8334 1203 8346 1231
rect 8151 1183 8154 1203
rect 8334 1183 8338 1203
rect 8398 1183 8404 1235
rect 7505 1167 7522 1183
rect 7578 1167 7604 1183
rect 7660 1167 7686 1183
rect 7742 1167 7768 1183
rect 7824 1167 7850 1183
rect 7906 1167 7932 1183
rect 7988 1167 8014 1183
rect 8070 1167 8095 1183
rect 8151 1167 8176 1183
rect 8232 1167 8257 1183
rect 8313 1167 8338 1183
rect 8394 1167 8404 1183
rect 7505 1115 7511 1167
rect 7758 1147 7768 1167
rect 7824 1147 7834 1167
rect 7563 1119 7576 1147
rect 7628 1119 7641 1147
rect 7693 1119 7706 1147
rect 7758 1119 7770 1147
rect 7822 1119 7834 1147
rect 7886 1119 7898 1147
rect 7950 1119 7962 1147
rect 8014 1119 8026 1147
rect 7758 1115 7768 1119
rect 7824 1115 7834 1119
rect 8078 1115 8090 1167
rect 8151 1147 8154 1167
rect 8334 1147 8338 1167
rect 8142 1119 8154 1147
rect 8206 1119 8218 1147
rect 8270 1119 8282 1147
rect 8334 1119 8346 1147
rect 8151 1115 8154 1119
rect 8334 1115 8338 1119
rect 8398 1115 8404 1167
rect 7505 1099 7522 1115
rect 7578 1099 7604 1115
rect 7660 1099 7686 1115
rect 7742 1099 7768 1115
rect 7824 1099 7850 1115
rect 7906 1099 7932 1115
rect 7988 1099 8014 1115
rect 8070 1099 8095 1115
rect 8151 1099 8176 1115
rect 8232 1099 8257 1115
rect 8313 1099 8338 1115
rect 8394 1099 8404 1115
rect 7505 1047 7511 1099
rect 7758 1063 7768 1099
rect 7824 1063 7834 1099
rect 7563 1047 7576 1063
rect 7628 1047 7641 1063
rect 7693 1047 7706 1063
rect 7758 1047 7770 1063
rect 7822 1047 7834 1063
rect 7886 1047 7898 1063
rect 7950 1047 7962 1063
rect 8014 1047 8026 1063
rect 8078 1047 8090 1099
rect 8151 1063 8154 1099
rect 8334 1063 8338 1099
rect 8142 1047 8154 1063
rect 8206 1047 8218 1063
rect 8270 1047 8282 1063
rect 8334 1047 8346 1063
rect 8398 1047 8404 1099
rect 7505 1035 8404 1047
rect 7505 1031 7522 1035
rect 7578 1031 7604 1035
rect 7660 1031 7686 1035
rect 7742 1031 7768 1035
rect 7824 1031 7850 1035
rect 7906 1031 7932 1035
rect 7988 1031 8014 1035
rect 8070 1031 8095 1035
rect 8151 1031 8176 1035
rect 8232 1031 8257 1035
rect 8313 1031 8338 1035
rect 8394 1031 8404 1035
rect 7505 979 7511 1031
rect 7758 979 7768 1031
rect 7824 979 7834 1031
rect 8078 979 8090 1031
rect 8151 979 8154 1031
rect 8334 979 8338 1031
rect 8398 979 8404 1031
rect 7505 975 8404 979
rect 19610 1412 19890 1452
rect 19891 1413 19892 1451
rect 19952 1413 19953 1451
rect 19954 1417 20118 1452
tri 20118 1417 20153 1452 sw
rect 19954 1412 20153 1417
rect 19610 1402 19669 1412
tri 19669 1402 19679 1412 nw
tri 19967 1402 19977 1412 ne
rect 19977 1402 20153 1412
rect 19610 1396 19662 1402
rect 3907 861 4804 862
rect 3907 809 3913 861
rect 3965 858 3977 861
rect 4029 858 4041 861
rect 4093 858 4105 861
rect 4157 858 4169 861
rect 3972 809 3977 858
rect 4157 809 4162 858
rect 4221 809 4233 861
rect 4285 858 4297 861
rect 4349 858 4361 861
rect 4413 858 4425 861
rect 4477 809 4489 861
rect 4541 858 4553 861
rect 4605 858 4617 861
rect 4669 858 4681 861
rect 4733 858 4746 861
rect 4546 809 4553 858
rect 4733 809 4739 858
rect 4798 809 4804 861
rect 3907 802 3916 809
rect 3972 802 3998 809
rect 4054 802 4080 809
rect 4136 802 4162 809
rect 4218 802 4244 809
rect 4300 802 4326 809
rect 4382 802 4408 809
rect 4464 802 4490 809
rect 4546 802 4573 809
rect 4629 802 4656 809
rect 4712 802 4739 809
rect 4795 802 4804 809
rect 3907 789 4804 802
rect 3907 737 3913 789
rect 3965 737 3977 789
rect 4029 737 4041 789
rect 4093 737 4105 789
rect 4157 737 4169 789
rect 4221 737 4233 789
rect 4285 737 4297 789
rect 4349 737 4361 789
rect 4413 737 4425 789
rect 4477 737 4489 789
rect 4541 737 4553 789
rect 4605 737 4617 789
rect 4669 737 4681 789
rect 4733 737 4746 789
rect 4798 737 4804 789
rect 3907 724 4804 737
rect 3907 717 3916 724
rect 3972 717 3998 724
rect 4054 717 4080 724
rect 4136 717 4162 724
rect 4218 717 4244 724
rect 4300 717 4326 724
rect 4382 717 4408 724
rect 4464 717 4490 724
rect 4546 717 4573 724
rect 4629 717 4656 724
rect 4712 717 4739 724
rect 4795 717 4804 724
rect 3907 665 3913 717
rect 3972 668 3977 717
rect 4157 668 4162 717
rect 3965 665 3977 668
rect 4029 665 4041 668
rect 4093 665 4105 668
rect 4157 665 4169 668
rect 4221 665 4233 717
rect 4285 665 4297 668
rect 4349 665 4361 668
rect 4413 665 4425 668
rect 4477 665 4489 717
rect 4546 668 4553 717
rect 4733 668 4739 717
rect 4541 665 4553 668
rect 4605 665 4617 668
rect 4669 665 4681 668
rect 4733 665 4746 668
rect 4798 665 4804 717
rect 3907 664 4804 665
rect 8550 861 9447 862
rect 8550 809 8556 861
rect 8608 858 8621 861
rect 8673 858 8685 861
rect 8737 858 8749 861
rect 8801 858 8813 861
rect 8615 809 8621 858
rect 8801 809 8808 858
rect 8865 809 8877 861
rect 8929 858 8941 861
rect 8993 858 9005 861
rect 9057 858 9069 861
rect 9121 809 9133 861
rect 9185 858 9197 861
rect 9249 858 9261 861
rect 9313 858 9325 861
rect 9377 858 9389 861
rect 9192 809 9197 858
rect 9377 809 9382 858
rect 9441 809 9447 861
rect 8550 802 8559 809
rect 8615 802 8642 809
rect 8698 802 8725 809
rect 8781 802 8808 809
rect 8864 802 8890 809
rect 8946 802 8972 809
rect 9028 802 9054 809
rect 9110 802 9136 809
rect 9192 802 9218 809
rect 9274 802 9300 809
rect 9356 802 9382 809
rect 9438 802 9447 809
rect 8550 789 9447 802
rect 8550 737 8556 789
rect 8608 737 8621 789
rect 8673 737 8685 789
rect 8737 737 8749 789
rect 8801 737 8813 789
rect 8865 737 8877 789
rect 8929 737 8941 789
rect 8993 737 9005 789
rect 9057 737 9069 789
rect 9121 737 9133 789
rect 9185 737 9197 789
rect 9249 737 9261 789
rect 9313 737 9325 789
rect 9377 737 9389 789
rect 9441 737 9447 789
rect 8550 724 9447 737
rect 8550 717 8559 724
rect 8615 717 8642 724
rect 8698 717 8725 724
rect 8781 717 8808 724
rect 8864 717 8890 724
rect 8946 717 8972 724
rect 9028 717 9054 724
rect 9110 717 9136 724
rect 9192 717 9218 724
rect 9274 717 9300 724
rect 9356 717 9382 724
rect 9438 717 9447 724
rect 8550 665 8556 717
rect 8615 668 8621 717
rect 8801 668 8808 717
rect 8608 665 8621 668
rect 8673 665 8685 668
rect 8737 665 8749 668
rect 8801 665 8813 668
rect 8865 665 8877 717
rect 8929 665 8941 668
rect 8993 665 9005 668
rect 9057 665 9069 668
rect 9121 665 9133 717
rect 9192 668 9197 717
rect 9377 668 9382 717
rect 9185 665 9197 668
rect 9249 665 9261 668
rect 9313 665 9325 668
rect 9377 665 9389 668
rect 9441 665 9447 717
rect 8550 664 9447 665
rect 5193 547 5645 551
rect 5193 495 5199 547
rect 5259 495 5263 547
rect 5379 495 5387 547
rect 5444 495 5457 547
rect 5639 495 5645 547
rect 5193 491 5203 495
rect 5259 491 5295 495
rect 5351 491 5387 495
rect 5443 491 5479 495
rect 5535 491 5572 495
rect 5628 491 5645 495
rect 5193 479 5645 491
rect 5193 427 5199 479
rect 5251 463 5263 479
rect 5315 463 5327 479
rect 5379 463 5392 479
rect 5259 427 5263 463
rect 5379 427 5387 463
rect 5444 427 5457 479
rect 5509 463 5522 479
rect 5574 463 5587 479
rect 5639 427 5645 479
rect 5193 411 5203 427
rect 5259 411 5295 427
rect 5351 411 5387 427
rect 5443 411 5479 427
rect 5535 411 5572 427
rect 5628 411 5645 427
rect 5193 359 5199 411
rect 5259 407 5263 411
rect 5379 407 5387 411
rect 5251 379 5263 407
rect 5315 379 5327 407
rect 5379 379 5392 407
rect 5259 359 5263 379
rect 5379 359 5387 379
rect 5444 359 5457 411
rect 5509 379 5522 407
rect 5574 379 5587 407
rect 5639 359 5645 411
rect 5193 343 5203 359
rect 5259 343 5295 359
rect 5351 343 5387 359
rect 5443 343 5479 359
rect 5535 343 5572 359
rect 5628 343 5645 359
rect 5193 291 5199 343
rect 5259 323 5263 343
rect 5379 323 5387 343
rect 5251 295 5263 323
rect 5315 295 5327 323
rect 5379 295 5392 323
rect 5259 291 5263 295
rect 5379 291 5387 295
rect 5444 291 5457 343
rect 5509 295 5522 323
rect 5574 295 5587 323
rect 5639 291 5645 343
rect 5193 275 5203 291
rect 5259 275 5295 291
rect 5351 275 5387 291
rect 5443 275 5479 291
rect 5535 275 5572 291
rect 5628 275 5645 291
rect 5193 223 5199 275
rect 5259 239 5263 275
rect 5379 239 5387 275
rect 5251 223 5263 239
rect 5315 223 5327 239
rect 5379 223 5392 239
rect 5444 223 5457 275
rect 5509 223 5522 239
rect 5574 223 5587 239
rect 5639 223 5645 275
rect 5193 211 5645 223
rect 5193 207 5203 211
rect 5259 207 5295 211
rect 5351 207 5387 211
rect 5443 207 5479 211
rect 5535 207 5572 211
rect 5628 207 5645 211
rect 5193 155 5199 207
rect 5259 155 5263 207
rect 5379 155 5387 207
rect 5444 155 5457 207
rect 5639 155 5645 207
rect 5193 151 5645 155
rect 7505 547 8404 551
rect 7505 495 7511 547
rect 7758 495 7768 547
rect 7824 495 7834 547
rect 8078 495 8090 547
rect 8151 495 8154 547
rect 8334 495 8338 547
rect 8398 495 8404 547
rect 7505 491 7522 495
rect 7578 491 7604 495
rect 7660 491 7686 495
rect 7742 491 7768 495
rect 7824 491 7850 495
rect 7906 491 7932 495
rect 7988 491 8014 495
rect 8070 491 8095 495
rect 8151 491 8176 495
rect 8232 491 8257 495
rect 8313 491 8338 495
rect 8394 491 8404 495
rect 7505 479 8404 491
rect 7505 427 7511 479
rect 7563 463 7576 479
rect 7628 463 7641 479
rect 7693 463 7706 479
rect 7758 463 7770 479
rect 7822 463 7834 479
rect 7886 463 7898 479
rect 7950 463 7962 479
rect 8014 463 8026 479
rect 7758 427 7768 463
rect 7824 427 7834 463
rect 8078 427 8090 479
rect 8142 463 8154 479
rect 8206 463 8218 479
rect 8270 463 8282 479
rect 8334 463 8346 479
rect 8151 427 8154 463
rect 8334 427 8338 463
rect 8398 427 8404 479
rect 7505 411 7522 427
rect 7578 411 7604 427
rect 7660 411 7686 427
rect 7742 411 7768 427
rect 7824 411 7850 427
rect 7906 411 7932 427
rect 7988 411 8014 427
rect 8070 411 8095 427
rect 8151 411 8176 427
rect 8232 411 8257 427
rect 8313 411 8338 427
rect 8394 411 8404 427
rect 7505 359 7511 411
rect 7758 407 7768 411
rect 7824 407 7834 411
rect 7563 379 7576 407
rect 7628 379 7641 407
rect 7693 379 7706 407
rect 7758 379 7770 407
rect 7822 379 7834 407
rect 7886 379 7898 407
rect 7950 379 7962 407
rect 8014 379 8026 407
rect 7758 359 7768 379
rect 7824 359 7834 379
rect 8078 359 8090 411
rect 8151 407 8154 411
rect 8334 407 8338 411
rect 8142 379 8154 407
rect 8206 379 8218 407
rect 8270 379 8282 407
rect 8334 379 8346 407
rect 8151 359 8154 379
rect 8334 359 8338 379
rect 8398 359 8404 411
rect 7505 343 7522 359
rect 7578 343 7604 359
rect 7660 343 7686 359
rect 7742 343 7768 359
rect 7824 343 7850 359
rect 7906 343 7932 359
rect 7988 343 8014 359
rect 8070 343 8095 359
rect 8151 343 8176 359
rect 8232 343 8257 359
rect 8313 343 8338 359
rect 8394 343 8404 359
rect 7505 291 7511 343
rect 7758 323 7768 343
rect 7824 323 7834 343
rect 7563 295 7576 323
rect 7628 295 7641 323
rect 7693 295 7706 323
rect 7758 295 7770 323
rect 7822 295 7834 323
rect 7886 295 7898 323
rect 7950 295 7962 323
rect 8014 295 8026 323
rect 7758 291 7768 295
rect 7824 291 7834 295
rect 8078 291 8090 343
rect 8151 323 8154 343
rect 8334 323 8338 343
rect 8142 295 8154 323
rect 8206 295 8218 323
rect 8270 295 8282 323
rect 8334 295 8346 323
rect 8151 291 8154 295
rect 8334 291 8338 295
rect 8398 291 8404 343
rect 7505 275 7522 291
rect 7578 275 7604 291
rect 7660 275 7686 291
rect 7742 275 7768 291
rect 7824 275 7850 291
rect 7906 275 7932 291
rect 7988 275 8014 291
rect 8070 275 8095 291
rect 8151 275 8176 291
rect 8232 275 8257 291
rect 8313 275 8338 291
rect 8394 275 8404 291
rect 7505 223 7511 275
rect 7758 239 7768 275
rect 7824 239 7834 275
rect 7563 223 7576 239
rect 7628 223 7641 239
rect 7693 223 7706 239
rect 7758 223 7770 239
rect 7822 223 7834 239
rect 7886 223 7898 239
rect 7950 223 7962 239
rect 8014 223 8026 239
rect 8078 223 8090 275
rect 8151 239 8154 275
rect 8334 239 8338 275
rect 8142 223 8154 239
rect 8206 223 8218 239
rect 8270 223 8282 239
rect 8334 223 8346 239
rect 8398 223 8404 275
rect 7505 211 8404 223
rect 7505 207 7522 211
rect 7578 207 7604 211
rect 7660 207 7686 211
rect 7742 207 7768 211
rect 7824 207 7850 211
rect 7906 207 7932 211
rect 7988 207 8014 211
rect 8070 207 8095 211
rect 8151 207 8176 211
rect 8232 207 8257 211
rect 8313 207 8338 211
rect 8394 207 8404 211
rect 7505 155 7511 207
rect 7758 155 7768 207
rect 7824 155 7834 207
rect 8078 155 8090 207
rect 8151 155 8154 207
rect 8334 155 8338 207
rect 8398 155 8404 207
rect 7505 151 8404 155
rect 3907 38 3916 39
rect 3972 38 3998 39
rect 4054 38 4080 39
rect 4136 38 4162 39
rect 4218 38 4244 39
rect 4300 38 4326 39
rect 4382 38 4408 39
rect 4464 38 4490 39
rect 4546 38 4573 39
rect 4629 38 4656 39
rect 4712 38 4739 39
rect 4795 38 4804 39
rect 3907 -14 3913 38
rect 3972 -14 3978 38
rect 4158 -14 4162 38
rect 4222 -14 4234 38
rect 4478 -14 4490 38
rect 4546 -14 4554 38
rect 4734 -14 4739 38
rect 4798 -14 4804 38
rect 3907 -17 3916 -14
rect 3972 -17 3998 -14
rect 4054 -17 4080 -14
rect 4136 -17 4162 -14
rect 4218 -17 4244 -14
rect 4300 -17 4326 -14
rect 4382 -17 4408 -14
rect 4464 -17 4490 -14
rect 4546 -17 4573 -14
rect 4629 -17 4656 -14
rect 4712 -17 4739 -14
rect 4795 -17 4804 -14
rect 3907 -34 4804 -17
rect 3907 -86 3913 -34
rect 3965 -86 3978 -34
rect 4030 -86 4042 -34
rect 4094 -86 4106 -34
rect 4158 -86 4170 -34
rect 4222 -86 4234 -34
rect 4286 -86 4298 -34
rect 4350 -86 4362 -34
rect 4414 -86 4426 -34
rect 4478 -86 4490 -34
rect 4542 -86 4554 -34
rect 4606 -86 4618 -34
rect 4670 -86 4682 -34
rect 4734 -86 4746 -34
rect 4798 -86 4804 -34
rect 3907 -95 4804 -86
rect 3907 -106 3916 -95
rect 3972 -106 3998 -95
rect 4054 -106 4080 -95
rect 4136 -106 4162 -95
rect 4218 -106 4244 -95
rect 4300 -106 4326 -95
rect 4382 -106 4408 -95
rect 4464 -106 4490 -95
rect 4546 -106 4573 -95
rect 4629 -106 4656 -95
rect 4712 -106 4739 -95
rect 4795 -106 4804 -95
rect 3907 -158 3913 -106
rect 3972 -151 3978 -106
rect 4158 -151 4162 -106
rect 3965 -158 3978 -151
rect 4030 -158 4042 -151
rect 4094 -158 4106 -151
rect 4158 -158 4170 -151
rect 4222 -158 4234 -106
rect 4286 -158 4298 -151
rect 4350 -158 4362 -151
rect 4414 -158 4426 -151
rect 4478 -158 4490 -106
rect 4546 -151 4554 -106
rect 4734 -151 4739 -106
rect 4542 -158 4554 -151
rect 4606 -158 4618 -151
rect 4670 -158 4682 -151
rect 4734 -158 4746 -151
rect 4798 -158 4804 -106
rect 8550 38 9447 39
rect 8550 -14 8556 38
rect 8608 35 8621 38
rect 8673 35 8685 38
rect 8737 35 8749 38
rect 8801 35 8813 38
rect 8615 -14 8621 35
rect 8801 -14 8808 35
rect 8865 -14 8877 38
rect 8929 35 8941 38
rect 8993 35 9005 38
rect 9057 35 9069 38
rect 9121 -14 9133 38
rect 9185 35 9197 38
rect 9249 35 9261 38
rect 9313 35 9325 38
rect 9377 35 9389 38
rect 9192 -14 9197 35
rect 9377 -14 9382 35
rect 9441 -14 9447 38
rect 8550 -21 8559 -14
rect 8615 -21 8642 -14
rect 8698 -21 8725 -14
rect 8781 -21 8808 -14
rect 8864 -21 8890 -14
rect 8946 -21 8972 -14
rect 9028 -21 9054 -14
rect 9110 -21 9136 -14
rect 9192 -21 9218 -14
rect 9274 -21 9300 -14
rect 9356 -21 9382 -14
rect 9438 -21 9447 -14
rect 8550 -34 9447 -21
rect 8550 -86 8556 -34
rect 8608 -86 8621 -34
rect 8673 -86 8685 -34
rect 8737 -86 8749 -34
rect 8801 -86 8813 -34
rect 8865 -86 8877 -34
rect 8929 -86 8941 -34
rect 8993 -86 9005 -34
rect 9057 -86 9069 -34
rect 9121 -86 9133 -34
rect 9185 -86 9197 -34
rect 9249 -86 9261 -34
rect 9313 -86 9325 -34
rect 9377 -86 9389 -34
rect 9441 -86 9447 -34
rect 8550 -99 9447 -86
rect 8550 -106 8559 -99
rect 8615 -106 8642 -99
rect 8698 -106 8725 -99
rect 8781 -106 8808 -99
rect 8864 -106 8890 -99
rect 8946 -106 8972 -99
rect 9028 -106 9054 -99
rect 9110 -106 9136 -99
rect 9192 -106 9218 -99
rect 9274 -106 9300 -99
rect 9356 -106 9382 -99
rect 9438 -106 9447 -99
rect 3907 -159 4804 -158
rect 6012 -211 6021 -155
rect 6077 -211 6103 -155
rect 6159 -211 6184 -155
rect 6240 -211 6265 -155
rect 6321 -211 6346 -155
rect 6402 -211 6411 -155
rect 6012 -229 6411 -211
rect 6012 -281 6018 -229
rect 6070 -239 6085 -229
rect 6137 -239 6152 -229
rect 6204 -239 6219 -229
rect 6271 -239 6286 -229
rect 6338 -239 6353 -229
rect 6077 -281 6085 -239
rect 6338 -281 6346 -239
rect 6405 -281 6411 -229
rect 6012 -295 6021 -281
rect 6077 -295 6103 -281
rect 6159 -295 6184 -281
rect 6240 -295 6265 -281
rect 6321 -295 6346 -281
rect 6402 -295 6411 -281
rect 6943 -211 6952 -155
rect 7008 -211 7034 -155
rect 7090 -211 7115 -155
rect 7171 -211 7196 -155
rect 7252 -211 7277 -155
rect 7333 -211 7342 -155
rect 8550 -158 8556 -106
rect 8615 -155 8621 -106
rect 8801 -155 8808 -106
rect 8608 -158 8621 -155
rect 8673 -158 8685 -155
rect 8737 -158 8749 -155
rect 8801 -158 8813 -155
rect 8865 -158 8877 -106
rect 8929 -158 8941 -155
rect 8993 -158 9005 -155
rect 9057 -158 9069 -155
rect 9121 -158 9133 -106
rect 9192 -155 9197 -106
rect 9377 -155 9382 -106
rect 9185 -158 9197 -155
rect 9249 -158 9261 -155
rect 9313 -158 9325 -155
rect 9377 -158 9389 -155
rect 9441 -158 9447 -106
rect 8550 -159 9447 -158
rect 9897 -10 9949 1374
rect 11434 1371 12333 1375
rect 11434 1319 11440 1371
rect 11500 1319 11504 1371
rect 11684 1319 11687 1371
rect 11748 1319 11760 1371
rect 12004 1319 12014 1371
rect 12070 1319 12080 1371
rect 12327 1319 12333 1371
rect 11434 1315 11444 1319
rect 11500 1315 11525 1319
rect 11581 1315 11606 1319
rect 11662 1315 11687 1319
rect 11743 1315 11768 1319
rect 11824 1315 11850 1319
rect 11906 1315 11932 1319
rect 11988 1315 12014 1319
rect 12070 1315 12096 1319
rect 12152 1315 12178 1319
rect 12234 1315 12260 1319
rect 12316 1315 12333 1319
rect 11434 1303 12333 1315
rect 11434 1251 11440 1303
rect 11492 1287 11504 1303
rect 11556 1287 11568 1303
rect 11620 1287 11632 1303
rect 11684 1287 11696 1303
rect 11500 1251 11504 1287
rect 11684 1251 11687 1287
rect 11748 1251 11760 1303
rect 11812 1287 11824 1303
rect 11876 1287 11888 1303
rect 11940 1287 11952 1303
rect 12004 1287 12016 1303
rect 12068 1287 12080 1303
rect 12132 1287 12145 1303
rect 12197 1287 12210 1303
rect 12262 1287 12275 1303
rect 12004 1251 12014 1287
rect 12070 1251 12080 1287
rect 12327 1251 12333 1303
rect 11434 1235 11444 1251
rect 11500 1235 11525 1251
rect 11581 1235 11606 1251
rect 11662 1235 11687 1251
rect 11743 1235 11768 1251
rect 11824 1235 11850 1251
rect 11906 1235 11932 1251
rect 11988 1235 12014 1251
rect 12070 1235 12096 1251
rect 12152 1235 12178 1251
rect 12234 1235 12260 1251
rect 12316 1235 12333 1251
rect 11434 1183 11440 1235
rect 11500 1231 11504 1235
rect 11684 1231 11687 1235
rect 11492 1203 11504 1231
rect 11556 1203 11568 1231
rect 11620 1203 11632 1231
rect 11684 1203 11696 1231
rect 11500 1183 11504 1203
rect 11684 1183 11687 1203
rect 11748 1183 11760 1235
rect 12004 1231 12014 1235
rect 12070 1231 12080 1235
rect 11812 1203 11824 1231
rect 11876 1203 11888 1231
rect 11940 1203 11952 1231
rect 12004 1203 12016 1231
rect 12068 1203 12080 1231
rect 12132 1203 12145 1231
rect 12197 1203 12210 1231
rect 12262 1203 12275 1231
rect 12004 1183 12014 1203
rect 12070 1183 12080 1203
rect 12327 1183 12333 1235
rect 11434 1167 11444 1183
rect 11500 1167 11525 1183
rect 11581 1167 11606 1183
rect 11662 1167 11687 1183
rect 11743 1167 11768 1183
rect 11824 1167 11850 1183
rect 11906 1167 11932 1183
rect 11988 1167 12014 1183
rect 12070 1167 12096 1183
rect 12152 1167 12178 1183
rect 12234 1167 12260 1183
rect 12316 1167 12333 1183
rect 11434 1115 11440 1167
rect 11500 1147 11504 1167
rect 11684 1147 11687 1167
rect 11492 1119 11504 1147
rect 11556 1119 11568 1147
rect 11620 1119 11632 1147
rect 11684 1119 11696 1147
rect 11500 1115 11504 1119
rect 11684 1115 11687 1119
rect 11748 1115 11760 1167
rect 12004 1147 12014 1167
rect 12070 1147 12080 1167
rect 11812 1119 11824 1147
rect 11876 1119 11888 1147
rect 11940 1119 11952 1147
rect 12004 1119 12016 1147
rect 12068 1119 12080 1147
rect 12132 1119 12145 1147
rect 12197 1119 12210 1147
rect 12262 1119 12275 1147
rect 12004 1115 12014 1119
rect 12070 1115 12080 1119
rect 12327 1115 12333 1167
rect 11434 1099 11444 1115
rect 11500 1099 11525 1115
rect 11581 1099 11606 1115
rect 11662 1099 11687 1115
rect 11743 1099 11768 1115
rect 11824 1099 11850 1115
rect 11906 1099 11932 1115
rect 11988 1099 12014 1115
rect 12070 1099 12096 1115
rect 12152 1099 12178 1115
rect 12234 1099 12260 1115
rect 12316 1099 12333 1115
rect 11434 1047 11440 1099
rect 11500 1063 11504 1099
rect 11684 1063 11687 1099
rect 11492 1047 11504 1063
rect 11556 1047 11568 1063
rect 11620 1047 11632 1063
rect 11684 1047 11696 1063
rect 11748 1047 11760 1099
rect 12004 1063 12014 1099
rect 12070 1063 12080 1099
rect 11812 1047 11824 1063
rect 11876 1047 11888 1063
rect 11940 1047 11952 1063
rect 12004 1047 12016 1063
rect 12068 1047 12080 1063
rect 12132 1047 12145 1063
rect 12197 1047 12210 1063
rect 12262 1047 12275 1063
rect 12327 1047 12333 1099
rect 11434 1035 12333 1047
rect 11434 1031 11444 1035
rect 11500 1031 11525 1035
rect 11581 1031 11606 1035
rect 11662 1031 11687 1035
rect 11743 1031 11768 1035
rect 11824 1031 11850 1035
rect 11906 1031 11932 1035
rect 11988 1031 12014 1035
rect 12070 1031 12096 1035
rect 12152 1031 12178 1035
rect 12234 1031 12260 1035
rect 12316 1031 12333 1035
rect 11434 979 11440 1031
rect 11500 979 11504 1031
rect 11684 979 11687 1031
rect 11748 979 11760 1031
rect 12004 979 12014 1031
rect 12070 979 12080 1031
rect 12327 979 12333 1031
rect 11434 975 12333 979
rect 13989 1371 14888 1375
rect 13989 1319 13995 1371
rect 14242 1319 14252 1371
rect 14308 1319 14318 1371
rect 14562 1319 14574 1371
rect 14635 1319 14638 1371
rect 14818 1319 14822 1371
rect 14882 1319 14888 1371
rect 13989 1315 14006 1319
rect 14062 1315 14088 1319
rect 14144 1315 14170 1319
rect 14226 1315 14252 1319
rect 14308 1315 14334 1319
rect 14390 1315 14416 1319
rect 14472 1315 14498 1319
rect 14554 1315 14579 1319
rect 14635 1315 14660 1319
rect 14716 1315 14741 1319
rect 14797 1315 14822 1319
rect 14878 1315 14888 1319
rect 13989 1303 14888 1315
rect 13989 1251 13995 1303
rect 14047 1287 14060 1303
rect 14112 1287 14125 1303
rect 14177 1287 14190 1303
rect 14242 1287 14254 1303
rect 14306 1287 14318 1303
rect 14370 1287 14382 1303
rect 14434 1287 14446 1303
rect 14498 1287 14510 1303
rect 14242 1251 14252 1287
rect 14308 1251 14318 1287
rect 14562 1251 14574 1303
rect 14626 1287 14638 1303
rect 14690 1287 14702 1303
rect 14754 1287 14766 1303
rect 14818 1287 14830 1303
rect 14635 1251 14638 1287
rect 14818 1251 14822 1287
rect 14882 1251 14888 1303
rect 13989 1235 14006 1251
rect 14062 1235 14088 1251
rect 14144 1235 14170 1251
rect 14226 1235 14252 1251
rect 14308 1235 14334 1251
rect 14390 1235 14416 1251
rect 14472 1235 14498 1251
rect 14554 1235 14579 1251
rect 14635 1235 14660 1251
rect 14716 1235 14741 1251
rect 14797 1235 14822 1251
rect 14878 1235 14888 1251
rect 13989 1183 13995 1235
rect 14242 1231 14252 1235
rect 14308 1231 14318 1235
rect 14047 1203 14060 1231
rect 14112 1203 14125 1231
rect 14177 1203 14190 1231
rect 14242 1203 14254 1231
rect 14306 1203 14318 1231
rect 14370 1203 14382 1231
rect 14434 1203 14446 1231
rect 14498 1203 14510 1231
rect 14242 1183 14252 1203
rect 14308 1183 14318 1203
rect 14562 1183 14574 1235
rect 14635 1231 14638 1235
rect 14818 1231 14822 1235
rect 14626 1203 14638 1231
rect 14690 1203 14702 1231
rect 14754 1203 14766 1231
rect 14818 1203 14830 1231
rect 14635 1183 14638 1203
rect 14818 1183 14822 1203
rect 14882 1183 14888 1235
rect 13989 1167 14006 1183
rect 14062 1167 14088 1183
rect 14144 1167 14170 1183
rect 14226 1167 14252 1183
rect 14308 1167 14334 1183
rect 14390 1167 14416 1183
rect 14472 1167 14498 1183
rect 14554 1167 14579 1183
rect 14635 1167 14660 1183
rect 14716 1167 14741 1183
rect 14797 1167 14822 1183
rect 14878 1167 14888 1183
rect 13989 1115 13995 1167
rect 14242 1147 14252 1167
rect 14308 1147 14318 1167
rect 14047 1119 14060 1147
rect 14112 1119 14125 1147
rect 14177 1119 14190 1147
rect 14242 1119 14254 1147
rect 14306 1119 14318 1147
rect 14370 1119 14382 1147
rect 14434 1119 14446 1147
rect 14498 1119 14510 1147
rect 14242 1115 14252 1119
rect 14308 1115 14318 1119
rect 14562 1115 14574 1167
rect 14635 1147 14638 1167
rect 14818 1147 14822 1167
rect 14626 1119 14638 1147
rect 14690 1119 14702 1147
rect 14754 1119 14766 1147
rect 14818 1119 14830 1147
rect 14635 1115 14638 1119
rect 14818 1115 14822 1119
rect 14882 1115 14888 1167
rect 13989 1099 14006 1115
rect 14062 1099 14088 1115
rect 14144 1099 14170 1115
rect 14226 1099 14252 1115
rect 14308 1099 14334 1115
rect 14390 1099 14416 1115
rect 14472 1099 14498 1115
rect 14554 1099 14579 1115
rect 14635 1099 14660 1115
rect 14716 1099 14741 1115
rect 14797 1099 14822 1115
rect 14878 1099 14888 1115
rect 13989 1047 13995 1099
rect 14242 1063 14252 1099
rect 14308 1063 14318 1099
rect 14047 1047 14060 1063
rect 14112 1047 14125 1063
rect 14177 1047 14190 1063
rect 14242 1047 14254 1063
rect 14306 1047 14318 1063
rect 14370 1047 14382 1063
rect 14434 1047 14446 1063
rect 14498 1047 14510 1063
rect 14562 1047 14574 1099
rect 14635 1063 14638 1099
rect 14818 1063 14822 1099
rect 14626 1047 14638 1063
rect 14690 1047 14702 1063
rect 14754 1047 14766 1063
rect 14818 1047 14830 1063
rect 14882 1047 14888 1099
rect 13989 1035 14888 1047
rect 13989 1031 14006 1035
rect 14062 1031 14088 1035
rect 14144 1031 14170 1035
rect 14226 1031 14252 1035
rect 14308 1031 14334 1035
rect 14390 1031 14416 1035
rect 14472 1031 14498 1035
rect 14554 1031 14579 1035
rect 14635 1031 14660 1035
rect 14716 1031 14741 1035
rect 14797 1031 14822 1035
rect 14878 1031 14888 1035
rect 13989 979 13995 1031
rect 14242 979 14252 1031
rect 14308 979 14318 1031
rect 14562 979 14574 1031
rect 14635 979 14638 1031
rect 14818 979 14822 1031
rect 14882 979 14888 1031
rect 13989 975 14888 979
rect 17918 1371 18817 1375
rect 17918 1319 17924 1371
rect 17984 1319 17988 1371
rect 18168 1319 18171 1371
rect 18232 1319 18244 1371
rect 18488 1319 18498 1371
rect 18554 1319 18564 1371
rect 18811 1319 18817 1371
rect 17918 1315 17928 1319
rect 17984 1315 18009 1319
rect 18065 1315 18090 1319
rect 18146 1315 18171 1319
rect 18227 1315 18252 1319
rect 18308 1315 18334 1319
rect 18390 1315 18416 1319
rect 18472 1315 18498 1319
rect 18554 1315 18580 1319
rect 18636 1315 18662 1319
rect 18718 1315 18744 1319
rect 18800 1315 18817 1319
rect 17918 1303 18817 1315
rect 17918 1251 17924 1303
rect 17976 1287 17988 1303
rect 18040 1287 18052 1303
rect 18104 1287 18116 1303
rect 18168 1287 18180 1303
rect 17984 1251 17988 1287
rect 18168 1251 18171 1287
rect 18232 1251 18244 1303
rect 18296 1287 18308 1303
rect 18360 1287 18372 1303
rect 18424 1287 18436 1303
rect 18488 1287 18500 1303
rect 18552 1287 18564 1303
rect 18616 1287 18629 1303
rect 18681 1287 18694 1303
rect 18746 1287 18759 1303
rect 18488 1251 18498 1287
rect 18554 1251 18564 1287
rect 18811 1251 18817 1303
rect 17918 1235 17928 1251
rect 17984 1235 18009 1251
rect 18065 1235 18090 1251
rect 18146 1235 18171 1251
rect 18227 1235 18252 1251
rect 18308 1235 18334 1251
rect 18390 1235 18416 1251
rect 18472 1235 18498 1251
rect 18554 1235 18580 1251
rect 18636 1235 18662 1251
rect 18718 1235 18744 1251
rect 18800 1235 18817 1251
rect 17918 1183 17924 1235
rect 17984 1231 17988 1235
rect 18168 1231 18171 1235
rect 17976 1203 17988 1231
rect 18040 1203 18052 1231
rect 18104 1203 18116 1231
rect 18168 1203 18180 1231
rect 17984 1183 17988 1203
rect 18168 1183 18171 1203
rect 18232 1183 18244 1235
rect 18488 1231 18498 1235
rect 18554 1231 18564 1235
rect 18296 1203 18308 1231
rect 18360 1203 18372 1231
rect 18424 1203 18436 1231
rect 18488 1203 18500 1231
rect 18552 1203 18564 1231
rect 18616 1203 18629 1231
rect 18681 1203 18694 1231
rect 18746 1203 18759 1231
rect 18488 1183 18498 1203
rect 18554 1183 18564 1203
rect 18811 1183 18817 1235
rect 17918 1167 17928 1183
rect 17984 1167 18009 1183
rect 18065 1167 18090 1183
rect 18146 1167 18171 1183
rect 18227 1167 18252 1183
rect 18308 1167 18334 1183
rect 18390 1167 18416 1183
rect 18472 1167 18498 1183
rect 18554 1167 18580 1183
rect 18636 1167 18662 1183
rect 18718 1167 18744 1183
rect 18800 1167 18817 1183
rect 17918 1115 17924 1167
rect 17984 1147 17988 1167
rect 18168 1147 18171 1167
rect 17976 1119 17988 1147
rect 18040 1119 18052 1147
rect 18104 1119 18116 1147
rect 18168 1119 18180 1147
rect 17984 1115 17988 1119
rect 18168 1115 18171 1119
rect 18232 1115 18244 1167
rect 18488 1147 18498 1167
rect 18554 1147 18564 1167
rect 18296 1119 18308 1147
rect 18360 1119 18372 1147
rect 18424 1119 18436 1147
rect 18488 1119 18500 1147
rect 18552 1119 18564 1147
rect 18616 1119 18629 1147
rect 18681 1119 18694 1147
rect 18746 1119 18759 1147
rect 18488 1115 18498 1119
rect 18554 1115 18564 1119
rect 18811 1115 18817 1167
tri 19662 1395 19669 1402 nw
tri 19977 1395 19984 1402 ne
rect 19984 1395 20153 1402
tri 19984 1379 20000 1395 ne
rect 20000 1379 20153 1395
tri 20072 1352 20099 1379 ne
rect 19610 1332 19662 1344
rect 19610 1258 19662 1280
rect 19611 1256 19661 1257
rect 19610 1196 19662 1256
rect 19611 1195 19661 1196
rect 19610 1190 19662 1194
rect 19759 1203 19811 1211
rect 19610 1151 19759 1190
rect 19610 1139 19811 1151
rect 19610 1132 19759 1139
rect 17918 1099 17928 1115
rect 17984 1099 18009 1115
rect 18065 1099 18090 1115
rect 18146 1099 18171 1115
rect 18227 1099 18252 1115
rect 18308 1099 18334 1115
rect 18390 1099 18416 1115
rect 18472 1099 18498 1115
rect 18554 1099 18580 1115
rect 18636 1099 18662 1115
rect 18718 1099 18744 1115
rect 18800 1099 18817 1115
rect 17918 1047 17924 1099
rect 17984 1063 17988 1099
rect 18168 1063 18171 1099
rect 17976 1047 17988 1063
rect 18040 1047 18052 1063
rect 18104 1047 18116 1063
rect 18168 1047 18180 1063
rect 18232 1047 18244 1099
rect 18488 1063 18498 1099
rect 18554 1063 18564 1099
rect 18296 1047 18308 1063
rect 18360 1047 18372 1063
rect 18424 1047 18436 1063
rect 18488 1047 18500 1063
rect 18552 1047 18564 1063
rect 18616 1047 18629 1063
rect 18681 1047 18694 1063
rect 18746 1047 18759 1063
rect 18811 1047 18817 1099
rect 19759 1081 19811 1087
rect 17918 1035 18817 1047
rect 20099 1035 20153 1379
tri 20153 1035 20176 1058 sw
rect 17918 1031 17928 1035
rect 17984 1031 18009 1035
rect 18065 1031 18090 1035
rect 18146 1031 18171 1035
rect 18227 1031 18252 1035
rect 18308 1031 18334 1035
rect 18390 1031 18416 1035
rect 18472 1031 18498 1035
rect 18554 1031 18580 1035
rect 18636 1031 18662 1035
rect 18718 1031 18744 1035
rect 18800 1031 18817 1035
rect 17918 979 17924 1031
rect 17984 979 17988 1031
rect 18168 979 18171 1031
rect 18232 979 18244 1031
rect 18488 979 18498 1031
rect 18554 979 18564 1031
rect 18811 979 18817 1031
rect 17918 975 18817 979
rect 19610 1027 20058 1035
rect 19662 975 20006 1027
rect 19610 963 20058 975
rect 19662 911 20006 963
rect 19610 905 20058 911
rect 20099 1027 20250 1035
rect 20099 975 20198 1027
rect 20099 963 20250 975
rect 20099 911 20198 963
rect 20099 905 20250 911
rect 10391 861 11288 862
rect 10391 809 10397 861
rect 10449 858 10461 861
rect 10513 858 10525 861
rect 10577 858 10589 861
rect 10641 858 10653 861
rect 10456 809 10461 858
rect 10641 809 10646 858
rect 10705 809 10717 861
rect 10769 858 10781 861
rect 10833 858 10845 861
rect 10897 858 10909 861
rect 10961 809 10973 861
rect 11025 858 11037 861
rect 11089 858 11101 861
rect 11153 858 11165 861
rect 11217 858 11230 861
rect 11030 809 11037 858
rect 11217 809 11223 858
rect 11282 809 11288 861
rect 10391 802 10400 809
rect 10456 802 10482 809
rect 10538 802 10564 809
rect 10620 802 10646 809
rect 10702 802 10728 809
rect 10784 802 10810 809
rect 10866 802 10892 809
rect 10948 802 10974 809
rect 11030 802 11057 809
rect 11113 802 11140 809
rect 11196 802 11223 809
rect 11279 802 11288 809
rect 10391 789 11288 802
rect 10391 737 10397 789
rect 10449 737 10461 789
rect 10513 737 10525 789
rect 10577 737 10589 789
rect 10641 737 10653 789
rect 10705 737 10717 789
rect 10769 737 10781 789
rect 10833 737 10845 789
rect 10897 737 10909 789
rect 10961 737 10973 789
rect 11025 737 11037 789
rect 11089 737 11101 789
rect 11153 737 11165 789
rect 11217 737 11230 789
rect 11282 737 11288 789
rect 10391 724 11288 737
rect 10391 717 10400 724
rect 10456 717 10482 724
rect 10538 717 10564 724
rect 10620 717 10646 724
rect 10702 717 10728 724
rect 10784 717 10810 724
rect 10866 717 10892 724
rect 10948 717 10974 724
rect 11030 717 11057 724
rect 11113 717 11140 724
rect 11196 717 11223 724
rect 11279 717 11288 724
rect 10391 665 10397 717
rect 10456 668 10461 717
rect 10641 668 10646 717
rect 10449 665 10461 668
rect 10513 665 10525 668
rect 10577 665 10589 668
rect 10641 665 10653 668
rect 10705 665 10717 717
rect 10769 665 10781 668
rect 10833 665 10845 668
rect 10897 665 10909 668
rect 10961 665 10973 717
rect 11030 668 11037 717
rect 11217 668 11223 717
rect 11025 665 11037 668
rect 11089 665 11101 668
rect 11153 665 11165 668
rect 11217 665 11230 668
rect 11282 665 11288 717
rect 10391 664 11288 665
rect 15034 861 15931 862
rect 15034 809 15040 861
rect 15092 858 15105 861
rect 15157 858 15169 861
rect 15221 858 15233 861
rect 15285 858 15297 861
rect 15099 809 15105 858
rect 15285 809 15292 858
rect 15349 809 15361 861
rect 15413 858 15425 861
rect 15477 858 15489 861
rect 15541 858 15553 861
rect 15605 809 15617 861
rect 15669 858 15681 861
rect 15733 858 15745 861
rect 15797 858 15809 861
rect 15861 858 15873 861
rect 15676 809 15681 858
rect 15861 809 15866 858
rect 15925 809 15931 861
rect 15034 802 15043 809
rect 15099 802 15126 809
rect 15182 802 15209 809
rect 15265 802 15292 809
rect 15348 802 15374 809
rect 15430 802 15456 809
rect 15512 802 15538 809
rect 15594 802 15620 809
rect 15676 802 15702 809
rect 15758 802 15784 809
rect 15840 802 15866 809
rect 15922 802 15931 809
rect 15034 789 15931 802
rect 15034 737 15040 789
rect 15092 737 15105 789
rect 15157 737 15169 789
rect 15221 737 15233 789
rect 15285 737 15297 789
rect 15349 737 15361 789
rect 15413 737 15425 789
rect 15477 737 15489 789
rect 15541 737 15553 789
rect 15605 737 15617 789
rect 15669 737 15681 789
rect 15733 737 15745 789
rect 15797 737 15809 789
rect 15861 737 15873 789
rect 15925 737 15931 789
rect 15034 724 15931 737
rect 15034 717 15043 724
rect 15099 717 15126 724
rect 15182 717 15209 724
rect 15265 717 15292 724
rect 15348 717 15374 724
rect 15430 717 15456 724
rect 15512 717 15538 724
rect 15594 717 15620 724
rect 15676 717 15702 724
rect 15758 717 15784 724
rect 15840 717 15866 724
rect 15922 717 15931 724
rect 15034 665 15040 717
rect 15099 668 15105 717
rect 15285 668 15292 717
rect 15092 665 15105 668
rect 15157 665 15169 668
rect 15221 665 15233 668
rect 15285 665 15297 668
rect 15349 665 15361 717
rect 15413 665 15425 668
rect 15477 665 15489 668
rect 15541 665 15553 668
rect 15605 665 15617 717
rect 15676 668 15681 717
rect 15861 668 15866 717
rect 15669 665 15681 668
rect 15733 665 15745 668
rect 15797 665 15809 668
rect 15861 665 15873 668
rect 15925 665 15931 717
rect 15034 664 15931 665
rect 16875 861 17772 862
rect 16875 809 16881 861
rect 16933 858 16945 861
rect 16997 858 17009 861
rect 17061 858 17073 861
rect 17125 858 17137 861
rect 16940 809 16945 858
rect 17125 809 17130 858
rect 17189 809 17201 861
rect 17253 858 17265 861
rect 17317 858 17329 861
rect 17381 858 17393 861
rect 17445 809 17457 861
rect 17509 858 17521 861
rect 17573 858 17585 861
rect 17637 858 17649 861
rect 17701 858 17714 861
rect 17514 809 17521 858
rect 17701 809 17707 858
rect 17766 809 17772 861
rect 16875 802 16884 809
rect 16940 802 16966 809
rect 17022 802 17048 809
rect 17104 802 17130 809
rect 17186 802 17212 809
rect 17268 802 17294 809
rect 17350 802 17376 809
rect 17432 802 17458 809
rect 17514 802 17541 809
rect 17597 802 17624 809
rect 17680 802 17707 809
rect 17763 802 17772 809
rect 16875 789 17772 802
rect 16875 737 16881 789
rect 16933 737 16945 789
rect 16997 737 17009 789
rect 17061 737 17073 789
rect 17125 737 17137 789
rect 17189 737 17201 789
rect 17253 737 17265 789
rect 17317 737 17329 789
rect 17381 737 17393 789
rect 17445 737 17457 789
rect 17509 737 17521 789
rect 17573 737 17585 789
rect 17637 737 17649 789
rect 17701 737 17714 789
rect 17766 737 17772 789
rect 16875 724 17772 737
rect 16875 717 16884 724
rect 16940 717 16966 724
rect 17022 717 17048 724
rect 17104 717 17130 724
rect 17186 717 17212 724
rect 17268 717 17294 724
rect 17350 717 17376 724
rect 17432 717 17458 724
rect 17514 717 17541 724
rect 17597 717 17624 724
rect 17680 717 17707 724
rect 17763 717 17772 724
rect 16875 665 16881 717
rect 16940 668 16945 717
rect 17125 668 17130 717
rect 16933 665 16945 668
rect 16997 665 17009 668
rect 17061 665 17073 668
rect 17125 665 17137 668
rect 17189 665 17201 717
rect 17253 665 17265 668
rect 17317 665 17329 668
rect 17381 665 17393 668
rect 17445 665 17457 717
rect 17514 668 17521 717
rect 17701 668 17707 717
rect 17509 665 17521 668
rect 17573 665 17585 668
rect 17637 665 17649 668
rect 17701 665 17714 668
rect 17766 665 17772 717
rect 16875 664 17772 665
rect 19610 615 20058 621
rect 19662 563 20006 615
rect 19610 551 20058 563
rect 11434 547 12333 551
rect 11434 495 11440 547
rect 11500 495 11504 547
rect 11684 495 11687 547
rect 11748 495 11760 547
rect 12004 495 12014 547
rect 12070 495 12080 547
rect 12327 495 12333 547
rect 11434 491 11444 495
rect 11500 491 11525 495
rect 11581 491 11606 495
rect 11662 491 11687 495
rect 11743 491 11768 495
rect 11824 491 11850 495
rect 11906 491 11932 495
rect 11988 491 12014 495
rect 12070 491 12096 495
rect 12152 491 12178 495
rect 12234 491 12260 495
rect 12316 491 12333 495
rect 11434 479 12333 491
rect 11434 427 11440 479
rect 11492 463 11504 479
rect 11556 463 11568 479
rect 11620 463 11632 479
rect 11684 463 11696 479
rect 11500 427 11504 463
rect 11684 427 11687 463
rect 11748 427 11760 479
rect 11812 463 11824 479
rect 11876 463 11888 479
rect 11940 463 11952 479
rect 12004 463 12016 479
rect 12068 463 12080 479
rect 12132 463 12145 479
rect 12197 463 12210 479
rect 12262 463 12275 479
rect 12004 427 12014 463
rect 12070 427 12080 463
rect 12327 427 12333 479
rect 11434 411 11444 427
rect 11500 411 11525 427
rect 11581 411 11606 427
rect 11662 411 11687 427
rect 11743 411 11768 427
rect 11824 411 11850 427
rect 11906 411 11932 427
rect 11988 411 12014 427
rect 12070 411 12096 427
rect 12152 411 12178 427
rect 12234 411 12260 427
rect 12316 411 12333 427
rect 11434 359 11440 411
rect 11500 407 11504 411
rect 11684 407 11687 411
rect 11492 379 11504 407
rect 11556 379 11568 407
rect 11620 379 11632 407
rect 11684 379 11696 407
rect 11500 359 11504 379
rect 11684 359 11687 379
rect 11748 359 11760 411
rect 12004 407 12014 411
rect 12070 407 12080 411
rect 11812 379 11824 407
rect 11876 379 11888 407
rect 11940 379 11952 407
rect 12004 379 12016 407
rect 12068 379 12080 407
rect 12132 379 12145 407
rect 12197 379 12210 407
rect 12262 379 12275 407
rect 12004 359 12014 379
rect 12070 359 12080 379
rect 12327 359 12333 411
rect 11434 343 11444 359
rect 11500 343 11525 359
rect 11581 343 11606 359
rect 11662 343 11687 359
rect 11743 343 11768 359
rect 11824 343 11850 359
rect 11906 343 11932 359
rect 11988 343 12014 359
rect 12070 343 12096 359
rect 12152 343 12178 359
rect 12234 343 12260 359
rect 12316 343 12333 359
rect 11434 291 11440 343
rect 11500 323 11504 343
rect 11684 323 11687 343
rect 11492 295 11504 323
rect 11556 295 11568 323
rect 11620 295 11632 323
rect 11684 295 11696 323
rect 11500 291 11504 295
rect 11684 291 11687 295
rect 11748 291 11760 343
rect 12004 323 12014 343
rect 12070 323 12080 343
rect 11812 295 11824 323
rect 11876 295 11888 323
rect 11940 295 11952 323
rect 12004 295 12016 323
rect 12068 295 12080 323
rect 12132 295 12145 323
rect 12197 295 12210 323
rect 12262 295 12275 323
rect 12004 291 12014 295
rect 12070 291 12080 295
rect 12327 291 12333 343
rect 11434 275 11444 291
rect 11500 275 11525 291
rect 11581 275 11606 291
rect 11662 275 11687 291
rect 11743 275 11768 291
rect 11824 275 11850 291
rect 11906 275 11932 291
rect 11988 275 12014 291
rect 12070 275 12096 291
rect 12152 275 12178 291
rect 12234 275 12260 291
rect 12316 275 12333 291
rect 11434 223 11440 275
rect 11500 239 11504 275
rect 11684 239 11687 275
rect 11492 223 11504 239
rect 11556 223 11568 239
rect 11620 223 11632 239
rect 11684 223 11696 239
rect 11748 223 11760 275
rect 12004 239 12014 275
rect 12070 239 12080 275
rect 11812 223 11824 239
rect 11876 223 11888 239
rect 11940 223 11952 239
rect 12004 223 12016 239
rect 12068 223 12080 239
rect 12132 223 12145 239
rect 12197 223 12210 239
rect 12262 223 12275 239
rect 12327 223 12333 275
rect 11434 211 12333 223
rect 11434 207 11444 211
rect 11500 207 11525 211
rect 11581 207 11606 211
rect 11662 207 11687 211
rect 11743 207 11768 211
rect 11824 207 11850 211
rect 11906 207 11932 211
rect 11988 207 12014 211
rect 12070 207 12096 211
rect 12152 207 12178 211
rect 12234 207 12260 211
rect 12316 207 12333 211
rect 11434 155 11440 207
rect 11500 155 11504 207
rect 11684 155 11687 207
rect 11748 155 11760 207
rect 12004 155 12014 207
rect 12070 155 12080 207
rect 12327 155 12333 207
rect 11434 151 12333 155
rect 13989 547 14888 551
rect 13989 495 13995 547
rect 14242 495 14252 547
rect 14308 495 14318 547
rect 14562 495 14574 547
rect 14635 495 14638 547
rect 14818 495 14822 547
rect 14882 495 14888 547
rect 13989 491 14006 495
rect 14062 491 14088 495
rect 14144 491 14170 495
rect 14226 491 14252 495
rect 14308 491 14334 495
rect 14390 491 14416 495
rect 14472 491 14498 495
rect 14554 491 14579 495
rect 14635 491 14660 495
rect 14716 491 14741 495
rect 14797 491 14822 495
rect 14878 491 14888 495
rect 13989 479 14888 491
rect 13989 427 13995 479
rect 14047 463 14060 479
rect 14112 463 14125 479
rect 14177 463 14190 479
rect 14242 463 14254 479
rect 14306 463 14318 479
rect 14370 463 14382 479
rect 14434 463 14446 479
rect 14498 463 14510 479
rect 14242 427 14252 463
rect 14308 427 14318 463
rect 14562 427 14574 479
rect 14626 463 14638 479
rect 14690 463 14702 479
rect 14754 463 14766 479
rect 14818 463 14830 479
rect 14635 427 14638 463
rect 14818 427 14822 463
rect 14882 427 14888 479
rect 13989 411 14006 427
rect 14062 411 14088 427
rect 14144 411 14170 427
rect 14226 411 14252 427
rect 14308 411 14334 427
rect 14390 411 14416 427
rect 14472 411 14498 427
rect 14554 411 14579 427
rect 14635 411 14660 427
rect 14716 411 14741 427
rect 14797 411 14822 427
rect 14878 411 14888 427
rect 13989 359 13995 411
rect 14242 407 14252 411
rect 14308 407 14318 411
rect 14047 379 14060 407
rect 14112 379 14125 407
rect 14177 379 14190 407
rect 14242 379 14254 407
rect 14306 379 14318 407
rect 14370 379 14382 407
rect 14434 379 14446 407
rect 14498 379 14510 407
rect 14242 359 14252 379
rect 14308 359 14318 379
rect 14562 359 14574 411
rect 14635 407 14638 411
rect 14818 407 14822 411
rect 14626 379 14638 407
rect 14690 379 14702 407
rect 14754 379 14766 407
rect 14818 379 14830 407
rect 14635 359 14638 379
rect 14818 359 14822 379
rect 14882 359 14888 411
rect 13989 343 14006 359
rect 14062 343 14088 359
rect 14144 343 14170 359
rect 14226 343 14252 359
rect 14308 343 14334 359
rect 14390 343 14416 359
rect 14472 343 14498 359
rect 14554 343 14579 359
rect 14635 343 14660 359
rect 14716 343 14741 359
rect 14797 343 14822 359
rect 14878 343 14888 359
rect 13989 291 13995 343
rect 14242 323 14252 343
rect 14308 323 14318 343
rect 14047 295 14060 323
rect 14112 295 14125 323
rect 14177 295 14190 323
rect 14242 295 14254 323
rect 14306 295 14318 323
rect 14370 295 14382 323
rect 14434 295 14446 323
rect 14498 295 14510 323
rect 14242 291 14252 295
rect 14308 291 14318 295
rect 14562 291 14574 343
rect 14635 323 14638 343
rect 14818 323 14822 343
rect 14626 295 14638 323
rect 14690 295 14702 323
rect 14754 295 14766 323
rect 14818 295 14830 323
rect 14635 291 14638 295
rect 14818 291 14822 295
rect 14882 291 14888 343
rect 13989 275 14006 291
rect 14062 275 14088 291
rect 14144 275 14170 291
rect 14226 275 14252 291
rect 14308 275 14334 291
rect 14390 275 14416 291
rect 14472 275 14498 291
rect 14554 275 14579 291
rect 14635 275 14660 291
rect 14716 275 14741 291
rect 14797 275 14822 291
rect 14878 275 14888 291
rect 13989 223 13995 275
rect 14242 239 14252 275
rect 14308 239 14318 275
rect 14047 223 14060 239
rect 14112 223 14125 239
rect 14177 223 14190 239
rect 14242 223 14254 239
rect 14306 223 14318 239
rect 14370 223 14382 239
rect 14434 223 14446 239
rect 14498 223 14510 239
rect 14562 223 14574 275
rect 14635 239 14638 275
rect 14818 239 14822 275
rect 14626 223 14638 239
rect 14690 223 14702 239
rect 14754 223 14766 239
rect 14818 223 14830 239
rect 14882 223 14888 275
rect 13989 211 14888 223
rect 13989 207 14006 211
rect 14062 207 14088 211
rect 14144 207 14170 211
rect 14226 207 14252 211
rect 14308 207 14334 211
rect 14390 207 14416 211
rect 14472 207 14498 211
rect 14554 207 14579 211
rect 14635 207 14660 211
rect 14716 207 14741 211
rect 14797 207 14822 211
rect 14878 207 14888 211
rect 13989 155 13995 207
rect 14242 155 14252 207
rect 14308 155 14318 207
rect 14562 155 14574 207
rect 14635 155 14638 207
rect 14818 155 14822 207
rect 14882 155 14888 207
rect 13989 151 14888 155
rect 17918 547 18817 551
rect 17918 495 17924 547
rect 17984 495 17988 547
rect 18168 495 18171 547
rect 18232 495 18244 547
rect 18488 495 18498 547
rect 18554 495 18564 547
rect 18811 495 18817 547
rect 17918 491 17928 495
rect 17984 491 18009 495
rect 18065 491 18090 495
rect 18146 491 18171 495
rect 18227 491 18252 495
rect 18308 491 18334 495
rect 18390 491 18416 495
rect 18472 491 18498 495
rect 18554 491 18580 495
rect 18636 491 18662 495
rect 18718 491 18744 495
rect 18800 491 18817 495
rect 19662 499 20006 551
rect 19610 493 20058 499
rect 17918 479 18817 491
rect 17918 427 17924 479
rect 17976 463 17988 479
rect 18040 463 18052 479
rect 18104 463 18116 479
rect 18168 463 18180 479
rect 17984 427 17988 463
rect 18168 427 18171 463
rect 18232 427 18244 479
rect 18296 463 18308 479
rect 18360 463 18372 479
rect 18424 463 18436 479
rect 18488 463 18500 479
rect 18552 463 18564 479
rect 18616 463 18629 479
rect 18681 463 18694 479
rect 18746 463 18759 479
rect 18488 427 18498 463
rect 18554 427 18564 463
rect 18811 427 18817 479
rect 17918 411 17928 427
rect 17984 411 18009 427
rect 18065 411 18090 427
rect 18146 411 18171 427
rect 18227 411 18252 427
rect 18308 411 18334 427
rect 18390 411 18416 427
rect 18472 411 18498 427
rect 18554 411 18580 427
rect 18636 411 18662 427
rect 18718 411 18744 427
rect 18800 411 18817 427
rect 17918 359 17924 411
rect 17984 407 17988 411
rect 18168 407 18171 411
rect 17976 379 17988 407
rect 18040 379 18052 407
rect 18104 379 18116 407
rect 18168 379 18180 407
rect 17984 359 17988 379
rect 18168 359 18171 379
rect 18232 359 18244 411
rect 18488 407 18498 411
rect 18554 407 18564 411
rect 18296 379 18308 407
rect 18360 379 18372 407
rect 18424 379 18436 407
rect 18488 379 18500 407
rect 18552 379 18564 407
rect 18616 379 18629 407
rect 18681 379 18694 407
rect 18746 379 18759 407
rect 18488 359 18498 379
rect 18554 359 18564 379
rect 18811 359 18817 411
rect 17918 343 17928 359
rect 17984 343 18009 359
rect 18065 343 18090 359
rect 18146 343 18171 359
rect 18227 343 18252 359
rect 18308 343 18334 359
rect 18390 343 18416 359
rect 18472 343 18498 359
rect 18554 343 18580 359
rect 18636 343 18662 359
rect 18718 343 18744 359
rect 18800 343 18817 359
rect 17918 291 17924 343
rect 17984 323 17988 343
rect 18168 323 18171 343
rect 17976 295 17988 323
rect 18040 295 18052 323
rect 18104 295 18116 323
rect 18168 295 18180 323
rect 17984 291 17988 295
rect 18168 291 18171 295
rect 18232 291 18244 343
rect 18488 323 18498 343
rect 18554 323 18564 343
rect 18296 295 18308 323
rect 18360 295 18372 323
rect 18424 295 18436 323
rect 18488 295 18500 323
rect 18552 295 18564 323
rect 18616 295 18629 323
rect 18681 295 18694 323
rect 18746 295 18759 323
rect 18488 291 18498 295
rect 18554 291 18564 295
rect 18811 291 18817 343
rect 17918 275 17928 291
rect 17984 275 18009 291
rect 18065 275 18090 291
rect 18146 275 18171 291
rect 18227 275 18252 291
rect 18308 275 18334 291
rect 18390 275 18416 291
rect 18472 275 18498 291
rect 18554 275 18580 291
rect 18636 275 18662 291
rect 18718 275 18744 291
rect 18800 275 18817 291
rect 17918 223 17924 275
rect 17984 239 17988 275
rect 18168 239 18171 275
rect 17976 223 17988 239
rect 18040 223 18052 239
rect 18104 223 18116 239
rect 18168 223 18180 239
rect 18232 223 18244 275
rect 18488 239 18498 275
rect 18554 239 18564 275
rect 18296 223 18308 239
rect 18360 223 18372 239
rect 18424 223 18436 239
rect 18488 223 18500 239
rect 18552 223 18564 239
rect 18616 223 18629 239
rect 18681 223 18694 239
rect 18746 223 18759 239
rect 18811 223 18817 275
tri 20004 240 20006 242 se
rect 20006 240 20058 242
rect 17918 211 18817 223
rect 17918 207 17928 211
rect 17984 207 18009 211
rect 18065 207 18090 211
rect 18146 207 18171 211
rect 18227 207 18252 211
rect 18308 207 18334 211
rect 18390 207 18416 211
rect 18472 207 18498 211
rect 18554 207 18580 211
rect 18636 207 18662 211
rect 18718 207 18744 211
rect 18800 207 18817 211
rect 17918 155 17924 207
rect 17984 155 17988 207
rect 18168 155 18171 207
rect 18232 155 18244 207
rect 18488 155 18498 207
rect 18554 155 18564 207
rect 18811 155 18817 207
rect 17918 151 18817 155
rect 19610 203 19890 240
rect 19662 200 19890 203
rect 19891 201 19892 239
rect 19952 201 19953 239
rect 19954 234 20058 240
rect 19954 200 20006 234
tri 19662 185 19677 200 nw
tri 19967 185 19982 200 ne
rect 19982 185 20006 200
tri 19982 182 19985 185 ne
rect 19985 182 20006 185
tri 19985 170 19997 182 ne
rect 19997 170 20058 182
tri 19997 161 20006 170 ne
rect 19610 139 19662 151
rect 20006 112 20058 118
rect 20430 222 20482 228
rect 20430 158 20482 170
rect 9898 -12 9948 -11
rect 9897 -72 9949 -12
rect 9898 -73 9948 -72
rect 6943 -229 7342 -211
rect 6943 -281 6949 -229
rect 7001 -239 7016 -229
rect 7068 -239 7083 -229
rect 7135 -239 7150 -229
rect 7202 -239 7217 -229
rect 7269 -239 7284 -229
rect 7008 -281 7016 -239
rect 7269 -281 7277 -239
rect 7336 -281 7342 -229
rect 6943 -295 6952 -281
rect 7008 -295 7034 -281
rect 7090 -295 7115 -281
rect 7171 -295 7196 -281
rect 7252 -295 7277 -281
rect 7333 -295 7342 -281
tri 9892 -293 9897 -288 se
rect 9897 -293 9949 -74
rect 10391 38 11288 39
rect 10391 -14 10397 38
rect 10449 35 10462 38
rect 10514 35 10526 38
rect 10578 35 10590 38
rect 10642 35 10654 38
rect 10456 -14 10462 35
rect 10642 -14 10646 35
rect 10706 -14 10718 38
rect 10770 35 10782 38
rect 10834 35 10846 38
rect 10898 35 10910 38
rect 10962 -14 10974 38
rect 11026 35 11038 38
rect 11090 35 11102 38
rect 11154 35 11166 38
rect 11218 35 11230 38
rect 11030 -14 11038 35
rect 11218 -14 11223 35
rect 11282 -14 11288 38
rect 15034 37 15931 38
rect 10391 -21 10400 -14
rect 10456 -21 10482 -14
rect 10538 -21 10564 -14
rect 10620 -21 10646 -14
rect 10702 -21 10728 -14
rect 10784 -21 10810 -14
rect 10866 -21 10892 -14
rect 10948 -21 10974 -14
rect 11030 -21 11057 -14
rect 11113 -21 11140 -14
rect 11196 -21 11223 -14
rect 11279 -21 11288 -14
rect 10391 -34 11288 -21
rect 10391 -86 10397 -34
rect 10449 -86 10462 -34
rect 10514 -86 10526 -34
rect 10578 -86 10590 -34
rect 10642 -86 10654 -34
rect 10706 -86 10718 -34
rect 10770 -86 10782 -34
rect 10834 -86 10846 -34
rect 10898 -86 10910 -34
rect 10962 -86 10974 -34
rect 11026 -86 11038 -34
rect 11090 -86 11102 -34
rect 11154 -86 11166 -34
rect 11218 -86 11230 -34
rect 11282 -86 11288 -34
rect 10391 -99 11288 -86
rect 10391 -106 10400 -99
rect 10456 -106 10482 -99
rect 10538 -106 10564 -99
rect 10620 -106 10646 -99
rect 10702 -106 10728 -99
rect 10784 -106 10810 -99
rect 10866 -106 10892 -99
rect 10948 -106 10974 -99
rect 11030 -106 11057 -99
rect 11113 -106 11140 -99
rect 11196 -106 11223 -99
rect 11279 -106 11288 -99
rect 10391 -158 10397 -106
rect 10456 -155 10462 -106
rect 10642 -155 10646 -106
rect 10449 -158 10462 -155
rect 10514 -158 10526 -155
rect 10578 -158 10590 -155
rect 10642 -158 10654 -155
rect 10706 -158 10718 -106
rect 10770 -158 10782 -155
rect 10834 -158 10846 -155
rect 10898 -158 10910 -155
rect 10962 -158 10974 -106
rect 11030 -155 11038 -106
rect 11218 -155 11223 -106
rect 11026 -158 11038 -155
rect 11090 -158 11102 -155
rect 11154 -158 11166 -155
rect 11218 -158 11230 -155
rect 11282 -158 11288 -106
rect 11915 -22 11924 34
rect 11980 -22 12005 34
rect 12061 -22 12086 34
rect 12142 -22 12167 34
rect 12223 -22 12249 34
rect 12305 -22 12331 34
rect 12387 -22 12396 34
rect 11915 -100 12396 -22
rect 11915 -156 11924 -100
rect 11980 -156 12005 -100
rect 12061 -156 12086 -100
rect 12142 -156 12167 -100
rect 12223 -156 12249 -100
rect 12305 -156 12331 -100
rect 12387 -156 12396 -100
rect 15034 -15 15040 37
rect 15092 34 15105 37
rect 15157 34 15169 37
rect 15221 34 15233 37
rect 15285 34 15297 37
rect 15099 -15 15105 34
rect 15285 -15 15292 34
rect 15349 -15 15361 37
rect 15413 34 15425 37
rect 15477 34 15489 37
rect 15541 34 15553 37
rect 15605 -15 15617 37
rect 15669 34 15681 37
rect 15733 34 15745 37
rect 15797 34 15809 37
rect 15861 34 15873 37
rect 15676 -15 15681 34
rect 15861 -15 15866 34
rect 15925 -15 15931 37
rect 15034 -22 15043 -15
rect 15099 -22 15126 -15
rect 15182 -22 15209 -15
rect 15265 -22 15292 -15
rect 15348 -22 15374 -15
rect 15430 -22 15456 -15
rect 15512 -22 15538 -15
rect 15594 -22 15620 -15
rect 15676 -22 15702 -15
rect 15758 -22 15784 -15
rect 15840 -22 15866 -15
rect 15922 -22 15931 -15
rect 15034 -35 15931 -22
rect 15034 -87 15040 -35
rect 15092 -87 15105 -35
rect 15157 -87 15169 -35
rect 15221 -87 15233 -35
rect 15285 -87 15297 -35
rect 15349 -87 15361 -35
rect 15413 -87 15425 -35
rect 15477 -87 15489 -35
rect 15541 -87 15553 -35
rect 15605 -87 15617 -35
rect 15669 -87 15681 -35
rect 15733 -87 15745 -35
rect 15797 -87 15809 -35
rect 15861 -87 15873 -35
rect 15925 -87 15931 -35
rect 15034 -100 15931 -87
rect 15034 -107 15043 -100
rect 15099 -107 15126 -100
rect 15182 -107 15209 -100
rect 15265 -107 15292 -100
rect 15348 -107 15374 -100
rect 15430 -107 15456 -100
rect 15512 -107 15538 -100
rect 15594 -107 15620 -100
rect 15676 -107 15702 -100
rect 15758 -107 15784 -100
rect 15840 -107 15866 -100
rect 15922 -107 15931 -100
rect 10391 -159 11288 -158
rect 12496 -211 12505 -155
rect 12561 -211 12587 -155
rect 12643 -211 12668 -155
rect 12724 -211 12749 -155
rect 12805 -211 12830 -155
rect 12886 -211 12895 -155
rect 12496 -228 12895 -211
rect 12496 -280 12502 -228
rect 12554 -239 12569 -228
rect 12621 -239 12636 -228
rect 12688 -239 12703 -228
rect 12755 -239 12770 -228
rect 12822 -239 12837 -228
rect 12561 -280 12569 -239
rect 12822 -280 12830 -239
rect 12889 -280 12895 -228
tri 9949 -293 9954 -288 sw
tri 9890 -295 9892 -293 se
rect 9892 -295 9954 -293
tri 9860 -325 9890 -295 se
rect 9890 -325 9954 -295
tri 9954 -325 9986 -293 sw
rect 12496 -295 12505 -280
rect 12561 -295 12587 -280
rect 12643 -295 12668 -280
rect 12724 -295 12749 -280
rect 12805 -295 12830 -280
rect 12886 -295 12895 -280
rect 13427 -211 13436 -155
rect 13492 -211 13518 -155
rect 13574 -211 13599 -155
rect 13655 -211 13680 -155
rect 13736 -211 13761 -155
rect 13817 -211 13826 -155
rect 15034 -159 15040 -107
rect 15099 -156 15105 -107
rect 15285 -156 15292 -107
rect 15092 -159 15105 -156
rect 15157 -159 15169 -156
rect 15221 -159 15233 -156
rect 15285 -159 15297 -156
rect 15349 -159 15361 -107
rect 15413 -159 15425 -156
rect 15477 -159 15489 -156
rect 15541 -159 15553 -156
rect 15605 -159 15617 -107
rect 15676 -156 15681 -107
rect 15861 -156 15866 -107
rect 15669 -159 15681 -156
rect 15733 -159 15745 -156
rect 15797 -159 15809 -156
rect 15861 -159 15873 -156
rect 15925 -159 15931 -107
rect 15034 -160 15931 -159
rect 16875 37 17772 38
rect 16875 -15 16881 37
rect 16933 34 16946 37
rect 16998 34 17010 37
rect 17062 34 17074 37
rect 17126 34 17138 37
rect 16940 -15 16946 34
rect 17126 -15 17133 34
rect 17190 -15 17202 37
rect 17254 34 17266 37
rect 17318 34 17330 37
rect 17382 34 17394 37
rect 17446 -15 17458 37
rect 17510 34 17522 37
rect 17574 34 17586 37
rect 17638 34 17650 37
rect 17702 34 17714 37
rect 17517 -15 17522 34
rect 17702 -15 17707 34
rect 17766 -15 17772 37
rect 16875 -22 16884 -15
rect 16940 -22 16967 -15
rect 17023 -22 17050 -15
rect 17106 -22 17133 -15
rect 17189 -22 17215 -15
rect 17271 -22 17297 -15
rect 17353 -22 17379 -15
rect 17435 -22 17461 -15
rect 17517 -22 17543 -15
rect 17599 -22 17625 -15
rect 17681 -22 17707 -15
rect 17763 -22 17772 -15
rect 16875 -35 17772 -22
rect 16875 -87 16881 -35
rect 16933 -87 16946 -35
rect 16998 -87 17010 -35
rect 17062 -87 17074 -35
rect 17126 -87 17138 -35
rect 17190 -87 17202 -35
rect 17254 -87 17266 -35
rect 17318 -87 17330 -35
rect 17382 -87 17394 -35
rect 17446 -87 17458 -35
rect 17510 -87 17522 -35
rect 17574 -87 17586 -35
rect 17638 -87 17650 -35
rect 17702 -87 17714 -35
rect 17766 -87 17772 -35
rect 16875 -100 17772 -87
rect 16875 -107 16884 -100
rect 16940 -107 16967 -100
rect 17023 -107 17050 -100
rect 17106 -107 17133 -100
rect 17189 -107 17215 -100
rect 17271 -107 17297 -100
rect 17353 -107 17379 -100
rect 17435 -107 17461 -100
rect 17517 -107 17543 -100
rect 17599 -107 17625 -100
rect 17681 -107 17707 -100
rect 17763 -107 17772 -100
rect 19610 30 19662 87
tri 20416 81 20430 95 se
rect 20430 81 20482 106
tri 22907 81 22930 104 se
rect 22930 81 23046 4619
tri 20406 71 20416 81 se
rect 20416 71 20482 81
rect 20006 63 20482 71
tri 22889 63 22907 81 se
rect 22907 63 23046 81
tri 20005 31 20006 32 se
tri 20004 30 20005 31 se
rect 20005 30 20006 31
tri 20003 29 20004 30 se
rect 20004 29 20006 30
rect 19611 28 19661 29
tri 20002 28 20003 29 se
rect 20003 28 20006 29
rect 19610 -32 19662 28
tri 19985 11 20002 28 se
rect 20002 11 20006 28
rect 20058 34 20482 63
rect 20058 11 20072 34
tri 19973 -1 19985 11 se
rect 19985 8 20072 11
tri 20072 8 20098 34 nw
tri 20404 8 20430 34 ne
rect 20430 8 20482 34
rect 22755 57 23046 63
rect 19985 -1 20058 8
tri 19964 -10 19973 -1 se
rect 19973 -10 20006 -1
rect 19611 -33 19661 -32
rect 19610 -48 19662 -34
rect 19759 -18 20006 -10
rect 19610 -70 19759 -48
rect 19811 -50 20006 -18
rect 19811 -53 19861 -50
tri 19861 -53 19864 -50 nw
tri 19973 -53 19976 -50 ne
rect 19976 -53 20006 -50
tri 20058 -6 20072 8 nw
rect 19811 -59 19855 -53
tri 19855 -59 19861 -53 nw
tri 19976 -59 19982 -53 ne
rect 19982 -59 20058 -53
rect 19811 -70 19813 -59
rect 19610 -82 19813 -70
rect 19610 -101 19759 -82
rect 16875 -159 16881 -107
rect 16940 -156 16946 -107
rect 17126 -156 17133 -107
rect 16933 -159 16946 -156
rect 16998 -159 17010 -156
rect 17062 -159 17074 -156
rect 17126 -159 17138 -156
rect 17190 -159 17202 -107
rect 17254 -159 17266 -156
rect 17318 -159 17330 -156
rect 17382 -159 17394 -156
rect 17446 -159 17458 -107
rect 17517 -156 17522 -107
rect 17702 -156 17707 -107
rect 17510 -159 17522 -156
rect 17574 -159 17586 -156
rect 17638 -159 17650 -156
rect 17702 -159 17714 -156
rect 17766 -159 17772 -107
rect 19811 -101 19813 -82
tri 19813 -101 19855 -59 nw
tri 19982 -83 20006 -59 ne
tri 19811 -103 19813 -101 nw
rect 19759 -140 19811 -134
rect 16875 -160 17772 -159
rect 13427 -229 13826 -211
rect 13427 -281 13433 -229
rect 13485 -239 13500 -229
rect 13552 -239 13567 -229
rect 13619 -239 13634 -229
rect 13686 -239 13701 -229
rect 13753 -239 13768 -229
rect 13492 -281 13500 -239
rect 13753 -281 13761 -239
rect 13820 -281 13826 -229
rect 13427 -295 13436 -281
rect 13492 -295 13518 -281
rect 13574 -295 13599 -281
rect 13655 -295 13680 -281
rect 13736 -295 13761 -281
rect 13817 -295 13826 -281
rect 19065 -211 19074 -155
rect 19130 -211 19154 -155
rect 19210 -211 19234 -155
rect 19290 -211 19314 -155
rect 19370 -211 19379 -155
rect 19065 -229 19379 -211
rect 19065 -281 19071 -229
rect 19123 -239 19155 -229
rect 19207 -239 19238 -229
rect 19290 -239 19321 -229
rect 19065 -295 19074 -281
rect 19130 -295 19154 -239
rect 19210 -295 19234 -239
rect 19290 -295 19314 -239
rect 19373 -281 19379 -229
rect 19370 -295 19379 -281
tri 19995 -295 20006 -284 se
rect 20006 -295 20058 -59
rect 22871 -16 23046 57
rect 22871 -59 22997 -16
rect 22755 -65 22997 -59
tri 22997 -65 23046 -16 nw
tri 19965 -325 19995 -295 se
rect 19995 -325 20058 -295
rect 3708 -469 3714 -417
rect 3766 -469 3778 -417
rect 3830 -469 3836 -417
tri 4053 -388 4116 -325 se
rect 4116 -377 20058 -325
rect 4116 -388 4127 -377
tri 4127 -388 4138 -377 nw
rect 4053 -399 4116 -388
tri 4116 -399 4127 -388 nw
tri 3497 -500 3502 -495 ne
rect 3502 -500 3549 -495
tri 3549 -500 3576 -473 sw
tri 4026 -500 4053 -473 se
rect 4053 -495 4105 -399
tri 4105 -410 4116 -399 nw
rect 4053 -500 4100 -495
tri 4100 -500 4105 -495 nw
tri 3502 -546 3548 -500 ne
rect 3548 -546 4054 -500
tri 4054 -546 4100 -500 nw
tri -899 -1926 -847 -1874 nw
tri -1035 -1994 -967 -1926 se
tri -967 -1994 -899 -1926 nw
tri -1103 -2062 -1035 -1994 se
tri -1035 -2062 -967 -1994 nw
tri -1171 -2130 -1103 -2062 se
tri -1103 -2130 -1035 -2062 nw
tri -1239 -2198 -1171 -2130 se
tri -1171 -2198 -1103 -2130 nw
tri -1307 -2266 -1239 -2198 se
tri -1239 -2266 -1171 -2198 nw
tri -1375 -2334 -1307 -2266 se
tri -1307 -2334 -1239 -2266 nw
tri -1379 -2338 -1375 -2334 se
rect -1375 -2338 -1311 -2334
tri -1311 -2338 -1307 -2334 nw
rect -1379 -2554 -1318 -2338
tri -1318 -2345 -1311 -2338 nw
rect 15039 -2810 15048 -2754
rect 15104 -2810 15129 -2754
rect 15185 -2810 15210 -2754
rect 15266 -2810 15291 -2754
rect 15347 -2810 15372 -2754
rect 15428 -2810 15453 -2754
rect 15509 -2810 15534 -2754
rect 15590 -2810 15614 -2754
rect 15670 -2810 15694 -2754
rect 15750 -2810 15774 -2754
rect 15830 -2810 15854 -2754
rect 15910 -2810 15919 -2754
rect 15039 -2862 15919 -2810
rect 15039 -2871 15048 -2862
rect 15104 -2871 15129 -2862
rect 15185 -2871 15210 -2862
rect 15266 -2871 15291 -2862
rect 15347 -2871 15372 -2862
rect 15428 -2871 15453 -2862
rect 15509 -2871 15534 -2862
rect 15590 -2871 15614 -2862
rect 15670 -2871 15694 -2862
rect 15750 -2871 15774 -2862
rect 15830 -2871 15854 -2862
rect 15910 -2871 15919 -2862
rect 15039 -2923 15045 -2871
rect 15104 -2918 15113 -2871
rect 15369 -2918 15372 -2871
rect 15097 -2923 15113 -2918
rect 15165 -2923 15181 -2918
rect 15233 -2923 15249 -2918
rect 15301 -2923 15317 -2918
rect 15369 -2923 15385 -2918
rect 15437 -2923 15453 -2871
rect 15509 -2918 15521 -2871
rect 15845 -2918 15854 -2871
rect 15505 -2923 15521 -2918
rect 15573 -2923 15589 -2918
rect 15641 -2923 15657 -2918
rect 15709 -2923 15725 -2918
rect 15777 -2923 15793 -2918
rect 15845 -2923 15861 -2918
rect 15913 -2923 15919 -2871
rect 16880 -2810 16889 -2754
rect 16945 -2810 16970 -2754
rect 17026 -2810 17051 -2754
rect 17107 -2810 17132 -2754
rect 17188 -2810 17213 -2754
rect 17269 -2810 17294 -2754
rect 17350 -2810 17375 -2754
rect 17431 -2810 17455 -2754
rect 17511 -2810 17535 -2754
rect 17591 -2810 17615 -2754
rect 17671 -2810 17695 -2754
rect 17751 -2810 17760 -2754
rect 16880 -2862 17760 -2810
rect 16880 -2871 16889 -2862
rect 16945 -2871 16970 -2862
rect 17026 -2871 17051 -2862
rect 17107 -2871 17132 -2862
rect 17188 -2871 17213 -2862
rect 17269 -2871 17294 -2862
rect 17350 -2871 17375 -2862
rect 17431 -2871 17455 -2862
rect 17511 -2871 17535 -2862
rect 17591 -2871 17615 -2862
rect 17671 -2871 17695 -2862
rect 17751 -2871 17760 -2862
rect 16880 -2923 16886 -2871
rect 16945 -2918 16954 -2871
rect 17210 -2918 17213 -2871
rect 16938 -2923 16954 -2918
rect 17006 -2923 17022 -2918
rect 17074 -2923 17090 -2918
rect 17142 -2923 17158 -2918
rect 17210 -2923 17226 -2918
rect 17278 -2923 17294 -2871
rect 17350 -2918 17362 -2871
rect 17686 -2918 17695 -2871
rect 17346 -2923 17362 -2918
rect 17414 -2923 17430 -2918
rect 17482 -2923 17498 -2918
rect 17550 -2923 17566 -2918
rect 17618 -2923 17634 -2918
rect 17686 -2923 17702 -2918
rect 17754 -2923 17760 -2871
<< rmetal2 >>
rect 50 240 52 241
rect 50 202 51 240
rect 50 201 52 202
rect 112 240 114 241
rect 113 202 114 240
rect 112 201 114 202
rect -1 120 1 121
rect 61 120 63 121
rect -1 82 0 120
rect 62 82 63 120
rect -1 81 1 82
rect 61 81 63 82
rect 19890 1451 19892 1452
rect 19890 1413 19891 1451
rect 19890 1412 19892 1413
rect 19952 1451 19954 1452
rect 19953 1413 19954 1451
rect 19952 1412 19954 1413
rect 19610 1257 19662 1258
rect 19610 1256 19611 1257
rect 19661 1256 19662 1257
rect 19610 1195 19611 1196
rect 19661 1195 19662 1196
rect 19610 1194 19662 1195
rect 19890 239 19892 240
rect 19890 201 19891 239
rect 19890 200 19892 201
rect 19952 239 19954 240
rect 19953 201 19954 239
rect 19952 200 19954 201
rect 9897 -11 9949 -10
rect 9897 -12 9898 -11
rect 9948 -12 9949 -11
rect 9897 -73 9898 -72
rect 9948 -73 9949 -72
rect 9897 -74 9949 -73
rect 19610 29 19662 30
rect 19610 28 19611 29
rect 19661 28 19662 29
rect 19610 -33 19611 -32
rect 19661 -33 19662 -32
rect 19610 -34 19662 -33
<< via2 >>
rect 19675 5499 19731 5501
rect 19755 5499 19811 5501
rect 19675 5447 19690 5499
rect 19690 5447 19731 5499
rect 19755 5447 19806 5499
rect 19806 5447 19811 5499
rect 19675 5445 19731 5447
rect 19755 5445 19811 5447
rect 3033 5079 3081 5128
rect 3081 5079 3089 5128
rect 3115 5079 3147 5128
rect 3147 5079 3161 5128
rect 3161 5079 3171 5128
rect 3197 5079 3213 5128
rect 3213 5079 3227 5128
rect 3227 5079 3253 5128
rect 3279 5079 3293 5128
rect 3293 5079 3335 5128
rect 3361 5079 3410 5128
rect 3410 5079 3417 5128
rect 3443 5079 3475 5128
rect 3475 5079 3488 5128
rect 3488 5079 3499 5128
rect 3525 5079 3540 5128
rect 3540 5079 3553 5128
rect 3553 5079 3581 5128
rect 3607 5079 3618 5128
rect 3618 5079 3663 5128
rect 3689 5079 3735 5128
rect 3735 5079 3745 5128
rect 3771 5079 3800 5128
rect 3800 5079 3813 5128
rect 3813 5079 3827 5128
rect 3853 5079 3865 5128
rect 3865 5079 3878 5128
rect 3878 5079 3909 5128
rect 3935 5079 3943 5128
rect 3943 5079 3991 5128
rect 4016 5079 4060 5128
rect 4060 5079 4072 5128
rect 4097 5079 4125 5128
rect 4125 5079 4138 5128
rect 4138 5079 4153 5128
rect 4178 5079 4190 5128
rect 4190 5079 4203 5128
rect 4203 5079 4234 5128
rect 4259 5079 4268 5128
rect 4268 5079 4315 5128
rect 3033 5072 3089 5079
rect 3115 5072 3171 5079
rect 3197 5072 3253 5079
rect 3279 5072 3335 5079
rect 3361 5072 3417 5079
rect 3443 5072 3499 5079
rect 3525 5072 3581 5079
rect 3607 5072 3663 5079
rect 3689 5072 3745 5079
rect 3771 5072 3827 5079
rect 3853 5072 3909 5079
rect 3935 5072 3991 5079
rect 4016 5072 4072 5079
rect 4097 5072 4153 5079
rect 4178 5072 4234 5079
rect 4259 5072 4315 5079
rect 3033 5015 3089 5020
rect 3115 5015 3171 5020
rect 3197 5015 3253 5020
rect 3279 5015 3335 5020
rect 3361 5015 3417 5020
rect 3443 5015 3499 5020
rect 3525 5015 3581 5020
rect 3607 5015 3663 5020
rect 3689 5015 3745 5020
rect 3771 5015 3827 5020
rect 3853 5015 3909 5020
rect 3935 5015 3991 5020
rect 4016 5015 4072 5020
rect 4097 5015 4153 5020
rect 4178 5015 4234 5020
rect 4259 5015 4315 5020
rect 3033 4964 3081 5015
rect 3081 4964 3089 5015
rect 3115 4964 3147 5015
rect 3147 4964 3161 5015
rect 3161 4964 3171 5015
rect 3197 4964 3213 5015
rect 3213 4964 3227 5015
rect 3227 4964 3253 5015
rect 3279 4964 3293 5015
rect 3293 4964 3335 5015
rect 3361 4964 3410 5015
rect 3410 4964 3417 5015
rect 3443 4964 3475 5015
rect 3475 4964 3488 5015
rect 3488 4964 3499 5015
rect 3525 4964 3540 5015
rect 3540 4964 3553 5015
rect 3553 4964 3581 5015
rect 3607 4964 3618 5015
rect 3618 4964 3663 5015
rect 3689 4964 3735 5015
rect 3735 4964 3745 5015
rect 3771 4964 3800 5015
rect 3800 4964 3813 5015
rect 3813 4964 3827 5015
rect 3853 4964 3865 5015
rect 3865 4964 3878 5015
rect 3878 4964 3909 5015
rect 3935 4964 3943 5015
rect 3943 4964 3991 5015
rect 4016 4964 4060 5015
rect 4060 4964 4072 5015
rect 4097 4964 4125 5015
rect 4125 4964 4138 5015
rect 4138 4964 4153 5015
rect 4178 4964 4190 5015
rect 4190 4964 4203 5015
rect 4203 4964 4234 5015
rect 4259 4964 4268 5015
rect 4268 4964 4315 5015
rect 9211 5079 9212 5128
rect 9212 5079 9226 5128
rect 9226 5079 9267 5128
rect 9296 5079 9344 5128
rect 9344 5079 9352 5128
rect 9381 5079 9410 5128
rect 9410 5079 9424 5128
rect 9424 5079 9437 5128
rect 9466 5079 9476 5128
rect 9476 5079 9490 5128
rect 9490 5079 9522 5128
rect 9550 5079 9556 5128
rect 9556 5079 9606 5128
rect 9211 5072 9267 5079
rect 9296 5072 9352 5079
rect 9381 5072 9437 5079
rect 9466 5072 9522 5079
rect 9550 5072 9606 5079
rect 9634 5072 9690 5128
rect 9718 5072 9774 5128
rect 9211 5015 9267 5020
rect 9296 5015 9352 5020
rect 9381 5015 9437 5020
rect 9466 5015 9522 5020
rect 9550 5015 9606 5020
rect 9211 4964 9212 5015
rect 9212 4964 9226 5015
rect 9226 4964 9267 5015
rect 9296 4964 9344 5015
rect 9344 4964 9352 5015
rect 9381 4964 9410 5015
rect 9410 4964 9424 5015
rect 9424 4964 9437 5015
rect 9466 4964 9476 5015
rect 9476 4964 9490 5015
rect 9490 4964 9522 5015
rect 9550 4964 9556 5015
rect 9556 4964 9606 5015
rect 9634 4964 9690 5020
rect 9718 4964 9774 5020
rect 11018 5079 11066 5128
rect 11066 5079 11074 5128
rect 11114 5079 11134 5128
rect 11134 5079 11150 5128
rect 11150 5079 11170 5128
rect 11209 5079 11217 5128
rect 11217 5079 11265 5128
rect 11018 5072 11074 5079
rect 11114 5072 11170 5079
rect 11209 5072 11265 5079
rect 11018 5015 11074 5020
rect 11114 5015 11170 5020
rect 11209 5015 11265 5020
rect 11018 4964 11066 5015
rect 11066 4964 11074 5015
rect 11114 4964 11134 5015
rect 11134 4964 11150 5015
rect 11150 4964 11170 5015
rect 11209 4964 11217 5015
rect 11217 4964 11265 5015
rect 15053 5079 15101 5128
rect 15101 5079 15109 5128
rect 15134 5079 15170 5128
rect 15170 5079 15187 5128
rect 15187 5079 15190 5128
rect 15215 5079 15239 5128
rect 15239 5079 15255 5128
rect 15255 5079 15271 5128
rect 15296 5079 15307 5128
rect 15307 5079 15323 5128
rect 15323 5079 15352 5128
rect 15377 5079 15391 5128
rect 15391 5079 15433 5128
rect 15458 5079 15459 5128
rect 15459 5079 15511 5128
rect 15511 5079 15514 5128
rect 15539 5079 15579 5128
rect 15579 5079 15595 5128
rect 15619 5079 15647 5128
rect 15647 5079 15663 5128
rect 15663 5079 15675 5128
rect 15699 5079 15715 5128
rect 15715 5079 15731 5128
rect 15731 5079 15755 5128
rect 15779 5079 15783 5128
rect 15783 5079 15799 5128
rect 15799 5079 15835 5128
rect 15859 5079 15867 5128
rect 15867 5079 15915 5128
rect 15053 5072 15109 5079
rect 15134 5072 15190 5079
rect 15215 5072 15271 5079
rect 15296 5072 15352 5079
rect 15377 5072 15433 5079
rect 15458 5072 15514 5079
rect 15539 5072 15595 5079
rect 15619 5072 15675 5079
rect 15699 5072 15755 5079
rect 15779 5072 15835 5079
rect 15859 5072 15915 5079
rect 15053 5015 15109 5020
rect 15134 5015 15190 5020
rect 15215 5015 15271 5020
rect 15296 5015 15352 5020
rect 15377 5015 15433 5020
rect 15458 5015 15514 5020
rect 15539 5015 15595 5020
rect 15619 5015 15675 5020
rect 15699 5015 15755 5020
rect 15779 5015 15835 5020
rect 15859 5015 15915 5020
rect 15053 4964 15101 5015
rect 15101 4964 15109 5015
rect 15134 4964 15170 5015
rect 15170 4964 15187 5015
rect 15187 4964 15190 5015
rect 15215 4964 15239 5015
rect 15239 4964 15255 5015
rect 15255 4964 15271 5015
rect 15296 4964 15307 5015
rect 15307 4964 15323 5015
rect 15323 4964 15352 5015
rect 15377 4964 15391 5015
rect 15391 4964 15433 5015
rect 15458 4964 15459 5015
rect 15459 4964 15511 5015
rect 15511 4964 15514 5015
rect 15539 4964 15579 5015
rect 15579 4964 15595 5015
rect 15619 4964 15647 5015
rect 15647 4964 15663 5015
rect 15663 4964 15675 5015
rect 15699 4964 15715 5015
rect 15715 4964 15731 5015
rect 15731 4964 15755 5015
rect 15779 4964 15783 5015
rect 15783 4964 15799 5015
rect 15799 4964 15835 5015
rect 15859 4964 15867 5015
rect 15867 4964 15915 5015
rect 16892 5079 16940 5128
rect 16940 5079 16948 5128
rect 16973 5079 17009 5128
rect 17009 5079 17026 5128
rect 17026 5079 17029 5128
rect 17054 5079 17078 5128
rect 17078 5079 17094 5128
rect 17094 5079 17110 5128
rect 17135 5079 17146 5128
rect 17146 5079 17162 5128
rect 17162 5079 17191 5128
rect 17216 5079 17230 5128
rect 17230 5079 17272 5128
rect 17297 5079 17298 5128
rect 17298 5079 17350 5128
rect 17350 5079 17353 5128
rect 17378 5079 17418 5128
rect 17418 5079 17434 5128
rect 17458 5079 17486 5128
rect 17486 5079 17502 5128
rect 17502 5079 17514 5128
rect 17538 5079 17554 5128
rect 17554 5079 17570 5128
rect 17570 5079 17594 5128
rect 17618 5079 17622 5128
rect 17622 5079 17638 5128
rect 17638 5079 17674 5128
rect 17698 5079 17706 5128
rect 17706 5079 17754 5128
rect 16892 5072 16948 5079
rect 16973 5072 17029 5079
rect 17054 5072 17110 5079
rect 17135 5072 17191 5079
rect 17216 5072 17272 5079
rect 17297 5072 17353 5079
rect 17378 5072 17434 5079
rect 17458 5072 17514 5079
rect 17538 5072 17594 5079
rect 17618 5072 17674 5079
rect 17698 5072 17754 5079
rect 16892 5015 16948 5020
rect 16973 5015 17029 5020
rect 17054 5015 17110 5020
rect 17135 5015 17191 5020
rect 17216 5015 17272 5020
rect 17297 5015 17353 5020
rect 17378 5015 17434 5020
rect 17458 5015 17514 5020
rect 17538 5015 17594 5020
rect 17618 5015 17674 5020
rect 17698 5015 17754 5020
rect 16892 4964 16940 5015
rect 16940 4964 16948 5015
rect 16973 4964 17009 5015
rect 17009 4964 17026 5015
rect 17026 4964 17029 5015
rect 17054 4964 17078 5015
rect 17078 4964 17094 5015
rect 17094 4964 17110 5015
rect 17135 4964 17146 5015
rect 17146 4964 17162 5015
rect 17162 4964 17191 5015
rect 17216 4964 17230 5015
rect 17230 4964 17272 5015
rect 17297 4964 17298 5015
rect 17298 4964 17350 5015
rect 17350 4964 17353 5015
rect 17378 4964 17418 5015
rect 17418 4964 17434 5015
rect 17458 4964 17486 5015
rect 17486 4964 17502 5015
rect 17502 4964 17514 5015
rect 17538 4964 17554 5015
rect 17554 4964 17570 5015
rect 17570 4964 17594 5015
rect 17618 4964 17622 5015
rect 17622 4964 17638 5015
rect 17638 4964 17674 5015
rect 17698 4964 17706 5015
rect 17706 4964 17754 5015
rect 19675 5079 19723 5128
rect 19723 5079 19731 5128
rect 19675 5072 19731 5079
rect 19755 5079 19762 5128
rect 19762 5079 19811 5128
rect 19755 5072 19811 5079
rect 19675 5015 19731 5020
rect 19675 4964 19723 5015
rect 19723 4964 19731 5015
rect 19755 5015 19811 5020
rect 19755 4964 19762 5015
rect 19762 4964 19811 5015
rect 647 4347 703 4351
rect 729 4347 785 4351
rect 811 4347 867 4351
rect 647 4295 649 4347
rect 649 4295 701 4347
rect 701 4295 703 4347
rect 729 4295 777 4347
rect 777 4295 785 4347
rect 811 4295 852 4347
rect 852 4295 867 4347
rect 892 4295 948 4351
rect 647 4215 649 4267
rect 649 4215 701 4267
rect 701 4215 703 4267
rect 729 4215 777 4267
rect 777 4215 785 4267
rect 811 4215 852 4267
rect 852 4215 867 4267
rect 647 4211 703 4215
rect 729 4211 785 4215
rect 811 4211 867 4215
rect 892 4211 948 4267
rect 6021 4347 6077 4351
rect 6103 4347 6159 4351
rect 6184 4347 6240 4351
rect 6265 4347 6321 4351
rect 6346 4347 6402 4351
rect 6021 4295 6070 4347
rect 6070 4295 6077 4347
rect 6103 4295 6137 4347
rect 6137 4295 6152 4347
rect 6152 4295 6159 4347
rect 6184 4295 6204 4347
rect 6204 4295 6219 4347
rect 6219 4295 6240 4347
rect 6265 4295 6271 4347
rect 6271 4295 6286 4347
rect 6286 4295 6321 4347
rect 6346 4295 6353 4347
rect 6353 4295 6402 4347
rect 6021 4215 6070 4267
rect 6070 4215 6077 4267
rect 6103 4215 6137 4267
rect 6137 4215 6152 4267
rect 6152 4215 6159 4267
rect 6184 4215 6204 4267
rect 6204 4215 6219 4267
rect 6219 4215 6240 4267
rect 6265 4215 6271 4267
rect 6271 4215 6286 4267
rect 6286 4215 6321 4267
rect 6346 4215 6353 4267
rect 6353 4215 6402 4267
rect 6021 4211 6077 4215
rect 6103 4211 6159 4215
rect 6184 4211 6240 4215
rect 6265 4211 6321 4215
rect 6346 4211 6402 4215
rect 6952 4347 7008 4351
rect 7034 4347 7090 4351
rect 7115 4347 7171 4351
rect 7196 4347 7252 4351
rect 7277 4347 7333 4351
rect 6952 4295 7001 4347
rect 7001 4295 7008 4347
rect 7034 4295 7068 4347
rect 7068 4295 7083 4347
rect 7083 4295 7090 4347
rect 7115 4295 7135 4347
rect 7135 4295 7150 4347
rect 7150 4295 7171 4347
rect 7196 4295 7202 4347
rect 7202 4295 7217 4347
rect 7217 4295 7252 4347
rect 7277 4295 7284 4347
rect 7284 4295 7333 4347
rect 6952 4215 7001 4267
rect 7001 4215 7008 4267
rect 7034 4215 7068 4267
rect 7068 4215 7083 4267
rect 7083 4215 7090 4267
rect 7115 4215 7135 4267
rect 7135 4215 7150 4267
rect 7150 4215 7171 4267
rect 7196 4215 7202 4267
rect 7202 4215 7217 4267
rect 7217 4215 7252 4267
rect 7277 4215 7284 4267
rect 7284 4215 7333 4267
rect 6952 4211 7008 4215
rect 7034 4211 7090 4215
rect 7115 4211 7171 4215
rect 7196 4211 7252 4215
rect 7277 4211 7333 4215
rect 12505 4347 12561 4351
rect 12587 4347 12643 4351
rect 12668 4347 12724 4351
rect 12749 4347 12805 4351
rect 12830 4347 12886 4351
rect 12505 4295 12554 4347
rect 12554 4295 12561 4347
rect 12587 4295 12621 4347
rect 12621 4295 12636 4347
rect 12636 4295 12643 4347
rect 12668 4295 12688 4347
rect 12688 4295 12703 4347
rect 12703 4295 12724 4347
rect 12749 4295 12755 4347
rect 12755 4295 12770 4347
rect 12770 4295 12805 4347
rect 12830 4295 12837 4347
rect 12837 4295 12886 4347
rect 12505 4215 12554 4267
rect 12554 4215 12561 4267
rect 12587 4215 12621 4267
rect 12621 4215 12636 4267
rect 12636 4215 12643 4267
rect 12668 4215 12688 4267
rect 12688 4215 12703 4267
rect 12703 4215 12724 4267
rect 12749 4215 12755 4267
rect 12755 4215 12770 4267
rect 12770 4215 12805 4267
rect 12830 4215 12837 4267
rect 12837 4215 12886 4267
rect 12505 4211 12561 4215
rect 12587 4211 12643 4215
rect 12668 4211 12724 4215
rect 12749 4211 12805 4215
rect 12830 4211 12886 4215
rect 13436 4347 13492 4351
rect 13518 4347 13574 4351
rect 13599 4347 13655 4351
rect 13680 4347 13736 4351
rect 13761 4347 13817 4351
rect 13436 4295 13485 4347
rect 13485 4295 13492 4347
rect 13518 4295 13552 4347
rect 13552 4295 13567 4347
rect 13567 4295 13574 4347
rect 13599 4295 13619 4347
rect 13619 4295 13634 4347
rect 13634 4295 13655 4347
rect 13680 4295 13686 4347
rect 13686 4295 13701 4347
rect 13701 4295 13736 4347
rect 13761 4295 13768 4347
rect 13768 4295 13817 4347
rect 13436 4215 13485 4267
rect 13485 4215 13492 4267
rect 13518 4215 13552 4267
rect 13552 4215 13567 4267
rect 13567 4215 13574 4267
rect 13599 4215 13619 4267
rect 13619 4215 13634 4267
rect 13634 4215 13655 4267
rect 13680 4215 13686 4267
rect 13686 4215 13701 4267
rect 13701 4215 13736 4267
rect 13761 4215 13768 4267
rect 13768 4215 13817 4267
rect 13436 4211 13492 4215
rect 13518 4211 13574 4215
rect 13599 4211 13655 4215
rect 13680 4211 13736 4215
rect 13761 4211 13817 4215
rect 19070 4347 19126 4351
rect 19070 4295 19119 4347
rect 19119 4295 19126 4347
rect 19152 4347 19208 4351
rect 19152 4295 19204 4347
rect 19204 4295 19208 4347
rect 19233 4347 19289 4351
rect 19233 4295 19237 4347
rect 19237 4295 19289 4347
rect 19314 4347 19370 4351
rect 19314 4295 19321 4347
rect 19321 4295 19370 4347
rect 19070 4215 19119 4267
rect 19119 4215 19126 4267
rect 19070 4211 19126 4215
rect 19152 4215 19204 4267
rect 19204 4215 19208 4267
rect 19152 4211 19208 4215
rect 19233 4215 19237 4267
rect 19237 4215 19289 4267
rect 19233 4211 19289 4215
rect 19314 4215 19321 4267
rect 19321 4215 19370 4267
rect 19314 4211 19370 4215
rect 647 2959 703 2963
rect 647 2907 696 2959
rect 696 2907 703 2959
rect 728 2959 784 2963
rect 728 2907 780 2959
rect 780 2907 784 2959
rect 808 2959 864 2963
rect 808 2907 812 2959
rect 812 2907 864 2959
rect 888 2959 944 2963
rect 888 2907 895 2959
rect 895 2907 944 2959
rect 647 2827 696 2879
rect 696 2827 703 2879
rect 647 2823 703 2827
rect 728 2827 780 2879
rect 780 2827 784 2879
rect 728 2823 784 2827
rect 808 2827 812 2879
rect 812 2827 864 2879
rect 808 2823 864 2827
rect 888 2827 895 2879
rect 895 2827 944 2879
rect 888 2823 944 2827
rect 6021 2959 6077 2963
rect 6103 2959 6159 2963
rect 6184 2959 6240 2963
rect 6265 2959 6321 2963
rect 6346 2959 6402 2963
rect 6021 2907 6070 2959
rect 6070 2907 6077 2959
rect 6103 2907 6137 2959
rect 6137 2907 6152 2959
rect 6152 2907 6159 2959
rect 6184 2907 6204 2959
rect 6204 2907 6219 2959
rect 6219 2907 6240 2959
rect 6265 2907 6271 2959
rect 6271 2907 6286 2959
rect 6286 2907 6321 2959
rect 6346 2907 6353 2959
rect 6353 2907 6402 2959
rect 6021 2827 6070 2879
rect 6070 2827 6077 2879
rect 6103 2827 6137 2879
rect 6137 2827 6152 2879
rect 6152 2827 6159 2879
rect 6184 2827 6204 2879
rect 6204 2827 6219 2879
rect 6219 2827 6240 2879
rect 6265 2827 6271 2879
rect 6271 2827 6286 2879
rect 6286 2827 6321 2879
rect 6346 2827 6353 2879
rect 6353 2827 6402 2879
rect 6021 2823 6077 2827
rect 6103 2823 6159 2827
rect 6184 2823 6240 2827
rect 6265 2823 6321 2827
rect 6346 2823 6402 2827
rect 6952 2959 7008 2963
rect 7034 2959 7090 2963
rect 7115 2959 7171 2963
rect 7196 2959 7252 2963
rect 7277 2959 7333 2963
rect 6952 2907 7001 2959
rect 7001 2907 7008 2959
rect 7034 2907 7068 2959
rect 7068 2907 7083 2959
rect 7083 2907 7090 2959
rect 7115 2907 7135 2959
rect 7135 2907 7150 2959
rect 7150 2907 7171 2959
rect 7196 2907 7202 2959
rect 7202 2907 7217 2959
rect 7217 2907 7252 2959
rect 7277 2907 7284 2959
rect 7284 2907 7333 2959
rect 6952 2827 7001 2879
rect 7001 2827 7008 2879
rect 7034 2827 7068 2879
rect 7068 2827 7083 2879
rect 7083 2827 7090 2879
rect 7115 2827 7135 2879
rect 7135 2827 7150 2879
rect 7150 2827 7171 2879
rect 7196 2827 7202 2879
rect 7202 2827 7217 2879
rect 7217 2827 7252 2879
rect 7277 2827 7284 2879
rect 7284 2827 7333 2879
rect 6952 2823 7008 2827
rect 7034 2823 7090 2827
rect 7115 2823 7171 2827
rect 7196 2823 7252 2827
rect 7277 2823 7333 2827
rect 12505 2959 12561 2963
rect 12587 2959 12643 2963
rect 12668 2959 12724 2963
rect 12749 2959 12805 2963
rect 12830 2959 12886 2963
rect 12505 2907 12554 2959
rect 12554 2907 12561 2959
rect 12587 2907 12621 2959
rect 12621 2907 12636 2959
rect 12636 2907 12643 2959
rect 12668 2907 12688 2959
rect 12688 2907 12703 2959
rect 12703 2907 12724 2959
rect 12749 2907 12755 2959
rect 12755 2907 12770 2959
rect 12770 2907 12805 2959
rect 12830 2907 12837 2959
rect 12837 2907 12886 2959
rect 12505 2827 12554 2879
rect 12554 2827 12561 2879
rect 12587 2827 12621 2879
rect 12621 2827 12636 2879
rect 12636 2827 12643 2879
rect 12668 2827 12688 2879
rect 12688 2827 12703 2879
rect 12703 2827 12724 2879
rect 12749 2827 12755 2879
rect 12755 2827 12770 2879
rect 12770 2827 12805 2879
rect 12830 2827 12837 2879
rect 12837 2827 12886 2879
rect 12505 2823 12561 2827
rect 12587 2823 12643 2827
rect 12668 2823 12724 2827
rect 12749 2823 12805 2827
rect 12830 2823 12886 2827
rect 13436 2959 13492 2963
rect 13518 2959 13574 2963
rect 13599 2959 13655 2963
rect 13680 2959 13736 2963
rect 13761 2959 13817 2963
rect 13436 2907 13485 2959
rect 13485 2907 13492 2959
rect 13518 2907 13552 2959
rect 13552 2907 13567 2959
rect 13567 2907 13574 2959
rect 13599 2907 13619 2959
rect 13619 2907 13634 2959
rect 13634 2907 13655 2959
rect 13680 2907 13686 2959
rect 13686 2907 13701 2959
rect 13701 2907 13736 2959
rect 13761 2907 13768 2959
rect 13768 2907 13817 2959
rect 13436 2827 13485 2879
rect 13485 2827 13492 2879
rect 13518 2827 13552 2879
rect 13552 2827 13567 2879
rect 13567 2827 13574 2879
rect 13599 2827 13619 2879
rect 13619 2827 13634 2879
rect 13634 2827 13655 2879
rect 13680 2827 13686 2879
rect 13686 2827 13701 2879
rect 13701 2827 13736 2879
rect 13761 2827 13768 2879
rect 13768 2827 13817 2879
rect 13436 2823 13492 2827
rect 13518 2823 13574 2827
rect 13599 2823 13655 2827
rect 13680 2823 13736 2827
rect 13761 2823 13817 2827
rect 19074 2959 19130 2963
rect 19074 2907 19123 2959
rect 19123 2907 19130 2959
rect 19154 2959 19210 2963
rect 19154 2907 19155 2959
rect 19155 2907 19207 2959
rect 19207 2907 19210 2959
rect 19234 2959 19290 2963
rect 19234 2907 19238 2959
rect 19238 2907 19290 2959
rect 19314 2959 19370 2963
rect 19314 2907 19321 2959
rect 19321 2907 19370 2959
rect 19074 2827 19123 2879
rect 19123 2827 19130 2879
rect 19074 2823 19130 2827
rect 19154 2827 19155 2879
rect 19155 2827 19207 2879
rect 19207 2827 19210 2879
rect 19154 2823 19210 2827
rect 19234 2827 19238 2879
rect 19238 2827 19290 2879
rect 19234 2823 19290 2827
rect 19314 2827 19321 2879
rect 19321 2827 19370 2879
rect 19314 2823 19370 2827
rect 647 2686 696 2738
rect 696 2686 703 2738
rect 647 2682 703 2686
rect 728 2686 780 2738
rect 780 2686 784 2738
rect 728 2682 784 2686
rect 808 2686 812 2738
rect 812 2686 864 2738
rect 808 2682 864 2686
rect 888 2686 895 2738
rect 895 2686 944 2738
rect 888 2682 944 2686
rect 647 2610 703 2614
rect 647 2558 696 2610
rect 696 2558 703 2610
rect 728 2610 784 2614
rect 728 2558 780 2610
rect 780 2558 784 2610
rect 808 2610 864 2614
rect 808 2558 812 2610
rect 812 2558 864 2610
rect 888 2610 944 2614
rect 888 2558 895 2610
rect 895 2558 944 2610
rect 6021 2686 6070 2738
rect 6070 2686 6077 2738
rect 6102 2686 6137 2738
rect 6137 2686 6152 2738
rect 6152 2686 6158 2738
rect 6183 2686 6204 2738
rect 6204 2686 6219 2738
rect 6219 2686 6239 2738
rect 6264 2686 6271 2738
rect 6271 2686 6286 2738
rect 6286 2686 6320 2738
rect 6346 2686 6353 2738
rect 6353 2686 6402 2738
rect 6021 2682 6077 2686
rect 6102 2682 6158 2686
rect 6183 2682 6239 2686
rect 6264 2682 6320 2686
rect 6346 2682 6402 2686
rect 6021 2610 6077 2614
rect 6102 2610 6158 2614
rect 6183 2610 6239 2614
rect 6264 2610 6320 2614
rect 6346 2610 6402 2614
rect 6021 2558 6070 2610
rect 6070 2558 6077 2610
rect 6102 2558 6137 2610
rect 6137 2558 6152 2610
rect 6152 2558 6158 2610
rect 6183 2558 6204 2610
rect 6204 2558 6219 2610
rect 6219 2558 6239 2610
rect 6264 2558 6271 2610
rect 6271 2558 6286 2610
rect 6286 2558 6320 2610
rect 6346 2558 6353 2610
rect 6353 2558 6402 2610
rect 6952 2686 7001 2738
rect 7001 2686 7008 2738
rect 7034 2686 7068 2738
rect 7068 2686 7083 2738
rect 7083 2686 7090 2738
rect 7115 2686 7135 2738
rect 7135 2686 7150 2738
rect 7150 2686 7171 2738
rect 7196 2686 7202 2738
rect 7202 2686 7217 2738
rect 7217 2686 7252 2738
rect 7277 2686 7284 2738
rect 7284 2686 7333 2738
rect 6952 2682 7008 2686
rect 7034 2682 7090 2686
rect 7115 2682 7171 2686
rect 7196 2682 7252 2686
rect 7277 2682 7333 2686
rect 6952 2610 7008 2614
rect 7034 2610 7090 2614
rect 7115 2610 7171 2614
rect 7196 2610 7252 2614
rect 7277 2610 7333 2614
rect 6952 2558 7001 2610
rect 7001 2558 7008 2610
rect 7034 2558 7068 2610
rect 7068 2558 7083 2610
rect 7083 2558 7090 2610
rect 7115 2558 7135 2610
rect 7135 2558 7150 2610
rect 7150 2558 7171 2610
rect 7196 2558 7202 2610
rect 7202 2558 7217 2610
rect 7217 2558 7252 2610
rect 7277 2558 7284 2610
rect 7284 2558 7333 2610
rect 12505 2686 12554 2738
rect 12554 2686 12561 2738
rect 12586 2686 12621 2738
rect 12621 2686 12636 2738
rect 12636 2686 12642 2738
rect 12667 2686 12688 2738
rect 12688 2686 12703 2738
rect 12703 2686 12723 2738
rect 12748 2686 12755 2738
rect 12755 2686 12770 2738
rect 12770 2686 12804 2738
rect 12830 2686 12837 2738
rect 12837 2686 12886 2738
rect 12505 2682 12561 2686
rect 12586 2682 12642 2686
rect 12667 2682 12723 2686
rect 12748 2682 12804 2686
rect 12830 2682 12886 2686
rect 12505 2610 12561 2614
rect 12586 2610 12642 2614
rect 12667 2610 12723 2614
rect 12748 2610 12804 2614
rect 12830 2610 12886 2614
rect 12505 2558 12554 2610
rect 12554 2558 12561 2610
rect 12586 2558 12621 2610
rect 12621 2558 12636 2610
rect 12636 2558 12642 2610
rect 12667 2558 12688 2610
rect 12688 2558 12703 2610
rect 12703 2558 12723 2610
rect 12748 2558 12755 2610
rect 12755 2558 12770 2610
rect 12770 2558 12804 2610
rect 12830 2558 12837 2610
rect 12837 2558 12886 2610
rect 13436 2686 13485 2738
rect 13485 2686 13492 2738
rect 13518 2686 13552 2738
rect 13552 2686 13567 2738
rect 13567 2686 13574 2738
rect 13599 2686 13619 2738
rect 13619 2686 13634 2738
rect 13634 2686 13655 2738
rect 13680 2686 13686 2738
rect 13686 2686 13701 2738
rect 13701 2686 13736 2738
rect 13761 2686 13768 2738
rect 13768 2686 13817 2738
rect 13436 2682 13492 2686
rect 13518 2682 13574 2686
rect 13599 2682 13655 2686
rect 13680 2682 13736 2686
rect 13761 2682 13817 2686
rect 13436 2610 13492 2614
rect 13518 2610 13574 2614
rect 13599 2610 13655 2614
rect 13680 2610 13736 2614
rect 13761 2610 13817 2614
rect 13436 2558 13485 2610
rect 13485 2558 13492 2610
rect 13518 2558 13552 2610
rect 13552 2558 13567 2610
rect 13567 2558 13574 2610
rect 13599 2558 13619 2610
rect 13619 2558 13634 2610
rect 13634 2558 13655 2610
rect 13680 2558 13686 2610
rect 13686 2558 13701 2610
rect 13701 2558 13736 2610
rect 13761 2558 13768 2610
rect 13768 2558 13817 2610
rect 19074 2686 19123 2738
rect 19123 2686 19130 2738
rect 19074 2682 19130 2686
rect 19154 2686 19206 2738
rect 19206 2686 19210 2738
rect 19154 2682 19210 2686
rect 19234 2686 19237 2738
rect 19237 2686 19289 2738
rect 19289 2686 19290 2738
rect 19234 2682 19290 2686
rect 19314 2686 19321 2738
rect 19321 2686 19370 2738
rect 19314 2682 19370 2686
rect 19074 2610 19130 2614
rect 19074 2558 19123 2610
rect 19123 2558 19130 2610
rect 19154 2610 19210 2614
rect 19154 2558 19206 2610
rect 19206 2558 19210 2610
rect 19234 2610 19290 2614
rect 19234 2558 19237 2610
rect 19237 2558 19289 2610
rect 19289 2558 19290 2610
rect 19314 2610 19370 2614
rect 19314 2558 19321 2610
rect 19321 2558 19370 2610
rect 1038 2385 1079 2437
rect 1079 2385 1092 2437
rect 1092 2385 1094 2437
rect 1120 2385 1144 2437
rect 1144 2385 1157 2437
rect 1157 2385 1176 2437
rect 1202 2385 1209 2437
rect 1209 2385 1222 2437
rect 1222 2385 1258 2437
rect 1284 2385 1286 2437
rect 1286 2385 1338 2437
rect 1338 2385 1340 2437
rect 1366 2385 1402 2437
rect 1402 2385 1414 2437
rect 1414 2385 1422 2437
rect 1448 2385 1466 2437
rect 1466 2385 1478 2437
rect 1478 2385 1504 2437
rect 1530 2385 1542 2437
rect 1542 2385 1586 2437
rect 1611 2385 1658 2437
rect 1658 2385 1667 2437
rect 1692 2385 1722 2437
rect 1722 2385 1734 2437
rect 1734 2385 1748 2437
rect 1773 2385 1786 2437
rect 1786 2385 1798 2437
rect 1798 2385 1829 2437
rect 1854 2385 1862 2437
rect 1862 2385 1910 2437
rect 1038 2381 1094 2385
rect 1120 2381 1176 2385
rect 1202 2381 1258 2385
rect 1284 2381 1340 2385
rect 1366 2381 1422 2385
rect 1448 2381 1504 2385
rect 1530 2381 1586 2385
rect 1611 2381 1667 2385
rect 1692 2381 1748 2385
rect 1773 2381 1829 2385
rect 1854 2381 1910 2385
rect 1038 2317 1079 2353
rect 1079 2317 1092 2353
rect 1092 2317 1094 2353
rect 1120 2317 1144 2353
rect 1144 2317 1157 2353
rect 1157 2317 1176 2353
rect 1202 2317 1209 2353
rect 1209 2317 1222 2353
rect 1222 2317 1258 2353
rect 1284 2317 1286 2353
rect 1286 2317 1338 2353
rect 1338 2317 1340 2353
rect 1366 2317 1402 2353
rect 1402 2317 1414 2353
rect 1414 2317 1422 2353
rect 1448 2317 1466 2353
rect 1466 2317 1478 2353
rect 1478 2317 1504 2353
rect 1530 2317 1542 2353
rect 1542 2317 1586 2353
rect 1611 2317 1658 2353
rect 1658 2317 1667 2353
rect 1692 2317 1722 2353
rect 1722 2317 1734 2353
rect 1734 2317 1748 2353
rect 1773 2317 1786 2353
rect 1786 2317 1798 2353
rect 1798 2317 1829 2353
rect 1854 2317 1862 2353
rect 1862 2317 1910 2353
rect 1038 2301 1094 2317
rect 1120 2301 1176 2317
rect 1202 2301 1258 2317
rect 1284 2301 1340 2317
rect 1366 2301 1422 2317
rect 1448 2301 1504 2317
rect 1530 2301 1586 2317
rect 1611 2301 1667 2317
rect 1692 2301 1748 2317
rect 1773 2301 1829 2317
rect 1854 2301 1910 2317
rect 1038 2297 1079 2301
rect 1079 2297 1092 2301
rect 1092 2297 1094 2301
rect 1120 2297 1144 2301
rect 1144 2297 1157 2301
rect 1157 2297 1176 2301
rect 1202 2297 1209 2301
rect 1209 2297 1222 2301
rect 1222 2297 1258 2301
rect 1284 2297 1286 2301
rect 1286 2297 1338 2301
rect 1338 2297 1340 2301
rect 1366 2297 1402 2301
rect 1402 2297 1414 2301
rect 1414 2297 1422 2301
rect 1448 2297 1466 2301
rect 1466 2297 1478 2301
rect 1478 2297 1504 2301
rect 1530 2297 1542 2301
rect 1542 2297 1586 2301
rect 1038 2249 1079 2269
rect 1079 2249 1092 2269
rect 1092 2249 1094 2269
rect 1120 2249 1144 2269
rect 1144 2249 1157 2269
rect 1157 2249 1176 2269
rect 1202 2249 1209 2269
rect 1209 2249 1222 2269
rect 1222 2249 1258 2269
rect 1284 2249 1286 2269
rect 1286 2249 1338 2269
rect 1338 2249 1340 2269
rect 1366 2249 1402 2269
rect 1402 2249 1414 2269
rect 1414 2249 1422 2269
rect 1448 2249 1466 2269
rect 1466 2249 1478 2269
rect 1478 2249 1504 2269
rect 1530 2249 1542 2269
rect 1542 2249 1586 2269
rect 1611 2297 1658 2301
rect 1658 2297 1667 2301
rect 1692 2297 1722 2301
rect 1722 2297 1734 2301
rect 1734 2297 1748 2301
rect 1773 2297 1786 2301
rect 1786 2297 1798 2301
rect 1798 2297 1829 2301
rect 1854 2297 1862 2301
rect 1862 2297 1910 2301
rect 1611 2249 1658 2269
rect 1658 2249 1667 2269
rect 1692 2249 1722 2269
rect 1722 2249 1734 2269
rect 1734 2249 1748 2269
rect 1773 2249 1786 2269
rect 1786 2249 1798 2269
rect 1798 2249 1829 2269
rect 1854 2249 1862 2269
rect 1862 2249 1910 2269
rect 1038 2233 1094 2249
rect 1120 2233 1176 2249
rect 1202 2233 1258 2249
rect 1284 2233 1340 2249
rect 1366 2233 1422 2249
rect 1448 2233 1504 2249
rect 1530 2233 1586 2249
rect 1611 2233 1667 2249
rect 1692 2233 1748 2249
rect 1773 2233 1829 2249
rect 1854 2233 1910 2249
rect 1038 2213 1079 2233
rect 1079 2213 1092 2233
rect 1092 2213 1094 2233
rect 1120 2213 1144 2233
rect 1144 2213 1157 2233
rect 1157 2213 1176 2233
rect 1202 2213 1209 2233
rect 1209 2213 1222 2233
rect 1222 2213 1258 2233
rect 1284 2213 1286 2233
rect 1286 2213 1338 2233
rect 1338 2213 1340 2233
rect 1366 2213 1402 2233
rect 1402 2213 1414 2233
rect 1414 2213 1422 2233
rect 1448 2213 1466 2233
rect 1466 2213 1478 2233
rect 1478 2213 1504 2233
rect 1530 2213 1542 2233
rect 1542 2213 1586 2233
rect 1038 2181 1079 2185
rect 1079 2181 1092 2185
rect 1092 2181 1094 2185
rect 1120 2181 1144 2185
rect 1144 2181 1157 2185
rect 1157 2181 1176 2185
rect 1202 2181 1209 2185
rect 1209 2181 1222 2185
rect 1222 2181 1258 2185
rect 1284 2181 1286 2185
rect 1286 2181 1338 2185
rect 1338 2181 1340 2185
rect 1366 2181 1402 2185
rect 1402 2181 1414 2185
rect 1414 2181 1422 2185
rect 1448 2181 1466 2185
rect 1466 2181 1478 2185
rect 1478 2181 1504 2185
rect 1530 2181 1542 2185
rect 1542 2181 1586 2185
rect 1611 2213 1658 2233
rect 1658 2213 1667 2233
rect 1692 2213 1722 2233
rect 1722 2213 1734 2233
rect 1734 2213 1748 2233
rect 1773 2213 1786 2233
rect 1786 2213 1798 2233
rect 1798 2213 1829 2233
rect 1854 2213 1862 2233
rect 1862 2213 1910 2233
rect 1611 2181 1658 2185
rect 1658 2181 1667 2185
rect 1692 2181 1722 2185
rect 1722 2181 1734 2185
rect 1734 2181 1748 2185
rect 1773 2181 1786 2185
rect 1786 2181 1798 2185
rect 1798 2181 1829 2185
rect 1854 2181 1862 2185
rect 1862 2181 1910 2185
rect 1038 2165 1094 2181
rect 1120 2165 1176 2181
rect 1202 2165 1258 2181
rect 1284 2165 1340 2181
rect 1366 2165 1422 2181
rect 1448 2165 1504 2181
rect 1530 2165 1586 2181
rect 1611 2165 1667 2181
rect 1692 2165 1748 2181
rect 1773 2165 1829 2181
rect 1854 2165 1910 2181
rect 1038 2129 1079 2165
rect 1079 2129 1092 2165
rect 1092 2129 1094 2165
rect 1120 2129 1144 2165
rect 1144 2129 1157 2165
rect 1157 2129 1176 2165
rect 1202 2129 1209 2165
rect 1209 2129 1222 2165
rect 1222 2129 1258 2165
rect 1284 2129 1286 2165
rect 1286 2129 1338 2165
rect 1338 2129 1340 2165
rect 1366 2129 1402 2165
rect 1402 2129 1414 2165
rect 1414 2129 1422 2165
rect 1448 2129 1466 2165
rect 1466 2129 1478 2165
rect 1478 2129 1504 2165
rect 1530 2129 1542 2165
rect 1542 2129 1586 2165
rect 1611 2129 1658 2165
rect 1658 2129 1667 2165
rect 1692 2129 1722 2165
rect 1722 2129 1734 2165
rect 1734 2129 1748 2165
rect 1773 2129 1786 2165
rect 1786 2129 1798 2165
rect 1798 2129 1829 2165
rect 1854 2129 1862 2165
rect 1862 2129 1910 2165
rect 1038 2097 1094 2101
rect 1120 2097 1176 2101
rect 1202 2097 1258 2101
rect 1284 2097 1340 2101
rect 1366 2097 1422 2101
rect 1448 2097 1504 2101
rect 1530 2097 1586 2101
rect 1611 2097 1667 2101
rect 1692 2097 1748 2101
rect 1773 2097 1829 2101
rect 1854 2097 1910 2101
rect 1038 2045 1079 2097
rect 1079 2045 1092 2097
rect 1092 2045 1094 2097
rect 1120 2045 1144 2097
rect 1144 2045 1157 2097
rect 1157 2045 1176 2097
rect 1202 2045 1209 2097
rect 1209 2045 1222 2097
rect 1222 2045 1258 2097
rect 1284 2045 1286 2097
rect 1286 2045 1338 2097
rect 1338 2045 1340 2097
rect 1366 2045 1402 2097
rect 1402 2045 1414 2097
rect 1414 2045 1422 2097
rect 1448 2045 1466 2097
rect 1466 2045 1478 2097
rect 1478 2045 1504 2097
rect 1530 2045 1542 2097
rect 1542 2045 1586 2097
rect 1611 2045 1658 2097
rect 1658 2045 1667 2097
rect 1692 2045 1722 2097
rect 1722 2045 1734 2097
rect 1734 2045 1748 2097
rect 1773 2045 1786 2097
rect 1786 2045 1798 2097
rect 1798 2045 1829 2097
rect 1854 2045 1862 2097
rect 1862 2045 1910 2097
rect 5203 2381 5259 2437
rect 5284 2381 5340 2437
rect 5366 2381 5422 2437
rect 5448 2381 5504 2437
rect 5530 2381 5586 2437
rect 5612 2381 5668 2437
rect 5694 2381 5750 2437
rect 5776 2381 5832 2437
rect 5203 2297 5259 2353
rect 5284 2297 5340 2353
rect 5366 2297 5422 2353
rect 5448 2297 5504 2353
rect 5530 2297 5586 2353
rect 5612 2297 5668 2353
rect 5694 2297 5750 2353
rect 5776 2297 5832 2353
rect 5203 2213 5259 2269
rect 5284 2213 5340 2269
rect 5366 2213 5422 2269
rect 5448 2213 5504 2269
rect 5530 2213 5586 2269
rect 5612 2213 5668 2269
rect 5694 2213 5750 2269
rect 5776 2213 5832 2269
rect 5203 2129 5259 2185
rect 5284 2129 5340 2185
rect 5366 2129 5422 2185
rect 5448 2129 5504 2185
rect 5530 2129 5586 2185
rect 5612 2129 5668 2185
rect 5694 2129 5750 2185
rect 5776 2129 5832 2185
rect 5203 2045 5259 2101
rect 5284 2045 5340 2101
rect 5366 2045 5422 2101
rect 5448 2045 5504 2101
rect 5530 2045 5586 2101
rect 5612 2045 5668 2101
rect 5694 2045 5750 2101
rect 5776 2045 5832 2101
rect 7522 2385 7563 2437
rect 7563 2385 7576 2437
rect 7576 2385 7578 2437
rect 7604 2385 7628 2437
rect 7628 2385 7641 2437
rect 7641 2385 7660 2437
rect 7686 2385 7693 2437
rect 7693 2385 7706 2437
rect 7706 2385 7742 2437
rect 7768 2385 7770 2437
rect 7770 2385 7822 2437
rect 7822 2385 7824 2437
rect 7850 2385 7886 2437
rect 7886 2385 7898 2437
rect 7898 2385 7906 2437
rect 7932 2385 7950 2437
rect 7950 2385 7962 2437
rect 7962 2385 7988 2437
rect 8014 2385 8026 2437
rect 8026 2385 8070 2437
rect 8095 2385 8142 2437
rect 8142 2385 8151 2437
rect 8176 2385 8206 2437
rect 8206 2385 8218 2437
rect 8218 2385 8232 2437
rect 8257 2385 8270 2437
rect 8270 2385 8282 2437
rect 8282 2385 8313 2437
rect 8338 2385 8346 2437
rect 8346 2385 8394 2437
rect 7522 2381 7578 2385
rect 7604 2381 7660 2385
rect 7686 2381 7742 2385
rect 7768 2381 7824 2385
rect 7850 2381 7906 2385
rect 7932 2381 7988 2385
rect 8014 2381 8070 2385
rect 8095 2381 8151 2385
rect 8176 2381 8232 2385
rect 8257 2381 8313 2385
rect 8338 2381 8394 2385
rect 7522 2317 7563 2353
rect 7563 2317 7576 2353
rect 7576 2317 7578 2353
rect 7604 2317 7628 2353
rect 7628 2317 7641 2353
rect 7641 2317 7660 2353
rect 7686 2317 7693 2353
rect 7693 2317 7706 2353
rect 7706 2317 7742 2353
rect 7768 2317 7770 2353
rect 7770 2317 7822 2353
rect 7822 2317 7824 2353
rect 7850 2317 7886 2353
rect 7886 2317 7898 2353
rect 7898 2317 7906 2353
rect 7932 2317 7950 2353
rect 7950 2317 7962 2353
rect 7962 2317 7988 2353
rect 8014 2317 8026 2353
rect 8026 2317 8070 2353
rect 8095 2317 8142 2353
rect 8142 2317 8151 2353
rect 8176 2317 8206 2353
rect 8206 2317 8218 2353
rect 8218 2317 8232 2353
rect 8257 2317 8270 2353
rect 8270 2317 8282 2353
rect 8282 2317 8313 2353
rect 8338 2317 8346 2353
rect 8346 2317 8394 2353
rect 7522 2301 7578 2317
rect 7604 2301 7660 2317
rect 7686 2301 7742 2317
rect 7768 2301 7824 2317
rect 7850 2301 7906 2317
rect 7932 2301 7988 2317
rect 8014 2301 8070 2317
rect 8095 2301 8151 2317
rect 8176 2301 8232 2317
rect 8257 2301 8313 2317
rect 8338 2301 8394 2317
rect 7522 2297 7563 2301
rect 7563 2297 7576 2301
rect 7576 2297 7578 2301
rect 7604 2297 7628 2301
rect 7628 2297 7641 2301
rect 7641 2297 7660 2301
rect 7686 2297 7693 2301
rect 7693 2297 7706 2301
rect 7706 2297 7742 2301
rect 7768 2297 7770 2301
rect 7770 2297 7822 2301
rect 7822 2297 7824 2301
rect 7850 2297 7886 2301
rect 7886 2297 7898 2301
rect 7898 2297 7906 2301
rect 7932 2297 7950 2301
rect 7950 2297 7962 2301
rect 7962 2297 7988 2301
rect 8014 2297 8026 2301
rect 8026 2297 8070 2301
rect 7522 2249 7563 2269
rect 7563 2249 7576 2269
rect 7576 2249 7578 2269
rect 7604 2249 7628 2269
rect 7628 2249 7641 2269
rect 7641 2249 7660 2269
rect 7686 2249 7693 2269
rect 7693 2249 7706 2269
rect 7706 2249 7742 2269
rect 7768 2249 7770 2269
rect 7770 2249 7822 2269
rect 7822 2249 7824 2269
rect 7850 2249 7886 2269
rect 7886 2249 7898 2269
rect 7898 2249 7906 2269
rect 7932 2249 7950 2269
rect 7950 2249 7962 2269
rect 7962 2249 7988 2269
rect 8014 2249 8026 2269
rect 8026 2249 8070 2269
rect 8095 2297 8142 2301
rect 8142 2297 8151 2301
rect 8176 2297 8206 2301
rect 8206 2297 8218 2301
rect 8218 2297 8232 2301
rect 8257 2297 8270 2301
rect 8270 2297 8282 2301
rect 8282 2297 8313 2301
rect 8338 2297 8346 2301
rect 8346 2297 8394 2301
rect 8095 2249 8142 2269
rect 8142 2249 8151 2269
rect 8176 2249 8206 2269
rect 8206 2249 8218 2269
rect 8218 2249 8232 2269
rect 8257 2249 8270 2269
rect 8270 2249 8282 2269
rect 8282 2249 8313 2269
rect 8338 2249 8346 2269
rect 8346 2249 8394 2269
rect 7522 2233 7578 2249
rect 7604 2233 7660 2249
rect 7686 2233 7742 2249
rect 7768 2233 7824 2249
rect 7850 2233 7906 2249
rect 7932 2233 7988 2249
rect 8014 2233 8070 2249
rect 8095 2233 8151 2249
rect 8176 2233 8232 2249
rect 8257 2233 8313 2249
rect 8338 2233 8394 2249
rect 7522 2213 7563 2233
rect 7563 2213 7576 2233
rect 7576 2213 7578 2233
rect 7604 2213 7628 2233
rect 7628 2213 7641 2233
rect 7641 2213 7660 2233
rect 7686 2213 7693 2233
rect 7693 2213 7706 2233
rect 7706 2213 7742 2233
rect 7768 2213 7770 2233
rect 7770 2213 7822 2233
rect 7822 2213 7824 2233
rect 7850 2213 7886 2233
rect 7886 2213 7898 2233
rect 7898 2213 7906 2233
rect 7932 2213 7950 2233
rect 7950 2213 7962 2233
rect 7962 2213 7988 2233
rect 8014 2213 8026 2233
rect 8026 2213 8070 2233
rect 7522 2181 7563 2185
rect 7563 2181 7576 2185
rect 7576 2181 7578 2185
rect 7604 2181 7628 2185
rect 7628 2181 7641 2185
rect 7641 2181 7660 2185
rect 7686 2181 7693 2185
rect 7693 2181 7706 2185
rect 7706 2181 7742 2185
rect 7768 2181 7770 2185
rect 7770 2181 7822 2185
rect 7822 2181 7824 2185
rect 7850 2181 7886 2185
rect 7886 2181 7898 2185
rect 7898 2181 7906 2185
rect 7932 2181 7950 2185
rect 7950 2181 7962 2185
rect 7962 2181 7988 2185
rect 8014 2181 8026 2185
rect 8026 2181 8070 2185
rect 8095 2213 8142 2233
rect 8142 2213 8151 2233
rect 8176 2213 8206 2233
rect 8206 2213 8218 2233
rect 8218 2213 8232 2233
rect 8257 2213 8270 2233
rect 8270 2213 8282 2233
rect 8282 2213 8313 2233
rect 8338 2213 8346 2233
rect 8346 2213 8394 2233
rect 8095 2181 8142 2185
rect 8142 2181 8151 2185
rect 8176 2181 8206 2185
rect 8206 2181 8218 2185
rect 8218 2181 8232 2185
rect 8257 2181 8270 2185
rect 8270 2181 8282 2185
rect 8282 2181 8313 2185
rect 8338 2181 8346 2185
rect 8346 2181 8394 2185
rect 7522 2165 7578 2181
rect 7604 2165 7660 2181
rect 7686 2165 7742 2181
rect 7768 2165 7824 2181
rect 7850 2165 7906 2181
rect 7932 2165 7988 2181
rect 8014 2165 8070 2181
rect 8095 2165 8151 2181
rect 8176 2165 8232 2181
rect 8257 2165 8313 2181
rect 8338 2165 8394 2181
rect 7522 2129 7563 2165
rect 7563 2129 7576 2165
rect 7576 2129 7578 2165
rect 7604 2129 7628 2165
rect 7628 2129 7641 2165
rect 7641 2129 7660 2165
rect 7686 2129 7693 2165
rect 7693 2129 7706 2165
rect 7706 2129 7742 2165
rect 7768 2129 7770 2165
rect 7770 2129 7822 2165
rect 7822 2129 7824 2165
rect 7850 2129 7886 2165
rect 7886 2129 7898 2165
rect 7898 2129 7906 2165
rect 7932 2129 7950 2165
rect 7950 2129 7962 2165
rect 7962 2129 7988 2165
rect 8014 2129 8026 2165
rect 8026 2129 8070 2165
rect 8095 2129 8142 2165
rect 8142 2129 8151 2165
rect 8176 2129 8206 2165
rect 8206 2129 8218 2165
rect 8218 2129 8232 2165
rect 8257 2129 8270 2165
rect 8270 2129 8282 2165
rect 8282 2129 8313 2165
rect 8338 2129 8346 2165
rect 8346 2129 8394 2165
rect 7522 2097 7578 2101
rect 7604 2097 7660 2101
rect 7686 2097 7742 2101
rect 7768 2097 7824 2101
rect 7850 2097 7906 2101
rect 7932 2097 7988 2101
rect 8014 2097 8070 2101
rect 8095 2097 8151 2101
rect 8176 2097 8232 2101
rect 8257 2097 8313 2101
rect 8338 2097 8394 2101
rect 7522 2045 7563 2097
rect 7563 2045 7576 2097
rect 7576 2045 7578 2097
rect 7604 2045 7628 2097
rect 7628 2045 7641 2097
rect 7641 2045 7660 2097
rect 7686 2045 7693 2097
rect 7693 2045 7706 2097
rect 7706 2045 7742 2097
rect 7768 2045 7770 2097
rect 7770 2045 7822 2097
rect 7822 2045 7824 2097
rect 7850 2045 7886 2097
rect 7886 2045 7898 2097
rect 7898 2045 7906 2097
rect 7932 2045 7950 2097
rect 7950 2045 7962 2097
rect 7962 2045 7988 2097
rect 8014 2045 8026 2097
rect 8026 2045 8070 2097
rect 8095 2045 8142 2097
rect 8142 2045 8151 2097
rect 8176 2045 8206 2097
rect 8206 2045 8218 2097
rect 8218 2045 8232 2097
rect 8257 2045 8270 2097
rect 8270 2045 8282 2097
rect 8282 2045 8313 2097
rect 8338 2045 8346 2097
rect 8346 2045 8394 2097
rect 11444 2385 11492 2437
rect 11492 2385 11500 2437
rect 11525 2385 11556 2437
rect 11556 2385 11568 2437
rect 11568 2385 11581 2437
rect 11606 2385 11620 2437
rect 11620 2385 11632 2437
rect 11632 2385 11662 2437
rect 11687 2385 11696 2437
rect 11696 2385 11743 2437
rect 11768 2385 11812 2437
rect 11812 2385 11824 2437
rect 11850 2385 11876 2437
rect 11876 2385 11888 2437
rect 11888 2385 11906 2437
rect 11932 2385 11940 2437
rect 11940 2385 11952 2437
rect 11952 2385 11988 2437
rect 12014 2385 12016 2437
rect 12016 2385 12068 2437
rect 12068 2385 12070 2437
rect 12096 2385 12132 2437
rect 12132 2385 12145 2437
rect 12145 2385 12152 2437
rect 12178 2385 12197 2437
rect 12197 2385 12210 2437
rect 12210 2385 12234 2437
rect 12260 2385 12262 2437
rect 12262 2385 12275 2437
rect 12275 2385 12316 2437
rect 11444 2381 11500 2385
rect 11525 2381 11581 2385
rect 11606 2381 11662 2385
rect 11687 2381 11743 2385
rect 11768 2381 11824 2385
rect 11850 2381 11906 2385
rect 11932 2381 11988 2385
rect 12014 2381 12070 2385
rect 12096 2381 12152 2385
rect 12178 2381 12234 2385
rect 12260 2381 12316 2385
rect 11444 2317 11492 2353
rect 11492 2317 11500 2353
rect 11525 2317 11556 2353
rect 11556 2317 11568 2353
rect 11568 2317 11581 2353
rect 11606 2317 11620 2353
rect 11620 2317 11632 2353
rect 11632 2317 11662 2353
rect 11687 2317 11696 2353
rect 11696 2317 11743 2353
rect 11768 2317 11812 2353
rect 11812 2317 11824 2353
rect 11850 2317 11876 2353
rect 11876 2317 11888 2353
rect 11888 2317 11906 2353
rect 11932 2317 11940 2353
rect 11940 2317 11952 2353
rect 11952 2317 11988 2353
rect 12014 2317 12016 2353
rect 12016 2317 12068 2353
rect 12068 2317 12070 2353
rect 12096 2317 12132 2353
rect 12132 2317 12145 2353
rect 12145 2317 12152 2353
rect 12178 2317 12197 2353
rect 12197 2317 12210 2353
rect 12210 2317 12234 2353
rect 12260 2317 12262 2353
rect 12262 2317 12275 2353
rect 12275 2317 12316 2353
rect 11444 2301 11500 2317
rect 11525 2301 11581 2317
rect 11606 2301 11662 2317
rect 11687 2301 11743 2317
rect 11768 2301 11824 2317
rect 11850 2301 11906 2317
rect 11932 2301 11988 2317
rect 12014 2301 12070 2317
rect 12096 2301 12152 2317
rect 12178 2301 12234 2317
rect 12260 2301 12316 2317
rect 11444 2297 11492 2301
rect 11492 2297 11500 2301
rect 11525 2297 11556 2301
rect 11556 2297 11568 2301
rect 11568 2297 11581 2301
rect 11606 2297 11620 2301
rect 11620 2297 11632 2301
rect 11632 2297 11662 2301
rect 11687 2297 11696 2301
rect 11696 2297 11743 2301
rect 11444 2249 11492 2269
rect 11492 2249 11500 2269
rect 11525 2249 11556 2269
rect 11556 2249 11568 2269
rect 11568 2249 11581 2269
rect 11606 2249 11620 2269
rect 11620 2249 11632 2269
rect 11632 2249 11662 2269
rect 11687 2249 11696 2269
rect 11696 2249 11743 2269
rect 11768 2297 11812 2301
rect 11812 2297 11824 2301
rect 11850 2297 11876 2301
rect 11876 2297 11888 2301
rect 11888 2297 11906 2301
rect 11932 2297 11940 2301
rect 11940 2297 11952 2301
rect 11952 2297 11988 2301
rect 12014 2297 12016 2301
rect 12016 2297 12068 2301
rect 12068 2297 12070 2301
rect 12096 2297 12132 2301
rect 12132 2297 12145 2301
rect 12145 2297 12152 2301
rect 12178 2297 12197 2301
rect 12197 2297 12210 2301
rect 12210 2297 12234 2301
rect 12260 2297 12262 2301
rect 12262 2297 12275 2301
rect 12275 2297 12316 2301
rect 11768 2249 11812 2269
rect 11812 2249 11824 2269
rect 11850 2249 11876 2269
rect 11876 2249 11888 2269
rect 11888 2249 11906 2269
rect 11932 2249 11940 2269
rect 11940 2249 11952 2269
rect 11952 2249 11988 2269
rect 12014 2249 12016 2269
rect 12016 2249 12068 2269
rect 12068 2249 12070 2269
rect 12096 2249 12132 2269
rect 12132 2249 12145 2269
rect 12145 2249 12152 2269
rect 12178 2249 12197 2269
rect 12197 2249 12210 2269
rect 12210 2249 12234 2269
rect 12260 2249 12262 2269
rect 12262 2249 12275 2269
rect 12275 2249 12316 2269
rect 11444 2233 11500 2249
rect 11525 2233 11581 2249
rect 11606 2233 11662 2249
rect 11687 2233 11743 2249
rect 11768 2233 11824 2249
rect 11850 2233 11906 2249
rect 11932 2233 11988 2249
rect 12014 2233 12070 2249
rect 12096 2233 12152 2249
rect 12178 2233 12234 2249
rect 12260 2233 12316 2249
rect 11444 2213 11492 2233
rect 11492 2213 11500 2233
rect 11525 2213 11556 2233
rect 11556 2213 11568 2233
rect 11568 2213 11581 2233
rect 11606 2213 11620 2233
rect 11620 2213 11632 2233
rect 11632 2213 11662 2233
rect 11687 2213 11696 2233
rect 11696 2213 11743 2233
rect 11444 2181 11492 2185
rect 11492 2181 11500 2185
rect 11525 2181 11556 2185
rect 11556 2181 11568 2185
rect 11568 2181 11581 2185
rect 11606 2181 11620 2185
rect 11620 2181 11632 2185
rect 11632 2181 11662 2185
rect 11687 2181 11696 2185
rect 11696 2181 11743 2185
rect 11768 2213 11812 2233
rect 11812 2213 11824 2233
rect 11850 2213 11876 2233
rect 11876 2213 11888 2233
rect 11888 2213 11906 2233
rect 11932 2213 11940 2233
rect 11940 2213 11952 2233
rect 11952 2213 11988 2233
rect 12014 2213 12016 2233
rect 12016 2213 12068 2233
rect 12068 2213 12070 2233
rect 12096 2213 12132 2233
rect 12132 2213 12145 2233
rect 12145 2213 12152 2233
rect 12178 2213 12197 2233
rect 12197 2213 12210 2233
rect 12210 2213 12234 2233
rect 12260 2213 12262 2233
rect 12262 2213 12275 2233
rect 12275 2213 12316 2233
rect 11768 2181 11812 2185
rect 11812 2181 11824 2185
rect 11850 2181 11876 2185
rect 11876 2181 11888 2185
rect 11888 2181 11906 2185
rect 11932 2181 11940 2185
rect 11940 2181 11952 2185
rect 11952 2181 11988 2185
rect 12014 2181 12016 2185
rect 12016 2181 12068 2185
rect 12068 2181 12070 2185
rect 12096 2181 12132 2185
rect 12132 2181 12145 2185
rect 12145 2181 12152 2185
rect 12178 2181 12197 2185
rect 12197 2181 12210 2185
rect 12210 2181 12234 2185
rect 12260 2181 12262 2185
rect 12262 2181 12275 2185
rect 12275 2181 12316 2185
rect 11444 2165 11500 2181
rect 11525 2165 11581 2181
rect 11606 2165 11662 2181
rect 11687 2165 11743 2181
rect 11768 2165 11824 2181
rect 11850 2165 11906 2181
rect 11932 2165 11988 2181
rect 12014 2165 12070 2181
rect 12096 2165 12152 2181
rect 12178 2165 12234 2181
rect 12260 2165 12316 2181
rect 11444 2129 11492 2165
rect 11492 2129 11500 2165
rect 11525 2129 11556 2165
rect 11556 2129 11568 2165
rect 11568 2129 11581 2165
rect 11606 2129 11620 2165
rect 11620 2129 11632 2165
rect 11632 2129 11662 2165
rect 11687 2129 11696 2165
rect 11696 2129 11743 2165
rect 11768 2129 11812 2165
rect 11812 2129 11824 2165
rect 11850 2129 11876 2165
rect 11876 2129 11888 2165
rect 11888 2129 11906 2165
rect 11932 2129 11940 2165
rect 11940 2129 11952 2165
rect 11952 2129 11988 2165
rect 12014 2129 12016 2165
rect 12016 2129 12068 2165
rect 12068 2129 12070 2165
rect 12096 2129 12132 2165
rect 12132 2129 12145 2165
rect 12145 2129 12152 2165
rect 12178 2129 12197 2165
rect 12197 2129 12210 2165
rect 12210 2129 12234 2165
rect 12260 2129 12262 2165
rect 12262 2129 12275 2165
rect 12275 2129 12316 2165
rect 11444 2097 11500 2101
rect 11525 2097 11581 2101
rect 11606 2097 11662 2101
rect 11687 2097 11743 2101
rect 11768 2097 11824 2101
rect 11850 2097 11906 2101
rect 11932 2097 11988 2101
rect 12014 2097 12070 2101
rect 12096 2097 12152 2101
rect 12178 2097 12234 2101
rect 12260 2097 12316 2101
rect 11444 2045 11492 2097
rect 11492 2045 11500 2097
rect 11525 2045 11556 2097
rect 11556 2045 11568 2097
rect 11568 2045 11581 2097
rect 11606 2045 11620 2097
rect 11620 2045 11632 2097
rect 11632 2045 11662 2097
rect 11687 2045 11696 2097
rect 11696 2045 11743 2097
rect 11768 2045 11812 2097
rect 11812 2045 11824 2097
rect 11850 2045 11876 2097
rect 11876 2045 11888 2097
rect 11888 2045 11906 2097
rect 11932 2045 11940 2097
rect 11940 2045 11952 2097
rect 11952 2045 11988 2097
rect 12014 2045 12016 2097
rect 12016 2045 12068 2097
rect 12068 2045 12070 2097
rect 12096 2045 12132 2097
rect 12132 2045 12145 2097
rect 12145 2045 12152 2097
rect 12178 2045 12197 2097
rect 12197 2045 12210 2097
rect 12210 2045 12234 2097
rect 12260 2045 12262 2097
rect 12262 2045 12275 2097
rect 12275 2045 12316 2097
rect 14006 2385 14047 2437
rect 14047 2385 14060 2437
rect 14060 2385 14062 2437
rect 14088 2385 14112 2437
rect 14112 2385 14125 2437
rect 14125 2385 14144 2437
rect 14170 2385 14177 2437
rect 14177 2385 14190 2437
rect 14190 2385 14226 2437
rect 14252 2385 14254 2437
rect 14254 2385 14306 2437
rect 14306 2385 14308 2437
rect 14334 2385 14370 2437
rect 14370 2385 14382 2437
rect 14382 2385 14390 2437
rect 14416 2385 14434 2437
rect 14434 2385 14446 2437
rect 14446 2385 14472 2437
rect 14498 2385 14510 2437
rect 14510 2385 14554 2437
rect 14579 2385 14626 2437
rect 14626 2385 14635 2437
rect 14660 2385 14690 2437
rect 14690 2385 14702 2437
rect 14702 2385 14716 2437
rect 14741 2385 14754 2437
rect 14754 2385 14766 2437
rect 14766 2385 14797 2437
rect 14822 2385 14830 2437
rect 14830 2385 14878 2437
rect 14006 2381 14062 2385
rect 14088 2381 14144 2385
rect 14170 2381 14226 2385
rect 14252 2381 14308 2385
rect 14334 2381 14390 2385
rect 14416 2381 14472 2385
rect 14498 2381 14554 2385
rect 14579 2381 14635 2385
rect 14660 2381 14716 2385
rect 14741 2381 14797 2385
rect 14822 2381 14878 2385
rect 14006 2317 14047 2353
rect 14047 2317 14060 2353
rect 14060 2317 14062 2353
rect 14088 2317 14112 2353
rect 14112 2317 14125 2353
rect 14125 2317 14144 2353
rect 14170 2317 14177 2353
rect 14177 2317 14190 2353
rect 14190 2317 14226 2353
rect 14252 2317 14254 2353
rect 14254 2317 14306 2353
rect 14306 2317 14308 2353
rect 14334 2317 14370 2353
rect 14370 2317 14382 2353
rect 14382 2317 14390 2353
rect 14416 2317 14434 2353
rect 14434 2317 14446 2353
rect 14446 2317 14472 2353
rect 14498 2317 14510 2353
rect 14510 2317 14554 2353
rect 14579 2317 14626 2353
rect 14626 2317 14635 2353
rect 14660 2317 14690 2353
rect 14690 2317 14702 2353
rect 14702 2317 14716 2353
rect 14741 2317 14754 2353
rect 14754 2317 14766 2353
rect 14766 2317 14797 2353
rect 14822 2317 14830 2353
rect 14830 2317 14878 2353
rect 14006 2301 14062 2317
rect 14088 2301 14144 2317
rect 14170 2301 14226 2317
rect 14252 2301 14308 2317
rect 14334 2301 14390 2317
rect 14416 2301 14472 2317
rect 14498 2301 14554 2317
rect 14579 2301 14635 2317
rect 14660 2301 14716 2317
rect 14741 2301 14797 2317
rect 14822 2301 14878 2317
rect 14006 2297 14047 2301
rect 14047 2297 14060 2301
rect 14060 2297 14062 2301
rect 14088 2297 14112 2301
rect 14112 2297 14125 2301
rect 14125 2297 14144 2301
rect 14170 2297 14177 2301
rect 14177 2297 14190 2301
rect 14190 2297 14226 2301
rect 14252 2297 14254 2301
rect 14254 2297 14306 2301
rect 14306 2297 14308 2301
rect 14334 2297 14370 2301
rect 14370 2297 14382 2301
rect 14382 2297 14390 2301
rect 14416 2297 14434 2301
rect 14434 2297 14446 2301
rect 14446 2297 14472 2301
rect 14498 2297 14510 2301
rect 14510 2297 14554 2301
rect 14006 2249 14047 2269
rect 14047 2249 14060 2269
rect 14060 2249 14062 2269
rect 14088 2249 14112 2269
rect 14112 2249 14125 2269
rect 14125 2249 14144 2269
rect 14170 2249 14177 2269
rect 14177 2249 14190 2269
rect 14190 2249 14226 2269
rect 14252 2249 14254 2269
rect 14254 2249 14306 2269
rect 14306 2249 14308 2269
rect 14334 2249 14370 2269
rect 14370 2249 14382 2269
rect 14382 2249 14390 2269
rect 14416 2249 14434 2269
rect 14434 2249 14446 2269
rect 14446 2249 14472 2269
rect 14498 2249 14510 2269
rect 14510 2249 14554 2269
rect 14579 2297 14626 2301
rect 14626 2297 14635 2301
rect 14660 2297 14690 2301
rect 14690 2297 14702 2301
rect 14702 2297 14716 2301
rect 14741 2297 14754 2301
rect 14754 2297 14766 2301
rect 14766 2297 14797 2301
rect 14822 2297 14830 2301
rect 14830 2297 14878 2301
rect 14579 2249 14626 2269
rect 14626 2249 14635 2269
rect 14660 2249 14690 2269
rect 14690 2249 14702 2269
rect 14702 2249 14716 2269
rect 14741 2249 14754 2269
rect 14754 2249 14766 2269
rect 14766 2249 14797 2269
rect 14822 2249 14830 2269
rect 14830 2249 14878 2269
rect 14006 2233 14062 2249
rect 14088 2233 14144 2249
rect 14170 2233 14226 2249
rect 14252 2233 14308 2249
rect 14334 2233 14390 2249
rect 14416 2233 14472 2249
rect 14498 2233 14554 2249
rect 14579 2233 14635 2249
rect 14660 2233 14716 2249
rect 14741 2233 14797 2249
rect 14822 2233 14878 2249
rect 14006 2213 14047 2233
rect 14047 2213 14060 2233
rect 14060 2213 14062 2233
rect 14088 2213 14112 2233
rect 14112 2213 14125 2233
rect 14125 2213 14144 2233
rect 14170 2213 14177 2233
rect 14177 2213 14190 2233
rect 14190 2213 14226 2233
rect 14252 2213 14254 2233
rect 14254 2213 14306 2233
rect 14306 2213 14308 2233
rect 14334 2213 14370 2233
rect 14370 2213 14382 2233
rect 14382 2213 14390 2233
rect 14416 2213 14434 2233
rect 14434 2213 14446 2233
rect 14446 2213 14472 2233
rect 14498 2213 14510 2233
rect 14510 2213 14554 2233
rect 14006 2181 14047 2185
rect 14047 2181 14060 2185
rect 14060 2181 14062 2185
rect 14088 2181 14112 2185
rect 14112 2181 14125 2185
rect 14125 2181 14144 2185
rect 14170 2181 14177 2185
rect 14177 2181 14190 2185
rect 14190 2181 14226 2185
rect 14252 2181 14254 2185
rect 14254 2181 14306 2185
rect 14306 2181 14308 2185
rect 14334 2181 14370 2185
rect 14370 2181 14382 2185
rect 14382 2181 14390 2185
rect 14416 2181 14434 2185
rect 14434 2181 14446 2185
rect 14446 2181 14472 2185
rect 14498 2181 14510 2185
rect 14510 2181 14554 2185
rect 14579 2213 14626 2233
rect 14626 2213 14635 2233
rect 14660 2213 14690 2233
rect 14690 2213 14702 2233
rect 14702 2213 14716 2233
rect 14741 2213 14754 2233
rect 14754 2213 14766 2233
rect 14766 2213 14797 2233
rect 14822 2213 14830 2233
rect 14830 2213 14878 2233
rect 14579 2181 14626 2185
rect 14626 2181 14635 2185
rect 14660 2181 14690 2185
rect 14690 2181 14702 2185
rect 14702 2181 14716 2185
rect 14741 2181 14754 2185
rect 14754 2181 14766 2185
rect 14766 2181 14797 2185
rect 14822 2181 14830 2185
rect 14830 2181 14878 2185
rect 14006 2165 14062 2181
rect 14088 2165 14144 2181
rect 14170 2165 14226 2181
rect 14252 2165 14308 2181
rect 14334 2165 14390 2181
rect 14416 2165 14472 2181
rect 14498 2165 14554 2181
rect 14579 2165 14635 2181
rect 14660 2165 14716 2181
rect 14741 2165 14797 2181
rect 14822 2165 14878 2181
rect 14006 2129 14047 2165
rect 14047 2129 14060 2165
rect 14060 2129 14062 2165
rect 14088 2129 14112 2165
rect 14112 2129 14125 2165
rect 14125 2129 14144 2165
rect 14170 2129 14177 2165
rect 14177 2129 14190 2165
rect 14190 2129 14226 2165
rect 14252 2129 14254 2165
rect 14254 2129 14306 2165
rect 14306 2129 14308 2165
rect 14334 2129 14370 2165
rect 14370 2129 14382 2165
rect 14382 2129 14390 2165
rect 14416 2129 14434 2165
rect 14434 2129 14446 2165
rect 14446 2129 14472 2165
rect 14498 2129 14510 2165
rect 14510 2129 14554 2165
rect 14579 2129 14626 2165
rect 14626 2129 14635 2165
rect 14660 2129 14690 2165
rect 14690 2129 14702 2165
rect 14702 2129 14716 2165
rect 14741 2129 14754 2165
rect 14754 2129 14766 2165
rect 14766 2129 14797 2165
rect 14822 2129 14830 2165
rect 14830 2129 14878 2165
rect 14006 2097 14062 2101
rect 14088 2097 14144 2101
rect 14170 2097 14226 2101
rect 14252 2097 14308 2101
rect 14334 2097 14390 2101
rect 14416 2097 14472 2101
rect 14498 2097 14554 2101
rect 14579 2097 14635 2101
rect 14660 2097 14716 2101
rect 14741 2097 14797 2101
rect 14822 2097 14878 2101
rect 14006 2045 14047 2097
rect 14047 2045 14060 2097
rect 14060 2045 14062 2097
rect 14088 2045 14112 2097
rect 14112 2045 14125 2097
rect 14125 2045 14144 2097
rect 14170 2045 14177 2097
rect 14177 2045 14190 2097
rect 14190 2045 14226 2097
rect 14252 2045 14254 2097
rect 14254 2045 14306 2097
rect 14306 2045 14308 2097
rect 14334 2045 14370 2097
rect 14370 2045 14382 2097
rect 14382 2045 14390 2097
rect 14416 2045 14434 2097
rect 14434 2045 14446 2097
rect 14446 2045 14472 2097
rect 14498 2045 14510 2097
rect 14510 2045 14554 2097
rect 14579 2045 14626 2097
rect 14626 2045 14635 2097
rect 14660 2045 14690 2097
rect 14690 2045 14702 2097
rect 14702 2045 14716 2097
rect 14741 2045 14754 2097
rect 14754 2045 14766 2097
rect 14766 2045 14797 2097
rect 14822 2045 14830 2097
rect 14830 2045 14878 2097
rect 17928 2385 17976 2437
rect 17976 2385 17984 2437
rect 18009 2385 18040 2437
rect 18040 2385 18052 2437
rect 18052 2385 18065 2437
rect 18090 2385 18104 2437
rect 18104 2385 18116 2437
rect 18116 2385 18146 2437
rect 18171 2385 18180 2437
rect 18180 2385 18227 2437
rect 18252 2385 18296 2437
rect 18296 2385 18308 2437
rect 18334 2385 18360 2437
rect 18360 2385 18372 2437
rect 18372 2385 18390 2437
rect 18416 2385 18424 2437
rect 18424 2385 18436 2437
rect 18436 2385 18472 2437
rect 18498 2385 18500 2437
rect 18500 2385 18552 2437
rect 18552 2385 18554 2437
rect 18580 2385 18616 2437
rect 18616 2385 18629 2437
rect 18629 2385 18636 2437
rect 18662 2385 18681 2437
rect 18681 2385 18694 2437
rect 18694 2385 18718 2437
rect 18744 2385 18746 2437
rect 18746 2385 18759 2437
rect 18759 2385 18800 2437
rect 17928 2381 17984 2385
rect 18009 2381 18065 2385
rect 18090 2381 18146 2385
rect 18171 2381 18227 2385
rect 18252 2381 18308 2385
rect 18334 2381 18390 2385
rect 18416 2381 18472 2385
rect 18498 2381 18554 2385
rect 18580 2381 18636 2385
rect 18662 2381 18718 2385
rect 18744 2381 18800 2385
rect 17928 2317 17976 2353
rect 17976 2317 17984 2353
rect 18009 2317 18040 2353
rect 18040 2317 18052 2353
rect 18052 2317 18065 2353
rect 18090 2317 18104 2353
rect 18104 2317 18116 2353
rect 18116 2317 18146 2353
rect 18171 2317 18180 2353
rect 18180 2317 18227 2353
rect 18252 2317 18296 2353
rect 18296 2317 18308 2353
rect 18334 2317 18360 2353
rect 18360 2317 18372 2353
rect 18372 2317 18390 2353
rect 18416 2317 18424 2353
rect 18424 2317 18436 2353
rect 18436 2317 18472 2353
rect 18498 2317 18500 2353
rect 18500 2317 18552 2353
rect 18552 2317 18554 2353
rect 18580 2317 18616 2353
rect 18616 2317 18629 2353
rect 18629 2317 18636 2353
rect 18662 2317 18681 2353
rect 18681 2317 18694 2353
rect 18694 2317 18718 2353
rect 18744 2317 18746 2353
rect 18746 2317 18759 2353
rect 18759 2317 18800 2353
rect 17928 2301 17984 2317
rect 18009 2301 18065 2317
rect 18090 2301 18146 2317
rect 18171 2301 18227 2317
rect 18252 2301 18308 2317
rect 18334 2301 18390 2317
rect 18416 2301 18472 2317
rect 18498 2301 18554 2317
rect 18580 2301 18636 2317
rect 18662 2301 18718 2317
rect 18744 2301 18800 2317
rect 17928 2297 17976 2301
rect 17976 2297 17984 2301
rect 18009 2297 18040 2301
rect 18040 2297 18052 2301
rect 18052 2297 18065 2301
rect 18090 2297 18104 2301
rect 18104 2297 18116 2301
rect 18116 2297 18146 2301
rect 18171 2297 18180 2301
rect 18180 2297 18227 2301
rect 17928 2249 17976 2269
rect 17976 2249 17984 2269
rect 18009 2249 18040 2269
rect 18040 2249 18052 2269
rect 18052 2249 18065 2269
rect 18090 2249 18104 2269
rect 18104 2249 18116 2269
rect 18116 2249 18146 2269
rect 18171 2249 18180 2269
rect 18180 2249 18227 2269
rect 18252 2297 18296 2301
rect 18296 2297 18308 2301
rect 18334 2297 18360 2301
rect 18360 2297 18372 2301
rect 18372 2297 18390 2301
rect 18416 2297 18424 2301
rect 18424 2297 18436 2301
rect 18436 2297 18472 2301
rect 18498 2297 18500 2301
rect 18500 2297 18552 2301
rect 18552 2297 18554 2301
rect 18580 2297 18616 2301
rect 18616 2297 18629 2301
rect 18629 2297 18636 2301
rect 18662 2297 18681 2301
rect 18681 2297 18694 2301
rect 18694 2297 18718 2301
rect 18744 2297 18746 2301
rect 18746 2297 18759 2301
rect 18759 2297 18800 2301
rect 18252 2249 18296 2269
rect 18296 2249 18308 2269
rect 18334 2249 18360 2269
rect 18360 2249 18372 2269
rect 18372 2249 18390 2269
rect 18416 2249 18424 2269
rect 18424 2249 18436 2269
rect 18436 2249 18472 2269
rect 18498 2249 18500 2269
rect 18500 2249 18552 2269
rect 18552 2249 18554 2269
rect 18580 2249 18616 2269
rect 18616 2249 18629 2269
rect 18629 2249 18636 2269
rect 18662 2249 18681 2269
rect 18681 2249 18694 2269
rect 18694 2249 18718 2269
rect 18744 2249 18746 2269
rect 18746 2249 18759 2269
rect 18759 2249 18800 2269
rect 17928 2233 17984 2249
rect 18009 2233 18065 2249
rect 18090 2233 18146 2249
rect 18171 2233 18227 2249
rect 18252 2233 18308 2249
rect 18334 2233 18390 2249
rect 18416 2233 18472 2249
rect 18498 2233 18554 2249
rect 18580 2233 18636 2249
rect 18662 2233 18718 2249
rect 18744 2233 18800 2249
rect 17928 2213 17976 2233
rect 17976 2213 17984 2233
rect 18009 2213 18040 2233
rect 18040 2213 18052 2233
rect 18052 2213 18065 2233
rect 18090 2213 18104 2233
rect 18104 2213 18116 2233
rect 18116 2213 18146 2233
rect 18171 2213 18180 2233
rect 18180 2213 18227 2233
rect 17928 2181 17976 2185
rect 17976 2181 17984 2185
rect 18009 2181 18040 2185
rect 18040 2181 18052 2185
rect 18052 2181 18065 2185
rect 18090 2181 18104 2185
rect 18104 2181 18116 2185
rect 18116 2181 18146 2185
rect 18171 2181 18180 2185
rect 18180 2181 18227 2185
rect 18252 2213 18296 2233
rect 18296 2213 18308 2233
rect 18334 2213 18360 2233
rect 18360 2213 18372 2233
rect 18372 2213 18390 2233
rect 18416 2213 18424 2233
rect 18424 2213 18436 2233
rect 18436 2213 18472 2233
rect 18498 2213 18500 2233
rect 18500 2213 18552 2233
rect 18552 2213 18554 2233
rect 18580 2213 18616 2233
rect 18616 2213 18629 2233
rect 18629 2213 18636 2233
rect 18662 2213 18681 2233
rect 18681 2213 18694 2233
rect 18694 2213 18718 2233
rect 18744 2213 18746 2233
rect 18746 2213 18759 2233
rect 18759 2213 18800 2233
rect 18252 2181 18296 2185
rect 18296 2181 18308 2185
rect 18334 2181 18360 2185
rect 18360 2181 18372 2185
rect 18372 2181 18390 2185
rect 18416 2181 18424 2185
rect 18424 2181 18436 2185
rect 18436 2181 18472 2185
rect 18498 2181 18500 2185
rect 18500 2181 18552 2185
rect 18552 2181 18554 2185
rect 18580 2181 18616 2185
rect 18616 2181 18629 2185
rect 18629 2181 18636 2185
rect 18662 2181 18681 2185
rect 18681 2181 18694 2185
rect 18694 2181 18718 2185
rect 18744 2181 18746 2185
rect 18746 2181 18759 2185
rect 18759 2181 18800 2185
rect 17928 2165 17984 2181
rect 18009 2165 18065 2181
rect 18090 2165 18146 2181
rect 18171 2165 18227 2181
rect 18252 2165 18308 2181
rect 18334 2165 18390 2181
rect 18416 2165 18472 2181
rect 18498 2165 18554 2181
rect 18580 2165 18636 2181
rect 18662 2165 18718 2181
rect 18744 2165 18800 2181
rect 17928 2129 17976 2165
rect 17976 2129 17984 2165
rect 18009 2129 18040 2165
rect 18040 2129 18052 2165
rect 18052 2129 18065 2165
rect 18090 2129 18104 2165
rect 18104 2129 18116 2165
rect 18116 2129 18146 2165
rect 18171 2129 18180 2165
rect 18180 2129 18227 2165
rect 18252 2129 18296 2165
rect 18296 2129 18308 2165
rect 18334 2129 18360 2165
rect 18360 2129 18372 2165
rect 18372 2129 18390 2165
rect 18416 2129 18424 2165
rect 18424 2129 18436 2165
rect 18436 2129 18472 2165
rect 18498 2129 18500 2165
rect 18500 2129 18552 2165
rect 18552 2129 18554 2165
rect 18580 2129 18616 2165
rect 18616 2129 18629 2165
rect 18629 2129 18636 2165
rect 18662 2129 18681 2165
rect 18681 2129 18694 2165
rect 18694 2129 18718 2165
rect 18744 2129 18746 2165
rect 18746 2129 18759 2165
rect 18759 2129 18800 2165
rect 17928 2097 17984 2101
rect 18009 2097 18065 2101
rect 18090 2097 18146 2101
rect 18171 2097 18227 2101
rect 18252 2097 18308 2101
rect 18334 2097 18390 2101
rect 18416 2097 18472 2101
rect 18498 2097 18554 2101
rect 18580 2097 18636 2101
rect 18662 2097 18718 2101
rect 18744 2097 18800 2101
rect 17928 2045 17976 2097
rect 17976 2045 17984 2097
rect 18009 2045 18040 2097
rect 18040 2045 18052 2097
rect 18052 2045 18065 2097
rect 18090 2045 18104 2097
rect 18104 2045 18116 2097
rect 18116 2045 18146 2097
rect 18171 2045 18180 2097
rect 18180 2045 18227 2097
rect 18252 2045 18296 2097
rect 18296 2045 18308 2097
rect 18334 2045 18360 2097
rect 18360 2045 18372 2097
rect 18372 2045 18390 2097
rect 18416 2045 18424 2097
rect 18424 2045 18436 2097
rect 18436 2045 18472 2097
rect 18498 2045 18500 2097
rect 18500 2045 18552 2097
rect 18552 2045 18554 2097
rect 18580 2045 18616 2097
rect 18616 2045 18629 2097
rect 18629 2045 18636 2097
rect 18662 2045 18681 2097
rect 18681 2045 18694 2097
rect 18694 2045 18718 2097
rect 18744 2045 18746 2097
rect 18746 2045 18759 2097
rect 18759 2045 18800 2097
rect 647 1867 696 1919
rect 696 1867 703 1919
rect 647 1863 703 1867
rect 728 1867 780 1919
rect 780 1867 784 1919
rect 728 1863 784 1867
rect 808 1867 812 1919
rect 812 1867 864 1919
rect 808 1863 864 1867
rect 888 1867 895 1919
rect 895 1867 944 1919
rect 888 1863 944 1867
rect 647 1791 703 1795
rect 647 1739 696 1791
rect 696 1739 703 1791
rect 728 1791 784 1795
rect 728 1739 780 1791
rect 780 1739 784 1791
rect 808 1791 864 1795
rect 808 1739 812 1791
rect 812 1739 864 1791
rect 888 1791 944 1795
rect 888 1739 895 1791
rect 895 1739 944 1791
rect 6021 1867 6070 1919
rect 6070 1867 6077 1919
rect 6102 1867 6137 1919
rect 6137 1867 6152 1919
rect 6152 1867 6158 1919
rect 6183 1867 6204 1919
rect 6204 1867 6219 1919
rect 6219 1867 6239 1919
rect 6264 1867 6271 1919
rect 6271 1867 6286 1919
rect 6286 1867 6320 1919
rect 6346 1867 6353 1919
rect 6353 1867 6402 1919
rect 6021 1863 6077 1867
rect 6102 1863 6158 1867
rect 6183 1863 6239 1867
rect 6264 1863 6320 1867
rect 6346 1863 6402 1867
rect 6021 1791 6077 1795
rect 6102 1791 6158 1795
rect 6183 1791 6239 1795
rect 6264 1791 6320 1795
rect 6346 1791 6402 1795
rect 6021 1739 6070 1791
rect 6070 1739 6077 1791
rect 6102 1739 6137 1791
rect 6137 1739 6152 1791
rect 6152 1739 6158 1791
rect 6183 1739 6204 1791
rect 6204 1739 6219 1791
rect 6219 1739 6239 1791
rect 6264 1739 6271 1791
rect 6271 1739 6286 1791
rect 6286 1739 6320 1791
rect 6346 1739 6353 1791
rect 6353 1739 6402 1791
rect 6952 1867 7001 1919
rect 7001 1867 7008 1919
rect 7034 1867 7068 1919
rect 7068 1867 7083 1919
rect 7083 1867 7090 1919
rect 7115 1867 7135 1919
rect 7135 1867 7150 1919
rect 7150 1867 7171 1919
rect 7196 1867 7202 1919
rect 7202 1867 7217 1919
rect 7217 1867 7252 1919
rect 7277 1867 7284 1919
rect 7284 1867 7333 1919
rect 6952 1863 7008 1867
rect 7034 1863 7090 1867
rect 7115 1863 7171 1867
rect 7196 1863 7252 1867
rect 7277 1863 7333 1867
rect 6952 1791 7008 1795
rect 7034 1791 7090 1795
rect 7115 1791 7171 1795
rect 7196 1791 7252 1795
rect 7277 1791 7333 1795
rect 6952 1739 7001 1791
rect 7001 1739 7008 1791
rect 7034 1739 7068 1791
rect 7068 1739 7083 1791
rect 7083 1739 7090 1791
rect 7115 1739 7135 1791
rect 7135 1739 7150 1791
rect 7150 1739 7171 1791
rect 7196 1739 7202 1791
rect 7202 1739 7217 1791
rect 7217 1739 7252 1791
rect 7277 1739 7284 1791
rect 7284 1739 7333 1791
rect 12505 1867 12554 1919
rect 12554 1867 12561 1919
rect 12586 1867 12621 1919
rect 12621 1867 12636 1919
rect 12636 1867 12642 1919
rect 12667 1867 12688 1919
rect 12688 1867 12703 1919
rect 12703 1867 12723 1919
rect 12748 1867 12755 1919
rect 12755 1867 12770 1919
rect 12770 1867 12804 1919
rect 12830 1867 12837 1919
rect 12837 1867 12886 1919
rect 12505 1863 12561 1867
rect 12586 1863 12642 1867
rect 12667 1863 12723 1867
rect 12748 1863 12804 1867
rect 12830 1863 12886 1867
rect 12505 1791 12561 1795
rect 12586 1791 12642 1795
rect 12667 1791 12723 1795
rect 12748 1791 12804 1795
rect 12830 1791 12886 1795
rect 12505 1739 12554 1791
rect 12554 1739 12561 1791
rect 12586 1739 12621 1791
rect 12621 1739 12636 1791
rect 12636 1739 12642 1791
rect 12667 1739 12688 1791
rect 12688 1739 12703 1791
rect 12703 1739 12723 1791
rect 12748 1739 12755 1791
rect 12755 1739 12770 1791
rect 12770 1739 12804 1791
rect 12830 1739 12837 1791
rect 12837 1739 12886 1791
rect 13436 1867 13485 1919
rect 13485 1867 13492 1919
rect 13518 1867 13552 1919
rect 13552 1867 13567 1919
rect 13567 1867 13574 1919
rect 13599 1867 13619 1919
rect 13619 1867 13634 1919
rect 13634 1867 13655 1919
rect 13680 1867 13686 1919
rect 13686 1867 13701 1919
rect 13701 1867 13736 1919
rect 13761 1867 13768 1919
rect 13768 1867 13817 1919
rect 13436 1863 13492 1867
rect 13518 1863 13574 1867
rect 13599 1863 13655 1867
rect 13680 1863 13736 1867
rect 13761 1863 13817 1867
rect 13436 1791 13492 1795
rect 13518 1791 13574 1795
rect 13599 1791 13655 1795
rect 13680 1791 13736 1795
rect 13761 1791 13817 1795
rect 13436 1739 13485 1791
rect 13485 1739 13492 1791
rect 13518 1739 13552 1791
rect 13552 1739 13567 1791
rect 13567 1739 13574 1791
rect 13599 1739 13619 1791
rect 13619 1739 13634 1791
rect 13634 1739 13655 1791
rect 13680 1739 13686 1791
rect 13686 1739 13701 1791
rect 13701 1739 13736 1791
rect 13761 1739 13768 1791
rect 13768 1739 13817 1791
rect 19074 1867 19123 1919
rect 19123 1867 19130 1919
rect 19074 1863 19130 1867
rect 19154 1867 19206 1919
rect 19206 1867 19210 1919
rect 19154 1863 19210 1867
rect 19234 1867 19237 1919
rect 19237 1867 19289 1919
rect 19289 1867 19290 1919
rect 19234 1863 19290 1867
rect 19314 1867 19321 1919
rect 19321 1867 19370 1919
rect 19314 1863 19370 1867
rect 19074 1791 19130 1795
rect 19074 1739 19123 1791
rect 19123 1739 19130 1791
rect 19154 1791 19210 1795
rect 19154 1739 19206 1791
rect 19206 1739 19210 1791
rect 19234 1791 19290 1795
rect 19234 1739 19237 1791
rect 19237 1739 19289 1791
rect 19289 1739 19290 1791
rect 19314 1791 19370 1795
rect 19314 1739 19321 1791
rect 19321 1739 19370 1791
rect 2680 1633 2729 1682
rect 2729 1633 2736 1682
rect 2766 1633 2796 1682
rect 2796 1633 2811 1682
rect 2811 1633 2822 1682
rect 2852 1633 2863 1682
rect 2863 1633 2878 1682
rect 2878 1633 2908 1682
rect 2938 1633 2945 1682
rect 2945 1633 2994 1682
rect 3024 1633 3064 1682
rect 3064 1633 3079 1682
rect 3079 1633 3080 1682
rect 3110 1633 3131 1682
rect 3131 1633 3146 1682
rect 3146 1633 3166 1682
rect 3196 1633 3198 1682
rect 3198 1633 3213 1682
rect 3213 1633 3252 1682
rect 3281 1633 3331 1682
rect 3331 1633 3337 1682
rect 3366 1633 3397 1682
rect 3397 1633 3411 1682
rect 3411 1633 3422 1682
rect 3451 1633 3463 1682
rect 3463 1633 3477 1682
rect 3477 1633 3507 1682
rect 3536 1633 3543 1682
rect 3543 1633 3592 1682
rect 2680 1626 2736 1633
rect 2766 1626 2822 1633
rect 2852 1626 2908 1633
rect 2938 1626 2994 1633
rect 3024 1626 3080 1633
rect 3110 1626 3166 1633
rect 3196 1626 3252 1633
rect 3281 1626 3337 1633
rect 3366 1626 3422 1633
rect 3451 1626 3507 1633
rect 3536 1626 3592 1633
rect 2680 1541 2736 1548
rect 2766 1541 2822 1548
rect 2852 1541 2908 1548
rect 2938 1541 2994 1548
rect 3024 1541 3080 1548
rect 3110 1541 3166 1548
rect 3196 1541 3252 1548
rect 3281 1541 3337 1548
rect 3366 1541 3422 1548
rect 3451 1541 3507 1548
rect 3536 1541 3592 1548
rect 2680 1492 2729 1541
rect 2729 1492 2736 1541
rect 2766 1492 2796 1541
rect 2796 1492 2811 1541
rect 2811 1492 2822 1541
rect 2852 1492 2863 1541
rect 2863 1492 2878 1541
rect 2878 1492 2908 1541
rect 2938 1492 2945 1541
rect 2945 1492 2994 1541
rect 3024 1492 3064 1541
rect 3064 1492 3079 1541
rect 3079 1492 3080 1541
rect 3110 1492 3131 1541
rect 3131 1492 3146 1541
rect 3146 1492 3166 1541
rect 3196 1492 3198 1541
rect 3198 1492 3213 1541
rect 3213 1492 3252 1541
rect 3281 1492 3331 1541
rect 3331 1492 3337 1541
rect 3366 1492 3397 1541
rect 3397 1492 3411 1541
rect 3411 1492 3422 1541
rect 3451 1492 3463 1541
rect 3463 1492 3477 1541
rect 3477 1492 3507 1541
rect 3536 1492 3543 1541
rect 3543 1492 3592 1541
rect 4885 1633 4934 1682
rect 4934 1633 4941 1682
rect 4885 1626 4941 1633
rect 4969 1633 4971 1682
rect 4971 1633 5023 1682
rect 5023 1633 5025 1682
rect 4969 1626 5025 1633
rect 5052 1633 5059 1682
rect 5059 1633 5108 1682
rect 5052 1626 5108 1633
rect 4885 1541 4941 1548
rect 4885 1492 4934 1541
rect 4934 1492 4941 1541
rect 4969 1541 5025 1548
rect 4969 1492 4971 1541
rect 4971 1492 5023 1541
rect 5023 1492 5025 1541
rect 5052 1541 5108 1548
rect 5052 1492 5059 1541
rect 5059 1492 5108 1541
rect 5722 1633 5772 1682
rect 5772 1633 5778 1682
rect 5871 1633 5878 1682
rect 5878 1633 5927 1682
rect 5722 1626 5778 1633
rect 5871 1626 5927 1633
rect 5722 1541 5778 1548
rect 5871 1541 5927 1548
rect 5722 1492 5772 1541
rect 5772 1492 5778 1541
rect 5871 1492 5878 1541
rect 5878 1492 5927 1541
rect 6496 1685 6552 1686
rect 6598 1685 6654 1686
rect 6700 1685 6756 1686
rect 6802 1685 6858 1686
rect 6496 1633 6497 1685
rect 6497 1633 6549 1685
rect 6549 1633 6552 1685
rect 6598 1633 6626 1685
rect 6626 1633 6651 1685
rect 6651 1633 6654 1685
rect 6700 1633 6703 1685
rect 6703 1633 6728 1685
rect 6728 1633 6756 1685
rect 6802 1633 6805 1685
rect 6805 1633 6857 1685
rect 6857 1633 6858 1685
rect 6496 1630 6552 1633
rect 6598 1630 6654 1633
rect 6700 1630 6756 1633
rect 6802 1630 6858 1633
rect 6496 1541 6552 1552
rect 6598 1541 6654 1552
rect 6700 1541 6756 1552
rect 6802 1541 6858 1552
rect 6496 1496 6497 1541
rect 6497 1496 6549 1541
rect 6549 1496 6552 1541
rect 6598 1496 6626 1541
rect 6626 1496 6651 1541
rect 6651 1496 6654 1541
rect 6700 1496 6703 1541
rect 6703 1496 6728 1541
rect 6728 1496 6756 1541
rect 6802 1496 6805 1541
rect 6805 1496 6857 1541
rect 6857 1496 6858 1541
rect 9528 1633 9577 1682
rect 9577 1633 9584 1682
rect 9624 1633 9644 1682
rect 9644 1633 9659 1682
rect 9659 1633 9680 1682
rect 9719 1633 9726 1682
rect 9726 1633 9775 1682
rect 9528 1626 9584 1633
rect 9624 1626 9680 1633
rect 9719 1626 9775 1633
rect 9528 1541 9584 1548
rect 9624 1541 9680 1548
rect 9719 1541 9775 1548
rect 9528 1492 9577 1541
rect 9577 1492 9584 1541
rect 9624 1492 9644 1541
rect 9644 1492 9659 1541
rect 9659 1492 9680 1541
rect 9719 1492 9726 1541
rect 9726 1492 9775 1541
rect 16406 1633 16455 1682
rect 16455 1633 16462 1682
rect 16488 1633 16523 1682
rect 16523 1633 16539 1682
rect 16539 1633 16544 1682
rect 16570 1633 16591 1682
rect 16591 1633 16607 1682
rect 16607 1633 16626 1682
rect 16652 1633 16659 1682
rect 16659 1633 16674 1682
rect 16674 1633 16708 1682
rect 16734 1633 16741 1682
rect 16741 1633 16790 1682
rect 16406 1626 16462 1633
rect 16488 1626 16544 1633
rect 16570 1626 16626 1633
rect 16652 1626 16708 1633
rect 16734 1626 16790 1633
rect 16406 1541 16462 1548
rect 16488 1541 16544 1548
rect 16570 1541 16626 1548
rect 16652 1541 16708 1548
rect 16734 1541 16790 1548
rect 16406 1492 16455 1541
rect 16455 1492 16462 1541
rect 16488 1492 16523 1541
rect 16523 1492 16539 1541
rect 16539 1492 16544 1541
rect 16570 1492 16591 1541
rect 16591 1492 16607 1541
rect 16607 1492 16626 1541
rect 16652 1492 16659 1541
rect 16659 1492 16674 1541
rect 16674 1492 16708 1541
rect 16734 1492 16741 1541
rect 16741 1492 16790 1541
rect 1038 1319 1079 1371
rect 1079 1319 1092 1371
rect 1092 1319 1094 1371
rect 1120 1319 1144 1371
rect 1144 1319 1157 1371
rect 1157 1319 1176 1371
rect 1202 1319 1209 1371
rect 1209 1319 1222 1371
rect 1222 1319 1258 1371
rect 1284 1319 1286 1371
rect 1286 1319 1338 1371
rect 1338 1319 1340 1371
rect 1366 1319 1402 1371
rect 1402 1319 1414 1371
rect 1414 1319 1422 1371
rect 1448 1319 1466 1371
rect 1466 1319 1478 1371
rect 1478 1319 1504 1371
rect 1530 1319 1542 1371
rect 1542 1319 1586 1371
rect 1611 1319 1658 1371
rect 1658 1319 1667 1371
rect 1692 1319 1722 1371
rect 1722 1319 1734 1371
rect 1734 1319 1748 1371
rect 1773 1319 1786 1371
rect 1786 1319 1798 1371
rect 1798 1319 1829 1371
rect 1854 1319 1862 1371
rect 1862 1319 1910 1371
rect 1038 1315 1094 1319
rect 1120 1315 1176 1319
rect 1202 1315 1258 1319
rect 1284 1315 1340 1319
rect 1366 1315 1422 1319
rect 1448 1315 1504 1319
rect 1530 1315 1586 1319
rect 1611 1315 1667 1319
rect 1692 1315 1748 1319
rect 1773 1315 1829 1319
rect 1854 1315 1910 1319
rect 1038 1251 1079 1287
rect 1079 1251 1092 1287
rect 1092 1251 1094 1287
rect 1120 1251 1144 1287
rect 1144 1251 1157 1287
rect 1157 1251 1176 1287
rect 1202 1251 1209 1287
rect 1209 1251 1222 1287
rect 1222 1251 1258 1287
rect 1284 1251 1286 1287
rect 1286 1251 1338 1287
rect 1338 1251 1340 1287
rect 1366 1251 1402 1287
rect 1402 1251 1414 1287
rect 1414 1251 1422 1287
rect 1448 1251 1466 1287
rect 1466 1251 1478 1287
rect 1478 1251 1504 1287
rect 1530 1251 1542 1287
rect 1542 1251 1586 1287
rect 1611 1251 1658 1287
rect 1658 1251 1667 1287
rect 1692 1251 1722 1287
rect 1722 1251 1734 1287
rect 1734 1251 1748 1287
rect 1773 1251 1786 1287
rect 1786 1251 1798 1287
rect 1798 1251 1829 1287
rect 1854 1251 1862 1287
rect 1862 1251 1910 1287
rect 1038 1235 1094 1251
rect 1120 1235 1176 1251
rect 1202 1235 1258 1251
rect 1284 1235 1340 1251
rect 1366 1235 1422 1251
rect 1448 1235 1504 1251
rect 1530 1235 1586 1251
rect 1611 1235 1667 1251
rect 1692 1235 1748 1251
rect 1773 1235 1829 1251
rect 1854 1235 1910 1251
rect 1038 1231 1079 1235
rect 1079 1231 1092 1235
rect 1092 1231 1094 1235
rect 1120 1231 1144 1235
rect 1144 1231 1157 1235
rect 1157 1231 1176 1235
rect 1202 1231 1209 1235
rect 1209 1231 1222 1235
rect 1222 1231 1258 1235
rect 1284 1231 1286 1235
rect 1286 1231 1338 1235
rect 1338 1231 1340 1235
rect 1366 1231 1402 1235
rect 1402 1231 1414 1235
rect 1414 1231 1422 1235
rect 1448 1231 1466 1235
rect 1466 1231 1478 1235
rect 1478 1231 1504 1235
rect 1530 1231 1542 1235
rect 1542 1231 1586 1235
rect 1038 1183 1079 1203
rect 1079 1183 1092 1203
rect 1092 1183 1094 1203
rect 1120 1183 1144 1203
rect 1144 1183 1157 1203
rect 1157 1183 1176 1203
rect 1202 1183 1209 1203
rect 1209 1183 1222 1203
rect 1222 1183 1258 1203
rect 1284 1183 1286 1203
rect 1286 1183 1338 1203
rect 1338 1183 1340 1203
rect 1366 1183 1402 1203
rect 1402 1183 1414 1203
rect 1414 1183 1422 1203
rect 1448 1183 1466 1203
rect 1466 1183 1478 1203
rect 1478 1183 1504 1203
rect 1530 1183 1542 1203
rect 1542 1183 1586 1203
rect 1611 1231 1658 1235
rect 1658 1231 1667 1235
rect 1692 1231 1722 1235
rect 1722 1231 1734 1235
rect 1734 1231 1748 1235
rect 1773 1231 1786 1235
rect 1786 1231 1798 1235
rect 1798 1231 1829 1235
rect 1854 1231 1862 1235
rect 1862 1231 1910 1235
rect 1611 1183 1658 1203
rect 1658 1183 1667 1203
rect 1692 1183 1722 1203
rect 1722 1183 1734 1203
rect 1734 1183 1748 1203
rect 1773 1183 1786 1203
rect 1786 1183 1798 1203
rect 1798 1183 1829 1203
rect 1854 1183 1862 1203
rect 1862 1183 1910 1203
rect 1038 1167 1094 1183
rect 1120 1167 1176 1183
rect 1202 1167 1258 1183
rect 1284 1167 1340 1183
rect 1366 1167 1422 1183
rect 1448 1167 1504 1183
rect 1530 1167 1586 1183
rect 1611 1167 1667 1183
rect 1692 1167 1748 1183
rect 1773 1167 1829 1183
rect 1854 1167 1910 1183
rect 1038 1147 1079 1167
rect 1079 1147 1092 1167
rect 1092 1147 1094 1167
rect 1120 1147 1144 1167
rect 1144 1147 1157 1167
rect 1157 1147 1176 1167
rect 1202 1147 1209 1167
rect 1209 1147 1222 1167
rect 1222 1147 1258 1167
rect 1284 1147 1286 1167
rect 1286 1147 1338 1167
rect 1338 1147 1340 1167
rect 1366 1147 1402 1167
rect 1402 1147 1414 1167
rect 1414 1147 1422 1167
rect 1448 1147 1466 1167
rect 1466 1147 1478 1167
rect 1478 1147 1504 1167
rect 1530 1147 1542 1167
rect 1542 1147 1586 1167
rect 1038 1115 1079 1119
rect 1079 1115 1092 1119
rect 1092 1115 1094 1119
rect 1120 1115 1144 1119
rect 1144 1115 1157 1119
rect 1157 1115 1176 1119
rect 1202 1115 1209 1119
rect 1209 1115 1222 1119
rect 1222 1115 1258 1119
rect 1284 1115 1286 1119
rect 1286 1115 1338 1119
rect 1338 1115 1340 1119
rect 1366 1115 1402 1119
rect 1402 1115 1414 1119
rect 1414 1115 1422 1119
rect 1448 1115 1466 1119
rect 1466 1115 1478 1119
rect 1478 1115 1504 1119
rect 1530 1115 1542 1119
rect 1542 1115 1586 1119
rect 1611 1147 1658 1167
rect 1658 1147 1667 1167
rect 1692 1147 1722 1167
rect 1722 1147 1734 1167
rect 1734 1147 1748 1167
rect 1773 1147 1786 1167
rect 1786 1147 1798 1167
rect 1798 1147 1829 1167
rect 1854 1147 1862 1167
rect 1862 1147 1910 1167
rect 1611 1115 1658 1119
rect 1658 1115 1667 1119
rect 1692 1115 1722 1119
rect 1722 1115 1734 1119
rect 1734 1115 1748 1119
rect 1773 1115 1786 1119
rect 1786 1115 1798 1119
rect 1798 1115 1829 1119
rect 1854 1115 1862 1119
rect 1862 1115 1910 1119
rect 1038 1099 1094 1115
rect 1120 1099 1176 1115
rect 1202 1099 1258 1115
rect 1284 1099 1340 1115
rect 1366 1099 1422 1115
rect 1448 1099 1504 1115
rect 1530 1099 1586 1115
rect 1611 1099 1667 1115
rect 1692 1099 1748 1115
rect 1773 1099 1829 1115
rect 1854 1099 1910 1115
rect 1038 1063 1079 1099
rect 1079 1063 1092 1099
rect 1092 1063 1094 1099
rect 1120 1063 1144 1099
rect 1144 1063 1157 1099
rect 1157 1063 1176 1099
rect 1202 1063 1209 1099
rect 1209 1063 1222 1099
rect 1222 1063 1258 1099
rect 1284 1063 1286 1099
rect 1286 1063 1338 1099
rect 1338 1063 1340 1099
rect 1366 1063 1402 1099
rect 1402 1063 1414 1099
rect 1414 1063 1422 1099
rect 1448 1063 1466 1099
rect 1466 1063 1478 1099
rect 1478 1063 1504 1099
rect 1530 1063 1542 1099
rect 1542 1063 1586 1099
rect 1611 1063 1658 1099
rect 1658 1063 1667 1099
rect 1692 1063 1722 1099
rect 1722 1063 1734 1099
rect 1734 1063 1748 1099
rect 1773 1063 1786 1099
rect 1786 1063 1798 1099
rect 1798 1063 1829 1099
rect 1854 1063 1862 1099
rect 1862 1063 1910 1099
rect 1038 1031 1094 1035
rect 1120 1031 1176 1035
rect 1202 1031 1258 1035
rect 1284 1031 1340 1035
rect 1366 1031 1422 1035
rect 1448 1031 1504 1035
rect 1530 1031 1586 1035
rect 1611 1031 1667 1035
rect 1692 1031 1748 1035
rect 1773 1031 1829 1035
rect 1854 1031 1910 1035
rect 1038 979 1079 1031
rect 1079 979 1092 1031
rect 1092 979 1094 1031
rect 1120 979 1144 1031
rect 1144 979 1157 1031
rect 1157 979 1176 1031
rect 1202 979 1209 1031
rect 1209 979 1222 1031
rect 1222 979 1258 1031
rect 1284 979 1286 1031
rect 1286 979 1338 1031
rect 1338 979 1340 1031
rect 1366 979 1402 1031
rect 1402 979 1414 1031
rect 1414 979 1422 1031
rect 1448 979 1466 1031
rect 1466 979 1478 1031
rect 1478 979 1504 1031
rect 1530 979 1542 1031
rect 1542 979 1586 1031
rect 1611 979 1658 1031
rect 1658 979 1667 1031
rect 1692 979 1722 1031
rect 1722 979 1734 1031
rect 1734 979 1748 1031
rect 1773 979 1786 1031
rect 1786 979 1798 1031
rect 1798 979 1829 1031
rect 1854 979 1862 1031
rect 1862 979 1910 1031
rect 1038 495 1079 547
rect 1079 495 1092 547
rect 1092 495 1094 547
rect 1120 495 1144 547
rect 1144 495 1157 547
rect 1157 495 1176 547
rect 1202 495 1209 547
rect 1209 495 1222 547
rect 1222 495 1258 547
rect 1284 495 1286 547
rect 1286 495 1338 547
rect 1338 495 1340 547
rect 1366 495 1402 547
rect 1402 495 1414 547
rect 1414 495 1422 547
rect 1448 495 1466 547
rect 1466 495 1478 547
rect 1478 495 1504 547
rect 1530 495 1542 547
rect 1542 495 1586 547
rect 1611 495 1658 547
rect 1658 495 1667 547
rect 1692 495 1722 547
rect 1722 495 1734 547
rect 1734 495 1748 547
rect 1773 495 1786 547
rect 1786 495 1798 547
rect 1798 495 1829 547
rect 1854 495 1862 547
rect 1862 495 1910 547
rect 1038 491 1094 495
rect 1120 491 1176 495
rect 1202 491 1258 495
rect 1284 491 1340 495
rect 1366 491 1422 495
rect 1448 491 1504 495
rect 1530 491 1586 495
rect 1611 491 1667 495
rect 1692 491 1748 495
rect 1773 491 1829 495
rect 1854 491 1910 495
rect 1038 427 1079 463
rect 1079 427 1092 463
rect 1092 427 1094 463
rect 1120 427 1144 463
rect 1144 427 1157 463
rect 1157 427 1176 463
rect 1202 427 1209 463
rect 1209 427 1222 463
rect 1222 427 1258 463
rect 1284 427 1286 463
rect 1286 427 1338 463
rect 1338 427 1340 463
rect 1366 427 1402 463
rect 1402 427 1414 463
rect 1414 427 1422 463
rect 1448 427 1466 463
rect 1466 427 1478 463
rect 1478 427 1504 463
rect 1530 427 1542 463
rect 1542 427 1586 463
rect 1611 427 1658 463
rect 1658 427 1667 463
rect 1692 427 1722 463
rect 1722 427 1734 463
rect 1734 427 1748 463
rect 1773 427 1786 463
rect 1786 427 1798 463
rect 1798 427 1829 463
rect 1854 427 1862 463
rect 1862 427 1910 463
rect 1038 411 1094 427
rect 1120 411 1176 427
rect 1202 411 1258 427
rect 1284 411 1340 427
rect 1366 411 1422 427
rect 1448 411 1504 427
rect 1530 411 1586 427
rect 1611 411 1667 427
rect 1692 411 1748 427
rect 1773 411 1829 427
rect 1854 411 1910 427
rect 1038 407 1079 411
rect 1079 407 1092 411
rect 1092 407 1094 411
rect 1120 407 1144 411
rect 1144 407 1157 411
rect 1157 407 1176 411
rect 1202 407 1209 411
rect 1209 407 1222 411
rect 1222 407 1258 411
rect 1284 407 1286 411
rect 1286 407 1338 411
rect 1338 407 1340 411
rect 1366 407 1402 411
rect 1402 407 1414 411
rect 1414 407 1422 411
rect 1448 407 1466 411
rect 1466 407 1478 411
rect 1478 407 1504 411
rect 1530 407 1542 411
rect 1542 407 1586 411
rect 1038 359 1079 379
rect 1079 359 1092 379
rect 1092 359 1094 379
rect 1120 359 1144 379
rect 1144 359 1157 379
rect 1157 359 1176 379
rect 1202 359 1209 379
rect 1209 359 1222 379
rect 1222 359 1258 379
rect 1284 359 1286 379
rect 1286 359 1338 379
rect 1338 359 1340 379
rect 1366 359 1402 379
rect 1402 359 1414 379
rect 1414 359 1422 379
rect 1448 359 1466 379
rect 1466 359 1478 379
rect 1478 359 1504 379
rect 1530 359 1542 379
rect 1542 359 1586 379
rect 1611 407 1658 411
rect 1658 407 1667 411
rect 1692 407 1722 411
rect 1722 407 1734 411
rect 1734 407 1748 411
rect 1773 407 1786 411
rect 1786 407 1798 411
rect 1798 407 1829 411
rect 1854 407 1862 411
rect 1862 407 1910 411
rect 1611 359 1658 379
rect 1658 359 1667 379
rect 1692 359 1722 379
rect 1722 359 1734 379
rect 1734 359 1748 379
rect 1773 359 1786 379
rect 1786 359 1798 379
rect 1798 359 1829 379
rect 1854 359 1862 379
rect 1862 359 1910 379
rect 1038 343 1094 359
rect 1120 343 1176 359
rect 1202 343 1258 359
rect 1284 343 1340 359
rect 1366 343 1422 359
rect 1448 343 1504 359
rect 1530 343 1586 359
rect 1611 343 1667 359
rect 1692 343 1748 359
rect 1773 343 1829 359
rect 1854 343 1910 359
rect 1038 323 1079 343
rect 1079 323 1092 343
rect 1092 323 1094 343
rect 1120 323 1144 343
rect 1144 323 1157 343
rect 1157 323 1176 343
rect 1202 323 1209 343
rect 1209 323 1222 343
rect 1222 323 1258 343
rect 1284 323 1286 343
rect 1286 323 1338 343
rect 1338 323 1340 343
rect 1366 323 1402 343
rect 1402 323 1414 343
rect 1414 323 1422 343
rect 1448 323 1466 343
rect 1466 323 1478 343
rect 1478 323 1504 343
rect 1530 323 1542 343
rect 1542 323 1586 343
rect 1038 291 1079 295
rect 1079 291 1092 295
rect 1092 291 1094 295
rect 1120 291 1144 295
rect 1144 291 1157 295
rect 1157 291 1176 295
rect 1202 291 1209 295
rect 1209 291 1222 295
rect 1222 291 1258 295
rect 1284 291 1286 295
rect 1286 291 1338 295
rect 1338 291 1340 295
rect 1366 291 1402 295
rect 1402 291 1414 295
rect 1414 291 1422 295
rect 1448 291 1466 295
rect 1466 291 1478 295
rect 1478 291 1504 295
rect 1530 291 1542 295
rect 1542 291 1586 295
rect 1611 323 1658 343
rect 1658 323 1667 343
rect 1692 323 1722 343
rect 1722 323 1734 343
rect 1734 323 1748 343
rect 1773 323 1786 343
rect 1786 323 1798 343
rect 1798 323 1829 343
rect 1854 323 1862 343
rect 1862 323 1910 343
rect 1611 291 1658 295
rect 1658 291 1667 295
rect 1692 291 1722 295
rect 1722 291 1734 295
rect 1734 291 1748 295
rect 1773 291 1786 295
rect 1786 291 1798 295
rect 1798 291 1829 295
rect 1854 291 1862 295
rect 1862 291 1910 295
rect 1038 275 1094 291
rect 1120 275 1176 291
rect 1202 275 1258 291
rect 1284 275 1340 291
rect 1366 275 1422 291
rect 1448 275 1504 291
rect 1530 275 1586 291
rect 1611 275 1667 291
rect 1692 275 1748 291
rect 1773 275 1829 291
rect 1854 275 1910 291
rect 1038 239 1079 275
rect 1079 239 1092 275
rect 1092 239 1094 275
rect 1120 239 1144 275
rect 1144 239 1157 275
rect 1157 239 1176 275
rect 1202 239 1209 275
rect 1209 239 1222 275
rect 1222 239 1258 275
rect 1284 239 1286 275
rect 1286 239 1338 275
rect 1338 239 1340 275
rect 1366 239 1402 275
rect 1402 239 1414 275
rect 1414 239 1422 275
rect 1448 239 1466 275
rect 1466 239 1478 275
rect 1478 239 1504 275
rect 1530 239 1542 275
rect 1542 239 1586 275
rect 1611 239 1658 275
rect 1658 239 1667 275
rect 1692 239 1722 275
rect 1722 239 1734 275
rect 1734 239 1748 275
rect 1773 239 1786 275
rect 1786 239 1798 275
rect 1798 239 1829 275
rect 1854 239 1862 275
rect 1862 239 1910 275
rect 1038 207 1094 211
rect 1120 207 1176 211
rect 1202 207 1258 211
rect 1284 207 1340 211
rect 1366 207 1422 211
rect 1448 207 1504 211
rect 1530 207 1586 211
rect 1611 207 1667 211
rect 1692 207 1748 211
rect 1773 207 1829 211
rect 1854 207 1910 211
rect 1038 155 1079 207
rect 1079 155 1092 207
rect 1092 155 1094 207
rect 1120 155 1144 207
rect 1144 155 1157 207
rect 1157 155 1176 207
rect 1202 155 1209 207
rect 1209 155 1222 207
rect 1222 155 1258 207
rect 1284 155 1286 207
rect 1286 155 1338 207
rect 1338 155 1340 207
rect 1366 155 1402 207
rect 1402 155 1414 207
rect 1414 155 1422 207
rect 1448 155 1466 207
rect 1466 155 1478 207
rect 1478 155 1504 207
rect 1530 155 1542 207
rect 1542 155 1586 207
rect 1611 155 1658 207
rect 1658 155 1667 207
rect 1692 155 1722 207
rect 1722 155 1734 207
rect 1734 155 1748 207
rect 1773 155 1786 207
rect 1786 155 1798 207
rect 1798 155 1829 207
rect 1854 155 1862 207
rect 1862 155 1910 207
rect 651 -211 707 -155
rect 770 -211 826 -155
rect 888 -211 944 -155
rect 651 -281 673 -239
rect 673 -281 707 -239
rect 770 -281 799 -239
rect 799 -281 821 -239
rect 821 -281 826 -239
rect 888 -281 895 -239
rect 895 -281 944 -239
rect 651 -295 707 -281
rect 770 -295 826 -281
rect 888 -295 944 -281
rect 5203 1319 5251 1371
rect 5251 1319 5259 1371
rect 5295 1319 5315 1371
rect 5315 1319 5327 1371
rect 5327 1319 5351 1371
rect 5387 1319 5392 1371
rect 5392 1319 5443 1371
rect 5479 1319 5509 1371
rect 5509 1319 5522 1371
rect 5522 1319 5535 1371
rect 5572 1319 5574 1371
rect 5574 1319 5587 1371
rect 5587 1319 5628 1371
rect 5203 1315 5259 1319
rect 5295 1315 5351 1319
rect 5387 1315 5443 1319
rect 5479 1315 5535 1319
rect 5572 1315 5628 1319
rect 5203 1251 5251 1287
rect 5251 1251 5259 1287
rect 5295 1251 5315 1287
rect 5315 1251 5327 1287
rect 5327 1251 5351 1287
rect 5387 1251 5392 1287
rect 5392 1251 5443 1287
rect 5479 1251 5509 1287
rect 5509 1251 5522 1287
rect 5522 1251 5535 1287
rect 5572 1251 5574 1287
rect 5574 1251 5587 1287
rect 5587 1251 5628 1287
rect 5203 1235 5259 1251
rect 5295 1235 5351 1251
rect 5387 1235 5443 1251
rect 5479 1235 5535 1251
rect 5572 1235 5628 1251
rect 5203 1231 5251 1235
rect 5251 1231 5259 1235
rect 5295 1231 5315 1235
rect 5315 1231 5327 1235
rect 5327 1231 5351 1235
rect 5387 1231 5392 1235
rect 5392 1231 5443 1235
rect 5203 1183 5251 1203
rect 5251 1183 5259 1203
rect 5295 1183 5315 1203
rect 5315 1183 5327 1203
rect 5327 1183 5351 1203
rect 5387 1183 5392 1203
rect 5392 1183 5443 1203
rect 5479 1231 5509 1235
rect 5509 1231 5522 1235
rect 5522 1231 5535 1235
rect 5572 1231 5574 1235
rect 5574 1231 5587 1235
rect 5587 1231 5628 1235
rect 5479 1183 5509 1203
rect 5509 1183 5522 1203
rect 5522 1183 5535 1203
rect 5572 1183 5574 1203
rect 5574 1183 5587 1203
rect 5587 1183 5628 1203
rect 5203 1167 5259 1183
rect 5295 1167 5351 1183
rect 5387 1167 5443 1183
rect 5479 1167 5535 1183
rect 5572 1167 5628 1183
rect 5203 1147 5251 1167
rect 5251 1147 5259 1167
rect 5295 1147 5315 1167
rect 5315 1147 5327 1167
rect 5327 1147 5351 1167
rect 5387 1147 5392 1167
rect 5392 1147 5443 1167
rect 5203 1115 5251 1119
rect 5251 1115 5259 1119
rect 5295 1115 5315 1119
rect 5315 1115 5327 1119
rect 5327 1115 5351 1119
rect 5387 1115 5392 1119
rect 5392 1115 5443 1119
rect 5479 1147 5509 1167
rect 5509 1147 5522 1167
rect 5522 1147 5535 1167
rect 5572 1147 5574 1167
rect 5574 1147 5587 1167
rect 5587 1147 5628 1167
rect 5479 1115 5509 1119
rect 5509 1115 5522 1119
rect 5522 1115 5535 1119
rect 5572 1115 5574 1119
rect 5574 1115 5587 1119
rect 5587 1115 5628 1119
rect 5203 1099 5259 1115
rect 5295 1099 5351 1115
rect 5387 1099 5443 1115
rect 5479 1099 5535 1115
rect 5572 1099 5628 1115
rect 5203 1063 5251 1099
rect 5251 1063 5259 1099
rect 5295 1063 5315 1099
rect 5315 1063 5327 1099
rect 5327 1063 5351 1099
rect 5387 1063 5392 1099
rect 5392 1063 5443 1099
rect 5479 1063 5509 1099
rect 5509 1063 5522 1099
rect 5522 1063 5535 1099
rect 5572 1063 5574 1099
rect 5574 1063 5587 1099
rect 5587 1063 5628 1099
rect 5203 1031 5259 1035
rect 5295 1031 5351 1035
rect 5387 1031 5443 1035
rect 5479 1031 5535 1035
rect 5572 1031 5628 1035
rect 5203 979 5251 1031
rect 5251 979 5259 1031
rect 5295 979 5315 1031
rect 5315 979 5327 1031
rect 5327 979 5351 1031
rect 5387 979 5392 1031
rect 5392 979 5443 1031
rect 5479 979 5509 1031
rect 5509 979 5522 1031
rect 5522 979 5535 1031
rect 5572 979 5574 1031
rect 5574 979 5587 1031
rect 5587 979 5628 1031
rect 7522 1319 7563 1371
rect 7563 1319 7576 1371
rect 7576 1319 7578 1371
rect 7604 1319 7628 1371
rect 7628 1319 7641 1371
rect 7641 1319 7660 1371
rect 7686 1319 7693 1371
rect 7693 1319 7706 1371
rect 7706 1319 7742 1371
rect 7768 1319 7770 1371
rect 7770 1319 7822 1371
rect 7822 1319 7824 1371
rect 7850 1319 7886 1371
rect 7886 1319 7898 1371
rect 7898 1319 7906 1371
rect 7932 1319 7950 1371
rect 7950 1319 7962 1371
rect 7962 1319 7988 1371
rect 8014 1319 8026 1371
rect 8026 1319 8070 1371
rect 8095 1319 8142 1371
rect 8142 1319 8151 1371
rect 8176 1319 8206 1371
rect 8206 1319 8218 1371
rect 8218 1319 8232 1371
rect 8257 1319 8270 1371
rect 8270 1319 8282 1371
rect 8282 1319 8313 1371
rect 8338 1319 8346 1371
rect 8346 1319 8394 1371
rect 7522 1315 7578 1319
rect 7604 1315 7660 1319
rect 7686 1315 7742 1319
rect 7768 1315 7824 1319
rect 7850 1315 7906 1319
rect 7932 1315 7988 1319
rect 8014 1315 8070 1319
rect 8095 1315 8151 1319
rect 8176 1315 8232 1319
rect 8257 1315 8313 1319
rect 8338 1315 8394 1319
rect 7522 1251 7563 1287
rect 7563 1251 7576 1287
rect 7576 1251 7578 1287
rect 7604 1251 7628 1287
rect 7628 1251 7641 1287
rect 7641 1251 7660 1287
rect 7686 1251 7693 1287
rect 7693 1251 7706 1287
rect 7706 1251 7742 1287
rect 7768 1251 7770 1287
rect 7770 1251 7822 1287
rect 7822 1251 7824 1287
rect 7850 1251 7886 1287
rect 7886 1251 7898 1287
rect 7898 1251 7906 1287
rect 7932 1251 7950 1287
rect 7950 1251 7962 1287
rect 7962 1251 7988 1287
rect 8014 1251 8026 1287
rect 8026 1251 8070 1287
rect 8095 1251 8142 1287
rect 8142 1251 8151 1287
rect 8176 1251 8206 1287
rect 8206 1251 8218 1287
rect 8218 1251 8232 1287
rect 8257 1251 8270 1287
rect 8270 1251 8282 1287
rect 8282 1251 8313 1287
rect 8338 1251 8346 1287
rect 8346 1251 8394 1287
rect 7522 1235 7578 1251
rect 7604 1235 7660 1251
rect 7686 1235 7742 1251
rect 7768 1235 7824 1251
rect 7850 1235 7906 1251
rect 7932 1235 7988 1251
rect 8014 1235 8070 1251
rect 8095 1235 8151 1251
rect 8176 1235 8232 1251
rect 8257 1235 8313 1251
rect 8338 1235 8394 1251
rect 7522 1231 7563 1235
rect 7563 1231 7576 1235
rect 7576 1231 7578 1235
rect 7604 1231 7628 1235
rect 7628 1231 7641 1235
rect 7641 1231 7660 1235
rect 7686 1231 7693 1235
rect 7693 1231 7706 1235
rect 7706 1231 7742 1235
rect 7768 1231 7770 1235
rect 7770 1231 7822 1235
rect 7822 1231 7824 1235
rect 7850 1231 7886 1235
rect 7886 1231 7898 1235
rect 7898 1231 7906 1235
rect 7932 1231 7950 1235
rect 7950 1231 7962 1235
rect 7962 1231 7988 1235
rect 8014 1231 8026 1235
rect 8026 1231 8070 1235
rect 7522 1183 7563 1203
rect 7563 1183 7576 1203
rect 7576 1183 7578 1203
rect 7604 1183 7628 1203
rect 7628 1183 7641 1203
rect 7641 1183 7660 1203
rect 7686 1183 7693 1203
rect 7693 1183 7706 1203
rect 7706 1183 7742 1203
rect 7768 1183 7770 1203
rect 7770 1183 7822 1203
rect 7822 1183 7824 1203
rect 7850 1183 7886 1203
rect 7886 1183 7898 1203
rect 7898 1183 7906 1203
rect 7932 1183 7950 1203
rect 7950 1183 7962 1203
rect 7962 1183 7988 1203
rect 8014 1183 8026 1203
rect 8026 1183 8070 1203
rect 8095 1231 8142 1235
rect 8142 1231 8151 1235
rect 8176 1231 8206 1235
rect 8206 1231 8218 1235
rect 8218 1231 8232 1235
rect 8257 1231 8270 1235
rect 8270 1231 8282 1235
rect 8282 1231 8313 1235
rect 8338 1231 8346 1235
rect 8346 1231 8394 1235
rect 8095 1183 8142 1203
rect 8142 1183 8151 1203
rect 8176 1183 8206 1203
rect 8206 1183 8218 1203
rect 8218 1183 8232 1203
rect 8257 1183 8270 1203
rect 8270 1183 8282 1203
rect 8282 1183 8313 1203
rect 8338 1183 8346 1203
rect 8346 1183 8394 1203
rect 7522 1167 7578 1183
rect 7604 1167 7660 1183
rect 7686 1167 7742 1183
rect 7768 1167 7824 1183
rect 7850 1167 7906 1183
rect 7932 1167 7988 1183
rect 8014 1167 8070 1183
rect 8095 1167 8151 1183
rect 8176 1167 8232 1183
rect 8257 1167 8313 1183
rect 8338 1167 8394 1183
rect 7522 1147 7563 1167
rect 7563 1147 7576 1167
rect 7576 1147 7578 1167
rect 7604 1147 7628 1167
rect 7628 1147 7641 1167
rect 7641 1147 7660 1167
rect 7686 1147 7693 1167
rect 7693 1147 7706 1167
rect 7706 1147 7742 1167
rect 7768 1147 7770 1167
rect 7770 1147 7822 1167
rect 7822 1147 7824 1167
rect 7850 1147 7886 1167
rect 7886 1147 7898 1167
rect 7898 1147 7906 1167
rect 7932 1147 7950 1167
rect 7950 1147 7962 1167
rect 7962 1147 7988 1167
rect 8014 1147 8026 1167
rect 8026 1147 8070 1167
rect 7522 1115 7563 1119
rect 7563 1115 7576 1119
rect 7576 1115 7578 1119
rect 7604 1115 7628 1119
rect 7628 1115 7641 1119
rect 7641 1115 7660 1119
rect 7686 1115 7693 1119
rect 7693 1115 7706 1119
rect 7706 1115 7742 1119
rect 7768 1115 7770 1119
rect 7770 1115 7822 1119
rect 7822 1115 7824 1119
rect 7850 1115 7886 1119
rect 7886 1115 7898 1119
rect 7898 1115 7906 1119
rect 7932 1115 7950 1119
rect 7950 1115 7962 1119
rect 7962 1115 7988 1119
rect 8014 1115 8026 1119
rect 8026 1115 8070 1119
rect 8095 1147 8142 1167
rect 8142 1147 8151 1167
rect 8176 1147 8206 1167
rect 8206 1147 8218 1167
rect 8218 1147 8232 1167
rect 8257 1147 8270 1167
rect 8270 1147 8282 1167
rect 8282 1147 8313 1167
rect 8338 1147 8346 1167
rect 8346 1147 8394 1167
rect 8095 1115 8142 1119
rect 8142 1115 8151 1119
rect 8176 1115 8206 1119
rect 8206 1115 8218 1119
rect 8218 1115 8232 1119
rect 8257 1115 8270 1119
rect 8270 1115 8282 1119
rect 8282 1115 8313 1119
rect 8338 1115 8346 1119
rect 8346 1115 8394 1119
rect 7522 1099 7578 1115
rect 7604 1099 7660 1115
rect 7686 1099 7742 1115
rect 7768 1099 7824 1115
rect 7850 1099 7906 1115
rect 7932 1099 7988 1115
rect 8014 1099 8070 1115
rect 8095 1099 8151 1115
rect 8176 1099 8232 1115
rect 8257 1099 8313 1115
rect 8338 1099 8394 1115
rect 7522 1063 7563 1099
rect 7563 1063 7576 1099
rect 7576 1063 7578 1099
rect 7604 1063 7628 1099
rect 7628 1063 7641 1099
rect 7641 1063 7660 1099
rect 7686 1063 7693 1099
rect 7693 1063 7706 1099
rect 7706 1063 7742 1099
rect 7768 1063 7770 1099
rect 7770 1063 7822 1099
rect 7822 1063 7824 1099
rect 7850 1063 7886 1099
rect 7886 1063 7898 1099
rect 7898 1063 7906 1099
rect 7932 1063 7950 1099
rect 7950 1063 7962 1099
rect 7962 1063 7988 1099
rect 8014 1063 8026 1099
rect 8026 1063 8070 1099
rect 8095 1063 8142 1099
rect 8142 1063 8151 1099
rect 8176 1063 8206 1099
rect 8206 1063 8218 1099
rect 8218 1063 8232 1099
rect 8257 1063 8270 1099
rect 8270 1063 8282 1099
rect 8282 1063 8313 1099
rect 8338 1063 8346 1099
rect 8346 1063 8394 1099
rect 7522 1031 7578 1035
rect 7604 1031 7660 1035
rect 7686 1031 7742 1035
rect 7768 1031 7824 1035
rect 7850 1031 7906 1035
rect 7932 1031 7988 1035
rect 8014 1031 8070 1035
rect 8095 1031 8151 1035
rect 8176 1031 8232 1035
rect 8257 1031 8313 1035
rect 8338 1031 8394 1035
rect 7522 979 7563 1031
rect 7563 979 7576 1031
rect 7576 979 7578 1031
rect 7604 979 7628 1031
rect 7628 979 7641 1031
rect 7641 979 7660 1031
rect 7686 979 7693 1031
rect 7693 979 7706 1031
rect 7706 979 7742 1031
rect 7768 979 7770 1031
rect 7770 979 7822 1031
rect 7822 979 7824 1031
rect 7850 979 7886 1031
rect 7886 979 7898 1031
rect 7898 979 7906 1031
rect 7932 979 7950 1031
rect 7950 979 7962 1031
rect 7962 979 7988 1031
rect 8014 979 8026 1031
rect 8026 979 8070 1031
rect 8095 979 8142 1031
rect 8142 979 8151 1031
rect 8176 979 8206 1031
rect 8206 979 8218 1031
rect 8218 979 8232 1031
rect 8257 979 8270 1031
rect 8270 979 8282 1031
rect 8282 979 8313 1031
rect 8338 979 8346 1031
rect 8346 979 8394 1031
rect 3916 809 3965 858
rect 3965 809 3972 858
rect 3998 809 4029 858
rect 4029 809 4041 858
rect 4041 809 4054 858
rect 4080 809 4093 858
rect 4093 809 4105 858
rect 4105 809 4136 858
rect 4162 809 4169 858
rect 4169 809 4218 858
rect 4244 809 4285 858
rect 4285 809 4297 858
rect 4297 809 4300 858
rect 4326 809 4349 858
rect 4349 809 4361 858
rect 4361 809 4382 858
rect 4408 809 4413 858
rect 4413 809 4425 858
rect 4425 809 4464 858
rect 4490 809 4541 858
rect 4541 809 4546 858
rect 4573 809 4605 858
rect 4605 809 4617 858
rect 4617 809 4629 858
rect 4656 809 4669 858
rect 4669 809 4681 858
rect 4681 809 4712 858
rect 4739 809 4746 858
rect 4746 809 4795 858
rect 3916 802 3972 809
rect 3998 802 4054 809
rect 4080 802 4136 809
rect 4162 802 4218 809
rect 4244 802 4300 809
rect 4326 802 4382 809
rect 4408 802 4464 809
rect 4490 802 4546 809
rect 4573 802 4629 809
rect 4656 802 4712 809
rect 4739 802 4795 809
rect 3916 717 3972 724
rect 3998 717 4054 724
rect 4080 717 4136 724
rect 4162 717 4218 724
rect 4244 717 4300 724
rect 4326 717 4382 724
rect 4408 717 4464 724
rect 4490 717 4546 724
rect 4573 717 4629 724
rect 4656 717 4712 724
rect 4739 717 4795 724
rect 3916 668 3965 717
rect 3965 668 3972 717
rect 3998 668 4029 717
rect 4029 668 4041 717
rect 4041 668 4054 717
rect 4080 668 4093 717
rect 4093 668 4105 717
rect 4105 668 4136 717
rect 4162 668 4169 717
rect 4169 668 4218 717
rect 4244 668 4285 717
rect 4285 668 4297 717
rect 4297 668 4300 717
rect 4326 668 4349 717
rect 4349 668 4361 717
rect 4361 668 4382 717
rect 4408 668 4413 717
rect 4413 668 4425 717
rect 4425 668 4464 717
rect 4490 668 4541 717
rect 4541 668 4546 717
rect 4573 668 4605 717
rect 4605 668 4617 717
rect 4617 668 4629 717
rect 4656 668 4669 717
rect 4669 668 4681 717
rect 4681 668 4712 717
rect 4739 668 4746 717
rect 4746 668 4795 717
rect 8559 809 8608 858
rect 8608 809 8615 858
rect 8642 809 8673 858
rect 8673 809 8685 858
rect 8685 809 8698 858
rect 8725 809 8737 858
rect 8737 809 8749 858
rect 8749 809 8781 858
rect 8808 809 8813 858
rect 8813 809 8864 858
rect 8890 809 8929 858
rect 8929 809 8941 858
rect 8941 809 8946 858
rect 8972 809 8993 858
rect 8993 809 9005 858
rect 9005 809 9028 858
rect 9054 809 9057 858
rect 9057 809 9069 858
rect 9069 809 9110 858
rect 9136 809 9185 858
rect 9185 809 9192 858
rect 9218 809 9249 858
rect 9249 809 9261 858
rect 9261 809 9274 858
rect 9300 809 9313 858
rect 9313 809 9325 858
rect 9325 809 9356 858
rect 9382 809 9389 858
rect 9389 809 9438 858
rect 8559 802 8615 809
rect 8642 802 8698 809
rect 8725 802 8781 809
rect 8808 802 8864 809
rect 8890 802 8946 809
rect 8972 802 9028 809
rect 9054 802 9110 809
rect 9136 802 9192 809
rect 9218 802 9274 809
rect 9300 802 9356 809
rect 9382 802 9438 809
rect 8559 717 8615 724
rect 8642 717 8698 724
rect 8725 717 8781 724
rect 8808 717 8864 724
rect 8890 717 8946 724
rect 8972 717 9028 724
rect 9054 717 9110 724
rect 9136 717 9192 724
rect 9218 717 9274 724
rect 9300 717 9356 724
rect 9382 717 9438 724
rect 8559 668 8608 717
rect 8608 668 8615 717
rect 8642 668 8673 717
rect 8673 668 8685 717
rect 8685 668 8698 717
rect 8725 668 8737 717
rect 8737 668 8749 717
rect 8749 668 8781 717
rect 8808 668 8813 717
rect 8813 668 8864 717
rect 8890 668 8929 717
rect 8929 668 8941 717
rect 8941 668 8946 717
rect 8972 668 8993 717
rect 8993 668 9005 717
rect 9005 668 9028 717
rect 9054 668 9057 717
rect 9057 668 9069 717
rect 9069 668 9110 717
rect 9136 668 9185 717
rect 9185 668 9192 717
rect 9218 668 9249 717
rect 9249 668 9261 717
rect 9261 668 9274 717
rect 9300 668 9313 717
rect 9313 668 9325 717
rect 9325 668 9356 717
rect 9382 668 9389 717
rect 9389 668 9438 717
rect 5203 495 5251 547
rect 5251 495 5259 547
rect 5295 495 5315 547
rect 5315 495 5327 547
rect 5327 495 5351 547
rect 5387 495 5392 547
rect 5392 495 5443 547
rect 5479 495 5509 547
rect 5509 495 5522 547
rect 5522 495 5535 547
rect 5572 495 5574 547
rect 5574 495 5587 547
rect 5587 495 5628 547
rect 5203 491 5259 495
rect 5295 491 5351 495
rect 5387 491 5443 495
rect 5479 491 5535 495
rect 5572 491 5628 495
rect 5203 427 5251 463
rect 5251 427 5259 463
rect 5295 427 5315 463
rect 5315 427 5327 463
rect 5327 427 5351 463
rect 5387 427 5392 463
rect 5392 427 5443 463
rect 5479 427 5509 463
rect 5509 427 5522 463
rect 5522 427 5535 463
rect 5572 427 5574 463
rect 5574 427 5587 463
rect 5587 427 5628 463
rect 5203 411 5259 427
rect 5295 411 5351 427
rect 5387 411 5443 427
rect 5479 411 5535 427
rect 5572 411 5628 427
rect 5203 407 5251 411
rect 5251 407 5259 411
rect 5295 407 5315 411
rect 5315 407 5327 411
rect 5327 407 5351 411
rect 5387 407 5392 411
rect 5392 407 5443 411
rect 5203 359 5251 379
rect 5251 359 5259 379
rect 5295 359 5315 379
rect 5315 359 5327 379
rect 5327 359 5351 379
rect 5387 359 5392 379
rect 5392 359 5443 379
rect 5479 407 5509 411
rect 5509 407 5522 411
rect 5522 407 5535 411
rect 5572 407 5574 411
rect 5574 407 5587 411
rect 5587 407 5628 411
rect 5479 359 5509 379
rect 5509 359 5522 379
rect 5522 359 5535 379
rect 5572 359 5574 379
rect 5574 359 5587 379
rect 5587 359 5628 379
rect 5203 343 5259 359
rect 5295 343 5351 359
rect 5387 343 5443 359
rect 5479 343 5535 359
rect 5572 343 5628 359
rect 5203 323 5251 343
rect 5251 323 5259 343
rect 5295 323 5315 343
rect 5315 323 5327 343
rect 5327 323 5351 343
rect 5387 323 5392 343
rect 5392 323 5443 343
rect 5203 291 5251 295
rect 5251 291 5259 295
rect 5295 291 5315 295
rect 5315 291 5327 295
rect 5327 291 5351 295
rect 5387 291 5392 295
rect 5392 291 5443 295
rect 5479 323 5509 343
rect 5509 323 5522 343
rect 5522 323 5535 343
rect 5572 323 5574 343
rect 5574 323 5587 343
rect 5587 323 5628 343
rect 5479 291 5509 295
rect 5509 291 5522 295
rect 5522 291 5535 295
rect 5572 291 5574 295
rect 5574 291 5587 295
rect 5587 291 5628 295
rect 5203 275 5259 291
rect 5295 275 5351 291
rect 5387 275 5443 291
rect 5479 275 5535 291
rect 5572 275 5628 291
rect 5203 239 5251 275
rect 5251 239 5259 275
rect 5295 239 5315 275
rect 5315 239 5327 275
rect 5327 239 5351 275
rect 5387 239 5392 275
rect 5392 239 5443 275
rect 5479 239 5509 275
rect 5509 239 5522 275
rect 5522 239 5535 275
rect 5572 239 5574 275
rect 5574 239 5587 275
rect 5587 239 5628 275
rect 5203 207 5259 211
rect 5295 207 5351 211
rect 5387 207 5443 211
rect 5479 207 5535 211
rect 5572 207 5628 211
rect 5203 155 5251 207
rect 5251 155 5259 207
rect 5295 155 5315 207
rect 5315 155 5327 207
rect 5327 155 5351 207
rect 5387 155 5392 207
rect 5392 155 5443 207
rect 5479 155 5509 207
rect 5509 155 5522 207
rect 5522 155 5535 207
rect 5572 155 5574 207
rect 5574 155 5587 207
rect 5587 155 5628 207
rect 7522 495 7563 547
rect 7563 495 7576 547
rect 7576 495 7578 547
rect 7604 495 7628 547
rect 7628 495 7641 547
rect 7641 495 7660 547
rect 7686 495 7693 547
rect 7693 495 7706 547
rect 7706 495 7742 547
rect 7768 495 7770 547
rect 7770 495 7822 547
rect 7822 495 7824 547
rect 7850 495 7886 547
rect 7886 495 7898 547
rect 7898 495 7906 547
rect 7932 495 7950 547
rect 7950 495 7962 547
rect 7962 495 7988 547
rect 8014 495 8026 547
rect 8026 495 8070 547
rect 8095 495 8142 547
rect 8142 495 8151 547
rect 8176 495 8206 547
rect 8206 495 8218 547
rect 8218 495 8232 547
rect 8257 495 8270 547
rect 8270 495 8282 547
rect 8282 495 8313 547
rect 8338 495 8346 547
rect 8346 495 8394 547
rect 7522 491 7578 495
rect 7604 491 7660 495
rect 7686 491 7742 495
rect 7768 491 7824 495
rect 7850 491 7906 495
rect 7932 491 7988 495
rect 8014 491 8070 495
rect 8095 491 8151 495
rect 8176 491 8232 495
rect 8257 491 8313 495
rect 8338 491 8394 495
rect 7522 427 7563 463
rect 7563 427 7576 463
rect 7576 427 7578 463
rect 7604 427 7628 463
rect 7628 427 7641 463
rect 7641 427 7660 463
rect 7686 427 7693 463
rect 7693 427 7706 463
rect 7706 427 7742 463
rect 7768 427 7770 463
rect 7770 427 7822 463
rect 7822 427 7824 463
rect 7850 427 7886 463
rect 7886 427 7898 463
rect 7898 427 7906 463
rect 7932 427 7950 463
rect 7950 427 7962 463
rect 7962 427 7988 463
rect 8014 427 8026 463
rect 8026 427 8070 463
rect 8095 427 8142 463
rect 8142 427 8151 463
rect 8176 427 8206 463
rect 8206 427 8218 463
rect 8218 427 8232 463
rect 8257 427 8270 463
rect 8270 427 8282 463
rect 8282 427 8313 463
rect 8338 427 8346 463
rect 8346 427 8394 463
rect 7522 411 7578 427
rect 7604 411 7660 427
rect 7686 411 7742 427
rect 7768 411 7824 427
rect 7850 411 7906 427
rect 7932 411 7988 427
rect 8014 411 8070 427
rect 8095 411 8151 427
rect 8176 411 8232 427
rect 8257 411 8313 427
rect 8338 411 8394 427
rect 7522 407 7563 411
rect 7563 407 7576 411
rect 7576 407 7578 411
rect 7604 407 7628 411
rect 7628 407 7641 411
rect 7641 407 7660 411
rect 7686 407 7693 411
rect 7693 407 7706 411
rect 7706 407 7742 411
rect 7768 407 7770 411
rect 7770 407 7822 411
rect 7822 407 7824 411
rect 7850 407 7886 411
rect 7886 407 7898 411
rect 7898 407 7906 411
rect 7932 407 7950 411
rect 7950 407 7962 411
rect 7962 407 7988 411
rect 8014 407 8026 411
rect 8026 407 8070 411
rect 7522 359 7563 379
rect 7563 359 7576 379
rect 7576 359 7578 379
rect 7604 359 7628 379
rect 7628 359 7641 379
rect 7641 359 7660 379
rect 7686 359 7693 379
rect 7693 359 7706 379
rect 7706 359 7742 379
rect 7768 359 7770 379
rect 7770 359 7822 379
rect 7822 359 7824 379
rect 7850 359 7886 379
rect 7886 359 7898 379
rect 7898 359 7906 379
rect 7932 359 7950 379
rect 7950 359 7962 379
rect 7962 359 7988 379
rect 8014 359 8026 379
rect 8026 359 8070 379
rect 8095 407 8142 411
rect 8142 407 8151 411
rect 8176 407 8206 411
rect 8206 407 8218 411
rect 8218 407 8232 411
rect 8257 407 8270 411
rect 8270 407 8282 411
rect 8282 407 8313 411
rect 8338 407 8346 411
rect 8346 407 8394 411
rect 8095 359 8142 379
rect 8142 359 8151 379
rect 8176 359 8206 379
rect 8206 359 8218 379
rect 8218 359 8232 379
rect 8257 359 8270 379
rect 8270 359 8282 379
rect 8282 359 8313 379
rect 8338 359 8346 379
rect 8346 359 8394 379
rect 7522 343 7578 359
rect 7604 343 7660 359
rect 7686 343 7742 359
rect 7768 343 7824 359
rect 7850 343 7906 359
rect 7932 343 7988 359
rect 8014 343 8070 359
rect 8095 343 8151 359
rect 8176 343 8232 359
rect 8257 343 8313 359
rect 8338 343 8394 359
rect 7522 323 7563 343
rect 7563 323 7576 343
rect 7576 323 7578 343
rect 7604 323 7628 343
rect 7628 323 7641 343
rect 7641 323 7660 343
rect 7686 323 7693 343
rect 7693 323 7706 343
rect 7706 323 7742 343
rect 7768 323 7770 343
rect 7770 323 7822 343
rect 7822 323 7824 343
rect 7850 323 7886 343
rect 7886 323 7898 343
rect 7898 323 7906 343
rect 7932 323 7950 343
rect 7950 323 7962 343
rect 7962 323 7988 343
rect 8014 323 8026 343
rect 8026 323 8070 343
rect 7522 291 7563 295
rect 7563 291 7576 295
rect 7576 291 7578 295
rect 7604 291 7628 295
rect 7628 291 7641 295
rect 7641 291 7660 295
rect 7686 291 7693 295
rect 7693 291 7706 295
rect 7706 291 7742 295
rect 7768 291 7770 295
rect 7770 291 7822 295
rect 7822 291 7824 295
rect 7850 291 7886 295
rect 7886 291 7898 295
rect 7898 291 7906 295
rect 7932 291 7950 295
rect 7950 291 7962 295
rect 7962 291 7988 295
rect 8014 291 8026 295
rect 8026 291 8070 295
rect 8095 323 8142 343
rect 8142 323 8151 343
rect 8176 323 8206 343
rect 8206 323 8218 343
rect 8218 323 8232 343
rect 8257 323 8270 343
rect 8270 323 8282 343
rect 8282 323 8313 343
rect 8338 323 8346 343
rect 8346 323 8394 343
rect 8095 291 8142 295
rect 8142 291 8151 295
rect 8176 291 8206 295
rect 8206 291 8218 295
rect 8218 291 8232 295
rect 8257 291 8270 295
rect 8270 291 8282 295
rect 8282 291 8313 295
rect 8338 291 8346 295
rect 8346 291 8394 295
rect 7522 275 7578 291
rect 7604 275 7660 291
rect 7686 275 7742 291
rect 7768 275 7824 291
rect 7850 275 7906 291
rect 7932 275 7988 291
rect 8014 275 8070 291
rect 8095 275 8151 291
rect 8176 275 8232 291
rect 8257 275 8313 291
rect 8338 275 8394 291
rect 7522 239 7563 275
rect 7563 239 7576 275
rect 7576 239 7578 275
rect 7604 239 7628 275
rect 7628 239 7641 275
rect 7641 239 7660 275
rect 7686 239 7693 275
rect 7693 239 7706 275
rect 7706 239 7742 275
rect 7768 239 7770 275
rect 7770 239 7822 275
rect 7822 239 7824 275
rect 7850 239 7886 275
rect 7886 239 7898 275
rect 7898 239 7906 275
rect 7932 239 7950 275
rect 7950 239 7962 275
rect 7962 239 7988 275
rect 8014 239 8026 275
rect 8026 239 8070 275
rect 8095 239 8142 275
rect 8142 239 8151 275
rect 8176 239 8206 275
rect 8206 239 8218 275
rect 8218 239 8232 275
rect 8257 239 8270 275
rect 8270 239 8282 275
rect 8282 239 8313 275
rect 8338 239 8346 275
rect 8346 239 8394 275
rect 7522 207 7578 211
rect 7604 207 7660 211
rect 7686 207 7742 211
rect 7768 207 7824 211
rect 7850 207 7906 211
rect 7932 207 7988 211
rect 8014 207 8070 211
rect 8095 207 8151 211
rect 8176 207 8232 211
rect 8257 207 8313 211
rect 8338 207 8394 211
rect 7522 155 7563 207
rect 7563 155 7576 207
rect 7576 155 7578 207
rect 7604 155 7628 207
rect 7628 155 7641 207
rect 7641 155 7660 207
rect 7686 155 7693 207
rect 7693 155 7706 207
rect 7706 155 7742 207
rect 7768 155 7770 207
rect 7770 155 7822 207
rect 7822 155 7824 207
rect 7850 155 7886 207
rect 7886 155 7898 207
rect 7898 155 7906 207
rect 7932 155 7950 207
rect 7950 155 7962 207
rect 7962 155 7988 207
rect 8014 155 8026 207
rect 8026 155 8070 207
rect 8095 155 8142 207
rect 8142 155 8151 207
rect 8176 155 8206 207
rect 8206 155 8218 207
rect 8218 155 8232 207
rect 8257 155 8270 207
rect 8270 155 8282 207
rect 8282 155 8313 207
rect 8338 155 8346 207
rect 8346 155 8394 207
rect 3916 38 3972 39
rect 3998 38 4054 39
rect 4080 38 4136 39
rect 4162 38 4218 39
rect 4244 38 4300 39
rect 4326 38 4382 39
rect 4408 38 4464 39
rect 4490 38 4546 39
rect 4573 38 4629 39
rect 4656 38 4712 39
rect 4739 38 4795 39
rect 3916 -14 3965 38
rect 3965 -14 3972 38
rect 3998 -14 4030 38
rect 4030 -14 4042 38
rect 4042 -14 4054 38
rect 4080 -14 4094 38
rect 4094 -14 4106 38
rect 4106 -14 4136 38
rect 4162 -14 4170 38
rect 4170 -14 4218 38
rect 4244 -14 4286 38
rect 4286 -14 4298 38
rect 4298 -14 4300 38
rect 4326 -14 4350 38
rect 4350 -14 4362 38
rect 4362 -14 4382 38
rect 4408 -14 4414 38
rect 4414 -14 4426 38
rect 4426 -14 4464 38
rect 4490 -14 4542 38
rect 4542 -14 4546 38
rect 4573 -14 4606 38
rect 4606 -14 4618 38
rect 4618 -14 4629 38
rect 4656 -14 4670 38
rect 4670 -14 4682 38
rect 4682 -14 4712 38
rect 4739 -14 4746 38
rect 4746 -14 4795 38
rect 3916 -17 3972 -14
rect 3998 -17 4054 -14
rect 4080 -17 4136 -14
rect 4162 -17 4218 -14
rect 4244 -17 4300 -14
rect 4326 -17 4382 -14
rect 4408 -17 4464 -14
rect 4490 -17 4546 -14
rect 4573 -17 4629 -14
rect 4656 -17 4712 -14
rect 4739 -17 4795 -14
rect 3916 -106 3972 -95
rect 3998 -106 4054 -95
rect 4080 -106 4136 -95
rect 4162 -106 4218 -95
rect 4244 -106 4300 -95
rect 4326 -106 4382 -95
rect 4408 -106 4464 -95
rect 4490 -106 4546 -95
rect 4573 -106 4629 -95
rect 4656 -106 4712 -95
rect 4739 -106 4795 -95
rect 3916 -151 3965 -106
rect 3965 -151 3972 -106
rect 3998 -151 4030 -106
rect 4030 -151 4042 -106
rect 4042 -151 4054 -106
rect 4080 -151 4094 -106
rect 4094 -151 4106 -106
rect 4106 -151 4136 -106
rect 4162 -151 4170 -106
rect 4170 -151 4218 -106
rect 4244 -151 4286 -106
rect 4286 -151 4298 -106
rect 4298 -151 4300 -106
rect 4326 -151 4350 -106
rect 4350 -151 4362 -106
rect 4362 -151 4382 -106
rect 4408 -151 4414 -106
rect 4414 -151 4426 -106
rect 4426 -151 4464 -106
rect 4490 -151 4542 -106
rect 4542 -151 4546 -106
rect 4573 -151 4606 -106
rect 4606 -151 4618 -106
rect 4618 -151 4629 -106
rect 4656 -151 4670 -106
rect 4670 -151 4682 -106
rect 4682 -151 4712 -106
rect 4739 -151 4746 -106
rect 4746 -151 4795 -106
rect 8559 -14 8608 35
rect 8608 -14 8615 35
rect 8642 -14 8673 35
rect 8673 -14 8685 35
rect 8685 -14 8698 35
rect 8725 -14 8737 35
rect 8737 -14 8749 35
rect 8749 -14 8781 35
rect 8808 -14 8813 35
rect 8813 -14 8864 35
rect 8890 -14 8929 35
rect 8929 -14 8941 35
rect 8941 -14 8946 35
rect 8972 -14 8993 35
rect 8993 -14 9005 35
rect 9005 -14 9028 35
rect 9054 -14 9057 35
rect 9057 -14 9069 35
rect 9069 -14 9110 35
rect 9136 -14 9185 35
rect 9185 -14 9192 35
rect 9218 -14 9249 35
rect 9249 -14 9261 35
rect 9261 -14 9274 35
rect 9300 -14 9313 35
rect 9313 -14 9325 35
rect 9325 -14 9356 35
rect 9382 -14 9389 35
rect 9389 -14 9438 35
rect 8559 -21 8615 -14
rect 8642 -21 8698 -14
rect 8725 -21 8781 -14
rect 8808 -21 8864 -14
rect 8890 -21 8946 -14
rect 8972 -21 9028 -14
rect 9054 -21 9110 -14
rect 9136 -21 9192 -14
rect 9218 -21 9274 -14
rect 9300 -21 9356 -14
rect 9382 -21 9438 -14
rect 8559 -106 8615 -99
rect 8642 -106 8698 -99
rect 8725 -106 8781 -99
rect 8808 -106 8864 -99
rect 8890 -106 8946 -99
rect 8972 -106 9028 -99
rect 9054 -106 9110 -99
rect 9136 -106 9192 -99
rect 9218 -106 9274 -99
rect 9300 -106 9356 -99
rect 9382 -106 9438 -99
rect 6021 -211 6077 -155
rect 6103 -211 6159 -155
rect 6184 -211 6240 -155
rect 6265 -211 6321 -155
rect 6346 -211 6402 -155
rect 6021 -281 6070 -239
rect 6070 -281 6077 -239
rect 6103 -281 6137 -239
rect 6137 -281 6152 -239
rect 6152 -281 6159 -239
rect 6184 -281 6204 -239
rect 6204 -281 6219 -239
rect 6219 -281 6240 -239
rect 6265 -281 6271 -239
rect 6271 -281 6286 -239
rect 6286 -281 6321 -239
rect 6346 -281 6353 -239
rect 6353 -281 6402 -239
rect 6021 -295 6077 -281
rect 6103 -295 6159 -281
rect 6184 -295 6240 -281
rect 6265 -295 6321 -281
rect 6346 -295 6402 -281
rect 6952 -211 7008 -155
rect 7034 -211 7090 -155
rect 7115 -211 7171 -155
rect 7196 -211 7252 -155
rect 7277 -211 7333 -155
rect 8559 -155 8608 -106
rect 8608 -155 8615 -106
rect 8642 -155 8673 -106
rect 8673 -155 8685 -106
rect 8685 -155 8698 -106
rect 8725 -155 8737 -106
rect 8737 -155 8749 -106
rect 8749 -155 8781 -106
rect 8808 -155 8813 -106
rect 8813 -155 8864 -106
rect 8890 -155 8929 -106
rect 8929 -155 8941 -106
rect 8941 -155 8946 -106
rect 8972 -155 8993 -106
rect 8993 -155 9005 -106
rect 9005 -155 9028 -106
rect 9054 -155 9057 -106
rect 9057 -155 9069 -106
rect 9069 -155 9110 -106
rect 9136 -155 9185 -106
rect 9185 -155 9192 -106
rect 9218 -155 9249 -106
rect 9249 -155 9261 -106
rect 9261 -155 9274 -106
rect 9300 -155 9313 -106
rect 9313 -155 9325 -106
rect 9325 -155 9356 -106
rect 9382 -155 9389 -106
rect 9389 -155 9438 -106
rect 11444 1319 11492 1371
rect 11492 1319 11500 1371
rect 11525 1319 11556 1371
rect 11556 1319 11568 1371
rect 11568 1319 11581 1371
rect 11606 1319 11620 1371
rect 11620 1319 11632 1371
rect 11632 1319 11662 1371
rect 11687 1319 11696 1371
rect 11696 1319 11743 1371
rect 11768 1319 11812 1371
rect 11812 1319 11824 1371
rect 11850 1319 11876 1371
rect 11876 1319 11888 1371
rect 11888 1319 11906 1371
rect 11932 1319 11940 1371
rect 11940 1319 11952 1371
rect 11952 1319 11988 1371
rect 12014 1319 12016 1371
rect 12016 1319 12068 1371
rect 12068 1319 12070 1371
rect 12096 1319 12132 1371
rect 12132 1319 12145 1371
rect 12145 1319 12152 1371
rect 12178 1319 12197 1371
rect 12197 1319 12210 1371
rect 12210 1319 12234 1371
rect 12260 1319 12262 1371
rect 12262 1319 12275 1371
rect 12275 1319 12316 1371
rect 11444 1315 11500 1319
rect 11525 1315 11581 1319
rect 11606 1315 11662 1319
rect 11687 1315 11743 1319
rect 11768 1315 11824 1319
rect 11850 1315 11906 1319
rect 11932 1315 11988 1319
rect 12014 1315 12070 1319
rect 12096 1315 12152 1319
rect 12178 1315 12234 1319
rect 12260 1315 12316 1319
rect 11444 1251 11492 1287
rect 11492 1251 11500 1287
rect 11525 1251 11556 1287
rect 11556 1251 11568 1287
rect 11568 1251 11581 1287
rect 11606 1251 11620 1287
rect 11620 1251 11632 1287
rect 11632 1251 11662 1287
rect 11687 1251 11696 1287
rect 11696 1251 11743 1287
rect 11768 1251 11812 1287
rect 11812 1251 11824 1287
rect 11850 1251 11876 1287
rect 11876 1251 11888 1287
rect 11888 1251 11906 1287
rect 11932 1251 11940 1287
rect 11940 1251 11952 1287
rect 11952 1251 11988 1287
rect 12014 1251 12016 1287
rect 12016 1251 12068 1287
rect 12068 1251 12070 1287
rect 12096 1251 12132 1287
rect 12132 1251 12145 1287
rect 12145 1251 12152 1287
rect 12178 1251 12197 1287
rect 12197 1251 12210 1287
rect 12210 1251 12234 1287
rect 12260 1251 12262 1287
rect 12262 1251 12275 1287
rect 12275 1251 12316 1287
rect 11444 1235 11500 1251
rect 11525 1235 11581 1251
rect 11606 1235 11662 1251
rect 11687 1235 11743 1251
rect 11768 1235 11824 1251
rect 11850 1235 11906 1251
rect 11932 1235 11988 1251
rect 12014 1235 12070 1251
rect 12096 1235 12152 1251
rect 12178 1235 12234 1251
rect 12260 1235 12316 1251
rect 11444 1231 11492 1235
rect 11492 1231 11500 1235
rect 11525 1231 11556 1235
rect 11556 1231 11568 1235
rect 11568 1231 11581 1235
rect 11606 1231 11620 1235
rect 11620 1231 11632 1235
rect 11632 1231 11662 1235
rect 11687 1231 11696 1235
rect 11696 1231 11743 1235
rect 11444 1183 11492 1203
rect 11492 1183 11500 1203
rect 11525 1183 11556 1203
rect 11556 1183 11568 1203
rect 11568 1183 11581 1203
rect 11606 1183 11620 1203
rect 11620 1183 11632 1203
rect 11632 1183 11662 1203
rect 11687 1183 11696 1203
rect 11696 1183 11743 1203
rect 11768 1231 11812 1235
rect 11812 1231 11824 1235
rect 11850 1231 11876 1235
rect 11876 1231 11888 1235
rect 11888 1231 11906 1235
rect 11932 1231 11940 1235
rect 11940 1231 11952 1235
rect 11952 1231 11988 1235
rect 12014 1231 12016 1235
rect 12016 1231 12068 1235
rect 12068 1231 12070 1235
rect 12096 1231 12132 1235
rect 12132 1231 12145 1235
rect 12145 1231 12152 1235
rect 12178 1231 12197 1235
rect 12197 1231 12210 1235
rect 12210 1231 12234 1235
rect 12260 1231 12262 1235
rect 12262 1231 12275 1235
rect 12275 1231 12316 1235
rect 11768 1183 11812 1203
rect 11812 1183 11824 1203
rect 11850 1183 11876 1203
rect 11876 1183 11888 1203
rect 11888 1183 11906 1203
rect 11932 1183 11940 1203
rect 11940 1183 11952 1203
rect 11952 1183 11988 1203
rect 12014 1183 12016 1203
rect 12016 1183 12068 1203
rect 12068 1183 12070 1203
rect 12096 1183 12132 1203
rect 12132 1183 12145 1203
rect 12145 1183 12152 1203
rect 12178 1183 12197 1203
rect 12197 1183 12210 1203
rect 12210 1183 12234 1203
rect 12260 1183 12262 1203
rect 12262 1183 12275 1203
rect 12275 1183 12316 1203
rect 11444 1167 11500 1183
rect 11525 1167 11581 1183
rect 11606 1167 11662 1183
rect 11687 1167 11743 1183
rect 11768 1167 11824 1183
rect 11850 1167 11906 1183
rect 11932 1167 11988 1183
rect 12014 1167 12070 1183
rect 12096 1167 12152 1183
rect 12178 1167 12234 1183
rect 12260 1167 12316 1183
rect 11444 1147 11492 1167
rect 11492 1147 11500 1167
rect 11525 1147 11556 1167
rect 11556 1147 11568 1167
rect 11568 1147 11581 1167
rect 11606 1147 11620 1167
rect 11620 1147 11632 1167
rect 11632 1147 11662 1167
rect 11687 1147 11696 1167
rect 11696 1147 11743 1167
rect 11444 1115 11492 1119
rect 11492 1115 11500 1119
rect 11525 1115 11556 1119
rect 11556 1115 11568 1119
rect 11568 1115 11581 1119
rect 11606 1115 11620 1119
rect 11620 1115 11632 1119
rect 11632 1115 11662 1119
rect 11687 1115 11696 1119
rect 11696 1115 11743 1119
rect 11768 1147 11812 1167
rect 11812 1147 11824 1167
rect 11850 1147 11876 1167
rect 11876 1147 11888 1167
rect 11888 1147 11906 1167
rect 11932 1147 11940 1167
rect 11940 1147 11952 1167
rect 11952 1147 11988 1167
rect 12014 1147 12016 1167
rect 12016 1147 12068 1167
rect 12068 1147 12070 1167
rect 12096 1147 12132 1167
rect 12132 1147 12145 1167
rect 12145 1147 12152 1167
rect 12178 1147 12197 1167
rect 12197 1147 12210 1167
rect 12210 1147 12234 1167
rect 12260 1147 12262 1167
rect 12262 1147 12275 1167
rect 12275 1147 12316 1167
rect 11768 1115 11812 1119
rect 11812 1115 11824 1119
rect 11850 1115 11876 1119
rect 11876 1115 11888 1119
rect 11888 1115 11906 1119
rect 11932 1115 11940 1119
rect 11940 1115 11952 1119
rect 11952 1115 11988 1119
rect 12014 1115 12016 1119
rect 12016 1115 12068 1119
rect 12068 1115 12070 1119
rect 12096 1115 12132 1119
rect 12132 1115 12145 1119
rect 12145 1115 12152 1119
rect 12178 1115 12197 1119
rect 12197 1115 12210 1119
rect 12210 1115 12234 1119
rect 12260 1115 12262 1119
rect 12262 1115 12275 1119
rect 12275 1115 12316 1119
rect 11444 1099 11500 1115
rect 11525 1099 11581 1115
rect 11606 1099 11662 1115
rect 11687 1099 11743 1115
rect 11768 1099 11824 1115
rect 11850 1099 11906 1115
rect 11932 1099 11988 1115
rect 12014 1099 12070 1115
rect 12096 1099 12152 1115
rect 12178 1099 12234 1115
rect 12260 1099 12316 1115
rect 11444 1063 11492 1099
rect 11492 1063 11500 1099
rect 11525 1063 11556 1099
rect 11556 1063 11568 1099
rect 11568 1063 11581 1099
rect 11606 1063 11620 1099
rect 11620 1063 11632 1099
rect 11632 1063 11662 1099
rect 11687 1063 11696 1099
rect 11696 1063 11743 1099
rect 11768 1063 11812 1099
rect 11812 1063 11824 1099
rect 11850 1063 11876 1099
rect 11876 1063 11888 1099
rect 11888 1063 11906 1099
rect 11932 1063 11940 1099
rect 11940 1063 11952 1099
rect 11952 1063 11988 1099
rect 12014 1063 12016 1099
rect 12016 1063 12068 1099
rect 12068 1063 12070 1099
rect 12096 1063 12132 1099
rect 12132 1063 12145 1099
rect 12145 1063 12152 1099
rect 12178 1063 12197 1099
rect 12197 1063 12210 1099
rect 12210 1063 12234 1099
rect 12260 1063 12262 1099
rect 12262 1063 12275 1099
rect 12275 1063 12316 1099
rect 11444 1031 11500 1035
rect 11525 1031 11581 1035
rect 11606 1031 11662 1035
rect 11687 1031 11743 1035
rect 11768 1031 11824 1035
rect 11850 1031 11906 1035
rect 11932 1031 11988 1035
rect 12014 1031 12070 1035
rect 12096 1031 12152 1035
rect 12178 1031 12234 1035
rect 12260 1031 12316 1035
rect 11444 979 11492 1031
rect 11492 979 11500 1031
rect 11525 979 11556 1031
rect 11556 979 11568 1031
rect 11568 979 11581 1031
rect 11606 979 11620 1031
rect 11620 979 11632 1031
rect 11632 979 11662 1031
rect 11687 979 11696 1031
rect 11696 979 11743 1031
rect 11768 979 11812 1031
rect 11812 979 11824 1031
rect 11850 979 11876 1031
rect 11876 979 11888 1031
rect 11888 979 11906 1031
rect 11932 979 11940 1031
rect 11940 979 11952 1031
rect 11952 979 11988 1031
rect 12014 979 12016 1031
rect 12016 979 12068 1031
rect 12068 979 12070 1031
rect 12096 979 12132 1031
rect 12132 979 12145 1031
rect 12145 979 12152 1031
rect 12178 979 12197 1031
rect 12197 979 12210 1031
rect 12210 979 12234 1031
rect 12260 979 12262 1031
rect 12262 979 12275 1031
rect 12275 979 12316 1031
rect 14006 1319 14047 1371
rect 14047 1319 14060 1371
rect 14060 1319 14062 1371
rect 14088 1319 14112 1371
rect 14112 1319 14125 1371
rect 14125 1319 14144 1371
rect 14170 1319 14177 1371
rect 14177 1319 14190 1371
rect 14190 1319 14226 1371
rect 14252 1319 14254 1371
rect 14254 1319 14306 1371
rect 14306 1319 14308 1371
rect 14334 1319 14370 1371
rect 14370 1319 14382 1371
rect 14382 1319 14390 1371
rect 14416 1319 14434 1371
rect 14434 1319 14446 1371
rect 14446 1319 14472 1371
rect 14498 1319 14510 1371
rect 14510 1319 14554 1371
rect 14579 1319 14626 1371
rect 14626 1319 14635 1371
rect 14660 1319 14690 1371
rect 14690 1319 14702 1371
rect 14702 1319 14716 1371
rect 14741 1319 14754 1371
rect 14754 1319 14766 1371
rect 14766 1319 14797 1371
rect 14822 1319 14830 1371
rect 14830 1319 14878 1371
rect 14006 1315 14062 1319
rect 14088 1315 14144 1319
rect 14170 1315 14226 1319
rect 14252 1315 14308 1319
rect 14334 1315 14390 1319
rect 14416 1315 14472 1319
rect 14498 1315 14554 1319
rect 14579 1315 14635 1319
rect 14660 1315 14716 1319
rect 14741 1315 14797 1319
rect 14822 1315 14878 1319
rect 14006 1251 14047 1287
rect 14047 1251 14060 1287
rect 14060 1251 14062 1287
rect 14088 1251 14112 1287
rect 14112 1251 14125 1287
rect 14125 1251 14144 1287
rect 14170 1251 14177 1287
rect 14177 1251 14190 1287
rect 14190 1251 14226 1287
rect 14252 1251 14254 1287
rect 14254 1251 14306 1287
rect 14306 1251 14308 1287
rect 14334 1251 14370 1287
rect 14370 1251 14382 1287
rect 14382 1251 14390 1287
rect 14416 1251 14434 1287
rect 14434 1251 14446 1287
rect 14446 1251 14472 1287
rect 14498 1251 14510 1287
rect 14510 1251 14554 1287
rect 14579 1251 14626 1287
rect 14626 1251 14635 1287
rect 14660 1251 14690 1287
rect 14690 1251 14702 1287
rect 14702 1251 14716 1287
rect 14741 1251 14754 1287
rect 14754 1251 14766 1287
rect 14766 1251 14797 1287
rect 14822 1251 14830 1287
rect 14830 1251 14878 1287
rect 14006 1235 14062 1251
rect 14088 1235 14144 1251
rect 14170 1235 14226 1251
rect 14252 1235 14308 1251
rect 14334 1235 14390 1251
rect 14416 1235 14472 1251
rect 14498 1235 14554 1251
rect 14579 1235 14635 1251
rect 14660 1235 14716 1251
rect 14741 1235 14797 1251
rect 14822 1235 14878 1251
rect 14006 1231 14047 1235
rect 14047 1231 14060 1235
rect 14060 1231 14062 1235
rect 14088 1231 14112 1235
rect 14112 1231 14125 1235
rect 14125 1231 14144 1235
rect 14170 1231 14177 1235
rect 14177 1231 14190 1235
rect 14190 1231 14226 1235
rect 14252 1231 14254 1235
rect 14254 1231 14306 1235
rect 14306 1231 14308 1235
rect 14334 1231 14370 1235
rect 14370 1231 14382 1235
rect 14382 1231 14390 1235
rect 14416 1231 14434 1235
rect 14434 1231 14446 1235
rect 14446 1231 14472 1235
rect 14498 1231 14510 1235
rect 14510 1231 14554 1235
rect 14006 1183 14047 1203
rect 14047 1183 14060 1203
rect 14060 1183 14062 1203
rect 14088 1183 14112 1203
rect 14112 1183 14125 1203
rect 14125 1183 14144 1203
rect 14170 1183 14177 1203
rect 14177 1183 14190 1203
rect 14190 1183 14226 1203
rect 14252 1183 14254 1203
rect 14254 1183 14306 1203
rect 14306 1183 14308 1203
rect 14334 1183 14370 1203
rect 14370 1183 14382 1203
rect 14382 1183 14390 1203
rect 14416 1183 14434 1203
rect 14434 1183 14446 1203
rect 14446 1183 14472 1203
rect 14498 1183 14510 1203
rect 14510 1183 14554 1203
rect 14579 1231 14626 1235
rect 14626 1231 14635 1235
rect 14660 1231 14690 1235
rect 14690 1231 14702 1235
rect 14702 1231 14716 1235
rect 14741 1231 14754 1235
rect 14754 1231 14766 1235
rect 14766 1231 14797 1235
rect 14822 1231 14830 1235
rect 14830 1231 14878 1235
rect 14579 1183 14626 1203
rect 14626 1183 14635 1203
rect 14660 1183 14690 1203
rect 14690 1183 14702 1203
rect 14702 1183 14716 1203
rect 14741 1183 14754 1203
rect 14754 1183 14766 1203
rect 14766 1183 14797 1203
rect 14822 1183 14830 1203
rect 14830 1183 14878 1203
rect 14006 1167 14062 1183
rect 14088 1167 14144 1183
rect 14170 1167 14226 1183
rect 14252 1167 14308 1183
rect 14334 1167 14390 1183
rect 14416 1167 14472 1183
rect 14498 1167 14554 1183
rect 14579 1167 14635 1183
rect 14660 1167 14716 1183
rect 14741 1167 14797 1183
rect 14822 1167 14878 1183
rect 14006 1147 14047 1167
rect 14047 1147 14060 1167
rect 14060 1147 14062 1167
rect 14088 1147 14112 1167
rect 14112 1147 14125 1167
rect 14125 1147 14144 1167
rect 14170 1147 14177 1167
rect 14177 1147 14190 1167
rect 14190 1147 14226 1167
rect 14252 1147 14254 1167
rect 14254 1147 14306 1167
rect 14306 1147 14308 1167
rect 14334 1147 14370 1167
rect 14370 1147 14382 1167
rect 14382 1147 14390 1167
rect 14416 1147 14434 1167
rect 14434 1147 14446 1167
rect 14446 1147 14472 1167
rect 14498 1147 14510 1167
rect 14510 1147 14554 1167
rect 14006 1115 14047 1119
rect 14047 1115 14060 1119
rect 14060 1115 14062 1119
rect 14088 1115 14112 1119
rect 14112 1115 14125 1119
rect 14125 1115 14144 1119
rect 14170 1115 14177 1119
rect 14177 1115 14190 1119
rect 14190 1115 14226 1119
rect 14252 1115 14254 1119
rect 14254 1115 14306 1119
rect 14306 1115 14308 1119
rect 14334 1115 14370 1119
rect 14370 1115 14382 1119
rect 14382 1115 14390 1119
rect 14416 1115 14434 1119
rect 14434 1115 14446 1119
rect 14446 1115 14472 1119
rect 14498 1115 14510 1119
rect 14510 1115 14554 1119
rect 14579 1147 14626 1167
rect 14626 1147 14635 1167
rect 14660 1147 14690 1167
rect 14690 1147 14702 1167
rect 14702 1147 14716 1167
rect 14741 1147 14754 1167
rect 14754 1147 14766 1167
rect 14766 1147 14797 1167
rect 14822 1147 14830 1167
rect 14830 1147 14878 1167
rect 14579 1115 14626 1119
rect 14626 1115 14635 1119
rect 14660 1115 14690 1119
rect 14690 1115 14702 1119
rect 14702 1115 14716 1119
rect 14741 1115 14754 1119
rect 14754 1115 14766 1119
rect 14766 1115 14797 1119
rect 14822 1115 14830 1119
rect 14830 1115 14878 1119
rect 14006 1099 14062 1115
rect 14088 1099 14144 1115
rect 14170 1099 14226 1115
rect 14252 1099 14308 1115
rect 14334 1099 14390 1115
rect 14416 1099 14472 1115
rect 14498 1099 14554 1115
rect 14579 1099 14635 1115
rect 14660 1099 14716 1115
rect 14741 1099 14797 1115
rect 14822 1099 14878 1115
rect 14006 1063 14047 1099
rect 14047 1063 14060 1099
rect 14060 1063 14062 1099
rect 14088 1063 14112 1099
rect 14112 1063 14125 1099
rect 14125 1063 14144 1099
rect 14170 1063 14177 1099
rect 14177 1063 14190 1099
rect 14190 1063 14226 1099
rect 14252 1063 14254 1099
rect 14254 1063 14306 1099
rect 14306 1063 14308 1099
rect 14334 1063 14370 1099
rect 14370 1063 14382 1099
rect 14382 1063 14390 1099
rect 14416 1063 14434 1099
rect 14434 1063 14446 1099
rect 14446 1063 14472 1099
rect 14498 1063 14510 1099
rect 14510 1063 14554 1099
rect 14579 1063 14626 1099
rect 14626 1063 14635 1099
rect 14660 1063 14690 1099
rect 14690 1063 14702 1099
rect 14702 1063 14716 1099
rect 14741 1063 14754 1099
rect 14754 1063 14766 1099
rect 14766 1063 14797 1099
rect 14822 1063 14830 1099
rect 14830 1063 14878 1099
rect 14006 1031 14062 1035
rect 14088 1031 14144 1035
rect 14170 1031 14226 1035
rect 14252 1031 14308 1035
rect 14334 1031 14390 1035
rect 14416 1031 14472 1035
rect 14498 1031 14554 1035
rect 14579 1031 14635 1035
rect 14660 1031 14716 1035
rect 14741 1031 14797 1035
rect 14822 1031 14878 1035
rect 14006 979 14047 1031
rect 14047 979 14060 1031
rect 14060 979 14062 1031
rect 14088 979 14112 1031
rect 14112 979 14125 1031
rect 14125 979 14144 1031
rect 14170 979 14177 1031
rect 14177 979 14190 1031
rect 14190 979 14226 1031
rect 14252 979 14254 1031
rect 14254 979 14306 1031
rect 14306 979 14308 1031
rect 14334 979 14370 1031
rect 14370 979 14382 1031
rect 14382 979 14390 1031
rect 14416 979 14434 1031
rect 14434 979 14446 1031
rect 14446 979 14472 1031
rect 14498 979 14510 1031
rect 14510 979 14554 1031
rect 14579 979 14626 1031
rect 14626 979 14635 1031
rect 14660 979 14690 1031
rect 14690 979 14702 1031
rect 14702 979 14716 1031
rect 14741 979 14754 1031
rect 14754 979 14766 1031
rect 14766 979 14797 1031
rect 14822 979 14830 1031
rect 14830 979 14878 1031
rect 17928 1319 17976 1371
rect 17976 1319 17984 1371
rect 18009 1319 18040 1371
rect 18040 1319 18052 1371
rect 18052 1319 18065 1371
rect 18090 1319 18104 1371
rect 18104 1319 18116 1371
rect 18116 1319 18146 1371
rect 18171 1319 18180 1371
rect 18180 1319 18227 1371
rect 18252 1319 18296 1371
rect 18296 1319 18308 1371
rect 18334 1319 18360 1371
rect 18360 1319 18372 1371
rect 18372 1319 18390 1371
rect 18416 1319 18424 1371
rect 18424 1319 18436 1371
rect 18436 1319 18472 1371
rect 18498 1319 18500 1371
rect 18500 1319 18552 1371
rect 18552 1319 18554 1371
rect 18580 1319 18616 1371
rect 18616 1319 18629 1371
rect 18629 1319 18636 1371
rect 18662 1319 18681 1371
rect 18681 1319 18694 1371
rect 18694 1319 18718 1371
rect 18744 1319 18746 1371
rect 18746 1319 18759 1371
rect 18759 1319 18800 1371
rect 17928 1315 17984 1319
rect 18009 1315 18065 1319
rect 18090 1315 18146 1319
rect 18171 1315 18227 1319
rect 18252 1315 18308 1319
rect 18334 1315 18390 1319
rect 18416 1315 18472 1319
rect 18498 1315 18554 1319
rect 18580 1315 18636 1319
rect 18662 1315 18718 1319
rect 18744 1315 18800 1319
rect 17928 1251 17976 1287
rect 17976 1251 17984 1287
rect 18009 1251 18040 1287
rect 18040 1251 18052 1287
rect 18052 1251 18065 1287
rect 18090 1251 18104 1287
rect 18104 1251 18116 1287
rect 18116 1251 18146 1287
rect 18171 1251 18180 1287
rect 18180 1251 18227 1287
rect 18252 1251 18296 1287
rect 18296 1251 18308 1287
rect 18334 1251 18360 1287
rect 18360 1251 18372 1287
rect 18372 1251 18390 1287
rect 18416 1251 18424 1287
rect 18424 1251 18436 1287
rect 18436 1251 18472 1287
rect 18498 1251 18500 1287
rect 18500 1251 18552 1287
rect 18552 1251 18554 1287
rect 18580 1251 18616 1287
rect 18616 1251 18629 1287
rect 18629 1251 18636 1287
rect 18662 1251 18681 1287
rect 18681 1251 18694 1287
rect 18694 1251 18718 1287
rect 18744 1251 18746 1287
rect 18746 1251 18759 1287
rect 18759 1251 18800 1287
rect 17928 1235 17984 1251
rect 18009 1235 18065 1251
rect 18090 1235 18146 1251
rect 18171 1235 18227 1251
rect 18252 1235 18308 1251
rect 18334 1235 18390 1251
rect 18416 1235 18472 1251
rect 18498 1235 18554 1251
rect 18580 1235 18636 1251
rect 18662 1235 18718 1251
rect 18744 1235 18800 1251
rect 17928 1231 17976 1235
rect 17976 1231 17984 1235
rect 18009 1231 18040 1235
rect 18040 1231 18052 1235
rect 18052 1231 18065 1235
rect 18090 1231 18104 1235
rect 18104 1231 18116 1235
rect 18116 1231 18146 1235
rect 18171 1231 18180 1235
rect 18180 1231 18227 1235
rect 17928 1183 17976 1203
rect 17976 1183 17984 1203
rect 18009 1183 18040 1203
rect 18040 1183 18052 1203
rect 18052 1183 18065 1203
rect 18090 1183 18104 1203
rect 18104 1183 18116 1203
rect 18116 1183 18146 1203
rect 18171 1183 18180 1203
rect 18180 1183 18227 1203
rect 18252 1231 18296 1235
rect 18296 1231 18308 1235
rect 18334 1231 18360 1235
rect 18360 1231 18372 1235
rect 18372 1231 18390 1235
rect 18416 1231 18424 1235
rect 18424 1231 18436 1235
rect 18436 1231 18472 1235
rect 18498 1231 18500 1235
rect 18500 1231 18552 1235
rect 18552 1231 18554 1235
rect 18580 1231 18616 1235
rect 18616 1231 18629 1235
rect 18629 1231 18636 1235
rect 18662 1231 18681 1235
rect 18681 1231 18694 1235
rect 18694 1231 18718 1235
rect 18744 1231 18746 1235
rect 18746 1231 18759 1235
rect 18759 1231 18800 1235
rect 18252 1183 18296 1203
rect 18296 1183 18308 1203
rect 18334 1183 18360 1203
rect 18360 1183 18372 1203
rect 18372 1183 18390 1203
rect 18416 1183 18424 1203
rect 18424 1183 18436 1203
rect 18436 1183 18472 1203
rect 18498 1183 18500 1203
rect 18500 1183 18552 1203
rect 18552 1183 18554 1203
rect 18580 1183 18616 1203
rect 18616 1183 18629 1203
rect 18629 1183 18636 1203
rect 18662 1183 18681 1203
rect 18681 1183 18694 1203
rect 18694 1183 18718 1203
rect 18744 1183 18746 1203
rect 18746 1183 18759 1203
rect 18759 1183 18800 1203
rect 17928 1167 17984 1183
rect 18009 1167 18065 1183
rect 18090 1167 18146 1183
rect 18171 1167 18227 1183
rect 18252 1167 18308 1183
rect 18334 1167 18390 1183
rect 18416 1167 18472 1183
rect 18498 1167 18554 1183
rect 18580 1167 18636 1183
rect 18662 1167 18718 1183
rect 18744 1167 18800 1183
rect 17928 1147 17976 1167
rect 17976 1147 17984 1167
rect 18009 1147 18040 1167
rect 18040 1147 18052 1167
rect 18052 1147 18065 1167
rect 18090 1147 18104 1167
rect 18104 1147 18116 1167
rect 18116 1147 18146 1167
rect 18171 1147 18180 1167
rect 18180 1147 18227 1167
rect 17928 1115 17976 1119
rect 17976 1115 17984 1119
rect 18009 1115 18040 1119
rect 18040 1115 18052 1119
rect 18052 1115 18065 1119
rect 18090 1115 18104 1119
rect 18104 1115 18116 1119
rect 18116 1115 18146 1119
rect 18171 1115 18180 1119
rect 18180 1115 18227 1119
rect 18252 1147 18296 1167
rect 18296 1147 18308 1167
rect 18334 1147 18360 1167
rect 18360 1147 18372 1167
rect 18372 1147 18390 1167
rect 18416 1147 18424 1167
rect 18424 1147 18436 1167
rect 18436 1147 18472 1167
rect 18498 1147 18500 1167
rect 18500 1147 18552 1167
rect 18552 1147 18554 1167
rect 18580 1147 18616 1167
rect 18616 1147 18629 1167
rect 18629 1147 18636 1167
rect 18662 1147 18681 1167
rect 18681 1147 18694 1167
rect 18694 1147 18718 1167
rect 18744 1147 18746 1167
rect 18746 1147 18759 1167
rect 18759 1147 18800 1167
rect 18252 1115 18296 1119
rect 18296 1115 18308 1119
rect 18334 1115 18360 1119
rect 18360 1115 18372 1119
rect 18372 1115 18390 1119
rect 18416 1115 18424 1119
rect 18424 1115 18436 1119
rect 18436 1115 18472 1119
rect 18498 1115 18500 1119
rect 18500 1115 18552 1119
rect 18552 1115 18554 1119
rect 18580 1115 18616 1119
rect 18616 1115 18629 1119
rect 18629 1115 18636 1119
rect 18662 1115 18681 1119
rect 18681 1115 18694 1119
rect 18694 1115 18718 1119
rect 18744 1115 18746 1119
rect 18746 1115 18759 1119
rect 18759 1115 18800 1119
rect 17928 1099 17984 1115
rect 18009 1099 18065 1115
rect 18090 1099 18146 1115
rect 18171 1099 18227 1115
rect 18252 1099 18308 1115
rect 18334 1099 18390 1115
rect 18416 1099 18472 1115
rect 18498 1099 18554 1115
rect 18580 1099 18636 1115
rect 18662 1099 18718 1115
rect 18744 1099 18800 1115
rect 17928 1063 17976 1099
rect 17976 1063 17984 1099
rect 18009 1063 18040 1099
rect 18040 1063 18052 1099
rect 18052 1063 18065 1099
rect 18090 1063 18104 1099
rect 18104 1063 18116 1099
rect 18116 1063 18146 1099
rect 18171 1063 18180 1099
rect 18180 1063 18227 1099
rect 18252 1063 18296 1099
rect 18296 1063 18308 1099
rect 18334 1063 18360 1099
rect 18360 1063 18372 1099
rect 18372 1063 18390 1099
rect 18416 1063 18424 1099
rect 18424 1063 18436 1099
rect 18436 1063 18472 1099
rect 18498 1063 18500 1099
rect 18500 1063 18552 1099
rect 18552 1063 18554 1099
rect 18580 1063 18616 1099
rect 18616 1063 18629 1099
rect 18629 1063 18636 1099
rect 18662 1063 18681 1099
rect 18681 1063 18694 1099
rect 18694 1063 18718 1099
rect 18744 1063 18746 1099
rect 18746 1063 18759 1099
rect 18759 1063 18800 1099
rect 17928 1031 17984 1035
rect 18009 1031 18065 1035
rect 18090 1031 18146 1035
rect 18171 1031 18227 1035
rect 18252 1031 18308 1035
rect 18334 1031 18390 1035
rect 18416 1031 18472 1035
rect 18498 1031 18554 1035
rect 18580 1031 18636 1035
rect 18662 1031 18718 1035
rect 18744 1031 18800 1035
rect 17928 979 17976 1031
rect 17976 979 17984 1031
rect 18009 979 18040 1031
rect 18040 979 18052 1031
rect 18052 979 18065 1031
rect 18090 979 18104 1031
rect 18104 979 18116 1031
rect 18116 979 18146 1031
rect 18171 979 18180 1031
rect 18180 979 18227 1031
rect 18252 979 18296 1031
rect 18296 979 18308 1031
rect 18334 979 18360 1031
rect 18360 979 18372 1031
rect 18372 979 18390 1031
rect 18416 979 18424 1031
rect 18424 979 18436 1031
rect 18436 979 18472 1031
rect 18498 979 18500 1031
rect 18500 979 18552 1031
rect 18552 979 18554 1031
rect 18580 979 18616 1031
rect 18616 979 18629 1031
rect 18629 979 18636 1031
rect 18662 979 18681 1031
rect 18681 979 18694 1031
rect 18694 979 18718 1031
rect 18744 979 18746 1031
rect 18746 979 18759 1031
rect 18759 979 18800 1031
rect 10400 809 10449 858
rect 10449 809 10456 858
rect 10482 809 10513 858
rect 10513 809 10525 858
rect 10525 809 10538 858
rect 10564 809 10577 858
rect 10577 809 10589 858
rect 10589 809 10620 858
rect 10646 809 10653 858
rect 10653 809 10702 858
rect 10728 809 10769 858
rect 10769 809 10781 858
rect 10781 809 10784 858
rect 10810 809 10833 858
rect 10833 809 10845 858
rect 10845 809 10866 858
rect 10892 809 10897 858
rect 10897 809 10909 858
rect 10909 809 10948 858
rect 10974 809 11025 858
rect 11025 809 11030 858
rect 11057 809 11089 858
rect 11089 809 11101 858
rect 11101 809 11113 858
rect 11140 809 11153 858
rect 11153 809 11165 858
rect 11165 809 11196 858
rect 11223 809 11230 858
rect 11230 809 11279 858
rect 10400 802 10456 809
rect 10482 802 10538 809
rect 10564 802 10620 809
rect 10646 802 10702 809
rect 10728 802 10784 809
rect 10810 802 10866 809
rect 10892 802 10948 809
rect 10974 802 11030 809
rect 11057 802 11113 809
rect 11140 802 11196 809
rect 11223 802 11279 809
rect 10400 717 10456 724
rect 10482 717 10538 724
rect 10564 717 10620 724
rect 10646 717 10702 724
rect 10728 717 10784 724
rect 10810 717 10866 724
rect 10892 717 10948 724
rect 10974 717 11030 724
rect 11057 717 11113 724
rect 11140 717 11196 724
rect 11223 717 11279 724
rect 10400 668 10449 717
rect 10449 668 10456 717
rect 10482 668 10513 717
rect 10513 668 10525 717
rect 10525 668 10538 717
rect 10564 668 10577 717
rect 10577 668 10589 717
rect 10589 668 10620 717
rect 10646 668 10653 717
rect 10653 668 10702 717
rect 10728 668 10769 717
rect 10769 668 10781 717
rect 10781 668 10784 717
rect 10810 668 10833 717
rect 10833 668 10845 717
rect 10845 668 10866 717
rect 10892 668 10897 717
rect 10897 668 10909 717
rect 10909 668 10948 717
rect 10974 668 11025 717
rect 11025 668 11030 717
rect 11057 668 11089 717
rect 11089 668 11101 717
rect 11101 668 11113 717
rect 11140 668 11153 717
rect 11153 668 11165 717
rect 11165 668 11196 717
rect 11223 668 11230 717
rect 11230 668 11279 717
rect 15043 809 15092 858
rect 15092 809 15099 858
rect 15126 809 15157 858
rect 15157 809 15169 858
rect 15169 809 15182 858
rect 15209 809 15221 858
rect 15221 809 15233 858
rect 15233 809 15265 858
rect 15292 809 15297 858
rect 15297 809 15348 858
rect 15374 809 15413 858
rect 15413 809 15425 858
rect 15425 809 15430 858
rect 15456 809 15477 858
rect 15477 809 15489 858
rect 15489 809 15512 858
rect 15538 809 15541 858
rect 15541 809 15553 858
rect 15553 809 15594 858
rect 15620 809 15669 858
rect 15669 809 15676 858
rect 15702 809 15733 858
rect 15733 809 15745 858
rect 15745 809 15758 858
rect 15784 809 15797 858
rect 15797 809 15809 858
rect 15809 809 15840 858
rect 15866 809 15873 858
rect 15873 809 15922 858
rect 15043 802 15099 809
rect 15126 802 15182 809
rect 15209 802 15265 809
rect 15292 802 15348 809
rect 15374 802 15430 809
rect 15456 802 15512 809
rect 15538 802 15594 809
rect 15620 802 15676 809
rect 15702 802 15758 809
rect 15784 802 15840 809
rect 15866 802 15922 809
rect 15043 717 15099 724
rect 15126 717 15182 724
rect 15209 717 15265 724
rect 15292 717 15348 724
rect 15374 717 15430 724
rect 15456 717 15512 724
rect 15538 717 15594 724
rect 15620 717 15676 724
rect 15702 717 15758 724
rect 15784 717 15840 724
rect 15866 717 15922 724
rect 15043 668 15092 717
rect 15092 668 15099 717
rect 15126 668 15157 717
rect 15157 668 15169 717
rect 15169 668 15182 717
rect 15209 668 15221 717
rect 15221 668 15233 717
rect 15233 668 15265 717
rect 15292 668 15297 717
rect 15297 668 15348 717
rect 15374 668 15413 717
rect 15413 668 15425 717
rect 15425 668 15430 717
rect 15456 668 15477 717
rect 15477 668 15489 717
rect 15489 668 15512 717
rect 15538 668 15541 717
rect 15541 668 15553 717
rect 15553 668 15594 717
rect 15620 668 15669 717
rect 15669 668 15676 717
rect 15702 668 15733 717
rect 15733 668 15745 717
rect 15745 668 15758 717
rect 15784 668 15797 717
rect 15797 668 15809 717
rect 15809 668 15840 717
rect 15866 668 15873 717
rect 15873 668 15922 717
rect 16884 809 16933 858
rect 16933 809 16940 858
rect 16966 809 16997 858
rect 16997 809 17009 858
rect 17009 809 17022 858
rect 17048 809 17061 858
rect 17061 809 17073 858
rect 17073 809 17104 858
rect 17130 809 17137 858
rect 17137 809 17186 858
rect 17212 809 17253 858
rect 17253 809 17265 858
rect 17265 809 17268 858
rect 17294 809 17317 858
rect 17317 809 17329 858
rect 17329 809 17350 858
rect 17376 809 17381 858
rect 17381 809 17393 858
rect 17393 809 17432 858
rect 17458 809 17509 858
rect 17509 809 17514 858
rect 17541 809 17573 858
rect 17573 809 17585 858
rect 17585 809 17597 858
rect 17624 809 17637 858
rect 17637 809 17649 858
rect 17649 809 17680 858
rect 17707 809 17714 858
rect 17714 809 17763 858
rect 16884 802 16940 809
rect 16966 802 17022 809
rect 17048 802 17104 809
rect 17130 802 17186 809
rect 17212 802 17268 809
rect 17294 802 17350 809
rect 17376 802 17432 809
rect 17458 802 17514 809
rect 17541 802 17597 809
rect 17624 802 17680 809
rect 17707 802 17763 809
rect 16884 717 16940 724
rect 16966 717 17022 724
rect 17048 717 17104 724
rect 17130 717 17186 724
rect 17212 717 17268 724
rect 17294 717 17350 724
rect 17376 717 17432 724
rect 17458 717 17514 724
rect 17541 717 17597 724
rect 17624 717 17680 724
rect 17707 717 17763 724
rect 16884 668 16933 717
rect 16933 668 16940 717
rect 16966 668 16997 717
rect 16997 668 17009 717
rect 17009 668 17022 717
rect 17048 668 17061 717
rect 17061 668 17073 717
rect 17073 668 17104 717
rect 17130 668 17137 717
rect 17137 668 17186 717
rect 17212 668 17253 717
rect 17253 668 17265 717
rect 17265 668 17268 717
rect 17294 668 17317 717
rect 17317 668 17329 717
rect 17329 668 17350 717
rect 17376 668 17381 717
rect 17381 668 17393 717
rect 17393 668 17432 717
rect 17458 668 17509 717
rect 17509 668 17514 717
rect 17541 668 17573 717
rect 17573 668 17585 717
rect 17585 668 17597 717
rect 17624 668 17637 717
rect 17637 668 17649 717
rect 17649 668 17680 717
rect 17707 668 17714 717
rect 17714 668 17763 717
rect 11444 495 11492 547
rect 11492 495 11500 547
rect 11525 495 11556 547
rect 11556 495 11568 547
rect 11568 495 11581 547
rect 11606 495 11620 547
rect 11620 495 11632 547
rect 11632 495 11662 547
rect 11687 495 11696 547
rect 11696 495 11743 547
rect 11768 495 11812 547
rect 11812 495 11824 547
rect 11850 495 11876 547
rect 11876 495 11888 547
rect 11888 495 11906 547
rect 11932 495 11940 547
rect 11940 495 11952 547
rect 11952 495 11988 547
rect 12014 495 12016 547
rect 12016 495 12068 547
rect 12068 495 12070 547
rect 12096 495 12132 547
rect 12132 495 12145 547
rect 12145 495 12152 547
rect 12178 495 12197 547
rect 12197 495 12210 547
rect 12210 495 12234 547
rect 12260 495 12262 547
rect 12262 495 12275 547
rect 12275 495 12316 547
rect 11444 491 11500 495
rect 11525 491 11581 495
rect 11606 491 11662 495
rect 11687 491 11743 495
rect 11768 491 11824 495
rect 11850 491 11906 495
rect 11932 491 11988 495
rect 12014 491 12070 495
rect 12096 491 12152 495
rect 12178 491 12234 495
rect 12260 491 12316 495
rect 11444 427 11492 463
rect 11492 427 11500 463
rect 11525 427 11556 463
rect 11556 427 11568 463
rect 11568 427 11581 463
rect 11606 427 11620 463
rect 11620 427 11632 463
rect 11632 427 11662 463
rect 11687 427 11696 463
rect 11696 427 11743 463
rect 11768 427 11812 463
rect 11812 427 11824 463
rect 11850 427 11876 463
rect 11876 427 11888 463
rect 11888 427 11906 463
rect 11932 427 11940 463
rect 11940 427 11952 463
rect 11952 427 11988 463
rect 12014 427 12016 463
rect 12016 427 12068 463
rect 12068 427 12070 463
rect 12096 427 12132 463
rect 12132 427 12145 463
rect 12145 427 12152 463
rect 12178 427 12197 463
rect 12197 427 12210 463
rect 12210 427 12234 463
rect 12260 427 12262 463
rect 12262 427 12275 463
rect 12275 427 12316 463
rect 11444 411 11500 427
rect 11525 411 11581 427
rect 11606 411 11662 427
rect 11687 411 11743 427
rect 11768 411 11824 427
rect 11850 411 11906 427
rect 11932 411 11988 427
rect 12014 411 12070 427
rect 12096 411 12152 427
rect 12178 411 12234 427
rect 12260 411 12316 427
rect 11444 407 11492 411
rect 11492 407 11500 411
rect 11525 407 11556 411
rect 11556 407 11568 411
rect 11568 407 11581 411
rect 11606 407 11620 411
rect 11620 407 11632 411
rect 11632 407 11662 411
rect 11687 407 11696 411
rect 11696 407 11743 411
rect 11444 359 11492 379
rect 11492 359 11500 379
rect 11525 359 11556 379
rect 11556 359 11568 379
rect 11568 359 11581 379
rect 11606 359 11620 379
rect 11620 359 11632 379
rect 11632 359 11662 379
rect 11687 359 11696 379
rect 11696 359 11743 379
rect 11768 407 11812 411
rect 11812 407 11824 411
rect 11850 407 11876 411
rect 11876 407 11888 411
rect 11888 407 11906 411
rect 11932 407 11940 411
rect 11940 407 11952 411
rect 11952 407 11988 411
rect 12014 407 12016 411
rect 12016 407 12068 411
rect 12068 407 12070 411
rect 12096 407 12132 411
rect 12132 407 12145 411
rect 12145 407 12152 411
rect 12178 407 12197 411
rect 12197 407 12210 411
rect 12210 407 12234 411
rect 12260 407 12262 411
rect 12262 407 12275 411
rect 12275 407 12316 411
rect 11768 359 11812 379
rect 11812 359 11824 379
rect 11850 359 11876 379
rect 11876 359 11888 379
rect 11888 359 11906 379
rect 11932 359 11940 379
rect 11940 359 11952 379
rect 11952 359 11988 379
rect 12014 359 12016 379
rect 12016 359 12068 379
rect 12068 359 12070 379
rect 12096 359 12132 379
rect 12132 359 12145 379
rect 12145 359 12152 379
rect 12178 359 12197 379
rect 12197 359 12210 379
rect 12210 359 12234 379
rect 12260 359 12262 379
rect 12262 359 12275 379
rect 12275 359 12316 379
rect 11444 343 11500 359
rect 11525 343 11581 359
rect 11606 343 11662 359
rect 11687 343 11743 359
rect 11768 343 11824 359
rect 11850 343 11906 359
rect 11932 343 11988 359
rect 12014 343 12070 359
rect 12096 343 12152 359
rect 12178 343 12234 359
rect 12260 343 12316 359
rect 11444 323 11492 343
rect 11492 323 11500 343
rect 11525 323 11556 343
rect 11556 323 11568 343
rect 11568 323 11581 343
rect 11606 323 11620 343
rect 11620 323 11632 343
rect 11632 323 11662 343
rect 11687 323 11696 343
rect 11696 323 11743 343
rect 11444 291 11492 295
rect 11492 291 11500 295
rect 11525 291 11556 295
rect 11556 291 11568 295
rect 11568 291 11581 295
rect 11606 291 11620 295
rect 11620 291 11632 295
rect 11632 291 11662 295
rect 11687 291 11696 295
rect 11696 291 11743 295
rect 11768 323 11812 343
rect 11812 323 11824 343
rect 11850 323 11876 343
rect 11876 323 11888 343
rect 11888 323 11906 343
rect 11932 323 11940 343
rect 11940 323 11952 343
rect 11952 323 11988 343
rect 12014 323 12016 343
rect 12016 323 12068 343
rect 12068 323 12070 343
rect 12096 323 12132 343
rect 12132 323 12145 343
rect 12145 323 12152 343
rect 12178 323 12197 343
rect 12197 323 12210 343
rect 12210 323 12234 343
rect 12260 323 12262 343
rect 12262 323 12275 343
rect 12275 323 12316 343
rect 11768 291 11812 295
rect 11812 291 11824 295
rect 11850 291 11876 295
rect 11876 291 11888 295
rect 11888 291 11906 295
rect 11932 291 11940 295
rect 11940 291 11952 295
rect 11952 291 11988 295
rect 12014 291 12016 295
rect 12016 291 12068 295
rect 12068 291 12070 295
rect 12096 291 12132 295
rect 12132 291 12145 295
rect 12145 291 12152 295
rect 12178 291 12197 295
rect 12197 291 12210 295
rect 12210 291 12234 295
rect 12260 291 12262 295
rect 12262 291 12275 295
rect 12275 291 12316 295
rect 11444 275 11500 291
rect 11525 275 11581 291
rect 11606 275 11662 291
rect 11687 275 11743 291
rect 11768 275 11824 291
rect 11850 275 11906 291
rect 11932 275 11988 291
rect 12014 275 12070 291
rect 12096 275 12152 291
rect 12178 275 12234 291
rect 12260 275 12316 291
rect 11444 239 11492 275
rect 11492 239 11500 275
rect 11525 239 11556 275
rect 11556 239 11568 275
rect 11568 239 11581 275
rect 11606 239 11620 275
rect 11620 239 11632 275
rect 11632 239 11662 275
rect 11687 239 11696 275
rect 11696 239 11743 275
rect 11768 239 11812 275
rect 11812 239 11824 275
rect 11850 239 11876 275
rect 11876 239 11888 275
rect 11888 239 11906 275
rect 11932 239 11940 275
rect 11940 239 11952 275
rect 11952 239 11988 275
rect 12014 239 12016 275
rect 12016 239 12068 275
rect 12068 239 12070 275
rect 12096 239 12132 275
rect 12132 239 12145 275
rect 12145 239 12152 275
rect 12178 239 12197 275
rect 12197 239 12210 275
rect 12210 239 12234 275
rect 12260 239 12262 275
rect 12262 239 12275 275
rect 12275 239 12316 275
rect 11444 207 11500 211
rect 11525 207 11581 211
rect 11606 207 11662 211
rect 11687 207 11743 211
rect 11768 207 11824 211
rect 11850 207 11906 211
rect 11932 207 11988 211
rect 12014 207 12070 211
rect 12096 207 12152 211
rect 12178 207 12234 211
rect 12260 207 12316 211
rect 11444 155 11492 207
rect 11492 155 11500 207
rect 11525 155 11556 207
rect 11556 155 11568 207
rect 11568 155 11581 207
rect 11606 155 11620 207
rect 11620 155 11632 207
rect 11632 155 11662 207
rect 11687 155 11696 207
rect 11696 155 11743 207
rect 11768 155 11812 207
rect 11812 155 11824 207
rect 11850 155 11876 207
rect 11876 155 11888 207
rect 11888 155 11906 207
rect 11932 155 11940 207
rect 11940 155 11952 207
rect 11952 155 11988 207
rect 12014 155 12016 207
rect 12016 155 12068 207
rect 12068 155 12070 207
rect 12096 155 12132 207
rect 12132 155 12145 207
rect 12145 155 12152 207
rect 12178 155 12197 207
rect 12197 155 12210 207
rect 12210 155 12234 207
rect 12260 155 12262 207
rect 12262 155 12275 207
rect 12275 155 12316 207
rect 14006 495 14047 547
rect 14047 495 14060 547
rect 14060 495 14062 547
rect 14088 495 14112 547
rect 14112 495 14125 547
rect 14125 495 14144 547
rect 14170 495 14177 547
rect 14177 495 14190 547
rect 14190 495 14226 547
rect 14252 495 14254 547
rect 14254 495 14306 547
rect 14306 495 14308 547
rect 14334 495 14370 547
rect 14370 495 14382 547
rect 14382 495 14390 547
rect 14416 495 14434 547
rect 14434 495 14446 547
rect 14446 495 14472 547
rect 14498 495 14510 547
rect 14510 495 14554 547
rect 14579 495 14626 547
rect 14626 495 14635 547
rect 14660 495 14690 547
rect 14690 495 14702 547
rect 14702 495 14716 547
rect 14741 495 14754 547
rect 14754 495 14766 547
rect 14766 495 14797 547
rect 14822 495 14830 547
rect 14830 495 14878 547
rect 14006 491 14062 495
rect 14088 491 14144 495
rect 14170 491 14226 495
rect 14252 491 14308 495
rect 14334 491 14390 495
rect 14416 491 14472 495
rect 14498 491 14554 495
rect 14579 491 14635 495
rect 14660 491 14716 495
rect 14741 491 14797 495
rect 14822 491 14878 495
rect 14006 427 14047 463
rect 14047 427 14060 463
rect 14060 427 14062 463
rect 14088 427 14112 463
rect 14112 427 14125 463
rect 14125 427 14144 463
rect 14170 427 14177 463
rect 14177 427 14190 463
rect 14190 427 14226 463
rect 14252 427 14254 463
rect 14254 427 14306 463
rect 14306 427 14308 463
rect 14334 427 14370 463
rect 14370 427 14382 463
rect 14382 427 14390 463
rect 14416 427 14434 463
rect 14434 427 14446 463
rect 14446 427 14472 463
rect 14498 427 14510 463
rect 14510 427 14554 463
rect 14579 427 14626 463
rect 14626 427 14635 463
rect 14660 427 14690 463
rect 14690 427 14702 463
rect 14702 427 14716 463
rect 14741 427 14754 463
rect 14754 427 14766 463
rect 14766 427 14797 463
rect 14822 427 14830 463
rect 14830 427 14878 463
rect 14006 411 14062 427
rect 14088 411 14144 427
rect 14170 411 14226 427
rect 14252 411 14308 427
rect 14334 411 14390 427
rect 14416 411 14472 427
rect 14498 411 14554 427
rect 14579 411 14635 427
rect 14660 411 14716 427
rect 14741 411 14797 427
rect 14822 411 14878 427
rect 14006 407 14047 411
rect 14047 407 14060 411
rect 14060 407 14062 411
rect 14088 407 14112 411
rect 14112 407 14125 411
rect 14125 407 14144 411
rect 14170 407 14177 411
rect 14177 407 14190 411
rect 14190 407 14226 411
rect 14252 407 14254 411
rect 14254 407 14306 411
rect 14306 407 14308 411
rect 14334 407 14370 411
rect 14370 407 14382 411
rect 14382 407 14390 411
rect 14416 407 14434 411
rect 14434 407 14446 411
rect 14446 407 14472 411
rect 14498 407 14510 411
rect 14510 407 14554 411
rect 14006 359 14047 379
rect 14047 359 14060 379
rect 14060 359 14062 379
rect 14088 359 14112 379
rect 14112 359 14125 379
rect 14125 359 14144 379
rect 14170 359 14177 379
rect 14177 359 14190 379
rect 14190 359 14226 379
rect 14252 359 14254 379
rect 14254 359 14306 379
rect 14306 359 14308 379
rect 14334 359 14370 379
rect 14370 359 14382 379
rect 14382 359 14390 379
rect 14416 359 14434 379
rect 14434 359 14446 379
rect 14446 359 14472 379
rect 14498 359 14510 379
rect 14510 359 14554 379
rect 14579 407 14626 411
rect 14626 407 14635 411
rect 14660 407 14690 411
rect 14690 407 14702 411
rect 14702 407 14716 411
rect 14741 407 14754 411
rect 14754 407 14766 411
rect 14766 407 14797 411
rect 14822 407 14830 411
rect 14830 407 14878 411
rect 14579 359 14626 379
rect 14626 359 14635 379
rect 14660 359 14690 379
rect 14690 359 14702 379
rect 14702 359 14716 379
rect 14741 359 14754 379
rect 14754 359 14766 379
rect 14766 359 14797 379
rect 14822 359 14830 379
rect 14830 359 14878 379
rect 14006 343 14062 359
rect 14088 343 14144 359
rect 14170 343 14226 359
rect 14252 343 14308 359
rect 14334 343 14390 359
rect 14416 343 14472 359
rect 14498 343 14554 359
rect 14579 343 14635 359
rect 14660 343 14716 359
rect 14741 343 14797 359
rect 14822 343 14878 359
rect 14006 323 14047 343
rect 14047 323 14060 343
rect 14060 323 14062 343
rect 14088 323 14112 343
rect 14112 323 14125 343
rect 14125 323 14144 343
rect 14170 323 14177 343
rect 14177 323 14190 343
rect 14190 323 14226 343
rect 14252 323 14254 343
rect 14254 323 14306 343
rect 14306 323 14308 343
rect 14334 323 14370 343
rect 14370 323 14382 343
rect 14382 323 14390 343
rect 14416 323 14434 343
rect 14434 323 14446 343
rect 14446 323 14472 343
rect 14498 323 14510 343
rect 14510 323 14554 343
rect 14006 291 14047 295
rect 14047 291 14060 295
rect 14060 291 14062 295
rect 14088 291 14112 295
rect 14112 291 14125 295
rect 14125 291 14144 295
rect 14170 291 14177 295
rect 14177 291 14190 295
rect 14190 291 14226 295
rect 14252 291 14254 295
rect 14254 291 14306 295
rect 14306 291 14308 295
rect 14334 291 14370 295
rect 14370 291 14382 295
rect 14382 291 14390 295
rect 14416 291 14434 295
rect 14434 291 14446 295
rect 14446 291 14472 295
rect 14498 291 14510 295
rect 14510 291 14554 295
rect 14579 323 14626 343
rect 14626 323 14635 343
rect 14660 323 14690 343
rect 14690 323 14702 343
rect 14702 323 14716 343
rect 14741 323 14754 343
rect 14754 323 14766 343
rect 14766 323 14797 343
rect 14822 323 14830 343
rect 14830 323 14878 343
rect 14579 291 14626 295
rect 14626 291 14635 295
rect 14660 291 14690 295
rect 14690 291 14702 295
rect 14702 291 14716 295
rect 14741 291 14754 295
rect 14754 291 14766 295
rect 14766 291 14797 295
rect 14822 291 14830 295
rect 14830 291 14878 295
rect 14006 275 14062 291
rect 14088 275 14144 291
rect 14170 275 14226 291
rect 14252 275 14308 291
rect 14334 275 14390 291
rect 14416 275 14472 291
rect 14498 275 14554 291
rect 14579 275 14635 291
rect 14660 275 14716 291
rect 14741 275 14797 291
rect 14822 275 14878 291
rect 14006 239 14047 275
rect 14047 239 14060 275
rect 14060 239 14062 275
rect 14088 239 14112 275
rect 14112 239 14125 275
rect 14125 239 14144 275
rect 14170 239 14177 275
rect 14177 239 14190 275
rect 14190 239 14226 275
rect 14252 239 14254 275
rect 14254 239 14306 275
rect 14306 239 14308 275
rect 14334 239 14370 275
rect 14370 239 14382 275
rect 14382 239 14390 275
rect 14416 239 14434 275
rect 14434 239 14446 275
rect 14446 239 14472 275
rect 14498 239 14510 275
rect 14510 239 14554 275
rect 14579 239 14626 275
rect 14626 239 14635 275
rect 14660 239 14690 275
rect 14690 239 14702 275
rect 14702 239 14716 275
rect 14741 239 14754 275
rect 14754 239 14766 275
rect 14766 239 14797 275
rect 14822 239 14830 275
rect 14830 239 14878 275
rect 14006 207 14062 211
rect 14088 207 14144 211
rect 14170 207 14226 211
rect 14252 207 14308 211
rect 14334 207 14390 211
rect 14416 207 14472 211
rect 14498 207 14554 211
rect 14579 207 14635 211
rect 14660 207 14716 211
rect 14741 207 14797 211
rect 14822 207 14878 211
rect 14006 155 14047 207
rect 14047 155 14060 207
rect 14060 155 14062 207
rect 14088 155 14112 207
rect 14112 155 14125 207
rect 14125 155 14144 207
rect 14170 155 14177 207
rect 14177 155 14190 207
rect 14190 155 14226 207
rect 14252 155 14254 207
rect 14254 155 14306 207
rect 14306 155 14308 207
rect 14334 155 14370 207
rect 14370 155 14382 207
rect 14382 155 14390 207
rect 14416 155 14434 207
rect 14434 155 14446 207
rect 14446 155 14472 207
rect 14498 155 14510 207
rect 14510 155 14554 207
rect 14579 155 14626 207
rect 14626 155 14635 207
rect 14660 155 14690 207
rect 14690 155 14702 207
rect 14702 155 14716 207
rect 14741 155 14754 207
rect 14754 155 14766 207
rect 14766 155 14797 207
rect 14822 155 14830 207
rect 14830 155 14878 207
rect 17928 495 17976 547
rect 17976 495 17984 547
rect 18009 495 18040 547
rect 18040 495 18052 547
rect 18052 495 18065 547
rect 18090 495 18104 547
rect 18104 495 18116 547
rect 18116 495 18146 547
rect 18171 495 18180 547
rect 18180 495 18227 547
rect 18252 495 18296 547
rect 18296 495 18308 547
rect 18334 495 18360 547
rect 18360 495 18372 547
rect 18372 495 18390 547
rect 18416 495 18424 547
rect 18424 495 18436 547
rect 18436 495 18472 547
rect 18498 495 18500 547
rect 18500 495 18552 547
rect 18552 495 18554 547
rect 18580 495 18616 547
rect 18616 495 18629 547
rect 18629 495 18636 547
rect 18662 495 18681 547
rect 18681 495 18694 547
rect 18694 495 18718 547
rect 18744 495 18746 547
rect 18746 495 18759 547
rect 18759 495 18800 547
rect 17928 491 17984 495
rect 18009 491 18065 495
rect 18090 491 18146 495
rect 18171 491 18227 495
rect 18252 491 18308 495
rect 18334 491 18390 495
rect 18416 491 18472 495
rect 18498 491 18554 495
rect 18580 491 18636 495
rect 18662 491 18718 495
rect 18744 491 18800 495
rect 17928 427 17976 463
rect 17976 427 17984 463
rect 18009 427 18040 463
rect 18040 427 18052 463
rect 18052 427 18065 463
rect 18090 427 18104 463
rect 18104 427 18116 463
rect 18116 427 18146 463
rect 18171 427 18180 463
rect 18180 427 18227 463
rect 18252 427 18296 463
rect 18296 427 18308 463
rect 18334 427 18360 463
rect 18360 427 18372 463
rect 18372 427 18390 463
rect 18416 427 18424 463
rect 18424 427 18436 463
rect 18436 427 18472 463
rect 18498 427 18500 463
rect 18500 427 18552 463
rect 18552 427 18554 463
rect 18580 427 18616 463
rect 18616 427 18629 463
rect 18629 427 18636 463
rect 18662 427 18681 463
rect 18681 427 18694 463
rect 18694 427 18718 463
rect 18744 427 18746 463
rect 18746 427 18759 463
rect 18759 427 18800 463
rect 17928 411 17984 427
rect 18009 411 18065 427
rect 18090 411 18146 427
rect 18171 411 18227 427
rect 18252 411 18308 427
rect 18334 411 18390 427
rect 18416 411 18472 427
rect 18498 411 18554 427
rect 18580 411 18636 427
rect 18662 411 18718 427
rect 18744 411 18800 427
rect 17928 407 17976 411
rect 17976 407 17984 411
rect 18009 407 18040 411
rect 18040 407 18052 411
rect 18052 407 18065 411
rect 18090 407 18104 411
rect 18104 407 18116 411
rect 18116 407 18146 411
rect 18171 407 18180 411
rect 18180 407 18227 411
rect 17928 359 17976 379
rect 17976 359 17984 379
rect 18009 359 18040 379
rect 18040 359 18052 379
rect 18052 359 18065 379
rect 18090 359 18104 379
rect 18104 359 18116 379
rect 18116 359 18146 379
rect 18171 359 18180 379
rect 18180 359 18227 379
rect 18252 407 18296 411
rect 18296 407 18308 411
rect 18334 407 18360 411
rect 18360 407 18372 411
rect 18372 407 18390 411
rect 18416 407 18424 411
rect 18424 407 18436 411
rect 18436 407 18472 411
rect 18498 407 18500 411
rect 18500 407 18552 411
rect 18552 407 18554 411
rect 18580 407 18616 411
rect 18616 407 18629 411
rect 18629 407 18636 411
rect 18662 407 18681 411
rect 18681 407 18694 411
rect 18694 407 18718 411
rect 18744 407 18746 411
rect 18746 407 18759 411
rect 18759 407 18800 411
rect 18252 359 18296 379
rect 18296 359 18308 379
rect 18334 359 18360 379
rect 18360 359 18372 379
rect 18372 359 18390 379
rect 18416 359 18424 379
rect 18424 359 18436 379
rect 18436 359 18472 379
rect 18498 359 18500 379
rect 18500 359 18552 379
rect 18552 359 18554 379
rect 18580 359 18616 379
rect 18616 359 18629 379
rect 18629 359 18636 379
rect 18662 359 18681 379
rect 18681 359 18694 379
rect 18694 359 18718 379
rect 18744 359 18746 379
rect 18746 359 18759 379
rect 18759 359 18800 379
rect 17928 343 17984 359
rect 18009 343 18065 359
rect 18090 343 18146 359
rect 18171 343 18227 359
rect 18252 343 18308 359
rect 18334 343 18390 359
rect 18416 343 18472 359
rect 18498 343 18554 359
rect 18580 343 18636 359
rect 18662 343 18718 359
rect 18744 343 18800 359
rect 17928 323 17976 343
rect 17976 323 17984 343
rect 18009 323 18040 343
rect 18040 323 18052 343
rect 18052 323 18065 343
rect 18090 323 18104 343
rect 18104 323 18116 343
rect 18116 323 18146 343
rect 18171 323 18180 343
rect 18180 323 18227 343
rect 17928 291 17976 295
rect 17976 291 17984 295
rect 18009 291 18040 295
rect 18040 291 18052 295
rect 18052 291 18065 295
rect 18090 291 18104 295
rect 18104 291 18116 295
rect 18116 291 18146 295
rect 18171 291 18180 295
rect 18180 291 18227 295
rect 18252 323 18296 343
rect 18296 323 18308 343
rect 18334 323 18360 343
rect 18360 323 18372 343
rect 18372 323 18390 343
rect 18416 323 18424 343
rect 18424 323 18436 343
rect 18436 323 18472 343
rect 18498 323 18500 343
rect 18500 323 18552 343
rect 18552 323 18554 343
rect 18580 323 18616 343
rect 18616 323 18629 343
rect 18629 323 18636 343
rect 18662 323 18681 343
rect 18681 323 18694 343
rect 18694 323 18718 343
rect 18744 323 18746 343
rect 18746 323 18759 343
rect 18759 323 18800 343
rect 18252 291 18296 295
rect 18296 291 18308 295
rect 18334 291 18360 295
rect 18360 291 18372 295
rect 18372 291 18390 295
rect 18416 291 18424 295
rect 18424 291 18436 295
rect 18436 291 18472 295
rect 18498 291 18500 295
rect 18500 291 18552 295
rect 18552 291 18554 295
rect 18580 291 18616 295
rect 18616 291 18629 295
rect 18629 291 18636 295
rect 18662 291 18681 295
rect 18681 291 18694 295
rect 18694 291 18718 295
rect 18744 291 18746 295
rect 18746 291 18759 295
rect 18759 291 18800 295
rect 17928 275 17984 291
rect 18009 275 18065 291
rect 18090 275 18146 291
rect 18171 275 18227 291
rect 18252 275 18308 291
rect 18334 275 18390 291
rect 18416 275 18472 291
rect 18498 275 18554 291
rect 18580 275 18636 291
rect 18662 275 18718 291
rect 18744 275 18800 291
rect 17928 239 17976 275
rect 17976 239 17984 275
rect 18009 239 18040 275
rect 18040 239 18052 275
rect 18052 239 18065 275
rect 18090 239 18104 275
rect 18104 239 18116 275
rect 18116 239 18146 275
rect 18171 239 18180 275
rect 18180 239 18227 275
rect 18252 239 18296 275
rect 18296 239 18308 275
rect 18334 239 18360 275
rect 18360 239 18372 275
rect 18372 239 18390 275
rect 18416 239 18424 275
rect 18424 239 18436 275
rect 18436 239 18472 275
rect 18498 239 18500 275
rect 18500 239 18552 275
rect 18552 239 18554 275
rect 18580 239 18616 275
rect 18616 239 18629 275
rect 18629 239 18636 275
rect 18662 239 18681 275
rect 18681 239 18694 275
rect 18694 239 18718 275
rect 18744 239 18746 275
rect 18746 239 18759 275
rect 18759 239 18800 275
rect 17928 207 17984 211
rect 18009 207 18065 211
rect 18090 207 18146 211
rect 18171 207 18227 211
rect 18252 207 18308 211
rect 18334 207 18390 211
rect 18416 207 18472 211
rect 18498 207 18554 211
rect 18580 207 18636 211
rect 18662 207 18718 211
rect 18744 207 18800 211
rect 17928 155 17976 207
rect 17976 155 17984 207
rect 18009 155 18040 207
rect 18040 155 18052 207
rect 18052 155 18065 207
rect 18090 155 18104 207
rect 18104 155 18116 207
rect 18116 155 18146 207
rect 18171 155 18180 207
rect 18180 155 18227 207
rect 18252 155 18296 207
rect 18296 155 18308 207
rect 18334 155 18360 207
rect 18360 155 18372 207
rect 18372 155 18390 207
rect 18416 155 18424 207
rect 18424 155 18436 207
rect 18436 155 18472 207
rect 18498 155 18500 207
rect 18500 155 18552 207
rect 18552 155 18554 207
rect 18580 155 18616 207
rect 18616 155 18629 207
rect 18629 155 18636 207
rect 18662 155 18681 207
rect 18681 155 18694 207
rect 18694 155 18718 207
rect 18744 155 18746 207
rect 18746 155 18759 207
rect 18759 155 18800 207
rect 6952 -281 7001 -239
rect 7001 -281 7008 -239
rect 7034 -281 7068 -239
rect 7068 -281 7083 -239
rect 7083 -281 7090 -239
rect 7115 -281 7135 -239
rect 7135 -281 7150 -239
rect 7150 -281 7171 -239
rect 7196 -281 7202 -239
rect 7202 -281 7217 -239
rect 7217 -281 7252 -239
rect 7277 -281 7284 -239
rect 7284 -281 7333 -239
rect 6952 -295 7008 -281
rect 7034 -295 7090 -281
rect 7115 -295 7171 -281
rect 7196 -295 7252 -281
rect 7277 -295 7333 -281
rect 10400 -14 10449 35
rect 10449 -14 10456 35
rect 10482 -14 10514 35
rect 10514 -14 10526 35
rect 10526 -14 10538 35
rect 10564 -14 10578 35
rect 10578 -14 10590 35
rect 10590 -14 10620 35
rect 10646 -14 10654 35
rect 10654 -14 10702 35
rect 10728 -14 10770 35
rect 10770 -14 10782 35
rect 10782 -14 10784 35
rect 10810 -14 10834 35
rect 10834 -14 10846 35
rect 10846 -14 10866 35
rect 10892 -14 10898 35
rect 10898 -14 10910 35
rect 10910 -14 10948 35
rect 10974 -14 11026 35
rect 11026 -14 11030 35
rect 11057 -14 11090 35
rect 11090 -14 11102 35
rect 11102 -14 11113 35
rect 11140 -14 11154 35
rect 11154 -14 11166 35
rect 11166 -14 11196 35
rect 11223 -14 11230 35
rect 11230 -14 11279 35
rect 10400 -21 10456 -14
rect 10482 -21 10538 -14
rect 10564 -21 10620 -14
rect 10646 -21 10702 -14
rect 10728 -21 10784 -14
rect 10810 -21 10866 -14
rect 10892 -21 10948 -14
rect 10974 -21 11030 -14
rect 11057 -21 11113 -14
rect 11140 -21 11196 -14
rect 11223 -21 11279 -14
rect 10400 -106 10456 -99
rect 10482 -106 10538 -99
rect 10564 -106 10620 -99
rect 10646 -106 10702 -99
rect 10728 -106 10784 -99
rect 10810 -106 10866 -99
rect 10892 -106 10948 -99
rect 10974 -106 11030 -99
rect 11057 -106 11113 -99
rect 11140 -106 11196 -99
rect 11223 -106 11279 -99
rect 10400 -155 10449 -106
rect 10449 -155 10456 -106
rect 10482 -155 10514 -106
rect 10514 -155 10526 -106
rect 10526 -155 10538 -106
rect 10564 -155 10578 -106
rect 10578 -155 10590 -106
rect 10590 -155 10620 -106
rect 10646 -155 10654 -106
rect 10654 -155 10702 -106
rect 10728 -155 10770 -106
rect 10770 -155 10782 -106
rect 10782 -155 10784 -106
rect 10810 -155 10834 -106
rect 10834 -155 10846 -106
rect 10846 -155 10866 -106
rect 10892 -155 10898 -106
rect 10898 -155 10910 -106
rect 10910 -155 10948 -106
rect 10974 -155 11026 -106
rect 11026 -155 11030 -106
rect 11057 -155 11090 -106
rect 11090 -155 11102 -106
rect 11102 -155 11113 -106
rect 11140 -155 11154 -106
rect 11154 -155 11166 -106
rect 11166 -155 11196 -106
rect 11223 -155 11230 -106
rect 11230 -155 11279 -106
rect 11924 -22 11980 34
rect 12005 -22 12061 34
rect 12086 -22 12142 34
rect 12167 -22 12223 34
rect 12249 -22 12305 34
rect 12331 -22 12387 34
rect 11924 -156 11980 -100
rect 12005 -156 12061 -100
rect 12086 -156 12142 -100
rect 12167 -156 12223 -100
rect 12249 -156 12305 -100
rect 12331 -156 12387 -100
rect 15043 -15 15092 34
rect 15092 -15 15099 34
rect 15126 -15 15157 34
rect 15157 -15 15169 34
rect 15169 -15 15182 34
rect 15209 -15 15221 34
rect 15221 -15 15233 34
rect 15233 -15 15265 34
rect 15292 -15 15297 34
rect 15297 -15 15348 34
rect 15374 -15 15413 34
rect 15413 -15 15425 34
rect 15425 -15 15430 34
rect 15456 -15 15477 34
rect 15477 -15 15489 34
rect 15489 -15 15512 34
rect 15538 -15 15541 34
rect 15541 -15 15553 34
rect 15553 -15 15594 34
rect 15620 -15 15669 34
rect 15669 -15 15676 34
rect 15702 -15 15733 34
rect 15733 -15 15745 34
rect 15745 -15 15758 34
rect 15784 -15 15797 34
rect 15797 -15 15809 34
rect 15809 -15 15840 34
rect 15866 -15 15873 34
rect 15873 -15 15922 34
rect 15043 -22 15099 -15
rect 15126 -22 15182 -15
rect 15209 -22 15265 -15
rect 15292 -22 15348 -15
rect 15374 -22 15430 -15
rect 15456 -22 15512 -15
rect 15538 -22 15594 -15
rect 15620 -22 15676 -15
rect 15702 -22 15758 -15
rect 15784 -22 15840 -15
rect 15866 -22 15922 -15
rect 15043 -107 15099 -100
rect 15126 -107 15182 -100
rect 15209 -107 15265 -100
rect 15292 -107 15348 -100
rect 15374 -107 15430 -100
rect 15456 -107 15512 -100
rect 15538 -107 15594 -100
rect 15620 -107 15676 -100
rect 15702 -107 15758 -100
rect 15784 -107 15840 -100
rect 15866 -107 15922 -100
rect 12505 -211 12561 -155
rect 12587 -211 12643 -155
rect 12668 -211 12724 -155
rect 12749 -211 12805 -155
rect 12830 -211 12886 -155
rect 12505 -280 12554 -239
rect 12554 -280 12561 -239
rect 12587 -280 12621 -239
rect 12621 -280 12636 -239
rect 12636 -280 12643 -239
rect 12668 -280 12688 -239
rect 12688 -280 12703 -239
rect 12703 -280 12724 -239
rect 12749 -280 12755 -239
rect 12755 -280 12770 -239
rect 12770 -280 12805 -239
rect 12830 -280 12837 -239
rect 12837 -280 12886 -239
rect 12505 -295 12561 -280
rect 12587 -295 12643 -280
rect 12668 -295 12724 -280
rect 12749 -295 12805 -280
rect 12830 -295 12886 -280
rect 13436 -211 13492 -155
rect 13518 -211 13574 -155
rect 13599 -211 13655 -155
rect 13680 -211 13736 -155
rect 13761 -211 13817 -155
rect 15043 -156 15092 -107
rect 15092 -156 15099 -107
rect 15126 -156 15157 -107
rect 15157 -156 15169 -107
rect 15169 -156 15182 -107
rect 15209 -156 15221 -107
rect 15221 -156 15233 -107
rect 15233 -156 15265 -107
rect 15292 -156 15297 -107
rect 15297 -156 15348 -107
rect 15374 -156 15413 -107
rect 15413 -156 15425 -107
rect 15425 -156 15430 -107
rect 15456 -156 15477 -107
rect 15477 -156 15489 -107
rect 15489 -156 15512 -107
rect 15538 -156 15541 -107
rect 15541 -156 15553 -107
rect 15553 -156 15594 -107
rect 15620 -156 15669 -107
rect 15669 -156 15676 -107
rect 15702 -156 15733 -107
rect 15733 -156 15745 -107
rect 15745 -156 15758 -107
rect 15784 -156 15797 -107
rect 15797 -156 15809 -107
rect 15809 -156 15840 -107
rect 15866 -156 15873 -107
rect 15873 -156 15922 -107
rect 16884 -15 16933 34
rect 16933 -15 16940 34
rect 16967 -15 16998 34
rect 16998 -15 17010 34
rect 17010 -15 17023 34
rect 17050 -15 17062 34
rect 17062 -15 17074 34
rect 17074 -15 17106 34
rect 17133 -15 17138 34
rect 17138 -15 17189 34
rect 17215 -15 17254 34
rect 17254 -15 17266 34
rect 17266 -15 17271 34
rect 17297 -15 17318 34
rect 17318 -15 17330 34
rect 17330 -15 17353 34
rect 17379 -15 17382 34
rect 17382 -15 17394 34
rect 17394 -15 17435 34
rect 17461 -15 17510 34
rect 17510 -15 17517 34
rect 17543 -15 17574 34
rect 17574 -15 17586 34
rect 17586 -15 17599 34
rect 17625 -15 17638 34
rect 17638 -15 17650 34
rect 17650 -15 17681 34
rect 17707 -15 17714 34
rect 17714 -15 17763 34
rect 16884 -22 16940 -15
rect 16967 -22 17023 -15
rect 17050 -22 17106 -15
rect 17133 -22 17189 -15
rect 17215 -22 17271 -15
rect 17297 -22 17353 -15
rect 17379 -22 17435 -15
rect 17461 -22 17517 -15
rect 17543 -22 17599 -15
rect 17625 -22 17681 -15
rect 17707 -22 17763 -15
rect 16884 -107 16940 -100
rect 16967 -107 17023 -100
rect 17050 -107 17106 -100
rect 17133 -107 17189 -100
rect 17215 -107 17271 -100
rect 17297 -107 17353 -100
rect 17379 -107 17435 -100
rect 17461 -107 17517 -100
rect 17543 -107 17599 -100
rect 17625 -107 17681 -100
rect 17707 -107 17763 -100
rect 16884 -156 16933 -107
rect 16933 -156 16940 -107
rect 16967 -156 16998 -107
rect 16998 -156 17010 -107
rect 17010 -156 17023 -107
rect 17050 -156 17062 -107
rect 17062 -156 17074 -107
rect 17074 -156 17106 -107
rect 17133 -156 17138 -107
rect 17138 -156 17189 -107
rect 17215 -156 17254 -107
rect 17254 -156 17266 -107
rect 17266 -156 17271 -107
rect 17297 -156 17318 -107
rect 17318 -156 17330 -107
rect 17330 -156 17353 -107
rect 17379 -156 17382 -107
rect 17382 -156 17394 -107
rect 17394 -156 17435 -107
rect 17461 -156 17510 -107
rect 17510 -156 17517 -107
rect 17543 -156 17574 -107
rect 17574 -156 17586 -107
rect 17586 -156 17599 -107
rect 17625 -156 17638 -107
rect 17638 -156 17650 -107
rect 17650 -156 17681 -107
rect 17707 -156 17714 -107
rect 17714 -156 17763 -107
rect 13436 -281 13485 -239
rect 13485 -281 13492 -239
rect 13518 -281 13552 -239
rect 13552 -281 13567 -239
rect 13567 -281 13574 -239
rect 13599 -281 13619 -239
rect 13619 -281 13634 -239
rect 13634 -281 13655 -239
rect 13680 -281 13686 -239
rect 13686 -281 13701 -239
rect 13701 -281 13736 -239
rect 13761 -281 13768 -239
rect 13768 -281 13817 -239
rect 13436 -295 13492 -281
rect 13518 -295 13574 -281
rect 13599 -295 13655 -281
rect 13680 -295 13736 -281
rect 13761 -295 13817 -281
rect 19074 -211 19130 -155
rect 19154 -211 19210 -155
rect 19234 -211 19290 -155
rect 19314 -211 19370 -155
rect 19074 -281 19123 -239
rect 19123 -281 19130 -239
rect 19074 -295 19130 -281
rect 19154 -281 19155 -239
rect 19155 -281 19207 -239
rect 19207 -281 19210 -239
rect 19154 -295 19210 -281
rect 19234 -281 19238 -239
rect 19238 -281 19290 -239
rect 19234 -295 19290 -281
rect 19314 -281 19321 -239
rect 19321 -281 19370 -239
rect 19314 -295 19370 -281
rect 15048 -2810 15104 -2754
rect 15129 -2810 15185 -2754
rect 15210 -2810 15266 -2754
rect 15291 -2810 15347 -2754
rect 15372 -2810 15428 -2754
rect 15453 -2810 15509 -2754
rect 15534 -2810 15590 -2754
rect 15614 -2810 15670 -2754
rect 15694 -2810 15750 -2754
rect 15774 -2810 15830 -2754
rect 15854 -2810 15910 -2754
rect 15048 -2871 15104 -2862
rect 15129 -2871 15185 -2862
rect 15210 -2871 15266 -2862
rect 15291 -2871 15347 -2862
rect 15372 -2871 15428 -2862
rect 15453 -2871 15509 -2862
rect 15534 -2871 15590 -2862
rect 15614 -2871 15670 -2862
rect 15694 -2871 15750 -2862
rect 15774 -2871 15830 -2862
rect 15854 -2871 15910 -2862
rect 15048 -2918 15097 -2871
rect 15097 -2918 15104 -2871
rect 15129 -2918 15165 -2871
rect 15165 -2918 15181 -2871
rect 15181 -2918 15185 -2871
rect 15210 -2918 15233 -2871
rect 15233 -2918 15249 -2871
rect 15249 -2918 15266 -2871
rect 15291 -2918 15301 -2871
rect 15301 -2918 15317 -2871
rect 15317 -2918 15347 -2871
rect 15372 -2918 15385 -2871
rect 15385 -2918 15428 -2871
rect 15453 -2918 15505 -2871
rect 15505 -2918 15509 -2871
rect 15534 -2918 15573 -2871
rect 15573 -2918 15589 -2871
rect 15589 -2918 15590 -2871
rect 15614 -2918 15641 -2871
rect 15641 -2918 15657 -2871
rect 15657 -2918 15670 -2871
rect 15694 -2918 15709 -2871
rect 15709 -2918 15725 -2871
rect 15725 -2918 15750 -2871
rect 15774 -2918 15777 -2871
rect 15777 -2918 15793 -2871
rect 15793 -2918 15830 -2871
rect 15854 -2918 15861 -2871
rect 15861 -2918 15910 -2871
rect 16889 -2810 16945 -2754
rect 16970 -2810 17026 -2754
rect 17051 -2810 17107 -2754
rect 17132 -2810 17188 -2754
rect 17213 -2810 17269 -2754
rect 17294 -2810 17350 -2754
rect 17375 -2810 17431 -2754
rect 17455 -2810 17511 -2754
rect 17535 -2810 17591 -2754
rect 17615 -2810 17671 -2754
rect 17695 -2810 17751 -2754
rect 16889 -2871 16945 -2862
rect 16970 -2871 17026 -2862
rect 17051 -2871 17107 -2862
rect 17132 -2871 17188 -2862
rect 17213 -2871 17269 -2862
rect 17294 -2871 17350 -2862
rect 17375 -2871 17431 -2862
rect 17455 -2871 17511 -2862
rect 17535 -2871 17591 -2862
rect 17615 -2871 17671 -2862
rect 17695 -2871 17751 -2862
rect 16889 -2918 16938 -2871
rect 16938 -2918 16945 -2871
rect 16970 -2918 17006 -2871
rect 17006 -2918 17022 -2871
rect 17022 -2918 17026 -2871
rect 17051 -2918 17074 -2871
rect 17074 -2918 17090 -2871
rect 17090 -2918 17107 -2871
rect 17132 -2918 17142 -2871
rect 17142 -2918 17158 -2871
rect 17158 -2918 17188 -2871
rect 17213 -2918 17226 -2871
rect 17226 -2918 17269 -2871
rect 17294 -2918 17346 -2871
rect 17346 -2918 17350 -2871
rect 17375 -2918 17414 -2871
rect 17414 -2918 17430 -2871
rect 17430 -2918 17431 -2871
rect 17455 -2918 17482 -2871
rect 17482 -2918 17498 -2871
rect 17498 -2918 17511 -2871
rect 17535 -2918 17550 -2871
rect 17550 -2918 17566 -2871
rect 17566 -2918 17591 -2871
rect 17615 -2918 17618 -2871
rect 17618 -2918 17634 -2871
rect 17634 -2918 17671 -2871
rect 17695 -2918 17702 -2871
rect 17702 -2918 17751 -2871
<< metal3 >>
rect 19670 5501 19816 5754
rect 19670 5445 19675 5501
rect 19731 5445 19755 5501
rect 19811 5445 19816 5501
rect 14001 5226 14883 5258
rect 3911 5133 4393 5135
rect 3028 5128 4393 5133
rect 3028 5072 3033 5128
rect 3089 5072 3115 5128
rect 3171 5072 3197 5128
rect 3253 5072 3279 5128
rect 3335 5072 3361 5128
rect 3417 5072 3443 5128
rect 3499 5072 3525 5128
rect 3581 5072 3607 5128
rect 3663 5072 3689 5128
rect 3745 5072 3771 5128
rect 3827 5072 3853 5128
rect 3909 5072 3935 5128
rect 3991 5072 4016 5128
rect 4072 5072 4097 5128
rect 4153 5072 4178 5128
rect 4234 5072 4259 5128
rect 4315 5072 4393 5128
rect 3028 5020 4393 5072
rect 3028 4964 3033 5020
rect 3089 4964 3115 5020
rect 3171 4964 3197 5020
rect 3253 4964 3279 5020
rect 3335 4964 3361 5020
rect 3417 4964 3443 5020
rect 3499 4964 3525 5020
rect 3581 4964 3607 5020
rect 3663 4964 3689 5020
rect 3745 4964 3771 5020
rect 3827 4964 3853 5020
rect 3909 4964 3935 5020
rect 3991 4964 4016 5020
rect 4072 4964 4097 5020
rect 4153 4964 4178 5020
rect 4234 4964 4259 5020
rect 4315 4964 4393 5020
rect 3028 4959 4393 4964
rect 1033 4792 1047 4856
rect 1111 4792 1135 4856
rect 1199 4792 1223 4856
rect 1287 4792 1311 4856
rect 1375 4792 1399 4856
rect 1463 4792 1487 4856
rect 1551 4792 1575 4856
rect 1639 4792 1662 4856
rect 1726 4792 1749 4856
rect 1813 4792 1836 4856
rect 1900 4792 1915 4856
rect 1033 4764 1915 4792
rect 1033 4700 1047 4764
rect 1111 4700 1135 4764
rect 1199 4700 1223 4764
rect 1287 4700 1311 4764
rect 1375 4700 1399 4764
rect 1463 4700 1487 4764
rect 1551 4700 1575 4764
rect 1639 4700 1662 4764
rect 1726 4700 1749 4764
rect 1813 4700 1836 4764
rect 1900 4700 1915 4764
rect 1033 4672 1915 4700
rect 1033 4608 1047 4672
rect 1111 4608 1135 4672
rect 1199 4608 1223 4672
rect 1287 4608 1311 4672
rect 1375 4608 1399 4672
rect 1463 4608 1487 4672
rect 1551 4608 1575 4672
rect 1639 4608 1662 4672
rect 1726 4608 1749 4672
rect 1813 4608 1836 4672
rect 1900 4608 1915 4672
rect 1033 4580 1915 4608
rect 1033 4516 1047 4580
rect 1111 4516 1135 4580
rect 1199 4516 1223 4580
rect 1287 4516 1311 4580
rect 1375 4516 1399 4580
rect 1463 4516 1487 4580
rect 1551 4516 1575 4580
rect 1639 4516 1662 4580
rect 1726 4516 1749 4580
rect 1813 4516 1836 4580
rect 1900 4516 1915 4580
rect 1033 4488 1915 4516
rect 1033 4424 1047 4488
rect 1111 4424 1135 4488
rect 1199 4424 1223 4488
rect 1287 4424 1311 4488
rect 1375 4424 1399 4488
rect 1463 4424 1487 4488
rect 1551 4424 1575 4488
rect 1639 4424 1662 4488
rect 1726 4424 1749 4488
rect 1813 4424 1836 4488
rect 1900 4424 1915 4488
rect 1033 4396 1915 4424
rect 642 4351 953 4376
rect 642 4295 647 4351
rect 703 4295 729 4351
rect 785 4295 811 4351
rect 867 4295 892 4351
rect 948 4295 953 4351
rect 642 4267 953 4295
rect 642 4211 647 4267
rect 703 4211 729 4267
rect 785 4211 811 4267
rect 867 4211 892 4267
rect 948 4211 953 4267
rect 642 2963 953 4211
rect 642 2907 647 2963
rect 703 2907 728 2963
rect 784 2907 808 2963
rect 864 2907 888 2963
rect 944 2907 953 2963
rect 642 2879 953 2907
rect 642 2823 647 2879
rect 703 2823 728 2879
rect 784 2823 808 2879
rect 864 2823 888 2879
rect 944 2823 953 2879
rect 642 2738 953 2823
rect 642 2682 647 2738
rect 703 2682 728 2738
rect 784 2682 808 2738
rect 864 2682 888 2738
rect 944 2682 953 2738
rect 642 2614 953 2682
rect 642 2558 647 2614
rect 703 2558 728 2614
rect 784 2558 808 2614
rect 864 2558 888 2614
rect 944 2558 953 2614
rect 642 1919 953 2558
rect 642 1863 647 1919
rect 703 1863 728 1919
rect 784 1863 808 1919
rect 864 1863 888 1919
rect 944 1863 953 1919
rect 642 1795 953 1863
rect 642 1739 647 1795
rect 703 1739 728 1795
rect 784 1739 808 1795
rect 864 1739 888 1795
rect 944 1739 953 1795
rect 642 -155 953 1739
rect 642 -211 651 -155
rect 707 -211 770 -155
rect 826 -211 888 -155
rect 944 -211 953 -155
rect 642 -239 953 -211
rect 642 -295 651 -239
rect 707 -295 770 -239
rect 826 -295 888 -239
rect 944 -295 953 -239
rect 642 -1785 953 -295
rect 1033 4332 1047 4396
rect 1111 4332 1135 4396
rect 1199 4332 1223 4396
rect 1287 4332 1311 4396
rect 1375 4332 1399 4396
rect 1463 4332 1487 4396
rect 1551 4332 1575 4396
rect 1639 4332 1662 4396
rect 1726 4332 1749 4396
rect 1813 4332 1836 4396
rect 1900 4332 1915 4396
rect 1033 2437 1915 4332
rect 1033 2381 1038 2437
rect 1094 2381 1120 2437
rect 1176 2381 1202 2437
rect 1258 2381 1284 2437
rect 1340 2381 1366 2437
rect 1422 2381 1448 2437
rect 1504 2381 1530 2437
rect 1586 2381 1611 2437
rect 1667 2381 1692 2437
rect 1748 2381 1773 2437
rect 1829 2381 1854 2437
rect 1910 2381 1915 2437
rect 1033 2353 1915 2381
rect 1033 2297 1038 2353
rect 1094 2297 1120 2353
rect 1176 2297 1202 2353
rect 1258 2297 1284 2353
rect 1340 2297 1366 2353
rect 1422 2297 1448 2353
rect 1504 2297 1530 2353
rect 1586 2297 1611 2353
rect 1667 2297 1692 2353
rect 1748 2297 1773 2353
rect 1829 2297 1854 2353
rect 1910 2297 1915 2353
rect 1033 2269 1915 2297
rect 1033 2213 1038 2269
rect 1094 2213 1120 2269
rect 1176 2213 1202 2269
rect 1258 2213 1284 2269
rect 1340 2213 1366 2269
rect 1422 2213 1448 2269
rect 1504 2213 1530 2269
rect 1586 2213 1611 2269
rect 1667 2213 1692 2269
rect 1748 2213 1773 2269
rect 1829 2213 1854 2269
rect 1910 2213 1915 2269
rect 1033 2185 1915 2213
rect 1033 2129 1038 2185
rect 1094 2129 1120 2185
rect 1176 2129 1202 2185
rect 1258 2129 1284 2185
rect 1340 2129 1366 2185
rect 1422 2129 1448 2185
rect 1504 2129 1530 2185
rect 1586 2129 1611 2185
rect 1667 2129 1692 2185
rect 1748 2129 1773 2185
rect 1829 2129 1854 2185
rect 1910 2129 1915 2185
rect 1033 2101 1915 2129
rect 1033 2045 1038 2101
rect 1094 2045 1120 2101
rect 1176 2045 1202 2101
rect 1258 2045 1284 2101
rect 1340 2045 1366 2101
rect 1422 2045 1448 2101
rect 1504 2045 1530 2101
rect 1586 2045 1611 2101
rect 1667 2045 1692 2101
rect 1748 2045 1773 2101
rect 1829 2045 1854 2101
rect 1910 2045 1915 2101
rect 1033 1371 1915 2045
rect 3911 3709 4393 4959
rect 9206 5128 9789 5135
rect 9206 5072 9211 5128
rect 9267 5072 9296 5128
rect 9352 5072 9381 5128
rect 9437 5072 9466 5128
rect 9522 5072 9550 5128
rect 9606 5072 9634 5128
rect 9690 5072 9718 5128
rect 9774 5072 9789 5128
rect 9206 5020 9789 5072
rect 9206 4964 9211 5020
rect 9267 4964 9296 5020
rect 9352 4964 9381 5020
rect 9437 4964 9466 5020
rect 9522 4964 9550 5020
rect 9606 4964 9634 5020
rect 9690 4964 9718 5020
rect 9774 4964 9789 5020
rect 4955 4856 5837 4862
rect 4707 4792 4713 4856
rect 4777 4792 4794 4856
rect 4858 4792 4875 4856
rect 4939 4792 4956 4856
rect 5020 4792 5037 4856
rect 5101 4792 5118 4856
rect 5182 4792 5198 4856
rect 5262 4792 5278 4856
rect 5342 4792 5358 4856
rect 5422 4792 5438 4856
rect 5502 4792 5518 4856
rect 5582 4792 5598 4856
rect 5662 4792 5678 4856
rect 5742 4792 5758 4856
rect 5822 4792 5837 4856
rect 4707 4764 5837 4792
rect 4707 4700 4713 4764
rect 4777 4700 4794 4764
rect 4858 4700 4875 4764
rect 4939 4700 4956 4764
rect 5020 4700 5037 4764
rect 5101 4700 5118 4764
rect 5182 4700 5198 4764
rect 5262 4700 5278 4764
rect 5342 4700 5358 4764
rect 5422 4700 5438 4764
rect 5502 4700 5518 4764
rect 5582 4700 5598 4764
rect 5662 4700 5678 4764
rect 5742 4700 5758 4764
rect 5822 4700 5837 4764
rect 4707 4672 5837 4700
rect 4707 4608 4713 4672
rect 4777 4608 4794 4672
rect 4858 4608 4875 4672
rect 4939 4608 4956 4672
rect 5020 4608 5037 4672
rect 5101 4608 5118 4672
rect 5182 4608 5198 4672
rect 5262 4608 5278 4672
rect 5342 4608 5358 4672
rect 5422 4608 5438 4672
rect 5502 4608 5518 4672
rect 5582 4608 5598 4672
rect 5662 4608 5678 4672
rect 5742 4608 5758 4672
rect 5822 4608 5837 4672
rect 4707 4580 5837 4608
rect 4707 4516 4713 4580
rect 4777 4516 4794 4580
rect 4858 4516 4875 4580
rect 4939 4516 4956 4580
rect 5020 4516 5037 4580
rect 5101 4516 5118 4580
rect 5182 4516 5198 4580
rect 5262 4516 5278 4580
rect 5342 4516 5358 4580
rect 5422 4516 5438 4580
rect 5502 4516 5518 4580
rect 5582 4516 5598 4580
rect 5662 4516 5678 4580
rect 5742 4516 5758 4580
rect 5822 4516 5837 4580
rect 4707 4488 5837 4516
rect 4707 4424 4713 4488
rect 4777 4424 4794 4488
rect 4858 4424 4875 4488
rect 4939 4424 4956 4488
rect 5020 4424 5037 4488
rect 5101 4424 5118 4488
rect 5182 4424 5198 4488
rect 5262 4424 5278 4488
rect 5342 4424 5358 4488
rect 5422 4424 5438 4488
rect 5502 4424 5518 4488
rect 5582 4424 5598 4488
rect 5662 4424 5678 4488
rect 5742 4424 5758 4488
rect 5822 4424 5837 4488
rect 4707 4396 5837 4424
rect 4707 4332 4713 4396
rect 4777 4332 4794 4396
rect 4858 4332 4875 4396
rect 4939 4332 4956 4396
rect 5020 4332 5037 4396
rect 5101 4332 5118 4396
rect 5182 4332 5198 4396
rect 5262 4332 5278 4396
rect 5342 4332 5358 4396
rect 5422 4332 5438 4396
rect 5502 4332 5518 4396
rect 5582 4332 5598 4396
rect 5662 4332 5678 4396
rect 5742 4332 5758 4396
rect 5822 4332 5837 4396
rect 7517 4856 8399 4862
rect 7517 4792 7531 4856
rect 7595 4792 7617 4856
rect 7681 4792 7703 4856
rect 7767 4792 7789 4856
rect 7853 4792 7875 4856
rect 7939 4792 7961 4856
rect 8025 4792 8047 4856
rect 8111 4792 8133 4856
rect 8197 4792 8219 4856
rect 8283 4792 8305 4856
rect 8369 4792 8391 4856
rect 8455 4792 8477 4856
rect 8541 4792 8563 4856
rect 8627 4792 8648 4856
rect 8712 4792 8718 4856
rect 7517 4764 8718 4792
rect 7517 4700 7531 4764
rect 7595 4700 7617 4764
rect 7681 4700 7703 4764
rect 7767 4700 7789 4764
rect 7853 4700 7875 4764
rect 7939 4700 7961 4764
rect 8025 4700 8047 4764
rect 8111 4700 8133 4764
rect 8197 4700 8219 4764
rect 8283 4700 8305 4764
rect 8369 4700 8391 4764
rect 8455 4700 8477 4764
rect 8541 4700 8563 4764
rect 8627 4700 8648 4764
rect 8712 4700 8718 4764
rect 7517 4672 8718 4700
rect 7517 4608 7531 4672
rect 7595 4608 7617 4672
rect 7681 4608 7703 4672
rect 7767 4608 7789 4672
rect 7853 4608 7875 4672
rect 7939 4608 7961 4672
rect 8025 4608 8047 4672
rect 8111 4608 8133 4672
rect 8197 4608 8219 4672
rect 8283 4608 8305 4672
rect 8369 4608 8391 4672
rect 8455 4608 8477 4672
rect 8541 4608 8563 4672
rect 8627 4608 8648 4672
rect 8712 4608 8718 4672
rect 7517 4580 8718 4608
rect 7517 4516 7531 4580
rect 7595 4516 7617 4580
rect 7681 4516 7703 4580
rect 7767 4516 7789 4580
rect 7853 4516 7875 4580
rect 7939 4516 7961 4580
rect 8025 4516 8047 4580
rect 8111 4516 8133 4580
rect 8197 4516 8219 4580
rect 8283 4516 8305 4580
rect 8369 4516 8391 4580
rect 8455 4516 8477 4580
rect 8541 4516 8563 4580
rect 8627 4516 8648 4580
rect 8712 4516 8718 4580
rect 7517 4488 8718 4516
rect 7517 4424 7531 4488
rect 7595 4424 7617 4488
rect 7681 4424 7703 4488
rect 7767 4424 7789 4488
rect 7853 4424 7875 4488
rect 7939 4424 7961 4488
rect 8025 4424 8047 4488
rect 8111 4424 8133 4488
rect 8197 4424 8219 4488
rect 8283 4424 8305 4488
rect 8369 4424 8391 4488
rect 8455 4424 8477 4488
rect 8541 4424 8563 4488
rect 8627 4424 8648 4488
rect 8712 4424 8718 4488
rect 7517 4396 8718 4424
tri 4393 3709 4800 4116 sw
rect 3911 2352 4800 3709
rect 1033 1315 1038 1371
rect 1094 1315 1120 1371
rect 1176 1315 1202 1371
rect 1258 1315 1284 1371
rect 1340 1315 1366 1371
rect 1422 1315 1448 1371
rect 1504 1315 1530 1371
rect 1586 1315 1611 1371
rect 1667 1315 1692 1371
rect 1748 1315 1773 1371
rect 1829 1315 1854 1371
rect 1910 1315 1915 1371
rect 1033 1287 1915 1315
rect 1033 1231 1038 1287
rect 1094 1231 1120 1287
rect 1176 1231 1202 1287
rect 1258 1231 1284 1287
rect 1340 1231 1366 1287
rect 1422 1231 1448 1287
rect 1504 1231 1530 1287
rect 1586 1231 1611 1287
rect 1667 1231 1692 1287
rect 1748 1231 1773 1287
rect 1829 1231 1854 1287
rect 1910 1231 1915 1287
rect 1033 1203 1915 1231
rect 1033 1147 1038 1203
rect 1094 1147 1120 1203
rect 1176 1147 1202 1203
rect 1258 1147 1284 1203
rect 1340 1147 1366 1203
rect 1422 1147 1448 1203
rect 1504 1147 1530 1203
rect 1586 1147 1611 1203
rect 1667 1147 1692 1203
rect 1748 1147 1773 1203
rect 1829 1147 1854 1203
rect 1910 1147 1915 1203
rect 1033 1119 1915 1147
rect 1033 1063 1038 1119
rect 1094 1063 1120 1119
rect 1176 1063 1202 1119
rect 1258 1063 1284 1119
rect 1340 1063 1366 1119
rect 1422 1063 1448 1119
rect 1504 1063 1530 1119
rect 1586 1063 1611 1119
rect 1667 1063 1692 1119
rect 1748 1063 1773 1119
rect 1829 1063 1854 1119
rect 1910 1063 1915 1119
rect 1033 1035 1915 1063
rect 1033 979 1038 1035
rect 1094 979 1120 1035
rect 1176 979 1202 1035
rect 1258 979 1284 1035
rect 1340 979 1366 1035
rect 1422 979 1448 1035
rect 1504 979 1530 1035
rect 1586 979 1611 1035
rect 1667 979 1692 1035
rect 1748 979 1773 1035
rect 1829 979 1854 1035
rect 1910 979 1915 1035
rect 1033 547 1915 979
rect 1033 491 1038 547
rect 1094 491 1120 547
rect 1176 491 1202 547
rect 1258 491 1284 547
rect 1340 491 1366 547
rect 1422 491 1448 547
rect 1504 491 1530 547
rect 1586 491 1611 547
rect 1667 491 1692 547
rect 1748 491 1773 547
rect 1829 491 1854 547
rect 1910 491 1915 547
rect 1033 463 1915 491
rect 1033 407 1038 463
rect 1094 407 1120 463
rect 1176 407 1202 463
rect 1258 407 1284 463
rect 1340 407 1366 463
rect 1422 407 1448 463
rect 1504 407 1530 463
rect 1586 407 1611 463
rect 1667 407 1692 463
rect 1748 407 1773 463
rect 1829 407 1854 463
rect 1910 407 1915 463
rect 1033 379 1915 407
rect 1033 323 1038 379
rect 1094 323 1120 379
rect 1176 323 1202 379
rect 1258 323 1284 379
rect 1340 323 1366 379
rect 1422 323 1448 379
rect 1504 323 1530 379
rect 1586 323 1611 379
rect 1667 323 1692 379
rect 1748 323 1773 379
rect 1829 323 1854 379
rect 1910 323 1915 379
rect 1033 295 1915 323
rect 1033 239 1038 295
rect 1094 239 1120 295
rect 1176 239 1202 295
rect 1258 239 1284 295
rect 1340 239 1366 295
rect 1422 239 1448 295
rect 1504 239 1530 295
rect 1586 239 1611 295
rect 1667 239 1692 295
rect 1748 239 1773 295
rect 1829 239 1854 295
rect 1910 239 1915 295
rect 1033 211 1915 239
rect 1033 155 1038 211
rect 1094 155 1120 211
rect 1176 155 1202 211
rect 1258 155 1284 211
rect 1340 155 1366 211
rect 1422 155 1448 211
rect 1504 155 1530 211
rect 1586 155 1611 211
rect 1667 155 1692 211
rect 1748 155 1773 211
rect 1829 155 1854 211
rect 1910 155 1915 211
rect 1033 -2645 1915 155
rect 2675 1682 3601 1687
rect 2675 1626 2680 1682
rect 2736 1626 2766 1682
rect 2822 1626 2852 1682
rect 2908 1626 2938 1682
rect 2994 1626 3024 1682
rect 3080 1626 3110 1682
rect 3166 1626 3196 1682
rect 3252 1626 3281 1682
rect 3337 1626 3366 1682
rect 3422 1626 3451 1682
rect 3507 1626 3536 1682
rect 3592 1626 3601 1682
rect 2675 1548 3601 1626
rect 2675 1492 2680 1548
rect 2736 1492 2766 1548
rect 2822 1492 2852 1548
rect 2908 1492 2938 1548
rect 2994 1492 3024 1548
rect 3080 1492 3110 1548
rect 3166 1492 3196 1548
rect 3252 1492 3281 1548
rect 3337 1492 3366 1548
rect 3422 1492 3451 1548
rect 3507 1492 3536 1548
rect 3592 1492 3601 1548
rect 2675 -3189 3601 1492
rect 3911 858 3924 2352
rect 4788 858 4800 2352
rect 4955 2437 5837 4332
rect 4955 2381 5203 2437
rect 5259 2381 5284 2437
rect 5340 2381 5366 2437
rect 5422 2381 5448 2437
rect 5504 2381 5530 2437
rect 5586 2381 5612 2437
rect 5668 2381 5694 2437
rect 5750 2381 5776 2437
rect 5832 2381 5837 2437
rect 4955 2353 5837 2381
rect 4955 2297 5203 2353
rect 5259 2297 5284 2353
rect 5340 2297 5366 2353
rect 5422 2297 5448 2353
rect 5504 2297 5530 2353
rect 5586 2297 5612 2353
rect 5668 2297 5694 2353
rect 5750 2297 5776 2353
rect 5832 2297 5837 2353
rect 4955 2269 5837 2297
rect 4955 2213 5203 2269
rect 5259 2213 5284 2269
rect 5340 2213 5366 2269
rect 5422 2213 5448 2269
rect 5504 2213 5530 2269
rect 5586 2213 5612 2269
rect 5668 2213 5694 2269
rect 5750 2213 5776 2269
rect 5832 2213 5837 2269
rect 4955 2185 5837 2213
rect 4955 2129 5203 2185
rect 5259 2129 5284 2185
rect 5340 2129 5366 2185
rect 5422 2129 5448 2185
rect 5504 2129 5530 2185
rect 5586 2129 5612 2185
rect 5668 2129 5694 2185
rect 5750 2129 5776 2185
rect 5832 2129 5837 2185
rect 4955 2101 5837 2129
rect 4955 2045 5203 2101
rect 5259 2045 5284 2101
rect 5340 2045 5366 2101
rect 5422 2045 5448 2101
rect 5504 2045 5530 2101
rect 5586 2045 5612 2101
rect 5668 2045 5694 2101
rect 5750 2045 5776 2101
rect 5832 2045 5837 2101
tri 4955 2038 4962 2045 ne
rect 4962 2038 5837 2045
tri 4962 1919 5081 2038 ne
rect 5081 2033 5837 2038
rect 5081 1919 5723 2033
tri 5723 1919 5837 2033 nw
rect 6012 4351 6411 4367
rect 6012 4295 6021 4351
rect 6077 4295 6103 4351
rect 6159 4295 6184 4351
rect 6240 4295 6265 4351
rect 6321 4295 6346 4351
rect 6402 4295 6411 4351
rect 6012 4267 6411 4295
rect 6012 4211 6021 4267
rect 6077 4211 6103 4267
rect 6159 4211 6184 4267
rect 6240 4211 6265 4267
rect 6321 4211 6346 4267
rect 6402 4211 6411 4267
rect 6012 2963 6411 4211
rect 6012 2907 6021 2963
rect 6077 2907 6103 2963
rect 6159 2907 6184 2963
rect 6240 2907 6265 2963
rect 6321 2907 6346 2963
rect 6402 2907 6411 2963
rect 6012 2879 6411 2907
rect 6012 2823 6021 2879
rect 6077 2823 6103 2879
rect 6159 2823 6184 2879
rect 6240 2823 6265 2879
rect 6321 2823 6346 2879
rect 6402 2823 6411 2879
rect 6012 2738 6411 2823
rect 6012 2682 6021 2738
rect 6077 2682 6102 2738
rect 6158 2682 6183 2738
rect 6239 2682 6264 2738
rect 6320 2682 6346 2738
rect 6402 2682 6411 2738
rect 6012 2614 6411 2682
rect 6012 2558 6021 2614
rect 6077 2558 6102 2614
rect 6158 2558 6183 2614
rect 6239 2558 6264 2614
rect 6320 2558 6346 2614
rect 6402 2558 6411 2614
rect 6012 1919 6411 2558
tri 5081 1863 5137 1919 ne
rect 5137 1863 5667 1919
tri 5667 1863 5723 1919 nw
rect 6012 1863 6021 1919
rect 6077 1863 6102 1919
rect 6158 1863 6183 1919
rect 6239 1863 6264 1919
rect 6320 1863 6346 1919
rect 6402 1863 6411 1919
tri 5137 1806 5194 1863 ne
rect 3911 802 3916 858
rect 4795 802 4800 858
rect 3911 724 3924 802
rect 4788 724 4800 802
rect 3911 668 3916 724
rect 4795 668 4800 724
rect 3911 39 3924 668
rect 4788 39 4800 668
rect 3911 -17 3916 39
rect 4795 -17 4800 39
rect 3911 -95 3924 -17
rect 4788 -95 4800 -17
rect 3911 -151 3916 -95
rect 4795 -151 4800 -95
rect 3911 -832 3924 -151
rect 4788 -832 4800 -151
rect 3911 -849 4800 -832
rect 3911 -913 3924 -849
rect 3988 -913 4004 -849
rect 4068 -913 4084 -849
rect 4148 -913 4164 -849
rect 4228 -913 4244 -849
rect 4308 -913 4324 -849
rect 4388 -913 4404 -849
rect 4468 -913 4484 -849
rect 4548 -913 4564 -849
rect 4628 -913 4644 -849
rect 4708 -913 4724 -849
rect 4788 -913 4800 -849
rect 3911 -930 4800 -913
rect 3911 -994 3924 -930
rect 3988 -994 4004 -930
rect 4068 -994 4084 -930
rect 4148 -994 4164 -930
rect 4228 -994 4244 -930
rect 4308 -994 4324 -930
rect 4388 -994 4404 -930
rect 4468 -994 4484 -930
rect 4548 -994 4564 -930
rect 4628 -994 4644 -930
rect 4708 -994 4724 -930
rect 4788 -994 4800 -930
rect 3911 -1011 4800 -994
rect 3911 -1075 3924 -1011
rect 3988 -1075 4004 -1011
rect 4068 -1075 4084 -1011
rect 4148 -1075 4164 -1011
rect 4228 -1075 4244 -1011
rect 4308 -1075 4324 -1011
rect 4388 -1075 4404 -1011
rect 4468 -1075 4484 -1011
rect 4548 -1075 4564 -1011
rect 4628 -1075 4644 -1011
rect 4708 -1075 4724 -1011
rect 4788 -1075 4800 -1011
rect 3911 -1092 4800 -1075
rect 3911 -1156 3924 -1092
rect 3988 -1156 4004 -1092
rect 4068 -1156 4084 -1092
rect 4148 -1156 4164 -1092
rect 4228 -1156 4244 -1092
rect 4308 -1156 4324 -1092
rect 4388 -1156 4404 -1092
rect 4468 -1156 4484 -1092
rect 4548 -1156 4564 -1092
rect 4628 -1156 4644 -1092
rect 4708 -1156 4724 -1092
rect 4788 -1156 4800 -1092
rect 3911 -1173 4800 -1156
rect 3911 -1237 3924 -1173
rect 3988 -1237 4004 -1173
rect 4068 -1237 4084 -1173
rect 4148 -1237 4164 -1173
rect 4228 -1237 4244 -1173
rect 4308 -1237 4324 -1173
rect 4388 -1237 4404 -1173
rect 4468 -1237 4484 -1173
rect 4548 -1237 4564 -1173
rect 4628 -1237 4644 -1173
rect 4708 -1237 4724 -1173
rect 4788 -1237 4800 -1173
rect 3911 -1254 4800 -1237
rect 3911 -1318 3924 -1254
rect 3988 -1318 4004 -1254
rect 4068 -1318 4084 -1254
rect 4148 -1318 4164 -1254
rect 4228 -1318 4244 -1254
rect 4308 -1318 4324 -1254
rect 4388 -1318 4404 -1254
rect 4468 -1318 4484 -1254
rect 4548 -1318 4564 -1254
rect 4628 -1318 4644 -1254
rect 4708 -1318 4724 -1254
rect 4788 -1318 4800 -1254
rect 3911 -1335 4800 -1318
rect 3911 -1399 3924 -1335
rect 3988 -1399 4004 -1335
rect 4068 -1399 4084 -1335
rect 4148 -1399 4164 -1335
rect 4228 -1399 4244 -1335
rect 4308 -1399 4324 -1335
rect 4388 -1399 4404 -1335
rect 4468 -1399 4484 -1335
rect 4548 -1399 4564 -1335
rect 4628 -1399 4644 -1335
rect 4708 -1399 4724 -1335
rect 4788 -1399 4800 -1335
rect 3911 -1416 4800 -1399
rect 3911 -1480 3924 -1416
rect 3988 -1480 4004 -1416
rect 4068 -1480 4084 -1416
rect 4148 -1480 4164 -1416
rect 4228 -1480 4244 -1416
rect 4308 -1480 4324 -1416
rect 4388 -1480 4404 -1416
rect 4468 -1480 4484 -1416
rect 4548 -1480 4564 -1416
rect 4628 -1480 4644 -1416
rect 4708 -1480 4724 -1416
rect 4788 -1480 4800 -1416
rect 3911 -1497 4800 -1480
rect 3911 -1561 3924 -1497
rect 3988 -1561 4004 -1497
rect 4068 -1561 4084 -1497
rect 4148 -1561 4164 -1497
rect 4228 -1561 4244 -1497
rect 4308 -1561 4324 -1497
rect 4388 -1561 4404 -1497
rect 4468 -1561 4484 -1497
rect 4548 -1561 4564 -1497
rect 4628 -1561 4644 -1497
rect 4708 -1561 4724 -1497
rect 4788 -1561 4800 -1497
rect 3911 -1578 4800 -1561
rect 3911 -1642 3924 -1578
rect 3988 -1642 4004 -1578
rect 4068 -1642 4084 -1578
rect 4148 -1642 4164 -1578
rect 4228 -1642 4244 -1578
rect 4308 -1642 4324 -1578
rect 4388 -1642 4404 -1578
rect 4468 -1642 4484 -1578
rect 4548 -1642 4564 -1578
rect 4628 -1642 4644 -1578
rect 4708 -1642 4724 -1578
rect 4788 -1642 4800 -1578
rect 3911 -1659 4800 -1642
rect 3911 -1723 3924 -1659
rect 3988 -1723 4004 -1659
rect 4068 -1723 4084 -1659
rect 4148 -1723 4164 -1659
rect 4228 -1723 4244 -1659
rect 4308 -1723 4324 -1659
rect 4388 -1723 4404 -1659
rect 4468 -1723 4484 -1659
rect 4548 -1723 4564 -1659
rect 4628 -1723 4644 -1659
rect 4708 -1723 4724 -1659
rect 4788 -1723 4800 -1659
rect 3911 -1740 4800 -1723
rect 3911 -1804 3924 -1740
rect 3988 -1804 4004 -1740
rect 4068 -1804 4084 -1740
rect 4148 -1804 4164 -1740
rect 4228 -1804 4244 -1740
rect 4308 -1804 4324 -1740
rect 4388 -1804 4404 -1740
rect 4468 -1804 4484 -1740
rect 4548 -1804 4564 -1740
rect 4628 -1804 4644 -1740
rect 4708 -1804 4724 -1740
rect 4788 -1804 4800 -1740
rect 3911 -1821 4800 -1804
rect 3911 -1885 3924 -1821
rect 3988 -1885 4004 -1821
rect 4068 -1885 4084 -1821
rect 4148 -1885 4164 -1821
rect 4228 -1885 4244 -1821
rect 4308 -1885 4324 -1821
rect 4388 -1885 4404 -1821
rect 4468 -1885 4484 -1821
rect 4548 -1885 4564 -1821
rect 4628 -1885 4644 -1821
rect 4708 -1885 4724 -1821
rect 4788 -1885 4800 -1821
rect 3911 -1902 4800 -1885
rect 3911 -1966 3924 -1902
rect 3988 -1966 4004 -1902
rect 4068 -1966 4084 -1902
rect 4148 -1966 4164 -1902
rect 4228 -1966 4244 -1902
rect 4308 -1966 4324 -1902
rect 4388 -1966 4404 -1902
rect 4468 -1966 4484 -1902
rect 4548 -1966 4564 -1902
rect 4628 -1966 4644 -1902
rect 4708 -1966 4724 -1902
rect 4788 -1966 4800 -1902
rect 3911 -1983 4800 -1966
rect 3911 -2047 3924 -1983
rect 3988 -2047 4004 -1983
rect 4068 -2047 4084 -1983
rect 4148 -2047 4164 -1983
rect 4228 -2047 4244 -1983
rect 4308 -2047 4324 -1983
rect 4388 -2047 4404 -1983
rect 4468 -2047 4484 -1983
rect 4548 -2047 4564 -1983
rect 4628 -2047 4644 -1983
rect 4708 -2047 4724 -1983
rect 4788 -2047 4800 -1983
rect 3911 -2064 4800 -2047
rect 3911 -2128 3924 -2064
rect 3988 -2128 4004 -2064
rect 4068 -2128 4084 -2064
rect 4148 -2128 4164 -2064
rect 4228 -2128 4244 -2064
rect 4308 -2128 4324 -2064
rect 4388 -2128 4404 -2064
rect 4468 -2128 4484 -2064
rect 4548 -2128 4564 -2064
rect 4628 -2128 4644 -2064
rect 4708 -2128 4724 -2064
rect 4788 -2128 4800 -2064
rect 3911 -2145 4800 -2128
rect 3911 -2209 3924 -2145
rect 3988 -2209 4004 -2145
rect 4068 -2209 4084 -2145
rect 4148 -2209 4164 -2145
rect 4228 -2209 4244 -2145
rect 4308 -2209 4324 -2145
rect 4388 -2209 4404 -2145
rect 4468 -2209 4484 -2145
rect 4548 -2209 4564 -2145
rect 4628 -2209 4644 -2145
rect 4708 -2209 4724 -2145
rect 4788 -2209 4800 -2145
rect 3911 -2226 4800 -2209
rect 3911 -2290 3924 -2226
rect 3988 -2290 4004 -2226
rect 4068 -2290 4084 -2226
rect 4148 -2290 4164 -2226
rect 4228 -2290 4244 -2226
rect 4308 -2290 4324 -2226
rect 4388 -2290 4404 -2226
rect 4468 -2290 4484 -2226
rect 4548 -2290 4564 -2226
rect 4628 -2290 4644 -2226
rect 4708 -2290 4724 -2226
rect 4788 -2290 4800 -2226
rect 3911 -2307 4800 -2290
rect 3911 -2371 3924 -2307
rect 3988 -2371 4004 -2307
rect 4068 -2371 4084 -2307
rect 4148 -2371 4164 -2307
rect 4228 -2371 4244 -2307
rect 4308 -2371 4324 -2307
rect 4388 -2371 4404 -2307
rect 4468 -2371 4484 -2307
rect 4548 -2371 4564 -2307
rect 4628 -2371 4644 -2307
rect 4708 -2371 4724 -2307
rect 4788 -2371 4800 -2307
rect 3911 -2388 4800 -2371
rect 3911 -2452 3924 -2388
rect 3988 -2452 4004 -2388
rect 4068 -2452 4084 -2388
rect 4148 -2452 4164 -2388
rect 4228 -2452 4244 -2388
rect 4308 -2452 4324 -2388
rect 4388 -2452 4404 -2388
rect 4468 -2452 4484 -2388
rect 4548 -2452 4564 -2388
rect 4628 -2452 4644 -2388
rect 4708 -2452 4724 -2388
rect 4788 -2452 4800 -2388
rect 3911 -2469 4800 -2452
rect 3911 -2533 3924 -2469
rect 3988 -2533 4004 -2469
rect 4068 -2533 4084 -2469
rect 4148 -2533 4164 -2469
rect 4228 -2533 4244 -2469
rect 4308 -2533 4324 -2469
rect 4388 -2533 4404 -2469
rect 4468 -2533 4484 -2469
rect 4548 -2533 4564 -2469
rect 4628 -2533 4644 -2469
rect 4708 -2533 4724 -2469
rect 4788 -2533 4800 -2469
rect 3911 -2550 4800 -2533
rect 3911 -2614 3924 -2550
rect 3988 -2614 4004 -2550
rect 4068 -2614 4084 -2550
rect 4148 -2614 4164 -2550
rect 4228 -2614 4244 -2550
rect 4308 -2614 4324 -2550
rect 4388 -2614 4404 -2550
rect 4468 -2614 4484 -2550
rect 4548 -2614 4564 -2550
rect 4628 -2614 4644 -2550
rect 4708 -2614 4724 -2550
rect 4788 -2614 4800 -2550
rect 3911 -2645 4800 -2614
tri 4035 -2754 4144 -2645 ne
rect 4144 -2754 4800 -2645
tri 4144 -2763 4153 -2754 ne
rect 4153 -2979 4800 -2754
rect 4880 1682 5113 1687
rect 4880 1626 4885 1682
rect 4941 1626 4969 1682
rect 5025 1626 5052 1682
rect 5108 1626 5113 1682
rect 4880 1548 5113 1626
rect 4880 1492 4885 1548
rect 4941 1492 4969 1548
rect 5025 1492 5052 1548
rect 5108 1492 5113 1548
rect 4880 -2936 5113 1492
rect 5194 1371 5637 1863
tri 5637 1833 5667 1863 nw
rect 6012 1795 6411 1863
rect 6012 1739 6021 1795
rect 6077 1739 6102 1795
rect 6158 1739 6183 1795
rect 6239 1739 6264 1795
rect 6320 1739 6346 1795
rect 6402 1739 6411 1795
rect 5194 1315 5203 1371
rect 5259 1315 5295 1371
rect 5351 1315 5387 1371
rect 5443 1315 5479 1371
rect 5535 1315 5572 1371
rect 5628 1315 5637 1371
rect 5194 1287 5637 1315
rect 5194 1231 5203 1287
rect 5259 1231 5295 1287
rect 5351 1231 5387 1287
rect 5443 1231 5479 1287
rect 5535 1231 5572 1287
rect 5628 1231 5637 1287
rect 5194 1203 5637 1231
rect 5194 1147 5203 1203
rect 5259 1147 5295 1203
rect 5351 1147 5387 1203
rect 5443 1147 5479 1203
rect 5535 1147 5572 1203
rect 5628 1147 5637 1203
rect 5194 1119 5637 1147
rect 5194 1063 5203 1119
rect 5259 1063 5295 1119
rect 5351 1063 5387 1119
rect 5443 1063 5479 1119
rect 5535 1063 5572 1119
rect 5628 1063 5637 1119
rect 5194 1035 5637 1063
rect 5194 979 5203 1035
rect 5259 979 5295 1035
rect 5351 979 5387 1035
rect 5443 979 5479 1035
rect 5535 979 5572 1035
rect 5628 979 5637 1035
rect 5194 547 5637 979
rect 5194 491 5203 547
rect 5259 491 5295 547
rect 5351 491 5387 547
rect 5443 491 5479 547
rect 5535 491 5572 547
rect 5628 491 5637 547
rect 5194 463 5637 491
rect 5194 407 5203 463
rect 5259 407 5295 463
rect 5351 407 5387 463
rect 5443 407 5479 463
rect 5535 407 5572 463
rect 5628 407 5637 463
rect 5194 379 5637 407
rect 5194 323 5203 379
rect 5259 323 5295 379
rect 5351 323 5387 379
rect 5443 323 5479 379
rect 5535 323 5572 379
rect 5628 323 5637 379
rect 5194 295 5637 323
rect 5194 239 5203 295
rect 5259 239 5295 295
rect 5351 239 5387 295
rect 5443 239 5479 295
rect 5535 239 5572 295
rect 5628 239 5637 295
rect 5194 211 5637 239
rect 5194 155 5203 211
rect 5259 155 5295 211
rect 5351 155 5387 211
rect 5443 155 5479 211
rect 5535 155 5572 211
rect 5628 155 5637 211
rect 5194 148 5637 155
rect 5717 1682 5932 1687
rect 5717 1626 5722 1682
rect 5778 1626 5871 1682
rect 5927 1626 5932 1682
rect 5717 1548 5932 1626
rect 5717 1492 5722 1548
rect 5778 1492 5871 1548
rect 5927 1492 5932 1548
rect 4880 -3000 4883 -2936
rect 4947 -3000 4963 -2936
rect 5027 -3000 5043 -2936
rect 5107 -3000 5113 -2936
rect 4880 -3027 5113 -3000
rect 4880 -3091 4883 -3027
rect 4947 -3091 4963 -3027
rect 5027 -3091 5043 -3027
rect 5107 -3091 5113 -3027
rect 4880 -3119 5113 -3091
rect 4880 -3183 4883 -3119
rect 4947 -3183 4963 -3119
rect 5027 -3183 5043 -3119
rect 5107 -3183 5113 -3119
rect 4880 -3211 5113 -3183
rect 4880 -3275 4883 -3211
rect 4947 -3275 4963 -3211
rect 5027 -3275 5043 -3211
rect 5107 -3275 5113 -3211
rect 4880 -3285 5113 -3275
rect 5717 -2930 5932 1492
rect 6012 -155 6411 1739
rect 6943 4351 7342 4367
rect 6943 4295 6952 4351
rect 7008 4295 7034 4351
rect 7090 4295 7115 4351
rect 7171 4295 7196 4351
rect 7252 4295 7277 4351
rect 7333 4295 7342 4351
rect 6943 4267 7342 4295
rect 6943 4211 6952 4267
rect 7008 4211 7034 4267
rect 7090 4211 7115 4267
rect 7171 4211 7196 4267
rect 7252 4211 7277 4267
rect 7333 4211 7342 4267
rect 6943 2963 7342 4211
rect 6943 2907 6952 2963
rect 7008 2907 7034 2963
rect 7090 2907 7115 2963
rect 7171 2907 7196 2963
rect 7252 2907 7277 2963
rect 7333 2907 7342 2963
rect 6943 2879 7342 2907
rect 6943 2823 6952 2879
rect 7008 2823 7034 2879
rect 7090 2823 7115 2879
rect 7171 2823 7196 2879
rect 7252 2823 7277 2879
rect 7333 2823 7342 2879
rect 6943 2738 7342 2823
rect 6943 2682 6952 2738
rect 7008 2682 7034 2738
rect 7090 2682 7115 2738
rect 7171 2682 7196 2738
rect 7252 2682 7277 2738
rect 7333 2682 7342 2738
rect 6943 2614 7342 2682
rect 6943 2558 6952 2614
rect 7008 2558 7034 2614
rect 7090 2558 7115 2614
rect 7171 2558 7196 2614
rect 7252 2558 7277 2614
rect 7333 2558 7342 2614
rect 6943 1919 7342 2558
rect 6943 1863 6952 1919
rect 7008 1863 7034 1919
rect 7090 1863 7115 1919
rect 7171 1863 7196 1919
rect 7252 1863 7277 1919
rect 7333 1863 7342 1919
rect 6943 1795 7342 1863
rect 6943 1739 6952 1795
rect 7008 1739 7034 1795
rect 7090 1739 7115 1795
rect 7171 1739 7196 1795
rect 7252 1739 7277 1795
rect 7333 1739 7342 1795
rect 6012 -211 6021 -155
rect 6077 -211 6103 -155
rect 6159 -211 6184 -155
rect 6240 -211 6265 -155
rect 6321 -211 6346 -155
rect 6402 -211 6411 -155
rect 6012 -239 6411 -211
rect 6012 -295 6021 -239
rect 6077 -295 6103 -239
rect 6159 -295 6184 -239
rect 6240 -295 6265 -239
rect 6321 -295 6346 -239
rect 6402 -295 6411 -239
rect 6012 -2423 6411 -295
rect 6491 1686 6863 1691
rect 6491 1630 6496 1686
rect 6552 1630 6598 1686
rect 6654 1630 6700 1686
rect 6756 1630 6802 1686
rect 6858 1630 6863 1686
rect 6491 1552 6863 1630
rect 6491 1496 6496 1552
rect 6552 1496 6598 1552
rect 6654 1496 6700 1552
rect 6756 1496 6802 1552
rect 6858 1496 6863 1552
tri 5932 -2930 5941 -2921 sw
rect 5717 -2936 5941 -2930
rect 5781 -3000 5797 -2936
rect 5861 -3000 5877 -2936
rect 5717 -3027 5941 -3000
rect 5781 -3091 5797 -3027
rect 5861 -3091 5877 -3027
rect 5717 -3119 5941 -3091
rect 5781 -3183 5797 -3119
rect 5861 -3183 5877 -3119
rect 5717 -3211 5941 -3183
rect 5781 -3275 5797 -3211
rect 5861 -3275 5877 -3211
rect 5717 -3281 5941 -3275
rect 6491 -2936 6863 1496
rect 6943 -155 7342 1739
rect 7517 4332 7531 4396
rect 7595 4332 7617 4396
rect 7681 4332 7703 4396
rect 7767 4332 7789 4396
rect 7853 4332 7875 4396
rect 7939 4332 7961 4396
rect 8025 4332 8047 4396
rect 8111 4332 8133 4396
rect 8197 4332 8219 4396
rect 8283 4332 8305 4396
rect 8369 4332 8391 4396
rect 8455 4332 8477 4396
rect 8541 4332 8563 4396
rect 8627 4332 8648 4396
rect 8712 4332 8718 4396
rect 7517 2437 8399 4332
tri 9155 4211 9206 4262 se
rect 9206 4211 9789 4964
rect 11008 5128 11284 5135
rect 11008 5072 11018 5128
rect 11074 5072 11114 5128
rect 11170 5072 11209 5128
rect 11265 5072 11284 5128
rect 11008 5020 11284 5072
rect 11008 4964 11018 5020
rect 11074 4964 11114 5020
rect 11170 4964 11209 5020
rect 11265 4964 11284 5020
tri 10997 4211 11008 4222 se
rect 11008 4211 11284 4964
tri 8779 3835 9155 4211 se
rect 9155 3835 9789 4211
rect 7517 2381 7522 2437
rect 7578 2381 7604 2437
rect 7660 2381 7686 2437
rect 7742 2381 7768 2437
rect 7824 2381 7850 2437
rect 7906 2381 7932 2437
rect 7988 2381 8014 2437
rect 8070 2381 8095 2437
rect 8151 2381 8176 2437
rect 8232 2381 8257 2437
rect 8313 2381 8338 2437
rect 8394 2381 8399 2437
rect 7517 2353 8399 2381
rect 7517 2297 7522 2353
rect 7578 2297 7604 2353
rect 7660 2297 7686 2353
rect 7742 2297 7768 2353
rect 7824 2297 7850 2353
rect 7906 2297 7932 2353
rect 7988 2297 8014 2353
rect 8070 2297 8095 2353
rect 8151 2297 8176 2353
rect 8232 2297 8257 2353
rect 8313 2297 8338 2353
rect 8394 2297 8399 2353
rect 7517 2269 8399 2297
rect 7517 2213 7522 2269
rect 7578 2213 7604 2269
rect 7660 2213 7686 2269
rect 7742 2213 7768 2269
rect 7824 2213 7850 2269
rect 7906 2213 7932 2269
rect 7988 2213 8014 2269
rect 8070 2213 8095 2269
rect 8151 2213 8176 2269
rect 8232 2213 8257 2269
rect 8313 2213 8338 2269
rect 8394 2213 8399 2269
rect 7517 2185 8399 2213
rect 7517 2129 7522 2185
rect 7578 2129 7604 2185
rect 7660 2129 7686 2185
rect 7742 2129 7768 2185
rect 7824 2129 7850 2185
rect 7906 2129 7932 2185
rect 7988 2129 8014 2185
rect 8070 2129 8095 2185
rect 8151 2129 8176 2185
rect 8232 2129 8257 2185
rect 8313 2129 8338 2185
rect 8394 2129 8399 2185
rect 7517 2101 8399 2129
rect 7517 2045 7522 2101
rect 7578 2045 7604 2101
rect 7660 2045 7686 2101
rect 7742 2045 7768 2101
rect 7824 2045 7850 2101
rect 7906 2045 7932 2101
rect 7988 2045 8014 2101
rect 8070 2045 8095 2101
rect 8151 2045 8176 2101
rect 8232 2045 8257 2101
rect 8313 2045 8338 2101
rect 8394 2045 8399 2101
rect 7517 1371 8399 2045
rect 7517 1315 7522 1371
rect 7578 1315 7604 1371
rect 7660 1315 7686 1371
rect 7742 1315 7768 1371
rect 7824 1315 7850 1371
rect 7906 1315 7932 1371
rect 7988 1315 8014 1371
rect 8070 1315 8095 1371
rect 8151 1315 8176 1371
rect 8232 1315 8257 1371
rect 8313 1315 8338 1371
rect 8394 1315 8399 1371
rect 7517 1287 8399 1315
rect 7517 1231 7522 1287
rect 7578 1231 7604 1287
rect 7660 1231 7686 1287
rect 7742 1231 7768 1287
rect 7824 1231 7850 1287
rect 7906 1231 7932 1287
rect 7988 1231 8014 1287
rect 8070 1231 8095 1287
rect 8151 1231 8176 1287
rect 8232 1231 8257 1287
rect 8313 1231 8338 1287
rect 8394 1231 8399 1287
rect 7517 1203 8399 1231
rect 7517 1147 7522 1203
rect 7578 1147 7604 1203
rect 7660 1147 7686 1203
rect 7742 1147 7768 1203
rect 7824 1147 7850 1203
rect 7906 1147 7932 1203
rect 7988 1147 8014 1203
rect 8070 1147 8095 1203
rect 8151 1147 8176 1203
rect 8232 1147 8257 1203
rect 8313 1147 8338 1203
rect 8394 1147 8399 1203
rect 7517 1119 8399 1147
rect 7517 1063 7522 1119
rect 7578 1063 7604 1119
rect 7660 1063 7686 1119
rect 7742 1063 7768 1119
rect 7824 1063 7850 1119
rect 7906 1063 7932 1119
rect 7988 1063 8014 1119
rect 8070 1063 8095 1119
rect 8151 1063 8176 1119
rect 8232 1063 8257 1119
rect 8313 1063 8338 1119
rect 8394 1063 8399 1119
rect 7517 1035 8399 1063
rect 7517 979 7522 1035
rect 7578 979 7604 1035
rect 7660 979 7686 1035
rect 7742 979 7768 1035
rect 7824 979 7850 1035
rect 7906 979 7932 1035
rect 7988 979 8014 1035
rect 8070 979 8095 1035
rect 8151 979 8176 1035
rect 8232 979 8257 1035
rect 8313 979 8338 1035
rect 8394 979 8399 1035
rect 7517 547 8399 979
rect 7517 491 7522 547
rect 7578 491 7604 547
rect 7660 491 7686 547
rect 7742 491 7768 547
rect 7824 491 7850 547
rect 7906 491 7932 547
rect 7988 491 8014 547
rect 8070 491 8095 547
rect 8151 491 8176 547
rect 8232 491 8257 547
rect 8313 491 8338 547
rect 8394 491 8399 547
rect 7517 463 8399 491
rect 7517 407 7522 463
rect 7578 407 7604 463
rect 7660 407 7686 463
rect 7742 407 7768 463
rect 7824 407 7850 463
rect 7906 407 7932 463
rect 7988 407 8014 463
rect 8070 407 8095 463
rect 8151 407 8176 463
rect 8232 407 8257 463
rect 8313 407 8338 463
rect 8394 407 8399 463
rect 7517 379 8399 407
rect 7517 323 7522 379
rect 7578 323 7604 379
rect 7660 323 7686 379
rect 7742 323 7768 379
rect 7824 323 7850 379
rect 7906 323 7932 379
rect 7988 323 8014 379
rect 8070 323 8095 379
rect 8151 323 8176 379
rect 8232 323 8257 379
rect 8313 323 8338 379
rect 8394 323 8399 379
rect 7517 295 8399 323
rect 7517 239 7522 295
rect 7578 239 7604 295
rect 7660 239 7686 295
rect 7742 239 7768 295
rect 7824 239 7850 295
rect 7906 239 7932 295
rect 7988 239 8014 295
rect 8070 239 8095 295
rect 8151 239 8176 295
rect 8232 239 8257 295
rect 8313 239 8338 295
rect 8394 239 8399 295
rect 7517 211 8399 239
rect 7517 155 7522 211
rect 7578 155 7604 211
rect 7660 155 7686 211
rect 7742 155 7768 211
rect 7824 155 7850 211
rect 7906 155 7932 211
rect 7988 155 8014 211
rect 8070 155 8095 211
rect 8151 155 8176 211
rect 8232 155 8257 211
rect 8313 155 8338 211
rect 8394 155 8399 211
rect 7517 148 8399 155
tri 8554 3610 8779 3835 se
rect 8779 3610 9443 3835
rect 8554 2352 9443 3610
tri 9443 3489 9789 3835 nw
tri 10395 3609 10997 4211 se
rect 10997 3609 11284 4211
rect 8554 858 8568 2352
rect 9432 858 9443 2352
rect 10395 2352 11284 3609
rect 8554 802 8559 858
rect 9438 802 9443 858
rect 8554 724 8568 802
rect 9432 724 9443 802
rect 8554 668 8559 724
rect 9438 668 9443 724
rect 6943 -211 6952 -155
rect 7008 -211 7034 -155
rect 7090 -211 7115 -155
rect 7171 -211 7196 -155
rect 7252 -211 7277 -155
rect 7333 -211 7342 -155
rect 6943 -239 7342 -211
rect 6943 -295 6952 -239
rect 7008 -295 7034 -239
rect 7090 -295 7115 -239
rect 7171 -295 7196 -239
rect 7252 -295 7277 -239
rect 7333 -295 7342 -239
rect 6943 -2423 7342 -295
rect 8554 35 8568 668
rect 9432 35 9443 668
rect 8554 -21 8559 35
rect 9438 -21 9443 35
rect 8554 -99 8568 -21
rect 9432 -99 9443 -21
rect 8554 -155 8559 -99
rect 9438 -155 9443 -99
rect 8554 -832 8568 -155
rect 9432 -832 9443 -155
rect 8554 -849 9443 -832
rect 8554 -913 8568 -849
rect 8632 -913 8648 -849
rect 8712 -913 8728 -849
rect 8792 -913 8808 -849
rect 8872 -913 8888 -849
rect 8952 -913 8968 -849
rect 9032 -913 9048 -849
rect 9112 -913 9128 -849
rect 9192 -913 9208 -849
rect 9272 -913 9288 -849
rect 9352 -913 9368 -849
rect 9432 -913 9443 -849
rect 8554 -930 9443 -913
rect 8554 -994 8568 -930
rect 8632 -994 8648 -930
rect 8712 -994 8728 -930
rect 8792 -994 8808 -930
rect 8872 -994 8888 -930
rect 8952 -994 8968 -930
rect 9032 -994 9048 -930
rect 9112 -994 9128 -930
rect 9192 -994 9208 -930
rect 9272 -994 9288 -930
rect 9352 -994 9368 -930
rect 9432 -994 9443 -930
rect 8554 -1011 9443 -994
rect 8554 -1075 8568 -1011
rect 8632 -1075 8648 -1011
rect 8712 -1075 8728 -1011
rect 8792 -1075 8808 -1011
rect 8872 -1075 8888 -1011
rect 8952 -1075 8968 -1011
rect 9032 -1075 9048 -1011
rect 9112 -1075 9128 -1011
rect 9192 -1075 9208 -1011
rect 9272 -1075 9288 -1011
rect 9352 -1075 9368 -1011
rect 9432 -1075 9443 -1011
rect 8554 -1092 9443 -1075
rect 8554 -1156 8568 -1092
rect 8632 -1156 8648 -1092
rect 8712 -1156 8728 -1092
rect 8792 -1156 8808 -1092
rect 8872 -1156 8888 -1092
rect 8952 -1156 8968 -1092
rect 9032 -1156 9048 -1092
rect 9112 -1156 9128 -1092
rect 9192 -1156 9208 -1092
rect 9272 -1156 9288 -1092
rect 9352 -1156 9368 -1092
rect 9432 -1156 9443 -1092
rect 8554 -1173 9443 -1156
rect 8554 -1237 8568 -1173
rect 8632 -1237 8648 -1173
rect 8712 -1237 8728 -1173
rect 8792 -1237 8808 -1173
rect 8872 -1237 8888 -1173
rect 8952 -1237 8968 -1173
rect 9032 -1237 9048 -1173
rect 9112 -1237 9128 -1173
rect 9192 -1237 9208 -1173
rect 9272 -1237 9288 -1173
rect 9352 -1237 9368 -1173
rect 9432 -1237 9443 -1173
rect 8554 -1254 9443 -1237
rect 8554 -1318 8568 -1254
rect 8632 -1318 8648 -1254
rect 8712 -1318 8728 -1254
rect 8792 -1318 8808 -1254
rect 8872 -1318 8888 -1254
rect 8952 -1318 8968 -1254
rect 9032 -1318 9048 -1254
rect 9112 -1318 9128 -1254
rect 9192 -1318 9208 -1254
rect 9272 -1318 9288 -1254
rect 9352 -1318 9368 -1254
rect 9432 -1318 9443 -1254
rect 8554 -1335 9443 -1318
rect 8554 -1399 8568 -1335
rect 8632 -1399 8648 -1335
rect 8712 -1399 8728 -1335
rect 8792 -1399 8808 -1335
rect 8872 -1399 8888 -1335
rect 8952 -1399 8968 -1335
rect 9032 -1399 9048 -1335
rect 9112 -1399 9128 -1335
rect 9192 -1399 9208 -1335
rect 9272 -1399 9288 -1335
rect 9352 -1399 9368 -1335
rect 9432 -1399 9443 -1335
rect 8554 -1416 9443 -1399
rect 8554 -1480 8568 -1416
rect 8632 -1480 8648 -1416
rect 8712 -1480 8728 -1416
rect 8792 -1480 8808 -1416
rect 8872 -1480 8888 -1416
rect 8952 -1480 8968 -1416
rect 9032 -1480 9048 -1416
rect 9112 -1480 9128 -1416
rect 9192 -1480 9208 -1416
rect 9272 -1480 9288 -1416
rect 9352 -1480 9368 -1416
rect 9432 -1480 9443 -1416
rect 8554 -1497 9443 -1480
rect 8554 -1561 8568 -1497
rect 8632 -1561 8648 -1497
rect 8712 -1561 8728 -1497
rect 8792 -1561 8808 -1497
rect 8872 -1561 8888 -1497
rect 8952 -1561 8968 -1497
rect 9032 -1561 9048 -1497
rect 9112 -1561 9128 -1497
rect 9192 -1561 9208 -1497
rect 9272 -1561 9288 -1497
rect 9352 -1561 9368 -1497
rect 9432 -1561 9443 -1497
rect 8554 -1578 9443 -1561
rect 8554 -1642 8568 -1578
rect 8632 -1642 8648 -1578
rect 8712 -1642 8728 -1578
rect 8792 -1642 8808 -1578
rect 8872 -1642 8888 -1578
rect 8952 -1642 8968 -1578
rect 9032 -1642 9048 -1578
rect 9112 -1642 9128 -1578
rect 9192 -1642 9208 -1578
rect 9272 -1642 9288 -1578
rect 9352 -1642 9368 -1578
rect 9432 -1642 9443 -1578
rect 8554 -1659 9443 -1642
rect 8554 -1723 8568 -1659
rect 8632 -1723 8648 -1659
rect 8712 -1723 8728 -1659
rect 8792 -1723 8808 -1659
rect 8872 -1723 8888 -1659
rect 8952 -1723 8968 -1659
rect 9032 -1723 9048 -1659
rect 9112 -1723 9128 -1659
rect 9192 -1723 9208 -1659
rect 9272 -1723 9288 -1659
rect 9352 -1723 9368 -1659
rect 9432 -1723 9443 -1659
rect 8554 -1740 9443 -1723
rect 8554 -1804 8568 -1740
rect 8632 -1804 8648 -1740
rect 8712 -1804 8728 -1740
rect 8792 -1804 8808 -1740
rect 8872 -1804 8888 -1740
rect 8952 -1804 8968 -1740
rect 9032 -1804 9048 -1740
rect 9112 -1804 9128 -1740
rect 9192 -1804 9208 -1740
rect 9272 -1804 9288 -1740
rect 9352 -1804 9368 -1740
rect 9432 -1804 9443 -1740
rect 8554 -1821 9443 -1804
rect 8554 -1885 8568 -1821
rect 8632 -1885 8648 -1821
rect 8712 -1885 8728 -1821
rect 8792 -1885 8808 -1821
rect 8872 -1885 8888 -1821
rect 8952 -1885 8968 -1821
rect 9032 -1885 9048 -1821
rect 9112 -1885 9128 -1821
rect 9192 -1885 9208 -1821
rect 9272 -1885 9288 -1821
rect 9352 -1885 9368 -1821
rect 9432 -1885 9443 -1821
rect 8554 -1902 9443 -1885
rect 8554 -1966 8568 -1902
rect 8632 -1966 8648 -1902
rect 8712 -1966 8728 -1902
rect 8792 -1966 8808 -1902
rect 8872 -1966 8888 -1902
rect 8952 -1966 8968 -1902
rect 9032 -1966 9048 -1902
rect 9112 -1966 9128 -1902
rect 9192 -1966 9208 -1902
rect 9272 -1966 9288 -1902
rect 9352 -1966 9368 -1902
rect 9432 -1966 9443 -1902
rect 8554 -1983 9443 -1966
rect 8554 -2047 8568 -1983
rect 8632 -2047 8648 -1983
rect 8712 -2047 8728 -1983
rect 8792 -2047 8808 -1983
rect 8872 -2047 8888 -1983
rect 8952 -2047 8968 -1983
rect 9032 -2047 9048 -1983
rect 9112 -2047 9128 -1983
rect 9192 -2047 9208 -1983
rect 9272 -2047 9288 -1983
rect 9352 -2047 9368 -1983
rect 9432 -2047 9443 -1983
rect 8554 -2064 9443 -2047
rect 8554 -2128 8568 -2064
rect 8632 -2128 8648 -2064
rect 8712 -2128 8728 -2064
rect 8792 -2128 8808 -2064
rect 8872 -2128 8888 -2064
rect 8952 -2128 8968 -2064
rect 9032 -2128 9048 -2064
rect 9112 -2128 9128 -2064
rect 9192 -2128 9208 -2064
rect 9272 -2128 9288 -2064
rect 9352 -2128 9368 -2064
rect 9432 -2128 9443 -2064
rect 8554 -2145 9443 -2128
rect 8554 -2209 8568 -2145
rect 8632 -2209 8648 -2145
rect 8712 -2209 8728 -2145
rect 8792 -2209 8808 -2145
rect 8872 -2209 8888 -2145
rect 8952 -2209 8968 -2145
rect 9032 -2209 9048 -2145
rect 9112 -2209 9128 -2145
rect 9192 -2209 9208 -2145
rect 9272 -2209 9288 -2145
rect 9352 -2209 9368 -2145
rect 9432 -2209 9443 -2145
rect 8554 -2226 9443 -2209
rect 8554 -2290 8568 -2226
rect 8632 -2290 8648 -2226
rect 8712 -2290 8728 -2226
rect 8792 -2290 8808 -2226
rect 8872 -2290 8888 -2226
rect 8952 -2290 8968 -2226
rect 9032 -2290 9048 -2226
rect 9112 -2290 9128 -2226
rect 9192 -2290 9208 -2226
rect 9272 -2290 9288 -2226
rect 9352 -2290 9368 -2226
rect 9432 -2290 9443 -2226
rect 8554 -2307 9443 -2290
rect 8554 -2371 8568 -2307
rect 8632 -2371 8648 -2307
rect 8712 -2371 8728 -2307
rect 8792 -2371 8808 -2307
rect 8872 -2371 8888 -2307
rect 8952 -2371 8968 -2307
rect 9032 -2371 9048 -2307
rect 9112 -2371 9128 -2307
rect 9192 -2371 9208 -2307
rect 9272 -2371 9288 -2307
rect 9352 -2371 9368 -2307
rect 9432 -2371 9443 -2307
rect 8554 -2388 9443 -2371
rect 8554 -2452 8568 -2388
rect 8632 -2452 8648 -2388
rect 8712 -2452 8728 -2388
rect 8792 -2452 8808 -2388
rect 8872 -2452 8888 -2388
rect 8952 -2452 8968 -2388
rect 9032 -2452 9048 -2388
rect 9112 -2452 9128 -2388
rect 9192 -2452 9208 -2388
rect 9272 -2452 9288 -2388
rect 9352 -2452 9368 -2388
rect 9432 -2452 9443 -2388
rect 8554 -2469 9443 -2452
rect 8554 -2533 8568 -2469
rect 8632 -2533 8648 -2469
rect 8712 -2533 8728 -2469
rect 8792 -2533 8808 -2469
rect 8872 -2533 8888 -2469
rect 8952 -2533 8968 -2469
rect 9032 -2533 9048 -2469
rect 9112 -2533 9128 -2469
rect 9192 -2533 9208 -2469
rect 9272 -2533 9288 -2469
rect 9352 -2533 9368 -2469
rect 9432 -2533 9443 -2469
rect 8554 -2550 9443 -2533
rect 8554 -2614 8568 -2550
rect 8632 -2614 8648 -2550
rect 8712 -2614 8728 -2550
rect 8792 -2614 8808 -2550
rect 8872 -2614 8888 -2550
rect 8952 -2614 8968 -2550
rect 9032 -2614 9048 -2550
rect 9112 -2614 9128 -2550
rect 9192 -2614 9208 -2550
rect 9272 -2614 9288 -2550
rect 9352 -2614 9368 -2550
rect 9432 -2614 9443 -2550
rect 8554 -2620 9443 -2614
rect 9523 1682 9780 1687
rect 9523 1626 9528 1682
rect 9584 1626 9624 1682
rect 9680 1626 9719 1682
rect 9775 1626 9780 1682
rect 9523 1548 9780 1626
rect 9523 1492 9528 1548
rect 9584 1492 9624 1548
rect 9680 1492 9719 1548
rect 9775 1492 9780 1548
rect 6491 -3000 6492 -2936
rect 6556 -3000 6594 -2936
rect 6658 -3000 6696 -2936
rect 6760 -3000 6798 -2936
rect 6862 -3000 6863 -2936
rect 6491 -3016 6863 -3000
rect 6491 -3080 6492 -3016
rect 6556 -3080 6594 -3016
rect 6658 -3080 6696 -3016
rect 6760 -3080 6798 -3016
rect 6862 -3080 6863 -3016
rect 6491 -3096 6863 -3080
rect 6491 -3160 6492 -3096
rect 6556 -3160 6594 -3096
rect 6658 -3160 6696 -3096
rect 6760 -3160 6798 -3096
rect 6862 -3160 6863 -3096
rect 6491 -3176 6863 -3160
rect 6491 -3240 6492 -3176
rect 6556 -3240 6594 -3176
rect 6658 -3240 6696 -3176
rect 6760 -3240 6798 -3176
rect 6862 -3240 6863 -3176
rect 6491 -3256 6863 -3240
rect 5717 -3285 5932 -3281
rect 6491 -3320 6492 -3256
rect 6556 -3320 6594 -3256
rect 6658 -3320 6696 -3256
rect 6760 -3320 6798 -3256
rect 6862 -3320 6863 -3256
rect 6491 -3337 6863 -3320
rect 6491 -3401 6492 -3337
rect 6556 -3401 6594 -3337
rect 6658 -3401 6696 -3337
rect 6760 -3401 6798 -3337
rect 6862 -3401 6863 -3337
rect 6491 -3418 6863 -3401
rect 6491 -3482 6492 -3418
rect 6556 -3482 6594 -3418
rect 6658 -3482 6696 -3418
rect 6760 -3482 6798 -3418
rect 6862 -3482 6863 -3418
rect 6491 -3499 6863 -3482
rect 6491 -3563 6492 -3499
rect 6556 -3563 6594 -3499
rect 6658 -3563 6696 -3499
rect 6760 -3563 6798 -3499
rect 6862 -3563 6863 -3499
rect 6491 -3580 6863 -3563
rect 6491 -3644 6492 -3580
rect 6556 -3644 6594 -3580
rect 6658 -3644 6696 -3580
rect 6760 -3644 6798 -3580
rect 6862 -3644 6863 -3580
rect 6491 -3661 6863 -3644
rect 6491 -3725 6492 -3661
rect 6556 -3725 6594 -3661
rect 6658 -3725 6696 -3661
rect 6760 -3725 6798 -3661
rect 6862 -3725 6863 -3661
rect 6491 -3742 6863 -3725
rect 9523 -2936 9780 1492
rect 10395 858 10407 2352
rect 11271 858 11284 2352
rect 10395 802 10400 858
rect 11279 802 11284 858
rect 10395 724 10407 802
rect 11271 724 11284 802
rect 10395 668 10400 724
rect 11279 668 11284 724
rect 10395 35 10407 668
rect 11271 35 11284 668
rect 11439 4856 12321 4863
rect 11439 4792 11453 4856
rect 11517 4792 11541 4856
rect 11605 4792 11629 4856
rect 11693 4792 11717 4856
rect 11781 4792 11805 4856
rect 11869 4792 11893 4856
rect 11957 4792 11981 4856
rect 12045 4792 12068 4856
rect 12132 4792 12155 4856
rect 12219 4792 12242 4856
rect 12306 4792 12321 4856
rect 11439 4764 12321 4792
rect 11439 4700 11453 4764
rect 11517 4700 11541 4764
rect 11605 4700 11629 4764
rect 11693 4700 11717 4764
rect 11781 4700 11805 4764
rect 11869 4700 11893 4764
rect 11957 4700 11981 4764
rect 12045 4700 12068 4764
rect 12132 4700 12155 4764
rect 12219 4700 12242 4764
rect 12306 4700 12321 4764
rect 11439 4672 12321 4700
rect 11439 4608 11453 4672
rect 11517 4608 11541 4672
rect 11605 4608 11629 4672
rect 11693 4608 11717 4672
rect 11781 4608 11805 4672
rect 11869 4608 11893 4672
rect 11957 4608 11981 4672
rect 12045 4608 12068 4672
rect 12132 4608 12155 4672
rect 12219 4608 12242 4672
rect 12306 4608 12321 4672
rect 11439 4580 12321 4608
rect 11439 4516 11453 4580
rect 11517 4516 11541 4580
rect 11605 4516 11629 4580
rect 11693 4516 11717 4580
rect 11781 4516 11805 4580
rect 11869 4516 11893 4580
rect 11957 4516 11981 4580
rect 12045 4516 12068 4580
rect 12132 4516 12155 4580
rect 12219 4516 12242 4580
rect 12306 4516 12321 4580
rect 11439 4488 12321 4516
rect 11439 4424 11453 4488
rect 11517 4424 11541 4488
rect 11605 4424 11629 4488
rect 11693 4424 11717 4488
rect 11781 4424 11805 4488
rect 11869 4424 11893 4488
rect 11957 4424 11981 4488
rect 12045 4424 12068 4488
rect 12132 4424 12155 4488
rect 12219 4424 12242 4488
rect 12306 4424 12321 4488
rect 11439 4396 12321 4424
rect 11439 4332 11453 4396
rect 11517 4332 11541 4396
rect 11605 4332 11629 4396
rect 11693 4332 11717 4396
rect 11781 4332 11805 4396
rect 11869 4332 11893 4396
rect 11957 4332 11981 4396
rect 12045 4332 12068 4396
rect 12132 4332 12155 4396
rect 12219 4332 12242 4396
rect 12306 4332 12321 4396
rect 11439 2437 12321 4332
rect 11439 2381 11444 2437
rect 11500 2381 11525 2437
rect 11581 2381 11606 2437
rect 11662 2381 11687 2437
rect 11743 2381 11768 2437
rect 11824 2381 11850 2437
rect 11906 2381 11932 2437
rect 11988 2381 12014 2437
rect 12070 2381 12096 2437
rect 12152 2381 12178 2437
rect 12234 2381 12260 2437
rect 12316 2381 12321 2437
rect 11439 2353 12321 2381
rect 11439 2297 11444 2353
rect 11500 2297 11525 2353
rect 11581 2297 11606 2353
rect 11662 2297 11687 2353
rect 11743 2297 11768 2353
rect 11824 2297 11850 2353
rect 11906 2297 11932 2353
rect 11988 2297 12014 2353
rect 12070 2297 12096 2353
rect 12152 2297 12178 2353
rect 12234 2297 12260 2353
rect 12316 2297 12321 2353
rect 11439 2269 12321 2297
rect 11439 2213 11444 2269
rect 11500 2213 11525 2269
rect 11581 2213 11606 2269
rect 11662 2213 11687 2269
rect 11743 2213 11768 2269
rect 11824 2213 11850 2269
rect 11906 2213 11932 2269
rect 11988 2213 12014 2269
rect 12070 2213 12096 2269
rect 12152 2213 12178 2269
rect 12234 2213 12260 2269
rect 12316 2213 12321 2269
rect 11439 2185 12321 2213
rect 11439 2129 11444 2185
rect 11500 2129 11525 2185
rect 11581 2129 11606 2185
rect 11662 2129 11687 2185
rect 11743 2129 11768 2185
rect 11824 2129 11850 2185
rect 11906 2129 11932 2185
rect 11988 2129 12014 2185
rect 12070 2129 12096 2185
rect 12152 2129 12178 2185
rect 12234 2129 12260 2185
rect 12316 2129 12321 2185
rect 11439 2101 12321 2129
rect 11439 2045 11444 2101
rect 11500 2045 11525 2101
rect 11581 2045 11606 2101
rect 11662 2045 11687 2101
rect 11743 2045 11768 2101
rect 11824 2045 11850 2101
rect 11906 2045 11932 2101
rect 11988 2045 12014 2101
rect 12070 2045 12096 2101
rect 12152 2045 12178 2101
rect 12234 2045 12260 2101
rect 12316 2045 12321 2101
rect 11439 1371 12321 2045
rect 11439 1315 11444 1371
rect 11500 1315 11525 1371
rect 11581 1315 11606 1371
rect 11662 1315 11687 1371
rect 11743 1315 11768 1371
rect 11824 1315 11850 1371
rect 11906 1315 11932 1371
rect 11988 1315 12014 1371
rect 12070 1315 12096 1371
rect 12152 1315 12178 1371
rect 12234 1315 12260 1371
rect 12316 1315 12321 1371
rect 11439 1287 12321 1315
rect 11439 1231 11444 1287
rect 11500 1231 11525 1287
rect 11581 1231 11606 1287
rect 11662 1231 11687 1287
rect 11743 1231 11768 1287
rect 11824 1231 11850 1287
rect 11906 1231 11932 1287
rect 11988 1231 12014 1287
rect 12070 1231 12096 1287
rect 12152 1231 12178 1287
rect 12234 1231 12260 1287
rect 12316 1231 12321 1287
rect 11439 1203 12321 1231
rect 11439 1147 11444 1203
rect 11500 1147 11525 1203
rect 11581 1147 11606 1203
rect 11662 1147 11687 1203
rect 11743 1147 11768 1203
rect 11824 1147 11850 1203
rect 11906 1147 11932 1203
rect 11988 1147 12014 1203
rect 12070 1147 12096 1203
rect 12152 1147 12178 1203
rect 12234 1147 12260 1203
rect 12316 1147 12321 1203
rect 11439 1119 12321 1147
rect 11439 1063 11444 1119
rect 11500 1063 11525 1119
rect 11581 1063 11606 1119
rect 11662 1063 11687 1119
rect 11743 1063 11768 1119
rect 11824 1063 11850 1119
rect 11906 1063 11932 1119
rect 11988 1063 12014 1119
rect 12070 1063 12096 1119
rect 12152 1063 12178 1119
rect 12234 1063 12260 1119
rect 12316 1063 12321 1119
rect 11439 1035 12321 1063
rect 11439 979 11444 1035
rect 11500 979 11525 1035
rect 11581 979 11606 1035
rect 11662 979 11687 1035
rect 11743 979 11768 1035
rect 11824 979 11850 1035
rect 11906 979 11932 1035
rect 11988 979 12014 1035
rect 12070 979 12096 1035
rect 12152 979 12178 1035
rect 12234 979 12260 1035
rect 12316 979 12321 1035
rect 11439 547 12321 979
rect 11439 491 11444 547
rect 11500 491 11525 547
rect 11581 491 11606 547
rect 11662 491 11687 547
rect 11743 491 11768 547
rect 11824 491 11850 547
rect 11906 491 11932 547
rect 11988 491 12014 547
rect 12070 491 12096 547
rect 12152 491 12178 547
rect 12234 491 12260 547
rect 12316 491 12321 547
rect 11439 463 12321 491
rect 11439 407 11444 463
rect 11500 407 11525 463
rect 11581 407 11606 463
rect 11662 407 11687 463
rect 11743 407 11768 463
rect 11824 407 11850 463
rect 11906 407 11932 463
rect 11988 407 12014 463
rect 12070 407 12096 463
rect 12152 407 12178 463
rect 12234 407 12260 463
rect 12316 407 12321 463
rect 11439 379 12321 407
rect 11439 323 11444 379
rect 11500 323 11525 379
rect 11581 323 11606 379
rect 11662 323 11687 379
rect 11743 323 11768 379
rect 11824 323 11850 379
rect 11906 323 11932 379
rect 11988 323 12014 379
rect 12070 323 12096 379
rect 12152 323 12178 379
rect 12234 323 12260 379
rect 12316 323 12321 379
rect 11439 295 12321 323
rect 11439 239 11444 295
rect 11500 239 11525 295
rect 11581 239 11606 295
rect 11662 239 11687 295
rect 11743 239 11768 295
rect 11824 239 11850 295
rect 11906 239 11932 295
rect 11988 239 12014 295
rect 12070 239 12096 295
rect 12152 239 12178 295
rect 12234 239 12260 295
rect 12316 239 12321 295
rect 11439 211 12321 239
rect 11439 155 11444 211
rect 11500 155 11525 211
rect 11581 155 11606 211
rect 11662 155 11687 211
rect 11743 155 11768 211
rect 11824 155 11850 211
rect 11906 155 11932 211
rect 11988 155 12014 211
rect 12070 155 12096 211
rect 12152 155 12178 211
rect 12234 155 12260 211
rect 12316 155 12321 211
rect 11439 147 12321 155
rect 12496 4351 12895 4367
rect 12496 4295 12505 4351
rect 12561 4295 12587 4351
rect 12643 4295 12668 4351
rect 12724 4295 12749 4351
rect 12805 4295 12830 4351
rect 12886 4295 12895 4351
rect 12496 4267 12895 4295
rect 12496 4211 12505 4267
rect 12561 4211 12587 4267
rect 12643 4211 12668 4267
rect 12724 4211 12749 4267
rect 12805 4211 12830 4267
rect 12886 4211 12895 4267
rect 12496 2963 12895 4211
rect 12496 2907 12505 2963
rect 12561 2907 12587 2963
rect 12643 2907 12668 2963
rect 12724 2907 12749 2963
rect 12805 2907 12830 2963
rect 12886 2907 12895 2963
rect 12496 2879 12895 2907
rect 12496 2823 12505 2879
rect 12561 2823 12587 2879
rect 12643 2823 12668 2879
rect 12724 2823 12749 2879
rect 12805 2823 12830 2879
rect 12886 2823 12895 2879
rect 12496 2738 12895 2823
rect 12496 2682 12505 2738
rect 12561 2682 12586 2738
rect 12642 2682 12667 2738
rect 12723 2682 12748 2738
rect 12804 2682 12830 2738
rect 12886 2682 12895 2738
rect 12496 2614 12895 2682
rect 12496 2558 12505 2614
rect 12561 2558 12586 2614
rect 12642 2558 12667 2614
rect 12723 2558 12748 2614
rect 12804 2558 12830 2614
rect 12886 2558 12895 2614
rect 12496 1919 12895 2558
rect 12496 1863 12505 1919
rect 12561 1863 12586 1919
rect 12642 1863 12667 1919
rect 12723 1863 12748 1919
rect 12804 1863 12830 1919
rect 12886 1863 12895 1919
rect 12496 1795 12895 1863
rect 12496 1739 12505 1795
rect 12561 1739 12586 1795
rect 12642 1739 12667 1795
rect 12723 1739 12748 1795
rect 12804 1739 12830 1795
rect 12886 1739 12895 1795
rect 10395 -21 10400 35
rect 11279 -21 11284 35
rect 10395 -99 10407 -21
rect 11271 -99 11284 -21
rect 10395 -155 10400 -99
rect 11279 -155 11284 -99
rect 10395 -832 10407 -155
rect 11271 -832 11284 -155
rect 10395 -849 11284 -832
rect 10395 -913 10407 -849
rect 10471 -913 10487 -849
rect 10551 -913 10567 -849
rect 10631 -913 10647 -849
rect 10711 -913 10727 -849
rect 10791 -913 10807 -849
rect 10871 -913 10887 -849
rect 10951 -913 10967 -849
rect 11031 -913 11047 -849
rect 11111 -913 11127 -849
rect 11191 -913 11207 -849
rect 11271 -913 11284 -849
rect 10395 -930 11284 -913
rect 10395 -994 10407 -930
rect 10471 -994 10487 -930
rect 10551 -994 10567 -930
rect 10631 -994 10647 -930
rect 10711 -994 10727 -930
rect 10791 -994 10807 -930
rect 10871 -994 10887 -930
rect 10951 -994 10967 -930
rect 11031 -994 11047 -930
rect 11111 -994 11127 -930
rect 11191 -994 11207 -930
rect 11271 -994 11284 -930
rect 10395 -1011 11284 -994
rect 10395 -1075 10407 -1011
rect 10471 -1075 10487 -1011
rect 10551 -1075 10567 -1011
rect 10631 -1075 10647 -1011
rect 10711 -1075 10727 -1011
rect 10791 -1075 10807 -1011
rect 10871 -1075 10887 -1011
rect 10951 -1075 10967 -1011
rect 11031 -1075 11047 -1011
rect 11111 -1075 11127 -1011
rect 11191 -1075 11207 -1011
rect 11271 -1075 11284 -1011
rect 10395 -1092 11284 -1075
rect 10395 -1156 10407 -1092
rect 10471 -1156 10487 -1092
rect 10551 -1156 10567 -1092
rect 10631 -1156 10647 -1092
rect 10711 -1156 10727 -1092
rect 10791 -1156 10807 -1092
rect 10871 -1156 10887 -1092
rect 10951 -1156 10967 -1092
rect 11031 -1156 11047 -1092
rect 11111 -1156 11127 -1092
rect 11191 -1156 11207 -1092
rect 11271 -1156 11284 -1092
rect 10395 -1173 11284 -1156
rect 10395 -1237 10407 -1173
rect 10471 -1237 10487 -1173
rect 10551 -1237 10567 -1173
rect 10631 -1237 10647 -1173
rect 10711 -1237 10727 -1173
rect 10791 -1237 10807 -1173
rect 10871 -1237 10887 -1173
rect 10951 -1237 10967 -1173
rect 11031 -1237 11047 -1173
rect 11111 -1237 11127 -1173
rect 11191 -1237 11207 -1173
rect 11271 -1237 11284 -1173
rect 10395 -1254 11284 -1237
rect 10395 -1318 10407 -1254
rect 10471 -1318 10487 -1254
rect 10551 -1318 10567 -1254
rect 10631 -1318 10647 -1254
rect 10711 -1318 10727 -1254
rect 10791 -1318 10807 -1254
rect 10871 -1318 10887 -1254
rect 10951 -1318 10967 -1254
rect 11031 -1318 11047 -1254
rect 11111 -1318 11127 -1254
rect 11191 -1318 11207 -1254
rect 11271 -1318 11284 -1254
rect 10395 -1335 11284 -1318
rect 10395 -1399 10407 -1335
rect 10471 -1399 10487 -1335
rect 10551 -1399 10567 -1335
rect 10631 -1399 10647 -1335
rect 10711 -1399 10727 -1335
rect 10791 -1399 10807 -1335
rect 10871 -1399 10887 -1335
rect 10951 -1399 10967 -1335
rect 11031 -1399 11047 -1335
rect 11111 -1399 11127 -1335
rect 11191 -1399 11207 -1335
rect 11271 -1399 11284 -1335
rect 10395 -1416 11284 -1399
rect 10395 -1480 10407 -1416
rect 10471 -1480 10487 -1416
rect 10551 -1480 10567 -1416
rect 10631 -1480 10647 -1416
rect 10711 -1480 10727 -1416
rect 10791 -1480 10807 -1416
rect 10871 -1480 10887 -1416
rect 10951 -1480 10967 -1416
rect 11031 -1480 11047 -1416
rect 11111 -1480 11127 -1416
rect 11191 -1480 11207 -1416
rect 11271 -1480 11284 -1416
rect 10395 -1497 11284 -1480
rect 10395 -1561 10407 -1497
rect 10471 -1561 10487 -1497
rect 10551 -1561 10567 -1497
rect 10631 -1561 10647 -1497
rect 10711 -1561 10727 -1497
rect 10791 -1561 10807 -1497
rect 10871 -1561 10887 -1497
rect 10951 -1561 10967 -1497
rect 11031 -1561 11047 -1497
rect 11111 -1561 11127 -1497
rect 11191 -1561 11207 -1497
rect 11271 -1561 11284 -1497
rect 10395 -1578 11284 -1561
rect 10395 -1642 10407 -1578
rect 10471 -1642 10487 -1578
rect 10551 -1642 10567 -1578
rect 10631 -1642 10647 -1578
rect 10711 -1642 10727 -1578
rect 10791 -1642 10807 -1578
rect 10871 -1642 10887 -1578
rect 10951 -1642 10967 -1578
rect 11031 -1642 11047 -1578
rect 11111 -1642 11127 -1578
rect 11191 -1642 11207 -1578
rect 11271 -1642 11284 -1578
rect 10395 -1659 11284 -1642
rect 10395 -1723 10407 -1659
rect 10471 -1723 10487 -1659
rect 10551 -1723 10567 -1659
rect 10631 -1723 10647 -1659
rect 10711 -1723 10727 -1659
rect 10791 -1723 10807 -1659
rect 10871 -1723 10887 -1659
rect 10951 -1723 10967 -1659
rect 11031 -1723 11047 -1659
rect 11111 -1723 11127 -1659
rect 11191 -1723 11207 -1659
rect 11271 -1723 11284 -1659
rect 10395 -1740 11284 -1723
rect 10395 -1804 10407 -1740
rect 10471 -1804 10487 -1740
rect 10551 -1804 10567 -1740
rect 10631 -1804 10647 -1740
rect 10711 -1804 10727 -1740
rect 10791 -1804 10807 -1740
rect 10871 -1804 10887 -1740
rect 10951 -1804 10967 -1740
rect 11031 -1804 11047 -1740
rect 11111 -1804 11127 -1740
rect 11191 -1804 11207 -1740
rect 11271 -1804 11284 -1740
rect 10395 -1821 11284 -1804
rect 10395 -1885 10407 -1821
rect 10471 -1885 10487 -1821
rect 10551 -1885 10567 -1821
rect 10631 -1885 10647 -1821
rect 10711 -1885 10727 -1821
rect 10791 -1885 10807 -1821
rect 10871 -1885 10887 -1821
rect 10951 -1885 10967 -1821
rect 11031 -1885 11047 -1821
rect 11111 -1885 11127 -1821
rect 11191 -1885 11207 -1821
rect 11271 -1885 11284 -1821
rect 10395 -1902 11284 -1885
rect 10395 -1966 10407 -1902
rect 10471 -1966 10487 -1902
rect 10551 -1966 10567 -1902
rect 10631 -1966 10647 -1902
rect 10711 -1966 10727 -1902
rect 10791 -1966 10807 -1902
rect 10871 -1966 10887 -1902
rect 10951 -1966 10967 -1902
rect 11031 -1966 11047 -1902
rect 11111 -1966 11127 -1902
rect 11191 -1966 11207 -1902
rect 11271 -1966 11284 -1902
rect 10395 -1983 11284 -1966
rect 10395 -2047 10407 -1983
rect 10471 -2047 10487 -1983
rect 10551 -2047 10567 -1983
rect 10631 -2047 10647 -1983
rect 10711 -2047 10727 -1983
rect 10791 -2047 10807 -1983
rect 10871 -2047 10887 -1983
rect 10951 -2047 10967 -1983
rect 11031 -2047 11047 -1983
rect 11111 -2047 11127 -1983
rect 11191 -2047 11207 -1983
rect 11271 -2047 11284 -1983
rect 10395 -2064 11284 -2047
rect 10395 -2128 10407 -2064
rect 10471 -2128 10487 -2064
rect 10551 -2128 10567 -2064
rect 10631 -2128 10647 -2064
rect 10711 -2128 10727 -2064
rect 10791 -2128 10807 -2064
rect 10871 -2128 10887 -2064
rect 10951 -2128 10967 -2064
rect 11031 -2128 11047 -2064
rect 11111 -2128 11127 -2064
rect 11191 -2128 11207 -2064
rect 11271 -2128 11284 -2064
rect 10395 -2145 11284 -2128
rect 10395 -2209 10407 -2145
rect 10471 -2209 10487 -2145
rect 10551 -2209 10567 -2145
rect 10631 -2209 10647 -2145
rect 10711 -2209 10727 -2145
rect 10791 -2209 10807 -2145
rect 10871 -2209 10887 -2145
rect 10951 -2209 10967 -2145
rect 11031 -2209 11047 -2145
rect 11111 -2209 11127 -2145
rect 11191 -2209 11207 -2145
rect 11271 -2209 11284 -2145
rect 10395 -2226 11284 -2209
rect 10395 -2290 10407 -2226
rect 10471 -2290 10487 -2226
rect 10551 -2290 10567 -2226
rect 10631 -2290 10647 -2226
rect 10711 -2290 10727 -2226
rect 10791 -2290 10807 -2226
rect 10871 -2290 10887 -2226
rect 10951 -2290 10967 -2226
rect 11031 -2290 11047 -2226
rect 11111 -2290 11127 -2226
rect 11191 -2290 11207 -2226
rect 11271 -2290 11284 -2226
rect 10395 -2307 11284 -2290
rect 10395 -2371 10407 -2307
rect 10471 -2371 10487 -2307
rect 10551 -2371 10567 -2307
rect 10631 -2371 10647 -2307
rect 10711 -2371 10727 -2307
rect 10791 -2371 10807 -2307
rect 10871 -2371 10887 -2307
rect 10951 -2371 10967 -2307
rect 11031 -2371 11047 -2307
rect 11111 -2371 11127 -2307
rect 11191 -2371 11207 -2307
rect 11271 -2371 11284 -2307
rect 10395 -2388 11284 -2371
rect 10395 -2452 10407 -2388
rect 10471 -2452 10487 -2388
rect 10551 -2452 10567 -2388
rect 10631 -2452 10647 -2388
rect 10711 -2452 10727 -2388
rect 10791 -2452 10807 -2388
rect 10871 -2452 10887 -2388
rect 10951 -2452 10967 -2388
rect 11031 -2452 11047 -2388
rect 11111 -2452 11127 -2388
rect 11191 -2452 11207 -2388
rect 11271 -2452 11284 -2388
rect 10395 -2469 11284 -2452
rect 10395 -2533 10407 -2469
rect 10471 -2533 10487 -2469
rect 10551 -2533 10567 -2469
rect 10631 -2533 10647 -2469
rect 10711 -2533 10727 -2469
rect 10791 -2533 10807 -2469
rect 10871 -2533 10887 -2469
rect 10951 -2533 10967 -2469
rect 11031 -2533 11047 -2469
rect 11111 -2533 11127 -2469
rect 11191 -2533 11207 -2469
rect 11271 -2533 11284 -2469
rect 10395 -2550 11284 -2533
rect 10395 -2614 10407 -2550
rect 10471 -2614 10487 -2550
rect 10551 -2614 10567 -2550
rect 10631 -2614 10647 -2550
rect 10711 -2614 10727 -2550
rect 10791 -2614 10807 -2550
rect 10871 -2614 10887 -2550
rect 10951 -2614 10967 -2550
rect 11031 -2614 11047 -2550
rect 11111 -2614 11127 -2550
rect 11191 -2614 11207 -2550
rect 11271 -2614 11284 -2550
rect 10395 -2620 11284 -2614
rect 11911 34 12396 39
rect 11911 -22 11924 34
rect 11980 -22 12005 34
rect 12061 -22 12086 34
rect 12142 -22 12167 34
rect 12223 -22 12249 34
rect 12305 -22 12331 34
rect 12387 -22 12396 34
rect 11911 -100 12396 -22
rect 11911 -156 11924 -100
rect 11980 -156 12005 -100
rect 12061 -156 12086 -100
rect 12142 -156 12167 -100
rect 12223 -156 12249 -100
rect 12305 -156 12331 -100
rect 12387 -156 12396 -100
rect 11911 -2620 12396 -156
rect 12496 -155 12895 1739
rect 12496 -211 12505 -155
rect 12561 -211 12587 -155
rect 12643 -211 12668 -155
rect 12724 -211 12749 -155
rect 12805 -211 12830 -155
rect 12886 -211 12895 -155
rect 12496 -239 12895 -211
rect 12496 -295 12505 -239
rect 12561 -295 12587 -239
rect 12643 -295 12668 -239
rect 12724 -295 12749 -239
rect 12805 -295 12830 -239
rect 12886 -295 12895 -239
rect 12496 -2423 12895 -295
rect 13427 4351 13826 4367
rect 13427 4295 13436 4351
rect 13492 4295 13518 4351
rect 13574 4295 13599 4351
rect 13655 4295 13680 4351
rect 13736 4295 13761 4351
rect 13817 4295 13826 4351
rect 13427 4267 13826 4295
rect 13427 4211 13436 4267
rect 13492 4211 13518 4267
rect 13574 4211 13599 4267
rect 13655 4211 13680 4267
rect 13736 4211 13761 4267
rect 13817 4211 13826 4267
rect 13427 2963 13826 4211
rect 13427 2907 13436 2963
rect 13492 2907 13518 2963
rect 13574 2907 13599 2963
rect 13655 2907 13680 2963
rect 13736 2907 13761 2963
rect 13817 2907 13826 2963
rect 13427 2879 13826 2907
rect 13427 2823 13436 2879
rect 13492 2823 13518 2879
rect 13574 2823 13599 2879
rect 13655 2823 13680 2879
rect 13736 2823 13761 2879
rect 13817 2823 13826 2879
rect 13427 2738 13826 2823
rect 13427 2682 13436 2738
rect 13492 2682 13518 2738
rect 13574 2682 13599 2738
rect 13655 2682 13680 2738
rect 13736 2682 13761 2738
rect 13817 2682 13826 2738
rect 13427 2614 13826 2682
rect 13427 2558 13436 2614
rect 13492 2558 13518 2614
rect 13574 2558 13599 2614
rect 13655 2558 13680 2614
rect 13736 2558 13761 2614
rect 13817 2558 13826 2614
rect 13427 1919 13826 2558
rect 13427 1863 13436 1919
rect 13492 1863 13518 1919
rect 13574 1863 13599 1919
rect 13655 1863 13680 1919
rect 13736 1863 13761 1919
rect 13817 1863 13826 1919
rect 13427 1795 13826 1863
rect 13427 1739 13436 1795
rect 13492 1739 13518 1795
rect 13574 1739 13599 1795
rect 13655 1739 13680 1795
rect 13736 1739 13761 1795
rect 13817 1739 13826 1795
rect 13427 -155 13826 1739
rect 13427 -211 13436 -155
rect 13492 -211 13518 -155
rect 13574 -211 13599 -155
rect 13655 -211 13680 -155
rect 13736 -211 13761 -155
rect 13817 -211 13826 -155
rect 13427 -239 13826 -211
rect 13427 -295 13436 -239
rect 13492 -295 13518 -239
rect 13574 -295 13599 -239
rect 13655 -295 13680 -239
rect 13736 -295 13761 -239
rect 13817 -295 13826 -239
rect 13427 -2423 13826 -295
rect 14001 4362 14014 5226
rect 14878 4362 14884 5226
rect 15038 5128 15927 5135
rect 15038 5072 15053 5128
rect 15109 5072 15134 5128
rect 15190 5072 15215 5128
rect 15271 5072 15296 5128
rect 15352 5072 15377 5128
rect 15433 5072 15458 5128
rect 15514 5072 15539 5128
rect 15595 5072 15619 5128
rect 15675 5072 15699 5128
rect 15755 5072 15779 5128
rect 15835 5072 15859 5128
rect 15915 5072 15927 5128
rect 15038 5020 15927 5072
rect 15038 4964 15053 5020
rect 15109 4964 15134 5020
rect 15190 4964 15215 5020
rect 15271 4964 15296 5020
rect 15352 4964 15377 5020
rect 15433 4964 15458 5020
rect 15514 4964 15539 5020
rect 15595 4964 15619 5020
rect 15675 4964 15699 5020
rect 15755 4964 15779 5020
rect 15835 4964 15859 5020
rect 15915 4964 15927 5020
rect 14001 2437 14883 4362
rect 14001 2381 14006 2437
rect 14062 2381 14088 2437
rect 14144 2381 14170 2437
rect 14226 2381 14252 2437
rect 14308 2381 14334 2437
rect 14390 2381 14416 2437
rect 14472 2381 14498 2437
rect 14554 2381 14579 2437
rect 14635 2381 14660 2437
rect 14716 2381 14741 2437
rect 14797 2381 14822 2437
rect 14878 2381 14883 2437
rect 14001 2353 14883 2381
rect 14001 2297 14006 2353
rect 14062 2297 14088 2353
rect 14144 2297 14170 2353
rect 14226 2297 14252 2353
rect 14308 2297 14334 2353
rect 14390 2297 14416 2353
rect 14472 2297 14498 2353
rect 14554 2297 14579 2353
rect 14635 2297 14660 2353
rect 14716 2297 14741 2353
rect 14797 2297 14822 2353
rect 14878 2297 14883 2353
rect 14001 2269 14883 2297
rect 14001 2213 14006 2269
rect 14062 2213 14088 2269
rect 14144 2213 14170 2269
rect 14226 2213 14252 2269
rect 14308 2213 14334 2269
rect 14390 2213 14416 2269
rect 14472 2213 14498 2269
rect 14554 2213 14579 2269
rect 14635 2213 14660 2269
rect 14716 2213 14741 2269
rect 14797 2213 14822 2269
rect 14878 2213 14883 2269
rect 14001 2185 14883 2213
rect 14001 2129 14006 2185
rect 14062 2129 14088 2185
rect 14144 2129 14170 2185
rect 14226 2129 14252 2185
rect 14308 2129 14334 2185
rect 14390 2129 14416 2185
rect 14472 2129 14498 2185
rect 14554 2129 14579 2185
rect 14635 2129 14660 2185
rect 14716 2129 14741 2185
rect 14797 2129 14822 2185
rect 14878 2129 14883 2185
rect 14001 2101 14883 2129
rect 14001 2045 14006 2101
rect 14062 2045 14088 2101
rect 14144 2045 14170 2101
rect 14226 2045 14252 2101
rect 14308 2045 14334 2101
rect 14390 2045 14416 2101
rect 14472 2045 14498 2101
rect 14554 2045 14579 2101
rect 14635 2045 14660 2101
rect 14716 2045 14741 2101
rect 14797 2045 14822 2101
rect 14878 2045 14883 2101
rect 14001 1371 14883 2045
rect 14001 1315 14006 1371
rect 14062 1315 14088 1371
rect 14144 1315 14170 1371
rect 14226 1315 14252 1371
rect 14308 1315 14334 1371
rect 14390 1315 14416 1371
rect 14472 1315 14498 1371
rect 14554 1315 14579 1371
rect 14635 1315 14660 1371
rect 14716 1315 14741 1371
rect 14797 1315 14822 1371
rect 14878 1315 14883 1371
rect 14001 1287 14883 1315
rect 14001 1231 14006 1287
rect 14062 1231 14088 1287
rect 14144 1231 14170 1287
rect 14226 1231 14252 1287
rect 14308 1231 14334 1287
rect 14390 1231 14416 1287
rect 14472 1231 14498 1287
rect 14554 1231 14579 1287
rect 14635 1231 14660 1287
rect 14716 1231 14741 1287
rect 14797 1231 14822 1287
rect 14878 1231 14883 1287
rect 14001 1203 14883 1231
rect 14001 1147 14006 1203
rect 14062 1147 14088 1203
rect 14144 1147 14170 1203
rect 14226 1147 14252 1203
rect 14308 1147 14334 1203
rect 14390 1147 14416 1203
rect 14472 1147 14498 1203
rect 14554 1147 14579 1203
rect 14635 1147 14660 1203
rect 14716 1147 14741 1203
rect 14797 1147 14822 1203
rect 14878 1147 14883 1203
rect 14001 1119 14883 1147
rect 14001 1063 14006 1119
rect 14062 1063 14088 1119
rect 14144 1063 14170 1119
rect 14226 1063 14252 1119
rect 14308 1063 14334 1119
rect 14390 1063 14416 1119
rect 14472 1063 14498 1119
rect 14554 1063 14579 1119
rect 14635 1063 14660 1119
rect 14716 1063 14741 1119
rect 14797 1063 14822 1119
rect 14878 1063 14883 1119
rect 14001 1035 14883 1063
rect 14001 979 14006 1035
rect 14062 979 14088 1035
rect 14144 979 14170 1035
rect 14226 979 14252 1035
rect 14308 979 14334 1035
rect 14390 979 14416 1035
rect 14472 979 14498 1035
rect 14554 979 14579 1035
rect 14635 979 14660 1035
rect 14716 979 14741 1035
rect 14797 979 14822 1035
rect 14878 979 14883 1035
rect 14001 547 14883 979
rect 14001 491 14006 547
rect 14062 491 14088 547
rect 14144 491 14170 547
rect 14226 491 14252 547
rect 14308 491 14334 547
rect 14390 491 14416 547
rect 14472 491 14498 547
rect 14554 491 14579 547
rect 14635 491 14660 547
rect 14716 491 14741 547
rect 14797 491 14822 547
rect 14878 491 14883 547
rect 14001 463 14883 491
rect 14001 407 14006 463
rect 14062 407 14088 463
rect 14144 407 14170 463
rect 14226 407 14252 463
rect 14308 407 14334 463
rect 14390 407 14416 463
rect 14472 407 14498 463
rect 14554 407 14579 463
rect 14635 407 14660 463
rect 14716 407 14741 463
rect 14797 407 14822 463
rect 14878 407 14883 463
rect 14001 379 14883 407
rect 14001 323 14006 379
rect 14062 323 14088 379
rect 14144 323 14170 379
rect 14226 323 14252 379
rect 14308 323 14334 379
rect 14390 323 14416 379
rect 14472 323 14498 379
rect 14554 323 14579 379
rect 14635 323 14660 379
rect 14716 323 14741 379
rect 14797 323 14822 379
rect 14878 323 14883 379
rect 14001 295 14883 323
rect 14001 239 14006 295
rect 14062 239 14088 295
rect 14144 239 14170 295
rect 14226 239 14252 295
rect 14308 239 14334 295
rect 14390 239 14416 295
rect 14472 239 14498 295
rect 14554 239 14579 295
rect 14635 239 14660 295
rect 14716 239 14741 295
rect 14797 239 14822 295
rect 14878 239 14883 295
rect 14001 211 14883 239
rect 14001 155 14006 211
rect 14062 155 14088 211
rect 14144 155 14170 211
rect 14226 155 14252 211
rect 14308 155 14334 211
rect 14390 155 14416 211
rect 14472 155 14498 211
rect 14554 155 14579 211
rect 14635 155 14660 211
rect 14716 155 14741 211
rect 14797 155 14822 211
rect 14878 155 14883 211
tri 12396 -2620 12449 -2567 sw
rect 11911 -2645 12449 -2620
tri 12449 -2645 12474 -2620 sw
rect 14001 -2645 14883 155
rect 15038 2352 15927 4964
rect 15038 858 15052 2352
rect 15916 858 15927 2352
rect 16879 5128 17768 5135
rect 16879 5072 16892 5128
rect 16948 5072 16973 5128
rect 17029 5072 17054 5128
rect 17110 5072 17135 5128
rect 17191 5072 17216 5128
rect 17272 5072 17297 5128
rect 17353 5072 17378 5128
rect 17434 5072 17458 5128
rect 17514 5072 17538 5128
rect 17594 5072 17618 5128
rect 17674 5072 17698 5128
rect 17754 5072 17768 5128
rect 16879 5020 17768 5072
rect 16879 4964 16892 5020
rect 16948 4964 16973 5020
rect 17029 4964 17054 5020
rect 17110 4964 17135 5020
rect 17191 4964 17216 5020
rect 17272 4964 17297 5020
rect 17353 4964 17378 5020
rect 17434 4964 17458 5020
rect 17514 4964 17538 5020
rect 17594 4964 17618 5020
rect 17674 4964 17698 5020
rect 17754 4964 17768 5020
rect 16879 2352 17768 4964
rect 17928 4362 17934 5226
rect 18798 4362 18804 5226
rect 19670 5128 19816 5445
rect 19670 5072 19675 5128
rect 19731 5072 19755 5128
rect 19811 5072 19816 5128
rect 19670 5020 19816 5072
rect 19670 4964 19675 5020
rect 19731 4964 19755 5020
rect 19811 4964 19816 5020
rect 19065 4351 19379 4367
rect 19065 4295 19070 4351
rect 19126 4295 19152 4351
rect 19208 4295 19233 4351
rect 19289 4295 19314 4351
rect 19370 4295 19379 4351
rect 19065 4267 19379 4295
rect 19065 4211 19070 4267
rect 19126 4211 19152 4267
rect 19208 4211 19233 4267
rect 19289 4211 19314 4267
rect 19370 4211 19379 4267
rect 19065 2963 19379 4211
rect 19065 2907 19074 2963
rect 19130 2907 19154 2963
rect 19210 2907 19234 2963
rect 19290 2907 19314 2963
rect 19370 2907 19379 2963
rect 19065 2879 19379 2907
rect 19065 2823 19074 2879
rect 19130 2823 19154 2879
rect 19210 2823 19234 2879
rect 19290 2823 19314 2879
rect 19370 2823 19379 2879
rect 15038 802 15043 858
rect 15922 802 15927 858
rect 15038 724 15052 802
rect 15916 724 15927 802
rect 15038 668 15043 724
rect 15922 668 15927 724
rect 15038 34 15052 668
rect 15916 34 15927 668
rect 15038 -22 15043 34
rect 15922 -22 15927 34
rect 15038 -100 15052 -22
rect 15916 -100 15927 -22
rect 15038 -156 15043 -100
rect 15922 -156 15927 -100
rect 15038 -832 15052 -156
rect 15916 -832 15927 -156
rect 15038 -849 15927 -832
rect 15038 -913 15052 -849
rect 15116 -913 15132 -849
rect 15196 -913 15212 -849
rect 15276 -913 15292 -849
rect 15356 -913 15372 -849
rect 15436 -913 15452 -849
rect 15516 -913 15532 -849
rect 15596 -913 15612 -849
rect 15676 -913 15692 -849
rect 15756 -913 15772 -849
rect 15836 -913 15852 -849
rect 15916 -913 15927 -849
rect 15038 -930 15927 -913
rect 15038 -994 15052 -930
rect 15116 -994 15132 -930
rect 15196 -994 15212 -930
rect 15276 -994 15292 -930
rect 15356 -994 15372 -930
rect 15436 -994 15452 -930
rect 15516 -994 15532 -930
rect 15596 -994 15612 -930
rect 15676 -994 15692 -930
rect 15756 -994 15772 -930
rect 15836 -994 15852 -930
rect 15916 -994 15927 -930
rect 15038 -1011 15927 -994
rect 15038 -1075 15052 -1011
rect 15116 -1075 15132 -1011
rect 15196 -1075 15212 -1011
rect 15276 -1075 15292 -1011
rect 15356 -1075 15372 -1011
rect 15436 -1075 15452 -1011
rect 15516 -1075 15532 -1011
rect 15596 -1075 15612 -1011
rect 15676 -1075 15692 -1011
rect 15756 -1075 15772 -1011
rect 15836 -1075 15852 -1011
rect 15916 -1075 15927 -1011
rect 15038 -1092 15927 -1075
rect 15038 -1156 15052 -1092
rect 15116 -1156 15132 -1092
rect 15196 -1156 15212 -1092
rect 15276 -1156 15292 -1092
rect 15356 -1156 15372 -1092
rect 15436 -1156 15452 -1092
rect 15516 -1156 15532 -1092
rect 15596 -1156 15612 -1092
rect 15676 -1156 15692 -1092
rect 15756 -1156 15772 -1092
rect 15836 -1156 15852 -1092
rect 15916 -1156 15927 -1092
rect 15038 -1173 15927 -1156
rect 15038 -1237 15052 -1173
rect 15116 -1237 15132 -1173
rect 15196 -1237 15212 -1173
rect 15276 -1237 15292 -1173
rect 15356 -1237 15372 -1173
rect 15436 -1237 15452 -1173
rect 15516 -1237 15532 -1173
rect 15596 -1237 15612 -1173
rect 15676 -1237 15692 -1173
rect 15756 -1237 15772 -1173
rect 15836 -1237 15852 -1173
rect 15916 -1237 15927 -1173
rect 15038 -1254 15927 -1237
rect 15038 -1318 15052 -1254
rect 15116 -1318 15132 -1254
rect 15196 -1318 15212 -1254
rect 15276 -1318 15292 -1254
rect 15356 -1318 15372 -1254
rect 15436 -1318 15452 -1254
rect 15516 -1318 15532 -1254
rect 15596 -1318 15612 -1254
rect 15676 -1318 15692 -1254
rect 15756 -1318 15772 -1254
rect 15836 -1318 15852 -1254
rect 15916 -1318 15927 -1254
rect 15038 -1335 15927 -1318
rect 15038 -1399 15052 -1335
rect 15116 -1399 15132 -1335
rect 15196 -1399 15212 -1335
rect 15276 -1399 15292 -1335
rect 15356 -1399 15372 -1335
rect 15436 -1399 15452 -1335
rect 15516 -1399 15532 -1335
rect 15596 -1399 15612 -1335
rect 15676 -1399 15692 -1335
rect 15756 -1399 15772 -1335
rect 15836 -1399 15852 -1335
rect 15916 -1399 15927 -1335
rect 15038 -1416 15927 -1399
rect 15038 -1480 15052 -1416
rect 15116 -1480 15132 -1416
rect 15196 -1480 15212 -1416
rect 15276 -1480 15292 -1416
rect 15356 -1480 15372 -1416
rect 15436 -1480 15452 -1416
rect 15516 -1480 15532 -1416
rect 15596 -1480 15612 -1416
rect 15676 -1480 15692 -1416
rect 15756 -1480 15772 -1416
rect 15836 -1480 15852 -1416
rect 15916 -1480 15927 -1416
rect 15038 -1497 15927 -1480
rect 15038 -1561 15052 -1497
rect 15116 -1561 15132 -1497
rect 15196 -1561 15212 -1497
rect 15276 -1561 15292 -1497
rect 15356 -1561 15372 -1497
rect 15436 -1561 15452 -1497
rect 15516 -1561 15532 -1497
rect 15596 -1561 15612 -1497
rect 15676 -1561 15692 -1497
rect 15756 -1561 15772 -1497
rect 15836 -1561 15852 -1497
rect 15916 -1561 15927 -1497
rect 15038 -1578 15927 -1561
rect 15038 -1642 15052 -1578
rect 15116 -1642 15132 -1578
rect 15196 -1642 15212 -1578
rect 15276 -1642 15292 -1578
rect 15356 -1642 15372 -1578
rect 15436 -1642 15452 -1578
rect 15516 -1642 15532 -1578
rect 15596 -1642 15612 -1578
rect 15676 -1642 15692 -1578
rect 15756 -1642 15772 -1578
rect 15836 -1642 15852 -1578
rect 15916 -1642 15927 -1578
rect 15038 -1659 15927 -1642
rect 15038 -1723 15052 -1659
rect 15116 -1723 15132 -1659
rect 15196 -1723 15212 -1659
rect 15276 -1723 15292 -1659
rect 15356 -1723 15372 -1659
rect 15436 -1723 15452 -1659
rect 15516 -1723 15532 -1659
rect 15596 -1723 15612 -1659
rect 15676 -1723 15692 -1659
rect 15756 -1723 15772 -1659
rect 15836 -1723 15852 -1659
rect 15916 -1723 15927 -1659
rect 15038 -1740 15927 -1723
rect 15038 -1804 15052 -1740
rect 15116 -1804 15132 -1740
rect 15196 -1804 15212 -1740
rect 15276 -1804 15292 -1740
rect 15356 -1804 15372 -1740
rect 15436 -1804 15452 -1740
rect 15516 -1804 15532 -1740
rect 15596 -1804 15612 -1740
rect 15676 -1804 15692 -1740
rect 15756 -1804 15772 -1740
rect 15836 -1804 15852 -1740
rect 15916 -1804 15927 -1740
rect 15038 -1821 15927 -1804
rect 15038 -1885 15052 -1821
rect 15116 -1885 15132 -1821
rect 15196 -1885 15212 -1821
rect 15276 -1885 15292 -1821
rect 15356 -1885 15372 -1821
rect 15436 -1885 15452 -1821
rect 15516 -1885 15532 -1821
rect 15596 -1885 15612 -1821
rect 15676 -1885 15692 -1821
rect 15756 -1885 15772 -1821
rect 15836 -1885 15852 -1821
rect 15916 -1885 15927 -1821
rect 15038 -1902 15927 -1885
rect 15038 -1966 15052 -1902
rect 15116 -1966 15132 -1902
rect 15196 -1966 15212 -1902
rect 15276 -1966 15292 -1902
rect 15356 -1966 15372 -1902
rect 15436 -1966 15452 -1902
rect 15516 -1966 15532 -1902
rect 15596 -1966 15612 -1902
rect 15676 -1966 15692 -1902
rect 15756 -1966 15772 -1902
rect 15836 -1966 15852 -1902
rect 15916 -1966 15927 -1902
rect 15038 -1983 15927 -1966
rect 15038 -2047 15052 -1983
rect 15116 -2047 15132 -1983
rect 15196 -2047 15212 -1983
rect 15276 -2047 15292 -1983
rect 15356 -2047 15372 -1983
rect 15436 -2047 15452 -1983
rect 15516 -2047 15532 -1983
rect 15596 -2047 15612 -1983
rect 15676 -2047 15692 -1983
rect 15756 -2047 15772 -1983
rect 15836 -2047 15852 -1983
rect 15916 -2047 15927 -1983
rect 15038 -2064 15927 -2047
rect 15038 -2128 15052 -2064
rect 15116 -2128 15132 -2064
rect 15196 -2128 15212 -2064
rect 15276 -2128 15292 -2064
rect 15356 -2128 15372 -2064
rect 15436 -2128 15452 -2064
rect 15516 -2128 15532 -2064
rect 15596 -2128 15612 -2064
rect 15676 -2128 15692 -2064
rect 15756 -2128 15772 -2064
rect 15836 -2128 15852 -2064
rect 15916 -2128 15927 -2064
rect 15038 -2145 15927 -2128
rect 15038 -2209 15052 -2145
rect 15116 -2209 15132 -2145
rect 15196 -2209 15212 -2145
rect 15276 -2209 15292 -2145
rect 15356 -2209 15372 -2145
rect 15436 -2209 15452 -2145
rect 15516 -2209 15532 -2145
rect 15596 -2209 15612 -2145
rect 15676 -2209 15692 -2145
rect 15756 -2209 15772 -2145
rect 15836 -2209 15852 -2145
rect 15916 -2209 15927 -2145
rect 15038 -2226 15927 -2209
rect 15038 -2290 15052 -2226
rect 15116 -2290 15132 -2226
rect 15196 -2290 15212 -2226
rect 15276 -2290 15292 -2226
rect 15356 -2290 15372 -2226
rect 15436 -2290 15452 -2226
rect 15516 -2290 15532 -2226
rect 15596 -2290 15612 -2226
rect 15676 -2290 15692 -2226
rect 15756 -2290 15772 -2226
rect 15836 -2290 15852 -2226
rect 15916 -2290 15927 -2226
rect 15038 -2307 15927 -2290
rect 15038 -2371 15052 -2307
rect 15116 -2371 15132 -2307
rect 15196 -2371 15212 -2307
rect 15276 -2371 15292 -2307
rect 15356 -2371 15372 -2307
rect 15436 -2371 15452 -2307
rect 15516 -2371 15532 -2307
rect 15596 -2371 15612 -2307
rect 15676 -2371 15692 -2307
rect 15756 -2371 15772 -2307
rect 15836 -2371 15852 -2307
rect 15916 -2371 15927 -2307
rect 15038 -2388 15927 -2371
rect 15038 -2452 15052 -2388
rect 15116 -2452 15132 -2388
rect 15196 -2452 15212 -2388
rect 15276 -2452 15292 -2388
rect 15356 -2452 15372 -2388
rect 15436 -2452 15452 -2388
rect 15516 -2452 15532 -2388
rect 15596 -2452 15612 -2388
rect 15676 -2452 15692 -2388
rect 15756 -2452 15772 -2388
rect 15836 -2452 15852 -2388
rect 15916 -2452 15927 -2388
rect 15038 -2469 15927 -2452
rect 15038 -2533 15052 -2469
rect 15116 -2533 15132 -2469
rect 15196 -2533 15212 -2469
rect 15276 -2533 15292 -2469
rect 15356 -2533 15372 -2469
rect 15436 -2533 15452 -2469
rect 15516 -2533 15532 -2469
rect 15596 -2533 15612 -2469
rect 15676 -2533 15692 -2469
rect 15756 -2533 15772 -2469
rect 15836 -2533 15852 -2469
rect 15916 -2533 15927 -2469
rect 15038 -2550 15927 -2533
rect 15038 -2614 15052 -2550
rect 15116 -2614 15132 -2550
rect 15196 -2614 15212 -2550
rect 15276 -2614 15292 -2550
rect 15356 -2614 15372 -2550
rect 15436 -2614 15452 -2550
rect 15516 -2614 15532 -2550
rect 15596 -2614 15612 -2550
rect 15676 -2614 15692 -2550
rect 15756 -2614 15772 -2550
rect 15836 -2614 15852 -2550
rect 15916 -2614 15927 -2550
rect 11911 -2754 12474 -2645
tri 12474 -2754 12583 -2645 sw
rect 15038 -2754 15927 -2614
rect 11911 -2810 12583 -2754
tri 12583 -2810 12639 -2754 sw
rect 15038 -2810 15048 -2754
rect 15104 -2810 15129 -2754
rect 15185 -2810 15210 -2754
rect 15266 -2810 15291 -2754
rect 15347 -2810 15372 -2754
rect 15428 -2810 15453 -2754
rect 15509 -2810 15534 -2754
rect 15590 -2810 15614 -2754
rect 15670 -2810 15694 -2754
rect 15750 -2810 15774 -2754
rect 15830 -2810 15854 -2754
rect 15910 -2810 15927 -2754
rect 11911 -2862 12639 -2810
tri 12639 -2862 12691 -2810 sw
rect 15038 -2862 15927 -2810
tri 11881 -2918 11911 -2888 se
rect 11911 -2918 12691 -2862
tri 12691 -2918 12747 -2862 sw
rect 15038 -2918 15048 -2862
rect 15104 -2918 15129 -2862
rect 15185 -2918 15210 -2862
rect 15266 -2918 15291 -2862
rect 15347 -2918 15372 -2862
rect 15428 -2918 15453 -2862
rect 15509 -2918 15534 -2862
rect 15590 -2918 15614 -2862
rect 15670 -2918 15694 -2862
rect 15750 -2918 15774 -2862
rect 15830 -2918 15854 -2862
rect 15910 -2918 15927 -2862
rect 9523 -3000 9540 -2936
rect 9604 -3000 9620 -2936
rect 9684 -3000 9700 -2936
rect 9764 -3000 9780 -2936
rect 9523 -3017 9780 -3000
rect 9523 -3081 9540 -3017
rect 9604 -3081 9620 -3017
rect 9684 -3081 9700 -3017
rect 9764 -3081 9780 -3017
rect 9523 -3098 9780 -3081
rect 9523 -3162 9540 -3098
rect 9604 -3162 9620 -3098
rect 9684 -3162 9700 -3098
rect 9764 -3162 9780 -3098
rect 9523 -3179 9780 -3162
rect 9523 -3243 9540 -3179
rect 9604 -3243 9620 -3179
rect 9684 -3243 9700 -3179
rect 9764 -3243 9780 -3179
rect 9523 -3260 9780 -3243
rect 9523 -3324 9540 -3260
rect 9604 -3324 9620 -3260
rect 9684 -3324 9700 -3260
rect 9764 -3324 9780 -3260
rect 9523 -3341 9780 -3324
rect 9523 -3405 9540 -3341
rect 9604 -3405 9620 -3341
rect 9684 -3405 9700 -3341
rect 9764 -3405 9780 -3341
rect 9523 -3423 9780 -3405
rect 9523 -3487 9540 -3423
rect 9604 -3487 9620 -3423
rect 9684 -3487 9700 -3423
rect 9764 -3487 9780 -3423
rect 9523 -3505 9780 -3487
rect 9523 -3569 9540 -3505
rect 9604 -3569 9620 -3505
rect 9684 -3569 9700 -3505
rect 9764 -3569 9780 -3505
rect 9523 -3587 9780 -3569
rect 9523 -3651 9540 -3587
rect 9604 -3651 9620 -3587
rect 9684 -3651 9700 -3587
rect 9764 -3651 9780 -3587
rect 9523 -3669 9780 -3651
rect 9523 -3733 9540 -3669
rect 9604 -3733 9620 -3669
rect 9684 -3733 9700 -3669
rect 9764 -3733 9780 -3669
rect 9523 -3739 9780 -3733
tri 11862 -2937 11881 -2918 se
rect 11881 -2937 12747 -2918
rect 11862 -2946 12747 -2937
tri 12747 -2946 12775 -2918 sw
rect 6491 -3806 6492 -3742
rect 6556 -3806 6594 -3742
rect 6658 -3806 6696 -3742
rect 6760 -3806 6798 -3742
rect 6862 -3806 6863 -3742
rect 6491 -3816 6863 -3806
rect 11862 -3816 12337 -2946
rect 15038 -3193 15927 -2918
rect 16397 1682 16799 1687
rect 16397 1626 16406 1682
rect 16462 1626 16488 1682
rect 16544 1626 16570 1682
rect 16626 1626 16652 1682
rect 16708 1626 16734 1682
rect 16790 1626 16799 1682
rect 16397 1548 16799 1626
rect 16397 1492 16406 1548
rect 16462 1492 16488 1548
rect 16544 1492 16570 1548
rect 16626 1492 16652 1548
rect 16708 1492 16734 1548
rect 16790 1492 16799 1548
rect 16397 -2936 16799 1492
rect 16397 -3320 16544 -2936
rect 16768 -3320 16799 -2936
rect 16879 858 16891 2352
rect 17755 858 17768 2352
rect 16879 802 16884 858
rect 17763 802 17768 858
rect 16879 724 16891 802
rect 17755 724 17768 802
rect 16879 668 16884 724
rect 17763 668 17768 724
rect 16879 34 16891 668
rect 17755 34 17768 668
rect 16879 -22 16884 34
rect 17763 -22 17768 34
rect 16879 -100 16891 -22
rect 17755 -100 17768 -22
rect 16879 -156 16884 -100
rect 17763 -156 17768 -100
rect 16879 -832 16891 -156
rect 17755 -832 17768 -156
rect 16879 -849 17768 -832
rect 16879 -913 16891 -849
rect 16955 -913 16971 -849
rect 17035 -913 17051 -849
rect 17115 -913 17131 -849
rect 17195 -913 17211 -849
rect 17275 -913 17291 -849
rect 17355 -913 17371 -849
rect 17435 -913 17451 -849
rect 17515 -913 17531 -849
rect 17595 -913 17611 -849
rect 17675 -913 17691 -849
rect 17755 -913 17768 -849
rect 16879 -930 17768 -913
rect 16879 -994 16891 -930
rect 16955 -994 16971 -930
rect 17035 -994 17051 -930
rect 17115 -994 17131 -930
rect 17195 -994 17211 -930
rect 17275 -994 17291 -930
rect 17355 -994 17371 -930
rect 17435 -994 17451 -930
rect 17515 -994 17531 -930
rect 17595 -994 17611 -930
rect 17675 -994 17691 -930
rect 17755 -994 17768 -930
rect 16879 -1011 17768 -994
rect 16879 -1075 16891 -1011
rect 16955 -1075 16971 -1011
rect 17035 -1075 17051 -1011
rect 17115 -1075 17131 -1011
rect 17195 -1075 17211 -1011
rect 17275 -1075 17291 -1011
rect 17355 -1075 17371 -1011
rect 17435 -1075 17451 -1011
rect 17515 -1075 17531 -1011
rect 17595 -1075 17611 -1011
rect 17675 -1075 17691 -1011
rect 17755 -1075 17768 -1011
rect 16879 -1092 17768 -1075
rect 16879 -1156 16891 -1092
rect 16955 -1156 16971 -1092
rect 17035 -1156 17051 -1092
rect 17115 -1156 17131 -1092
rect 17195 -1156 17211 -1092
rect 17275 -1156 17291 -1092
rect 17355 -1156 17371 -1092
rect 17435 -1156 17451 -1092
rect 17515 -1156 17531 -1092
rect 17595 -1156 17611 -1092
rect 17675 -1156 17691 -1092
rect 17755 -1156 17768 -1092
rect 16879 -1173 17768 -1156
rect 16879 -1237 16891 -1173
rect 16955 -1237 16971 -1173
rect 17035 -1237 17051 -1173
rect 17115 -1237 17131 -1173
rect 17195 -1237 17211 -1173
rect 17275 -1237 17291 -1173
rect 17355 -1237 17371 -1173
rect 17435 -1237 17451 -1173
rect 17515 -1237 17531 -1173
rect 17595 -1237 17611 -1173
rect 17675 -1237 17691 -1173
rect 17755 -1237 17768 -1173
rect 16879 -1254 17768 -1237
rect 16879 -1318 16891 -1254
rect 16955 -1318 16971 -1254
rect 17035 -1318 17051 -1254
rect 17115 -1318 17131 -1254
rect 17195 -1318 17211 -1254
rect 17275 -1318 17291 -1254
rect 17355 -1318 17371 -1254
rect 17435 -1318 17451 -1254
rect 17515 -1318 17531 -1254
rect 17595 -1318 17611 -1254
rect 17675 -1318 17691 -1254
rect 17755 -1318 17768 -1254
rect 16879 -1335 17768 -1318
rect 16879 -1399 16891 -1335
rect 16955 -1399 16971 -1335
rect 17035 -1399 17051 -1335
rect 17115 -1399 17131 -1335
rect 17195 -1399 17211 -1335
rect 17275 -1399 17291 -1335
rect 17355 -1399 17371 -1335
rect 17435 -1399 17451 -1335
rect 17515 -1399 17531 -1335
rect 17595 -1399 17611 -1335
rect 17675 -1399 17691 -1335
rect 17755 -1399 17768 -1335
rect 16879 -1416 17768 -1399
rect 16879 -1480 16891 -1416
rect 16955 -1480 16971 -1416
rect 17035 -1480 17051 -1416
rect 17115 -1480 17131 -1416
rect 17195 -1480 17211 -1416
rect 17275 -1480 17291 -1416
rect 17355 -1480 17371 -1416
rect 17435 -1480 17451 -1416
rect 17515 -1480 17531 -1416
rect 17595 -1480 17611 -1416
rect 17675 -1480 17691 -1416
rect 17755 -1480 17768 -1416
rect 16879 -1497 17768 -1480
rect 16879 -1561 16891 -1497
rect 16955 -1561 16971 -1497
rect 17035 -1561 17051 -1497
rect 17115 -1561 17131 -1497
rect 17195 -1561 17211 -1497
rect 17275 -1561 17291 -1497
rect 17355 -1561 17371 -1497
rect 17435 -1561 17451 -1497
rect 17515 -1561 17531 -1497
rect 17595 -1561 17611 -1497
rect 17675 -1561 17691 -1497
rect 17755 -1561 17768 -1497
rect 16879 -1578 17768 -1561
rect 16879 -1642 16891 -1578
rect 16955 -1642 16971 -1578
rect 17035 -1642 17051 -1578
rect 17115 -1642 17131 -1578
rect 17195 -1642 17211 -1578
rect 17275 -1642 17291 -1578
rect 17355 -1642 17371 -1578
rect 17435 -1642 17451 -1578
rect 17515 -1642 17531 -1578
rect 17595 -1642 17611 -1578
rect 17675 -1642 17691 -1578
rect 17755 -1642 17768 -1578
rect 16879 -1659 17768 -1642
rect 16879 -1723 16891 -1659
rect 16955 -1723 16971 -1659
rect 17035 -1723 17051 -1659
rect 17115 -1723 17131 -1659
rect 17195 -1723 17211 -1659
rect 17275 -1723 17291 -1659
rect 17355 -1723 17371 -1659
rect 17435 -1723 17451 -1659
rect 17515 -1723 17531 -1659
rect 17595 -1723 17611 -1659
rect 17675 -1723 17691 -1659
rect 17755 -1723 17768 -1659
rect 16879 -1740 17768 -1723
rect 16879 -1804 16891 -1740
rect 16955 -1804 16971 -1740
rect 17035 -1804 17051 -1740
rect 17115 -1804 17131 -1740
rect 17195 -1804 17211 -1740
rect 17275 -1804 17291 -1740
rect 17355 -1804 17371 -1740
rect 17435 -1804 17451 -1740
rect 17515 -1804 17531 -1740
rect 17595 -1804 17611 -1740
rect 17675 -1804 17691 -1740
rect 17755 -1804 17768 -1740
rect 16879 -1821 17768 -1804
rect 16879 -1885 16891 -1821
rect 16955 -1885 16971 -1821
rect 17035 -1885 17051 -1821
rect 17115 -1885 17131 -1821
rect 17195 -1885 17211 -1821
rect 17275 -1885 17291 -1821
rect 17355 -1885 17371 -1821
rect 17435 -1885 17451 -1821
rect 17515 -1885 17531 -1821
rect 17595 -1885 17611 -1821
rect 17675 -1885 17691 -1821
rect 17755 -1885 17768 -1821
rect 16879 -1902 17768 -1885
rect 16879 -1966 16891 -1902
rect 16955 -1966 16971 -1902
rect 17035 -1966 17051 -1902
rect 17115 -1966 17131 -1902
rect 17195 -1966 17211 -1902
rect 17275 -1966 17291 -1902
rect 17355 -1966 17371 -1902
rect 17435 -1966 17451 -1902
rect 17515 -1966 17531 -1902
rect 17595 -1966 17611 -1902
rect 17675 -1966 17691 -1902
rect 17755 -1966 17768 -1902
rect 16879 -1983 17768 -1966
rect 16879 -2047 16891 -1983
rect 16955 -2047 16971 -1983
rect 17035 -2047 17051 -1983
rect 17115 -2047 17131 -1983
rect 17195 -2047 17211 -1983
rect 17275 -2047 17291 -1983
rect 17355 -2047 17371 -1983
rect 17435 -2047 17451 -1983
rect 17515 -2047 17531 -1983
rect 17595 -2047 17611 -1983
rect 17675 -2047 17691 -1983
rect 17755 -2047 17768 -1983
rect 16879 -2064 17768 -2047
rect 16879 -2128 16891 -2064
rect 16955 -2128 16971 -2064
rect 17035 -2128 17051 -2064
rect 17115 -2128 17131 -2064
rect 17195 -2128 17211 -2064
rect 17275 -2128 17291 -2064
rect 17355 -2128 17371 -2064
rect 17435 -2128 17451 -2064
rect 17515 -2128 17531 -2064
rect 17595 -2128 17611 -2064
rect 17675 -2128 17691 -2064
rect 17755 -2128 17768 -2064
rect 16879 -2145 17768 -2128
rect 16879 -2209 16891 -2145
rect 16955 -2209 16971 -2145
rect 17035 -2209 17051 -2145
rect 17115 -2209 17131 -2145
rect 17195 -2209 17211 -2145
rect 17275 -2209 17291 -2145
rect 17355 -2209 17371 -2145
rect 17435 -2209 17451 -2145
rect 17515 -2209 17531 -2145
rect 17595 -2209 17611 -2145
rect 17675 -2209 17691 -2145
rect 17755 -2209 17768 -2145
rect 16879 -2226 17768 -2209
rect 16879 -2290 16891 -2226
rect 16955 -2290 16971 -2226
rect 17035 -2290 17051 -2226
rect 17115 -2290 17131 -2226
rect 17195 -2290 17211 -2226
rect 17275 -2290 17291 -2226
rect 17355 -2290 17371 -2226
rect 17435 -2290 17451 -2226
rect 17515 -2290 17531 -2226
rect 17595 -2290 17611 -2226
rect 17675 -2290 17691 -2226
rect 17755 -2290 17768 -2226
rect 16879 -2307 17768 -2290
rect 16879 -2371 16891 -2307
rect 16955 -2371 16971 -2307
rect 17035 -2371 17051 -2307
rect 17115 -2371 17131 -2307
rect 17195 -2371 17211 -2307
rect 17275 -2371 17291 -2307
rect 17355 -2371 17371 -2307
rect 17435 -2371 17451 -2307
rect 17515 -2371 17531 -2307
rect 17595 -2371 17611 -2307
rect 17675 -2371 17691 -2307
rect 17755 -2371 17768 -2307
rect 16879 -2388 17768 -2371
rect 16879 -2452 16891 -2388
rect 16955 -2452 16971 -2388
rect 17035 -2452 17051 -2388
rect 17115 -2452 17131 -2388
rect 17195 -2452 17211 -2388
rect 17275 -2452 17291 -2388
rect 17355 -2452 17371 -2388
rect 17435 -2452 17451 -2388
rect 17515 -2452 17531 -2388
rect 17595 -2452 17611 -2388
rect 17675 -2452 17691 -2388
rect 17755 -2452 17768 -2388
rect 16879 -2469 17768 -2452
rect 16879 -2533 16891 -2469
rect 16955 -2533 16971 -2469
rect 17035 -2533 17051 -2469
rect 17115 -2533 17131 -2469
rect 17195 -2533 17211 -2469
rect 17275 -2533 17291 -2469
rect 17355 -2533 17371 -2469
rect 17435 -2533 17451 -2469
rect 17515 -2533 17531 -2469
rect 17595 -2533 17611 -2469
rect 17675 -2533 17691 -2469
rect 17755 -2533 17768 -2469
rect 16879 -2550 17768 -2533
rect 16879 -2614 16891 -2550
rect 16955 -2614 16971 -2550
rect 17035 -2614 17051 -2550
rect 17115 -2614 17131 -2550
rect 17195 -2614 17211 -2550
rect 17275 -2614 17291 -2550
rect 17355 -2614 17371 -2550
rect 17435 -2614 17451 -2550
rect 17515 -2614 17531 -2550
rect 17595 -2614 17611 -2550
rect 17675 -2614 17691 -2550
rect 17755 -2614 17768 -2550
rect 16879 -2754 17768 -2614
rect 16879 -2810 16889 -2754
rect 16945 -2810 16970 -2754
rect 17026 -2810 17051 -2754
rect 17107 -2810 17132 -2754
rect 17188 -2810 17213 -2754
rect 17269 -2810 17294 -2754
rect 17350 -2810 17375 -2754
rect 17431 -2810 17455 -2754
rect 17511 -2810 17535 -2754
rect 17591 -2810 17615 -2754
rect 17671 -2810 17695 -2754
rect 17751 -2810 17768 -2754
rect 16879 -2862 17768 -2810
rect 16879 -2918 16889 -2862
rect 16945 -2918 16970 -2862
rect 17026 -2918 17051 -2862
rect 17107 -2918 17132 -2862
rect 17188 -2918 17213 -2862
rect 17269 -2918 17294 -2862
rect 17350 -2918 17375 -2862
rect 17431 -2918 17455 -2862
rect 17511 -2918 17535 -2862
rect 17591 -2918 17615 -2862
rect 17671 -2918 17695 -2862
rect 17751 -2918 17768 -2862
rect 17923 2437 18805 2751
rect 17923 2381 17928 2437
rect 17984 2381 18009 2437
rect 18065 2381 18090 2437
rect 18146 2381 18171 2437
rect 18227 2381 18252 2437
rect 18308 2381 18334 2437
rect 18390 2381 18416 2437
rect 18472 2381 18498 2437
rect 18554 2381 18580 2437
rect 18636 2381 18662 2437
rect 18718 2381 18744 2437
rect 18800 2381 18805 2437
rect 17923 2353 18805 2381
rect 17923 2297 17928 2353
rect 17984 2297 18009 2353
rect 18065 2297 18090 2353
rect 18146 2297 18171 2353
rect 18227 2297 18252 2353
rect 18308 2297 18334 2353
rect 18390 2297 18416 2353
rect 18472 2297 18498 2353
rect 18554 2297 18580 2353
rect 18636 2297 18662 2353
rect 18718 2297 18744 2353
rect 18800 2297 18805 2353
rect 17923 2269 18805 2297
rect 17923 2213 17928 2269
rect 17984 2213 18009 2269
rect 18065 2213 18090 2269
rect 18146 2213 18171 2269
rect 18227 2213 18252 2269
rect 18308 2213 18334 2269
rect 18390 2213 18416 2269
rect 18472 2213 18498 2269
rect 18554 2213 18580 2269
rect 18636 2213 18662 2269
rect 18718 2213 18744 2269
rect 18800 2213 18805 2269
rect 17923 2185 18805 2213
rect 17923 2129 17928 2185
rect 17984 2129 18009 2185
rect 18065 2129 18090 2185
rect 18146 2129 18171 2185
rect 18227 2129 18252 2185
rect 18308 2129 18334 2185
rect 18390 2129 18416 2185
rect 18472 2129 18498 2185
rect 18554 2129 18580 2185
rect 18636 2129 18662 2185
rect 18718 2129 18744 2185
rect 18800 2129 18805 2185
rect 17923 2101 18805 2129
rect 17923 2045 17928 2101
rect 17984 2045 18009 2101
rect 18065 2045 18090 2101
rect 18146 2045 18171 2101
rect 18227 2045 18252 2101
rect 18308 2045 18334 2101
rect 18390 2045 18416 2101
rect 18472 2045 18498 2101
rect 18554 2045 18580 2101
rect 18636 2045 18662 2101
rect 18718 2045 18744 2101
rect 18800 2045 18805 2101
rect 17923 1371 18805 2045
rect 17923 1315 17928 1371
rect 17984 1315 18009 1371
rect 18065 1315 18090 1371
rect 18146 1315 18171 1371
rect 18227 1315 18252 1371
rect 18308 1315 18334 1371
rect 18390 1315 18416 1371
rect 18472 1315 18498 1371
rect 18554 1315 18580 1371
rect 18636 1315 18662 1371
rect 18718 1315 18744 1371
rect 18800 1315 18805 1371
rect 17923 1287 18805 1315
rect 17923 1231 17928 1287
rect 17984 1231 18009 1287
rect 18065 1231 18090 1287
rect 18146 1231 18171 1287
rect 18227 1231 18252 1287
rect 18308 1231 18334 1287
rect 18390 1231 18416 1287
rect 18472 1231 18498 1287
rect 18554 1231 18580 1287
rect 18636 1231 18662 1287
rect 18718 1231 18744 1287
rect 18800 1231 18805 1287
rect 17923 1203 18805 1231
rect 17923 1147 17928 1203
rect 17984 1147 18009 1203
rect 18065 1147 18090 1203
rect 18146 1147 18171 1203
rect 18227 1147 18252 1203
rect 18308 1147 18334 1203
rect 18390 1147 18416 1203
rect 18472 1147 18498 1203
rect 18554 1147 18580 1203
rect 18636 1147 18662 1203
rect 18718 1147 18744 1203
rect 18800 1147 18805 1203
rect 17923 1119 18805 1147
rect 17923 1063 17928 1119
rect 17984 1063 18009 1119
rect 18065 1063 18090 1119
rect 18146 1063 18171 1119
rect 18227 1063 18252 1119
rect 18308 1063 18334 1119
rect 18390 1063 18416 1119
rect 18472 1063 18498 1119
rect 18554 1063 18580 1119
rect 18636 1063 18662 1119
rect 18718 1063 18744 1119
rect 18800 1063 18805 1119
rect 17923 1035 18805 1063
rect 17923 979 17928 1035
rect 17984 979 18009 1035
rect 18065 979 18090 1035
rect 18146 979 18171 1035
rect 18227 979 18252 1035
rect 18308 979 18334 1035
rect 18390 979 18416 1035
rect 18472 979 18498 1035
rect 18554 979 18580 1035
rect 18636 979 18662 1035
rect 18718 979 18744 1035
rect 18800 979 18805 1035
rect 17923 547 18805 979
rect 17923 491 17928 547
rect 17984 491 18009 547
rect 18065 491 18090 547
rect 18146 491 18171 547
rect 18227 491 18252 547
rect 18308 491 18334 547
rect 18390 491 18416 547
rect 18472 491 18498 547
rect 18554 491 18580 547
rect 18636 491 18662 547
rect 18718 491 18744 547
rect 18800 491 18805 547
rect 17923 463 18805 491
rect 17923 407 17928 463
rect 17984 407 18009 463
rect 18065 407 18090 463
rect 18146 407 18171 463
rect 18227 407 18252 463
rect 18308 407 18334 463
rect 18390 407 18416 463
rect 18472 407 18498 463
rect 18554 407 18580 463
rect 18636 407 18662 463
rect 18718 407 18744 463
rect 18800 407 18805 463
rect 17923 379 18805 407
rect 17923 323 17928 379
rect 17984 323 18009 379
rect 18065 323 18090 379
rect 18146 323 18171 379
rect 18227 323 18252 379
rect 18308 323 18334 379
rect 18390 323 18416 379
rect 18472 323 18498 379
rect 18554 323 18580 379
rect 18636 323 18662 379
rect 18718 323 18744 379
rect 18800 323 18805 379
rect 17923 295 18805 323
rect 17923 239 17928 295
rect 17984 239 18009 295
rect 18065 239 18090 295
rect 18146 239 18171 295
rect 18227 239 18252 295
rect 18308 239 18334 295
rect 18390 239 18416 295
rect 18472 239 18498 295
rect 18554 239 18580 295
rect 18636 239 18662 295
rect 18718 239 18744 295
rect 18800 239 18805 295
rect 17923 211 18805 239
rect 17923 155 17928 211
rect 17984 155 18009 211
rect 18065 155 18090 211
rect 18146 155 18171 211
rect 18227 155 18252 211
rect 18308 155 18334 211
rect 18390 155 18416 211
rect 18472 155 18498 211
rect 18554 155 18580 211
rect 18636 155 18662 211
rect 18718 155 18744 211
rect 18800 155 18805 211
rect 17923 -2874 18805 155
rect 19065 2738 19379 2823
rect 19065 2682 19074 2738
rect 19130 2682 19154 2738
rect 19210 2682 19234 2738
rect 19290 2682 19314 2738
rect 19370 2682 19379 2738
rect 19065 2614 19379 2682
rect 19065 2558 19074 2614
rect 19130 2558 19154 2614
rect 19210 2558 19234 2614
rect 19290 2558 19314 2614
rect 19370 2558 19379 2614
rect 19065 1919 19379 2558
rect 19065 1863 19074 1919
rect 19130 1863 19154 1919
rect 19210 1863 19234 1919
rect 19290 1863 19314 1919
rect 19370 1863 19379 1919
rect 19065 1795 19379 1863
rect 19065 1739 19074 1795
rect 19130 1739 19154 1795
rect 19210 1739 19234 1795
rect 19290 1739 19314 1795
rect 19370 1739 19379 1795
rect 19065 -155 19379 1739
rect 19670 -89 19816 4964
rect 19065 -211 19074 -155
rect 19130 -211 19154 -155
rect 19210 -211 19234 -155
rect 19290 -211 19314 -155
rect 19370 -211 19379 -155
rect 19065 -239 19379 -211
rect 19065 -295 19074 -239
rect 19130 -295 19154 -239
rect 19210 -295 19234 -239
rect 19290 -295 19314 -239
rect 19370 -295 19379 -239
rect 19065 -2423 19379 -295
rect 16879 -3196 17768 -2918
rect 16397 -3337 16799 -3320
rect 16397 -3401 16544 -3337
rect 16608 -3401 16624 -3337
rect 16688 -3401 16704 -3337
rect 16768 -3401 16799 -3337
rect 16397 -3418 16799 -3401
rect 16397 -3482 16544 -3418
rect 16608 -3482 16624 -3418
rect 16688 -3482 16704 -3418
rect 16768 -3482 16799 -3418
rect 16397 -3499 16799 -3482
rect 16397 -3563 16544 -3499
rect 16608 -3563 16624 -3499
rect 16688 -3563 16704 -3499
rect 16768 -3563 16799 -3499
rect 16397 -3580 16799 -3563
rect 16397 -3644 16544 -3580
rect 16608 -3644 16624 -3580
rect 16688 -3644 16704 -3580
rect 16768 -3644 16799 -3580
rect 16397 -3661 16799 -3644
rect 16397 -3725 16544 -3661
rect 16608 -3725 16624 -3661
rect 16688 -3725 16704 -3661
rect 16768 -3725 16799 -3661
rect 16397 -3742 16799 -3725
rect 16397 -3806 16544 -3742
rect 16608 -3806 16624 -3742
rect 16688 -3806 16704 -3742
rect 16768 -3806 16799 -3742
rect 16397 -3816 16799 -3806
<< via3 >>
rect 1047 4792 1111 4856
rect 1135 4792 1199 4856
rect 1223 4792 1287 4856
rect 1311 4792 1375 4856
rect 1399 4792 1463 4856
rect 1487 4792 1551 4856
rect 1575 4792 1639 4856
rect 1662 4792 1726 4856
rect 1749 4792 1813 4856
rect 1836 4792 1900 4856
rect 1047 4700 1111 4764
rect 1135 4700 1199 4764
rect 1223 4700 1287 4764
rect 1311 4700 1375 4764
rect 1399 4700 1463 4764
rect 1487 4700 1551 4764
rect 1575 4700 1639 4764
rect 1662 4700 1726 4764
rect 1749 4700 1813 4764
rect 1836 4700 1900 4764
rect 1047 4608 1111 4672
rect 1135 4608 1199 4672
rect 1223 4608 1287 4672
rect 1311 4608 1375 4672
rect 1399 4608 1463 4672
rect 1487 4608 1551 4672
rect 1575 4608 1639 4672
rect 1662 4608 1726 4672
rect 1749 4608 1813 4672
rect 1836 4608 1900 4672
rect 1047 4516 1111 4580
rect 1135 4516 1199 4580
rect 1223 4516 1287 4580
rect 1311 4516 1375 4580
rect 1399 4516 1463 4580
rect 1487 4516 1551 4580
rect 1575 4516 1639 4580
rect 1662 4516 1726 4580
rect 1749 4516 1813 4580
rect 1836 4516 1900 4580
rect 1047 4424 1111 4488
rect 1135 4424 1199 4488
rect 1223 4424 1287 4488
rect 1311 4424 1375 4488
rect 1399 4424 1463 4488
rect 1487 4424 1551 4488
rect 1575 4424 1639 4488
rect 1662 4424 1726 4488
rect 1749 4424 1813 4488
rect 1836 4424 1900 4488
rect 1047 4332 1111 4396
rect 1135 4332 1199 4396
rect 1223 4332 1287 4396
rect 1311 4332 1375 4396
rect 1399 4332 1463 4396
rect 1487 4332 1551 4396
rect 1575 4332 1639 4396
rect 1662 4332 1726 4396
rect 1749 4332 1813 4396
rect 1836 4332 1900 4396
rect 4713 4792 4777 4856
rect 4794 4792 4858 4856
rect 4875 4792 4939 4856
rect 4956 4792 5020 4856
rect 5037 4792 5101 4856
rect 5118 4792 5182 4856
rect 5198 4792 5262 4856
rect 5278 4792 5342 4856
rect 5358 4792 5422 4856
rect 5438 4792 5502 4856
rect 5518 4792 5582 4856
rect 5598 4792 5662 4856
rect 5678 4792 5742 4856
rect 5758 4792 5822 4856
rect 4713 4700 4777 4764
rect 4794 4700 4858 4764
rect 4875 4700 4939 4764
rect 4956 4700 5020 4764
rect 5037 4700 5101 4764
rect 5118 4700 5182 4764
rect 5198 4700 5262 4764
rect 5278 4700 5342 4764
rect 5358 4700 5422 4764
rect 5438 4700 5502 4764
rect 5518 4700 5582 4764
rect 5598 4700 5662 4764
rect 5678 4700 5742 4764
rect 5758 4700 5822 4764
rect 4713 4608 4777 4672
rect 4794 4608 4858 4672
rect 4875 4608 4939 4672
rect 4956 4608 5020 4672
rect 5037 4608 5101 4672
rect 5118 4608 5182 4672
rect 5198 4608 5262 4672
rect 5278 4608 5342 4672
rect 5358 4608 5422 4672
rect 5438 4608 5502 4672
rect 5518 4608 5582 4672
rect 5598 4608 5662 4672
rect 5678 4608 5742 4672
rect 5758 4608 5822 4672
rect 4713 4516 4777 4580
rect 4794 4516 4858 4580
rect 4875 4516 4939 4580
rect 4956 4516 5020 4580
rect 5037 4516 5101 4580
rect 5118 4516 5182 4580
rect 5198 4516 5262 4580
rect 5278 4516 5342 4580
rect 5358 4516 5422 4580
rect 5438 4516 5502 4580
rect 5518 4516 5582 4580
rect 5598 4516 5662 4580
rect 5678 4516 5742 4580
rect 5758 4516 5822 4580
rect 4713 4424 4777 4488
rect 4794 4424 4858 4488
rect 4875 4424 4939 4488
rect 4956 4424 5020 4488
rect 5037 4424 5101 4488
rect 5118 4424 5182 4488
rect 5198 4424 5262 4488
rect 5278 4424 5342 4488
rect 5358 4424 5422 4488
rect 5438 4424 5502 4488
rect 5518 4424 5582 4488
rect 5598 4424 5662 4488
rect 5678 4424 5742 4488
rect 5758 4424 5822 4488
rect 4713 4332 4777 4396
rect 4794 4332 4858 4396
rect 4875 4332 4939 4396
rect 4956 4332 5020 4396
rect 5037 4332 5101 4396
rect 5118 4332 5182 4396
rect 5198 4332 5262 4396
rect 5278 4332 5342 4396
rect 5358 4332 5422 4396
rect 5438 4332 5502 4396
rect 5518 4332 5582 4396
rect 5598 4332 5662 4396
rect 5678 4332 5742 4396
rect 5758 4332 5822 4396
rect 7531 4792 7595 4856
rect 7617 4792 7681 4856
rect 7703 4792 7767 4856
rect 7789 4792 7853 4856
rect 7875 4792 7939 4856
rect 7961 4792 8025 4856
rect 8047 4792 8111 4856
rect 8133 4792 8197 4856
rect 8219 4792 8283 4856
rect 8305 4792 8369 4856
rect 8391 4792 8455 4856
rect 8477 4792 8541 4856
rect 8563 4792 8627 4856
rect 8648 4792 8712 4856
rect 7531 4700 7595 4764
rect 7617 4700 7681 4764
rect 7703 4700 7767 4764
rect 7789 4700 7853 4764
rect 7875 4700 7939 4764
rect 7961 4700 8025 4764
rect 8047 4700 8111 4764
rect 8133 4700 8197 4764
rect 8219 4700 8283 4764
rect 8305 4700 8369 4764
rect 8391 4700 8455 4764
rect 8477 4700 8541 4764
rect 8563 4700 8627 4764
rect 8648 4700 8712 4764
rect 7531 4608 7595 4672
rect 7617 4608 7681 4672
rect 7703 4608 7767 4672
rect 7789 4608 7853 4672
rect 7875 4608 7939 4672
rect 7961 4608 8025 4672
rect 8047 4608 8111 4672
rect 8133 4608 8197 4672
rect 8219 4608 8283 4672
rect 8305 4608 8369 4672
rect 8391 4608 8455 4672
rect 8477 4608 8541 4672
rect 8563 4608 8627 4672
rect 8648 4608 8712 4672
rect 7531 4516 7595 4580
rect 7617 4516 7681 4580
rect 7703 4516 7767 4580
rect 7789 4516 7853 4580
rect 7875 4516 7939 4580
rect 7961 4516 8025 4580
rect 8047 4516 8111 4580
rect 8133 4516 8197 4580
rect 8219 4516 8283 4580
rect 8305 4516 8369 4580
rect 8391 4516 8455 4580
rect 8477 4516 8541 4580
rect 8563 4516 8627 4580
rect 8648 4516 8712 4580
rect 7531 4424 7595 4488
rect 7617 4424 7681 4488
rect 7703 4424 7767 4488
rect 7789 4424 7853 4488
rect 7875 4424 7939 4488
rect 7961 4424 8025 4488
rect 8047 4424 8111 4488
rect 8133 4424 8197 4488
rect 8219 4424 8283 4488
rect 8305 4424 8369 4488
rect 8391 4424 8455 4488
rect 8477 4424 8541 4488
rect 8563 4424 8627 4488
rect 8648 4424 8712 4488
rect 3924 858 4788 2352
rect 3924 802 3972 858
rect 3972 802 3998 858
rect 3998 802 4054 858
rect 4054 802 4080 858
rect 4080 802 4136 858
rect 4136 802 4162 858
rect 4162 802 4218 858
rect 4218 802 4244 858
rect 4244 802 4300 858
rect 4300 802 4326 858
rect 4326 802 4382 858
rect 4382 802 4408 858
rect 4408 802 4464 858
rect 4464 802 4490 858
rect 4490 802 4546 858
rect 4546 802 4573 858
rect 4573 802 4629 858
rect 4629 802 4656 858
rect 4656 802 4712 858
rect 4712 802 4739 858
rect 4739 802 4788 858
rect 3924 724 4788 802
rect 3924 668 3972 724
rect 3972 668 3998 724
rect 3998 668 4054 724
rect 4054 668 4080 724
rect 4080 668 4136 724
rect 4136 668 4162 724
rect 4162 668 4218 724
rect 4218 668 4244 724
rect 4244 668 4300 724
rect 4300 668 4326 724
rect 4326 668 4382 724
rect 4382 668 4408 724
rect 4408 668 4464 724
rect 4464 668 4490 724
rect 4490 668 4546 724
rect 4546 668 4573 724
rect 4573 668 4629 724
rect 4629 668 4656 724
rect 4656 668 4712 724
rect 4712 668 4739 724
rect 4739 668 4788 724
rect 3924 39 4788 668
rect 3924 -17 3972 39
rect 3972 -17 3998 39
rect 3998 -17 4054 39
rect 4054 -17 4080 39
rect 4080 -17 4136 39
rect 4136 -17 4162 39
rect 4162 -17 4218 39
rect 4218 -17 4244 39
rect 4244 -17 4300 39
rect 4300 -17 4326 39
rect 4326 -17 4382 39
rect 4382 -17 4408 39
rect 4408 -17 4464 39
rect 4464 -17 4490 39
rect 4490 -17 4546 39
rect 4546 -17 4573 39
rect 4573 -17 4629 39
rect 4629 -17 4656 39
rect 4656 -17 4712 39
rect 4712 -17 4739 39
rect 4739 -17 4788 39
rect 3924 -95 4788 -17
rect 3924 -151 3972 -95
rect 3972 -151 3998 -95
rect 3998 -151 4054 -95
rect 4054 -151 4080 -95
rect 4080 -151 4136 -95
rect 4136 -151 4162 -95
rect 4162 -151 4218 -95
rect 4218 -151 4244 -95
rect 4244 -151 4300 -95
rect 4300 -151 4326 -95
rect 4326 -151 4382 -95
rect 4382 -151 4408 -95
rect 4408 -151 4464 -95
rect 4464 -151 4490 -95
rect 4490 -151 4546 -95
rect 4546 -151 4573 -95
rect 4573 -151 4629 -95
rect 4629 -151 4656 -95
rect 4656 -151 4712 -95
rect 4712 -151 4739 -95
rect 4739 -151 4788 -95
rect 3924 -832 4788 -151
rect 3924 -913 3988 -849
rect 4004 -913 4068 -849
rect 4084 -913 4148 -849
rect 4164 -913 4228 -849
rect 4244 -913 4308 -849
rect 4324 -913 4388 -849
rect 4404 -913 4468 -849
rect 4484 -913 4548 -849
rect 4564 -913 4628 -849
rect 4644 -913 4708 -849
rect 4724 -913 4788 -849
rect 3924 -994 3988 -930
rect 4004 -994 4068 -930
rect 4084 -994 4148 -930
rect 4164 -994 4228 -930
rect 4244 -994 4308 -930
rect 4324 -994 4388 -930
rect 4404 -994 4468 -930
rect 4484 -994 4548 -930
rect 4564 -994 4628 -930
rect 4644 -994 4708 -930
rect 4724 -994 4788 -930
rect 3924 -1075 3988 -1011
rect 4004 -1075 4068 -1011
rect 4084 -1075 4148 -1011
rect 4164 -1075 4228 -1011
rect 4244 -1075 4308 -1011
rect 4324 -1075 4388 -1011
rect 4404 -1075 4468 -1011
rect 4484 -1075 4548 -1011
rect 4564 -1075 4628 -1011
rect 4644 -1075 4708 -1011
rect 4724 -1075 4788 -1011
rect 3924 -1156 3988 -1092
rect 4004 -1156 4068 -1092
rect 4084 -1156 4148 -1092
rect 4164 -1156 4228 -1092
rect 4244 -1156 4308 -1092
rect 4324 -1156 4388 -1092
rect 4404 -1156 4468 -1092
rect 4484 -1156 4548 -1092
rect 4564 -1156 4628 -1092
rect 4644 -1156 4708 -1092
rect 4724 -1156 4788 -1092
rect 3924 -1237 3988 -1173
rect 4004 -1237 4068 -1173
rect 4084 -1237 4148 -1173
rect 4164 -1237 4228 -1173
rect 4244 -1237 4308 -1173
rect 4324 -1237 4388 -1173
rect 4404 -1237 4468 -1173
rect 4484 -1237 4548 -1173
rect 4564 -1237 4628 -1173
rect 4644 -1237 4708 -1173
rect 4724 -1237 4788 -1173
rect 3924 -1318 3988 -1254
rect 4004 -1318 4068 -1254
rect 4084 -1318 4148 -1254
rect 4164 -1318 4228 -1254
rect 4244 -1318 4308 -1254
rect 4324 -1318 4388 -1254
rect 4404 -1318 4468 -1254
rect 4484 -1318 4548 -1254
rect 4564 -1318 4628 -1254
rect 4644 -1318 4708 -1254
rect 4724 -1318 4788 -1254
rect 3924 -1399 3988 -1335
rect 4004 -1399 4068 -1335
rect 4084 -1399 4148 -1335
rect 4164 -1399 4228 -1335
rect 4244 -1399 4308 -1335
rect 4324 -1399 4388 -1335
rect 4404 -1399 4468 -1335
rect 4484 -1399 4548 -1335
rect 4564 -1399 4628 -1335
rect 4644 -1399 4708 -1335
rect 4724 -1399 4788 -1335
rect 3924 -1480 3988 -1416
rect 4004 -1480 4068 -1416
rect 4084 -1480 4148 -1416
rect 4164 -1480 4228 -1416
rect 4244 -1480 4308 -1416
rect 4324 -1480 4388 -1416
rect 4404 -1480 4468 -1416
rect 4484 -1480 4548 -1416
rect 4564 -1480 4628 -1416
rect 4644 -1480 4708 -1416
rect 4724 -1480 4788 -1416
rect 3924 -1561 3988 -1497
rect 4004 -1561 4068 -1497
rect 4084 -1561 4148 -1497
rect 4164 -1561 4228 -1497
rect 4244 -1561 4308 -1497
rect 4324 -1561 4388 -1497
rect 4404 -1561 4468 -1497
rect 4484 -1561 4548 -1497
rect 4564 -1561 4628 -1497
rect 4644 -1561 4708 -1497
rect 4724 -1561 4788 -1497
rect 3924 -1642 3988 -1578
rect 4004 -1642 4068 -1578
rect 4084 -1642 4148 -1578
rect 4164 -1642 4228 -1578
rect 4244 -1642 4308 -1578
rect 4324 -1642 4388 -1578
rect 4404 -1642 4468 -1578
rect 4484 -1642 4548 -1578
rect 4564 -1642 4628 -1578
rect 4644 -1642 4708 -1578
rect 4724 -1642 4788 -1578
rect 3924 -1723 3988 -1659
rect 4004 -1723 4068 -1659
rect 4084 -1723 4148 -1659
rect 4164 -1723 4228 -1659
rect 4244 -1723 4308 -1659
rect 4324 -1723 4388 -1659
rect 4404 -1723 4468 -1659
rect 4484 -1723 4548 -1659
rect 4564 -1723 4628 -1659
rect 4644 -1723 4708 -1659
rect 4724 -1723 4788 -1659
rect 3924 -1804 3988 -1740
rect 4004 -1804 4068 -1740
rect 4084 -1804 4148 -1740
rect 4164 -1804 4228 -1740
rect 4244 -1804 4308 -1740
rect 4324 -1804 4388 -1740
rect 4404 -1804 4468 -1740
rect 4484 -1804 4548 -1740
rect 4564 -1804 4628 -1740
rect 4644 -1804 4708 -1740
rect 4724 -1804 4788 -1740
rect 3924 -1885 3988 -1821
rect 4004 -1885 4068 -1821
rect 4084 -1885 4148 -1821
rect 4164 -1885 4228 -1821
rect 4244 -1885 4308 -1821
rect 4324 -1885 4388 -1821
rect 4404 -1885 4468 -1821
rect 4484 -1885 4548 -1821
rect 4564 -1885 4628 -1821
rect 4644 -1885 4708 -1821
rect 4724 -1885 4788 -1821
rect 3924 -1966 3988 -1902
rect 4004 -1966 4068 -1902
rect 4084 -1966 4148 -1902
rect 4164 -1966 4228 -1902
rect 4244 -1966 4308 -1902
rect 4324 -1966 4388 -1902
rect 4404 -1966 4468 -1902
rect 4484 -1966 4548 -1902
rect 4564 -1966 4628 -1902
rect 4644 -1966 4708 -1902
rect 4724 -1966 4788 -1902
rect 3924 -2047 3988 -1983
rect 4004 -2047 4068 -1983
rect 4084 -2047 4148 -1983
rect 4164 -2047 4228 -1983
rect 4244 -2047 4308 -1983
rect 4324 -2047 4388 -1983
rect 4404 -2047 4468 -1983
rect 4484 -2047 4548 -1983
rect 4564 -2047 4628 -1983
rect 4644 -2047 4708 -1983
rect 4724 -2047 4788 -1983
rect 3924 -2128 3988 -2064
rect 4004 -2128 4068 -2064
rect 4084 -2128 4148 -2064
rect 4164 -2128 4228 -2064
rect 4244 -2128 4308 -2064
rect 4324 -2128 4388 -2064
rect 4404 -2128 4468 -2064
rect 4484 -2128 4548 -2064
rect 4564 -2128 4628 -2064
rect 4644 -2128 4708 -2064
rect 4724 -2128 4788 -2064
rect 3924 -2209 3988 -2145
rect 4004 -2209 4068 -2145
rect 4084 -2209 4148 -2145
rect 4164 -2209 4228 -2145
rect 4244 -2209 4308 -2145
rect 4324 -2209 4388 -2145
rect 4404 -2209 4468 -2145
rect 4484 -2209 4548 -2145
rect 4564 -2209 4628 -2145
rect 4644 -2209 4708 -2145
rect 4724 -2209 4788 -2145
rect 3924 -2290 3988 -2226
rect 4004 -2290 4068 -2226
rect 4084 -2290 4148 -2226
rect 4164 -2290 4228 -2226
rect 4244 -2290 4308 -2226
rect 4324 -2290 4388 -2226
rect 4404 -2290 4468 -2226
rect 4484 -2290 4548 -2226
rect 4564 -2290 4628 -2226
rect 4644 -2290 4708 -2226
rect 4724 -2290 4788 -2226
rect 3924 -2371 3988 -2307
rect 4004 -2371 4068 -2307
rect 4084 -2371 4148 -2307
rect 4164 -2371 4228 -2307
rect 4244 -2371 4308 -2307
rect 4324 -2371 4388 -2307
rect 4404 -2371 4468 -2307
rect 4484 -2371 4548 -2307
rect 4564 -2371 4628 -2307
rect 4644 -2371 4708 -2307
rect 4724 -2371 4788 -2307
rect 3924 -2452 3988 -2388
rect 4004 -2452 4068 -2388
rect 4084 -2452 4148 -2388
rect 4164 -2452 4228 -2388
rect 4244 -2452 4308 -2388
rect 4324 -2452 4388 -2388
rect 4404 -2452 4468 -2388
rect 4484 -2452 4548 -2388
rect 4564 -2452 4628 -2388
rect 4644 -2452 4708 -2388
rect 4724 -2452 4788 -2388
rect 3924 -2533 3988 -2469
rect 4004 -2533 4068 -2469
rect 4084 -2533 4148 -2469
rect 4164 -2533 4228 -2469
rect 4244 -2533 4308 -2469
rect 4324 -2533 4388 -2469
rect 4404 -2533 4468 -2469
rect 4484 -2533 4548 -2469
rect 4564 -2533 4628 -2469
rect 4644 -2533 4708 -2469
rect 4724 -2533 4788 -2469
rect 3924 -2614 3988 -2550
rect 4004 -2614 4068 -2550
rect 4084 -2614 4148 -2550
rect 4164 -2614 4228 -2550
rect 4244 -2614 4308 -2550
rect 4324 -2614 4388 -2550
rect 4404 -2614 4468 -2550
rect 4484 -2614 4548 -2550
rect 4564 -2614 4628 -2550
rect 4644 -2614 4708 -2550
rect 4724 -2614 4788 -2550
rect 4883 -3000 4947 -2936
rect 4963 -3000 5027 -2936
rect 5043 -3000 5107 -2936
rect 4883 -3091 4947 -3027
rect 4963 -3091 5027 -3027
rect 5043 -3091 5107 -3027
rect 4883 -3183 4947 -3119
rect 4963 -3183 5027 -3119
rect 5043 -3183 5107 -3119
rect 4883 -3275 4947 -3211
rect 4963 -3275 5027 -3211
rect 5043 -3275 5107 -3211
rect 5717 -3000 5781 -2936
rect 5797 -3000 5861 -2936
rect 5877 -3000 5941 -2936
rect 5717 -3091 5781 -3027
rect 5797 -3091 5861 -3027
rect 5877 -3091 5941 -3027
rect 5717 -3183 5781 -3119
rect 5797 -3183 5861 -3119
rect 5877 -3183 5941 -3119
rect 5717 -3275 5781 -3211
rect 5797 -3275 5861 -3211
rect 5877 -3275 5941 -3211
rect 7531 4332 7595 4396
rect 7617 4332 7681 4396
rect 7703 4332 7767 4396
rect 7789 4332 7853 4396
rect 7875 4332 7939 4396
rect 7961 4332 8025 4396
rect 8047 4332 8111 4396
rect 8133 4332 8197 4396
rect 8219 4332 8283 4396
rect 8305 4332 8369 4396
rect 8391 4332 8455 4396
rect 8477 4332 8541 4396
rect 8563 4332 8627 4396
rect 8648 4332 8712 4396
rect 8568 858 9432 2352
rect 8568 802 8615 858
rect 8615 802 8642 858
rect 8642 802 8698 858
rect 8698 802 8725 858
rect 8725 802 8781 858
rect 8781 802 8808 858
rect 8808 802 8864 858
rect 8864 802 8890 858
rect 8890 802 8946 858
rect 8946 802 8972 858
rect 8972 802 9028 858
rect 9028 802 9054 858
rect 9054 802 9110 858
rect 9110 802 9136 858
rect 9136 802 9192 858
rect 9192 802 9218 858
rect 9218 802 9274 858
rect 9274 802 9300 858
rect 9300 802 9356 858
rect 9356 802 9382 858
rect 9382 802 9432 858
rect 8568 724 9432 802
rect 8568 668 8615 724
rect 8615 668 8642 724
rect 8642 668 8698 724
rect 8698 668 8725 724
rect 8725 668 8781 724
rect 8781 668 8808 724
rect 8808 668 8864 724
rect 8864 668 8890 724
rect 8890 668 8946 724
rect 8946 668 8972 724
rect 8972 668 9028 724
rect 9028 668 9054 724
rect 9054 668 9110 724
rect 9110 668 9136 724
rect 9136 668 9192 724
rect 9192 668 9218 724
rect 9218 668 9274 724
rect 9274 668 9300 724
rect 9300 668 9356 724
rect 9356 668 9382 724
rect 9382 668 9432 724
rect 8568 35 9432 668
rect 8568 -21 8615 35
rect 8615 -21 8642 35
rect 8642 -21 8698 35
rect 8698 -21 8725 35
rect 8725 -21 8781 35
rect 8781 -21 8808 35
rect 8808 -21 8864 35
rect 8864 -21 8890 35
rect 8890 -21 8946 35
rect 8946 -21 8972 35
rect 8972 -21 9028 35
rect 9028 -21 9054 35
rect 9054 -21 9110 35
rect 9110 -21 9136 35
rect 9136 -21 9192 35
rect 9192 -21 9218 35
rect 9218 -21 9274 35
rect 9274 -21 9300 35
rect 9300 -21 9356 35
rect 9356 -21 9382 35
rect 9382 -21 9432 35
rect 8568 -99 9432 -21
rect 8568 -155 8615 -99
rect 8615 -155 8642 -99
rect 8642 -155 8698 -99
rect 8698 -155 8725 -99
rect 8725 -155 8781 -99
rect 8781 -155 8808 -99
rect 8808 -155 8864 -99
rect 8864 -155 8890 -99
rect 8890 -155 8946 -99
rect 8946 -155 8972 -99
rect 8972 -155 9028 -99
rect 9028 -155 9054 -99
rect 9054 -155 9110 -99
rect 9110 -155 9136 -99
rect 9136 -155 9192 -99
rect 9192 -155 9218 -99
rect 9218 -155 9274 -99
rect 9274 -155 9300 -99
rect 9300 -155 9356 -99
rect 9356 -155 9382 -99
rect 9382 -155 9432 -99
rect 8568 -832 9432 -155
rect 8568 -913 8632 -849
rect 8648 -913 8712 -849
rect 8728 -913 8792 -849
rect 8808 -913 8872 -849
rect 8888 -913 8952 -849
rect 8968 -913 9032 -849
rect 9048 -913 9112 -849
rect 9128 -913 9192 -849
rect 9208 -913 9272 -849
rect 9288 -913 9352 -849
rect 9368 -913 9432 -849
rect 8568 -994 8632 -930
rect 8648 -994 8712 -930
rect 8728 -994 8792 -930
rect 8808 -994 8872 -930
rect 8888 -994 8952 -930
rect 8968 -994 9032 -930
rect 9048 -994 9112 -930
rect 9128 -994 9192 -930
rect 9208 -994 9272 -930
rect 9288 -994 9352 -930
rect 9368 -994 9432 -930
rect 8568 -1075 8632 -1011
rect 8648 -1075 8712 -1011
rect 8728 -1075 8792 -1011
rect 8808 -1075 8872 -1011
rect 8888 -1075 8952 -1011
rect 8968 -1075 9032 -1011
rect 9048 -1075 9112 -1011
rect 9128 -1075 9192 -1011
rect 9208 -1075 9272 -1011
rect 9288 -1075 9352 -1011
rect 9368 -1075 9432 -1011
rect 8568 -1156 8632 -1092
rect 8648 -1156 8712 -1092
rect 8728 -1156 8792 -1092
rect 8808 -1156 8872 -1092
rect 8888 -1156 8952 -1092
rect 8968 -1156 9032 -1092
rect 9048 -1156 9112 -1092
rect 9128 -1156 9192 -1092
rect 9208 -1156 9272 -1092
rect 9288 -1156 9352 -1092
rect 9368 -1156 9432 -1092
rect 8568 -1237 8632 -1173
rect 8648 -1237 8712 -1173
rect 8728 -1237 8792 -1173
rect 8808 -1237 8872 -1173
rect 8888 -1237 8952 -1173
rect 8968 -1237 9032 -1173
rect 9048 -1237 9112 -1173
rect 9128 -1237 9192 -1173
rect 9208 -1237 9272 -1173
rect 9288 -1237 9352 -1173
rect 9368 -1237 9432 -1173
rect 8568 -1318 8632 -1254
rect 8648 -1318 8712 -1254
rect 8728 -1318 8792 -1254
rect 8808 -1318 8872 -1254
rect 8888 -1318 8952 -1254
rect 8968 -1318 9032 -1254
rect 9048 -1318 9112 -1254
rect 9128 -1318 9192 -1254
rect 9208 -1318 9272 -1254
rect 9288 -1318 9352 -1254
rect 9368 -1318 9432 -1254
rect 8568 -1399 8632 -1335
rect 8648 -1399 8712 -1335
rect 8728 -1399 8792 -1335
rect 8808 -1399 8872 -1335
rect 8888 -1399 8952 -1335
rect 8968 -1399 9032 -1335
rect 9048 -1399 9112 -1335
rect 9128 -1399 9192 -1335
rect 9208 -1399 9272 -1335
rect 9288 -1399 9352 -1335
rect 9368 -1399 9432 -1335
rect 8568 -1480 8632 -1416
rect 8648 -1480 8712 -1416
rect 8728 -1480 8792 -1416
rect 8808 -1480 8872 -1416
rect 8888 -1480 8952 -1416
rect 8968 -1480 9032 -1416
rect 9048 -1480 9112 -1416
rect 9128 -1480 9192 -1416
rect 9208 -1480 9272 -1416
rect 9288 -1480 9352 -1416
rect 9368 -1480 9432 -1416
rect 8568 -1561 8632 -1497
rect 8648 -1561 8712 -1497
rect 8728 -1561 8792 -1497
rect 8808 -1561 8872 -1497
rect 8888 -1561 8952 -1497
rect 8968 -1561 9032 -1497
rect 9048 -1561 9112 -1497
rect 9128 -1561 9192 -1497
rect 9208 -1561 9272 -1497
rect 9288 -1561 9352 -1497
rect 9368 -1561 9432 -1497
rect 8568 -1642 8632 -1578
rect 8648 -1642 8712 -1578
rect 8728 -1642 8792 -1578
rect 8808 -1642 8872 -1578
rect 8888 -1642 8952 -1578
rect 8968 -1642 9032 -1578
rect 9048 -1642 9112 -1578
rect 9128 -1642 9192 -1578
rect 9208 -1642 9272 -1578
rect 9288 -1642 9352 -1578
rect 9368 -1642 9432 -1578
rect 8568 -1723 8632 -1659
rect 8648 -1723 8712 -1659
rect 8728 -1723 8792 -1659
rect 8808 -1723 8872 -1659
rect 8888 -1723 8952 -1659
rect 8968 -1723 9032 -1659
rect 9048 -1723 9112 -1659
rect 9128 -1723 9192 -1659
rect 9208 -1723 9272 -1659
rect 9288 -1723 9352 -1659
rect 9368 -1723 9432 -1659
rect 8568 -1804 8632 -1740
rect 8648 -1804 8712 -1740
rect 8728 -1804 8792 -1740
rect 8808 -1804 8872 -1740
rect 8888 -1804 8952 -1740
rect 8968 -1804 9032 -1740
rect 9048 -1804 9112 -1740
rect 9128 -1804 9192 -1740
rect 9208 -1804 9272 -1740
rect 9288 -1804 9352 -1740
rect 9368 -1804 9432 -1740
rect 8568 -1885 8632 -1821
rect 8648 -1885 8712 -1821
rect 8728 -1885 8792 -1821
rect 8808 -1885 8872 -1821
rect 8888 -1885 8952 -1821
rect 8968 -1885 9032 -1821
rect 9048 -1885 9112 -1821
rect 9128 -1885 9192 -1821
rect 9208 -1885 9272 -1821
rect 9288 -1885 9352 -1821
rect 9368 -1885 9432 -1821
rect 8568 -1966 8632 -1902
rect 8648 -1966 8712 -1902
rect 8728 -1966 8792 -1902
rect 8808 -1966 8872 -1902
rect 8888 -1966 8952 -1902
rect 8968 -1966 9032 -1902
rect 9048 -1966 9112 -1902
rect 9128 -1966 9192 -1902
rect 9208 -1966 9272 -1902
rect 9288 -1966 9352 -1902
rect 9368 -1966 9432 -1902
rect 8568 -2047 8632 -1983
rect 8648 -2047 8712 -1983
rect 8728 -2047 8792 -1983
rect 8808 -2047 8872 -1983
rect 8888 -2047 8952 -1983
rect 8968 -2047 9032 -1983
rect 9048 -2047 9112 -1983
rect 9128 -2047 9192 -1983
rect 9208 -2047 9272 -1983
rect 9288 -2047 9352 -1983
rect 9368 -2047 9432 -1983
rect 8568 -2128 8632 -2064
rect 8648 -2128 8712 -2064
rect 8728 -2128 8792 -2064
rect 8808 -2128 8872 -2064
rect 8888 -2128 8952 -2064
rect 8968 -2128 9032 -2064
rect 9048 -2128 9112 -2064
rect 9128 -2128 9192 -2064
rect 9208 -2128 9272 -2064
rect 9288 -2128 9352 -2064
rect 9368 -2128 9432 -2064
rect 8568 -2209 8632 -2145
rect 8648 -2209 8712 -2145
rect 8728 -2209 8792 -2145
rect 8808 -2209 8872 -2145
rect 8888 -2209 8952 -2145
rect 8968 -2209 9032 -2145
rect 9048 -2209 9112 -2145
rect 9128 -2209 9192 -2145
rect 9208 -2209 9272 -2145
rect 9288 -2209 9352 -2145
rect 9368 -2209 9432 -2145
rect 8568 -2290 8632 -2226
rect 8648 -2290 8712 -2226
rect 8728 -2290 8792 -2226
rect 8808 -2290 8872 -2226
rect 8888 -2290 8952 -2226
rect 8968 -2290 9032 -2226
rect 9048 -2290 9112 -2226
rect 9128 -2290 9192 -2226
rect 9208 -2290 9272 -2226
rect 9288 -2290 9352 -2226
rect 9368 -2290 9432 -2226
rect 8568 -2371 8632 -2307
rect 8648 -2371 8712 -2307
rect 8728 -2371 8792 -2307
rect 8808 -2371 8872 -2307
rect 8888 -2371 8952 -2307
rect 8968 -2371 9032 -2307
rect 9048 -2371 9112 -2307
rect 9128 -2371 9192 -2307
rect 9208 -2371 9272 -2307
rect 9288 -2371 9352 -2307
rect 9368 -2371 9432 -2307
rect 8568 -2452 8632 -2388
rect 8648 -2452 8712 -2388
rect 8728 -2452 8792 -2388
rect 8808 -2452 8872 -2388
rect 8888 -2452 8952 -2388
rect 8968 -2452 9032 -2388
rect 9048 -2452 9112 -2388
rect 9128 -2452 9192 -2388
rect 9208 -2452 9272 -2388
rect 9288 -2452 9352 -2388
rect 9368 -2452 9432 -2388
rect 8568 -2533 8632 -2469
rect 8648 -2533 8712 -2469
rect 8728 -2533 8792 -2469
rect 8808 -2533 8872 -2469
rect 8888 -2533 8952 -2469
rect 8968 -2533 9032 -2469
rect 9048 -2533 9112 -2469
rect 9128 -2533 9192 -2469
rect 9208 -2533 9272 -2469
rect 9288 -2533 9352 -2469
rect 9368 -2533 9432 -2469
rect 8568 -2614 8632 -2550
rect 8648 -2614 8712 -2550
rect 8728 -2614 8792 -2550
rect 8808 -2614 8872 -2550
rect 8888 -2614 8952 -2550
rect 8968 -2614 9032 -2550
rect 9048 -2614 9112 -2550
rect 9128 -2614 9192 -2550
rect 9208 -2614 9272 -2550
rect 9288 -2614 9352 -2550
rect 9368 -2614 9432 -2550
rect 6492 -3000 6556 -2936
rect 6594 -3000 6658 -2936
rect 6696 -3000 6760 -2936
rect 6798 -3000 6862 -2936
rect 6492 -3080 6556 -3016
rect 6594 -3080 6658 -3016
rect 6696 -3080 6760 -3016
rect 6798 -3080 6862 -3016
rect 6492 -3160 6556 -3096
rect 6594 -3160 6658 -3096
rect 6696 -3160 6760 -3096
rect 6798 -3160 6862 -3096
rect 6492 -3240 6556 -3176
rect 6594 -3240 6658 -3176
rect 6696 -3240 6760 -3176
rect 6798 -3240 6862 -3176
rect 6492 -3320 6556 -3256
rect 6594 -3320 6658 -3256
rect 6696 -3320 6760 -3256
rect 6798 -3320 6862 -3256
rect 6492 -3401 6556 -3337
rect 6594 -3401 6658 -3337
rect 6696 -3401 6760 -3337
rect 6798 -3401 6862 -3337
rect 6492 -3482 6556 -3418
rect 6594 -3482 6658 -3418
rect 6696 -3482 6760 -3418
rect 6798 -3482 6862 -3418
rect 6492 -3563 6556 -3499
rect 6594 -3563 6658 -3499
rect 6696 -3563 6760 -3499
rect 6798 -3563 6862 -3499
rect 6492 -3644 6556 -3580
rect 6594 -3644 6658 -3580
rect 6696 -3644 6760 -3580
rect 6798 -3644 6862 -3580
rect 6492 -3725 6556 -3661
rect 6594 -3725 6658 -3661
rect 6696 -3725 6760 -3661
rect 6798 -3725 6862 -3661
rect 10407 858 11271 2352
rect 10407 802 10456 858
rect 10456 802 10482 858
rect 10482 802 10538 858
rect 10538 802 10564 858
rect 10564 802 10620 858
rect 10620 802 10646 858
rect 10646 802 10702 858
rect 10702 802 10728 858
rect 10728 802 10784 858
rect 10784 802 10810 858
rect 10810 802 10866 858
rect 10866 802 10892 858
rect 10892 802 10948 858
rect 10948 802 10974 858
rect 10974 802 11030 858
rect 11030 802 11057 858
rect 11057 802 11113 858
rect 11113 802 11140 858
rect 11140 802 11196 858
rect 11196 802 11223 858
rect 11223 802 11271 858
rect 10407 724 11271 802
rect 10407 668 10456 724
rect 10456 668 10482 724
rect 10482 668 10538 724
rect 10538 668 10564 724
rect 10564 668 10620 724
rect 10620 668 10646 724
rect 10646 668 10702 724
rect 10702 668 10728 724
rect 10728 668 10784 724
rect 10784 668 10810 724
rect 10810 668 10866 724
rect 10866 668 10892 724
rect 10892 668 10948 724
rect 10948 668 10974 724
rect 10974 668 11030 724
rect 11030 668 11057 724
rect 11057 668 11113 724
rect 11113 668 11140 724
rect 11140 668 11196 724
rect 11196 668 11223 724
rect 11223 668 11271 724
rect 10407 35 11271 668
rect 11453 4792 11517 4856
rect 11541 4792 11605 4856
rect 11629 4792 11693 4856
rect 11717 4792 11781 4856
rect 11805 4792 11869 4856
rect 11893 4792 11957 4856
rect 11981 4792 12045 4856
rect 12068 4792 12132 4856
rect 12155 4792 12219 4856
rect 12242 4792 12306 4856
rect 11453 4700 11517 4764
rect 11541 4700 11605 4764
rect 11629 4700 11693 4764
rect 11717 4700 11781 4764
rect 11805 4700 11869 4764
rect 11893 4700 11957 4764
rect 11981 4700 12045 4764
rect 12068 4700 12132 4764
rect 12155 4700 12219 4764
rect 12242 4700 12306 4764
rect 11453 4608 11517 4672
rect 11541 4608 11605 4672
rect 11629 4608 11693 4672
rect 11717 4608 11781 4672
rect 11805 4608 11869 4672
rect 11893 4608 11957 4672
rect 11981 4608 12045 4672
rect 12068 4608 12132 4672
rect 12155 4608 12219 4672
rect 12242 4608 12306 4672
rect 11453 4516 11517 4580
rect 11541 4516 11605 4580
rect 11629 4516 11693 4580
rect 11717 4516 11781 4580
rect 11805 4516 11869 4580
rect 11893 4516 11957 4580
rect 11981 4516 12045 4580
rect 12068 4516 12132 4580
rect 12155 4516 12219 4580
rect 12242 4516 12306 4580
rect 11453 4424 11517 4488
rect 11541 4424 11605 4488
rect 11629 4424 11693 4488
rect 11717 4424 11781 4488
rect 11805 4424 11869 4488
rect 11893 4424 11957 4488
rect 11981 4424 12045 4488
rect 12068 4424 12132 4488
rect 12155 4424 12219 4488
rect 12242 4424 12306 4488
rect 11453 4332 11517 4396
rect 11541 4332 11605 4396
rect 11629 4332 11693 4396
rect 11717 4332 11781 4396
rect 11805 4332 11869 4396
rect 11893 4332 11957 4396
rect 11981 4332 12045 4396
rect 12068 4332 12132 4396
rect 12155 4332 12219 4396
rect 12242 4332 12306 4396
rect 10407 -21 10456 35
rect 10456 -21 10482 35
rect 10482 -21 10538 35
rect 10538 -21 10564 35
rect 10564 -21 10620 35
rect 10620 -21 10646 35
rect 10646 -21 10702 35
rect 10702 -21 10728 35
rect 10728 -21 10784 35
rect 10784 -21 10810 35
rect 10810 -21 10866 35
rect 10866 -21 10892 35
rect 10892 -21 10948 35
rect 10948 -21 10974 35
rect 10974 -21 11030 35
rect 11030 -21 11057 35
rect 11057 -21 11113 35
rect 11113 -21 11140 35
rect 11140 -21 11196 35
rect 11196 -21 11223 35
rect 11223 -21 11271 35
rect 10407 -99 11271 -21
rect 10407 -155 10456 -99
rect 10456 -155 10482 -99
rect 10482 -155 10538 -99
rect 10538 -155 10564 -99
rect 10564 -155 10620 -99
rect 10620 -155 10646 -99
rect 10646 -155 10702 -99
rect 10702 -155 10728 -99
rect 10728 -155 10784 -99
rect 10784 -155 10810 -99
rect 10810 -155 10866 -99
rect 10866 -155 10892 -99
rect 10892 -155 10948 -99
rect 10948 -155 10974 -99
rect 10974 -155 11030 -99
rect 11030 -155 11057 -99
rect 11057 -155 11113 -99
rect 11113 -155 11140 -99
rect 11140 -155 11196 -99
rect 11196 -155 11223 -99
rect 11223 -155 11271 -99
rect 10407 -832 11271 -155
rect 10407 -913 10471 -849
rect 10487 -913 10551 -849
rect 10567 -913 10631 -849
rect 10647 -913 10711 -849
rect 10727 -913 10791 -849
rect 10807 -913 10871 -849
rect 10887 -913 10951 -849
rect 10967 -913 11031 -849
rect 11047 -913 11111 -849
rect 11127 -913 11191 -849
rect 11207 -913 11271 -849
rect 10407 -994 10471 -930
rect 10487 -994 10551 -930
rect 10567 -994 10631 -930
rect 10647 -994 10711 -930
rect 10727 -994 10791 -930
rect 10807 -994 10871 -930
rect 10887 -994 10951 -930
rect 10967 -994 11031 -930
rect 11047 -994 11111 -930
rect 11127 -994 11191 -930
rect 11207 -994 11271 -930
rect 10407 -1075 10471 -1011
rect 10487 -1075 10551 -1011
rect 10567 -1075 10631 -1011
rect 10647 -1075 10711 -1011
rect 10727 -1075 10791 -1011
rect 10807 -1075 10871 -1011
rect 10887 -1075 10951 -1011
rect 10967 -1075 11031 -1011
rect 11047 -1075 11111 -1011
rect 11127 -1075 11191 -1011
rect 11207 -1075 11271 -1011
rect 10407 -1156 10471 -1092
rect 10487 -1156 10551 -1092
rect 10567 -1156 10631 -1092
rect 10647 -1156 10711 -1092
rect 10727 -1156 10791 -1092
rect 10807 -1156 10871 -1092
rect 10887 -1156 10951 -1092
rect 10967 -1156 11031 -1092
rect 11047 -1156 11111 -1092
rect 11127 -1156 11191 -1092
rect 11207 -1156 11271 -1092
rect 10407 -1237 10471 -1173
rect 10487 -1237 10551 -1173
rect 10567 -1237 10631 -1173
rect 10647 -1237 10711 -1173
rect 10727 -1237 10791 -1173
rect 10807 -1237 10871 -1173
rect 10887 -1237 10951 -1173
rect 10967 -1237 11031 -1173
rect 11047 -1237 11111 -1173
rect 11127 -1237 11191 -1173
rect 11207 -1237 11271 -1173
rect 10407 -1318 10471 -1254
rect 10487 -1318 10551 -1254
rect 10567 -1318 10631 -1254
rect 10647 -1318 10711 -1254
rect 10727 -1318 10791 -1254
rect 10807 -1318 10871 -1254
rect 10887 -1318 10951 -1254
rect 10967 -1318 11031 -1254
rect 11047 -1318 11111 -1254
rect 11127 -1318 11191 -1254
rect 11207 -1318 11271 -1254
rect 10407 -1399 10471 -1335
rect 10487 -1399 10551 -1335
rect 10567 -1399 10631 -1335
rect 10647 -1399 10711 -1335
rect 10727 -1399 10791 -1335
rect 10807 -1399 10871 -1335
rect 10887 -1399 10951 -1335
rect 10967 -1399 11031 -1335
rect 11047 -1399 11111 -1335
rect 11127 -1399 11191 -1335
rect 11207 -1399 11271 -1335
rect 10407 -1480 10471 -1416
rect 10487 -1480 10551 -1416
rect 10567 -1480 10631 -1416
rect 10647 -1480 10711 -1416
rect 10727 -1480 10791 -1416
rect 10807 -1480 10871 -1416
rect 10887 -1480 10951 -1416
rect 10967 -1480 11031 -1416
rect 11047 -1480 11111 -1416
rect 11127 -1480 11191 -1416
rect 11207 -1480 11271 -1416
rect 10407 -1561 10471 -1497
rect 10487 -1561 10551 -1497
rect 10567 -1561 10631 -1497
rect 10647 -1561 10711 -1497
rect 10727 -1561 10791 -1497
rect 10807 -1561 10871 -1497
rect 10887 -1561 10951 -1497
rect 10967 -1561 11031 -1497
rect 11047 -1561 11111 -1497
rect 11127 -1561 11191 -1497
rect 11207 -1561 11271 -1497
rect 10407 -1642 10471 -1578
rect 10487 -1642 10551 -1578
rect 10567 -1642 10631 -1578
rect 10647 -1642 10711 -1578
rect 10727 -1642 10791 -1578
rect 10807 -1642 10871 -1578
rect 10887 -1642 10951 -1578
rect 10967 -1642 11031 -1578
rect 11047 -1642 11111 -1578
rect 11127 -1642 11191 -1578
rect 11207 -1642 11271 -1578
rect 10407 -1723 10471 -1659
rect 10487 -1723 10551 -1659
rect 10567 -1723 10631 -1659
rect 10647 -1723 10711 -1659
rect 10727 -1723 10791 -1659
rect 10807 -1723 10871 -1659
rect 10887 -1723 10951 -1659
rect 10967 -1723 11031 -1659
rect 11047 -1723 11111 -1659
rect 11127 -1723 11191 -1659
rect 11207 -1723 11271 -1659
rect 10407 -1804 10471 -1740
rect 10487 -1804 10551 -1740
rect 10567 -1804 10631 -1740
rect 10647 -1804 10711 -1740
rect 10727 -1804 10791 -1740
rect 10807 -1804 10871 -1740
rect 10887 -1804 10951 -1740
rect 10967 -1804 11031 -1740
rect 11047 -1804 11111 -1740
rect 11127 -1804 11191 -1740
rect 11207 -1804 11271 -1740
rect 10407 -1885 10471 -1821
rect 10487 -1885 10551 -1821
rect 10567 -1885 10631 -1821
rect 10647 -1885 10711 -1821
rect 10727 -1885 10791 -1821
rect 10807 -1885 10871 -1821
rect 10887 -1885 10951 -1821
rect 10967 -1885 11031 -1821
rect 11047 -1885 11111 -1821
rect 11127 -1885 11191 -1821
rect 11207 -1885 11271 -1821
rect 10407 -1966 10471 -1902
rect 10487 -1966 10551 -1902
rect 10567 -1966 10631 -1902
rect 10647 -1966 10711 -1902
rect 10727 -1966 10791 -1902
rect 10807 -1966 10871 -1902
rect 10887 -1966 10951 -1902
rect 10967 -1966 11031 -1902
rect 11047 -1966 11111 -1902
rect 11127 -1966 11191 -1902
rect 11207 -1966 11271 -1902
rect 10407 -2047 10471 -1983
rect 10487 -2047 10551 -1983
rect 10567 -2047 10631 -1983
rect 10647 -2047 10711 -1983
rect 10727 -2047 10791 -1983
rect 10807 -2047 10871 -1983
rect 10887 -2047 10951 -1983
rect 10967 -2047 11031 -1983
rect 11047 -2047 11111 -1983
rect 11127 -2047 11191 -1983
rect 11207 -2047 11271 -1983
rect 10407 -2128 10471 -2064
rect 10487 -2128 10551 -2064
rect 10567 -2128 10631 -2064
rect 10647 -2128 10711 -2064
rect 10727 -2128 10791 -2064
rect 10807 -2128 10871 -2064
rect 10887 -2128 10951 -2064
rect 10967 -2128 11031 -2064
rect 11047 -2128 11111 -2064
rect 11127 -2128 11191 -2064
rect 11207 -2128 11271 -2064
rect 10407 -2209 10471 -2145
rect 10487 -2209 10551 -2145
rect 10567 -2209 10631 -2145
rect 10647 -2209 10711 -2145
rect 10727 -2209 10791 -2145
rect 10807 -2209 10871 -2145
rect 10887 -2209 10951 -2145
rect 10967 -2209 11031 -2145
rect 11047 -2209 11111 -2145
rect 11127 -2209 11191 -2145
rect 11207 -2209 11271 -2145
rect 10407 -2290 10471 -2226
rect 10487 -2290 10551 -2226
rect 10567 -2290 10631 -2226
rect 10647 -2290 10711 -2226
rect 10727 -2290 10791 -2226
rect 10807 -2290 10871 -2226
rect 10887 -2290 10951 -2226
rect 10967 -2290 11031 -2226
rect 11047 -2290 11111 -2226
rect 11127 -2290 11191 -2226
rect 11207 -2290 11271 -2226
rect 10407 -2371 10471 -2307
rect 10487 -2371 10551 -2307
rect 10567 -2371 10631 -2307
rect 10647 -2371 10711 -2307
rect 10727 -2371 10791 -2307
rect 10807 -2371 10871 -2307
rect 10887 -2371 10951 -2307
rect 10967 -2371 11031 -2307
rect 11047 -2371 11111 -2307
rect 11127 -2371 11191 -2307
rect 11207 -2371 11271 -2307
rect 10407 -2452 10471 -2388
rect 10487 -2452 10551 -2388
rect 10567 -2452 10631 -2388
rect 10647 -2452 10711 -2388
rect 10727 -2452 10791 -2388
rect 10807 -2452 10871 -2388
rect 10887 -2452 10951 -2388
rect 10967 -2452 11031 -2388
rect 11047 -2452 11111 -2388
rect 11127 -2452 11191 -2388
rect 11207 -2452 11271 -2388
rect 10407 -2533 10471 -2469
rect 10487 -2533 10551 -2469
rect 10567 -2533 10631 -2469
rect 10647 -2533 10711 -2469
rect 10727 -2533 10791 -2469
rect 10807 -2533 10871 -2469
rect 10887 -2533 10951 -2469
rect 10967 -2533 11031 -2469
rect 11047 -2533 11111 -2469
rect 11127 -2533 11191 -2469
rect 11207 -2533 11271 -2469
rect 10407 -2614 10471 -2550
rect 10487 -2614 10551 -2550
rect 10567 -2614 10631 -2550
rect 10647 -2614 10711 -2550
rect 10727 -2614 10791 -2550
rect 10807 -2614 10871 -2550
rect 10887 -2614 10951 -2550
rect 10967 -2614 11031 -2550
rect 11047 -2614 11111 -2550
rect 11127 -2614 11191 -2550
rect 11207 -2614 11271 -2550
rect 14014 4362 14878 5226
rect 15052 858 15916 2352
rect 17934 4362 18798 5226
rect 15052 802 15099 858
rect 15099 802 15126 858
rect 15126 802 15182 858
rect 15182 802 15209 858
rect 15209 802 15265 858
rect 15265 802 15292 858
rect 15292 802 15348 858
rect 15348 802 15374 858
rect 15374 802 15430 858
rect 15430 802 15456 858
rect 15456 802 15512 858
rect 15512 802 15538 858
rect 15538 802 15594 858
rect 15594 802 15620 858
rect 15620 802 15676 858
rect 15676 802 15702 858
rect 15702 802 15758 858
rect 15758 802 15784 858
rect 15784 802 15840 858
rect 15840 802 15866 858
rect 15866 802 15916 858
rect 15052 724 15916 802
rect 15052 668 15099 724
rect 15099 668 15126 724
rect 15126 668 15182 724
rect 15182 668 15209 724
rect 15209 668 15265 724
rect 15265 668 15292 724
rect 15292 668 15348 724
rect 15348 668 15374 724
rect 15374 668 15430 724
rect 15430 668 15456 724
rect 15456 668 15512 724
rect 15512 668 15538 724
rect 15538 668 15594 724
rect 15594 668 15620 724
rect 15620 668 15676 724
rect 15676 668 15702 724
rect 15702 668 15758 724
rect 15758 668 15784 724
rect 15784 668 15840 724
rect 15840 668 15866 724
rect 15866 668 15916 724
rect 15052 34 15916 668
rect 15052 -22 15099 34
rect 15099 -22 15126 34
rect 15126 -22 15182 34
rect 15182 -22 15209 34
rect 15209 -22 15265 34
rect 15265 -22 15292 34
rect 15292 -22 15348 34
rect 15348 -22 15374 34
rect 15374 -22 15430 34
rect 15430 -22 15456 34
rect 15456 -22 15512 34
rect 15512 -22 15538 34
rect 15538 -22 15594 34
rect 15594 -22 15620 34
rect 15620 -22 15676 34
rect 15676 -22 15702 34
rect 15702 -22 15758 34
rect 15758 -22 15784 34
rect 15784 -22 15840 34
rect 15840 -22 15866 34
rect 15866 -22 15916 34
rect 15052 -100 15916 -22
rect 15052 -156 15099 -100
rect 15099 -156 15126 -100
rect 15126 -156 15182 -100
rect 15182 -156 15209 -100
rect 15209 -156 15265 -100
rect 15265 -156 15292 -100
rect 15292 -156 15348 -100
rect 15348 -156 15374 -100
rect 15374 -156 15430 -100
rect 15430 -156 15456 -100
rect 15456 -156 15512 -100
rect 15512 -156 15538 -100
rect 15538 -156 15594 -100
rect 15594 -156 15620 -100
rect 15620 -156 15676 -100
rect 15676 -156 15702 -100
rect 15702 -156 15758 -100
rect 15758 -156 15784 -100
rect 15784 -156 15840 -100
rect 15840 -156 15866 -100
rect 15866 -156 15916 -100
rect 15052 -832 15916 -156
rect 15052 -913 15116 -849
rect 15132 -913 15196 -849
rect 15212 -913 15276 -849
rect 15292 -913 15356 -849
rect 15372 -913 15436 -849
rect 15452 -913 15516 -849
rect 15532 -913 15596 -849
rect 15612 -913 15676 -849
rect 15692 -913 15756 -849
rect 15772 -913 15836 -849
rect 15852 -913 15916 -849
rect 15052 -994 15116 -930
rect 15132 -994 15196 -930
rect 15212 -994 15276 -930
rect 15292 -994 15356 -930
rect 15372 -994 15436 -930
rect 15452 -994 15516 -930
rect 15532 -994 15596 -930
rect 15612 -994 15676 -930
rect 15692 -994 15756 -930
rect 15772 -994 15836 -930
rect 15852 -994 15916 -930
rect 15052 -1075 15116 -1011
rect 15132 -1075 15196 -1011
rect 15212 -1075 15276 -1011
rect 15292 -1075 15356 -1011
rect 15372 -1075 15436 -1011
rect 15452 -1075 15516 -1011
rect 15532 -1075 15596 -1011
rect 15612 -1075 15676 -1011
rect 15692 -1075 15756 -1011
rect 15772 -1075 15836 -1011
rect 15852 -1075 15916 -1011
rect 15052 -1156 15116 -1092
rect 15132 -1156 15196 -1092
rect 15212 -1156 15276 -1092
rect 15292 -1156 15356 -1092
rect 15372 -1156 15436 -1092
rect 15452 -1156 15516 -1092
rect 15532 -1156 15596 -1092
rect 15612 -1156 15676 -1092
rect 15692 -1156 15756 -1092
rect 15772 -1156 15836 -1092
rect 15852 -1156 15916 -1092
rect 15052 -1237 15116 -1173
rect 15132 -1237 15196 -1173
rect 15212 -1237 15276 -1173
rect 15292 -1237 15356 -1173
rect 15372 -1237 15436 -1173
rect 15452 -1237 15516 -1173
rect 15532 -1237 15596 -1173
rect 15612 -1237 15676 -1173
rect 15692 -1237 15756 -1173
rect 15772 -1237 15836 -1173
rect 15852 -1237 15916 -1173
rect 15052 -1318 15116 -1254
rect 15132 -1318 15196 -1254
rect 15212 -1318 15276 -1254
rect 15292 -1318 15356 -1254
rect 15372 -1318 15436 -1254
rect 15452 -1318 15516 -1254
rect 15532 -1318 15596 -1254
rect 15612 -1318 15676 -1254
rect 15692 -1318 15756 -1254
rect 15772 -1318 15836 -1254
rect 15852 -1318 15916 -1254
rect 15052 -1399 15116 -1335
rect 15132 -1399 15196 -1335
rect 15212 -1399 15276 -1335
rect 15292 -1399 15356 -1335
rect 15372 -1399 15436 -1335
rect 15452 -1399 15516 -1335
rect 15532 -1399 15596 -1335
rect 15612 -1399 15676 -1335
rect 15692 -1399 15756 -1335
rect 15772 -1399 15836 -1335
rect 15852 -1399 15916 -1335
rect 15052 -1480 15116 -1416
rect 15132 -1480 15196 -1416
rect 15212 -1480 15276 -1416
rect 15292 -1480 15356 -1416
rect 15372 -1480 15436 -1416
rect 15452 -1480 15516 -1416
rect 15532 -1480 15596 -1416
rect 15612 -1480 15676 -1416
rect 15692 -1480 15756 -1416
rect 15772 -1480 15836 -1416
rect 15852 -1480 15916 -1416
rect 15052 -1561 15116 -1497
rect 15132 -1561 15196 -1497
rect 15212 -1561 15276 -1497
rect 15292 -1561 15356 -1497
rect 15372 -1561 15436 -1497
rect 15452 -1561 15516 -1497
rect 15532 -1561 15596 -1497
rect 15612 -1561 15676 -1497
rect 15692 -1561 15756 -1497
rect 15772 -1561 15836 -1497
rect 15852 -1561 15916 -1497
rect 15052 -1642 15116 -1578
rect 15132 -1642 15196 -1578
rect 15212 -1642 15276 -1578
rect 15292 -1642 15356 -1578
rect 15372 -1642 15436 -1578
rect 15452 -1642 15516 -1578
rect 15532 -1642 15596 -1578
rect 15612 -1642 15676 -1578
rect 15692 -1642 15756 -1578
rect 15772 -1642 15836 -1578
rect 15852 -1642 15916 -1578
rect 15052 -1723 15116 -1659
rect 15132 -1723 15196 -1659
rect 15212 -1723 15276 -1659
rect 15292 -1723 15356 -1659
rect 15372 -1723 15436 -1659
rect 15452 -1723 15516 -1659
rect 15532 -1723 15596 -1659
rect 15612 -1723 15676 -1659
rect 15692 -1723 15756 -1659
rect 15772 -1723 15836 -1659
rect 15852 -1723 15916 -1659
rect 15052 -1804 15116 -1740
rect 15132 -1804 15196 -1740
rect 15212 -1804 15276 -1740
rect 15292 -1804 15356 -1740
rect 15372 -1804 15436 -1740
rect 15452 -1804 15516 -1740
rect 15532 -1804 15596 -1740
rect 15612 -1804 15676 -1740
rect 15692 -1804 15756 -1740
rect 15772 -1804 15836 -1740
rect 15852 -1804 15916 -1740
rect 15052 -1885 15116 -1821
rect 15132 -1885 15196 -1821
rect 15212 -1885 15276 -1821
rect 15292 -1885 15356 -1821
rect 15372 -1885 15436 -1821
rect 15452 -1885 15516 -1821
rect 15532 -1885 15596 -1821
rect 15612 -1885 15676 -1821
rect 15692 -1885 15756 -1821
rect 15772 -1885 15836 -1821
rect 15852 -1885 15916 -1821
rect 15052 -1966 15116 -1902
rect 15132 -1966 15196 -1902
rect 15212 -1966 15276 -1902
rect 15292 -1966 15356 -1902
rect 15372 -1966 15436 -1902
rect 15452 -1966 15516 -1902
rect 15532 -1966 15596 -1902
rect 15612 -1966 15676 -1902
rect 15692 -1966 15756 -1902
rect 15772 -1966 15836 -1902
rect 15852 -1966 15916 -1902
rect 15052 -2047 15116 -1983
rect 15132 -2047 15196 -1983
rect 15212 -2047 15276 -1983
rect 15292 -2047 15356 -1983
rect 15372 -2047 15436 -1983
rect 15452 -2047 15516 -1983
rect 15532 -2047 15596 -1983
rect 15612 -2047 15676 -1983
rect 15692 -2047 15756 -1983
rect 15772 -2047 15836 -1983
rect 15852 -2047 15916 -1983
rect 15052 -2128 15116 -2064
rect 15132 -2128 15196 -2064
rect 15212 -2128 15276 -2064
rect 15292 -2128 15356 -2064
rect 15372 -2128 15436 -2064
rect 15452 -2128 15516 -2064
rect 15532 -2128 15596 -2064
rect 15612 -2128 15676 -2064
rect 15692 -2128 15756 -2064
rect 15772 -2128 15836 -2064
rect 15852 -2128 15916 -2064
rect 15052 -2209 15116 -2145
rect 15132 -2209 15196 -2145
rect 15212 -2209 15276 -2145
rect 15292 -2209 15356 -2145
rect 15372 -2209 15436 -2145
rect 15452 -2209 15516 -2145
rect 15532 -2209 15596 -2145
rect 15612 -2209 15676 -2145
rect 15692 -2209 15756 -2145
rect 15772 -2209 15836 -2145
rect 15852 -2209 15916 -2145
rect 15052 -2290 15116 -2226
rect 15132 -2290 15196 -2226
rect 15212 -2290 15276 -2226
rect 15292 -2290 15356 -2226
rect 15372 -2290 15436 -2226
rect 15452 -2290 15516 -2226
rect 15532 -2290 15596 -2226
rect 15612 -2290 15676 -2226
rect 15692 -2290 15756 -2226
rect 15772 -2290 15836 -2226
rect 15852 -2290 15916 -2226
rect 15052 -2371 15116 -2307
rect 15132 -2371 15196 -2307
rect 15212 -2371 15276 -2307
rect 15292 -2371 15356 -2307
rect 15372 -2371 15436 -2307
rect 15452 -2371 15516 -2307
rect 15532 -2371 15596 -2307
rect 15612 -2371 15676 -2307
rect 15692 -2371 15756 -2307
rect 15772 -2371 15836 -2307
rect 15852 -2371 15916 -2307
rect 15052 -2452 15116 -2388
rect 15132 -2452 15196 -2388
rect 15212 -2452 15276 -2388
rect 15292 -2452 15356 -2388
rect 15372 -2452 15436 -2388
rect 15452 -2452 15516 -2388
rect 15532 -2452 15596 -2388
rect 15612 -2452 15676 -2388
rect 15692 -2452 15756 -2388
rect 15772 -2452 15836 -2388
rect 15852 -2452 15916 -2388
rect 15052 -2533 15116 -2469
rect 15132 -2533 15196 -2469
rect 15212 -2533 15276 -2469
rect 15292 -2533 15356 -2469
rect 15372 -2533 15436 -2469
rect 15452 -2533 15516 -2469
rect 15532 -2533 15596 -2469
rect 15612 -2533 15676 -2469
rect 15692 -2533 15756 -2469
rect 15772 -2533 15836 -2469
rect 15852 -2533 15916 -2469
rect 15052 -2614 15116 -2550
rect 15132 -2614 15196 -2550
rect 15212 -2614 15276 -2550
rect 15292 -2614 15356 -2550
rect 15372 -2614 15436 -2550
rect 15452 -2614 15516 -2550
rect 15532 -2614 15596 -2550
rect 15612 -2614 15676 -2550
rect 15692 -2614 15756 -2550
rect 15772 -2614 15836 -2550
rect 15852 -2614 15916 -2550
rect 9540 -3000 9604 -2936
rect 9620 -3000 9684 -2936
rect 9700 -3000 9764 -2936
rect 9540 -3081 9604 -3017
rect 9620 -3081 9684 -3017
rect 9700 -3081 9764 -3017
rect 9540 -3162 9604 -3098
rect 9620 -3162 9684 -3098
rect 9700 -3162 9764 -3098
rect 9540 -3243 9604 -3179
rect 9620 -3243 9684 -3179
rect 9700 -3243 9764 -3179
rect 9540 -3324 9604 -3260
rect 9620 -3324 9684 -3260
rect 9700 -3324 9764 -3260
rect 9540 -3405 9604 -3341
rect 9620 -3405 9684 -3341
rect 9700 -3405 9764 -3341
rect 9540 -3487 9604 -3423
rect 9620 -3487 9684 -3423
rect 9700 -3487 9764 -3423
rect 9540 -3569 9604 -3505
rect 9620 -3569 9684 -3505
rect 9700 -3569 9764 -3505
rect 9540 -3651 9604 -3587
rect 9620 -3651 9684 -3587
rect 9700 -3651 9764 -3587
rect 9540 -3733 9604 -3669
rect 9620 -3733 9684 -3669
rect 9700 -3733 9764 -3669
rect 6492 -3806 6556 -3742
rect 6594 -3806 6658 -3742
rect 6696 -3806 6760 -3742
rect 6798 -3806 6862 -3742
rect 16544 -3320 16768 -2936
rect 16891 858 17755 2352
rect 16891 802 16940 858
rect 16940 802 16966 858
rect 16966 802 17022 858
rect 17022 802 17048 858
rect 17048 802 17104 858
rect 17104 802 17130 858
rect 17130 802 17186 858
rect 17186 802 17212 858
rect 17212 802 17268 858
rect 17268 802 17294 858
rect 17294 802 17350 858
rect 17350 802 17376 858
rect 17376 802 17432 858
rect 17432 802 17458 858
rect 17458 802 17514 858
rect 17514 802 17541 858
rect 17541 802 17597 858
rect 17597 802 17624 858
rect 17624 802 17680 858
rect 17680 802 17707 858
rect 17707 802 17755 858
rect 16891 724 17755 802
rect 16891 668 16940 724
rect 16940 668 16966 724
rect 16966 668 17022 724
rect 17022 668 17048 724
rect 17048 668 17104 724
rect 17104 668 17130 724
rect 17130 668 17186 724
rect 17186 668 17212 724
rect 17212 668 17268 724
rect 17268 668 17294 724
rect 17294 668 17350 724
rect 17350 668 17376 724
rect 17376 668 17432 724
rect 17432 668 17458 724
rect 17458 668 17514 724
rect 17514 668 17541 724
rect 17541 668 17597 724
rect 17597 668 17624 724
rect 17624 668 17680 724
rect 17680 668 17707 724
rect 17707 668 17755 724
rect 16891 34 17755 668
rect 16891 -22 16940 34
rect 16940 -22 16967 34
rect 16967 -22 17023 34
rect 17023 -22 17050 34
rect 17050 -22 17106 34
rect 17106 -22 17133 34
rect 17133 -22 17189 34
rect 17189 -22 17215 34
rect 17215 -22 17271 34
rect 17271 -22 17297 34
rect 17297 -22 17353 34
rect 17353 -22 17379 34
rect 17379 -22 17435 34
rect 17435 -22 17461 34
rect 17461 -22 17517 34
rect 17517 -22 17543 34
rect 17543 -22 17599 34
rect 17599 -22 17625 34
rect 17625 -22 17681 34
rect 17681 -22 17707 34
rect 17707 -22 17755 34
rect 16891 -100 17755 -22
rect 16891 -156 16940 -100
rect 16940 -156 16967 -100
rect 16967 -156 17023 -100
rect 17023 -156 17050 -100
rect 17050 -156 17106 -100
rect 17106 -156 17133 -100
rect 17133 -156 17189 -100
rect 17189 -156 17215 -100
rect 17215 -156 17271 -100
rect 17271 -156 17297 -100
rect 17297 -156 17353 -100
rect 17353 -156 17379 -100
rect 17379 -156 17435 -100
rect 17435 -156 17461 -100
rect 17461 -156 17517 -100
rect 17517 -156 17543 -100
rect 17543 -156 17599 -100
rect 17599 -156 17625 -100
rect 17625 -156 17681 -100
rect 17681 -156 17707 -100
rect 17707 -156 17755 -100
rect 16891 -832 17755 -156
rect 16891 -913 16955 -849
rect 16971 -913 17035 -849
rect 17051 -913 17115 -849
rect 17131 -913 17195 -849
rect 17211 -913 17275 -849
rect 17291 -913 17355 -849
rect 17371 -913 17435 -849
rect 17451 -913 17515 -849
rect 17531 -913 17595 -849
rect 17611 -913 17675 -849
rect 17691 -913 17755 -849
rect 16891 -994 16955 -930
rect 16971 -994 17035 -930
rect 17051 -994 17115 -930
rect 17131 -994 17195 -930
rect 17211 -994 17275 -930
rect 17291 -994 17355 -930
rect 17371 -994 17435 -930
rect 17451 -994 17515 -930
rect 17531 -994 17595 -930
rect 17611 -994 17675 -930
rect 17691 -994 17755 -930
rect 16891 -1075 16955 -1011
rect 16971 -1075 17035 -1011
rect 17051 -1075 17115 -1011
rect 17131 -1075 17195 -1011
rect 17211 -1075 17275 -1011
rect 17291 -1075 17355 -1011
rect 17371 -1075 17435 -1011
rect 17451 -1075 17515 -1011
rect 17531 -1075 17595 -1011
rect 17611 -1075 17675 -1011
rect 17691 -1075 17755 -1011
rect 16891 -1156 16955 -1092
rect 16971 -1156 17035 -1092
rect 17051 -1156 17115 -1092
rect 17131 -1156 17195 -1092
rect 17211 -1156 17275 -1092
rect 17291 -1156 17355 -1092
rect 17371 -1156 17435 -1092
rect 17451 -1156 17515 -1092
rect 17531 -1156 17595 -1092
rect 17611 -1156 17675 -1092
rect 17691 -1156 17755 -1092
rect 16891 -1237 16955 -1173
rect 16971 -1237 17035 -1173
rect 17051 -1237 17115 -1173
rect 17131 -1237 17195 -1173
rect 17211 -1237 17275 -1173
rect 17291 -1237 17355 -1173
rect 17371 -1237 17435 -1173
rect 17451 -1237 17515 -1173
rect 17531 -1237 17595 -1173
rect 17611 -1237 17675 -1173
rect 17691 -1237 17755 -1173
rect 16891 -1318 16955 -1254
rect 16971 -1318 17035 -1254
rect 17051 -1318 17115 -1254
rect 17131 -1318 17195 -1254
rect 17211 -1318 17275 -1254
rect 17291 -1318 17355 -1254
rect 17371 -1318 17435 -1254
rect 17451 -1318 17515 -1254
rect 17531 -1318 17595 -1254
rect 17611 -1318 17675 -1254
rect 17691 -1318 17755 -1254
rect 16891 -1399 16955 -1335
rect 16971 -1399 17035 -1335
rect 17051 -1399 17115 -1335
rect 17131 -1399 17195 -1335
rect 17211 -1399 17275 -1335
rect 17291 -1399 17355 -1335
rect 17371 -1399 17435 -1335
rect 17451 -1399 17515 -1335
rect 17531 -1399 17595 -1335
rect 17611 -1399 17675 -1335
rect 17691 -1399 17755 -1335
rect 16891 -1480 16955 -1416
rect 16971 -1480 17035 -1416
rect 17051 -1480 17115 -1416
rect 17131 -1480 17195 -1416
rect 17211 -1480 17275 -1416
rect 17291 -1480 17355 -1416
rect 17371 -1480 17435 -1416
rect 17451 -1480 17515 -1416
rect 17531 -1480 17595 -1416
rect 17611 -1480 17675 -1416
rect 17691 -1480 17755 -1416
rect 16891 -1561 16955 -1497
rect 16971 -1561 17035 -1497
rect 17051 -1561 17115 -1497
rect 17131 -1561 17195 -1497
rect 17211 -1561 17275 -1497
rect 17291 -1561 17355 -1497
rect 17371 -1561 17435 -1497
rect 17451 -1561 17515 -1497
rect 17531 -1561 17595 -1497
rect 17611 -1561 17675 -1497
rect 17691 -1561 17755 -1497
rect 16891 -1642 16955 -1578
rect 16971 -1642 17035 -1578
rect 17051 -1642 17115 -1578
rect 17131 -1642 17195 -1578
rect 17211 -1642 17275 -1578
rect 17291 -1642 17355 -1578
rect 17371 -1642 17435 -1578
rect 17451 -1642 17515 -1578
rect 17531 -1642 17595 -1578
rect 17611 -1642 17675 -1578
rect 17691 -1642 17755 -1578
rect 16891 -1723 16955 -1659
rect 16971 -1723 17035 -1659
rect 17051 -1723 17115 -1659
rect 17131 -1723 17195 -1659
rect 17211 -1723 17275 -1659
rect 17291 -1723 17355 -1659
rect 17371 -1723 17435 -1659
rect 17451 -1723 17515 -1659
rect 17531 -1723 17595 -1659
rect 17611 -1723 17675 -1659
rect 17691 -1723 17755 -1659
rect 16891 -1804 16955 -1740
rect 16971 -1804 17035 -1740
rect 17051 -1804 17115 -1740
rect 17131 -1804 17195 -1740
rect 17211 -1804 17275 -1740
rect 17291 -1804 17355 -1740
rect 17371 -1804 17435 -1740
rect 17451 -1804 17515 -1740
rect 17531 -1804 17595 -1740
rect 17611 -1804 17675 -1740
rect 17691 -1804 17755 -1740
rect 16891 -1885 16955 -1821
rect 16971 -1885 17035 -1821
rect 17051 -1885 17115 -1821
rect 17131 -1885 17195 -1821
rect 17211 -1885 17275 -1821
rect 17291 -1885 17355 -1821
rect 17371 -1885 17435 -1821
rect 17451 -1885 17515 -1821
rect 17531 -1885 17595 -1821
rect 17611 -1885 17675 -1821
rect 17691 -1885 17755 -1821
rect 16891 -1966 16955 -1902
rect 16971 -1966 17035 -1902
rect 17051 -1966 17115 -1902
rect 17131 -1966 17195 -1902
rect 17211 -1966 17275 -1902
rect 17291 -1966 17355 -1902
rect 17371 -1966 17435 -1902
rect 17451 -1966 17515 -1902
rect 17531 -1966 17595 -1902
rect 17611 -1966 17675 -1902
rect 17691 -1966 17755 -1902
rect 16891 -2047 16955 -1983
rect 16971 -2047 17035 -1983
rect 17051 -2047 17115 -1983
rect 17131 -2047 17195 -1983
rect 17211 -2047 17275 -1983
rect 17291 -2047 17355 -1983
rect 17371 -2047 17435 -1983
rect 17451 -2047 17515 -1983
rect 17531 -2047 17595 -1983
rect 17611 -2047 17675 -1983
rect 17691 -2047 17755 -1983
rect 16891 -2128 16955 -2064
rect 16971 -2128 17035 -2064
rect 17051 -2128 17115 -2064
rect 17131 -2128 17195 -2064
rect 17211 -2128 17275 -2064
rect 17291 -2128 17355 -2064
rect 17371 -2128 17435 -2064
rect 17451 -2128 17515 -2064
rect 17531 -2128 17595 -2064
rect 17611 -2128 17675 -2064
rect 17691 -2128 17755 -2064
rect 16891 -2209 16955 -2145
rect 16971 -2209 17035 -2145
rect 17051 -2209 17115 -2145
rect 17131 -2209 17195 -2145
rect 17211 -2209 17275 -2145
rect 17291 -2209 17355 -2145
rect 17371 -2209 17435 -2145
rect 17451 -2209 17515 -2145
rect 17531 -2209 17595 -2145
rect 17611 -2209 17675 -2145
rect 17691 -2209 17755 -2145
rect 16891 -2290 16955 -2226
rect 16971 -2290 17035 -2226
rect 17051 -2290 17115 -2226
rect 17131 -2290 17195 -2226
rect 17211 -2290 17275 -2226
rect 17291 -2290 17355 -2226
rect 17371 -2290 17435 -2226
rect 17451 -2290 17515 -2226
rect 17531 -2290 17595 -2226
rect 17611 -2290 17675 -2226
rect 17691 -2290 17755 -2226
rect 16891 -2371 16955 -2307
rect 16971 -2371 17035 -2307
rect 17051 -2371 17115 -2307
rect 17131 -2371 17195 -2307
rect 17211 -2371 17275 -2307
rect 17291 -2371 17355 -2307
rect 17371 -2371 17435 -2307
rect 17451 -2371 17515 -2307
rect 17531 -2371 17595 -2307
rect 17611 -2371 17675 -2307
rect 17691 -2371 17755 -2307
rect 16891 -2452 16955 -2388
rect 16971 -2452 17035 -2388
rect 17051 -2452 17115 -2388
rect 17131 -2452 17195 -2388
rect 17211 -2452 17275 -2388
rect 17291 -2452 17355 -2388
rect 17371 -2452 17435 -2388
rect 17451 -2452 17515 -2388
rect 17531 -2452 17595 -2388
rect 17611 -2452 17675 -2388
rect 17691 -2452 17755 -2388
rect 16891 -2533 16955 -2469
rect 16971 -2533 17035 -2469
rect 17051 -2533 17115 -2469
rect 17131 -2533 17195 -2469
rect 17211 -2533 17275 -2469
rect 17291 -2533 17355 -2469
rect 17371 -2533 17435 -2469
rect 17451 -2533 17515 -2469
rect 17531 -2533 17595 -2469
rect 17611 -2533 17675 -2469
rect 17691 -2533 17755 -2469
rect 16891 -2614 16955 -2550
rect 16971 -2614 17035 -2550
rect 17051 -2614 17115 -2550
rect 17131 -2614 17195 -2550
rect 17211 -2614 17275 -2550
rect 17291 -2614 17355 -2550
rect 17371 -2614 17435 -2550
rect 17451 -2614 17515 -2550
rect 17531 -2614 17595 -2550
rect 17611 -2614 17675 -2550
rect 17691 -2614 17755 -2550
rect 16544 -3401 16608 -3337
rect 16624 -3401 16688 -3337
rect 16704 -3401 16768 -3337
rect 16544 -3482 16608 -3418
rect 16624 -3482 16688 -3418
rect 16704 -3482 16768 -3418
rect 16544 -3563 16608 -3499
rect 16624 -3563 16688 -3499
rect 16704 -3563 16768 -3499
rect 16544 -3644 16608 -3580
rect 16624 -3644 16688 -3580
rect 16704 -3644 16768 -3580
rect 16544 -3725 16608 -3661
rect 16624 -3725 16688 -3661
rect 16704 -3725 16768 -3661
rect 16544 -3806 16608 -3742
rect 16624 -3806 16688 -3742
rect 16704 -3806 16768 -3742
<< metal4 >>
tri 13098 5258 13469 5629 se
rect 13469 5258 14233 5629
tri 14233 5258 14604 5629 sw
tri 13066 5226 13098 5258 se
rect 13098 5226 18805 5258
tri 12703 4863 13066 5226 se
rect 13066 4863 14014 5226
rect 1033 4856 14014 4863
rect 1033 4792 1047 4856
rect 1111 4792 1135 4856
rect 1199 4792 1223 4856
rect 1287 4792 1311 4856
rect 1375 4792 1399 4856
rect 1463 4792 1487 4856
rect 1551 4792 1575 4856
rect 1639 4792 1662 4856
rect 1726 4792 1749 4856
rect 1813 4792 1836 4856
rect 1900 4792 4713 4856
rect 4777 4792 4794 4856
rect 4858 4792 4875 4856
rect 4939 4792 4956 4856
rect 5020 4792 5037 4856
rect 5101 4792 5118 4856
rect 5182 4792 5198 4856
rect 5262 4792 5278 4856
rect 5342 4792 5358 4856
rect 5422 4792 5438 4856
rect 5502 4792 5518 4856
rect 5582 4792 5598 4856
rect 5662 4792 5678 4856
rect 5742 4792 5758 4856
rect 5822 4792 7531 4856
rect 7595 4792 7617 4856
rect 7681 4792 7703 4856
rect 7767 4792 7789 4856
rect 7853 4792 7875 4856
rect 7939 4792 7961 4856
rect 8025 4792 8047 4856
rect 8111 4792 8133 4856
rect 8197 4792 8219 4856
rect 8283 4792 8305 4856
rect 8369 4792 8391 4856
rect 8455 4792 8477 4856
rect 8541 4792 8563 4856
rect 8627 4792 8648 4856
rect 8712 4792 11453 4856
rect 11517 4792 11541 4856
rect 11605 4792 11629 4856
rect 11693 4792 11717 4856
rect 11781 4792 11805 4856
rect 11869 4792 11893 4856
rect 11957 4792 11981 4856
rect 12045 4792 12068 4856
rect 12132 4792 12155 4856
rect 12219 4792 12242 4856
rect 12306 4792 14014 4856
rect 1033 4764 14014 4792
rect 1033 4700 1047 4764
rect 1111 4700 1135 4764
rect 1199 4700 1223 4764
rect 1287 4700 1311 4764
rect 1375 4700 1399 4764
rect 1463 4700 1487 4764
rect 1551 4700 1575 4764
rect 1639 4700 1662 4764
rect 1726 4700 1749 4764
rect 1813 4700 1836 4764
rect 1900 4700 4713 4764
rect 4777 4700 4794 4764
rect 4858 4700 4875 4764
rect 4939 4700 4956 4764
rect 5020 4700 5037 4764
rect 5101 4700 5118 4764
rect 5182 4700 5198 4764
rect 5262 4700 5278 4764
rect 5342 4700 5358 4764
rect 5422 4700 5438 4764
rect 5502 4700 5518 4764
rect 5582 4700 5598 4764
rect 5662 4700 5678 4764
rect 5742 4700 5758 4764
rect 5822 4700 7531 4764
rect 7595 4700 7617 4764
rect 7681 4700 7703 4764
rect 7767 4700 7789 4764
rect 7853 4700 7875 4764
rect 7939 4700 7961 4764
rect 8025 4700 8047 4764
rect 8111 4700 8133 4764
rect 8197 4700 8219 4764
rect 8283 4700 8305 4764
rect 8369 4700 8391 4764
rect 8455 4700 8477 4764
rect 8541 4700 8563 4764
rect 8627 4700 8648 4764
rect 8712 4700 11453 4764
rect 11517 4700 11541 4764
rect 11605 4700 11629 4764
rect 11693 4700 11717 4764
rect 11781 4700 11805 4764
rect 11869 4700 11893 4764
rect 11957 4700 11981 4764
rect 12045 4700 12068 4764
rect 12132 4700 12155 4764
rect 12219 4700 12242 4764
rect 12306 4700 14014 4764
rect 1033 4672 14014 4700
rect 1033 4608 1047 4672
rect 1111 4608 1135 4672
rect 1199 4608 1223 4672
rect 1287 4608 1311 4672
rect 1375 4608 1399 4672
rect 1463 4608 1487 4672
rect 1551 4608 1575 4672
rect 1639 4608 1662 4672
rect 1726 4608 1749 4672
rect 1813 4608 1836 4672
rect 1900 4608 4713 4672
rect 4777 4608 4794 4672
rect 4858 4608 4875 4672
rect 4939 4608 4956 4672
rect 5020 4608 5037 4672
rect 5101 4608 5118 4672
rect 5182 4608 5198 4672
rect 5262 4608 5278 4672
rect 5342 4608 5358 4672
rect 5422 4608 5438 4672
rect 5502 4608 5518 4672
rect 5582 4608 5598 4672
rect 5662 4608 5678 4672
rect 5742 4608 5758 4672
rect 5822 4608 7531 4672
rect 7595 4608 7617 4672
rect 7681 4608 7703 4672
rect 7767 4608 7789 4672
rect 7853 4608 7875 4672
rect 7939 4608 7961 4672
rect 8025 4608 8047 4672
rect 8111 4608 8133 4672
rect 8197 4608 8219 4672
rect 8283 4608 8305 4672
rect 8369 4608 8391 4672
rect 8455 4608 8477 4672
rect 8541 4608 8563 4672
rect 8627 4608 8648 4672
rect 8712 4608 11453 4672
rect 11517 4608 11541 4672
rect 11605 4608 11629 4672
rect 11693 4608 11717 4672
rect 11781 4608 11805 4672
rect 11869 4608 11893 4672
rect 11957 4608 11981 4672
rect 12045 4608 12068 4672
rect 12132 4608 12155 4672
rect 12219 4608 12242 4672
rect 12306 4608 14014 4672
rect 1033 4580 14014 4608
rect 1033 4516 1047 4580
rect 1111 4516 1135 4580
rect 1199 4516 1223 4580
rect 1287 4516 1311 4580
rect 1375 4516 1399 4580
rect 1463 4516 1487 4580
rect 1551 4516 1575 4580
rect 1639 4516 1662 4580
rect 1726 4516 1749 4580
rect 1813 4516 1836 4580
rect 1900 4516 4713 4580
rect 4777 4516 4794 4580
rect 4858 4516 4875 4580
rect 4939 4516 4956 4580
rect 5020 4516 5037 4580
rect 5101 4516 5118 4580
rect 5182 4516 5198 4580
rect 5262 4516 5278 4580
rect 5342 4516 5358 4580
rect 5422 4516 5438 4580
rect 5502 4516 5518 4580
rect 5582 4516 5598 4580
rect 5662 4516 5678 4580
rect 5742 4516 5758 4580
rect 5822 4516 7531 4580
rect 7595 4516 7617 4580
rect 7681 4516 7703 4580
rect 7767 4516 7789 4580
rect 7853 4516 7875 4580
rect 7939 4516 7961 4580
rect 8025 4516 8047 4580
rect 8111 4516 8133 4580
rect 8197 4516 8219 4580
rect 8283 4516 8305 4580
rect 8369 4516 8391 4580
rect 8455 4516 8477 4580
rect 8541 4516 8563 4580
rect 8627 4516 8648 4580
rect 8712 4516 11453 4580
rect 11517 4516 11541 4580
rect 11605 4516 11629 4580
rect 11693 4516 11717 4580
rect 11781 4516 11805 4580
rect 11869 4516 11893 4580
rect 11957 4516 11981 4580
rect 12045 4516 12068 4580
rect 12132 4516 12155 4580
rect 12219 4516 12242 4580
rect 12306 4516 14014 4580
rect 1033 4488 14014 4516
rect 1033 4424 1047 4488
rect 1111 4424 1135 4488
rect 1199 4424 1223 4488
rect 1287 4424 1311 4488
rect 1375 4424 1399 4488
rect 1463 4424 1487 4488
rect 1551 4424 1575 4488
rect 1639 4424 1662 4488
rect 1726 4424 1749 4488
rect 1813 4424 1836 4488
rect 1900 4424 4713 4488
rect 4777 4424 4794 4488
rect 4858 4424 4875 4488
rect 4939 4424 4956 4488
rect 5020 4424 5037 4488
rect 5101 4424 5118 4488
rect 5182 4424 5198 4488
rect 5262 4424 5278 4488
rect 5342 4424 5358 4488
rect 5422 4424 5438 4488
rect 5502 4424 5518 4488
rect 5582 4424 5598 4488
rect 5662 4424 5678 4488
rect 5742 4424 5758 4488
rect 5822 4424 7531 4488
rect 7595 4424 7617 4488
rect 7681 4424 7703 4488
rect 7767 4424 7789 4488
rect 7853 4424 7875 4488
rect 7939 4424 7961 4488
rect 8025 4424 8047 4488
rect 8111 4424 8133 4488
rect 8197 4424 8219 4488
rect 8283 4424 8305 4488
rect 8369 4424 8391 4488
rect 8455 4424 8477 4488
rect 8541 4424 8563 4488
rect 8627 4424 8648 4488
rect 8712 4424 11453 4488
rect 11517 4424 11541 4488
rect 11605 4424 11629 4488
rect 11693 4424 11717 4488
rect 11781 4424 11805 4488
rect 11869 4424 11893 4488
rect 11957 4424 11981 4488
rect 12045 4424 12068 4488
rect 12132 4424 12155 4488
rect 12219 4424 12242 4488
rect 12306 4424 14014 4488
rect 1033 4396 14014 4424
rect 1033 4332 1047 4396
rect 1111 4332 1135 4396
rect 1199 4332 1223 4396
rect 1287 4332 1311 4396
rect 1375 4332 1399 4396
rect 1463 4332 1487 4396
rect 1551 4332 1575 4396
rect 1639 4332 1662 4396
rect 1726 4332 1749 4396
rect 1813 4332 1836 4396
rect 1900 4332 4713 4396
rect 4777 4332 4794 4396
rect 4858 4332 4875 4396
rect 4939 4332 4956 4396
rect 5020 4332 5037 4396
rect 5101 4332 5118 4396
rect 5182 4332 5198 4396
rect 5262 4332 5278 4396
rect 5342 4332 5358 4396
rect 5422 4332 5438 4396
rect 5502 4332 5518 4396
rect 5582 4332 5598 4396
rect 5662 4332 5678 4396
rect 5742 4332 5758 4396
rect 5822 4332 7531 4396
rect 7595 4332 7617 4396
rect 7681 4332 7703 4396
rect 7767 4332 7789 4396
rect 7853 4332 7875 4396
rect 7939 4332 7961 4396
rect 8025 4332 8047 4396
rect 8111 4332 8133 4396
rect 8197 4332 8219 4396
rect 8283 4332 8305 4396
rect 8369 4332 8391 4396
rect 8455 4332 8477 4396
rect 8541 4332 8563 4396
rect 8627 4332 8648 4396
rect 8712 4332 11453 4396
rect 11517 4332 11541 4396
rect 11605 4332 11629 4396
rect 11693 4332 11717 4396
rect 11781 4332 11805 4396
rect 11869 4332 11893 4396
rect 11957 4332 11981 4396
rect 12045 4332 12068 4396
rect 12132 4332 12155 4396
rect 12219 4332 12242 4396
rect 12306 4362 14014 4396
rect 14878 4362 17934 5226
rect 18798 4362 18805 5226
rect 12306 4332 18805 4362
rect 1033 4323 18805 4332
rect 2080 2352 17760 2353
rect 2080 -832 3924 2352
rect 4788 -832 8568 2352
rect 9432 -832 10407 2352
rect 11271 -832 15052 2352
rect 15916 -832 16891 2352
rect 17755 -832 17760 2352
rect 2080 -849 17760 -832
rect 2080 -913 3924 -849
rect 3988 -913 4004 -849
rect 4068 -913 4084 -849
rect 4148 -913 4164 -849
rect 4228 -913 4244 -849
rect 4308 -913 4324 -849
rect 4388 -913 4404 -849
rect 4468 -913 4484 -849
rect 4548 -913 4564 -849
rect 4628 -913 4644 -849
rect 4708 -913 4724 -849
rect 4788 -913 8568 -849
rect 8632 -913 8648 -849
rect 8712 -913 8728 -849
rect 8792 -913 8808 -849
rect 8872 -913 8888 -849
rect 8952 -913 8968 -849
rect 9032 -913 9048 -849
rect 9112 -913 9128 -849
rect 9192 -913 9208 -849
rect 9272 -913 9288 -849
rect 9352 -913 9368 -849
rect 9432 -913 10407 -849
rect 10471 -913 10487 -849
rect 10551 -913 10567 -849
rect 10631 -913 10647 -849
rect 10711 -913 10727 -849
rect 10791 -913 10807 -849
rect 10871 -913 10887 -849
rect 10951 -913 10967 -849
rect 11031 -913 11047 -849
rect 11111 -913 11127 -849
rect 11191 -913 11207 -849
rect 11271 -913 15052 -849
rect 15116 -913 15132 -849
rect 15196 -913 15212 -849
rect 15276 -913 15292 -849
rect 15356 -913 15372 -849
rect 15436 -913 15452 -849
rect 15516 -913 15532 -849
rect 15596 -913 15612 -849
rect 15676 -913 15692 -849
rect 15756 -913 15772 -849
rect 15836 -913 15852 -849
rect 15916 -913 16891 -849
rect 16955 -913 16971 -849
rect 17035 -913 17051 -849
rect 17115 -913 17131 -849
rect 17195 -913 17211 -849
rect 17275 -913 17291 -849
rect 17355 -913 17371 -849
rect 17435 -913 17451 -849
rect 17515 -913 17531 -849
rect 17595 -913 17611 -849
rect 17675 -913 17691 -849
rect 17755 -913 17760 -849
rect 2080 -930 17760 -913
rect 2080 -994 3924 -930
rect 3988 -994 4004 -930
rect 4068 -994 4084 -930
rect 4148 -994 4164 -930
rect 4228 -994 4244 -930
rect 4308 -994 4324 -930
rect 4388 -994 4404 -930
rect 4468 -994 4484 -930
rect 4548 -994 4564 -930
rect 4628 -994 4644 -930
rect 4708 -994 4724 -930
rect 4788 -994 8568 -930
rect 8632 -994 8648 -930
rect 8712 -994 8728 -930
rect 8792 -994 8808 -930
rect 8872 -994 8888 -930
rect 8952 -994 8968 -930
rect 9032 -994 9048 -930
rect 9112 -994 9128 -930
rect 9192 -994 9208 -930
rect 9272 -994 9288 -930
rect 9352 -994 9368 -930
rect 9432 -994 10407 -930
rect 10471 -994 10487 -930
rect 10551 -994 10567 -930
rect 10631 -994 10647 -930
rect 10711 -994 10727 -930
rect 10791 -994 10807 -930
rect 10871 -994 10887 -930
rect 10951 -994 10967 -930
rect 11031 -994 11047 -930
rect 11111 -994 11127 -930
rect 11191 -994 11207 -930
rect 11271 -994 15052 -930
rect 15116 -994 15132 -930
rect 15196 -994 15212 -930
rect 15276 -994 15292 -930
rect 15356 -994 15372 -930
rect 15436 -994 15452 -930
rect 15516 -994 15532 -930
rect 15596 -994 15612 -930
rect 15676 -994 15692 -930
rect 15756 -994 15772 -930
rect 15836 -994 15852 -930
rect 15916 -994 16891 -930
rect 16955 -994 16971 -930
rect 17035 -994 17051 -930
rect 17115 -994 17131 -930
rect 17195 -994 17211 -930
rect 17275 -994 17291 -930
rect 17355 -994 17371 -930
rect 17435 -994 17451 -930
rect 17515 -994 17531 -930
rect 17595 -994 17611 -930
rect 17675 -994 17691 -930
rect 17755 -994 17760 -930
rect 2080 -1011 17760 -994
rect 2080 -1075 3924 -1011
rect 3988 -1075 4004 -1011
rect 4068 -1075 4084 -1011
rect 4148 -1075 4164 -1011
rect 4228 -1075 4244 -1011
rect 4308 -1075 4324 -1011
rect 4388 -1075 4404 -1011
rect 4468 -1075 4484 -1011
rect 4548 -1075 4564 -1011
rect 4628 -1075 4644 -1011
rect 4708 -1075 4724 -1011
rect 4788 -1075 8568 -1011
rect 8632 -1075 8648 -1011
rect 8712 -1075 8728 -1011
rect 8792 -1075 8808 -1011
rect 8872 -1075 8888 -1011
rect 8952 -1075 8968 -1011
rect 9032 -1075 9048 -1011
rect 9112 -1075 9128 -1011
rect 9192 -1075 9208 -1011
rect 9272 -1075 9288 -1011
rect 9352 -1075 9368 -1011
rect 9432 -1075 10407 -1011
rect 10471 -1075 10487 -1011
rect 10551 -1075 10567 -1011
rect 10631 -1075 10647 -1011
rect 10711 -1075 10727 -1011
rect 10791 -1075 10807 -1011
rect 10871 -1075 10887 -1011
rect 10951 -1075 10967 -1011
rect 11031 -1075 11047 -1011
rect 11111 -1075 11127 -1011
rect 11191 -1075 11207 -1011
rect 11271 -1075 15052 -1011
rect 15116 -1075 15132 -1011
rect 15196 -1075 15212 -1011
rect 15276 -1075 15292 -1011
rect 15356 -1075 15372 -1011
rect 15436 -1075 15452 -1011
rect 15516 -1075 15532 -1011
rect 15596 -1075 15612 -1011
rect 15676 -1075 15692 -1011
rect 15756 -1075 15772 -1011
rect 15836 -1075 15852 -1011
rect 15916 -1075 16891 -1011
rect 16955 -1075 16971 -1011
rect 17035 -1075 17051 -1011
rect 17115 -1075 17131 -1011
rect 17195 -1075 17211 -1011
rect 17275 -1075 17291 -1011
rect 17355 -1075 17371 -1011
rect 17435 -1075 17451 -1011
rect 17515 -1075 17531 -1011
rect 17595 -1075 17611 -1011
rect 17675 -1075 17691 -1011
rect 17755 -1075 17760 -1011
rect 2080 -1092 17760 -1075
rect 2080 -1156 3924 -1092
rect 3988 -1156 4004 -1092
rect 4068 -1156 4084 -1092
rect 4148 -1156 4164 -1092
rect 4228 -1156 4244 -1092
rect 4308 -1156 4324 -1092
rect 4388 -1156 4404 -1092
rect 4468 -1156 4484 -1092
rect 4548 -1156 4564 -1092
rect 4628 -1156 4644 -1092
rect 4708 -1156 4724 -1092
rect 4788 -1156 8568 -1092
rect 8632 -1156 8648 -1092
rect 8712 -1156 8728 -1092
rect 8792 -1156 8808 -1092
rect 8872 -1156 8888 -1092
rect 8952 -1156 8968 -1092
rect 9032 -1156 9048 -1092
rect 9112 -1156 9128 -1092
rect 9192 -1156 9208 -1092
rect 9272 -1156 9288 -1092
rect 9352 -1156 9368 -1092
rect 9432 -1156 10407 -1092
rect 10471 -1156 10487 -1092
rect 10551 -1156 10567 -1092
rect 10631 -1156 10647 -1092
rect 10711 -1156 10727 -1092
rect 10791 -1156 10807 -1092
rect 10871 -1156 10887 -1092
rect 10951 -1156 10967 -1092
rect 11031 -1156 11047 -1092
rect 11111 -1156 11127 -1092
rect 11191 -1156 11207 -1092
rect 11271 -1156 15052 -1092
rect 15116 -1156 15132 -1092
rect 15196 -1156 15212 -1092
rect 15276 -1156 15292 -1092
rect 15356 -1156 15372 -1092
rect 15436 -1156 15452 -1092
rect 15516 -1156 15532 -1092
rect 15596 -1156 15612 -1092
rect 15676 -1156 15692 -1092
rect 15756 -1156 15772 -1092
rect 15836 -1156 15852 -1092
rect 15916 -1156 16891 -1092
rect 16955 -1156 16971 -1092
rect 17035 -1156 17051 -1092
rect 17115 -1156 17131 -1092
rect 17195 -1156 17211 -1092
rect 17275 -1156 17291 -1092
rect 17355 -1156 17371 -1092
rect 17435 -1156 17451 -1092
rect 17515 -1156 17531 -1092
rect 17595 -1156 17611 -1092
rect 17675 -1156 17691 -1092
rect 17755 -1156 17760 -1092
rect 2080 -1173 17760 -1156
rect 2080 -1237 3924 -1173
rect 3988 -1237 4004 -1173
rect 4068 -1237 4084 -1173
rect 4148 -1237 4164 -1173
rect 4228 -1237 4244 -1173
rect 4308 -1237 4324 -1173
rect 4388 -1237 4404 -1173
rect 4468 -1237 4484 -1173
rect 4548 -1237 4564 -1173
rect 4628 -1237 4644 -1173
rect 4708 -1237 4724 -1173
rect 4788 -1237 8568 -1173
rect 8632 -1237 8648 -1173
rect 8712 -1237 8728 -1173
rect 8792 -1237 8808 -1173
rect 8872 -1237 8888 -1173
rect 8952 -1237 8968 -1173
rect 9032 -1237 9048 -1173
rect 9112 -1237 9128 -1173
rect 9192 -1237 9208 -1173
rect 9272 -1237 9288 -1173
rect 9352 -1237 9368 -1173
rect 9432 -1237 10407 -1173
rect 10471 -1237 10487 -1173
rect 10551 -1237 10567 -1173
rect 10631 -1237 10647 -1173
rect 10711 -1237 10727 -1173
rect 10791 -1237 10807 -1173
rect 10871 -1237 10887 -1173
rect 10951 -1237 10967 -1173
rect 11031 -1237 11047 -1173
rect 11111 -1237 11127 -1173
rect 11191 -1237 11207 -1173
rect 11271 -1237 15052 -1173
rect 15116 -1237 15132 -1173
rect 15196 -1237 15212 -1173
rect 15276 -1237 15292 -1173
rect 15356 -1237 15372 -1173
rect 15436 -1237 15452 -1173
rect 15516 -1237 15532 -1173
rect 15596 -1237 15612 -1173
rect 15676 -1237 15692 -1173
rect 15756 -1237 15772 -1173
rect 15836 -1237 15852 -1173
rect 15916 -1237 16891 -1173
rect 16955 -1237 16971 -1173
rect 17035 -1237 17051 -1173
rect 17115 -1237 17131 -1173
rect 17195 -1237 17211 -1173
rect 17275 -1237 17291 -1173
rect 17355 -1237 17371 -1173
rect 17435 -1237 17451 -1173
rect 17515 -1237 17531 -1173
rect 17595 -1237 17611 -1173
rect 17675 -1237 17691 -1173
rect 17755 -1237 17760 -1173
rect 2080 -1254 17760 -1237
rect 2080 -1318 3924 -1254
rect 3988 -1318 4004 -1254
rect 4068 -1318 4084 -1254
rect 4148 -1318 4164 -1254
rect 4228 -1318 4244 -1254
rect 4308 -1318 4324 -1254
rect 4388 -1318 4404 -1254
rect 4468 -1318 4484 -1254
rect 4548 -1318 4564 -1254
rect 4628 -1318 4644 -1254
rect 4708 -1318 4724 -1254
rect 4788 -1318 8568 -1254
rect 8632 -1318 8648 -1254
rect 8712 -1318 8728 -1254
rect 8792 -1318 8808 -1254
rect 8872 -1318 8888 -1254
rect 8952 -1318 8968 -1254
rect 9032 -1318 9048 -1254
rect 9112 -1318 9128 -1254
rect 9192 -1318 9208 -1254
rect 9272 -1318 9288 -1254
rect 9352 -1318 9368 -1254
rect 9432 -1318 10407 -1254
rect 10471 -1318 10487 -1254
rect 10551 -1318 10567 -1254
rect 10631 -1318 10647 -1254
rect 10711 -1318 10727 -1254
rect 10791 -1318 10807 -1254
rect 10871 -1318 10887 -1254
rect 10951 -1318 10967 -1254
rect 11031 -1318 11047 -1254
rect 11111 -1318 11127 -1254
rect 11191 -1318 11207 -1254
rect 11271 -1318 15052 -1254
rect 15116 -1318 15132 -1254
rect 15196 -1318 15212 -1254
rect 15276 -1318 15292 -1254
rect 15356 -1318 15372 -1254
rect 15436 -1318 15452 -1254
rect 15516 -1318 15532 -1254
rect 15596 -1318 15612 -1254
rect 15676 -1318 15692 -1254
rect 15756 -1318 15772 -1254
rect 15836 -1318 15852 -1254
rect 15916 -1318 16891 -1254
rect 16955 -1318 16971 -1254
rect 17035 -1318 17051 -1254
rect 17115 -1318 17131 -1254
rect 17195 -1318 17211 -1254
rect 17275 -1318 17291 -1254
rect 17355 -1318 17371 -1254
rect 17435 -1318 17451 -1254
rect 17515 -1318 17531 -1254
rect 17595 -1318 17611 -1254
rect 17675 -1318 17691 -1254
rect 17755 -1318 17760 -1254
rect 2080 -1335 17760 -1318
rect 2080 -1399 3924 -1335
rect 3988 -1399 4004 -1335
rect 4068 -1399 4084 -1335
rect 4148 -1399 4164 -1335
rect 4228 -1399 4244 -1335
rect 4308 -1399 4324 -1335
rect 4388 -1399 4404 -1335
rect 4468 -1399 4484 -1335
rect 4548 -1399 4564 -1335
rect 4628 -1399 4644 -1335
rect 4708 -1399 4724 -1335
rect 4788 -1399 8568 -1335
rect 8632 -1399 8648 -1335
rect 8712 -1399 8728 -1335
rect 8792 -1399 8808 -1335
rect 8872 -1399 8888 -1335
rect 8952 -1399 8968 -1335
rect 9032 -1399 9048 -1335
rect 9112 -1399 9128 -1335
rect 9192 -1399 9208 -1335
rect 9272 -1399 9288 -1335
rect 9352 -1399 9368 -1335
rect 9432 -1399 10407 -1335
rect 10471 -1399 10487 -1335
rect 10551 -1399 10567 -1335
rect 10631 -1399 10647 -1335
rect 10711 -1399 10727 -1335
rect 10791 -1399 10807 -1335
rect 10871 -1399 10887 -1335
rect 10951 -1399 10967 -1335
rect 11031 -1399 11047 -1335
rect 11111 -1399 11127 -1335
rect 11191 -1399 11207 -1335
rect 11271 -1399 15052 -1335
rect 15116 -1399 15132 -1335
rect 15196 -1399 15212 -1335
rect 15276 -1399 15292 -1335
rect 15356 -1399 15372 -1335
rect 15436 -1399 15452 -1335
rect 15516 -1399 15532 -1335
rect 15596 -1399 15612 -1335
rect 15676 -1399 15692 -1335
rect 15756 -1399 15772 -1335
rect 15836 -1399 15852 -1335
rect 15916 -1399 16891 -1335
rect 16955 -1399 16971 -1335
rect 17035 -1399 17051 -1335
rect 17115 -1399 17131 -1335
rect 17195 -1399 17211 -1335
rect 17275 -1399 17291 -1335
rect 17355 -1399 17371 -1335
rect 17435 -1399 17451 -1335
rect 17515 -1399 17531 -1335
rect 17595 -1399 17611 -1335
rect 17675 -1399 17691 -1335
rect 17755 -1399 17760 -1335
rect 2080 -1416 17760 -1399
rect 2080 -1480 3924 -1416
rect 3988 -1480 4004 -1416
rect 4068 -1480 4084 -1416
rect 4148 -1480 4164 -1416
rect 4228 -1480 4244 -1416
rect 4308 -1480 4324 -1416
rect 4388 -1480 4404 -1416
rect 4468 -1480 4484 -1416
rect 4548 -1480 4564 -1416
rect 4628 -1480 4644 -1416
rect 4708 -1480 4724 -1416
rect 4788 -1480 8568 -1416
rect 8632 -1480 8648 -1416
rect 8712 -1480 8728 -1416
rect 8792 -1480 8808 -1416
rect 8872 -1480 8888 -1416
rect 8952 -1480 8968 -1416
rect 9032 -1480 9048 -1416
rect 9112 -1480 9128 -1416
rect 9192 -1480 9208 -1416
rect 9272 -1480 9288 -1416
rect 9352 -1480 9368 -1416
rect 9432 -1480 10407 -1416
rect 10471 -1480 10487 -1416
rect 10551 -1480 10567 -1416
rect 10631 -1480 10647 -1416
rect 10711 -1480 10727 -1416
rect 10791 -1480 10807 -1416
rect 10871 -1480 10887 -1416
rect 10951 -1480 10967 -1416
rect 11031 -1480 11047 -1416
rect 11111 -1480 11127 -1416
rect 11191 -1480 11207 -1416
rect 11271 -1480 15052 -1416
rect 15116 -1480 15132 -1416
rect 15196 -1480 15212 -1416
rect 15276 -1480 15292 -1416
rect 15356 -1480 15372 -1416
rect 15436 -1480 15452 -1416
rect 15516 -1480 15532 -1416
rect 15596 -1480 15612 -1416
rect 15676 -1480 15692 -1416
rect 15756 -1480 15772 -1416
rect 15836 -1480 15852 -1416
rect 15916 -1480 16891 -1416
rect 16955 -1480 16971 -1416
rect 17035 -1480 17051 -1416
rect 17115 -1480 17131 -1416
rect 17195 -1480 17211 -1416
rect 17275 -1480 17291 -1416
rect 17355 -1480 17371 -1416
rect 17435 -1480 17451 -1416
rect 17515 -1480 17531 -1416
rect 17595 -1480 17611 -1416
rect 17675 -1480 17691 -1416
rect 17755 -1480 17760 -1416
rect 2080 -1497 17760 -1480
rect 2080 -1561 3924 -1497
rect 3988 -1561 4004 -1497
rect 4068 -1561 4084 -1497
rect 4148 -1561 4164 -1497
rect 4228 -1561 4244 -1497
rect 4308 -1561 4324 -1497
rect 4388 -1561 4404 -1497
rect 4468 -1561 4484 -1497
rect 4548 -1561 4564 -1497
rect 4628 -1561 4644 -1497
rect 4708 -1561 4724 -1497
rect 4788 -1561 8568 -1497
rect 8632 -1561 8648 -1497
rect 8712 -1561 8728 -1497
rect 8792 -1561 8808 -1497
rect 8872 -1561 8888 -1497
rect 8952 -1561 8968 -1497
rect 9032 -1561 9048 -1497
rect 9112 -1561 9128 -1497
rect 9192 -1561 9208 -1497
rect 9272 -1561 9288 -1497
rect 9352 -1561 9368 -1497
rect 9432 -1561 10407 -1497
rect 10471 -1561 10487 -1497
rect 10551 -1561 10567 -1497
rect 10631 -1561 10647 -1497
rect 10711 -1561 10727 -1497
rect 10791 -1561 10807 -1497
rect 10871 -1561 10887 -1497
rect 10951 -1561 10967 -1497
rect 11031 -1561 11047 -1497
rect 11111 -1561 11127 -1497
rect 11191 -1561 11207 -1497
rect 11271 -1561 15052 -1497
rect 15116 -1561 15132 -1497
rect 15196 -1561 15212 -1497
rect 15276 -1561 15292 -1497
rect 15356 -1561 15372 -1497
rect 15436 -1561 15452 -1497
rect 15516 -1561 15532 -1497
rect 15596 -1561 15612 -1497
rect 15676 -1561 15692 -1497
rect 15756 -1561 15772 -1497
rect 15836 -1561 15852 -1497
rect 15916 -1561 16891 -1497
rect 16955 -1561 16971 -1497
rect 17035 -1561 17051 -1497
rect 17115 -1561 17131 -1497
rect 17195 -1561 17211 -1497
rect 17275 -1561 17291 -1497
rect 17355 -1561 17371 -1497
rect 17435 -1561 17451 -1497
rect 17515 -1561 17531 -1497
rect 17595 -1561 17611 -1497
rect 17675 -1561 17691 -1497
rect 17755 -1561 17760 -1497
rect 2080 -1578 17760 -1561
rect 2080 -1642 3924 -1578
rect 3988 -1642 4004 -1578
rect 4068 -1642 4084 -1578
rect 4148 -1642 4164 -1578
rect 4228 -1642 4244 -1578
rect 4308 -1642 4324 -1578
rect 4388 -1642 4404 -1578
rect 4468 -1642 4484 -1578
rect 4548 -1642 4564 -1578
rect 4628 -1642 4644 -1578
rect 4708 -1642 4724 -1578
rect 4788 -1642 8568 -1578
rect 8632 -1642 8648 -1578
rect 8712 -1642 8728 -1578
rect 8792 -1642 8808 -1578
rect 8872 -1642 8888 -1578
rect 8952 -1642 8968 -1578
rect 9032 -1642 9048 -1578
rect 9112 -1642 9128 -1578
rect 9192 -1642 9208 -1578
rect 9272 -1642 9288 -1578
rect 9352 -1642 9368 -1578
rect 9432 -1642 10407 -1578
rect 10471 -1642 10487 -1578
rect 10551 -1642 10567 -1578
rect 10631 -1642 10647 -1578
rect 10711 -1642 10727 -1578
rect 10791 -1642 10807 -1578
rect 10871 -1642 10887 -1578
rect 10951 -1642 10967 -1578
rect 11031 -1642 11047 -1578
rect 11111 -1642 11127 -1578
rect 11191 -1642 11207 -1578
rect 11271 -1642 15052 -1578
rect 15116 -1642 15132 -1578
rect 15196 -1642 15212 -1578
rect 15276 -1642 15292 -1578
rect 15356 -1642 15372 -1578
rect 15436 -1642 15452 -1578
rect 15516 -1642 15532 -1578
rect 15596 -1642 15612 -1578
rect 15676 -1642 15692 -1578
rect 15756 -1642 15772 -1578
rect 15836 -1642 15852 -1578
rect 15916 -1642 16891 -1578
rect 16955 -1642 16971 -1578
rect 17035 -1642 17051 -1578
rect 17115 -1642 17131 -1578
rect 17195 -1642 17211 -1578
rect 17275 -1642 17291 -1578
rect 17355 -1642 17371 -1578
rect 17435 -1642 17451 -1578
rect 17515 -1642 17531 -1578
rect 17595 -1642 17611 -1578
rect 17675 -1642 17691 -1578
rect 17755 -1642 17760 -1578
rect 2080 -1659 17760 -1642
rect 2080 -1723 3924 -1659
rect 3988 -1723 4004 -1659
rect 4068 -1723 4084 -1659
rect 4148 -1723 4164 -1659
rect 4228 -1723 4244 -1659
rect 4308 -1723 4324 -1659
rect 4388 -1723 4404 -1659
rect 4468 -1723 4484 -1659
rect 4548 -1723 4564 -1659
rect 4628 -1723 4644 -1659
rect 4708 -1723 4724 -1659
rect 4788 -1723 8568 -1659
rect 8632 -1723 8648 -1659
rect 8712 -1723 8728 -1659
rect 8792 -1723 8808 -1659
rect 8872 -1723 8888 -1659
rect 8952 -1723 8968 -1659
rect 9032 -1723 9048 -1659
rect 9112 -1723 9128 -1659
rect 9192 -1723 9208 -1659
rect 9272 -1723 9288 -1659
rect 9352 -1723 9368 -1659
rect 9432 -1723 10407 -1659
rect 10471 -1723 10487 -1659
rect 10551 -1723 10567 -1659
rect 10631 -1723 10647 -1659
rect 10711 -1723 10727 -1659
rect 10791 -1723 10807 -1659
rect 10871 -1723 10887 -1659
rect 10951 -1723 10967 -1659
rect 11031 -1723 11047 -1659
rect 11111 -1723 11127 -1659
rect 11191 -1723 11207 -1659
rect 11271 -1723 15052 -1659
rect 15116 -1723 15132 -1659
rect 15196 -1723 15212 -1659
rect 15276 -1723 15292 -1659
rect 15356 -1723 15372 -1659
rect 15436 -1723 15452 -1659
rect 15516 -1723 15532 -1659
rect 15596 -1723 15612 -1659
rect 15676 -1723 15692 -1659
rect 15756 -1723 15772 -1659
rect 15836 -1723 15852 -1659
rect 15916 -1723 16891 -1659
rect 16955 -1723 16971 -1659
rect 17035 -1723 17051 -1659
rect 17115 -1723 17131 -1659
rect 17195 -1723 17211 -1659
rect 17275 -1723 17291 -1659
rect 17355 -1723 17371 -1659
rect 17435 -1723 17451 -1659
rect 17515 -1723 17531 -1659
rect 17595 -1723 17611 -1659
rect 17675 -1723 17691 -1659
rect 17755 -1723 17760 -1659
rect 2080 -1740 17760 -1723
rect 2080 -1804 3924 -1740
rect 3988 -1804 4004 -1740
rect 4068 -1804 4084 -1740
rect 4148 -1804 4164 -1740
rect 4228 -1804 4244 -1740
rect 4308 -1804 4324 -1740
rect 4388 -1804 4404 -1740
rect 4468 -1804 4484 -1740
rect 4548 -1804 4564 -1740
rect 4628 -1804 4644 -1740
rect 4708 -1804 4724 -1740
rect 4788 -1804 8568 -1740
rect 8632 -1804 8648 -1740
rect 8712 -1804 8728 -1740
rect 8792 -1804 8808 -1740
rect 8872 -1804 8888 -1740
rect 8952 -1804 8968 -1740
rect 9032 -1804 9048 -1740
rect 9112 -1804 9128 -1740
rect 9192 -1804 9208 -1740
rect 9272 -1804 9288 -1740
rect 9352 -1804 9368 -1740
rect 9432 -1804 10407 -1740
rect 10471 -1804 10487 -1740
rect 10551 -1804 10567 -1740
rect 10631 -1804 10647 -1740
rect 10711 -1804 10727 -1740
rect 10791 -1804 10807 -1740
rect 10871 -1804 10887 -1740
rect 10951 -1804 10967 -1740
rect 11031 -1804 11047 -1740
rect 11111 -1804 11127 -1740
rect 11191 -1804 11207 -1740
rect 11271 -1804 15052 -1740
rect 15116 -1804 15132 -1740
rect 15196 -1804 15212 -1740
rect 15276 -1804 15292 -1740
rect 15356 -1804 15372 -1740
rect 15436 -1804 15452 -1740
rect 15516 -1804 15532 -1740
rect 15596 -1804 15612 -1740
rect 15676 -1804 15692 -1740
rect 15756 -1804 15772 -1740
rect 15836 -1804 15852 -1740
rect 15916 -1804 16891 -1740
rect 16955 -1804 16971 -1740
rect 17035 -1804 17051 -1740
rect 17115 -1804 17131 -1740
rect 17195 -1804 17211 -1740
rect 17275 -1804 17291 -1740
rect 17355 -1804 17371 -1740
rect 17435 -1804 17451 -1740
rect 17515 -1804 17531 -1740
rect 17595 -1804 17611 -1740
rect 17675 -1804 17691 -1740
rect 17755 -1804 17760 -1740
rect 2080 -1821 17760 -1804
rect 2080 -1885 3924 -1821
rect 3988 -1885 4004 -1821
rect 4068 -1885 4084 -1821
rect 4148 -1885 4164 -1821
rect 4228 -1885 4244 -1821
rect 4308 -1885 4324 -1821
rect 4388 -1885 4404 -1821
rect 4468 -1885 4484 -1821
rect 4548 -1885 4564 -1821
rect 4628 -1885 4644 -1821
rect 4708 -1885 4724 -1821
rect 4788 -1885 8568 -1821
rect 8632 -1885 8648 -1821
rect 8712 -1885 8728 -1821
rect 8792 -1885 8808 -1821
rect 8872 -1885 8888 -1821
rect 8952 -1885 8968 -1821
rect 9032 -1885 9048 -1821
rect 9112 -1885 9128 -1821
rect 9192 -1885 9208 -1821
rect 9272 -1885 9288 -1821
rect 9352 -1885 9368 -1821
rect 9432 -1885 10407 -1821
rect 10471 -1885 10487 -1821
rect 10551 -1885 10567 -1821
rect 10631 -1885 10647 -1821
rect 10711 -1885 10727 -1821
rect 10791 -1885 10807 -1821
rect 10871 -1885 10887 -1821
rect 10951 -1885 10967 -1821
rect 11031 -1885 11047 -1821
rect 11111 -1885 11127 -1821
rect 11191 -1885 11207 -1821
rect 11271 -1885 15052 -1821
rect 15116 -1885 15132 -1821
rect 15196 -1885 15212 -1821
rect 15276 -1885 15292 -1821
rect 15356 -1885 15372 -1821
rect 15436 -1885 15452 -1821
rect 15516 -1885 15532 -1821
rect 15596 -1885 15612 -1821
rect 15676 -1885 15692 -1821
rect 15756 -1885 15772 -1821
rect 15836 -1885 15852 -1821
rect 15916 -1885 16891 -1821
rect 16955 -1885 16971 -1821
rect 17035 -1885 17051 -1821
rect 17115 -1885 17131 -1821
rect 17195 -1885 17211 -1821
rect 17275 -1885 17291 -1821
rect 17355 -1885 17371 -1821
rect 17435 -1885 17451 -1821
rect 17515 -1885 17531 -1821
rect 17595 -1885 17611 -1821
rect 17675 -1885 17691 -1821
rect 17755 -1885 17760 -1821
rect 2080 -1902 17760 -1885
rect 2080 -1966 3924 -1902
rect 3988 -1966 4004 -1902
rect 4068 -1966 4084 -1902
rect 4148 -1966 4164 -1902
rect 4228 -1966 4244 -1902
rect 4308 -1966 4324 -1902
rect 4388 -1966 4404 -1902
rect 4468 -1966 4484 -1902
rect 4548 -1966 4564 -1902
rect 4628 -1966 4644 -1902
rect 4708 -1966 4724 -1902
rect 4788 -1966 8568 -1902
rect 8632 -1966 8648 -1902
rect 8712 -1966 8728 -1902
rect 8792 -1966 8808 -1902
rect 8872 -1966 8888 -1902
rect 8952 -1966 8968 -1902
rect 9032 -1966 9048 -1902
rect 9112 -1966 9128 -1902
rect 9192 -1966 9208 -1902
rect 9272 -1966 9288 -1902
rect 9352 -1966 9368 -1902
rect 9432 -1966 10407 -1902
rect 10471 -1966 10487 -1902
rect 10551 -1966 10567 -1902
rect 10631 -1966 10647 -1902
rect 10711 -1966 10727 -1902
rect 10791 -1966 10807 -1902
rect 10871 -1966 10887 -1902
rect 10951 -1966 10967 -1902
rect 11031 -1966 11047 -1902
rect 11111 -1966 11127 -1902
rect 11191 -1966 11207 -1902
rect 11271 -1966 15052 -1902
rect 15116 -1966 15132 -1902
rect 15196 -1966 15212 -1902
rect 15276 -1966 15292 -1902
rect 15356 -1966 15372 -1902
rect 15436 -1966 15452 -1902
rect 15516 -1966 15532 -1902
rect 15596 -1966 15612 -1902
rect 15676 -1966 15692 -1902
rect 15756 -1966 15772 -1902
rect 15836 -1966 15852 -1902
rect 15916 -1966 16891 -1902
rect 16955 -1966 16971 -1902
rect 17035 -1966 17051 -1902
rect 17115 -1966 17131 -1902
rect 17195 -1966 17211 -1902
rect 17275 -1966 17291 -1902
rect 17355 -1966 17371 -1902
rect 17435 -1966 17451 -1902
rect 17515 -1966 17531 -1902
rect 17595 -1966 17611 -1902
rect 17675 -1966 17691 -1902
rect 17755 -1966 17760 -1902
rect 2080 -1983 17760 -1966
rect 2080 -2047 3924 -1983
rect 3988 -2047 4004 -1983
rect 4068 -2047 4084 -1983
rect 4148 -2047 4164 -1983
rect 4228 -2047 4244 -1983
rect 4308 -2047 4324 -1983
rect 4388 -2047 4404 -1983
rect 4468 -2047 4484 -1983
rect 4548 -2047 4564 -1983
rect 4628 -2047 4644 -1983
rect 4708 -2047 4724 -1983
rect 4788 -2047 8568 -1983
rect 8632 -2047 8648 -1983
rect 8712 -2047 8728 -1983
rect 8792 -2047 8808 -1983
rect 8872 -2047 8888 -1983
rect 8952 -2047 8968 -1983
rect 9032 -2047 9048 -1983
rect 9112 -2047 9128 -1983
rect 9192 -2047 9208 -1983
rect 9272 -2047 9288 -1983
rect 9352 -2047 9368 -1983
rect 9432 -2047 10407 -1983
rect 10471 -2047 10487 -1983
rect 10551 -2047 10567 -1983
rect 10631 -2047 10647 -1983
rect 10711 -2047 10727 -1983
rect 10791 -2047 10807 -1983
rect 10871 -2047 10887 -1983
rect 10951 -2047 10967 -1983
rect 11031 -2047 11047 -1983
rect 11111 -2047 11127 -1983
rect 11191 -2047 11207 -1983
rect 11271 -2047 15052 -1983
rect 15116 -2047 15132 -1983
rect 15196 -2047 15212 -1983
rect 15276 -2047 15292 -1983
rect 15356 -2047 15372 -1983
rect 15436 -2047 15452 -1983
rect 15516 -2047 15532 -1983
rect 15596 -2047 15612 -1983
rect 15676 -2047 15692 -1983
rect 15756 -2047 15772 -1983
rect 15836 -2047 15852 -1983
rect 15916 -2047 16891 -1983
rect 16955 -2047 16971 -1983
rect 17035 -2047 17051 -1983
rect 17115 -2047 17131 -1983
rect 17195 -2047 17211 -1983
rect 17275 -2047 17291 -1983
rect 17355 -2047 17371 -1983
rect 17435 -2047 17451 -1983
rect 17515 -2047 17531 -1983
rect 17595 -2047 17611 -1983
rect 17675 -2047 17691 -1983
rect 17755 -2047 17760 -1983
rect 2080 -2064 17760 -2047
rect 2080 -2128 3924 -2064
rect 3988 -2128 4004 -2064
rect 4068 -2128 4084 -2064
rect 4148 -2128 4164 -2064
rect 4228 -2128 4244 -2064
rect 4308 -2128 4324 -2064
rect 4388 -2128 4404 -2064
rect 4468 -2128 4484 -2064
rect 4548 -2128 4564 -2064
rect 4628 -2128 4644 -2064
rect 4708 -2128 4724 -2064
rect 4788 -2128 8568 -2064
rect 8632 -2128 8648 -2064
rect 8712 -2128 8728 -2064
rect 8792 -2128 8808 -2064
rect 8872 -2128 8888 -2064
rect 8952 -2128 8968 -2064
rect 9032 -2128 9048 -2064
rect 9112 -2128 9128 -2064
rect 9192 -2128 9208 -2064
rect 9272 -2128 9288 -2064
rect 9352 -2128 9368 -2064
rect 9432 -2128 10407 -2064
rect 10471 -2128 10487 -2064
rect 10551 -2128 10567 -2064
rect 10631 -2128 10647 -2064
rect 10711 -2128 10727 -2064
rect 10791 -2128 10807 -2064
rect 10871 -2128 10887 -2064
rect 10951 -2128 10967 -2064
rect 11031 -2128 11047 -2064
rect 11111 -2128 11127 -2064
rect 11191 -2128 11207 -2064
rect 11271 -2128 15052 -2064
rect 15116 -2128 15132 -2064
rect 15196 -2128 15212 -2064
rect 15276 -2128 15292 -2064
rect 15356 -2128 15372 -2064
rect 15436 -2128 15452 -2064
rect 15516 -2128 15532 -2064
rect 15596 -2128 15612 -2064
rect 15676 -2128 15692 -2064
rect 15756 -2128 15772 -2064
rect 15836 -2128 15852 -2064
rect 15916 -2128 16891 -2064
rect 16955 -2128 16971 -2064
rect 17035 -2128 17051 -2064
rect 17115 -2128 17131 -2064
rect 17195 -2128 17211 -2064
rect 17275 -2128 17291 -2064
rect 17355 -2128 17371 -2064
rect 17435 -2128 17451 -2064
rect 17515 -2128 17531 -2064
rect 17595 -2128 17611 -2064
rect 17675 -2128 17691 -2064
rect 17755 -2128 17760 -2064
rect 2080 -2145 17760 -2128
rect 2080 -2209 3924 -2145
rect 3988 -2209 4004 -2145
rect 4068 -2209 4084 -2145
rect 4148 -2209 4164 -2145
rect 4228 -2209 4244 -2145
rect 4308 -2209 4324 -2145
rect 4388 -2209 4404 -2145
rect 4468 -2209 4484 -2145
rect 4548 -2209 4564 -2145
rect 4628 -2209 4644 -2145
rect 4708 -2209 4724 -2145
rect 4788 -2209 8568 -2145
rect 8632 -2209 8648 -2145
rect 8712 -2209 8728 -2145
rect 8792 -2209 8808 -2145
rect 8872 -2209 8888 -2145
rect 8952 -2209 8968 -2145
rect 9032 -2209 9048 -2145
rect 9112 -2209 9128 -2145
rect 9192 -2209 9208 -2145
rect 9272 -2209 9288 -2145
rect 9352 -2209 9368 -2145
rect 9432 -2209 10407 -2145
rect 10471 -2209 10487 -2145
rect 10551 -2209 10567 -2145
rect 10631 -2209 10647 -2145
rect 10711 -2209 10727 -2145
rect 10791 -2209 10807 -2145
rect 10871 -2209 10887 -2145
rect 10951 -2209 10967 -2145
rect 11031 -2209 11047 -2145
rect 11111 -2209 11127 -2145
rect 11191 -2209 11207 -2145
rect 11271 -2209 15052 -2145
rect 15116 -2209 15132 -2145
rect 15196 -2209 15212 -2145
rect 15276 -2209 15292 -2145
rect 15356 -2209 15372 -2145
rect 15436 -2209 15452 -2145
rect 15516 -2209 15532 -2145
rect 15596 -2209 15612 -2145
rect 15676 -2209 15692 -2145
rect 15756 -2209 15772 -2145
rect 15836 -2209 15852 -2145
rect 15916 -2209 16891 -2145
rect 16955 -2209 16971 -2145
rect 17035 -2209 17051 -2145
rect 17115 -2209 17131 -2145
rect 17195 -2209 17211 -2145
rect 17275 -2209 17291 -2145
rect 17355 -2209 17371 -2145
rect 17435 -2209 17451 -2145
rect 17515 -2209 17531 -2145
rect 17595 -2209 17611 -2145
rect 17675 -2209 17691 -2145
rect 17755 -2209 17760 -2145
rect 2080 -2226 17760 -2209
rect 2080 -2290 3924 -2226
rect 3988 -2290 4004 -2226
rect 4068 -2290 4084 -2226
rect 4148 -2290 4164 -2226
rect 4228 -2290 4244 -2226
rect 4308 -2290 4324 -2226
rect 4388 -2290 4404 -2226
rect 4468 -2290 4484 -2226
rect 4548 -2290 4564 -2226
rect 4628 -2290 4644 -2226
rect 4708 -2290 4724 -2226
rect 4788 -2290 8568 -2226
rect 8632 -2290 8648 -2226
rect 8712 -2290 8728 -2226
rect 8792 -2290 8808 -2226
rect 8872 -2290 8888 -2226
rect 8952 -2290 8968 -2226
rect 9032 -2290 9048 -2226
rect 9112 -2290 9128 -2226
rect 9192 -2290 9208 -2226
rect 9272 -2290 9288 -2226
rect 9352 -2290 9368 -2226
rect 9432 -2290 10407 -2226
rect 10471 -2290 10487 -2226
rect 10551 -2290 10567 -2226
rect 10631 -2290 10647 -2226
rect 10711 -2290 10727 -2226
rect 10791 -2290 10807 -2226
rect 10871 -2290 10887 -2226
rect 10951 -2290 10967 -2226
rect 11031 -2290 11047 -2226
rect 11111 -2290 11127 -2226
rect 11191 -2290 11207 -2226
rect 11271 -2290 15052 -2226
rect 15116 -2290 15132 -2226
rect 15196 -2290 15212 -2226
rect 15276 -2290 15292 -2226
rect 15356 -2290 15372 -2226
rect 15436 -2290 15452 -2226
rect 15516 -2290 15532 -2226
rect 15596 -2290 15612 -2226
rect 15676 -2290 15692 -2226
rect 15756 -2290 15772 -2226
rect 15836 -2290 15852 -2226
rect 15916 -2290 16891 -2226
rect 16955 -2290 16971 -2226
rect 17035 -2290 17051 -2226
rect 17115 -2290 17131 -2226
rect 17195 -2290 17211 -2226
rect 17275 -2290 17291 -2226
rect 17355 -2290 17371 -2226
rect 17435 -2290 17451 -2226
rect 17515 -2290 17531 -2226
rect 17595 -2290 17611 -2226
rect 17675 -2290 17691 -2226
rect 17755 -2290 17760 -2226
rect 2080 -2307 17760 -2290
rect 2080 -2371 3924 -2307
rect 3988 -2371 4004 -2307
rect 4068 -2371 4084 -2307
rect 4148 -2371 4164 -2307
rect 4228 -2371 4244 -2307
rect 4308 -2371 4324 -2307
rect 4388 -2371 4404 -2307
rect 4468 -2371 4484 -2307
rect 4548 -2371 4564 -2307
rect 4628 -2371 4644 -2307
rect 4708 -2371 4724 -2307
rect 4788 -2371 8568 -2307
rect 8632 -2371 8648 -2307
rect 8712 -2371 8728 -2307
rect 8792 -2371 8808 -2307
rect 8872 -2371 8888 -2307
rect 8952 -2371 8968 -2307
rect 9032 -2371 9048 -2307
rect 9112 -2371 9128 -2307
rect 9192 -2371 9208 -2307
rect 9272 -2371 9288 -2307
rect 9352 -2371 9368 -2307
rect 9432 -2371 10407 -2307
rect 10471 -2371 10487 -2307
rect 10551 -2371 10567 -2307
rect 10631 -2371 10647 -2307
rect 10711 -2371 10727 -2307
rect 10791 -2371 10807 -2307
rect 10871 -2371 10887 -2307
rect 10951 -2371 10967 -2307
rect 11031 -2371 11047 -2307
rect 11111 -2371 11127 -2307
rect 11191 -2371 11207 -2307
rect 11271 -2371 15052 -2307
rect 15116 -2371 15132 -2307
rect 15196 -2371 15212 -2307
rect 15276 -2371 15292 -2307
rect 15356 -2371 15372 -2307
rect 15436 -2371 15452 -2307
rect 15516 -2371 15532 -2307
rect 15596 -2371 15612 -2307
rect 15676 -2371 15692 -2307
rect 15756 -2371 15772 -2307
rect 15836 -2371 15852 -2307
rect 15916 -2371 16891 -2307
rect 16955 -2371 16971 -2307
rect 17035 -2371 17051 -2307
rect 17115 -2371 17131 -2307
rect 17195 -2371 17211 -2307
rect 17275 -2371 17291 -2307
rect 17355 -2371 17371 -2307
rect 17435 -2371 17451 -2307
rect 17515 -2371 17531 -2307
rect 17595 -2371 17611 -2307
rect 17675 -2371 17691 -2307
rect 17755 -2371 17760 -2307
rect 2080 -2388 17760 -2371
rect 2080 -2452 3924 -2388
rect 3988 -2452 4004 -2388
rect 4068 -2452 4084 -2388
rect 4148 -2452 4164 -2388
rect 4228 -2452 4244 -2388
rect 4308 -2452 4324 -2388
rect 4388 -2452 4404 -2388
rect 4468 -2452 4484 -2388
rect 4548 -2452 4564 -2388
rect 4628 -2452 4644 -2388
rect 4708 -2452 4724 -2388
rect 4788 -2452 8568 -2388
rect 8632 -2452 8648 -2388
rect 8712 -2452 8728 -2388
rect 8792 -2452 8808 -2388
rect 8872 -2452 8888 -2388
rect 8952 -2452 8968 -2388
rect 9032 -2452 9048 -2388
rect 9112 -2452 9128 -2388
rect 9192 -2452 9208 -2388
rect 9272 -2452 9288 -2388
rect 9352 -2452 9368 -2388
rect 9432 -2452 10407 -2388
rect 10471 -2452 10487 -2388
rect 10551 -2452 10567 -2388
rect 10631 -2452 10647 -2388
rect 10711 -2452 10727 -2388
rect 10791 -2452 10807 -2388
rect 10871 -2452 10887 -2388
rect 10951 -2452 10967 -2388
rect 11031 -2452 11047 -2388
rect 11111 -2452 11127 -2388
rect 11191 -2452 11207 -2388
rect 11271 -2452 15052 -2388
rect 15116 -2452 15132 -2388
rect 15196 -2452 15212 -2388
rect 15276 -2452 15292 -2388
rect 15356 -2452 15372 -2388
rect 15436 -2452 15452 -2388
rect 15516 -2452 15532 -2388
rect 15596 -2452 15612 -2388
rect 15676 -2452 15692 -2388
rect 15756 -2452 15772 -2388
rect 15836 -2452 15852 -2388
rect 15916 -2452 16891 -2388
rect 16955 -2452 16971 -2388
rect 17035 -2452 17051 -2388
rect 17115 -2452 17131 -2388
rect 17195 -2452 17211 -2388
rect 17275 -2452 17291 -2388
rect 17355 -2452 17371 -2388
rect 17435 -2452 17451 -2388
rect 17515 -2452 17531 -2388
rect 17595 -2452 17611 -2388
rect 17675 -2452 17691 -2388
rect 17755 -2452 17760 -2388
rect 2080 -2469 17760 -2452
rect 2080 -2533 3924 -2469
rect 3988 -2533 4004 -2469
rect 4068 -2533 4084 -2469
rect 4148 -2533 4164 -2469
rect 4228 -2533 4244 -2469
rect 4308 -2533 4324 -2469
rect 4388 -2533 4404 -2469
rect 4468 -2533 4484 -2469
rect 4548 -2533 4564 -2469
rect 4628 -2533 4644 -2469
rect 4708 -2533 4724 -2469
rect 4788 -2533 8568 -2469
rect 8632 -2533 8648 -2469
rect 8712 -2533 8728 -2469
rect 8792 -2533 8808 -2469
rect 8872 -2533 8888 -2469
rect 8952 -2533 8968 -2469
rect 9032 -2533 9048 -2469
rect 9112 -2533 9128 -2469
rect 9192 -2533 9208 -2469
rect 9272 -2533 9288 -2469
rect 9352 -2533 9368 -2469
rect 9432 -2533 10407 -2469
rect 10471 -2533 10487 -2469
rect 10551 -2533 10567 -2469
rect 10631 -2533 10647 -2469
rect 10711 -2533 10727 -2469
rect 10791 -2533 10807 -2469
rect 10871 -2533 10887 -2469
rect 10951 -2533 10967 -2469
rect 11031 -2533 11047 -2469
rect 11111 -2533 11127 -2469
rect 11191 -2533 11207 -2469
rect 11271 -2533 15052 -2469
rect 15116 -2533 15132 -2469
rect 15196 -2533 15212 -2469
rect 15276 -2533 15292 -2469
rect 15356 -2533 15372 -2469
rect 15436 -2533 15452 -2469
rect 15516 -2533 15532 -2469
rect 15596 -2533 15612 -2469
rect 15676 -2533 15692 -2469
rect 15756 -2533 15772 -2469
rect 15836 -2533 15852 -2469
rect 15916 -2533 16891 -2469
rect 16955 -2533 16971 -2469
rect 17035 -2533 17051 -2469
rect 17115 -2533 17131 -2469
rect 17195 -2533 17211 -2469
rect 17275 -2533 17291 -2469
rect 17355 -2533 17371 -2469
rect 17435 -2533 17451 -2469
rect 17515 -2533 17531 -2469
rect 17595 -2533 17611 -2469
rect 17675 -2533 17691 -2469
rect 17755 -2533 17760 -2469
rect 2080 -2550 17760 -2533
rect 2080 -2614 3924 -2550
rect 3988 -2614 4004 -2550
rect 4068 -2614 4084 -2550
rect 4148 -2614 4164 -2550
rect 4228 -2614 4244 -2550
rect 4308 -2614 4324 -2550
rect 4388 -2614 4404 -2550
rect 4468 -2614 4484 -2550
rect 4548 -2614 4564 -2550
rect 4628 -2614 4644 -2550
rect 4708 -2614 4724 -2550
rect 4788 -2614 8568 -2550
rect 8632 -2614 8648 -2550
rect 8712 -2614 8728 -2550
rect 8792 -2614 8808 -2550
rect 8872 -2614 8888 -2550
rect 8952 -2614 8968 -2550
rect 9032 -2614 9048 -2550
rect 9112 -2614 9128 -2550
rect 9192 -2614 9208 -2550
rect 9272 -2614 9288 -2550
rect 9352 -2614 9368 -2550
rect 9432 -2614 10407 -2550
rect 10471 -2614 10487 -2550
rect 10551 -2614 10567 -2550
rect 10631 -2614 10647 -2550
rect 10711 -2614 10727 -2550
rect 10791 -2614 10807 -2550
rect 10871 -2614 10887 -2550
rect 10951 -2614 10967 -2550
rect 11031 -2614 11047 -2550
rect 11111 -2614 11127 -2550
rect 11191 -2614 11207 -2550
rect 11271 -2614 15052 -2550
rect 15116 -2614 15132 -2550
rect 15196 -2614 15212 -2550
rect 15276 -2614 15292 -2550
rect 15356 -2614 15372 -2550
rect 15436 -2614 15452 -2550
rect 15516 -2614 15532 -2550
rect 15596 -2614 15612 -2550
rect 15676 -2614 15692 -2550
rect 15756 -2614 15772 -2550
rect 15836 -2614 15852 -2550
rect 15916 -2614 16891 -2550
rect 16955 -2614 16971 -2550
rect 17035 -2614 17051 -2550
rect 17115 -2614 17131 -2550
rect 17195 -2614 17211 -2550
rect 17275 -2614 17291 -2550
rect 17355 -2614 17371 -2550
rect 17435 -2614 17451 -2550
rect 17515 -2614 17531 -2550
rect 17595 -2614 17611 -2550
rect 17675 -2614 17691 -2550
rect 17755 -2614 17760 -2550
rect 2080 -2615 17760 -2614
rect 4882 -2936 5108 -2935
rect 4882 -3000 4883 -2936
rect 4947 -3000 4963 -2936
rect 5027 -3000 5043 -2936
rect 5107 -3000 5108 -2936
rect 4882 -3027 5108 -3000
rect 4882 -3091 4883 -3027
rect 4947 -3091 4963 -3027
rect 5027 -3091 5043 -3027
rect 5107 -3091 5108 -3027
rect 4882 -3119 5108 -3091
rect 4882 -3183 4883 -3119
rect 4947 -3183 4963 -3119
rect 5027 -3183 5043 -3119
rect 5107 -3183 5108 -3119
rect 4882 -3211 5108 -3183
rect 4882 -3275 4883 -3211
rect 4947 -3275 4963 -3211
rect 5027 -3275 5043 -3211
rect 5107 -3275 5108 -3211
rect 4882 -3276 5108 -3275
rect 5716 -2936 5942 -2935
rect 5716 -3000 5717 -2936
rect 5781 -3000 5797 -2936
rect 5861 -3000 5877 -2936
rect 5941 -3000 5942 -2936
rect 5716 -3027 5942 -3000
rect 5716 -3091 5717 -3027
rect 5781 -3091 5797 -3027
rect 5861 -3091 5877 -3027
rect 5941 -3091 5942 -3027
rect 5716 -3119 5942 -3091
rect 5716 -3183 5717 -3119
rect 5781 -3183 5797 -3119
rect 5861 -3183 5877 -3119
rect 5941 -3183 5942 -3119
rect 5716 -3211 5942 -3183
rect 5716 -3275 5717 -3211
rect 5781 -3275 5797 -3211
rect 5861 -3275 5877 -3211
rect 5941 -3275 5942 -3211
rect 5716 -3276 5942 -3275
rect 6490 -2936 6864 -2935
rect 6490 -3000 6492 -2936
rect 6556 -3000 6594 -2936
rect 6658 -3000 6696 -2936
rect 6760 -3000 6798 -2936
rect 6862 -3000 6864 -2936
rect 6490 -3016 6864 -3000
rect 6490 -3080 6492 -3016
rect 6556 -3080 6594 -3016
rect 6658 -3080 6696 -3016
rect 6760 -3080 6798 -3016
rect 6862 -3080 6864 -3016
rect 6490 -3096 6864 -3080
rect 6490 -3160 6492 -3096
rect 6556 -3160 6594 -3096
rect 6658 -3160 6696 -3096
rect 6760 -3160 6798 -3096
rect 6862 -3160 6864 -3096
rect 6490 -3176 6864 -3160
rect 6490 -3240 6492 -3176
rect 6556 -3240 6594 -3176
rect 6658 -3240 6696 -3176
rect 6760 -3240 6798 -3176
rect 6862 -3240 6864 -3176
rect 6490 -3256 6864 -3240
rect 6490 -3320 6492 -3256
rect 6556 -3320 6594 -3256
rect 6658 -3320 6696 -3256
rect 6760 -3320 6798 -3256
rect 6862 -3320 6864 -3256
rect 6490 -3337 6864 -3320
rect 6490 -3401 6492 -3337
rect 6556 -3401 6594 -3337
rect 6658 -3401 6696 -3337
rect 6760 -3401 6798 -3337
rect 6862 -3401 6864 -3337
rect 6490 -3418 6864 -3401
rect 6490 -3482 6492 -3418
rect 6556 -3482 6594 -3418
rect 6658 -3482 6696 -3418
rect 6760 -3482 6798 -3418
rect 6862 -3482 6864 -3418
rect 6490 -3499 6864 -3482
rect 6490 -3563 6492 -3499
rect 6556 -3563 6594 -3499
rect 6658 -3563 6696 -3499
rect 6760 -3563 6798 -3499
rect 6862 -3563 6864 -3499
rect 6490 -3580 6864 -3563
rect 6490 -3644 6492 -3580
rect 6556 -3644 6594 -3580
rect 6658 -3644 6696 -3580
rect 6760 -3644 6798 -3580
rect 6862 -3644 6864 -3580
rect 6490 -3661 6864 -3644
rect 6490 -3725 6492 -3661
rect 6556 -3725 6594 -3661
rect 6658 -3725 6696 -3661
rect 6760 -3725 6798 -3661
rect 6862 -3725 6864 -3661
rect 6490 -3742 6864 -3725
rect 9539 -2936 9765 -2935
rect 9539 -3000 9540 -2936
rect 9604 -3000 9620 -2936
rect 9684 -3000 9700 -2936
rect 9764 -3000 9765 -2936
rect 9539 -3017 9765 -3000
rect 9539 -3081 9540 -3017
rect 9604 -3081 9620 -3017
rect 9684 -3081 9700 -3017
rect 9764 -3081 9765 -3017
rect 9539 -3098 9765 -3081
rect 9539 -3162 9540 -3098
rect 9604 -3162 9620 -3098
rect 9684 -3162 9700 -3098
rect 9764 -3162 9765 -3098
rect 9539 -3179 9765 -3162
rect 9539 -3243 9540 -3179
rect 9604 -3243 9620 -3179
rect 9684 -3243 9700 -3179
rect 9764 -3243 9765 -3179
rect 9539 -3260 9765 -3243
rect 9539 -3324 9540 -3260
rect 9604 -3324 9620 -3260
rect 9684 -3324 9700 -3260
rect 9764 -3324 9765 -3260
rect 9539 -3341 9765 -3324
rect 9539 -3405 9540 -3341
rect 9604 -3405 9620 -3341
rect 9684 -3405 9700 -3341
rect 9764 -3405 9765 -3341
rect 9539 -3423 9765 -3405
rect 9539 -3487 9540 -3423
rect 9604 -3487 9620 -3423
rect 9684 -3487 9700 -3423
rect 9764 -3487 9765 -3423
rect 9539 -3505 9765 -3487
rect 9539 -3569 9540 -3505
rect 9604 -3569 9620 -3505
rect 9684 -3569 9700 -3505
rect 9764 -3569 9765 -3505
rect 9539 -3587 9765 -3569
rect 9539 -3651 9540 -3587
rect 9604 -3651 9620 -3587
rect 9684 -3651 9700 -3587
rect 9764 -3651 9765 -3587
rect 9539 -3669 9765 -3651
rect 9539 -3733 9540 -3669
rect 9604 -3733 9620 -3669
rect 9684 -3733 9700 -3669
rect 9764 -3733 9765 -3669
rect 9539 -3734 9765 -3733
rect 16543 -2936 16769 -2935
rect 16543 -3320 16544 -2936
rect 16768 -3320 16769 -2936
rect 16543 -3337 16769 -3320
rect 16543 -3401 16544 -3337
rect 16608 -3401 16624 -3337
rect 16688 -3401 16704 -3337
rect 16768 -3401 16769 -3337
rect 16543 -3418 16769 -3401
rect 16543 -3482 16544 -3418
rect 16608 -3482 16624 -3418
rect 16688 -3482 16704 -3418
rect 16768 -3482 16769 -3418
rect 16543 -3499 16769 -3482
rect 16543 -3563 16544 -3499
rect 16608 -3563 16624 -3499
rect 16688 -3563 16704 -3499
rect 16768 -3563 16769 -3499
rect 16543 -3580 16769 -3563
rect 16543 -3644 16544 -3580
rect 16608 -3644 16624 -3580
rect 16688 -3644 16704 -3580
rect 16768 -3644 16769 -3580
rect 16543 -3661 16769 -3644
rect 16543 -3725 16544 -3661
rect 16608 -3725 16624 -3661
rect 16688 -3725 16704 -3661
rect 16768 -3725 16769 -3661
rect 6490 -3806 6492 -3742
rect 6556 -3806 6594 -3742
rect 6658 -3806 6696 -3742
rect 6760 -3806 6798 -3742
rect 6862 -3806 6864 -3742
rect 6490 -3807 6864 -3806
rect 16543 -3742 16769 -3725
rect 16543 -3806 16544 -3742
rect 16608 -3806 16624 -3742
rect 16688 -3806 16704 -3742
rect 16768 -3806 16769 -3742
rect 16543 -3807 16769 -3806
use sky130_fd_io__gpio_ovtv2_hotswap_guardrings  sky130_fd_io__gpio_ovtv2_hotswap_guardrings_0
timestamp 1707688321
transform 1 0 -2942 0 1 -3349
box 0 0 26980 8664
use sky130_fd_io__tk_em1o_cdns_5595914180840  sky130_fd_io__tk_em1o_cdns_5595914180840_0
timestamp 1707688321
transform -1 0 6764 0 1 1406
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_5595914180843  sky130_fd_io__tk_em2o_cdns_5595914180843_0
timestamp 1707688321
transform -1 0 20006 0 -1 240
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_5595914180843  sky130_fd_io__tk_em2o_cdns_5595914180843_1
timestamp 1707688321
transform -1 0 20006 0 -1 1452
box 0 0 1 1
use sky130_fd_io__tk_em2o_cdns_5595914180843  sky130_fd_io__tk_em2o_cdns_5595914180843_2
timestamp 1707688321
transform 1 0 -2 0 -1 241
box 0 0 1 1
use sky130_fd_io__tk_em2s_cdns_5595914180841  sky130_fd_io__tk_em2s_cdns_5595914180841_0
timestamp 1707688321
transform 0 -1 19662 1 0 1142
box 0 0 1 1
use sky130_fd_io__tk_em2s_cdns_5595914180841  sky130_fd_io__tk_em2s_cdns_5595914180841_1
timestamp 1707688321
transform 0 -1 19662 1 0 -86
box 0 0 1 1
use sky130_fd_io__tk_em2s_cdns_5595914180841  sky130_fd_io__tk_em2s_cdns_5595914180841_2
timestamp 1707688321
transform 0 1 9897 1 0 -126
box 0 0 1 1
use sky130_fd_io__tk_em2s_cdns_5595914180842  sky130_fd_io__tk_em2s_cdns_5595914180842_0
timestamp 1707688321
transform 1 0 -53 0 -1 121
box 0 0 1 1
use sky130_fd_pr__nfet_01v8__example_5595914180834  sky130_fd_pr__nfet_01v8__example_5595914180834_0
timestamp 1707688321
transform 1 0 -1552 0 1 11787
box -1 0 257 1
use sky130_fd_pr__nfet_01v8__example_5595914180834  sky130_fd_pr__nfet_01v8__example_5595914180834_1
timestamp 1707688321
transform 1 0 -1552 0 -1 11655
box -1 0 257 1
use sky130_fd_pr__nfet_01v8__example_5595914180834  sky130_fd_pr__nfet_01v8__example_5595914180834_2
timestamp 1707688321
transform 1 0 -1552 0 1 10323
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_5595914180837  sky130_fd_pr__pfet_01v8__example_5595914180837_0
timestamp 1707688321
transform 1 0 -1596 0 -1 2025
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_5595914180837  sky130_fd_pr__pfet_01v8__example_5595914180837_1
timestamp 1707688321
transform 1 0 -1153 0 -1 2831
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_5595914180837  sky130_fd_pr__pfet_01v8__example_5595914180837_2
timestamp 1707688321
transform 1 0 -1596 0 -1 2831
box -1 0 257 1
use sky130_fd_pr__res_generic_po__example_5595914180838  sky130_fd_pr__res_generic_po__example_5595914180838_0
timestamp 1707688321
transform -1 0 21839 0 1 5424
box 15 17 2025 18
use sky130_fd_pr__res_generic_po__example_5595914180838  sky130_fd_pr__res_generic_po__example_5595914180838_1
timestamp 1707688321
transform -1 0 21796 0 1 6051
box 15 17 2025 18
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_0
timestamp 1707688321
transform 1 0 19638 0 1 6068
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_1
timestamp 1707688321
transform -1 0 21914 0 1 6068
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_2
timestamp 1707688321
transform -1 0 21923 0 1 5868
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_3
timestamp 1707688321
transform 1 0 19647 0 1 5868
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_4
timestamp 1707688321
transform -1 0 21914 0 1 5642
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_5
timestamp 1707688321
transform 1 0 19638 0 1 5642
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_6
timestamp 1707688321
transform -1 0 21957 0 1 5441
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_7
timestamp 1707688321
transform 1 0 19681 0 1 5441
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_0
timestamp 1707688321
transform -1 0 9957 0 1 902
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_1
timestamp 1707688321
transform -1 0 16441 0 1 78
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_2
timestamp 1707688321
transform -1 0 16441 0 -1 624
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_3
timestamp 1707688321
transform -1 0 13200 0 1 902
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_4
timestamp 1707688321
transform 1 0 19606 0 1 902
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_5
timestamp 1707688321
transform -1 0 232 0 -1 1448
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_6
timestamp 1707688321
transform -1 0 3473 0 -1 1448
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_7
timestamp 1707688321
transform -1 0 9957 0 -1 1448
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_8
timestamp 1707688321
transform -1 0 6715 0 1 902
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_9
timestamp 1707688321
transform -1 0 232 0 1 902
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_10
timestamp 1707688321
transform 1 0 19606 0 -1 1036
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_11
timestamp 1707688321
transform 1 0 19606 0 1 1314
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_12
timestamp 1707688321
transform -1 0 3473 0 -1 1036
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_13
timestamp 1707688321
transform -1 0 232 0 -1 624
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_14
timestamp 1707688321
transform -1 0 13199 0 -1 624
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_15
timestamp 1707688321
transform -1 0 9957 0 -1 624
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_16
timestamp 1707688321
transform -1 0 6715 0 -1 624
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_17
timestamp 1707688321
transform -1 0 3473 0 -1 624
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_18
timestamp 1707688321
transform -1 0 232 0 1 78
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_19
timestamp 1707688321
transform -1 0 3473 0 1 78
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_20
timestamp 1707688321
transform -1 0 9957 0 1 78
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_21
timestamp 1707688321
transform 1 0 19606 0 1 78
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_22
timestamp 1707688321
transform 1 0 19606 0 1 490
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_23
timestamp 1707688321
transform -1 0 16442 0 -1 1448
box 0 0 1 1
<< labels >>
flabel locali s -1538 2073 -1477 2121 3 FreeSans 200 0 0 0 PGHS_H[4]
port 1 nsew
flabel locali s -1028 2879 -978 2927 3 FreeSans 200 0 0 0 PGHS_H[3]
port 2 nsew
flabel locali s -1529 2879 -1484 2927 3 FreeSans 200 0 0 0 PGHS_H[2]
port 3 nsew
flabel metal3 s 18064 258 18628 471 3 FreeSans 200 0 0 0 PAD
port 4 nsew
flabel metal2 s -1084 2980 -1032 3030 3 FreeSans 200 0 0 0 PU_H_N[3]
port 5 nsew
flabel metal2 s -1360 2878 -1308 2933 3 FreeSans 200 0 0 0 PU_H_N[2]
port 6 nsew
flabel metal2 s -1636 1954 -1585 2032 3 FreeSans 200 0 0 0 PU_CSD_H
port 7 nsew
flabel metal1 s -877 7562 -698 7726 3 FreeSans 200 0 0 0 VDDIO
port 8 nsew
flabel metal1 s 19858 4225 19950 4344 3 FreeSans 520 90 0 0 VPB_DRVR
port 9 nsew
flabel metal1 s 6569 1538 6764 1632 3 FreeSans 200 0 0 0 VDDIO_AMX
port 10 nsew
flabel metal1 s -544 749 -434 875 3 FreeSans 200 0 0 0 PUG_H[4]
port 11 nsew
flabel metal1 s -506 2356 -456 2406 3 FreeSans 200 0 0 0 PUG_H[3]
port 12 nsew
flabel metal1 s -495 2523 -447 2573 3 FreeSans 200 0 0 0 PUG_H[2]
port 13 nsew
flabel metal1 s 21420 5415 21539 5532 3 FreeSans 200 0 0 0 TIE_HI_ESD
port 14 nsew
flabel metal1 s -1152 10966 -1069 11093 3 FreeSans 200 0 0 0 VSSIO
port 15 nsew
flabel metal1 s -2190 -2789 -2049 -2651 3 FreeSans 200 0 0 0 VSSD
port 16 nsew
flabel metal1 s -2635 -3184 -2456 -3020 3 FreeSans 200 0 0 0 VDDIO
port 8 nsew
flabel metal1 s -1525 11996 -1479 12047 3 FreeSans 200 0 0 0 NGHS_H[4]
port 17 nsew
flabel metal1 s -1524 11260 -1479 11301 3 FreeSans 200 0 0 0 NGHS_H[3]
port 18 nsew
flabel metal1 s -1525 10850 -1479 10892 3 FreeSans 200 0 0 0 NGHS_H[2]
port 19 nsew
flabel comment s 20827 6110 20827 6110 0 FreeSans 440 180 0 0 LEAKER
flabel comment s -105 -195 -105 -195 0 FreeSans 200 90 0 0 TIE_HI_VPBDRVR
flabel comment s -602 1435 -602 1435 0 FreeSans 200 90 0 0 <4>
flabel comment s 20026 1516 20026 1516 0 FreeSans 200 180 0 0 <3>
flabel comment s 20035 -183 20035 -183 0 FreeSans 200 90 0 0 TIE_HI_VPBDRVR
flabel comment s 20870 5483 20870 5483 0 FreeSans 440 180 0 0 LEAKER
flabel comment s -198 1470 -198 1470 0 FreeSans 200 90 0 0 <2>
flabel comment s 22098 18 22098 18 0 FreeSans 400 0 0 0 TIE_HI_VPBDRVR
<< properties >>
string GDS_END 75999870
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 74818954
<< end >>
