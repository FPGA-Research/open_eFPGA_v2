magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -68 -144 35034 84
<< ndiff >>
rect -42 46 0 58
rect -42 12 -34 46
rect -42 0 0 12
rect -42 -72 0 -60
rect -42 -106 -34 -72
rect -42 -118 0 -106
<< ndiffc >>
rect -34 12 0 46
rect -34 -106 0 -72
<< ndiffres >>
rect 0 0 35008 58
rect 34950 -60 35008 0
rect 0 -118 35008 -60
<< locali >>
rect -34 46 0 62
rect -34 -4 0 12
rect -34 -72 0 -56
rect -34 -122 0 -106
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_0
timestamp 1707688321
transform 1 0 -42 0 1 -118
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_1
timestamp 1707688321
transform 1 0 -42 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 24809284
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 24808480
<< end >>
