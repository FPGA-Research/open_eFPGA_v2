magic
tech sky130B
timestamp 1707688321
<< viali >>
rect 0 0 161 89
<< metal1 >>
rect -6 89 167 92
rect -6 0 0 89
rect 161 0 167 89
rect -6 -3 167 0
<< properties >>
string GDS_END 95663146
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 95662054
<< end >>
