magic
tech sky130A
timestamp 1707688321
<< viali >>
rect 0 0 53 377
<< metal1 >>
rect -6 377 59 380
rect -6 0 0 377
rect 53 0 59 377
rect -6 -3 59 0
<< properties >>
string GDS_END 94936628
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 94935088
<< end >>
