magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -38 287 2706 582
rect -38 261 977 287
rect 1440 261 2706 287
<< pwell >>
rect 1034 157 1427 229
rect 1680 157 1864 201
rect 2449 157 2639 203
rect 1 93 2639 157
rect 1 21 993 93
rect 1287 21 2639 93
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 351 47 381 131
rect 423 47 453 131
rect 611 47 641 131
rect 699 47 729 131
rect 801 47 831 131
rect 885 47 915 131
rect 1112 119 1142 203
rect 1196 119 1226 203
rect 1268 119 1298 203
rect 1443 47 1473 119
rect 1531 47 1561 119
rect 1637 47 1667 131
rect 1756 47 1786 175
rect 1944 47 1974 131
rect 2041 47 2071 119
rect 2147 47 2177 119
rect 2242 47 2272 131
rect 2430 47 2460 131
rect 2527 47 2557 177
<< scpmoshvt >>
rect 79 363 109 491
rect 163 363 193 491
rect 351 369 381 497
rect 423 369 453 497
rect 611 369 641 497
rect 699 369 729 497
rect 801 369 831 497
rect 893 369 923 497
rect 1092 369 1122 497
rect 1201 369 1231 497
rect 1297 369 1327 497
rect 1416 413 1446 497
rect 1507 413 1537 497
rect 1610 413 1640 497
rect 1742 347 1772 497
rect 1930 413 1960 497
rect 2021 413 2051 497
rect 2105 413 2135 497
rect 2219 413 2249 497
rect 2430 369 2460 497
rect 2527 297 2557 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 299 100 351 131
rect 299 66 307 100
rect 341 66 351 100
rect 299 47 351 66
rect 381 47 423 131
rect 453 93 505 131
rect 453 59 463 93
rect 497 59 505 93
rect 453 47 505 59
rect 559 119 611 131
rect 559 85 567 119
rect 601 85 611 119
rect 559 47 611 85
rect 641 106 699 131
rect 641 72 653 106
rect 687 72 699 106
rect 641 47 699 72
rect 729 47 801 131
rect 831 106 885 131
rect 831 72 841 106
rect 875 72 885 106
rect 831 47 885 72
rect 915 106 967 131
rect 915 72 925 106
rect 959 72 967 106
rect 915 47 967 72
rect 1060 167 1112 203
rect 1060 133 1068 167
rect 1102 133 1112 167
rect 1060 119 1112 133
rect 1142 165 1196 203
rect 1142 131 1152 165
rect 1186 131 1196 165
rect 1142 119 1196 131
rect 1226 119 1268 203
rect 1298 180 1401 203
rect 1298 146 1310 180
rect 1344 146 1401 180
rect 1298 119 1401 146
rect 1706 131 1756 175
rect 1587 119 1637 131
rect 1313 99 1443 119
rect 1313 65 1377 99
rect 1411 65 1443 99
rect 1313 47 1443 65
rect 1473 99 1531 119
rect 1473 65 1483 99
rect 1517 65 1531 99
rect 1473 47 1531 65
rect 1561 47 1637 119
rect 1667 101 1756 131
rect 1667 67 1678 101
rect 1712 67 1756 101
rect 1667 47 1756 67
rect 1786 163 1838 175
rect 1786 129 1796 163
rect 1830 129 1838 163
rect 1786 95 1838 129
rect 1786 61 1796 95
rect 1830 61 1838 95
rect 1786 47 1838 61
rect 1892 107 1944 131
rect 1892 73 1900 107
rect 1934 73 1944 107
rect 1892 47 1944 73
rect 1974 119 2024 131
rect 2475 164 2527 177
rect 2475 131 2483 164
rect 2192 119 2242 131
rect 1974 47 2041 119
rect 2071 104 2147 119
rect 2071 70 2084 104
rect 2118 70 2147 104
rect 2071 47 2147 70
rect 2177 47 2242 119
rect 2272 107 2324 131
rect 2272 73 2282 107
rect 2316 73 2324 107
rect 2272 47 2324 73
rect 2378 94 2430 131
rect 2378 60 2386 94
rect 2420 60 2430 94
rect 2378 47 2430 60
rect 2460 130 2483 131
rect 2517 130 2527 164
rect 2460 96 2527 130
rect 2460 62 2483 96
rect 2517 62 2527 96
rect 2460 47 2527 62
rect 2557 164 2613 177
rect 2557 130 2569 164
rect 2603 130 2613 164
rect 2557 96 2613 130
rect 2557 62 2569 96
rect 2603 62 2613 96
rect 2557 47 2613 62
<< pdiff >>
rect 27 477 79 491
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 363 79 375
rect 109 461 163 491
rect 109 427 119 461
rect 153 427 163 461
rect 109 363 163 427
rect 193 477 245 491
rect 193 443 203 477
rect 237 443 245 477
rect 193 409 245 443
rect 193 375 203 409
rect 237 375 245 409
rect 193 363 245 375
rect 299 485 351 497
rect 299 451 307 485
rect 341 451 351 485
rect 299 415 351 451
rect 299 381 307 415
rect 341 381 351 415
rect 299 369 351 381
rect 381 369 423 497
rect 453 485 505 497
rect 453 451 463 485
rect 497 451 505 485
rect 453 417 505 451
rect 453 383 463 417
rect 497 383 505 417
rect 453 369 505 383
rect 559 485 611 497
rect 559 451 567 485
rect 601 451 611 485
rect 559 415 611 451
rect 559 381 567 415
rect 601 381 611 415
rect 559 369 611 381
rect 641 485 699 497
rect 641 451 653 485
rect 687 451 699 485
rect 641 415 699 451
rect 641 381 653 415
rect 687 381 699 415
rect 641 369 699 381
rect 729 369 801 497
rect 831 485 893 497
rect 831 451 841 485
rect 875 451 893 485
rect 831 417 893 451
rect 831 383 841 417
rect 875 383 893 417
rect 831 369 893 383
rect 923 485 985 497
rect 923 451 943 485
rect 977 451 985 485
rect 923 417 985 451
rect 923 383 943 417
rect 977 383 985 417
rect 923 369 985 383
rect 1039 485 1092 497
rect 1039 451 1047 485
rect 1081 451 1092 485
rect 1039 417 1092 451
rect 1039 383 1047 417
rect 1081 383 1092 417
rect 1039 369 1092 383
rect 1122 485 1201 497
rect 1122 451 1144 485
rect 1178 451 1201 485
rect 1122 369 1201 451
rect 1231 369 1297 497
rect 1327 485 1416 497
rect 1327 451 1351 485
rect 1385 451 1416 485
rect 1327 417 1416 451
rect 1327 383 1351 417
rect 1385 413 1416 417
rect 1446 472 1507 497
rect 1446 438 1459 472
rect 1493 438 1507 472
rect 1446 413 1507 438
rect 1537 413 1610 497
rect 1640 485 1742 497
rect 1640 451 1692 485
rect 1726 451 1742 485
rect 1640 417 1742 451
rect 1640 413 1692 417
rect 1385 383 1401 413
rect 1327 369 1401 383
rect 1655 383 1692 413
rect 1726 383 1742 417
rect 1655 347 1742 383
rect 1772 485 1824 497
rect 1772 451 1782 485
rect 1816 451 1824 485
rect 1772 393 1824 451
rect 1878 472 1930 497
rect 1878 438 1886 472
rect 1920 438 1930 472
rect 1878 413 1930 438
rect 1960 413 2021 497
rect 2051 469 2105 497
rect 2051 435 2061 469
rect 2095 435 2105 469
rect 2051 413 2105 435
rect 2135 413 2219 497
rect 2249 477 2302 497
rect 2249 443 2260 477
rect 2294 443 2302 477
rect 2249 413 2302 443
rect 2376 485 2430 497
rect 2376 451 2384 485
rect 2418 451 2430 485
rect 2376 415 2430 451
rect 1772 359 1782 393
rect 1816 359 1824 393
rect 1772 347 1824 359
rect 2376 381 2384 415
rect 2418 381 2430 415
rect 2376 369 2430 381
rect 2460 479 2527 497
rect 2460 445 2483 479
rect 2517 445 2527 479
rect 2460 411 2527 445
rect 2460 377 2483 411
rect 2517 377 2527 411
rect 2460 369 2527 377
rect 2475 343 2527 369
rect 2475 309 2483 343
rect 2517 309 2527 343
rect 2475 297 2527 309
rect 2557 479 2613 497
rect 2557 445 2569 479
rect 2603 445 2613 479
rect 2557 411 2613 445
rect 2557 377 2569 411
rect 2603 377 2613 411
rect 2557 343 2613 377
rect 2557 309 2569 343
rect 2603 309 2613 343
rect 2557 297 2613 309
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 307 66 341 100
rect 463 59 497 93
rect 567 85 601 119
rect 653 72 687 106
rect 841 72 875 106
rect 925 72 959 106
rect 1068 133 1102 167
rect 1152 131 1186 165
rect 1310 146 1344 180
rect 1377 65 1411 99
rect 1483 65 1517 99
rect 1678 67 1712 101
rect 1796 129 1830 163
rect 1796 61 1830 95
rect 1900 73 1934 107
rect 2084 70 2118 104
rect 2282 73 2316 107
rect 2386 60 2420 94
rect 2483 130 2517 164
rect 2483 62 2517 96
rect 2569 130 2603 164
rect 2569 62 2603 96
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 427 153 461
rect 203 443 237 477
rect 203 375 237 409
rect 307 451 341 485
rect 307 381 341 415
rect 463 451 497 485
rect 463 383 497 417
rect 567 451 601 485
rect 567 381 601 415
rect 653 451 687 485
rect 653 381 687 415
rect 841 451 875 485
rect 841 383 875 417
rect 943 451 977 485
rect 943 383 977 417
rect 1047 451 1081 485
rect 1047 383 1081 417
rect 1144 451 1178 485
rect 1351 451 1385 485
rect 1351 383 1385 417
rect 1459 438 1493 472
rect 1692 451 1726 485
rect 1692 383 1726 417
rect 1782 451 1816 485
rect 1886 438 1920 472
rect 2061 435 2095 469
rect 2260 443 2294 477
rect 2384 451 2418 485
rect 1782 359 1816 393
rect 2384 381 2418 415
rect 2483 445 2517 479
rect 2483 377 2517 411
rect 2483 309 2517 343
rect 2569 445 2603 479
rect 2569 377 2603 411
rect 2569 309 2603 343
<< poly >>
rect 79 491 109 517
rect 163 491 193 517
rect 351 497 381 523
rect 423 497 453 523
rect 611 497 641 523
rect 699 497 729 523
rect 801 497 831 523
rect 893 497 923 523
rect 1092 497 1122 523
rect 1201 497 1231 523
rect 1297 497 1327 523
rect 1416 497 1446 523
rect 1507 497 1537 523
rect 1610 497 1640 523
rect 1742 497 1772 523
rect 1930 497 1960 523
rect 2021 497 2051 523
rect 2105 497 2135 523
rect 2219 497 2249 523
rect 2430 497 2460 523
rect 2527 497 2557 523
rect 79 348 109 363
rect 47 318 109 348
rect 47 265 77 318
rect 163 274 193 363
rect 351 330 381 369
rect 423 354 453 369
rect 423 343 549 354
rect 23 249 77 265
rect 23 215 33 249
rect 67 215 77 249
rect 119 264 193 274
rect 119 230 135 264
rect 169 230 193 264
rect 119 220 193 230
rect 23 199 77 215
rect 47 176 77 199
rect 47 146 109 176
rect 79 131 109 146
rect 163 131 193 220
rect 323 314 383 330
rect 425 324 549 343
rect 323 280 339 314
rect 373 280 383 314
rect 323 246 383 280
rect 483 321 549 324
rect 483 287 499 321
rect 533 287 549 321
rect 483 277 549 287
rect 611 322 641 369
rect 699 322 729 369
rect 801 330 831 369
rect 611 292 729 322
rect 791 314 845 330
rect 323 212 339 246
rect 373 212 383 246
rect 323 196 383 212
rect 425 219 491 235
rect 351 131 381 196
rect 425 185 441 219
rect 475 200 491 219
rect 611 200 641 292
rect 791 280 801 314
rect 835 280 845 314
rect 893 315 923 369
rect 1092 315 1122 369
rect 1201 337 1231 369
rect 1297 337 1327 369
rect 893 305 1122 315
rect 893 285 1007 305
rect 791 264 845 280
rect 991 271 1007 285
rect 1041 271 1122 305
rect 1177 321 1231 337
rect 1177 287 1187 321
rect 1221 287 1231 321
rect 1177 271 1231 287
rect 1273 321 1327 337
rect 1273 287 1283 321
rect 1317 287 1327 321
rect 1416 297 1446 413
rect 1507 381 1537 413
rect 1507 365 1568 381
rect 1507 331 1524 365
rect 1558 331 1568 365
rect 1507 315 1568 331
rect 1273 271 1327 287
rect 1403 287 1469 297
rect 475 185 641 200
rect 425 176 641 185
rect 423 170 641 176
rect 423 162 491 170
rect 423 131 453 162
rect 611 131 641 170
rect 683 219 737 235
rect 683 185 693 219
rect 727 185 737 219
rect 683 169 737 185
rect 699 131 729 169
rect 801 131 831 264
rect 991 261 1122 271
rect 1092 247 1122 261
rect 1092 218 1142 247
rect 1112 203 1142 218
rect 1196 203 1226 271
rect 1403 253 1419 287
rect 1453 273 1469 287
rect 1453 253 1561 273
rect 1403 243 1561 253
rect 1268 203 1298 229
rect 885 153 1029 183
rect 885 131 915 153
rect 999 101 1029 153
rect 1423 191 1489 201
rect 1423 157 1439 191
rect 1473 157 1489 191
rect 1423 147 1489 157
rect 1443 119 1473 147
rect 1531 119 1561 243
rect 1610 213 1640 413
rect 1742 309 1772 347
rect 1682 299 1772 309
rect 1682 265 1698 299
rect 1732 265 1772 299
rect 1930 275 1960 413
rect 2021 315 2051 413
rect 2105 375 2135 413
rect 2219 381 2249 413
rect 2104 365 2170 375
rect 2104 331 2120 365
rect 2154 331 2170 365
rect 2104 321 2170 331
rect 2219 365 2300 381
rect 2219 331 2256 365
rect 2290 331 2300 365
rect 2219 315 2300 331
rect 1682 255 1772 265
rect 1742 220 1772 255
rect 1905 259 1960 275
rect 1905 225 1915 259
rect 1949 225 1960 259
rect 2008 299 2062 315
rect 2008 265 2018 299
rect 2052 279 2062 299
rect 2052 265 2177 279
rect 2008 249 2177 265
rect 1610 203 1684 213
rect 1610 169 1634 203
rect 1668 169 1684 203
rect 1742 190 1786 220
rect 1756 175 1786 190
rect 1905 209 1960 225
rect 1905 179 1974 209
rect 1610 159 1684 169
rect 1637 131 1667 159
rect 999 85 1053 101
rect 999 51 1009 85
rect 1043 51 1053 85
rect 79 21 109 47
rect 163 21 193 47
rect 351 21 381 47
rect 423 21 453 47
rect 611 21 641 47
rect 699 21 729 47
rect 801 21 831 47
rect 885 21 915 47
rect 999 35 1053 51
rect 1112 51 1142 119
rect 1196 93 1226 119
rect 1268 51 1298 119
rect 1112 21 1298 51
rect 1944 131 1974 179
rect 2041 191 2105 207
rect 2041 157 2061 191
rect 2095 157 2105 191
rect 2041 141 2105 157
rect 2041 119 2071 141
rect 2147 119 2177 249
rect 2242 131 2272 315
rect 2430 265 2460 369
rect 2527 265 2557 297
rect 2318 249 2557 265
rect 2318 215 2328 249
rect 2362 215 2557 249
rect 2318 199 2557 215
rect 2430 131 2460 199
rect 2527 177 2557 199
rect 1443 21 1473 47
rect 1531 21 1561 47
rect 1637 21 1667 47
rect 1756 21 1786 47
rect 1944 21 1974 47
rect 2041 21 2071 47
rect 2147 21 2177 47
rect 2242 21 2272 47
rect 2430 21 2460 47
rect 2527 21 2557 47
<< polycont >>
rect 33 215 67 249
rect 135 230 169 264
rect 339 280 373 314
rect 499 287 533 321
rect 339 212 373 246
rect 441 185 475 219
rect 801 280 835 314
rect 1007 271 1041 305
rect 1187 287 1221 321
rect 1283 287 1317 321
rect 1524 331 1558 365
rect 693 185 727 219
rect 1419 253 1453 287
rect 1439 157 1473 191
rect 1698 265 1732 299
rect 2120 331 2154 365
rect 2256 331 2290 365
rect 1915 225 1949 259
rect 2018 265 2052 299
rect 1634 169 1668 203
rect 1009 51 1043 85
rect 2061 157 2095 191
rect 2328 215 2362 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2668 561
rect 35 477 69 493
rect 35 409 69 443
rect 103 461 169 527
rect 103 427 119 461
rect 153 427 169 461
rect 203 477 237 493
rect 203 409 237 443
rect 69 391 169 393
rect 69 375 127 391
rect 35 359 127 375
rect 123 357 127 359
rect 161 357 169 391
rect 19 249 89 325
rect 19 215 33 249
rect 67 215 89 249
rect 19 195 89 215
rect 123 264 169 357
rect 123 230 135 264
rect 123 161 169 230
rect 35 127 169 161
rect 203 323 237 375
rect 35 119 69 127
rect 203 119 237 289
rect 35 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 203 69 237 85
rect 271 485 357 493
rect 271 451 307 485
rect 341 451 357 485
rect 271 415 357 451
rect 271 381 307 415
rect 341 381 357 415
rect 271 378 357 381
rect 447 485 513 527
rect 653 485 692 527
rect 447 451 463 485
rect 497 451 513 485
rect 447 417 513 451
rect 447 383 463 417
rect 497 383 513 417
rect 447 378 513 383
rect 551 451 567 485
rect 601 451 617 485
rect 551 415 617 451
rect 551 381 567 415
rect 601 381 617 415
rect 271 119 305 378
rect 551 344 617 381
rect 687 451 692 485
rect 653 415 692 451
rect 687 381 692 415
rect 653 365 692 381
rect 825 485 891 493
rect 825 451 841 485
rect 875 451 891 485
rect 825 417 891 451
rect 927 485 993 493
rect 927 451 943 485
rect 977 451 993 485
rect 927 442 993 451
rect 825 383 841 417
rect 875 404 891 417
rect 937 417 993 442
rect 875 383 903 404
rect 825 364 903 383
rect 339 314 383 344
rect 373 280 383 314
rect 339 246 383 280
rect 499 321 617 344
rect 533 287 617 321
rect 373 212 383 246
rect 339 153 383 212
rect 422 237 465 274
rect 499 271 617 287
rect 422 219 513 237
rect 422 185 441 219
rect 475 185 513 219
rect 422 153 513 185
rect 556 235 617 271
rect 761 314 835 330
rect 761 280 801 314
rect 761 264 835 280
rect 556 219 727 235
rect 556 185 693 219
rect 556 169 727 185
rect 761 187 795 264
rect 869 230 903 364
rect 556 119 601 169
rect 761 137 795 153
rect 829 196 903 230
rect 937 383 943 417
rect 977 383 993 417
rect 937 357 993 383
rect 1031 485 1099 493
rect 1031 451 1047 485
rect 1081 451 1099 485
rect 1031 417 1099 451
rect 1133 485 1202 527
rect 1133 451 1144 485
rect 1178 451 1202 485
rect 1133 435 1202 451
rect 1335 485 1401 493
rect 1335 451 1351 485
rect 1385 451 1401 485
rect 1685 485 1732 527
rect 1335 430 1401 451
rect 1443 472 1651 475
rect 1443 438 1459 472
rect 1493 438 1651 472
rect 1443 435 1651 438
rect 1031 383 1047 417
rect 1081 401 1099 417
rect 1351 417 1401 430
rect 1081 383 1317 401
rect 1031 367 1317 383
rect 305 100 357 103
rect 305 85 307 100
rect 103 17 169 59
rect 271 66 307 85
rect 341 66 357 100
rect 271 51 357 66
rect 447 93 513 103
rect 447 59 463 93
rect 497 59 513 93
rect 447 17 513 59
rect 556 85 567 119
rect 556 51 601 85
rect 637 106 703 122
rect 637 72 653 106
rect 687 72 703 106
rect 637 17 703 72
rect 829 119 883 196
rect 937 165 971 357
rect 1005 305 1050 323
rect 1005 271 1007 305
rect 1041 271 1050 305
rect 1005 221 1050 271
rect 1084 187 1118 367
rect 1152 321 1243 333
rect 1152 287 1187 321
rect 1221 287 1243 321
rect 1152 221 1243 287
rect 1277 321 1317 367
rect 1277 287 1283 321
rect 1277 271 1317 287
rect 1385 383 1401 417
rect 1351 373 1401 383
rect 1490 391 1583 401
rect 1351 237 1385 373
rect 1490 357 1502 391
rect 1536 365 1583 391
rect 829 85 837 119
rect 871 106 883 119
rect 829 72 841 85
rect 875 72 883 106
rect 829 51 883 72
rect 919 129 971 165
rect 1052 167 1118 187
rect 1052 133 1068 167
rect 1102 133 1118 167
rect 919 119 959 129
rect 919 85 923 119
rect 957 106 959 119
rect 1052 103 1118 133
rect 919 72 925 85
rect 919 51 959 72
rect 993 85 1118 103
rect 993 51 1009 85
rect 1043 51 1118 85
rect 1152 165 1202 181
rect 1186 131 1202 165
rect 1152 17 1202 131
rect 1303 180 1385 237
rect 1419 323 1456 344
rect 1419 289 1420 323
rect 1454 289 1456 323
rect 1419 287 1456 289
rect 1453 253 1456 287
rect 1419 225 1456 253
rect 1490 191 1524 357
rect 1558 331 1583 365
rect 1617 315 1651 435
rect 1685 451 1692 485
rect 1726 451 1732 485
rect 1685 417 1732 451
rect 1685 383 1692 417
rect 1726 383 1732 417
rect 1685 367 1732 383
rect 1766 485 1832 493
rect 1766 451 1782 485
rect 1816 451 1832 485
rect 1766 393 1832 451
rect 1874 472 1932 527
rect 1874 438 1886 472
rect 1920 438 1932 472
rect 2256 477 2308 527
rect 1874 421 1932 438
rect 2045 469 2222 471
rect 2045 435 2061 469
rect 2095 435 2222 469
rect 2045 433 2222 435
rect 1766 359 1782 393
rect 1816 359 1832 393
rect 1617 299 1732 315
rect 1617 297 1698 299
rect 1303 146 1310 180
rect 1344 146 1385 180
rect 1423 157 1439 191
rect 1473 157 1524 191
rect 1423 147 1524 157
rect 1562 265 1698 297
rect 1562 263 1732 265
rect 1303 119 1385 146
rect 1303 85 1306 119
rect 1340 113 1385 119
rect 1562 113 1596 263
rect 1698 249 1732 263
rect 1766 275 1832 359
rect 2018 391 2056 393
rect 2018 357 2020 391
rect 2054 357 2056 391
rect 2018 299 2056 357
rect 1766 259 1949 275
rect 1766 225 1915 259
rect 2052 265 2056 299
rect 2018 249 2056 265
rect 2090 365 2154 399
rect 2090 331 2120 365
rect 2090 323 2154 331
rect 2090 289 2104 323
rect 2138 289 2154 323
rect 1634 213 1674 219
rect 1766 213 1949 225
rect 1634 209 1949 213
rect 1634 203 1847 209
rect 2090 207 2154 289
rect 1668 169 1847 203
rect 1634 163 1847 169
rect 1634 153 1796 163
rect 1340 99 1427 113
rect 1340 85 1377 99
rect 1303 65 1377 85
rect 1411 65 1427 99
rect 1303 51 1427 65
rect 1461 99 1596 113
rect 1766 129 1796 153
rect 1830 129 1847 163
rect 2061 191 2154 207
rect 2095 157 2154 191
rect 2061 141 2154 157
rect 2188 265 2222 433
rect 2256 443 2260 477
rect 2294 443 2308 477
rect 2256 427 2308 443
rect 2368 485 2436 493
rect 2368 451 2384 485
rect 2418 451 2436 485
rect 2368 415 2436 451
rect 2368 381 2384 415
rect 2418 381 2436 415
rect 2256 365 2436 381
rect 2290 331 2436 365
rect 2256 306 2436 331
rect 2188 249 2362 265
rect 2188 215 2328 249
rect 2188 199 2362 215
rect 1461 65 1483 99
rect 1517 65 1596 99
rect 1461 51 1596 65
rect 1649 101 1728 112
rect 1649 67 1678 101
rect 1712 67 1728 101
rect 1649 17 1728 67
rect 1766 95 1847 129
rect 1766 61 1796 95
rect 1830 61 1847 95
rect 1766 51 1847 61
rect 1893 107 1948 123
rect 2188 107 2222 199
rect 2398 187 2436 306
rect 2470 479 2519 527
rect 2470 445 2483 479
rect 2517 445 2519 479
rect 2470 411 2519 445
rect 2470 377 2483 411
rect 2517 377 2519 411
rect 2470 343 2519 377
rect 2470 309 2483 343
rect 2517 309 2519 343
rect 2470 293 2519 309
rect 2553 479 2619 484
rect 2553 445 2569 479
rect 2603 445 2619 479
rect 2553 411 2619 445
rect 2553 377 2569 411
rect 2603 377 2619 411
rect 2553 343 2619 377
rect 2553 309 2569 343
rect 2603 309 2619 343
rect 2398 165 2400 187
rect 2370 153 2400 165
rect 2434 153 2436 187
rect 1893 73 1900 107
rect 1934 73 1948 107
rect 1893 17 1948 73
rect 2065 104 2222 107
rect 2065 70 2084 104
rect 2118 70 2222 104
rect 2065 66 2222 70
rect 2270 107 2333 123
rect 2270 73 2282 107
rect 2316 73 2333 107
rect 2270 17 2333 73
rect 2370 94 2436 153
rect 2370 60 2386 94
rect 2420 60 2436 94
rect 2470 164 2519 180
rect 2470 130 2483 164
rect 2517 130 2519 164
rect 2470 96 2519 130
rect 2470 62 2483 96
rect 2517 62 2519 96
rect 2470 17 2519 62
rect 2553 164 2619 309
rect 2553 130 2569 164
rect 2603 130 2619 164
rect 2553 96 2619 130
rect 2553 62 2569 96
rect 2603 62 2619 96
rect 2553 61 2619 62
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2668 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 2605 527 2639 561
rect 127 357 161 391
rect 203 289 237 323
rect 271 85 305 119
rect 761 153 795 187
rect 1502 365 1536 391
rect 1502 357 1524 365
rect 1524 357 1536 365
rect 837 106 871 119
rect 837 85 841 106
rect 841 85 871 106
rect 923 106 957 119
rect 923 85 925 106
rect 925 85 957 106
rect 1420 289 1454 323
rect 1306 85 1340 119
rect 2020 357 2054 391
rect 2104 289 2138 323
rect 2400 153 2434 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
rect 2605 -17 2639 17
<< metal1 >>
rect 0 561 2668 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2605 561
rect 2639 527 2668 561
rect 0 496 2668 527
rect 115 391 173 397
rect 115 357 127 391
rect 161 388 173 391
rect 1490 391 1548 397
rect 1490 388 1502 391
rect 161 360 1502 388
rect 161 357 173 360
rect 115 351 173 357
rect 1490 357 1502 360
rect 1536 388 1548 391
rect 2008 391 2066 397
rect 2008 388 2020 391
rect 1536 360 2020 388
rect 1536 357 1548 360
rect 1490 351 1548 357
rect 2008 357 2020 360
rect 2054 357 2066 391
rect 2008 351 2066 357
rect 191 323 249 329
rect 191 289 203 323
rect 237 320 249 323
rect 1408 323 1466 329
rect 1408 320 1420 323
rect 237 292 1420 320
rect 237 289 249 292
rect 191 283 249 289
rect 1408 289 1420 292
rect 1454 320 1466 323
rect 2092 323 2150 329
rect 2092 320 2104 323
rect 1454 292 2104 320
rect 1454 289 1466 292
rect 1408 283 1466 289
rect 2092 289 2104 292
rect 2138 289 2150 323
rect 2092 283 2150 289
rect 749 187 807 193
rect 749 153 761 187
rect 795 184 807 187
rect 2388 187 2446 193
rect 2388 184 2400 187
rect 795 156 2400 184
rect 795 153 807 156
rect 749 147 807 153
rect 2388 153 2400 156
rect 2434 153 2446 187
rect 2388 147 2446 153
rect 259 119 317 125
rect 259 85 271 119
rect 305 116 317 119
rect 825 119 883 125
rect 825 116 837 119
rect 305 85 837 116
rect 871 85 883 119
rect 259 79 883 85
rect 911 119 969 125
rect 911 85 923 119
rect 957 116 969 119
rect 1294 119 1352 125
rect 1294 116 1306 119
rect 957 85 1306 116
rect 1340 85 1352 119
rect 911 79 1352 85
rect 0 17 2668 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2605 17
rect 2639 -17 2668 17
rect 0 -48 2668 -17
<< labels >>
rlabel comment s 0 0 0 0 4 sedfxtp_1
flabel comment s 1433 304 1433 304 0 FreeSans 200 0 0 0 clkpos
flabel comment s 1520 374 1520 374 0 FreeSans 200 0 0 0 clkneg
flabel comment s 2417 174 2417 174 0 FreeSans 200 0 0 0 q1
flabel comment s 219 304 219 304 0 FreeSans 200 0 0 0 clkpos
flabel comment s 147 374 147 374 0 FreeSans 200 0 0 0 clkneg
flabel comment s 623 209 623 209 0 FreeSans 200 0 0 0 deneg
flabel comment s 939 104 939 104 0 FreeSans 200 0 0 0 db
flabel comment s 780 174 780 174 0 FreeSans 200 0 0 0 q1
flabel comment s 2120 304 2120 304 0 FreeSans 200 0 0 0 clkpos
flabel comment s 2037 374 2037 374 0 FreeSans 200 0 0 0 clkneg
flabel comment s 1343 104 1343 104 0 FreeSans 200 0 0 0 db
flabel comment s 2205 269 2205 269 0 FreeSans 200 0 0 0 S0
flabel comment s 1099 344 1099 344 0 FreeSans 200 0 0 0 sceneg
flabel comment s 1716 269 1716 269 0 FreeSans 200 0 0 0 M0
flabel comment s 1802 269 1802 269 0 FreeSans 200 0 0 0 M1
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel locali s 29 221 63 255 0 FreeSans 400 0 0 0 CLK
port 1 nsew clock input
flabel locali s 1179 221 1213 255 0 FreeSans 400 0 0 0 SCD
port 4 nsew signal input
flabel locali s 426 153 460 187 0 FreeSans 400 0 0 0 DE
port 3 nsew signal input
flabel locali s 344 221 378 255 0 FreeSans 400 0 0 0 D
port 2 nsew signal input
flabel locali s 2565 221 2599 255 0 FreeSans 400 0 0 0 Q
port 10 nsew signal output
flabel locali s 1011 289 1045 323 0 FreeSans 400 0 0 0 SCE
port 5 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
flabel pwell s 29 -17 63 17 0 FreeSans 400 0 0 0 VNB
port 7 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
rlabel metal1 s 0 -48 2668 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 2668 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2668 544
string GDS_END 512704
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 491556
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
