magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 1 21 557 203
rect 29 -17 63 21
<< locali >>
rect 103 357 173 417
rect 17 199 69 265
rect 103 161 137 357
rect 171 285 251 323
rect 171 199 205 285
rect 246 215 319 251
rect 103 127 233 161
rect 183 59 233 127
rect 281 153 319 215
rect 361 199 433 265
rect 467 203 550 265
rect 281 69 341 153
rect 393 83 433 199
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 17 451 269 493
rect 17 367 69 451
rect 219 391 269 451
rect 311 427 361 527
rect 403 391 437 493
rect 219 357 437 391
rect 403 349 437 357
rect 471 299 539 527
rect 19 17 85 93
rect 471 17 539 161
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 281 69 341 153 6 A1
port 1 nsew signal input
rlabel locali s 281 153 319 215 6 A1
port 1 nsew signal input
rlabel locali s 246 215 319 251 6 A1
port 1 nsew signal input
rlabel locali s 393 83 433 199 6 A2
port 2 nsew signal input
rlabel locali s 361 199 433 265 6 A2
port 2 nsew signal input
rlabel locali s 467 203 550 265 6 A3
port 3 nsew signal input
rlabel locali s 171 199 205 285 6 B1
port 4 nsew signal input
rlabel locali s 171 285 251 323 6 B1
port 4 nsew signal input
rlabel locali s 17 199 69 265 6 B2
port 5 nsew signal input
rlabel metal1 s 0 -48 644 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1 21 557 203 6 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 682 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 183 59 233 127 6 Y
port 10 nsew signal output
rlabel locali s 103 127 233 161 6 Y
port 10 nsew signal output
rlabel locali s 103 161 137 357 6 Y
port 10 nsew signal output
rlabel locali s 103 357 173 417 6 Y
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 644 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3473666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3467700
<< end >>
