magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -122 -66 378 666
<< mvpmos >>
rect 0 0 100 600
rect 156 0 256 600
<< mvpdiff >>
rect -50 0 0 600
rect 256 0 306 600
<< poly >>
rect 0 600 100 632
rect 0 -32 100 0
rect 156 600 256 632
rect 156 -32 256 0
<< locali >>
rect -45 -4 -11 538
rect 111 -4 145 538
rect 267 -4 301 538
use DFL1sd2_CDNS_5246887918535  DFL1sd2_CDNS_5246887918535_0
timestamp 1707688321
transform 1 0 100 0 1 0
box -36 -36 92 636
use hvDFL1sd2_CDNS_52468879185138  hvDFL1sd2_CDNS_52468879185138_0
timestamp 1707688321
transform -1 0 0 0 1 0
box -36 -36 92 636
use hvDFL1sd2_CDNS_52468879185138  hvDFL1sd2_CDNS_52468879185138_1
timestamp 1707688321
transform 1 0 256 0 1 0
box -36 -36 92 636
<< labels >>
flabel comment s -28 267 -28 267 0 FreeSans 300 0 0 0 D
flabel comment s 128 267 128 267 0 FreeSans 300 0 0 0 S
flabel comment s 284 267 284 267 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 85598764
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85597246
<< end >>
