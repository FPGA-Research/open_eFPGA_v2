magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect 0 1854 3426 1950
rect 0 1152 136 1854
rect 3290 1582 3426 1854
rect 3338 1552 3426 1582
rect 0 1122 1516 1152
<< pwell >>
rect 278 10 364 1062
rect 1214 10 1300 1062
<< mvpsubdiff >>
rect 304 1012 338 1036
rect 304 941 338 978
rect 304 870 338 907
rect 304 799 338 836
rect 304 728 338 765
rect 304 657 338 694
rect 304 586 338 623
rect 304 515 338 552
rect 304 444 338 481
rect 304 374 338 410
rect 304 304 338 340
rect 304 234 338 270
rect 304 164 338 200
rect 304 94 338 130
rect 304 36 338 60
rect 1240 1012 1274 1036
rect 1240 941 1274 978
rect 1240 870 1274 907
rect 1240 799 1274 836
rect 1240 728 1274 765
rect 1240 657 1274 694
rect 1240 586 1274 623
rect 1240 515 1274 552
rect 1240 444 1274 481
rect 1240 374 1274 410
rect 1240 304 1274 340
rect 1240 234 1274 270
rect 1240 164 1274 200
rect 1240 94 1274 130
rect 1240 36 1274 60
<< mvnsubdiff >>
rect 66 1794 100 1818
rect 66 1725 100 1760
rect 66 1656 100 1691
rect 66 1587 100 1622
rect 3326 1794 3360 1818
rect 3326 1676 3360 1760
rect 3326 1618 3360 1642
rect 66 1518 100 1553
rect 66 1450 100 1484
rect 66 1382 100 1416
rect 66 1314 100 1348
rect 66 1246 100 1280
rect 66 1188 100 1212
<< mvpsubdiffcont >>
rect 304 978 338 1012
rect 304 907 338 941
rect 304 836 338 870
rect 304 765 338 799
rect 304 694 338 728
rect 304 623 338 657
rect 304 552 338 586
rect 304 481 338 515
rect 304 410 338 444
rect 304 340 338 374
rect 304 270 338 304
rect 304 200 338 234
rect 304 130 338 164
rect 304 60 338 94
rect 1240 978 1274 1012
rect 1240 907 1274 941
rect 1240 836 1274 870
rect 1240 765 1274 799
rect 1240 694 1274 728
rect 1240 623 1274 657
rect 1240 552 1274 586
rect 1240 481 1274 515
rect 1240 410 1274 444
rect 1240 340 1274 374
rect 1240 270 1274 304
rect 1240 200 1274 234
rect 1240 130 1274 164
rect 1240 60 1274 94
<< mvnsubdiffcont >>
rect 66 1760 100 1794
rect 66 1691 100 1725
rect 66 1622 100 1656
rect 3326 1760 3360 1794
rect 3326 1642 3360 1676
rect 66 1553 100 1587
rect 66 1484 100 1518
rect 66 1416 100 1450
rect 66 1348 100 1382
rect 66 1280 100 1314
rect 66 1212 100 1246
<< poly >>
rect 207 1844 775 1916
rect 939 1900 1141 1916
rect 939 1866 955 1900
rect 989 1866 1023 1900
rect 1057 1866 1091 1900
rect 1125 1866 1141 1900
rect 939 1844 1141 1866
rect 1197 1900 1399 1916
rect 1197 1866 1213 1900
rect 1247 1866 1281 1900
rect 1315 1866 1349 1900
rect 1383 1866 1399 1900
rect 1197 1844 1399 1866
rect 1563 1844 2363 1916
rect 2419 1844 3219 1916
rect 207 1150 775 1202
rect 207 1062 937 1150
rect 993 1118 1127 1134
rect 993 1084 1009 1118
rect 1043 1084 1077 1118
rect 1111 1084 1127 1118
rect 993 1062 1127 1084
<< polycont >>
rect 955 1866 989 1900
rect 1023 1866 1057 1900
rect 1091 1866 1125 1900
rect 1213 1866 1247 1900
rect 1281 1866 1315 1900
rect 1349 1866 1383 1900
rect 1009 1084 1043 1118
rect 1077 1084 1111 1118
<< locali >>
rect 939 1866 955 1900
rect 989 1866 1023 1900
rect 1057 1866 1091 1900
rect 1125 1866 1141 1900
rect 1197 1866 1213 1900
rect 1247 1866 1281 1900
rect 1315 1866 1349 1900
rect 1383 1866 1399 1900
rect 66 1794 100 1818
rect 977 1816 1107 1866
rect 977 1782 989 1816
rect 1023 1782 1061 1816
rect 1095 1782 1107 1816
rect 1234 1816 1364 1866
rect 1234 1782 1246 1816
rect 1280 1782 1318 1816
rect 1352 1782 1364 1816
rect 1510 1782 1548 1816
rect 3264 1794 3360 1822
rect 66 1728 100 1760
rect 3264 1760 3326 1794
rect 3264 1728 3360 1760
rect 66 1656 100 1691
rect 66 1587 100 1622
rect 1152 1652 1186 1690
rect 3346 1676 3360 1728
rect 3346 1622 3360 1642
rect 3264 1620 3360 1622
rect 3326 1618 3360 1620
rect 66 1518 100 1553
rect 630 1534 668 1568
rect 930 1534 968 1568
rect 66 1450 100 1484
rect 318 1460 356 1494
rect 1370 1460 1408 1494
rect 66 1382 100 1416
rect 66 1314 100 1348
rect 66 1246 100 1280
rect 162 1246 196 1280
rect 474 1246 508 1280
rect 786 1246 820 1280
rect 162 1212 820 1246
rect 66 1188 100 1212
rect 220 1158 898 1168
rect 220 1124 233 1158
rect 267 1124 305 1158
rect 339 1124 377 1158
rect 411 1124 449 1158
rect 483 1124 521 1158
rect 555 1124 593 1158
rect 627 1124 665 1158
rect 699 1124 898 1158
rect 220 1084 898 1124
rect 993 1158 1127 1164
rect 993 1124 1006 1158
rect 1040 1124 1078 1158
rect 1112 1124 1127 1158
rect 993 1118 1127 1124
rect 993 1084 1009 1118
rect 1043 1084 1077 1118
rect 1111 1084 1127 1118
rect 304 1012 338 1036
rect 304 941 338 978
rect 304 870 338 907
rect 1240 1012 1274 1036
rect 1240 941 1274 978
rect 1240 870 1274 907
rect 304 799 338 836
rect 454 820 492 854
rect 768 820 806 854
rect 1086 820 1124 854
rect 304 728 338 765
rect 304 657 338 694
rect 304 586 338 623
rect 1240 799 1274 836
rect 1240 728 1274 765
rect 1240 657 1274 694
rect 1240 586 1274 623
rect 304 515 338 518
rect 304 480 338 481
rect 304 444 338 446
rect 304 408 338 410
rect 596 480 630 518
rect 596 408 630 446
rect 948 480 982 518
rect 948 408 982 446
rect 1240 515 1274 518
rect 1240 480 1274 481
rect 1240 444 1274 446
rect 1240 408 1274 410
rect 304 304 338 340
rect 304 234 338 270
rect 304 164 338 200
rect 304 94 338 130
rect 304 36 338 60
rect 1240 304 1274 340
rect 1240 234 1274 270
rect 1240 164 1274 200
rect 1240 94 1274 130
rect 1240 36 1274 60
<< viali >>
rect 989 1782 1023 1816
rect 1061 1782 1095 1816
rect 1246 1782 1280 1816
rect 1318 1782 1352 1816
rect 1476 1782 1510 1816
rect 1548 1782 1582 1816
rect 66 1725 100 1728
rect 66 1694 100 1725
rect 66 1622 100 1656
rect 1152 1690 1186 1724
rect 1152 1618 1186 1652
rect 3240 1676 3346 1728
rect 3240 1642 3326 1676
rect 3326 1642 3346 1676
rect 3240 1622 3346 1642
rect 596 1534 630 1568
rect 668 1534 702 1568
rect 896 1534 930 1568
rect 968 1534 1002 1568
rect 284 1460 318 1494
rect 356 1460 390 1494
rect 1336 1460 1370 1494
rect 1408 1460 1442 1494
rect 233 1124 267 1158
rect 305 1124 339 1158
rect 377 1124 411 1158
rect 449 1124 483 1158
rect 521 1124 555 1158
rect 593 1124 627 1158
rect 665 1124 699 1158
rect 1006 1124 1040 1158
rect 1078 1124 1112 1158
rect 420 820 454 854
rect 492 820 526 854
rect 734 820 768 854
rect 806 820 840 854
rect 1052 820 1086 854
rect 1124 820 1158 854
rect 304 518 338 552
rect 304 446 338 480
rect 304 374 338 408
rect 596 518 630 552
rect 596 446 630 480
rect 596 374 630 408
rect 948 518 982 552
rect 948 446 982 480
rect 948 374 982 408
rect 1240 518 1274 552
rect 1240 446 1274 480
rect 1240 374 1274 408
<< metal1 >>
rect -227 1861 -221 1913
rect -169 1861 -157 1913
rect -105 1861 2353 1913
rect 2408 1861 2414 1913
rect 2466 1861 2478 1913
rect 2530 1861 3197 1913
rect 977 1816 1107 1822
rect 977 1782 989 1816
rect 1023 1782 1061 1816
rect 1095 1782 1107 1816
rect 977 1776 1107 1782
rect 1234 1816 1364 1822
rect 1234 1782 1246 1816
rect 1280 1782 1318 1816
rect 1352 1782 1364 1816
rect 1234 1776 1364 1782
rect 1464 1776 1470 1828
rect 1522 1776 1534 1828
rect 1586 1776 1594 1828
rect 0 1728 3426 1748
rect 0 1694 66 1728
rect 100 1724 3240 1728
rect 100 1694 1152 1724
rect 0 1690 1152 1694
rect 1186 1690 3240 1724
rect 0 1656 3240 1690
rect 0 1622 66 1656
rect 100 1652 3240 1656
rect 100 1622 1152 1652
rect 0 1618 1152 1622
rect 1186 1622 3240 1652
rect 3346 1622 3426 1728
rect 1186 1618 3426 1622
rect 0 1602 3426 1618
rect 584 1568 1014 1574
rect 584 1534 596 1568
rect 630 1534 668 1568
rect 702 1534 896 1568
rect 930 1534 968 1568
rect 1002 1534 1014 1568
rect 584 1528 1014 1534
rect 272 1494 1454 1500
rect 272 1460 284 1494
rect 318 1460 356 1494
rect 390 1460 1336 1494
rect 1370 1460 1408 1494
rect 1442 1460 1454 1494
rect 272 1454 1454 1460
rect -231 1204 -179 1210
tri -179 1198 -171 1206 sw
rect 150 1198 1470 1250
rect 1522 1198 1534 1250
rect 1586 1198 1592 1250
rect 2408 1240 2460 1246
rect -179 1170 -171 1198
tri -171 1170 -143 1198 sw
tri 2389 1170 2408 1189 se
rect 2408 1176 2460 1188
rect -179 1158 711 1170
tri 2383 1164 2389 1170 se
rect 2389 1164 2408 1170
rect -179 1152 233 1158
rect -231 1140 233 1152
rect -179 1124 233 1140
rect 267 1124 305 1158
rect 339 1124 377 1158
rect 411 1124 449 1158
rect 483 1124 521 1158
rect 555 1124 593 1158
rect 627 1124 665 1158
rect 699 1124 711 1158
rect -179 1118 711 1124
rect 993 1158 2408 1164
rect 993 1124 1006 1158
rect 1040 1124 1078 1158
rect 1112 1124 2408 1158
rect 993 1118 2460 1124
rect -231 1082 -179 1088
tri -179 1082 -143 1118 nw
rect 177 888 3426 1090
rect 408 854 1470 860
rect 408 820 420 854
rect 454 820 492 854
rect 526 820 734 854
rect 768 820 806 854
rect 840 820 1052 854
rect 1086 820 1124 854
rect 1158 820 1470 854
rect 408 808 1470 820
rect 1522 808 1534 860
rect 1586 808 1592 860
rect 0 552 1400 564
rect 0 518 304 552
rect 338 518 596 552
rect 630 518 948 552
rect 982 518 1240 552
rect 1274 519 1400 552
tri 1400 519 1445 564 sw
tri 1611 519 1656 564 se
rect 1656 519 3426 564
rect 1274 518 3426 519
rect 0 480 3426 518
rect 0 446 304 480
rect 338 446 596 480
rect 630 446 948 480
rect 982 446 1240 480
rect 1274 446 3426 480
rect 0 408 3426 446
rect 0 374 304 408
rect 338 374 596 408
rect 630 374 948 408
rect 982 374 1240 408
rect 1274 374 3426 408
rect 0 362 3426 374
<< via1 >>
rect -221 1861 -169 1913
rect -157 1861 -105 1913
rect 2414 1861 2466 1913
rect 2478 1861 2530 1913
rect 1470 1816 1522 1828
rect 1470 1782 1476 1816
rect 1476 1782 1510 1816
rect 1510 1782 1522 1816
rect 1470 1776 1522 1782
rect 1534 1816 1586 1828
rect 1534 1782 1548 1816
rect 1548 1782 1582 1816
rect 1582 1782 1586 1816
rect 1534 1776 1586 1782
rect -231 1152 -179 1204
rect 1470 1198 1522 1250
rect 1534 1198 1586 1250
rect 2408 1188 2460 1240
rect -231 1088 -179 1140
rect 2408 1124 2460 1176
rect 1470 808 1522 860
rect 1534 808 1586 860
<< metal2 >>
rect -227 1861 -221 1913
rect -169 1861 -157 1913
rect -105 1861 -99 1913
tri -307 1404 -227 1484 se
rect -227 1430 -99 1861
rect 2408 1861 2414 1913
rect 2466 1861 2478 1913
rect 2530 1861 2536 1913
rect -227 1404 -125 1430
tri -125 1404 -99 1430 nw
rect 1464 1776 1470 1828
rect 1522 1776 1534 1828
rect 1586 1776 1592 1828
rect -307 1204 -179 1404
tri -179 1350 -125 1404 nw
rect -307 1152 -231 1204
rect -307 1140 -179 1152
rect -307 1118 -231 1140
rect -231 1082 -179 1088
rect 1464 1250 1592 1776
rect 1464 1198 1470 1250
rect 1522 1198 1534 1250
rect 1586 1198 1592 1250
rect 1464 860 1592 1198
rect 2408 1240 2460 1861
tri 2460 1836 2485 1861 nw
rect 2408 1176 2460 1188
rect 2408 1118 2460 1124
rect 1464 808 1470 860
rect 1522 808 1534 860
rect 1586 808 1592 860
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1707688321
transform 0 -1 1186 -1 0 1724
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1707688321
transform 0 1 66 -1 0 1728
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1707688321
transform -1 0 526 0 1 820
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1707688321
transform -1 0 840 0 1 820
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1707688321
transform -1 0 1158 0 1 820
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1707688321
transform -1 0 1002 0 1 1534
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1707688321
transform -1 0 702 0 1 1534
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1707688321
transform -1 0 1442 0 1 1460
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1707688321
transform -1 0 390 0 1 1460
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_9
timestamp 1707688321
transform -1 0 1582 0 1 1782
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_10
timestamp 1707688321
transform -1 0 1352 0 1 1782
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_11
timestamp 1707688321
transform -1 0 1095 0 1 1782
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_12
timestamp 1707688321
transform -1 0 1112 0 1 1124
box 0 0 1 1
use L1M1_CDNS_5246887918559  L1M1_CDNS_5246887918559_0
timestamp 1707688321
transform 0 1 3240 -1 0 1728
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1707688321
transform 0 1 948 -1 0 552
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1707688321
transform 0 1 596 -1 0 552
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_2
timestamp 1707688321
transform 0 1 304 -1 0 552
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_3
timestamp 1707688321
transform 0 1 1240 -1 0 552
box 0 0 1 1
use L1M1_CDNS_52468879185194  L1M1_CDNS_52468879185194_0
timestamp 1707688321
transform -1 0 2341 0 1 1867
box -12 -6 766 40
use L1M1_CDNS_52468879185194  L1M1_CDNS_52468879185194_1
timestamp 1707688321
transform -1 0 3185 0 1 1867
box -12 -6 766 40
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_0
timestamp 1707688321
transform 1 0 221 0 1 1867
box -12 -6 550 40
use L1M1_CDNS_52468879185316  L1M1_CDNS_52468879185316_0
timestamp 1707688321
transform 1 0 162 0 1 1204
box -12 -6 622 40
use L1M1_CDNS_52468879185337  L1M1_CDNS_52468879185337_0
timestamp 1707688321
transform 1 0 233 0 1 1124
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1707688321
transform 0 -1 2460 -1 0 1246
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1707688321
transform 0 -1 -179 -1 0 1210
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1707688321
transform -1 0 1592 0 1 1776
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1707688321
transform -1 0 2536 0 1 1861
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1707688321
transform 1 0 1464 0 -1 1250
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_5
timestamp 1707688321
transform 1 0 -227 0 -1 1913
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_6
timestamp 1707688321
transform 1 0 1464 0 -1 860
box 0 0 1 1
use nfet_CDNS_52468879185343  nfet_CDNS_52468879185343_0
timestamp 1707688321
transform 1 0 993 0 -1 1036
box -79 -26 199 1026
use nfet_CDNS_524688791851403  nfet_CDNS_524688791851403_0
timestamp 1707688321
transform -1 0 937 0 -1 1036
box -79 -26 551 1026
use pfet_CDNS_52468879185323  pfet_CDNS_52468879185323_0
timestamp 1707688321
transform -1 0 1141 0 -1 1818
box -119 -66 319 666
use pfet_CDNS_52468879185323  pfet_CDNS_52468879185323_1
timestamp 1707688321
transform 1 0 1197 0 -1 1818
box -119 -66 319 666
use pfet_CDNS_52468879185324  pfet_CDNS_52468879185324_0
timestamp 1707688321
transform -1 0 463 0 -1 1818
box -119 -66 375 666
use pfet_CDNS_52468879185324  pfet_CDNS_52468879185324_1
timestamp 1707688321
transform 1 0 519 0 -1 1818
box -119 -66 375 666
use pfet_CDNS_52468879185325  pfet_CDNS_52468879185325_0
timestamp 1707688321
transform -1 0 3219 0 -1 1818
box -119 -66 1775 266
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1707688321
transform 0 1 993 -1 0 1134
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_0
timestamp 1707688321
transform 0 -1 1399 -1 0 1916
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_1
timestamp 1707688321
transform 0 1 939 -1 0 1916
box 0 0 1 1
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_0
timestamp 1707688321
transform 0 -1 3180 1 0 1850
box 0 0 66 746
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_1
timestamp 1707688321
transform 0 -1 2341 1 0 1850
box 0 0 66 746
use PYL1_CDNS_52468879185318  PYL1_CDNS_52468879185318_0
timestamp 1707688321
transform 0 -1 764 -1 0 1916
box 0 0 66 542
use PYL1_CDNS_52468879185370  PYL1_CDNS_52468879185370_0
timestamp 1707688321
transform 0 -1 898 -1 0 1134
box 0 0 66 678
<< labels >>
flabel comment s 2386 1810 2386 1810 0 FreeSans 300 90 0 0 int_slow
flabel comment s 1021 1913 1021 1913 0 FreeSans 300 0 0 0 en_fast_n<0>
flabel comment s 1337 1917 1337 1917 0 FreeSans 300 0 0 0 en_fast_n<1>
flabel comment s 1947 1924 1947 1924 0 FreeSans 300 0 0 0 drvlo_h_n
flabel comment s 536 844 536 844 0 FreeSans 300 0 0 0 pd_h
flabel comment s 438 1232 438 1232 0 FreeSans 300 0 0 0 pd_h
flabel comment s 1038 1484 1038 1484 0 FreeSans 300 0 0 0 intnr1
flabel comment s 869 1562 869 1562 0 FreeSans 300 0 0 0 intnr0
flabel comment s 565 1149 565 1149 3 FreeSans 300 180 0 0 drvlo_h_n
flabel comment s 3094 1686 3094 1686 0 FreeSans 300 0 0 0 vcc_io
flabel comment s 2630 1917 2630 1917 0 FreeSans 300 0 0 0 pden_h_n
flabel metal1 s 1081 1118 1127 1164 7 FreeSans 300 180 0 0 pden_h_n
port 1 nsew
flabel metal1 s 1545 1198 1592 1250 7 FreeSans 300 180 0 0 pd_h
port 2 nsew
flabel metal1 s 1234 1776 1282 1822 7 FreeSans 300 180 0 0 en_fast_n<1>
port 3 nsew
flabel metal1 s 977 1776 1023 1822 3 FreeSans 300 180 0 0 en_fast_n<0>
port 6 nsew
flabel metal1 s 209 1861 255 1913 3 FreeSans 300 180 0 0 drvlo_h_n
port 7 nsew
flabel metal1 s 3386 888 3426 1090 7 FreeSans 300 180 0 0 vcc_io
port 4 nsew
flabel metal1 s 177 888 217 1090 3 FreeSans 300 180 0 0 vcc_io
port 4 nsew
flabel metal1 s 0 362 40 564 3 FreeSans 300 180 0 0 vgnd_io
port 5 nsew
flabel metal1 s 0 1602 40 1748 3 FreeSans 300 180 0 0 vcc_io
port 4 nsew
flabel metal1 s 3386 362 3426 564 7 FreeSans 300 180 0 0 vgnd_io
port 5 nsew
flabel metal1 s 3386 1602 3426 1748 7 FreeSans 300 180 0 0 vcc_io
port 4 nsew
<< properties >>
string GDS_END 87871034
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87859750
string path 2.075 46.100 2.075 29.050 
<< end >>
