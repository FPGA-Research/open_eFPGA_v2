magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect 303 365 5779 4484
<< pwell >>
rect 144 4653 5974 4780
rect 144 4558 6144 4653
rect 5922 222 6144 4558
rect 144 0 6144 222
<< mvpsubdiff >>
rect 170 4720 194 4754
rect 228 4720 263 4754
rect 297 4720 332 4754
rect 366 4720 401 4754
rect 435 4720 470 4754
rect 504 4720 539 4754
rect 573 4720 608 4754
rect 642 4720 677 4754
rect 711 4720 746 4754
rect 780 4720 815 4754
rect 849 4720 884 4754
rect 918 4720 953 4754
rect 987 4720 1022 4754
rect 1056 4720 1091 4754
rect 1125 4720 1160 4754
rect 1194 4720 1229 4754
rect 1263 4720 1298 4754
rect 1332 4720 1367 4754
rect 1401 4720 1436 4754
rect 1470 4720 1505 4754
rect 1539 4720 1574 4754
rect 1608 4720 1643 4754
rect 1677 4720 1712 4754
rect 1746 4720 1781 4754
rect 1815 4720 1850 4754
rect 1884 4720 1919 4754
rect 1953 4720 1988 4754
rect 2022 4720 2057 4754
rect 2091 4720 2126 4754
rect 2160 4720 2195 4754
rect 2229 4720 2264 4754
rect 2298 4720 2333 4754
rect 2367 4720 2402 4754
rect 2436 4720 2471 4754
rect 2505 4720 2540 4754
rect 2574 4720 2609 4754
rect 2643 4720 2678 4754
rect 2712 4720 2747 4754
rect 2781 4720 2816 4754
rect 2850 4720 2885 4754
rect 2919 4720 2954 4754
rect 2988 4720 3023 4754
rect 3057 4720 3092 4754
rect 3126 4720 3161 4754
rect 3195 4720 3230 4754
rect 3264 4720 3299 4754
rect 3333 4720 3368 4754
rect 3402 4720 3437 4754
rect 3471 4720 3506 4754
rect 3540 4720 3575 4754
rect 3609 4720 3644 4754
rect 3678 4720 3713 4754
rect 3747 4720 3782 4754
rect 170 4686 3782 4720
rect 170 4652 194 4686
rect 228 4652 263 4686
rect 297 4652 332 4686
rect 366 4652 401 4686
rect 435 4652 470 4686
rect 504 4652 539 4686
rect 573 4652 608 4686
rect 642 4652 677 4686
rect 711 4652 746 4686
rect 780 4652 815 4686
rect 849 4652 884 4686
rect 918 4652 953 4686
rect 987 4652 1022 4686
rect 1056 4652 1091 4686
rect 1125 4652 1160 4686
rect 1194 4652 1229 4686
rect 1263 4652 1298 4686
rect 1332 4652 1367 4686
rect 1401 4652 1436 4686
rect 1470 4652 1505 4686
rect 1539 4652 1574 4686
rect 1608 4652 1643 4686
rect 1677 4652 1712 4686
rect 1746 4652 1781 4686
rect 1815 4652 1850 4686
rect 1884 4652 1919 4686
rect 1953 4652 1988 4686
rect 2022 4652 2057 4686
rect 2091 4652 2126 4686
rect 2160 4652 2195 4686
rect 2229 4652 2264 4686
rect 2298 4652 2333 4686
rect 2367 4652 2402 4686
rect 2436 4652 2471 4686
rect 2505 4652 2540 4686
rect 2574 4652 2609 4686
rect 2643 4652 2678 4686
rect 2712 4652 2747 4686
rect 2781 4652 2816 4686
rect 2850 4652 2885 4686
rect 2919 4652 2954 4686
rect 2988 4652 3023 4686
rect 3057 4652 3092 4686
rect 3126 4652 3161 4686
rect 3195 4652 3230 4686
rect 3264 4652 3299 4686
rect 3333 4652 3368 4686
rect 3402 4652 3437 4686
rect 3471 4652 3506 4686
rect 3540 4652 3575 4686
rect 3609 4652 3644 4686
rect 3678 4652 3713 4686
rect 3747 4652 3782 4686
rect 170 4618 3782 4652
rect 170 4584 194 4618
rect 228 4584 263 4618
rect 297 4584 332 4618
rect 366 4584 401 4618
rect 435 4584 470 4618
rect 504 4584 539 4618
rect 573 4584 608 4618
rect 642 4584 677 4618
rect 711 4584 746 4618
rect 780 4584 815 4618
rect 849 4584 884 4618
rect 918 4584 953 4618
rect 987 4584 1022 4618
rect 1056 4584 1091 4618
rect 1125 4584 1160 4618
rect 1194 4584 1229 4618
rect 1263 4584 1298 4618
rect 1332 4584 1367 4618
rect 1401 4584 1436 4618
rect 1470 4584 1505 4618
rect 1539 4584 1574 4618
rect 1608 4584 1643 4618
rect 1677 4584 1712 4618
rect 1746 4584 1781 4618
rect 1815 4584 1850 4618
rect 1884 4584 1919 4618
rect 1953 4584 1988 4618
rect 2022 4584 2057 4618
rect 2091 4584 2126 4618
rect 2160 4584 2195 4618
rect 2229 4584 2264 4618
rect 2298 4584 2333 4618
rect 2367 4584 2402 4618
rect 2436 4584 2471 4618
rect 2505 4584 2540 4618
rect 2574 4584 2609 4618
rect 2643 4584 2678 4618
rect 2712 4584 2747 4618
rect 2781 4584 2816 4618
rect 2850 4584 2885 4618
rect 2919 4584 2954 4618
rect 2988 4584 3023 4618
rect 3057 4584 3092 4618
rect 3126 4584 3161 4618
rect 3195 4584 3230 4618
rect 3264 4584 3299 4618
rect 3333 4584 3368 4618
rect 3402 4584 3437 4618
rect 3471 4584 3506 4618
rect 3540 4584 3575 4618
rect 3609 4584 3644 4618
rect 3678 4584 3713 4618
rect 3747 4584 3782 4618
rect 5924 4627 5948 4754
rect 5924 4584 6118 4627
rect 5948 4582 6118 4584
rect 5948 4548 6084 4582
rect 170 26 204 196
rect 5882 162 5948 196
rect 5882 128 6016 162
rect 5950 94 6016 128
rect 5950 60 6084 94
rect 5950 26 5984 60
rect 6018 26 6118 60
<< mvnsubdiff >>
rect 370 4355 5712 4398
rect 370 4321 470 4355
rect 504 4321 539 4355
rect 573 4321 608 4355
rect 642 4321 677 4355
rect 711 4321 746 4355
rect 780 4321 815 4355
rect 849 4321 884 4355
rect 918 4321 953 4355
rect 987 4321 1022 4355
rect 1056 4321 1091 4355
rect 1125 4321 1160 4355
rect 1194 4321 1229 4355
rect 1263 4321 1298 4355
rect 1332 4321 1367 4355
rect 1401 4321 1436 4355
rect 1470 4321 1505 4355
rect 1539 4321 1574 4355
rect 1608 4321 1643 4355
rect 1677 4321 1712 4355
rect 1746 4321 1781 4355
rect 1815 4321 1850 4355
rect 1884 4321 1919 4355
rect 1953 4321 1988 4355
rect 2022 4321 2057 4355
rect 2091 4321 2126 4355
rect 2160 4321 2195 4355
rect 2229 4321 2264 4355
rect 2298 4321 2333 4355
rect 2367 4321 2402 4355
rect 2436 4321 2471 4355
rect 370 4287 2471 4321
rect 370 4253 470 4287
rect 504 4253 539 4287
rect 573 4253 608 4287
rect 642 4253 677 4287
rect 711 4253 746 4287
rect 780 4253 815 4287
rect 849 4253 884 4287
rect 918 4253 953 4287
rect 987 4253 1022 4287
rect 1056 4253 1091 4287
rect 1125 4253 1160 4287
rect 1194 4253 1229 4287
rect 1263 4253 1298 4287
rect 1332 4253 1367 4287
rect 1401 4253 1436 4287
rect 1470 4253 1505 4287
rect 1539 4253 1574 4287
rect 1608 4253 1643 4287
rect 1677 4253 1712 4287
rect 1746 4253 1781 4287
rect 1815 4253 1850 4287
rect 1884 4253 1919 4287
rect 1953 4253 1988 4287
rect 2022 4253 2057 4287
rect 2091 4253 2126 4287
rect 2160 4253 2195 4287
rect 2229 4253 2264 4287
rect 2298 4253 2333 4287
rect 2367 4253 2402 4287
rect 2436 4253 2471 4287
rect 370 4219 2471 4253
rect 370 4185 470 4219
rect 504 4185 539 4219
rect 573 4185 608 4219
rect 642 4185 677 4219
rect 711 4185 746 4219
rect 780 4185 815 4219
rect 849 4185 884 4219
rect 918 4185 953 4219
rect 987 4185 1022 4219
rect 1056 4185 1091 4219
rect 1125 4185 1160 4219
rect 1194 4185 1229 4219
rect 1263 4185 1298 4219
rect 1332 4185 1367 4219
rect 1401 4185 1436 4219
rect 1470 4185 1505 4219
rect 1539 4185 1574 4219
rect 1608 4185 1643 4219
rect 1677 4185 1712 4219
rect 1746 4185 1781 4219
rect 1815 4185 1850 4219
rect 1884 4185 1919 4219
rect 1953 4185 1988 4219
rect 2022 4185 2057 4219
rect 2091 4185 2126 4219
rect 2160 4185 2195 4219
rect 2229 4185 2264 4219
rect 2298 4185 2333 4219
rect 2367 4185 2402 4219
rect 2436 4185 2471 4219
rect 370 4151 2471 4185
rect 370 4117 470 4151
rect 504 4117 539 4151
rect 573 4117 608 4151
rect 642 4117 677 4151
rect 711 4117 746 4151
rect 780 4117 815 4151
rect 849 4117 884 4151
rect 918 4117 953 4151
rect 987 4117 1022 4151
rect 1056 4117 1091 4151
rect 1125 4117 1160 4151
rect 1194 4117 1229 4151
rect 1263 4117 1298 4151
rect 1332 4117 1367 4151
rect 1401 4117 1436 4151
rect 1470 4117 1505 4151
rect 1539 4117 1574 4151
rect 1608 4117 1643 4151
rect 1677 4117 1712 4151
rect 1746 4117 1781 4151
rect 1815 4117 1850 4151
rect 1884 4117 1919 4151
rect 1953 4117 1988 4151
rect 2022 4117 2057 4151
rect 2091 4117 2126 4151
rect 2160 4117 2195 4151
rect 2229 4117 2264 4151
rect 2298 4117 2333 4151
rect 2367 4117 2402 4151
rect 2436 4117 2471 4151
rect 5633 4117 5712 4355
rect 370 4032 5712 4117
rect 370 3998 472 4032
rect 5402 3998 5437 4032
rect 5471 3998 5506 4032
rect 5540 3998 5575 4032
rect 5609 3998 5644 4032
rect 5678 3998 5712 4032
rect 404 3964 472 3998
rect 5368 3964 5712 3998
rect 370 3930 438 3964
rect 5368 3930 5403 3964
rect 5437 3930 5472 3964
rect 5506 3930 5541 3964
rect 5575 3930 5610 3964
rect 5644 3930 5712 3964
rect 370 3929 506 3930
rect 404 3895 506 3929
rect 370 3894 506 3895
rect 370 3860 438 3894
rect 472 3862 506 3894
rect 5300 3896 5610 3930
rect 5300 3862 5335 3896
rect 5369 3862 5404 3896
rect 5438 3862 5473 3896
rect 5507 3862 5542 3896
rect 472 3860 540 3862
rect 404 3826 540 3860
rect 370 3824 506 3826
rect 370 3791 438 3824
rect 404 3790 438 3791
rect 472 3792 506 3824
rect 472 3790 540 3792
rect 404 3757 540 3790
rect 370 3756 540 3757
rect 370 3754 506 3756
rect 370 3722 438 3754
rect 404 3720 438 3722
rect 472 3722 506 3754
rect 472 3720 540 3722
rect 404 3688 540 3720
rect 370 3686 540 3688
rect 370 3684 506 3686
rect 370 3653 438 3684
rect 404 3650 438 3653
rect 472 3652 506 3684
rect 472 3650 540 3652
rect 404 3619 540 3650
rect 370 3616 540 3619
rect 370 3614 506 3616
rect 370 3584 438 3614
rect 404 3580 438 3584
rect 472 3582 506 3614
rect 472 3580 540 3582
rect 404 3550 540 3580
rect 370 3546 540 3550
rect 370 3544 506 3546
rect 370 3515 438 3544
rect 404 3510 438 3515
rect 472 3512 506 3544
rect 472 3510 540 3512
rect 404 3481 540 3510
rect 370 3476 540 3481
rect 370 3474 506 3476
rect 370 3446 438 3474
rect 404 3440 438 3446
rect 472 3442 506 3474
rect 472 3440 540 3442
rect 404 3412 540 3440
rect 370 3406 540 3412
rect 370 3404 506 3406
rect 370 3377 438 3404
rect 404 3370 438 3377
rect 472 3372 506 3404
rect 472 3370 540 3372
rect 404 3343 540 3370
rect 370 3336 540 3343
rect 370 3334 506 3336
rect 370 3308 438 3334
rect 404 3300 438 3308
rect 472 3302 506 3334
rect 472 3300 540 3302
rect 404 3274 540 3300
rect 370 3266 540 3274
rect 370 3264 506 3266
rect 370 3239 438 3264
rect 404 3230 438 3239
rect 472 3232 506 3264
rect 472 3230 540 3232
rect 404 3205 540 3230
rect 370 3196 540 3205
rect 370 3194 506 3196
rect 370 3170 438 3194
rect 404 3160 438 3170
rect 472 3162 506 3194
rect 472 3160 540 3162
rect 404 3136 540 3160
rect 370 3126 540 3136
rect 370 3124 506 3126
rect 370 3101 438 3124
rect 404 3090 438 3101
rect 472 3092 506 3124
rect 472 3090 540 3092
rect 404 3067 540 3090
rect 370 3056 540 3067
rect 370 3054 506 3056
rect 370 3032 438 3054
rect 404 3020 438 3032
rect 472 3022 506 3054
rect 472 3020 540 3022
rect 404 2998 540 3020
rect 370 2986 540 2998
rect 370 2984 506 2986
rect 370 2963 438 2984
rect 404 2950 438 2963
rect 472 2952 506 2984
rect 472 2950 540 2952
rect 404 2929 540 2950
rect 370 2916 540 2929
rect 370 2914 506 2916
rect 370 2894 438 2914
rect 404 2880 438 2894
rect 472 2882 506 2914
rect 472 2880 540 2882
rect 404 2860 540 2880
rect 370 2846 540 2860
rect 370 2844 506 2846
rect 370 2825 438 2844
rect 404 2810 438 2825
rect 472 2812 506 2844
rect 472 2810 540 2812
rect 404 2791 540 2810
rect 370 2776 540 2791
rect 370 2774 506 2776
rect 370 2756 438 2774
rect 404 2740 438 2756
rect 472 2742 506 2774
rect 472 2740 540 2742
rect 404 2722 540 2740
rect 370 2706 540 2722
rect 370 2704 506 2706
rect 370 2687 438 2704
rect 404 2670 438 2687
rect 472 2672 506 2704
rect 472 2670 540 2672
rect 404 2653 540 2670
rect 370 2636 540 2653
rect 370 2634 506 2636
rect 370 2618 438 2634
rect 404 2600 438 2618
rect 472 2602 506 2634
rect 472 2600 540 2602
rect 404 2584 540 2600
rect 370 2566 540 2584
rect 370 2564 506 2566
rect 370 2549 438 2564
rect 404 2530 438 2549
rect 472 2532 506 2564
rect 472 2530 540 2532
rect 404 2515 540 2530
rect 370 2496 540 2515
rect 370 2494 506 2496
rect 370 2480 438 2494
rect 404 2460 438 2480
rect 472 2462 506 2494
rect 472 2460 540 2462
rect 404 2446 540 2460
rect 370 2426 540 2446
rect 370 2424 506 2426
rect 370 2411 438 2424
rect 404 2390 438 2411
rect 472 2392 506 2424
rect 472 2390 540 2392
rect 404 2377 540 2390
rect 370 2356 540 2377
rect 370 2354 506 2356
rect 370 2342 438 2354
rect 404 2320 438 2342
rect 472 2322 506 2354
rect 472 2320 540 2322
rect 404 2308 540 2320
rect 370 2286 540 2308
rect 370 2284 506 2286
rect 370 2273 438 2284
rect 404 2250 438 2273
rect 472 2252 506 2284
rect 472 2250 540 2252
rect 404 2239 540 2250
rect 370 2216 540 2239
rect 370 2214 506 2216
rect 370 2204 438 2214
rect 404 2180 438 2204
rect 472 2182 506 2214
rect 472 2180 540 2182
rect 404 2170 540 2180
rect 370 2146 540 2170
rect 370 2144 506 2146
rect 370 2135 438 2144
rect 404 2110 438 2135
rect 472 2112 506 2144
rect 472 2110 540 2112
rect 404 2101 540 2110
rect 370 2076 540 2101
rect 370 2075 506 2076
rect 370 2066 438 2075
rect 404 2041 438 2066
rect 472 2042 506 2075
rect 472 2041 540 2042
rect 404 2032 540 2041
rect 370 2006 540 2032
rect 370 1997 438 2006
rect 404 1972 438 1997
rect 472 1972 506 2006
rect 404 1963 540 1972
rect 370 1937 540 1963
rect 370 1929 438 1937
rect 404 1903 438 1929
rect 472 1903 506 1937
rect 404 1895 540 1903
rect 370 1868 540 1895
rect 370 1861 438 1868
rect 404 1834 438 1861
rect 472 1834 506 1868
rect 404 1827 540 1834
rect 370 1799 540 1827
rect 370 1793 438 1799
rect 404 1765 438 1793
rect 472 1765 506 1799
rect 404 1759 540 1765
rect 370 1730 540 1759
rect 370 1725 438 1730
rect 404 1696 438 1725
rect 472 1696 506 1730
rect 404 1691 540 1696
rect 370 1661 540 1691
rect 370 1657 438 1661
rect 404 1627 438 1657
rect 472 1627 506 1661
rect 404 1623 540 1627
rect 370 1592 540 1623
rect 370 1589 438 1592
rect 404 1558 438 1589
rect 472 1558 506 1592
rect 404 1555 540 1558
rect 370 1523 540 1555
rect 370 1521 438 1523
rect 404 1489 438 1521
rect 472 1489 506 1523
rect 404 1487 540 1489
rect 370 1454 540 1487
rect 370 1453 438 1454
rect 404 1420 438 1453
rect 472 1420 506 1454
rect 404 1419 540 1420
rect 370 1385 540 1419
rect 404 1351 438 1385
rect 472 1351 506 1385
rect 370 1283 540 1351
rect 404 1249 438 1283
rect 472 1249 506 1283
rect 370 1214 540 1249
rect 370 1212 438 1214
rect 404 1178 438 1212
rect 370 1141 438 1178
rect 404 1107 438 1141
rect 370 1070 438 1107
rect 404 1036 438 1070
rect 370 999 438 1036
rect 404 965 438 999
rect 370 928 438 965
rect 404 894 438 928
rect 370 857 438 894
rect 404 823 438 857
rect 370 786 438 823
rect 404 752 438 786
rect 370 715 438 752
rect 404 681 438 715
rect 370 644 438 681
rect 404 610 438 644
rect 370 573 438 610
rect 404 568 438 573
rect 5542 2603 5610 2638
rect 5576 2570 5610 2603
rect 5576 2569 5678 2570
rect 5542 2536 5678 2569
rect 5542 2535 5712 2536
rect 5542 2534 5610 2535
rect 5576 2501 5610 2534
rect 5644 2501 5712 2535
rect 5576 2500 5678 2501
rect 5542 2467 5678 2500
rect 5542 2466 5712 2467
rect 5542 2465 5610 2466
rect 5576 2432 5610 2465
rect 5644 2432 5712 2466
rect 5576 2431 5678 2432
rect 5542 2398 5678 2431
rect 5542 2397 5712 2398
rect 5542 2396 5610 2397
rect 5576 2363 5610 2396
rect 5644 2363 5712 2397
rect 5576 2362 5678 2363
rect 5542 2329 5678 2362
rect 5542 2328 5712 2329
rect 5542 2327 5610 2328
rect 5576 2294 5610 2327
rect 5644 2294 5712 2328
rect 5576 2293 5678 2294
rect 5542 2260 5678 2293
rect 5542 2259 5712 2260
rect 5542 2258 5610 2259
rect 5576 2225 5610 2258
rect 5644 2225 5712 2259
rect 5576 2224 5678 2225
rect 5542 2191 5678 2224
rect 5542 2190 5712 2191
rect 5542 2189 5610 2190
rect 5576 2156 5610 2189
rect 5644 2156 5712 2190
rect 5576 2155 5678 2156
rect 5542 2122 5678 2155
rect 5542 2121 5712 2122
rect 5542 2120 5610 2121
rect 5576 2087 5610 2120
rect 5644 2087 5712 2121
rect 5576 2086 5678 2087
rect 5542 2053 5678 2086
rect 5542 2052 5712 2053
rect 5542 2051 5610 2052
rect 5576 2018 5610 2051
rect 5644 2018 5712 2052
rect 5576 2017 5678 2018
rect 5542 1984 5678 2017
rect 5542 1983 5712 1984
rect 5542 1982 5610 1983
rect 5576 1949 5610 1982
rect 5644 1949 5712 1983
rect 5576 1948 5678 1949
rect 5542 1915 5678 1948
rect 5542 1914 5712 1915
rect 5542 1913 5610 1914
rect 5576 1880 5610 1913
rect 5644 1880 5712 1914
rect 5576 1879 5678 1880
rect 5542 1846 5678 1879
rect 5542 1845 5712 1846
rect 5542 1844 5610 1845
rect 5576 1811 5610 1844
rect 5644 1811 5712 1845
rect 5576 1810 5678 1811
rect 5542 1777 5678 1810
rect 5542 1776 5712 1777
rect 5542 1775 5610 1776
rect 5576 1742 5610 1775
rect 5644 1742 5712 1776
rect 5576 1741 5678 1742
rect 5542 1708 5678 1741
rect 5542 1707 5712 1708
rect 5542 1706 5610 1707
rect 5576 1673 5610 1706
rect 5644 1673 5712 1707
rect 5576 1672 5678 1673
rect 5542 1639 5678 1672
rect 5542 1638 5712 1639
rect 5542 1637 5610 1638
rect 5576 1604 5610 1637
rect 5644 1604 5712 1638
rect 5576 1603 5678 1604
rect 5542 1570 5678 1603
rect 5542 1569 5712 1570
rect 5542 1568 5610 1569
rect 5576 1535 5610 1568
rect 5644 1535 5712 1569
rect 5576 1534 5678 1535
rect 5542 1501 5678 1534
rect 5542 1500 5712 1501
rect 5542 1499 5610 1500
rect 5576 1466 5610 1499
rect 5644 1466 5712 1500
rect 5576 1465 5678 1466
rect 5542 1432 5678 1465
rect 5542 1431 5712 1432
rect 5542 1430 5610 1431
rect 5576 1397 5610 1430
rect 5644 1397 5712 1431
rect 5576 1396 5678 1397
rect 5542 1363 5678 1396
rect 5542 1362 5712 1363
rect 5542 1361 5610 1362
rect 5576 1328 5610 1361
rect 5644 1328 5712 1362
rect 5576 1327 5678 1328
rect 5542 1294 5678 1327
rect 5542 1293 5712 1294
rect 5542 1292 5610 1293
rect 5576 1259 5610 1292
rect 5644 1259 5712 1293
rect 5576 1258 5678 1259
rect 5542 1225 5678 1258
rect 5542 1224 5712 1225
rect 5542 1223 5610 1224
rect 5576 1190 5610 1223
rect 5644 1190 5712 1224
rect 5576 1189 5678 1190
rect 5542 1156 5678 1189
rect 5542 1155 5712 1156
rect 5542 1154 5610 1155
rect 5576 1121 5610 1154
rect 5644 1121 5712 1155
rect 5576 1120 5678 1121
rect 5542 1087 5678 1120
rect 5542 1086 5712 1087
rect 5542 1085 5610 1086
rect 5576 1052 5610 1085
rect 5644 1052 5712 1086
rect 5576 1051 5678 1052
rect 5542 1018 5678 1051
rect 5542 1017 5712 1018
rect 5542 1016 5610 1017
rect 5576 983 5610 1016
rect 5644 983 5712 1017
rect 5576 982 5678 983
rect 5542 949 5678 982
rect 5542 948 5712 949
rect 5542 947 5610 948
rect 5576 914 5610 947
rect 5644 914 5712 948
rect 5576 913 5678 914
rect 5542 880 5678 913
rect 5542 879 5712 880
rect 5542 878 5610 879
rect 5576 845 5610 878
rect 5644 845 5712 879
rect 5576 844 5678 845
rect 5542 811 5678 844
rect 5542 810 5712 811
rect 5542 809 5610 810
rect 5576 776 5610 809
rect 5644 776 5712 810
rect 5576 775 5678 776
rect 5542 742 5678 775
rect 5542 741 5712 742
rect 5542 740 5610 741
rect 5576 707 5610 740
rect 5644 707 5712 741
rect 5576 706 5678 707
rect 5542 673 5678 706
rect 5542 672 5712 673
rect 5542 671 5610 672
rect 5576 638 5610 671
rect 5644 638 5712 672
rect 5576 637 5678 638
rect 5542 604 5678 637
rect 5542 603 5712 604
rect 5542 602 5610 603
rect 540 568 575 602
rect 609 568 644 602
rect 678 568 713 602
rect 747 568 782 602
rect 404 539 782 568
rect 370 534 782 539
rect 5576 569 5610 602
rect 5644 569 5712 603
rect 5576 535 5678 569
rect 5576 534 5712 535
rect 370 500 438 534
rect 472 500 507 534
rect 541 500 576 534
rect 610 500 645 534
rect 679 500 714 534
rect 5644 500 5712 534
rect 370 466 714 500
rect 5610 466 5678 500
rect 370 432 404 466
rect 438 432 473 466
rect 507 432 542 466
rect 576 432 611 466
rect 645 432 680 466
rect 5610 432 5712 466
<< nsubdiffcont >>
rect 506 3722 540 3724
rect 506 3652 540 3686
rect 506 3582 540 3616
rect 506 3512 540 3546
rect 506 3442 540 3476
rect 506 3372 540 3406
rect 506 3302 540 3336
rect 506 3232 540 3266
rect 506 3162 540 3196
rect 506 3092 540 3126
rect 506 3022 540 3056
rect 506 2952 540 2986
rect 506 2882 540 2916
rect 506 2812 540 2846
rect 506 2742 540 2776
rect 506 2672 540 2706
rect 506 2602 540 2636
rect 506 2532 540 2566
rect 506 2462 540 2496
rect 506 2392 540 2426
rect 506 2322 540 2356
rect 506 2252 540 2286
rect 506 2182 540 2216
rect 506 2112 540 2146
rect 506 2042 540 2076
rect 506 1972 540 2006
rect 506 1903 540 1937
rect 506 1834 540 1868
rect 506 1765 540 1799
rect 506 1696 540 1730
rect 506 1627 540 1661
rect 506 1558 540 1592
rect 506 1489 540 1523
rect 506 1420 540 1454
rect 506 1351 540 1385
rect 506 1249 540 1283
rect 506 1180 540 1214
rect 506 1112 540 1146
rect 506 1044 540 1078
rect 506 976 540 1010
rect 506 908 540 942
rect 506 840 540 874
rect 506 772 540 806
rect 506 724 540 738
rect 5542 3658 5576 3692
rect 5542 3590 5576 3624
rect 5542 3522 5576 3556
rect 5542 3454 5576 3488
rect 5542 3386 5576 3420
rect 5542 3318 5576 3352
rect 5542 3250 5576 3284
rect 5542 3182 5576 3216
rect 5542 3114 5576 3148
rect 5542 3046 5576 3080
rect 5542 2978 5576 3012
rect 5542 2910 5576 2944
rect 5542 2842 5576 2876
rect 5542 2774 5576 2808
rect 5542 2706 5576 2740
rect 5542 2638 5576 2672
rect 5542 2569 5576 2603
rect 5542 2500 5576 2534
rect 5542 2431 5576 2465
rect 5542 2362 5576 2396
rect 5542 2293 5576 2327
rect 5542 2224 5576 2258
rect 5542 2155 5576 2189
rect 5542 2086 5576 2120
rect 5542 2017 5576 2051
rect 5542 1948 5576 1982
rect 5542 1879 5576 1913
rect 5542 1810 5576 1844
rect 5542 1741 5576 1775
rect 5542 1672 5576 1706
rect 5542 1603 5576 1637
rect 5542 1534 5576 1568
rect 5542 1465 5576 1499
rect 5542 1396 5576 1430
rect 5542 1327 5576 1361
rect 5542 1258 5576 1292
rect 5542 1189 5576 1223
rect 5542 1120 5576 1154
rect 5542 1051 5576 1085
rect 5542 982 5576 1016
rect 5542 913 5576 947
rect 5542 844 5576 878
rect 5542 775 5576 809
rect 5542 724 5576 740
<< mvpsubdiffcont >>
rect 194 4720 228 4754
rect 263 4720 297 4754
rect 332 4720 366 4754
rect 401 4720 435 4754
rect 470 4720 504 4754
rect 539 4720 573 4754
rect 608 4720 642 4754
rect 677 4720 711 4754
rect 746 4720 780 4754
rect 815 4720 849 4754
rect 884 4720 918 4754
rect 953 4720 987 4754
rect 1022 4720 1056 4754
rect 1091 4720 1125 4754
rect 1160 4720 1194 4754
rect 1229 4720 1263 4754
rect 1298 4720 1332 4754
rect 1367 4720 1401 4754
rect 1436 4720 1470 4754
rect 1505 4720 1539 4754
rect 1574 4720 1608 4754
rect 1643 4720 1677 4754
rect 1712 4720 1746 4754
rect 1781 4720 1815 4754
rect 1850 4720 1884 4754
rect 1919 4720 1953 4754
rect 1988 4720 2022 4754
rect 2057 4720 2091 4754
rect 2126 4720 2160 4754
rect 2195 4720 2229 4754
rect 2264 4720 2298 4754
rect 2333 4720 2367 4754
rect 2402 4720 2436 4754
rect 2471 4720 2505 4754
rect 2540 4720 2574 4754
rect 2609 4720 2643 4754
rect 2678 4720 2712 4754
rect 2747 4720 2781 4754
rect 2816 4720 2850 4754
rect 2885 4720 2919 4754
rect 2954 4720 2988 4754
rect 3023 4720 3057 4754
rect 3092 4720 3126 4754
rect 3161 4720 3195 4754
rect 3230 4720 3264 4754
rect 3299 4720 3333 4754
rect 3368 4720 3402 4754
rect 3437 4720 3471 4754
rect 3506 4720 3540 4754
rect 3575 4720 3609 4754
rect 3644 4720 3678 4754
rect 3713 4720 3747 4754
rect 194 4652 228 4686
rect 263 4652 297 4686
rect 332 4652 366 4686
rect 401 4652 435 4686
rect 470 4652 504 4686
rect 539 4652 573 4686
rect 608 4652 642 4686
rect 677 4652 711 4686
rect 746 4652 780 4686
rect 815 4652 849 4686
rect 884 4652 918 4686
rect 953 4652 987 4686
rect 1022 4652 1056 4686
rect 1091 4652 1125 4686
rect 1160 4652 1194 4686
rect 1229 4652 1263 4686
rect 1298 4652 1332 4686
rect 1367 4652 1401 4686
rect 1436 4652 1470 4686
rect 1505 4652 1539 4686
rect 1574 4652 1608 4686
rect 1643 4652 1677 4686
rect 1712 4652 1746 4686
rect 1781 4652 1815 4686
rect 1850 4652 1884 4686
rect 1919 4652 1953 4686
rect 1988 4652 2022 4686
rect 2057 4652 2091 4686
rect 2126 4652 2160 4686
rect 2195 4652 2229 4686
rect 2264 4652 2298 4686
rect 2333 4652 2367 4686
rect 2402 4652 2436 4686
rect 2471 4652 2505 4686
rect 2540 4652 2574 4686
rect 2609 4652 2643 4686
rect 2678 4652 2712 4686
rect 2747 4652 2781 4686
rect 2816 4652 2850 4686
rect 2885 4652 2919 4686
rect 2954 4652 2988 4686
rect 3023 4652 3057 4686
rect 3092 4652 3126 4686
rect 3161 4652 3195 4686
rect 3230 4652 3264 4686
rect 3299 4652 3333 4686
rect 3368 4652 3402 4686
rect 3437 4652 3471 4686
rect 3506 4652 3540 4686
rect 3575 4652 3609 4686
rect 3644 4652 3678 4686
rect 3713 4652 3747 4686
rect 194 4584 228 4618
rect 263 4584 297 4618
rect 332 4584 366 4618
rect 401 4584 435 4618
rect 470 4584 504 4618
rect 539 4584 573 4618
rect 608 4584 642 4618
rect 677 4584 711 4618
rect 746 4584 780 4618
rect 815 4584 849 4618
rect 884 4584 918 4618
rect 953 4584 987 4618
rect 1022 4584 1056 4618
rect 1091 4584 1125 4618
rect 1160 4584 1194 4618
rect 1229 4584 1263 4618
rect 1298 4584 1332 4618
rect 1367 4584 1401 4618
rect 1436 4584 1470 4618
rect 1505 4584 1539 4618
rect 1574 4584 1608 4618
rect 1643 4584 1677 4618
rect 1712 4584 1746 4618
rect 1781 4584 1815 4618
rect 1850 4584 1884 4618
rect 1919 4584 1953 4618
rect 1988 4584 2022 4618
rect 2057 4584 2091 4618
rect 2126 4584 2160 4618
rect 2195 4584 2229 4618
rect 2264 4584 2298 4618
rect 2333 4584 2367 4618
rect 2402 4584 2436 4618
rect 2471 4584 2505 4618
rect 2540 4584 2574 4618
rect 2609 4584 2643 4618
rect 2678 4584 2712 4618
rect 2747 4584 2781 4618
rect 2816 4584 2850 4618
rect 2885 4584 2919 4618
rect 2954 4584 2988 4618
rect 3023 4584 3057 4618
rect 3092 4584 3126 4618
rect 3161 4584 3195 4618
rect 3230 4584 3264 4618
rect 3299 4584 3333 4618
rect 3368 4584 3402 4618
rect 3437 4584 3471 4618
rect 3506 4584 3540 4618
rect 3575 4584 3609 4618
rect 3644 4584 3678 4618
rect 3713 4584 3747 4618
rect 3782 4584 5924 4754
rect 6084 4548 6118 4582
rect 204 128 5882 196
rect 5948 162 6118 4548
rect 204 26 5950 128
rect 6016 94 6118 162
rect 6084 60 6118 94
rect 5984 26 6018 60
<< mvnsubdiffcont >>
rect 470 4321 504 4355
rect 539 4321 573 4355
rect 608 4321 642 4355
rect 677 4321 711 4355
rect 746 4321 780 4355
rect 815 4321 849 4355
rect 884 4321 918 4355
rect 953 4321 987 4355
rect 1022 4321 1056 4355
rect 1091 4321 1125 4355
rect 1160 4321 1194 4355
rect 1229 4321 1263 4355
rect 1298 4321 1332 4355
rect 1367 4321 1401 4355
rect 1436 4321 1470 4355
rect 1505 4321 1539 4355
rect 1574 4321 1608 4355
rect 1643 4321 1677 4355
rect 1712 4321 1746 4355
rect 1781 4321 1815 4355
rect 1850 4321 1884 4355
rect 1919 4321 1953 4355
rect 1988 4321 2022 4355
rect 2057 4321 2091 4355
rect 2126 4321 2160 4355
rect 2195 4321 2229 4355
rect 2264 4321 2298 4355
rect 2333 4321 2367 4355
rect 2402 4321 2436 4355
rect 470 4253 504 4287
rect 539 4253 573 4287
rect 608 4253 642 4287
rect 677 4253 711 4287
rect 746 4253 780 4287
rect 815 4253 849 4287
rect 884 4253 918 4287
rect 953 4253 987 4287
rect 1022 4253 1056 4287
rect 1091 4253 1125 4287
rect 1160 4253 1194 4287
rect 1229 4253 1263 4287
rect 1298 4253 1332 4287
rect 1367 4253 1401 4287
rect 1436 4253 1470 4287
rect 1505 4253 1539 4287
rect 1574 4253 1608 4287
rect 1643 4253 1677 4287
rect 1712 4253 1746 4287
rect 1781 4253 1815 4287
rect 1850 4253 1884 4287
rect 1919 4253 1953 4287
rect 1988 4253 2022 4287
rect 2057 4253 2091 4287
rect 2126 4253 2160 4287
rect 2195 4253 2229 4287
rect 2264 4253 2298 4287
rect 2333 4253 2367 4287
rect 2402 4253 2436 4287
rect 470 4185 504 4219
rect 539 4185 573 4219
rect 608 4185 642 4219
rect 677 4185 711 4219
rect 746 4185 780 4219
rect 815 4185 849 4219
rect 884 4185 918 4219
rect 953 4185 987 4219
rect 1022 4185 1056 4219
rect 1091 4185 1125 4219
rect 1160 4185 1194 4219
rect 1229 4185 1263 4219
rect 1298 4185 1332 4219
rect 1367 4185 1401 4219
rect 1436 4185 1470 4219
rect 1505 4185 1539 4219
rect 1574 4185 1608 4219
rect 1643 4185 1677 4219
rect 1712 4185 1746 4219
rect 1781 4185 1815 4219
rect 1850 4185 1884 4219
rect 1919 4185 1953 4219
rect 1988 4185 2022 4219
rect 2057 4185 2091 4219
rect 2126 4185 2160 4219
rect 2195 4185 2229 4219
rect 2264 4185 2298 4219
rect 2333 4185 2367 4219
rect 2402 4185 2436 4219
rect 470 4117 504 4151
rect 539 4117 573 4151
rect 608 4117 642 4151
rect 677 4117 711 4151
rect 746 4117 780 4151
rect 815 4117 849 4151
rect 884 4117 918 4151
rect 953 4117 987 4151
rect 1022 4117 1056 4151
rect 1091 4117 1125 4151
rect 1160 4117 1194 4151
rect 1229 4117 1263 4151
rect 1298 4117 1332 4151
rect 1367 4117 1401 4151
rect 1436 4117 1470 4151
rect 1505 4117 1539 4151
rect 1574 4117 1608 4151
rect 1643 4117 1677 4151
rect 1712 4117 1746 4151
rect 1781 4117 1815 4151
rect 1850 4117 1884 4151
rect 1919 4117 1953 4151
rect 1988 4117 2022 4151
rect 2057 4117 2091 4151
rect 2126 4117 2160 4151
rect 2195 4117 2229 4151
rect 2264 4117 2298 4151
rect 2333 4117 2367 4151
rect 2402 4117 2436 4151
rect 2471 4117 5633 4355
rect 472 3998 5402 4032
rect 5437 3998 5471 4032
rect 5506 3998 5540 4032
rect 5575 3998 5609 4032
rect 5644 3998 5678 4032
rect 370 3964 404 3998
rect 472 3964 5368 3998
rect 438 3930 5368 3964
rect 5403 3930 5437 3964
rect 5472 3930 5506 3964
rect 5541 3930 5575 3964
rect 5610 3930 5644 3964
rect 370 3895 404 3929
rect 438 3860 472 3894
rect 506 3862 5300 3930
rect 5610 3896 5712 3930
rect 5335 3862 5369 3896
rect 5404 3862 5438 3896
rect 5473 3862 5507 3896
rect 370 3826 404 3860
rect 370 3757 404 3791
rect 438 3790 472 3824
rect 506 3792 540 3826
rect 370 3688 404 3722
rect 438 3720 472 3754
rect 506 3724 540 3756
rect 370 3619 404 3653
rect 438 3650 472 3684
rect 370 3550 404 3584
rect 438 3580 472 3614
rect 370 3481 404 3515
rect 438 3510 472 3544
rect 370 3412 404 3446
rect 438 3440 472 3474
rect 370 3343 404 3377
rect 438 3370 472 3404
rect 370 3274 404 3308
rect 438 3300 472 3334
rect 370 3205 404 3239
rect 438 3230 472 3264
rect 370 3136 404 3170
rect 438 3160 472 3194
rect 370 3067 404 3101
rect 438 3090 472 3124
rect 370 2998 404 3032
rect 438 3020 472 3054
rect 370 2929 404 2963
rect 438 2950 472 2984
rect 370 2860 404 2894
rect 438 2880 472 2914
rect 370 2791 404 2825
rect 438 2810 472 2844
rect 370 2722 404 2756
rect 438 2740 472 2774
rect 370 2653 404 2687
rect 438 2670 472 2704
rect 370 2584 404 2618
rect 438 2600 472 2634
rect 370 2515 404 2549
rect 438 2530 472 2564
rect 370 2446 404 2480
rect 438 2460 472 2494
rect 370 2377 404 2411
rect 438 2390 472 2424
rect 370 2308 404 2342
rect 438 2320 472 2354
rect 370 2239 404 2273
rect 438 2250 472 2284
rect 370 2170 404 2204
rect 438 2180 472 2214
rect 370 2101 404 2135
rect 438 2110 472 2144
rect 370 2032 404 2066
rect 438 2041 472 2075
rect 370 1963 404 1997
rect 438 1972 472 2006
rect 370 1895 404 1929
rect 438 1903 472 1937
rect 370 1827 404 1861
rect 438 1834 472 1868
rect 370 1759 404 1793
rect 438 1765 472 1799
rect 370 1691 404 1725
rect 438 1696 472 1730
rect 370 1623 404 1657
rect 438 1627 472 1661
rect 370 1555 404 1589
rect 438 1558 472 1592
rect 370 1487 404 1521
rect 438 1489 472 1523
rect 370 1419 404 1453
rect 438 1420 472 1454
rect 370 1351 404 1385
rect 438 1351 472 1385
rect 370 1249 404 1283
rect 438 1249 472 1283
rect 370 1178 404 1212
rect 438 1180 506 1214
rect 438 1146 540 1180
rect 370 1107 404 1141
rect 438 1112 506 1146
rect 438 1078 540 1112
rect 370 1036 404 1070
rect 438 1044 506 1078
rect 438 1010 540 1044
rect 370 965 404 999
rect 438 976 506 1010
rect 438 942 540 976
rect 370 894 404 928
rect 438 908 506 942
rect 438 874 540 908
rect 370 823 404 857
rect 438 840 506 874
rect 438 806 540 840
rect 370 752 404 786
rect 438 772 506 806
rect 438 738 540 772
rect 438 724 506 738
rect 370 681 404 715
rect 370 610 404 644
rect 370 539 404 573
rect 438 568 540 724
rect 5542 3692 5712 3896
rect 5576 3658 5712 3692
rect 5542 3624 5712 3658
rect 5576 3590 5712 3624
rect 5542 3556 5712 3590
rect 5576 3522 5712 3556
rect 5542 3488 5712 3522
rect 5576 3454 5712 3488
rect 5542 3420 5712 3454
rect 5576 3386 5712 3420
rect 5542 3352 5712 3386
rect 5576 3318 5712 3352
rect 5542 3284 5712 3318
rect 5576 3250 5712 3284
rect 5542 3216 5712 3250
rect 5576 3182 5712 3216
rect 5542 3148 5712 3182
rect 5576 3114 5712 3148
rect 5542 3080 5712 3114
rect 5576 3046 5712 3080
rect 5542 3012 5712 3046
rect 5576 2978 5712 3012
rect 5542 2944 5712 2978
rect 5576 2910 5712 2944
rect 5542 2876 5712 2910
rect 5576 2842 5712 2876
rect 5542 2808 5712 2842
rect 5576 2774 5712 2808
rect 5542 2740 5712 2774
rect 5576 2706 5712 2740
rect 5542 2672 5712 2706
rect 5576 2638 5712 2672
rect 5610 2570 5712 2638
rect 5678 2536 5712 2570
rect 5610 2501 5644 2535
rect 5678 2467 5712 2501
rect 5610 2432 5644 2466
rect 5678 2398 5712 2432
rect 5610 2363 5644 2397
rect 5678 2329 5712 2363
rect 5610 2294 5644 2328
rect 5678 2260 5712 2294
rect 5610 2225 5644 2259
rect 5678 2191 5712 2225
rect 5610 2156 5644 2190
rect 5678 2122 5712 2156
rect 5610 2087 5644 2121
rect 5678 2053 5712 2087
rect 5610 2018 5644 2052
rect 5678 1984 5712 2018
rect 5610 1949 5644 1983
rect 5678 1915 5712 1949
rect 5610 1880 5644 1914
rect 5678 1846 5712 1880
rect 5610 1811 5644 1845
rect 5678 1777 5712 1811
rect 5610 1742 5644 1776
rect 5678 1708 5712 1742
rect 5610 1673 5644 1707
rect 5678 1639 5712 1673
rect 5610 1604 5644 1638
rect 5678 1570 5712 1604
rect 5610 1535 5644 1569
rect 5678 1501 5712 1535
rect 5610 1466 5644 1500
rect 5678 1432 5712 1466
rect 5610 1397 5644 1431
rect 5678 1363 5712 1397
rect 5610 1328 5644 1362
rect 5678 1294 5712 1328
rect 5610 1259 5644 1293
rect 5678 1225 5712 1259
rect 5610 1190 5644 1224
rect 5678 1156 5712 1190
rect 5610 1121 5644 1155
rect 5678 1087 5712 1121
rect 5610 1052 5644 1086
rect 5678 1018 5712 1052
rect 5610 983 5644 1017
rect 5678 949 5712 983
rect 5610 914 5644 948
rect 5678 880 5712 914
rect 5610 845 5644 879
rect 5678 811 5712 845
rect 5610 776 5644 810
rect 5678 742 5712 776
rect 5542 706 5576 724
rect 5610 707 5644 741
rect 5678 673 5712 707
rect 5542 637 5576 671
rect 5610 638 5644 672
rect 5678 604 5712 638
rect 575 568 609 602
rect 644 568 678 602
rect 713 568 747 602
rect 782 534 5576 602
rect 5610 569 5644 603
rect 5678 535 5712 569
rect 438 500 472 534
rect 507 500 541 534
rect 576 500 610 534
rect 645 500 679 534
rect 714 500 5644 534
rect 714 466 5610 500
rect 5678 466 5712 500
rect 404 432 438 466
rect 473 432 507 466
rect 542 432 576 466
rect 611 432 645 466
rect 680 432 5610 466
<< poly >>
rect 687 3806 1255 3822
rect 687 3772 703 3806
rect 737 3772 774 3806
rect 808 3772 845 3806
rect 879 3772 917 3806
rect 951 3772 989 3806
rect 1023 3772 1061 3806
rect 1095 3772 1133 3806
rect 1167 3772 1205 3806
rect 1239 3772 1255 3806
rect 687 3750 1255 3772
rect 1515 3806 2083 3822
rect 1515 3772 1531 3806
rect 1565 3772 1602 3806
rect 1636 3772 1673 3806
rect 1707 3772 1745 3806
rect 1779 3772 1817 3806
rect 1851 3772 1889 3806
rect 1923 3772 1961 3806
rect 1995 3772 2033 3806
rect 2067 3772 2083 3806
rect 1515 3750 2083 3772
rect 2343 3806 2911 3822
rect 2343 3772 2359 3806
rect 2393 3772 2430 3806
rect 2464 3772 2501 3806
rect 2535 3772 2573 3806
rect 2607 3772 2645 3806
rect 2679 3772 2717 3806
rect 2751 3772 2789 3806
rect 2823 3772 2861 3806
rect 2895 3772 2911 3806
rect 2343 3750 2911 3772
rect 3171 3806 3739 3822
rect 3171 3772 3187 3806
rect 3221 3772 3258 3806
rect 3292 3772 3329 3806
rect 3363 3772 3401 3806
rect 3435 3772 3473 3806
rect 3507 3772 3545 3806
rect 3579 3772 3617 3806
rect 3651 3772 3689 3806
rect 3723 3772 3739 3806
rect 3171 3750 3739 3772
rect 3998 3806 4567 3822
rect 3998 3772 4014 3806
rect 4048 3772 4085 3806
rect 4119 3772 4157 3806
rect 4191 3772 4229 3806
rect 4263 3772 4301 3806
rect 4335 3772 4373 3806
rect 4407 3772 4445 3806
rect 4479 3772 4517 3806
rect 4551 3772 4567 3806
rect 3998 3756 4567 3772
rect 3999 3750 4567 3756
rect 4827 3806 5395 3822
rect 4827 3772 4843 3806
rect 4877 3772 4914 3806
rect 4948 3772 4985 3806
rect 5019 3772 5057 3806
rect 5091 3772 5129 3806
rect 5163 3772 5201 3806
rect 5235 3772 5273 3806
rect 5307 3772 5345 3806
rect 5379 3772 5395 3806
rect 4827 3750 5395 3772
rect 687 676 1255 698
rect 687 642 703 676
rect 737 642 774 676
rect 808 642 845 676
rect 879 642 917 676
rect 951 642 989 676
rect 1023 642 1061 676
rect 1095 642 1133 676
rect 1167 642 1205 676
rect 1239 642 1255 676
rect 687 626 1255 642
rect 1515 676 2083 698
rect 1515 642 1531 676
rect 1565 642 1602 676
rect 1636 642 1673 676
rect 1707 642 1745 676
rect 1779 642 1817 676
rect 1851 642 1889 676
rect 1923 642 1961 676
rect 1995 642 2033 676
rect 2067 642 2083 676
rect 1515 626 2083 642
rect 2343 676 2911 698
rect 2343 642 2359 676
rect 2393 642 2430 676
rect 2464 642 2501 676
rect 2535 642 2573 676
rect 2607 642 2645 676
rect 2679 642 2717 676
rect 2751 642 2789 676
rect 2823 642 2861 676
rect 2895 642 2911 676
rect 2343 626 2911 642
rect 3171 676 3739 698
rect 3171 642 3187 676
rect 3221 642 3258 676
rect 3292 642 3329 676
rect 3363 642 3401 676
rect 3435 642 3473 676
rect 3507 642 3545 676
rect 3579 642 3617 676
rect 3651 642 3689 676
rect 3723 642 3739 676
rect 3171 626 3739 642
rect 3999 676 4567 698
rect 3999 642 4015 676
rect 4049 642 4086 676
rect 4120 642 4157 676
rect 4191 642 4229 676
rect 4263 642 4301 676
rect 4335 642 4373 676
rect 4407 642 4445 676
rect 4479 642 4517 676
rect 4551 642 4567 676
rect 3999 626 4567 642
rect 4827 676 5395 698
rect 4827 642 4843 676
rect 4877 642 4914 676
rect 4948 642 4985 676
rect 5019 642 5057 676
rect 5091 642 5129 676
rect 5163 642 5201 676
rect 5235 642 5273 676
rect 5307 642 5345 676
rect 5379 642 5395 676
rect 4827 626 5395 642
<< polycont >>
rect 703 3772 737 3806
rect 774 3772 808 3806
rect 845 3772 879 3806
rect 917 3772 951 3806
rect 989 3772 1023 3806
rect 1061 3772 1095 3806
rect 1133 3772 1167 3806
rect 1205 3772 1239 3806
rect 1531 3772 1565 3806
rect 1602 3772 1636 3806
rect 1673 3772 1707 3806
rect 1745 3772 1779 3806
rect 1817 3772 1851 3806
rect 1889 3772 1923 3806
rect 1961 3772 1995 3806
rect 2033 3772 2067 3806
rect 2359 3772 2393 3806
rect 2430 3772 2464 3806
rect 2501 3772 2535 3806
rect 2573 3772 2607 3806
rect 2645 3772 2679 3806
rect 2717 3772 2751 3806
rect 2789 3772 2823 3806
rect 2861 3772 2895 3806
rect 3187 3772 3221 3806
rect 3258 3772 3292 3806
rect 3329 3772 3363 3806
rect 3401 3772 3435 3806
rect 3473 3772 3507 3806
rect 3545 3772 3579 3806
rect 3617 3772 3651 3806
rect 3689 3772 3723 3806
rect 4014 3772 4048 3806
rect 4085 3772 4119 3806
rect 4157 3772 4191 3806
rect 4229 3772 4263 3806
rect 4301 3772 4335 3806
rect 4373 3772 4407 3806
rect 4445 3772 4479 3806
rect 4517 3772 4551 3806
rect 4843 3772 4877 3806
rect 4914 3772 4948 3806
rect 4985 3772 5019 3806
rect 5057 3772 5091 3806
rect 5129 3772 5163 3806
rect 5201 3772 5235 3806
rect 5273 3772 5307 3806
rect 5345 3772 5379 3806
rect 703 642 737 676
rect 774 642 808 676
rect 845 642 879 676
rect 917 642 951 676
rect 989 642 1023 676
rect 1061 642 1095 676
rect 1133 642 1167 676
rect 1205 642 1239 676
rect 1531 642 1565 676
rect 1602 642 1636 676
rect 1673 642 1707 676
rect 1745 642 1779 676
rect 1817 642 1851 676
rect 1889 642 1923 676
rect 1961 642 1995 676
rect 2033 642 2067 676
rect 2359 642 2393 676
rect 2430 642 2464 676
rect 2501 642 2535 676
rect 2573 642 2607 676
rect 2645 642 2679 676
rect 2717 642 2751 676
rect 2789 642 2823 676
rect 2861 642 2895 676
rect 3187 642 3221 676
rect 3258 642 3292 676
rect 3329 642 3363 676
rect 3401 642 3435 676
rect 3473 642 3507 676
rect 3545 642 3579 676
rect 3617 642 3651 676
rect 3689 642 3723 676
rect 4015 642 4049 676
rect 4086 642 4120 676
rect 4157 642 4191 676
rect 4229 642 4263 676
rect 4301 642 4335 676
rect 4373 642 4407 676
rect 4445 642 4479 676
rect 4517 642 4551 676
rect 4843 642 4877 676
rect 4914 642 4948 676
rect 4985 642 5019 676
rect 5057 642 5091 676
rect 5129 642 5163 676
rect 5201 642 5235 676
rect 5273 642 5307 676
rect 5345 642 5379 676
<< locali >>
rect 170 4720 194 4754
rect 228 4734 263 4754
rect 297 4734 332 4754
rect 366 4734 401 4754
rect 435 4734 470 4754
rect 504 4734 539 4754
rect 243 4720 263 4734
rect 316 4720 332 4734
rect 389 4720 401 4734
rect 462 4720 470 4734
rect 535 4720 539 4734
rect 573 4734 608 4754
rect 573 4720 574 4734
rect 170 4700 209 4720
rect 243 4700 282 4720
rect 316 4700 355 4720
rect 389 4700 428 4720
rect 462 4700 501 4720
rect 535 4700 574 4720
rect 642 4734 677 4754
rect 711 4734 746 4754
rect 780 4734 815 4754
rect 849 4734 884 4754
rect 918 4734 953 4754
rect 987 4734 1022 4754
rect 1056 4734 1091 4754
rect 1125 4734 1160 4754
rect 642 4720 647 4734
rect 711 4720 720 4734
rect 780 4720 793 4734
rect 849 4720 866 4734
rect 918 4720 939 4734
rect 987 4720 1012 4734
rect 1056 4720 1085 4734
rect 1125 4720 1158 4734
rect 1194 4720 1229 4754
rect 1263 4734 1298 4754
rect 1332 4734 1367 4754
rect 1401 4734 1436 4754
rect 1470 4734 1505 4754
rect 1539 4734 1574 4754
rect 1608 4734 1643 4754
rect 1677 4734 1712 4754
rect 1746 4734 1781 4754
rect 1265 4720 1298 4734
rect 1338 4720 1367 4734
rect 1411 4720 1436 4734
rect 1484 4720 1505 4734
rect 1557 4720 1574 4734
rect 1630 4720 1643 4734
rect 1703 4720 1712 4734
rect 1776 4720 1781 4734
rect 1815 4734 1850 4754
rect 608 4700 647 4720
rect 681 4700 720 4720
rect 754 4700 793 4720
rect 827 4700 866 4720
rect 900 4700 939 4720
rect 973 4700 1012 4720
rect 1046 4700 1085 4720
rect 1119 4700 1158 4720
rect 1192 4700 1231 4720
rect 1265 4700 1304 4720
rect 1338 4700 1377 4720
rect 1411 4700 1450 4720
rect 1484 4700 1523 4720
rect 1557 4700 1596 4720
rect 1630 4700 1669 4720
rect 1703 4700 1742 4720
rect 1776 4700 1815 4720
rect 1849 4720 1850 4734
rect 1884 4734 1919 4754
rect 1953 4734 1988 4754
rect 2022 4734 2057 4754
rect 2091 4734 2126 4754
rect 2160 4734 2195 4754
rect 2229 4734 2264 4754
rect 2298 4734 2333 4754
rect 2367 4734 2402 4754
rect 1884 4720 1888 4734
rect 1953 4720 1961 4734
rect 2022 4720 2034 4734
rect 2091 4720 2107 4734
rect 2160 4720 2180 4734
rect 2229 4720 2253 4734
rect 2298 4720 2326 4734
rect 2367 4720 2399 4734
rect 2436 4720 2471 4754
rect 2505 4734 2540 4754
rect 2574 4734 2609 4754
rect 2643 4734 2678 4754
rect 2712 4734 2747 4754
rect 2781 4734 2816 4754
rect 2850 4734 2885 4754
rect 2919 4734 2954 4754
rect 2988 4734 3023 4754
rect 3057 4734 3092 4754
rect 2506 4720 2540 4734
rect 2579 4720 2609 4734
rect 2652 4720 2678 4734
rect 2725 4720 2747 4734
rect 2798 4720 2816 4734
rect 2871 4720 2885 4734
rect 2944 4720 2954 4734
rect 3017 4720 3023 4734
rect 3090 4720 3092 4734
rect 3126 4734 3161 4754
rect 3195 4734 3230 4754
rect 3264 4734 3299 4754
rect 3333 4734 3368 4754
rect 3402 4734 3437 4754
rect 3471 4734 3506 4754
rect 3540 4734 3575 4754
rect 3609 4734 3644 4754
rect 3126 4720 3129 4734
rect 3195 4720 3202 4734
rect 3264 4720 3275 4734
rect 3333 4720 3348 4734
rect 3402 4720 3421 4734
rect 3471 4720 3494 4734
rect 3540 4720 3567 4734
rect 3609 4720 3640 4734
rect 3678 4720 3713 4754
rect 1849 4700 1888 4720
rect 1922 4700 1961 4720
rect 1995 4700 2034 4720
rect 2068 4700 2107 4720
rect 2141 4700 2180 4720
rect 2214 4700 2253 4720
rect 2287 4700 2326 4720
rect 2360 4700 2399 4720
rect 2433 4700 2472 4720
rect 2506 4700 2545 4720
rect 2579 4700 2618 4720
rect 2652 4700 2691 4720
rect 2725 4700 2764 4720
rect 2798 4700 2837 4720
rect 2871 4700 2910 4720
rect 2944 4700 2983 4720
rect 3017 4700 3056 4720
rect 3090 4700 3129 4720
rect 3163 4700 3202 4720
rect 3236 4700 3275 4720
rect 3309 4700 3348 4720
rect 3382 4700 3421 4720
rect 3455 4700 3494 4720
rect 3528 4700 3567 4720
rect 3601 4700 3640 4720
rect 3674 4700 3713 4720
rect 3747 4700 3782 4754
rect 170 4686 3782 4700
rect 170 4652 194 4686
rect 228 4662 263 4686
rect 297 4662 332 4686
rect 366 4662 401 4686
rect 435 4662 470 4686
rect 504 4662 539 4686
rect 243 4652 263 4662
rect 316 4652 332 4662
rect 389 4652 401 4662
rect 462 4652 470 4662
rect 535 4652 539 4662
rect 573 4662 608 4686
rect 573 4652 574 4662
rect 170 4628 209 4652
rect 243 4628 282 4652
rect 316 4628 355 4652
rect 389 4628 428 4652
rect 462 4628 501 4652
rect 535 4628 574 4652
rect 642 4662 677 4686
rect 711 4662 746 4686
rect 780 4662 815 4686
rect 849 4662 884 4686
rect 918 4662 953 4686
rect 987 4662 1022 4686
rect 1056 4662 1091 4686
rect 1125 4662 1160 4686
rect 642 4652 647 4662
rect 711 4652 720 4662
rect 780 4652 793 4662
rect 849 4652 866 4662
rect 918 4652 939 4662
rect 987 4652 1012 4662
rect 1056 4652 1085 4662
rect 1125 4652 1158 4662
rect 1194 4652 1229 4686
rect 1263 4662 1298 4686
rect 1332 4662 1367 4686
rect 1401 4662 1436 4686
rect 1470 4662 1505 4686
rect 1539 4662 1574 4686
rect 1608 4662 1643 4686
rect 1677 4662 1712 4686
rect 1746 4662 1781 4686
rect 1265 4652 1298 4662
rect 1338 4652 1367 4662
rect 1411 4652 1436 4662
rect 1484 4652 1505 4662
rect 1557 4652 1574 4662
rect 1630 4652 1643 4662
rect 1703 4652 1712 4662
rect 1776 4652 1781 4662
rect 1815 4662 1850 4686
rect 608 4628 647 4652
rect 681 4628 720 4652
rect 754 4628 793 4652
rect 827 4628 866 4652
rect 900 4628 939 4652
rect 973 4628 1012 4652
rect 1046 4628 1085 4652
rect 1119 4628 1158 4652
rect 1192 4628 1231 4652
rect 1265 4628 1304 4652
rect 1338 4628 1377 4652
rect 1411 4628 1450 4652
rect 1484 4628 1523 4652
rect 1557 4628 1596 4652
rect 1630 4628 1669 4652
rect 1703 4628 1742 4652
rect 1776 4628 1815 4652
rect 1849 4652 1850 4662
rect 1884 4662 1919 4686
rect 1953 4662 1988 4686
rect 2022 4662 2057 4686
rect 2091 4662 2126 4686
rect 2160 4662 2195 4686
rect 2229 4662 2264 4686
rect 2298 4662 2333 4686
rect 2367 4662 2402 4686
rect 1884 4652 1888 4662
rect 1953 4652 1961 4662
rect 2022 4652 2034 4662
rect 2091 4652 2107 4662
rect 2160 4652 2180 4662
rect 2229 4652 2253 4662
rect 2298 4652 2326 4662
rect 2367 4652 2399 4662
rect 2436 4652 2471 4686
rect 2505 4662 2540 4686
rect 2574 4662 2609 4686
rect 2643 4662 2678 4686
rect 2712 4662 2747 4686
rect 2781 4662 2816 4686
rect 2850 4662 2885 4686
rect 2919 4662 2954 4686
rect 2988 4662 3023 4686
rect 3057 4662 3092 4686
rect 2506 4652 2540 4662
rect 2579 4652 2609 4662
rect 2652 4652 2678 4662
rect 2725 4652 2747 4662
rect 2798 4652 2816 4662
rect 2871 4652 2885 4662
rect 2944 4652 2954 4662
rect 3017 4652 3023 4662
rect 3090 4652 3092 4662
rect 3126 4662 3161 4686
rect 3195 4662 3230 4686
rect 3264 4662 3299 4686
rect 3333 4662 3368 4686
rect 3402 4662 3437 4686
rect 3471 4662 3506 4686
rect 3540 4662 3575 4686
rect 3609 4662 3644 4686
rect 3126 4652 3129 4662
rect 3195 4652 3202 4662
rect 3264 4652 3275 4662
rect 3333 4652 3348 4662
rect 3402 4652 3421 4662
rect 3471 4652 3494 4662
rect 3540 4652 3567 4662
rect 3609 4652 3640 4662
rect 3678 4652 3713 4686
rect 1849 4628 1888 4652
rect 1922 4628 1961 4652
rect 1995 4628 2034 4652
rect 2068 4628 2107 4652
rect 2141 4628 2180 4652
rect 2214 4628 2253 4652
rect 2287 4628 2326 4652
rect 2360 4628 2399 4652
rect 2433 4628 2472 4652
rect 2506 4628 2545 4652
rect 2579 4628 2618 4652
rect 2652 4628 2691 4652
rect 2725 4628 2764 4652
rect 2798 4628 2837 4652
rect 2871 4628 2910 4652
rect 2944 4628 2983 4652
rect 3017 4628 3056 4652
rect 3090 4628 3129 4652
rect 3163 4628 3202 4652
rect 3236 4628 3275 4652
rect 3309 4628 3348 4652
rect 3382 4628 3421 4652
rect 3455 4628 3494 4652
rect 3528 4628 3567 4652
rect 3601 4628 3640 4652
rect 3674 4628 3713 4652
rect 3747 4628 3782 4686
rect 170 4618 3782 4628
rect 170 4584 194 4618
rect 228 4584 263 4618
rect 297 4584 332 4618
rect 366 4584 401 4618
rect 435 4584 470 4618
rect 504 4584 539 4618
rect 573 4584 608 4618
rect 642 4584 677 4618
rect 711 4584 746 4618
rect 780 4584 815 4618
rect 849 4584 884 4618
rect 918 4584 953 4618
rect 987 4584 1022 4618
rect 1056 4584 1091 4618
rect 1125 4584 1160 4618
rect 1194 4584 1229 4618
rect 1263 4584 1298 4618
rect 1332 4584 1367 4618
rect 1401 4584 1436 4618
rect 1470 4584 1505 4618
rect 1539 4584 1574 4618
rect 1608 4584 1643 4618
rect 1677 4584 1712 4618
rect 1746 4584 1781 4618
rect 1815 4584 1850 4618
rect 1884 4584 1919 4618
rect 1953 4584 1988 4618
rect 2022 4584 2057 4618
rect 2091 4584 2126 4618
rect 2160 4584 2195 4618
rect 2229 4584 2264 4618
rect 2298 4584 2333 4618
rect 2367 4584 2402 4618
rect 2436 4584 2471 4618
rect 2505 4584 2540 4618
rect 2574 4584 2609 4618
rect 2643 4584 2678 4618
rect 2712 4584 2747 4618
rect 2781 4584 2816 4618
rect 2850 4584 2885 4618
rect 2919 4584 2954 4618
rect 2988 4584 3023 4618
rect 3057 4584 3092 4618
rect 3126 4584 3161 4618
rect 3195 4584 3230 4618
rect 3264 4584 3299 4618
rect 3333 4584 3368 4618
rect 3402 4584 3437 4618
rect 3471 4584 3506 4618
rect 3540 4584 3575 4618
rect 3609 4584 3644 4618
rect 3678 4584 3713 4618
rect 3747 4584 3782 4618
rect 5924 4627 5948 4754
rect 5924 4612 6118 4627
rect 5924 4584 5980 4612
rect 5948 4548 5980 4584
rect 6086 4582 6118 4612
rect 370 4355 5712 4398
rect 370 4321 470 4355
rect 504 4321 539 4355
rect 573 4321 608 4355
rect 642 4321 677 4355
rect 711 4321 746 4355
rect 780 4321 815 4355
rect 849 4321 884 4355
rect 918 4321 953 4355
rect 987 4321 1022 4355
rect 1056 4321 1091 4355
rect 1125 4321 1160 4355
rect 1194 4321 1229 4355
rect 1263 4321 1298 4355
rect 1332 4321 1367 4355
rect 1401 4321 1436 4355
rect 1470 4321 1505 4355
rect 1539 4321 1574 4355
rect 1608 4321 1643 4355
rect 1677 4321 1712 4355
rect 1746 4321 1781 4355
rect 1815 4321 1850 4355
rect 1884 4321 1919 4355
rect 1953 4321 1988 4355
rect 2022 4321 2057 4355
rect 2091 4321 2126 4355
rect 2160 4321 2195 4355
rect 2229 4321 2264 4355
rect 2298 4321 2333 4355
rect 2367 4321 2402 4355
rect 2436 4321 2471 4355
rect 370 4288 2471 4321
rect 5633 4288 5712 4355
rect 370 4254 382 4288
rect 416 4254 455 4288
rect 489 4287 528 4288
rect 562 4287 601 4288
rect 635 4287 674 4288
rect 708 4287 747 4288
rect 781 4287 820 4288
rect 854 4287 893 4288
rect 927 4287 966 4288
rect 1000 4287 1039 4288
rect 1073 4287 1112 4288
rect 1146 4287 1185 4288
rect 1219 4287 1258 4288
rect 1292 4287 1331 4288
rect 1365 4287 1404 4288
rect 1438 4287 1477 4288
rect 1511 4287 1550 4288
rect 1584 4287 1623 4288
rect 1657 4287 1696 4288
rect 1730 4287 1769 4288
rect 1803 4287 1842 4288
rect 1876 4287 1915 4288
rect 1949 4287 1988 4288
rect 2022 4287 2061 4288
rect 2095 4287 2134 4288
rect 2168 4287 2207 4288
rect 2241 4287 2280 4288
rect 2314 4287 2353 4288
rect 2387 4287 2426 4288
rect 504 4254 528 4287
rect 573 4254 601 4287
rect 642 4254 674 4287
rect 370 4253 470 4254
rect 504 4253 539 4254
rect 573 4253 608 4254
rect 642 4253 677 4254
rect 711 4253 746 4287
rect 781 4254 815 4287
rect 854 4254 884 4287
rect 927 4254 953 4287
rect 1000 4254 1022 4287
rect 1073 4254 1091 4287
rect 1146 4254 1160 4287
rect 1219 4254 1229 4287
rect 1292 4254 1298 4287
rect 1365 4254 1367 4287
rect 780 4253 815 4254
rect 849 4253 884 4254
rect 918 4253 953 4254
rect 987 4253 1022 4254
rect 1056 4253 1091 4254
rect 1125 4253 1160 4254
rect 1194 4253 1229 4254
rect 1263 4253 1298 4254
rect 1332 4253 1367 4254
rect 1401 4254 1404 4287
rect 1470 4254 1477 4287
rect 1539 4254 1550 4287
rect 1608 4254 1623 4287
rect 1677 4254 1696 4287
rect 1746 4254 1769 4287
rect 1815 4254 1842 4287
rect 1884 4254 1915 4287
rect 1401 4253 1436 4254
rect 1470 4253 1505 4254
rect 1539 4253 1574 4254
rect 1608 4253 1643 4254
rect 1677 4253 1712 4254
rect 1746 4253 1781 4254
rect 1815 4253 1850 4254
rect 1884 4253 1919 4254
rect 1953 4253 1988 4287
rect 2022 4253 2057 4287
rect 2095 4254 2126 4287
rect 2168 4254 2195 4287
rect 2241 4254 2264 4287
rect 2314 4254 2333 4287
rect 2387 4254 2402 4287
rect 2091 4253 2126 4254
rect 2160 4253 2195 4254
rect 2229 4253 2264 4254
rect 2298 4253 2333 4254
rect 2367 4253 2402 4254
rect 370 4219 2426 4253
rect 370 4216 470 4219
rect 504 4216 539 4219
rect 573 4216 608 4219
rect 642 4216 677 4219
rect 370 4182 382 4216
rect 416 4182 455 4216
rect 504 4185 528 4216
rect 573 4185 601 4216
rect 642 4185 674 4216
rect 711 4185 746 4219
rect 780 4216 815 4219
rect 849 4216 884 4219
rect 918 4216 953 4219
rect 987 4216 1022 4219
rect 1056 4216 1091 4219
rect 1125 4216 1160 4219
rect 1194 4216 1229 4219
rect 1263 4216 1298 4219
rect 1332 4216 1367 4219
rect 781 4185 815 4216
rect 854 4185 884 4216
rect 927 4185 953 4216
rect 1000 4185 1022 4216
rect 1073 4185 1091 4216
rect 1146 4185 1160 4216
rect 1219 4185 1229 4216
rect 1292 4185 1298 4216
rect 1365 4185 1367 4216
rect 1401 4216 1436 4219
rect 1470 4216 1505 4219
rect 1539 4216 1574 4219
rect 1608 4216 1643 4219
rect 1677 4216 1712 4219
rect 1746 4216 1781 4219
rect 1815 4216 1850 4219
rect 1884 4216 1919 4219
rect 1401 4185 1404 4216
rect 1470 4185 1477 4216
rect 1539 4185 1550 4216
rect 1608 4185 1623 4216
rect 1677 4185 1696 4216
rect 1746 4185 1769 4216
rect 1815 4185 1842 4216
rect 1884 4185 1915 4216
rect 1953 4185 1988 4219
rect 2022 4185 2057 4219
rect 2091 4216 2126 4219
rect 2160 4216 2195 4219
rect 2229 4216 2264 4219
rect 2298 4216 2333 4219
rect 2367 4216 2402 4219
rect 2095 4185 2126 4216
rect 2168 4185 2195 4216
rect 2241 4185 2264 4216
rect 2314 4185 2333 4216
rect 2387 4185 2402 4216
rect 489 4182 528 4185
rect 562 4182 601 4185
rect 635 4182 674 4185
rect 708 4182 747 4185
rect 781 4182 820 4185
rect 854 4182 893 4185
rect 927 4182 966 4185
rect 1000 4182 1039 4185
rect 1073 4182 1112 4185
rect 1146 4182 1185 4185
rect 1219 4182 1258 4185
rect 1292 4182 1331 4185
rect 1365 4182 1404 4185
rect 1438 4182 1477 4185
rect 1511 4182 1550 4185
rect 1584 4182 1623 4185
rect 1657 4182 1696 4185
rect 1730 4182 1769 4185
rect 1803 4182 1842 4185
rect 1876 4182 1915 4185
rect 1949 4182 1988 4185
rect 2022 4182 2061 4185
rect 2095 4182 2134 4185
rect 2168 4182 2207 4185
rect 2241 4182 2280 4185
rect 2314 4182 2353 4185
rect 2387 4182 2426 4185
rect 370 4151 2426 4182
rect 370 4144 470 4151
rect 504 4144 539 4151
rect 573 4144 608 4151
rect 642 4144 677 4151
rect 370 4110 382 4144
rect 416 4110 455 4144
rect 504 4117 528 4144
rect 573 4117 601 4144
rect 642 4117 674 4144
rect 711 4117 746 4151
rect 780 4144 815 4151
rect 849 4144 884 4151
rect 918 4144 953 4151
rect 987 4144 1022 4151
rect 1056 4144 1091 4151
rect 1125 4144 1160 4151
rect 1194 4144 1229 4151
rect 1263 4144 1298 4151
rect 1332 4144 1367 4151
rect 781 4117 815 4144
rect 854 4117 884 4144
rect 927 4117 953 4144
rect 1000 4117 1022 4144
rect 1073 4117 1091 4144
rect 1146 4117 1160 4144
rect 1219 4117 1229 4144
rect 1292 4117 1298 4144
rect 1365 4117 1367 4144
rect 1401 4144 1436 4151
rect 1470 4144 1505 4151
rect 1539 4144 1574 4151
rect 1608 4144 1643 4151
rect 1677 4144 1712 4151
rect 1746 4144 1781 4151
rect 1815 4144 1850 4151
rect 1884 4144 1919 4151
rect 1401 4117 1404 4144
rect 1470 4117 1477 4144
rect 1539 4117 1550 4144
rect 1608 4117 1623 4144
rect 1677 4117 1696 4144
rect 1746 4117 1769 4144
rect 1815 4117 1842 4144
rect 1884 4117 1915 4144
rect 1953 4117 1988 4151
rect 2022 4117 2057 4151
rect 2091 4144 2126 4151
rect 2160 4144 2195 4151
rect 2229 4144 2264 4151
rect 2298 4144 2333 4151
rect 2367 4144 2402 4151
rect 2095 4117 2126 4144
rect 2168 4117 2195 4144
rect 2241 4117 2264 4144
rect 2314 4117 2333 4144
rect 2387 4117 2402 4144
rect 489 4110 528 4117
rect 562 4110 601 4117
rect 635 4110 674 4117
rect 708 4110 747 4117
rect 781 4110 820 4117
rect 854 4110 893 4117
rect 927 4110 966 4117
rect 1000 4110 1039 4117
rect 1073 4110 1112 4117
rect 1146 4110 1185 4117
rect 1219 4110 1258 4117
rect 1292 4110 1331 4117
rect 1365 4110 1404 4117
rect 1438 4110 1477 4117
rect 1511 4110 1550 4117
rect 1584 4110 1623 4117
rect 1657 4110 1696 4117
rect 1730 4110 1769 4117
rect 1803 4110 1842 4117
rect 1876 4110 1915 4117
rect 1949 4110 1988 4117
rect 2022 4110 2061 4117
rect 2095 4110 2134 4117
rect 2168 4110 2207 4117
rect 2241 4110 2280 4117
rect 2314 4110 2353 4117
rect 2387 4110 2426 4117
rect 370 4072 2426 4110
rect 370 4038 382 4072
rect 416 4038 455 4072
rect 489 4038 528 4072
rect 562 4038 601 4072
rect 635 4038 674 4072
rect 708 4038 747 4072
rect 781 4038 820 4072
rect 854 4038 893 4072
rect 927 4038 966 4072
rect 1000 4038 1039 4072
rect 1073 4038 1112 4072
rect 1146 4038 1185 4072
rect 1219 4038 1258 4072
rect 1292 4038 1331 4072
rect 1365 4038 1404 4072
rect 1438 4038 1477 4072
rect 1511 4038 1550 4072
rect 1584 4038 1623 4072
rect 1657 4038 1696 4072
rect 1730 4038 1769 4072
rect 1803 4038 1842 4072
rect 1876 4038 1915 4072
rect 1949 4038 1988 4072
rect 2022 4038 2061 4072
rect 2095 4038 2134 4072
rect 2168 4038 2207 4072
rect 2241 4038 2280 4072
rect 2314 4038 2353 4072
rect 2387 4038 2426 4072
rect 5700 4038 5712 4288
rect 370 4032 2426 4038
rect 3334 4032 5125 4038
rect 5231 4032 5712 4038
rect 370 3998 472 4032
rect 404 3964 472 3998
rect 370 3930 438 3964
rect 370 3929 506 3930
rect 404 3895 506 3929
rect 370 3894 506 3895
rect 5402 4000 5437 4032
rect 5422 3998 5437 4000
rect 5471 4000 5506 4032
rect 5471 3998 5484 4000
rect 5540 3998 5575 4032
rect 5609 3998 5644 4032
rect 5678 3998 5712 4032
rect 5368 3966 5388 3998
rect 5422 3966 5484 3998
rect 5518 3966 5712 3998
rect 5368 3964 5712 3966
rect 5368 3930 5403 3964
rect 5437 3930 5472 3964
rect 5506 3930 5541 3964
rect 5575 3930 5610 3964
rect 5644 3930 5712 3964
rect 5300 3928 5610 3930
rect 5315 3896 5365 3928
rect 5399 3896 5450 3928
rect 5484 3896 5610 3928
rect 5315 3894 5335 3896
rect 5399 3894 5404 3896
rect 370 3860 438 3894
rect 472 3862 506 3894
rect 5300 3862 5335 3894
rect 5369 3862 5404 3894
rect 5438 3894 5450 3896
rect 5438 3862 5473 3894
rect 5507 3890 5542 3896
rect 5507 3862 5522 3890
rect 472 3860 526 3862
rect 404 3855 526 3860
rect 560 3855 632 3862
rect 404 3850 598 3855
rect 488 3826 598 3850
rect 370 3791 382 3826
rect 488 3792 506 3826
rect 540 3821 598 3826
rect 540 3816 632 3821
rect 488 3782 526 3792
rect 560 3782 632 3816
rect 370 3722 382 3757
rect 488 3756 598 3782
rect 488 3724 506 3756
rect 540 3748 598 3756
rect 721 3806 763 3818
rect 797 3806 839 3818
rect 873 3806 915 3818
rect 949 3806 991 3818
rect 1025 3806 1067 3818
rect 1101 3806 1144 3818
rect 1178 3806 1221 3818
rect 737 3784 763 3806
rect 808 3784 839 3806
rect 879 3784 915 3806
rect 687 3772 703 3784
rect 737 3772 774 3784
rect 808 3772 845 3784
rect 879 3772 917 3784
rect 951 3772 989 3806
rect 1025 3784 1061 3806
rect 1101 3784 1133 3806
rect 1178 3784 1205 3806
rect 1023 3772 1061 3784
rect 1095 3772 1133 3784
rect 1167 3772 1205 3784
rect 1239 3772 1255 3784
rect 540 3743 632 3748
rect 488 3709 526 3724
rect 560 3709 632 3743
rect 1289 3738 1481 3862
rect 1549 3806 1591 3818
rect 1625 3806 1667 3818
rect 1701 3806 1743 3818
rect 1777 3806 1819 3818
rect 1853 3806 1895 3818
rect 1929 3806 1972 3818
rect 2006 3806 2049 3818
rect 1565 3784 1591 3806
rect 1636 3784 1667 3806
rect 1707 3784 1743 3806
rect 1515 3772 1531 3784
rect 1565 3772 1602 3784
rect 1636 3772 1673 3784
rect 1707 3772 1745 3784
rect 1779 3772 1817 3806
rect 1853 3784 1889 3806
rect 1929 3784 1961 3806
rect 2006 3784 2033 3806
rect 1851 3772 1889 3784
rect 1923 3772 1961 3784
rect 1995 3772 2033 3784
rect 2067 3772 2083 3784
rect 2117 3738 2309 3862
rect 2377 3806 2419 3818
rect 2453 3806 2495 3818
rect 2529 3806 2571 3818
rect 2605 3806 2647 3818
rect 2681 3806 2723 3818
rect 2757 3806 2800 3818
rect 2834 3806 2877 3818
rect 2393 3784 2419 3806
rect 2464 3784 2495 3806
rect 2535 3784 2571 3806
rect 2343 3772 2359 3784
rect 2393 3772 2430 3784
rect 2464 3772 2501 3784
rect 2535 3772 2573 3784
rect 2607 3772 2645 3806
rect 2681 3784 2717 3806
rect 2757 3784 2789 3806
rect 2834 3784 2861 3806
rect 2679 3772 2717 3784
rect 2751 3772 2789 3784
rect 2823 3772 2861 3784
rect 2895 3772 2911 3784
rect 370 3653 382 3688
rect 488 3675 598 3709
rect 488 3670 632 3675
rect 488 3636 526 3670
rect 560 3636 632 3670
rect 370 3584 382 3619
rect 488 3602 598 3636
rect 488 3597 632 3602
rect 488 3563 526 3597
rect 560 3563 632 3597
rect 370 3515 382 3550
rect 488 3529 598 3563
rect 488 3524 632 3529
rect 488 3490 526 3524
rect 560 3490 632 3524
rect 370 3446 382 3481
rect 488 3456 598 3490
rect 488 3451 632 3456
rect 488 3417 526 3451
rect 560 3417 632 3451
rect 370 3377 382 3412
rect 488 3383 598 3417
rect 488 3378 632 3383
rect 488 3344 526 3378
rect 560 3344 632 3378
rect 370 3308 382 3343
rect 488 3310 598 3344
rect 488 3305 632 3310
rect 370 3239 382 3274
rect 488 3271 526 3305
rect 560 3271 632 3305
rect 488 3237 598 3271
rect 488 3232 632 3237
rect 370 3170 382 3205
rect 488 3198 526 3232
rect 560 3198 632 3232
rect 488 3164 598 3198
rect 488 3159 632 3164
rect 370 3101 382 3136
rect 488 3125 526 3159
rect 560 3125 632 3159
rect 488 3091 598 3125
rect 488 3086 632 3091
rect 370 3032 382 3067
rect 488 3052 526 3086
rect 560 3052 632 3086
rect 488 3018 598 3052
rect 488 3013 632 3018
rect 370 2963 382 2998
rect 488 2979 526 3013
rect 560 2979 632 3013
rect 488 2952 598 2979
rect 404 2950 438 2952
rect 472 2950 598 2952
rect 404 2945 598 2950
rect 404 2940 632 2945
rect 404 2929 526 2940
rect 370 2914 526 2929
rect 370 2913 438 2914
rect 472 2913 526 2914
rect 370 2894 382 2913
rect 416 2880 438 2913
rect 488 2906 526 2913
rect 560 2906 632 2940
rect 416 2879 454 2880
rect 488 2879 598 2906
rect 404 2872 598 2879
rect 404 2867 632 2872
rect 404 2860 526 2867
rect 370 2844 526 2860
rect 370 2840 438 2844
rect 472 2840 526 2844
rect 370 2825 382 2840
rect 416 2810 438 2840
rect 488 2833 526 2840
rect 560 2833 632 2867
rect 416 2806 454 2810
rect 488 2806 598 2833
rect 404 2799 598 2806
rect 404 2794 632 2799
rect 404 2791 526 2794
rect 370 2774 526 2791
rect 370 2767 438 2774
rect 472 2767 526 2774
rect 370 2756 382 2767
rect 416 2740 438 2767
rect 488 2760 526 2767
rect 560 2760 632 2794
rect 416 2733 454 2740
rect 488 2733 598 2760
rect 404 2726 598 2733
rect 404 2722 632 2726
rect 370 2721 632 2722
rect 370 2704 526 2721
rect 370 2694 438 2704
rect 472 2694 526 2704
rect 370 2687 382 2694
rect 416 2670 438 2694
rect 488 2687 526 2694
rect 560 2687 632 2721
rect 416 2660 454 2670
rect 488 2660 598 2687
rect 404 2653 598 2660
rect 370 2648 632 2653
rect 370 2634 526 2648
rect 370 2621 438 2634
rect 472 2621 526 2634
rect 370 2618 382 2621
rect 416 2600 438 2621
rect 488 2614 526 2621
rect 560 2614 632 2648
rect 416 2587 454 2600
rect 488 2587 598 2614
rect 404 2584 598 2587
rect 370 2580 598 2584
rect 370 2575 632 2580
rect 370 2564 526 2575
rect 370 2549 438 2564
rect 404 2548 438 2549
rect 472 2548 526 2564
rect 416 2530 438 2548
rect 488 2541 526 2548
rect 560 2541 632 2575
rect 370 2514 382 2515
rect 416 2514 454 2530
rect 488 2514 598 2541
rect 370 2507 598 2514
rect 370 2502 632 2507
rect 370 2494 526 2502
rect 370 2480 438 2494
rect 404 2475 438 2480
rect 472 2475 526 2494
rect 416 2460 438 2475
rect 488 2468 526 2475
rect 560 2468 632 2502
rect 370 2441 382 2446
rect 416 2441 454 2460
rect 488 2441 598 2468
rect 370 2434 598 2441
rect 370 2429 632 2434
rect 370 2424 526 2429
rect 370 2411 438 2424
rect 404 2402 438 2411
rect 472 2402 526 2424
rect 416 2390 438 2402
rect 488 2395 526 2402
rect 560 2395 632 2429
rect 370 2368 382 2377
rect 416 2368 454 2390
rect 488 2368 598 2395
rect 370 2361 598 2368
rect 370 2356 632 2361
rect 370 2354 526 2356
rect 370 2342 438 2354
rect 404 2329 438 2342
rect 472 2329 526 2354
rect 416 2320 438 2329
rect 488 2322 526 2329
rect 560 2322 632 2356
rect 370 2295 382 2308
rect 416 2295 454 2320
rect 488 2295 598 2322
rect 370 2288 598 2295
rect 370 2284 632 2288
rect 370 2273 438 2284
rect 404 2256 438 2273
rect 472 2283 632 2284
rect 472 2256 526 2283
rect 416 2250 438 2256
rect 370 2222 382 2239
rect 416 2222 454 2250
rect 488 2249 526 2256
rect 560 2249 632 2283
rect 1289 3728 1297 3738
rect 954 3665 988 3704
rect 954 3592 988 3631
rect 954 3520 988 3558
rect 954 3448 988 3486
rect 954 3376 988 3414
rect 954 3304 988 3342
rect 954 3232 988 3270
rect 954 3160 988 3198
rect 954 3088 988 3126
rect 954 3016 988 3054
rect 954 2944 988 2982
rect 954 2872 988 2910
rect 954 2800 988 2838
rect 954 2728 988 2766
rect 954 2656 988 2694
rect 954 2584 988 2622
rect 954 2512 988 2550
rect 954 2440 988 2478
rect 954 2368 988 2406
rect 954 2296 988 2334
rect 1331 3704 1369 3738
rect 1403 3704 1441 3738
rect 1475 3728 1481 3738
rect 1297 3665 1475 3704
rect 1331 3631 1369 3665
rect 1403 3631 1441 3665
rect 1297 3592 1475 3631
rect 2117 3728 2124 3738
rect 1782 3665 1816 3704
rect 1782 3592 1816 3631
rect 1782 3520 1816 3558
rect 1782 3448 1816 3486
rect 1782 3376 1816 3414
rect 1782 3304 1816 3342
rect 1782 3232 1816 3270
rect 1782 3160 1816 3198
rect 1782 3088 1816 3126
rect 1782 3016 1816 3054
rect 1782 2944 1816 2982
rect 1782 2872 1816 2910
rect 1782 2800 1816 2838
rect 1782 2728 1816 2766
rect 1782 2656 1816 2694
rect 1782 2584 1816 2622
rect 1782 2512 1816 2550
rect 1782 2440 1816 2478
rect 1782 2368 1816 2406
rect 1782 2296 1816 2334
rect 2158 3704 2196 3738
rect 2230 3704 2268 3738
rect 2302 3728 2309 3738
rect 2124 3665 2302 3704
rect 2158 3631 2196 3665
rect 2230 3631 2268 3665
rect 2124 3592 2302 3631
rect 2610 3665 2644 3704
rect 2610 3592 2644 3631
rect 2610 3520 2644 3558
rect 2610 3448 2644 3486
rect 2610 3376 2644 3414
rect 2610 3304 2644 3342
rect 2610 3232 2644 3270
rect 2610 3160 2644 3198
rect 2610 3088 2644 3126
rect 2610 3016 2644 3054
rect 2610 2944 2644 2982
rect 2610 2872 2644 2910
rect 2610 2800 2644 2838
rect 2610 2728 2644 2766
rect 2610 2656 2644 2694
rect 2610 2584 2644 2622
rect 2610 2512 2644 2550
rect 2610 2440 2644 2478
rect 2610 2368 2644 2406
rect 2610 2296 2644 2334
rect 488 2222 598 2249
rect 370 2215 598 2222
rect 370 2214 632 2215
rect 370 2204 438 2214
rect 404 2183 438 2204
rect 472 2210 632 2214
rect 472 2183 526 2210
rect 416 2180 438 2183
rect 370 2149 382 2170
rect 416 2149 454 2180
rect 488 2176 526 2183
rect 560 2176 632 2210
rect 488 2149 598 2176
rect 370 2144 598 2149
rect 370 2135 438 2144
rect 404 2110 438 2135
rect 472 2142 598 2144
rect 472 2137 632 2142
rect 472 2110 526 2137
rect 370 2076 382 2101
rect 416 2076 454 2110
rect 488 2103 526 2110
rect 560 2103 632 2137
rect 488 2076 598 2103
rect 370 2075 598 2076
rect 370 2066 438 2075
rect 404 2041 438 2066
rect 472 2069 598 2075
rect 472 2064 632 2069
rect 472 2041 526 2064
rect 404 2037 526 2041
rect 370 2003 382 2032
rect 416 2006 454 2037
rect 488 2030 526 2037
rect 560 2030 632 2064
rect 416 2003 438 2006
rect 488 2003 598 2030
rect 370 1997 438 2003
rect 404 1972 438 1997
rect 472 1996 598 2003
rect 472 1991 632 1996
rect 472 1972 526 1991
rect 404 1964 526 1972
rect 370 1930 382 1963
rect 416 1937 454 1964
rect 488 1957 526 1964
rect 560 1957 632 1991
rect 416 1930 438 1937
rect 488 1930 598 1957
rect 370 1929 438 1930
rect 404 1903 438 1929
rect 472 1923 598 1930
rect 472 1918 632 1923
rect 472 1903 526 1918
rect 404 1895 526 1903
rect 370 1891 526 1895
rect 370 1861 382 1891
rect 416 1868 454 1891
rect 488 1884 526 1891
rect 560 1884 632 1918
rect 416 1857 438 1868
rect 488 1857 598 1884
rect 404 1834 438 1857
rect 472 1850 598 1857
rect 472 1845 632 1850
rect 472 1834 526 1845
rect 404 1827 526 1834
rect 370 1818 526 1827
rect 370 1793 382 1818
rect 416 1799 454 1818
rect 488 1811 526 1818
rect 560 1811 632 1845
rect 416 1784 438 1799
rect 488 1784 598 1811
rect 404 1765 438 1784
rect 472 1777 598 1784
rect 472 1772 632 1777
rect 472 1765 526 1772
rect 404 1759 526 1765
rect 370 1745 526 1759
rect 370 1725 382 1745
rect 416 1730 454 1745
rect 488 1738 526 1745
rect 560 1738 632 1772
rect 416 1711 438 1730
rect 488 1711 598 1738
rect 404 1696 438 1711
rect 472 1704 598 1711
rect 472 1699 632 1704
rect 472 1696 526 1699
rect 404 1691 526 1696
rect 370 1672 526 1691
rect 370 1657 382 1672
rect 416 1661 454 1672
rect 488 1665 526 1672
rect 560 1665 632 1699
rect 416 1638 438 1661
rect 488 1638 598 1665
rect 404 1627 438 1638
rect 472 1631 598 1638
rect 472 1627 632 1631
rect 404 1626 632 1627
rect 404 1623 526 1626
rect 370 1599 526 1623
rect 370 1589 382 1599
rect 416 1592 454 1599
rect 488 1592 526 1599
rect 560 1592 632 1626
rect 416 1565 438 1592
rect 488 1565 598 1592
rect 404 1558 438 1565
rect 472 1558 598 1565
rect 404 1555 632 1558
rect 370 1553 632 1555
rect 370 1526 526 1553
rect 370 1521 382 1526
rect 416 1523 454 1526
rect 416 1492 438 1523
rect 488 1519 526 1526
rect 560 1519 632 1553
rect 488 1492 598 1519
rect 404 1489 438 1492
rect 472 1489 598 1492
rect 404 1487 598 1489
rect 370 1485 598 1487
rect 370 1480 632 1485
rect 370 1454 526 1480
rect 370 1453 438 1454
rect 472 1453 526 1454
rect 416 1420 438 1453
rect 488 1446 526 1453
rect 560 1446 632 1480
rect 416 1419 454 1420
rect 488 1419 598 1446
rect 370 1412 598 1419
rect 370 1407 632 1412
rect 370 1385 526 1407
rect 404 1380 438 1385
rect 472 1380 526 1385
rect 416 1351 438 1380
rect 488 1373 526 1380
rect 560 1373 632 1407
rect 370 1346 382 1351
rect 416 1346 454 1351
rect 488 1346 598 1373
rect 370 1339 598 1346
rect 370 1334 632 1339
rect 370 1307 526 1334
rect 370 1283 382 1307
rect 416 1283 454 1307
rect 488 1300 526 1307
rect 560 1300 632 1334
rect 416 1273 438 1283
rect 488 1273 598 1300
rect 404 1249 438 1273
rect 472 1266 598 1273
rect 472 1261 632 1266
rect 472 1249 526 1261
rect 370 1234 526 1249
rect 370 1212 382 1234
rect 416 1214 454 1234
rect 488 1227 526 1234
rect 560 1227 632 1261
rect 488 1214 598 1227
rect 416 1200 438 1214
rect 404 1178 438 1200
rect 506 1193 598 1214
rect 506 1188 632 1193
rect 506 1180 526 1188
rect 370 1161 438 1178
rect 370 1141 382 1161
rect 416 1127 438 1161
rect 560 1154 632 1188
rect 540 1146 598 1154
rect 404 1107 438 1127
rect 506 1120 598 1146
rect 506 1115 632 1120
rect 506 1112 526 1115
rect 370 1088 438 1107
rect 370 1070 382 1088
rect 416 1054 438 1088
rect 560 1081 632 1115
rect 540 1078 598 1081
rect 404 1036 438 1054
rect 506 1047 598 1078
rect 506 1044 632 1047
rect 540 1042 632 1044
rect 370 1015 438 1036
rect 370 999 382 1015
rect 416 981 438 1015
rect 506 1008 526 1010
rect 560 1008 632 1042
rect 404 965 438 981
rect 506 976 598 1008
rect 540 974 598 976
rect 540 969 632 974
rect 370 942 438 965
rect 370 928 382 942
rect 416 908 438 942
rect 506 935 526 942
rect 560 935 632 969
rect 506 908 598 935
rect 404 894 438 908
rect 540 901 598 908
rect 540 896 632 901
rect 370 869 438 894
rect 370 857 382 869
rect 416 835 438 869
rect 506 862 526 874
rect 560 862 632 896
rect 506 840 598 862
rect 404 823 438 835
rect 540 828 598 840
rect 540 824 632 828
rect 370 796 438 823
rect 370 786 382 796
rect 416 762 438 796
rect 506 790 526 806
rect 560 790 632 824
rect 506 789 632 790
rect 506 772 598 789
rect 404 752 438 762
rect 540 755 598 772
rect 540 752 632 755
rect 370 723 438 752
rect 506 724 526 738
rect 370 715 382 723
rect 416 689 438 723
rect 560 718 632 752
rect 798 2137 832 2176
rect 798 2064 832 2103
rect 798 1992 832 2030
rect 798 1920 832 1958
rect 798 1848 832 1886
rect 798 1776 832 1814
rect 798 1704 832 1742
rect 798 1632 832 1670
rect 798 1560 832 1598
rect 798 1488 832 1526
rect 798 1416 832 1454
rect 798 1344 832 1382
rect 798 1272 832 1310
rect 798 1200 832 1238
rect 798 1128 832 1166
rect 798 1056 832 1094
rect 798 984 832 1022
rect 798 912 832 950
rect 798 840 832 878
rect 798 768 832 806
rect 1110 2137 1144 2176
rect 1110 2064 1144 2103
rect 1110 1992 1144 2030
rect 1110 1920 1144 1958
rect 1110 1848 1144 1886
rect 1110 1776 1144 1814
rect 1110 1704 1144 1742
rect 1110 1632 1144 1670
rect 1110 1560 1144 1598
rect 1110 1488 1144 1526
rect 1110 1416 1144 1454
rect 1110 1344 1144 1382
rect 1110 1272 1144 1310
rect 1110 1200 1144 1238
rect 1110 1128 1144 1166
rect 1110 1056 1144 1094
rect 1110 984 1144 1022
rect 1110 912 1144 950
rect 1110 840 1144 878
rect 1110 768 1144 806
rect 1626 2137 1660 2176
rect 1626 2064 1660 2103
rect 1626 1992 1660 2030
rect 1626 1920 1660 1958
rect 1626 1848 1660 1886
rect 1626 1776 1660 1814
rect 1626 1704 1660 1742
rect 1626 1632 1660 1670
rect 1626 1560 1660 1598
rect 1626 1488 1660 1526
rect 1626 1416 1660 1454
rect 1626 1344 1660 1382
rect 1626 1272 1660 1310
rect 1626 1200 1660 1238
rect 1626 1128 1660 1166
rect 1626 1056 1660 1094
rect 1626 984 1660 1022
rect 1626 912 1660 950
rect 1626 840 1660 878
rect 1626 768 1660 806
rect 540 716 632 718
rect 404 681 438 689
rect 370 650 438 681
rect 540 682 598 716
rect 540 680 632 682
rect 370 644 382 650
rect 416 616 438 650
rect 560 646 632 680
rect 540 643 632 646
rect 404 610 438 616
rect 370 573 438 610
rect 540 609 598 643
rect 687 642 688 676
rect 737 642 764 676
rect 808 642 840 676
rect 879 642 916 676
rect 951 642 989 676
rect 1026 642 1061 676
rect 1102 642 1133 676
rect 1178 642 1205 676
rect 540 608 632 609
rect 560 602 632 608
rect 1289 602 1481 738
rect 1938 2137 1972 2176
rect 1938 2064 1972 2103
rect 1938 1992 1972 2030
rect 1938 1920 1972 1958
rect 1938 1848 1972 1886
rect 1938 1776 1972 1814
rect 1938 1704 1972 1742
rect 1938 1632 1972 1670
rect 1938 1560 1972 1598
rect 1938 1488 1972 1526
rect 1938 1416 1972 1454
rect 1938 1344 1972 1382
rect 1938 1272 1972 1310
rect 1938 1200 1972 1238
rect 1938 1128 1972 1166
rect 1938 1056 1972 1094
rect 1938 984 1972 1022
rect 1938 912 1972 950
rect 1938 840 1972 878
rect 1938 768 1972 806
rect 2454 2137 2488 2176
rect 2454 2064 2488 2103
rect 2454 1992 2488 2030
rect 2454 1920 2488 1958
rect 2454 1848 2488 1886
rect 2454 1776 2488 1814
rect 2454 1704 2488 1742
rect 2454 1632 2488 1670
rect 2454 1560 2488 1598
rect 2454 1488 2488 1526
rect 2454 1416 2488 1454
rect 2454 1344 2488 1382
rect 2454 1272 2488 1310
rect 2454 1200 2488 1238
rect 2454 1128 2488 1166
rect 2454 1056 2488 1094
rect 2454 984 2488 1022
rect 2454 912 2488 950
rect 2454 840 2488 878
rect 2454 768 2488 806
rect 1515 642 1516 676
rect 1565 642 1592 676
rect 1636 642 1668 676
rect 1707 642 1744 676
rect 1779 642 1817 676
rect 1854 642 1889 676
rect 1930 642 1961 676
rect 2006 642 2033 676
rect 2117 602 2309 738
rect 2766 2137 2800 2176
rect 2766 2064 2800 2103
rect 2766 1992 2800 2030
rect 2766 1920 2800 1958
rect 2766 1848 2800 1886
rect 2766 1776 2800 1814
rect 2766 1704 2800 1742
rect 2766 1632 2800 1670
rect 2766 1560 2800 1598
rect 2766 1488 2800 1526
rect 2766 1416 2800 1454
rect 2766 1344 2800 1382
rect 2766 1272 2800 1310
rect 2766 1200 2800 1238
rect 2766 1128 2800 1166
rect 2766 1056 2800 1094
rect 2766 984 2800 1022
rect 2766 912 2800 950
rect 2766 840 2800 878
rect 2766 768 2800 806
rect 2834 676 2888 3772
rect 2945 3738 3137 3862
rect 3205 3806 3247 3818
rect 3281 3806 3323 3818
rect 3357 3806 3399 3818
rect 3433 3806 3475 3818
rect 3509 3806 3551 3818
rect 3585 3806 3628 3818
rect 3662 3806 3705 3818
rect 3221 3784 3247 3806
rect 3292 3784 3323 3806
rect 3363 3784 3399 3806
rect 3171 3772 3187 3784
rect 3221 3772 3258 3784
rect 3292 3772 3329 3784
rect 3363 3772 3401 3784
rect 3435 3772 3473 3806
rect 3509 3784 3545 3806
rect 3585 3784 3617 3806
rect 3662 3784 3689 3806
rect 3507 3772 3545 3784
rect 3579 3772 3617 3784
rect 3651 3772 3689 3784
rect 3723 3772 3739 3784
rect 2945 3728 2952 3738
rect 2986 3704 3024 3738
rect 3058 3704 3096 3738
rect 3130 3728 3137 3738
rect 2952 3665 3130 3704
rect 2986 3631 3024 3665
rect 3058 3631 3096 3665
rect 2952 3592 3130 3631
rect 2343 642 2344 676
rect 2393 642 2420 676
rect 2464 642 2496 676
rect 2535 642 2572 676
rect 2607 642 2645 676
rect 2682 642 2717 676
rect 2758 642 2789 676
rect 2834 642 2861 676
rect 2945 602 3137 738
rect 3194 676 3248 3772
rect 3773 3738 3964 3862
rect 4032 3806 4074 3818
rect 4108 3806 4150 3818
rect 4184 3806 4226 3818
rect 4260 3806 4302 3818
rect 4336 3806 4379 3818
rect 4413 3806 4456 3818
rect 4490 3806 4533 3818
rect 4048 3784 4074 3806
rect 4119 3784 4150 3806
rect 4191 3784 4226 3806
rect 3998 3772 4014 3784
rect 4048 3772 4085 3784
rect 4119 3772 4157 3784
rect 4191 3772 4229 3784
rect 4263 3772 4301 3806
rect 4336 3784 4373 3806
rect 4413 3784 4445 3806
rect 4490 3784 4517 3806
rect 4335 3772 4373 3784
rect 4407 3772 4445 3784
rect 4479 3772 4517 3784
rect 4551 3772 4567 3784
rect 4601 3738 4793 3862
rect 5450 3856 5522 3862
rect 5450 3855 5542 3856
rect 5484 3850 5542 3855
rect 5484 3821 5522 3850
rect 4861 3806 4903 3818
rect 4937 3806 4979 3818
rect 5013 3806 5055 3818
rect 5089 3806 5131 3818
rect 5165 3806 5207 3818
rect 5241 3806 5284 3818
rect 5318 3806 5361 3818
rect 4877 3784 4903 3806
rect 4948 3784 4979 3806
rect 5019 3784 5055 3806
rect 4827 3772 4843 3784
rect 4877 3772 4914 3784
rect 4948 3772 4985 3784
rect 5019 3772 5057 3784
rect 5091 3772 5129 3806
rect 5165 3784 5201 3806
rect 5241 3784 5273 3806
rect 5318 3784 5345 3806
rect 5163 3772 5201 3784
rect 5235 3772 5273 3784
rect 5307 3772 5345 3784
rect 5379 3772 5395 3784
rect 5450 3782 5522 3821
rect 5484 3748 5522 3782
rect 3773 3728 3781 3738
rect 3438 3665 3472 3704
rect 3438 3592 3472 3631
rect 3438 3520 3472 3558
rect 3438 3448 3472 3486
rect 3438 3376 3472 3414
rect 3438 3304 3472 3342
rect 3438 3232 3472 3270
rect 3438 3160 3472 3198
rect 3438 3088 3472 3126
rect 3438 3016 3472 3054
rect 3438 2944 3472 2982
rect 3438 2872 3472 2910
rect 3438 2800 3472 2838
rect 3438 2728 3472 2766
rect 3438 2656 3472 2694
rect 3438 2584 3472 2622
rect 3438 2512 3472 2550
rect 3438 2440 3472 2478
rect 3438 2368 3472 2406
rect 3438 2296 3472 2334
rect 3815 3704 3853 3738
rect 3887 3704 3925 3738
rect 3959 3728 3964 3738
rect 3781 3665 3959 3704
rect 3815 3631 3853 3665
rect 3887 3631 3925 3665
rect 3781 3592 3959 3631
rect 4601 3728 4608 3738
rect 4266 3665 4300 3704
rect 4266 3592 4300 3631
rect 4266 3520 4300 3558
rect 4266 3448 4300 3486
rect 4266 3376 4300 3414
rect 4266 3304 4300 3342
rect 4266 3232 4300 3270
rect 4266 3160 4300 3198
rect 4266 3088 4300 3126
rect 4266 3016 4300 3054
rect 4266 2944 4300 2982
rect 4266 2872 4300 2910
rect 4266 2800 4300 2838
rect 4266 2728 4300 2766
rect 4266 2656 4300 2694
rect 4266 2584 4300 2622
rect 4266 2512 4300 2550
rect 4266 2440 4300 2478
rect 4266 2368 4300 2406
rect 4266 2296 4300 2334
rect 4642 3704 4680 3738
rect 4714 3704 4752 3738
rect 4786 3728 4793 3738
rect 4608 3665 4786 3704
rect 4642 3631 4680 3665
rect 4714 3631 4752 3665
rect 4608 3592 4786 3631
rect 5094 3665 5128 3704
rect 5094 3592 5128 3631
rect 5094 3520 5128 3558
rect 5094 3448 5128 3486
rect 5094 3376 5128 3414
rect 5094 3304 5128 3342
rect 5094 3232 5128 3270
rect 5094 3160 5128 3198
rect 5094 3088 5128 3126
rect 5094 3016 5128 3054
rect 5094 2944 5128 2982
rect 5094 2872 5128 2910
rect 5094 2800 5128 2838
rect 5094 2728 5128 2766
rect 5094 2656 5128 2694
rect 5094 2584 5128 2622
rect 5094 2512 5128 2550
rect 5094 2440 5128 2478
rect 5094 2368 5128 2406
rect 5094 2296 5128 2334
rect 5450 3709 5522 3748
rect 5484 3675 5522 3709
rect 5450 3636 5522 3675
rect 5484 3602 5522 3636
rect 5450 3568 5522 3602
rect 5450 3563 5542 3568
rect 5484 3556 5542 3563
rect 5484 3529 5576 3556
rect 5450 3495 5522 3529
rect 5556 3522 5576 3529
rect 5450 3490 5542 3495
rect 5484 3488 5542 3490
rect 5484 3456 5576 3488
rect 5450 3422 5522 3456
rect 5556 3454 5576 3456
rect 5450 3420 5542 3422
rect 5450 3417 5576 3420
rect 5484 3386 5576 3417
rect 5484 3383 5542 3386
rect 5450 3349 5522 3383
rect 5556 3349 5576 3352
rect 5450 3344 5576 3349
rect 5484 3318 5576 3344
rect 5484 3310 5542 3318
rect 5450 3276 5522 3310
rect 5556 3276 5576 3284
rect 5450 3271 5576 3276
rect 5484 3250 5576 3271
rect 5484 3237 5542 3250
rect 5450 3203 5522 3237
rect 5556 3203 5576 3216
rect 5450 3198 5576 3203
rect 5484 3182 5576 3198
rect 5484 3164 5542 3182
rect 5450 3130 5522 3164
rect 5556 3130 5576 3148
rect 5450 3125 5576 3130
rect 5484 3114 5576 3125
rect 5484 3091 5542 3114
rect 5450 3057 5522 3091
rect 5556 3057 5576 3080
rect 5450 3052 5576 3057
rect 5484 3046 5576 3052
rect 5484 3018 5542 3046
rect 5450 2984 5522 3018
rect 5556 2984 5576 3012
rect 5450 2979 5576 2984
rect 5484 2978 5576 2979
rect 5484 2945 5542 2978
rect 5450 2911 5522 2945
rect 5556 2911 5576 2944
rect 5450 2910 5576 2911
rect 5450 2906 5542 2910
rect 5484 2876 5542 2906
rect 5484 2872 5576 2876
rect 5450 2838 5522 2872
rect 5556 2842 5576 2872
rect 5450 2833 5542 2838
rect 5484 2808 5542 2833
rect 5484 2799 5576 2808
rect 5450 2765 5522 2799
rect 5556 2774 5576 2799
rect 5450 2760 5542 2765
rect 5484 2740 5542 2760
rect 5484 2726 5576 2740
rect 5450 2692 5522 2726
rect 5556 2706 5576 2726
rect 5450 2687 5542 2692
rect 5484 2672 5542 2687
rect 5484 2653 5576 2672
rect 5450 2619 5522 2653
rect 5556 2638 5576 2653
rect 5556 2621 5610 2638
rect 5556 2619 5594 2621
rect 5450 2614 5594 2619
rect 5484 2587 5594 2614
rect 5484 2580 5610 2587
rect 5450 2546 5522 2580
rect 5556 2570 5610 2580
rect 5556 2548 5678 2570
rect 5556 2546 5594 2548
rect 5450 2541 5594 2546
rect 5484 2514 5594 2541
rect 5628 2535 5666 2548
rect 5644 2514 5666 2535
rect 5700 2514 5712 2536
rect 5484 2507 5610 2514
rect 5450 2473 5522 2507
rect 5556 2501 5610 2507
rect 5644 2501 5712 2514
rect 5556 2475 5678 2501
rect 5556 2473 5594 2475
rect 5450 2468 5594 2473
rect 5484 2441 5594 2468
rect 5628 2466 5666 2475
rect 5644 2441 5666 2466
rect 5700 2441 5712 2467
rect 5484 2434 5610 2441
rect 5450 2400 5522 2434
rect 5556 2432 5610 2434
rect 5644 2432 5712 2441
rect 5556 2402 5678 2432
rect 5556 2400 5594 2402
rect 5450 2395 5594 2400
rect 5628 2397 5666 2402
rect 5484 2368 5594 2395
rect 5644 2368 5666 2397
rect 5700 2368 5712 2398
rect 5484 2363 5610 2368
rect 5644 2363 5712 2368
rect 5484 2361 5678 2363
rect 5450 2327 5522 2361
rect 5556 2329 5678 2361
rect 5556 2327 5594 2329
rect 5628 2328 5666 2329
rect 5450 2322 5594 2327
rect 5484 2295 5594 2322
rect 5644 2295 5666 2328
rect 5700 2295 5712 2329
rect 5484 2294 5610 2295
rect 5644 2294 5712 2295
rect 5484 2288 5678 2294
rect 5450 2254 5522 2288
rect 5556 2260 5678 2288
rect 5556 2259 5712 2260
rect 5556 2256 5610 2259
rect 5644 2256 5712 2259
rect 5556 2254 5594 2256
rect 5450 2249 5594 2254
rect 5484 2222 5594 2249
rect 5644 2225 5666 2256
rect 5700 2225 5712 2256
rect 5628 2222 5666 2225
rect 5484 2215 5678 2222
rect 3282 2137 3316 2176
rect 3282 2064 3316 2103
rect 3282 1992 3316 2030
rect 3282 1920 3316 1958
rect 3282 1848 3316 1886
rect 3282 1776 3316 1814
rect 3282 1704 3316 1742
rect 3282 1632 3316 1670
rect 3282 1560 3316 1598
rect 3282 1488 3316 1526
rect 3282 1416 3316 1454
rect 3282 1344 3316 1382
rect 3282 1272 3316 1310
rect 3282 1200 3316 1238
rect 3282 1128 3316 1166
rect 3282 1056 3316 1094
rect 3282 984 3316 1022
rect 3282 912 3316 950
rect 3282 840 3316 878
rect 3282 768 3316 806
rect 3594 2137 3628 2176
rect 3594 2064 3628 2103
rect 3594 1992 3628 2030
rect 3594 1920 3628 1958
rect 3594 1848 3628 1886
rect 3594 1776 3628 1814
rect 3594 1704 3628 1742
rect 3594 1632 3628 1670
rect 3594 1560 3628 1598
rect 3594 1488 3628 1526
rect 3594 1416 3628 1454
rect 3594 1344 3628 1382
rect 3594 1272 3628 1310
rect 3594 1200 3628 1238
rect 3594 1128 3628 1166
rect 3594 1056 3628 1094
rect 3594 984 3628 1022
rect 3594 912 3628 950
rect 3594 840 3628 878
rect 3594 768 3628 806
rect 4110 2137 4144 2176
rect 4110 2064 4144 2103
rect 4110 1992 4144 2030
rect 4110 1920 4144 1958
rect 4110 1848 4144 1886
rect 4110 1776 4144 1814
rect 4110 1704 4144 1742
rect 4110 1632 4144 1670
rect 4110 1560 4144 1598
rect 4110 1488 4144 1526
rect 4110 1416 4144 1454
rect 4110 1344 4144 1382
rect 4110 1272 4144 1310
rect 4110 1200 4144 1238
rect 4110 1128 4144 1166
rect 4110 1056 4144 1094
rect 4110 984 4144 1022
rect 4110 912 4144 950
rect 4110 840 4144 878
rect 4110 768 4144 806
rect 3171 642 3172 676
rect 3221 642 3248 676
rect 3292 642 3324 676
rect 3363 642 3400 676
rect 3435 642 3473 676
rect 3510 642 3545 676
rect 3586 642 3617 676
rect 3662 642 3689 676
rect 3773 602 3965 738
rect 4422 2137 4456 2176
rect 4422 2064 4456 2103
rect 4422 1992 4456 2030
rect 4422 1920 4456 1958
rect 4422 1848 4456 1886
rect 4422 1776 4456 1814
rect 4422 1704 4456 1742
rect 4422 1632 4456 1670
rect 4422 1560 4456 1598
rect 4422 1488 4456 1526
rect 4422 1416 4456 1454
rect 4422 1344 4456 1382
rect 4422 1272 4456 1310
rect 4422 1200 4456 1238
rect 4422 1128 4456 1166
rect 4422 1056 4456 1094
rect 4422 984 4456 1022
rect 4422 912 4456 950
rect 4422 840 4456 878
rect 4422 768 4456 806
rect 4938 2137 4972 2176
rect 4938 2064 4972 2103
rect 4938 1992 4972 2030
rect 4938 1920 4972 1958
rect 4938 1848 4972 1886
rect 4938 1776 4972 1814
rect 4938 1704 4972 1742
rect 4938 1632 4972 1670
rect 4938 1560 4972 1598
rect 4938 1488 4972 1526
rect 4938 1416 4972 1454
rect 4938 1344 4972 1382
rect 4938 1272 4972 1310
rect 4938 1200 4972 1238
rect 4938 1128 4972 1166
rect 4938 1056 4972 1094
rect 4938 984 4972 1022
rect 4938 912 4972 950
rect 4938 840 4972 878
rect 4938 768 4972 806
rect 3999 642 4000 676
rect 4049 642 4076 676
rect 4120 642 4152 676
rect 4191 642 4228 676
rect 4263 642 4301 676
rect 4338 642 4373 676
rect 4414 642 4445 676
rect 4490 642 4517 676
rect 4601 602 4793 738
rect 5250 2137 5284 2176
rect 5250 2064 5284 2103
rect 5250 1992 5284 2030
rect 5250 1920 5284 1958
rect 5250 1848 5284 1886
rect 5250 1776 5284 1814
rect 5250 1704 5284 1742
rect 5250 1632 5284 1670
rect 5250 1560 5284 1598
rect 5250 1488 5284 1526
rect 5250 1416 5284 1454
rect 5250 1344 5284 1382
rect 5250 1272 5284 1310
rect 5250 1200 5284 1238
rect 5250 1128 5284 1166
rect 5250 1056 5284 1094
rect 5250 984 5284 1022
rect 5250 912 5284 950
rect 5250 840 5284 878
rect 5250 768 5284 806
rect 5450 2181 5522 2215
rect 5556 2191 5678 2215
rect 5556 2190 5712 2191
rect 5556 2183 5610 2190
rect 5644 2183 5712 2190
rect 5556 2181 5594 2183
rect 5450 2176 5594 2181
rect 5484 2149 5594 2176
rect 5644 2156 5666 2183
rect 5700 2156 5712 2183
rect 5628 2149 5666 2156
rect 5484 2142 5678 2149
rect 5450 2108 5522 2142
rect 5556 2122 5678 2142
rect 5556 2121 5712 2122
rect 5556 2110 5610 2121
rect 5644 2110 5712 2121
rect 5556 2108 5594 2110
rect 5450 2103 5594 2108
rect 5484 2076 5594 2103
rect 5644 2087 5666 2110
rect 5700 2087 5712 2110
rect 5628 2076 5666 2087
rect 5484 2069 5678 2076
rect 5450 2035 5522 2069
rect 5556 2053 5678 2069
rect 5556 2052 5712 2053
rect 5556 2037 5610 2052
rect 5644 2037 5712 2052
rect 5556 2035 5594 2037
rect 5450 2030 5594 2035
rect 5484 2003 5594 2030
rect 5644 2018 5666 2037
rect 5700 2018 5712 2037
rect 5628 2003 5666 2018
rect 5484 1996 5678 2003
rect 5450 1962 5522 1996
rect 5556 1984 5678 1996
rect 5556 1983 5712 1984
rect 5556 1964 5610 1983
rect 5644 1964 5712 1983
rect 5556 1962 5594 1964
rect 5450 1957 5594 1962
rect 5484 1930 5594 1957
rect 5644 1949 5666 1964
rect 5700 1949 5712 1964
rect 5628 1930 5666 1949
rect 5484 1923 5678 1930
rect 5450 1889 5522 1923
rect 5556 1915 5678 1923
rect 5556 1914 5712 1915
rect 5556 1891 5610 1914
rect 5644 1891 5712 1914
rect 5556 1889 5594 1891
rect 5450 1884 5594 1889
rect 5484 1857 5594 1884
rect 5644 1880 5666 1891
rect 5700 1880 5712 1891
rect 5628 1857 5666 1880
rect 5484 1850 5678 1857
rect 5450 1816 5522 1850
rect 5556 1846 5678 1850
rect 5556 1845 5712 1846
rect 5556 1818 5610 1845
rect 5644 1818 5712 1845
rect 5556 1816 5594 1818
rect 5450 1811 5594 1816
rect 5644 1811 5666 1818
rect 5700 1811 5712 1818
rect 5484 1784 5594 1811
rect 5628 1784 5666 1811
rect 5484 1777 5678 1784
rect 5450 1743 5522 1777
rect 5556 1776 5712 1777
rect 5556 1745 5610 1776
rect 5644 1745 5712 1776
rect 5556 1743 5594 1745
rect 5450 1738 5594 1743
rect 5644 1742 5666 1745
rect 5700 1742 5712 1745
rect 5484 1711 5594 1738
rect 5628 1711 5666 1742
rect 5484 1708 5678 1711
rect 5484 1707 5712 1708
rect 5484 1704 5610 1707
rect 5450 1670 5522 1704
rect 5556 1673 5610 1704
rect 5644 1673 5712 1707
rect 5556 1672 5678 1673
rect 5556 1670 5594 1672
rect 5450 1665 5594 1670
rect 5484 1638 5594 1665
rect 5628 1638 5666 1672
rect 5700 1638 5712 1639
rect 5484 1631 5610 1638
rect 5450 1597 5522 1631
rect 5556 1604 5610 1631
rect 5644 1604 5712 1638
rect 5556 1599 5678 1604
rect 5556 1597 5594 1599
rect 5450 1592 5594 1597
rect 5484 1565 5594 1592
rect 5628 1569 5666 1599
rect 5644 1565 5666 1569
rect 5700 1565 5712 1570
rect 5484 1558 5610 1565
rect 5450 1524 5522 1558
rect 5556 1535 5610 1558
rect 5644 1535 5712 1565
rect 5556 1526 5678 1535
rect 5556 1524 5594 1526
rect 5450 1519 5594 1524
rect 5484 1492 5594 1519
rect 5628 1500 5666 1526
rect 5644 1492 5666 1500
rect 5700 1492 5712 1501
rect 5484 1485 5610 1492
rect 5450 1451 5522 1485
rect 5556 1466 5610 1485
rect 5644 1466 5712 1492
rect 5556 1453 5678 1466
rect 5556 1451 5594 1453
rect 5450 1446 5594 1451
rect 5484 1419 5594 1446
rect 5628 1431 5666 1453
rect 5644 1419 5666 1431
rect 5700 1419 5712 1432
rect 5484 1412 5610 1419
rect 5450 1378 5522 1412
rect 5556 1397 5610 1412
rect 5644 1397 5712 1419
rect 5556 1380 5678 1397
rect 5556 1378 5594 1380
rect 5450 1373 5594 1378
rect 5484 1346 5594 1373
rect 5628 1362 5666 1380
rect 5644 1346 5666 1362
rect 5700 1346 5712 1363
rect 5484 1339 5610 1346
rect 5450 1305 5522 1339
rect 5556 1328 5610 1339
rect 5644 1328 5712 1346
rect 5556 1307 5678 1328
rect 5556 1305 5594 1307
rect 5450 1300 5594 1305
rect 5484 1273 5594 1300
rect 5628 1293 5666 1307
rect 5644 1273 5666 1293
rect 5700 1273 5712 1294
rect 5484 1266 5610 1273
rect 5450 1232 5522 1266
rect 5556 1259 5610 1266
rect 5644 1259 5712 1273
rect 5556 1234 5678 1259
rect 5556 1232 5594 1234
rect 5450 1227 5594 1232
rect 5484 1200 5594 1227
rect 5628 1224 5666 1234
rect 5644 1200 5666 1224
rect 5700 1200 5712 1225
rect 5484 1193 5610 1200
rect 5450 1159 5522 1193
rect 5556 1190 5610 1193
rect 5644 1190 5712 1200
rect 5556 1161 5678 1190
rect 5556 1159 5594 1161
rect 5450 1154 5594 1159
rect 5628 1155 5666 1161
rect 5484 1127 5594 1154
rect 5644 1127 5666 1155
rect 5700 1127 5712 1156
rect 5484 1121 5610 1127
rect 5644 1121 5712 1127
rect 5484 1120 5678 1121
rect 5450 1086 5522 1120
rect 5556 1088 5678 1120
rect 5556 1086 5594 1088
rect 5628 1086 5666 1088
rect 5450 1081 5594 1086
rect 5484 1054 5594 1081
rect 5644 1054 5666 1086
rect 5700 1054 5712 1087
rect 5484 1052 5610 1054
rect 5644 1052 5712 1054
rect 5484 1047 5678 1052
rect 5450 1013 5522 1047
rect 5556 1018 5678 1047
rect 5556 1017 5712 1018
rect 5556 1015 5610 1017
rect 5644 1015 5712 1017
rect 5556 1013 5594 1015
rect 5450 1008 5594 1013
rect 5484 981 5594 1008
rect 5644 983 5666 1015
rect 5700 983 5712 1015
rect 5628 981 5666 983
rect 5484 974 5678 981
rect 5450 940 5522 974
rect 5556 949 5678 974
rect 5556 948 5712 949
rect 5556 942 5610 948
rect 5644 942 5712 948
rect 5556 940 5594 942
rect 5450 935 5594 940
rect 5484 908 5594 935
rect 5644 914 5666 942
rect 5700 914 5712 942
rect 5628 908 5666 914
rect 5484 901 5678 908
rect 5450 867 5522 901
rect 5556 880 5678 901
rect 5556 879 5712 880
rect 5556 869 5610 879
rect 5644 869 5712 879
rect 5556 867 5594 869
rect 5450 862 5594 867
rect 5484 835 5594 862
rect 5644 845 5666 869
rect 5700 845 5712 869
rect 5628 835 5666 845
rect 5484 828 5678 835
rect 5450 794 5522 828
rect 5556 811 5678 828
rect 5556 810 5712 811
rect 5556 796 5610 810
rect 5644 796 5712 810
rect 5556 794 5594 796
rect 5450 789 5594 794
rect 5484 762 5594 789
rect 5644 776 5666 796
rect 5700 776 5712 796
rect 5628 762 5666 776
rect 5484 755 5678 762
rect 5450 721 5522 755
rect 5556 742 5678 755
rect 5556 741 5712 742
rect 5556 724 5610 741
rect 5576 723 5610 724
rect 5644 723 5712 741
rect 5450 716 5542 721
rect 5484 706 5542 716
rect 5576 706 5594 723
rect 5644 707 5666 723
rect 5700 707 5712 723
rect 5484 689 5594 706
rect 5628 689 5666 707
rect 5484 682 5678 689
rect 4827 642 4828 676
rect 4877 642 4904 676
rect 4948 642 4980 676
rect 5019 642 5056 676
rect 5091 642 5129 676
rect 5166 642 5201 676
rect 5242 642 5273 676
rect 5318 642 5345 676
rect 5450 648 5522 682
rect 5556 673 5678 682
rect 5556 672 5712 673
rect 5556 671 5610 672
rect 5576 650 5610 671
rect 5644 650 5712 672
rect 5450 643 5542 648
rect 5484 637 5542 643
rect 5576 637 5594 650
rect 5644 638 5666 650
rect 5700 638 5712 650
rect 5484 616 5594 637
rect 5628 616 5666 638
rect 5484 609 5678 616
rect 5450 602 5522 609
rect 5556 604 5678 609
rect 5556 603 5712 604
rect 5556 602 5610 603
rect 560 574 575 602
rect 404 568 438 573
rect 540 568 575 574
rect 609 570 644 602
rect 678 570 713 602
rect 747 570 782 602
rect 632 568 644 570
rect 705 568 713 570
rect 404 539 598 568
rect 370 536 598 539
rect 632 536 671 568
rect 705 536 744 568
rect 778 536 782 570
rect 370 534 782 536
rect 370 500 438 534
rect 472 500 507 534
rect 541 500 576 534
rect 610 500 645 534
rect 679 500 714 534
rect 370 498 714 500
rect 370 466 564 498
rect 598 466 637 498
rect 671 466 710 498
rect 370 432 404 466
rect 438 432 473 466
rect 507 432 542 466
rect 598 464 611 466
rect 671 464 680 466
rect 5576 569 5610 602
rect 5644 569 5712 603
rect 5576 535 5678 569
rect 5576 534 5712 535
rect 5644 500 5712 534
rect 5610 466 5678 500
rect 576 432 611 464
rect 645 432 680 464
rect 5610 432 5712 466
rect 170 164 204 196
rect 5882 164 5948 196
rect 170 130 174 164
rect 170 92 204 130
rect 5976 130 5980 162
rect 6014 130 6016 162
rect 170 58 174 92
rect 5976 94 6016 130
rect 5976 60 6084 94
rect 5976 58 5984 60
rect 170 26 204 58
rect 5950 26 5984 58
rect 6018 26 6118 60
<< viali >>
rect 209 4720 228 4734
rect 228 4720 243 4734
rect 282 4720 297 4734
rect 297 4720 316 4734
rect 355 4720 366 4734
rect 366 4720 389 4734
rect 428 4720 435 4734
rect 435 4720 462 4734
rect 501 4720 504 4734
rect 504 4720 535 4734
rect 209 4700 243 4720
rect 282 4700 316 4720
rect 355 4700 389 4720
rect 428 4700 462 4720
rect 501 4700 535 4720
rect 574 4700 608 4734
rect 647 4720 677 4734
rect 677 4720 681 4734
rect 720 4720 746 4734
rect 746 4720 754 4734
rect 793 4720 815 4734
rect 815 4720 827 4734
rect 866 4720 884 4734
rect 884 4720 900 4734
rect 939 4720 953 4734
rect 953 4720 973 4734
rect 1012 4720 1022 4734
rect 1022 4720 1046 4734
rect 1085 4720 1091 4734
rect 1091 4720 1119 4734
rect 1158 4720 1160 4734
rect 1160 4720 1192 4734
rect 1231 4720 1263 4734
rect 1263 4720 1265 4734
rect 1304 4720 1332 4734
rect 1332 4720 1338 4734
rect 1377 4720 1401 4734
rect 1401 4720 1411 4734
rect 1450 4720 1470 4734
rect 1470 4720 1484 4734
rect 1523 4720 1539 4734
rect 1539 4720 1557 4734
rect 1596 4720 1608 4734
rect 1608 4720 1630 4734
rect 1669 4720 1677 4734
rect 1677 4720 1703 4734
rect 1742 4720 1746 4734
rect 1746 4720 1776 4734
rect 647 4700 681 4720
rect 720 4700 754 4720
rect 793 4700 827 4720
rect 866 4700 900 4720
rect 939 4700 973 4720
rect 1012 4700 1046 4720
rect 1085 4700 1119 4720
rect 1158 4700 1192 4720
rect 1231 4700 1265 4720
rect 1304 4700 1338 4720
rect 1377 4700 1411 4720
rect 1450 4700 1484 4720
rect 1523 4700 1557 4720
rect 1596 4700 1630 4720
rect 1669 4700 1703 4720
rect 1742 4700 1776 4720
rect 1815 4700 1849 4734
rect 1888 4720 1919 4734
rect 1919 4720 1922 4734
rect 1961 4720 1988 4734
rect 1988 4720 1995 4734
rect 2034 4720 2057 4734
rect 2057 4720 2068 4734
rect 2107 4720 2126 4734
rect 2126 4720 2141 4734
rect 2180 4720 2195 4734
rect 2195 4720 2214 4734
rect 2253 4720 2264 4734
rect 2264 4720 2287 4734
rect 2326 4720 2333 4734
rect 2333 4720 2360 4734
rect 2399 4720 2402 4734
rect 2402 4720 2433 4734
rect 2472 4720 2505 4734
rect 2505 4720 2506 4734
rect 2545 4720 2574 4734
rect 2574 4720 2579 4734
rect 2618 4720 2643 4734
rect 2643 4720 2652 4734
rect 2691 4720 2712 4734
rect 2712 4720 2725 4734
rect 2764 4720 2781 4734
rect 2781 4720 2798 4734
rect 2837 4720 2850 4734
rect 2850 4720 2871 4734
rect 2910 4720 2919 4734
rect 2919 4720 2944 4734
rect 2983 4720 2988 4734
rect 2988 4720 3017 4734
rect 3056 4720 3057 4734
rect 3057 4720 3090 4734
rect 3129 4720 3161 4734
rect 3161 4720 3163 4734
rect 3202 4720 3230 4734
rect 3230 4720 3236 4734
rect 3275 4720 3299 4734
rect 3299 4720 3309 4734
rect 3348 4720 3368 4734
rect 3368 4720 3382 4734
rect 3421 4720 3437 4734
rect 3437 4720 3455 4734
rect 3494 4720 3506 4734
rect 3506 4720 3528 4734
rect 3567 4720 3575 4734
rect 3575 4720 3601 4734
rect 3640 4720 3644 4734
rect 3644 4720 3674 4734
rect 3713 4720 3747 4734
rect 1888 4700 1922 4720
rect 1961 4700 1995 4720
rect 2034 4700 2068 4720
rect 2107 4700 2141 4720
rect 2180 4700 2214 4720
rect 2253 4700 2287 4720
rect 2326 4700 2360 4720
rect 2399 4700 2433 4720
rect 2472 4700 2506 4720
rect 2545 4700 2579 4720
rect 2618 4700 2652 4720
rect 2691 4700 2725 4720
rect 2764 4700 2798 4720
rect 2837 4700 2871 4720
rect 2910 4700 2944 4720
rect 2983 4700 3017 4720
rect 3056 4700 3090 4720
rect 3129 4700 3163 4720
rect 3202 4700 3236 4720
rect 3275 4700 3309 4720
rect 3348 4700 3382 4720
rect 3421 4700 3455 4720
rect 3494 4700 3528 4720
rect 3567 4700 3601 4720
rect 3640 4700 3674 4720
rect 3713 4700 3747 4720
rect 3786 4700 3820 4734
rect 3859 4700 3893 4734
rect 3932 4700 3966 4734
rect 4005 4700 4039 4734
rect 4078 4700 4112 4734
rect 4151 4700 4185 4734
rect 4224 4700 4258 4734
rect 4297 4700 4331 4734
rect 4370 4700 4404 4734
rect 4443 4700 4477 4734
rect 4516 4700 4550 4734
rect 4589 4700 4623 4734
rect 4662 4700 4696 4734
rect 4735 4700 4769 4734
rect 4808 4700 4842 4734
rect 4881 4700 4915 4734
rect 209 4652 228 4662
rect 228 4652 243 4662
rect 282 4652 297 4662
rect 297 4652 316 4662
rect 355 4652 366 4662
rect 366 4652 389 4662
rect 428 4652 435 4662
rect 435 4652 462 4662
rect 501 4652 504 4662
rect 504 4652 535 4662
rect 209 4628 243 4652
rect 282 4628 316 4652
rect 355 4628 389 4652
rect 428 4628 462 4652
rect 501 4628 535 4652
rect 574 4628 608 4662
rect 647 4652 677 4662
rect 677 4652 681 4662
rect 720 4652 746 4662
rect 746 4652 754 4662
rect 793 4652 815 4662
rect 815 4652 827 4662
rect 866 4652 884 4662
rect 884 4652 900 4662
rect 939 4652 953 4662
rect 953 4652 973 4662
rect 1012 4652 1022 4662
rect 1022 4652 1046 4662
rect 1085 4652 1091 4662
rect 1091 4652 1119 4662
rect 1158 4652 1160 4662
rect 1160 4652 1192 4662
rect 1231 4652 1263 4662
rect 1263 4652 1265 4662
rect 1304 4652 1332 4662
rect 1332 4652 1338 4662
rect 1377 4652 1401 4662
rect 1401 4652 1411 4662
rect 1450 4652 1470 4662
rect 1470 4652 1484 4662
rect 1523 4652 1539 4662
rect 1539 4652 1557 4662
rect 1596 4652 1608 4662
rect 1608 4652 1630 4662
rect 1669 4652 1677 4662
rect 1677 4652 1703 4662
rect 1742 4652 1746 4662
rect 1746 4652 1776 4662
rect 647 4628 681 4652
rect 720 4628 754 4652
rect 793 4628 827 4652
rect 866 4628 900 4652
rect 939 4628 973 4652
rect 1012 4628 1046 4652
rect 1085 4628 1119 4652
rect 1158 4628 1192 4652
rect 1231 4628 1265 4652
rect 1304 4628 1338 4652
rect 1377 4628 1411 4652
rect 1450 4628 1484 4652
rect 1523 4628 1557 4652
rect 1596 4628 1630 4652
rect 1669 4628 1703 4652
rect 1742 4628 1776 4652
rect 1815 4628 1849 4662
rect 1888 4652 1919 4662
rect 1919 4652 1922 4662
rect 1961 4652 1988 4662
rect 1988 4652 1995 4662
rect 2034 4652 2057 4662
rect 2057 4652 2068 4662
rect 2107 4652 2126 4662
rect 2126 4652 2141 4662
rect 2180 4652 2195 4662
rect 2195 4652 2214 4662
rect 2253 4652 2264 4662
rect 2264 4652 2287 4662
rect 2326 4652 2333 4662
rect 2333 4652 2360 4662
rect 2399 4652 2402 4662
rect 2402 4652 2433 4662
rect 2472 4652 2505 4662
rect 2505 4652 2506 4662
rect 2545 4652 2574 4662
rect 2574 4652 2579 4662
rect 2618 4652 2643 4662
rect 2643 4652 2652 4662
rect 2691 4652 2712 4662
rect 2712 4652 2725 4662
rect 2764 4652 2781 4662
rect 2781 4652 2798 4662
rect 2837 4652 2850 4662
rect 2850 4652 2871 4662
rect 2910 4652 2919 4662
rect 2919 4652 2944 4662
rect 2983 4652 2988 4662
rect 2988 4652 3017 4662
rect 3056 4652 3057 4662
rect 3057 4652 3090 4662
rect 3129 4652 3161 4662
rect 3161 4652 3163 4662
rect 3202 4652 3230 4662
rect 3230 4652 3236 4662
rect 3275 4652 3299 4662
rect 3299 4652 3309 4662
rect 3348 4652 3368 4662
rect 3368 4652 3382 4662
rect 3421 4652 3437 4662
rect 3437 4652 3455 4662
rect 3494 4652 3506 4662
rect 3506 4652 3528 4662
rect 3567 4652 3575 4662
rect 3575 4652 3601 4662
rect 3640 4652 3644 4662
rect 3644 4652 3674 4662
rect 3713 4652 3747 4662
rect 1888 4628 1922 4652
rect 1961 4628 1995 4652
rect 2034 4628 2068 4652
rect 2107 4628 2141 4652
rect 2180 4628 2214 4652
rect 2253 4628 2287 4652
rect 2326 4628 2360 4652
rect 2399 4628 2433 4652
rect 2472 4628 2506 4652
rect 2545 4628 2579 4652
rect 2618 4628 2652 4652
rect 2691 4628 2725 4652
rect 2764 4628 2798 4652
rect 2837 4628 2871 4652
rect 2910 4628 2944 4652
rect 2983 4628 3017 4652
rect 3056 4628 3090 4652
rect 3129 4628 3163 4652
rect 3202 4628 3236 4652
rect 3275 4628 3309 4652
rect 3348 4628 3382 4652
rect 3421 4628 3455 4652
rect 3494 4628 3528 4652
rect 3567 4628 3601 4652
rect 3640 4628 3674 4652
rect 3713 4628 3747 4652
rect 3786 4628 3820 4662
rect 3859 4628 3893 4662
rect 3932 4628 3966 4662
rect 4005 4628 4039 4662
rect 4078 4628 4112 4662
rect 4151 4628 4185 4662
rect 4224 4628 4258 4662
rect 4297 4628 4331 4662
rect 4370 4628 4404 4662
rect 4443 4628 4477 4662
rect 4516 4628 4550 4662
rect 4589 4628 4623 4662
rect 4662 4628 4696 4662
rect 4735 4628 4769 4662
rect 4808 4628 4842 4662
rect 4881 4628 4915 4662
rect 4954 4628 5924 4734
rect 5980 4582 6086 4612
rect 5980 4548 6084 4582
rect 6084 4548 6086 4582
rect 382 4254 416 4288
rect 455 4287 489 4288
rect 528 4287 562 4288
rect 601 4287 635 4288
rect 674 4287 708 4288
rect 747 4287 781 4288
rect 820 4287 854 4288
rect 893 4287 927 4288
rect 966 4287 1000 4288
rect 1039 4287 1073 4288
rect 1112 4287 1146 4288
rect 1185 4287 1219 4288
rect 1258 4287 1292 4288
rect 1331 4287 1365 4288
rect 1404 4287 1438 4288
rect 1477 4287 1511 4288
rect 1550 4287 1584 4288
rect 1623 4287 1657 4288
rect 1696 4287 1730 4288
rect 1769 4287 1803 4288
rect 1842 4287 1876 4288
rect 1915 4287 1949 4288
rect 1988 4287 2022 4288
rect 2061 4287 2095 4288
rect 2134 4287 2168 4288
rect 2207 4287 2241 4288
rect 2280 4287 2314 4288
rect 2353 4287 2387 4288
rect 2426 4287 2471 4288
rect 455 4254 470 4287
rect 470 4254 489 4287
rect 528 4254 539 4287
rect 539 4254 562 4287
rect 601 4254 608 4287
rect 608 4254 635 4287
rect 674 4254 677 4287
rect 677 4254 708 4287
rect 747 4254 780 4287
rect 780 4254 781 4287
rect 820 4254 849 4287
rect 849 4254 854 4287
rect 893 4254 918 4287
rect 918 4254 927 4287
rect 966 4254 987 4287
rect 987 4254 1000 4287
rect 1039 4254 1056 4287
rect 1056 4254 1073 4287
rect 1112 4254 1125 4287
rect 1125 4254 1146 4287
rect 1185 4254 1194 4287
rect 1194 4254 1219 4287
rect 1258 4254 1263 4287
rect 1263 4254 1292 4287
rect 1331 4254 1332 4287
rect 1332 4254 1365 4287
rect 1404 4254 1436 4287
rect 1436 4254 1438 4287
rect 1477 4254 1505 4287
rect 1505 4254 1511 4287
rect 1550 4254 1574 4287
rect 1574 4254 1584 4287
rect 1623 4254 1643 4287
rect 1643 4254 1657 4287
rect 1696 4254 1712 4287
rect 1712 4254 1730 4287
rect 1769 4254 1781 4287
rect 1781 4254 1803 4287
rect 1842 4254 1850 4287
rect 1850 4254 1876 4287
rect 1915 4254 1919 4287
rect 1919 4254 1949 4287
rect 1988 4254 2022 4287
rect 2061 4254 2091 4287
rect 2091 4254 2095 4287
rect 2134 4254 2160 4287
rect 2160 4254 2168 4287
rect 2207 4254 2229 4287
rect 2229 4254 2241 4287
rect 2280 4254 2298 4287
rect 2298 4254 2314 4287
rect 2353 4254 2367 4287
rect 2367 4254 2387 4287
rect 2426 4253 2436 4287
rect 2436 4253 2471 4287
rect 2426 4219 2471 4253
rect 382 4182 416 4216
rect 455 4185 470 4216
rect 470 4185 489 4216
rect 528 4185 539 4216
rect 539 4185 562 4216
rect 601 4185 608 4216
rect 608 4185 635 4216
rect 674 4185 677 4216
rect 677 4185 708 4216
rect 747 4185 780 4216
rect 780 4185 781 4216
rect 820 4185 849 4216
rect 849 4185 854 4216
rect 893 4185 918 4216
rect 918 4185 927 4216
rect 966 4185 987 4216
rect 987 4185 1000 4216
rect 1039 4185 1056 4216
rect 1056 4185 1073 4216
rect 1112 4185 1125 4216
rect 1125 4185 1146 4216
rect 1185 4185 1194 4216
rect 1194 4185 1219 4216
rect 1258 4185 1263 4216
rect 1263 4185 1292 4216
rect 1331 4185 1332 4216
rect 1332 4185 1365 4216
rect 1404 4185 1436 4216
rect 1436 4185 1438 4216
rect 1477 4185 1505 4216
rect 1505 4185 1511 4216
rect 1550 4185 1574 4216
rect 1574 4185 1584 4216
rect 1623 4185 1643 4216
rect 1643 4185 1657 4216
rect 1696 4185 1712 4216
rect 1712 4185 1730 4216
rect 1769 4185 1781 4216
rect 1781 4185 1803 4216
rect 1842 4185 1850 4216
rect 1850 4185 1876 4216
rect 1915 4185 1919 4216
rect 1919 4185 1949 4216
rect 1988 4185 2022 4216
rect 2061 4185 2091 4216
rect 2091 4185 2095 4216
rect 2134 4185 2160 4216
rect 2160 4185 2168 4216
rect 2207 4185 2229 4216
rect 2229 4185 2241 4216
rect 2280 4185 2298 4216
rect 2298 4185 2314 4216
rect 2353 4185 2367 4216
rect 2367 4185 2387 4216
rect 2426 4185 2436 4219
rect 2436 4185 2471 4219
rect 455 4182 489 4185
rect 528 4182 562 4185
rect 601 4182 635 4185
rect 674 4182 708 4185
rect 747 4182 781 4185
rect 820 4182 854 4185
rect 893 4182 927 4185
rect 966 4182 1000 4185
rect 1039 4182 1073 4185
rect 1112 4182 1146 4185
rect 1185 4182 1219 4185
rect 1258 4182 1292 4185
rect 1331 4182 1365 4185
rect 1404 4182 1438 4185
rect 1477 4182 1511 4185
rect 1550 4182 1584 4185
rect 1623 4182 1657 4185
rect 1696 4182 1730 4185
rect 1769 4182 1803 4185
rect 1842 4182 1876 4185
rect 1915 4182 1949 4185
rect 1988 4182 2022 4185
rect 2061 4182 2095 4185
rect 2134 4182 2168 4185
rect 2207 4182 2241 4185
rect 2280 4182 2314 4185
rect 2353 4182 2387 4185
rect 2426 4151 2471 4185
rect 382 4110 416 4144
rect 455 4117 470 4144
rect 470 4117 489 4144
rect 528 4117 539 4144
rect 539 4117 562 4144
rect 601 4117 608 4144
rect 608 4117 635 4144
rect 674 4117 677 4144
rect 677 4117 708 4144
rect 747 4117 780 4144
rect 780 4117 781 4144
rect 820 4117 849 4144
rect 849 4117 854 4144
rect 893 4117 918 4144
rect 918 4117 927 4144
rect 966 4117 987 4144
rect 987 4117 1000 4144
rect 1039 4117 1056 4144
rect 1056 4117 1073 4144
rect 1112 4117 1125 4144
rect 1125 4117 1146 4144
rect 1185 4117 1194 4144
rect 1194 4117 1219 4144
rect 1258 4117 1263 4144
rect 1263 4117 1292 4144
rect 1331 4117 1332 4144
rect 1332 4117 1365 4144
rect 1404 4117 1436 4144
rect 1436 4117 1438 4144
rect 1477 4117 1505 4144
rect 1505 4117 1511 4144
rect 1550 4117 1574 4144
rect 1574 4117 1584 4144
rect 1623 4117 1643 4144
rect 1643 4117 1657 4144
rect 1696 4117 1712 4144
rect 1712 4117 1730 4144
rect 1769 4117 1781 4144
rect 1781 4117 1803 4144
rect 1842 4117 1850 4144
rect 1850 4117 1876 4144
rect 1915 4117 1919 4144
rect 1919 4117 1949 4144
rect 1988 4117 2022 4144
rect 2061 4117 2091 4144
rect 2091 4117 2095 4144
rect 2134 4117 2160 4144
rect 2160 4117 2168 4144
rect 2207 4117 2229 4144
rect 2229 4117 2241 4144
rect 2280 4117 2298 4144
rect 2298 4117 2314 4144
rect 2353 4117 2367 4144
rect 2367 4117 2387 4144
rect 2426 4117 2436 4151
rect 2436 4117 2471 4151
rect 2471 4117 5633 4288
rect 5633 4117 5700 4288
rect 455 4110 489 4117
rect 528 4110 562 4117
rect 601 4110 635 4117
rect 674 4110 708 4117
rect 747 4110 781 4117
rect 820 4110 854 4117
rect 893 4110 927 4117
rect 966 4110 1000 4117
rect 1039 4110 1073 4117
rect 1112 4110 1146 4117
rect 1185 4110 1219 4117
rect 1258 4110 1292 4117
rect 1331 4110 1365 4117
rect 1404 4110 1438 4117
rect 1477 4110 1511 4117
rect 1550 4110 1584 4117
rect 1623 4110 1657 4117
rect 1696 4110 1730 4117
rect 1769 4110 1803 4117
rect 1842 4110 1876 4117
rect 1915 4110 1949 4117
rect 1988 4110 2022 4117
rect 2061 4110 2095 4117
rect 2134 4110 2168 4117
rect 2207 4110 2241 4117
rect 2280 4110 2314 4117
rect 2353 4110 2387 4117
rect 382 4038 416 4072
rect 455 4038 489 4072
rect 528 4038 562 4072
rect 601 4038 635 4072
rect 674 4038 708 4072
rect 747 4038 781 4072
rect 820 4038 854 4072
rect 893 4038 927 4072
rect 966 4038 1000 4072
rect 1039 4038 1073 4072
rect 1112 4038 1146 4072
rect 1185 4038 1219 4072
rect 1258 4038 1292 4072
rect 1331 4038 1365 4072
rect 1404 4038 1438 4072
rect 1477 4038 1511 4072
rect 1550 4038 1584 4072
rect 1623 4038 1657 4072
rect 1696 4038 1730 4072
rect 1769 4038 1803 4072
rect 1842 4038 1876 4072
rect 1915 4038 1949 4072
rect 1988 4038 2022 4072
rect 2061 4038 2095 4072
rect 2134 4038 2168 4072
rect 2207 4038 2241 4072
rect 2280 4038 2314 4072
rect 2353 4038 2387 4072
rect 2426 4038 5700 4117
rect 2426 4032 3334 4038
rect 5125 4032 5231 4038
rect 636 3966 670 4000
rect 708 3966 742 4000
rect 780 3966 814 4000
rect 852 3966 886 4000
rect 924 3966 958 4000
rect 996 3966 1030 4000
rect 1068 3966 1102 4000
rect 1140 3966 1174 4000
rect 1212 3966 1246 4000
rect 1284 3966 1318 4000
rect 1356 3966 1390 4000
rect 1428 3966 1462 4000
rect 1500 3966 1534 4000
rect 1572 3966 1606 4000
rect 1644 3966 1678 4000
rect 1716 3966 1750 4000
rect 1788 3966 1822 4000
rect 1860 3966 1894 4000
rect 1932 3966 1966 4000
rect 2004 3966 2038 4000
rect 2076 3966 2110 4000
rect 2148 3966 2182 4000
rect 2220 3966 2254 4000
rect 2292 3966 2326 4000
rect 2364 3966 2398 4000
rect 2426 3966 3334 4032
rect 3373 3966 3407 4000
rect 3446 3966 3480 4000
rect 3519 3966 3553 4000
rect 3592 3966 3626 4000
rect 3665 3966 3699 4000
rect 3738 3966 3772 4000
rect 3811 3966 3845 4000
rect 3884 3966 3918 4000
rect 3957 3966 3991 4000
rect 4030 3966 4064 4000
rect 4103 3966 4137 4000
rect 4176 3966 4210 4000
rect 4249 3966 4283 4000
rect 4322 3966 4356 4000
rect 4395 3966 4429 4000
rect 4468 3966 4502 4000
rect 4541 3966 4575 4000
rect 4614 3966 4648 4000
rect 4687 3966 4721 4000
rect 4760 3966 4794 4000
rect 4833 3966 4867 4000
rect 4906 3966 4940 4000
rect 4979 3966 5013 4000
rect 5052 3966 5086 4000
rect 526 3928 560 3962
rect 598 3894 632 3928
rect 671 3894 705 3928
rect 744 3894 778 3928
rect 817 3894 851 3928
rect 890 3894 924 3928
rect 963 3894 997 3928
rect 1036 3894 1070 3928
rect 1109 3894 1143 3928
rect 1182 3894 1216 3928
rect 1255 3894 1289 3928
rect 1328 3894 1362 3928
rect 1401 3894 1435 3928
rect 1474 3894 1508 3928
rect 1547 3894 1581 3928
rect 1620 3894 1654 3928
rect 1693 3894 1727 3928
rect 1766 3894 1800 3928
rect 1839 3894 1873 3928
rect 1912 3894 1946 3928
rect 1985 3894 2019 3928
rect 2058 3894 2092 3928
rect 2131 3894 2165 3928
rect 2204 3894 2238 3928
rect 2277 3894 2311 3928
rect 2350 3894 2384 3928
rect 2423 3894 2457 3928
rect 2496 3894 2530 3928
rect 2569 3894 2603 3928
rect 2642 3894 2676 3928
rect 2715 3894 2749 3928
rect 2788 3894 2822 3928
rect 2861 3894 2895 3928
rect 2934 3894 2968 3928
rect 3007 3894 3041 3928
rect 3080 3894 3114 3928
rect 3153 3894 3187 3928
rect 3226 3894 3260 3928
rect 3299 3894 3333 3928
rect 3372 3894 3406 3928
rect 3445 3894 3479 3928
rect 3518 3894 3552 3928
rect 3591 3894 3625 3928
rect 3664 3894 3698 3928
rect 3737 3894 3771 3928
rect 3810 3894 3844 3928
rect 3883 3894 3917 3928
rect 3956 3894 3990 3928
rect 4029 3894 4063 3928
rect 4102 3894 4136 3928
rect 4175 3894 4209 3928
rect 4248 3894 4282 3928
rect 4321 3894 4355 3928
rect 4394 3894 4428 3928
rect 4467 3894 4501 3928
rect 4540 3894 4574 3928
rect 4613 3894 4647 3928
rect 4686 3894 4720 3928
rect 4759 3894 4793 3928
rect 4832 3894 4866 3928
rect 4905 3894 4939 3928
rect 4978 3894 5012 3928
rect 5051 3894 5085 3928
rect 5125 3894 5231 4032
rect 5292 3966 5326 4000
rect 5388 3998 5402 4000
rect 5402 3998 5422 4000
rect 5484 3998 5506 4000
rect 5506 3998 5518 4000
rect 5388 3966 5422 3998
rect 5484 3966 5518 3998
rect 5281 3894 5300 3928
rect 5300 3894 5315 3928
rect 5365 3896 5399 3928
rect 5450 3896 5484 3928
rect 5365 3894 5369 3896
rect 5369 3894 5399 3896
rect 526 3862 560 3889
rect 5450 3894 5473 3896
rect 5473 3894 5484 3896
rect 526 3855 560 3862
rect 382 3826 404 3850
rect 404 3826 488 3850
rect 382 3824 488 3826
rect 382 3791 438 3824
rect 382 3757 404 3791
rect 404 3790 438 3791
rect 438 3790 472 3824
rect 472 3790 488 3824
rect 598 3821 632 3855
rect 526 3792 540 3816
rect 540 3792 560 3816
rect 404 3757 488 3790
rect 526 3782 560 3792
rect 382 3754 488 3757
rect 382 3722 438 3754
rect 382 3688 404 3722
rect 404 3720 438 3722
rect 438 3720 472 3754
rect 472 3720 488 3754
rect 598 3748 632 3782
rect 687 3806 721 3818
rect 763 3806 797 3818
rect 839 3806 873 3818
rect 915 3806 949 3818
rect 991 3806 1025 3818
rect 1067 3806 1101 3818
rect 1144 3806 1178 3818
rect 1221 3806 1255 3818
rect 687 3784 703 3806
rect 703 3784 721 3806
rect 763 3784 774 3806
rect 774 3784 797 3806
rect 839 3784 845 3806
rect 845 3784 873 3806
rect 915 3784 917 3806
rect 917 3784 949 3806
rect 991 3784 1023 3806
rect 1023 3784 1025 3806
rect 1067 3784 1095 3806
rect 1095 3784 1101 3806
rect 1144 3784 1167 3806
rect 1167 3784 1178 3806
rect 1221 3784 1239 3806
rect 1239 3784 1255 3806
rect 526 3724 540 3743
rect 540 3724 560 3743
rect 404 3688 488 3720
rect 526 3709 560 3724
rect 1515 3806 1549 3818
rect 1591 3806 1625 3818
rect 1667 3806 1701 3818
rect 1743 3806 1777 3818
rect 1819 3806 1853 3818
rect 1895 3806 1929 3818
rect 1972 3806 2006 3818
rect 2049 3806 2083 3818
rect 1515 3784 1531 3806
rect 1531 3784 1549 3806
rect 1591 3784 1602 3806
rect 1602 3784 1625 3806
rect 1667 3784 1673 3806
rect 1673 3784 1701 3806
rect 1743 3784 1745 3806
rect 1745 3784 1777 3806
rect 1819 3784 1851 3806
rect 1851 3784 1853 3806
rect 1895 3784 1923 3806
rect 1923 3784 1929 3806
rect 1972 3784 1995 3806
rect 1995 3784 2006 3806
rect 2049 3784 2067 3806
rect 2067 3784 2083 3806
rect 2343 3806 2377 3818
rect 2419 3806 2453 3818
rect 2495 3806 2529 3818
rect 2571 3806 2605 3818
rect 2647 3806 2681 3818
rect 2723 3806 2757 3818
rect 2800 3806 2834 3818
rect 2877 3806 2911 3818
rect 2343 3784 2359 3806
rect 2359 3784 2377 3806
rect 2419 3784 2430 3806
rect 2430 3784 2453 3806
rect 2495 3784 2501 3806
rect 2501 3784 2529 3806
rect 2571 3784 2573 3806
rect 2573 3784 2605 3806
rect 2647 3784 2679 3806
rect 2679 3784 2681 3806
rect 2723 3784 2751 3806
rect 2751 3784 2757 3806
rect 2800 3784 2823 3806
rect 2823 3784 2834 3806
rect 2877 3784 2895 3806
rect 2895 3784 2911 3806
rect 382 3684 488 3688
rect 382 3653 438 3684
rect 382 3619 404 3653
rect 404 3650 438 3653
rect 438 3650 472 3684
rect 472 3650 488 3684
rect 598 3675 632 3709
rect 404 3619 488 3650
rect 526 3636 560 3670
rect 382 3614 488 3619
rect 382 3584 438 3614
rect 382 3550 404 3584
rect 404 3580 438 3584
rect 438 3580 472 3614
rect 472 3580 488 3614
rect 598 3602 632 3636
rect 404 3550 488 3580
rect 526 3563 560 3597
rect 382 3544 488 3550
rect 382 3515 438 3544
rect 382 3481 404 3515
rect 404 3510 438 3515
rect 438 3510 472 3544
rect 472 3510 488 3544
rect 598 3529 632 3563
rect 404 3481 488 3510
rect 526 3490 560 3524
rect 382 3474 488 3481
rect 382 3446 438 3474
rect 382 3412 404 3446
rect 404 3440 438 3446
rect 438 3440 472 3474
rect 472 3440 488 3474
rect 598 3456 632 3490
rect 404 3412 488 3440
rect 526 3417 560 3451
rect 382 3404 488 3412
rect 382 3377 438 3404
rect 382 3343 404 3377
rect 404 3370 438 3377
rect 438 3370 472 3404
rect 472 3370 488 3404
rect 598 3383 632 3417
rect 404 3343 488 3370
rect 526 3344 560 3378
rect 382 3334 488 3343
rect 382 3308 438 3334
rect 382 3274 404 3308
rect 404 3300 438 3308
rect 438 3300 472 3334
rect 472 3300 488 3334
rect 598 3310 632 3344
rect 404 3274 488 3300
rect 382 3264 488 3274
rect 526 3271 560 3305
rect 382 3239 438 3264
rect 382 3205 404 3239
rect 404 3230 438 3239
rect 438 3230 472 3264
rect 472 3230 488 3264
rect 598 3237 632 3271
rect 404 3205 488 3230
rect 382 3194 488 3205
rect 526 3198 560 3232
rect 382 3170 438 3194
rect 382 3136 404 3170
rect 404 3160 438 3170
rect 438 3160 472 3194
rect 472 3160 488 3194
rect 598 3164 632 3198
rect 404 3136 488 3160
rect 382 3124 488 3136
rect 526 3125 560 3159
rect 382 3101 438 3124
rect 382 3067 404 3101
rect 404 3090 438 3101
rect 438 3090 472 3124
rect 472 3090 488 3124
rect 598 3091 632 3125
rect 404 3067 488 3090
rect 382 3054 488 3067
rect 382 3032 438 3054
rect 382 2998 404 3032
rect 404 3020 438 3032
rect 438 3020 472 3054
rect 472 3020 488 3054
rect 526 3052 560 3086
rect 404 2998 488 3020
rect 598 3018 632 3052
rect 382 2984 488 2998
rect 382 2963 438 2984
rect 382 2952 404 2963
rect 404 2952 438 2963
rect 438 2952 472 2984
rect 472 2952 488 2984
rect 526 2979 560 3013
rect 598 2945 632 2979
rect 382 2894 416 2913
rect 382 2879 404 2894
rect 404 2879 416 2894
rect 454 2880 472 2913
rect 472 2880 488 2913
rect 526 2906 560 2940
rect 454 2879 488 2880
rect 598 2872 632 2906
rect 382 2825 416 2840
rect 382 2806 404 2825
rect 404 2806 416 2825
rect 454 2810 472 2840
rect 472 2810 488 2840
rect 526 2833 560 2867
rect 454 2806 488 2810
rect 598 2799 632 2833
rect 382 2756 416 2767
rect 382 2733 404 2756
rect 404 2733 416 2756
rect 454 2740 472 2767
rect 472 2740 488 2767
rect 526 2760 560 2794
rect 454 2733 488 2740
rect 598 2726 632 2760
rect 382 2687 416 2694
rect 382 2660 404 2687
rect 404 2660 416 2687
rect 454 2670 472 2694
rect 472 2670 488 2694
rect 526 2687 560 2721
rect 454 2660 488 2670
rect 598 2653 632 2687
rect 382 2618 416 2621
rect 382 2587 404 2618
rect 404 2587 416 2618
rect 454 2600 472 2621
rect 472 2600 488 2621
rect 526 2614 560 2648
rect 454 2587 488 2600
rect 598 2580 632 2614
rect 382 2515 404 2548
rect 404 2515 416 2548
rect 454 2530 472 2548
rect 472 2530 488 2548
rect 526 2541 560 2575
rect 382 2514 416 2515
rect 454 2514 488 2530
rect 598 2507 632 2541
rect 382 2446 404 2475
rect 404 2446 416 2475
rect 454 2460 472 2475
rect 472 2460 488 2475
rect 526 2468 560 2502
rect 382 2441 416 2446
rect 454 2441 488 2460
rect 598 2434 632 2468
rect 382 2377 404 2402
rect 404 2377 416 2402
rect 454 2390 472 2402
rect 472 2390 488 2402
rect 526 2395 560 2429
rect 382 2368 416 2377
rect 454 2368 488 2390
rect 598 2361 632 2395
rect 382 2308 404 2329
rect 404 2308 416 2329
rect 454 2320 472 2329
rect 472 2320 488 2329
rect 526 2322 560 2356
rect 382 2295 416 2308
rect 454 2295 488 2320
rect 598 2288 632 2322
rect 382 2239 404 2256
rect 404 2239 416 2256
rect 454 2250 472 2256
rect 472 2250 488 2256
rect 382 2222 416 2239
rect 454 2222 488 2250
rect 526 2249 560 2283
rect 954 3704 988 3738
rect 954 3631 988 3665
rect 954 3558 988 3592
rect 954 3486 988 3520
rect 954 3414 988 3448
rect 954 3342 988 3376
rect 954 3270 988 3304
rect 954 3198 988 3232
rect 954 3126 988 3160
rect 954 3054 988 3088
rect 954 2982 988 3016
rect 954 2910 988 2944
rect 954 2838 988 2872
rect 954 2766 988 2800
rect 954 2694 988 2728
rect 954 2622 988 2656
rect 954 2550 988 2584
rect 954 2478 988 2512
rect 954 2406 988 2440
rect 954 2334 988 2368
rect 954 2262 988 2296
rect 1297 3704 1331 3738
rect 1369 3704 1403 3738
rect 1441 3704 1475 3738
rect 1297 3631 1331 3665
rect 1369 3631 1403 3665
rect 1441 3631 1475 3665
rect 1297 2262 1475 3592
rect 1782 3704 1816 3738
rect 1782 3631 1816 3665
rect 1782 3558 1816 3592
rect 1782 3486 1816 3520
rect 1782 3414 1816 3448
rect 1782 3342 1816 3376
rect 1782 3270 1816 3304
rect 1782 3198 1816 3232
rect 1782 3126 1816 3160
rect 1782 3054 1816 3088
rect 1782 2982 1816 3016
rect 1782 2910 1816 2944
rect 1782 2838 1816 2872
rect 1782 2766 1816 2800
rect 1782 2694 1816 2728
rect 1782 2622 1816 2656
rect 1782 2550 1816 2584
rect 1782 2478 1816 2512
rect 1782 2406 1816 2440
rect 1782 2334 1816 2368
rect 1782 2262 1816 2296
rect 2124 3704 2158 3738
rect 2196 3704 2230 3738
rect 2268 3704 2302 3738
rect 2124 3631 2158 3665
rect 2196 3631 2230 3665
rect 2268 3631 2302 3665
rect 2124 2262 2302 3592
rect 2610 3704 2644 3738
rect 2610 3631 2644 3665
rect 2610 3558 2644 3592
rect 2610 3486 2644 3520
rect 2610 3414 2644 3448
rect 2610 3342 2644 3376
rect 2610 3270 2644 3304
rect 2610 3198 2644 3232
rect 2610 3126 2644 3160
rect 2610 3054 2644 3088
rect 2610 2982 2644 3016
rect 2610 2910 2644 2944
rect 2610 2838 2644 2872
rect 2610 2766 2644 2800
rect 2610 2694 2644 2728
rect 2610 2622 2644 2656
rect 2610 2550 2644 2584
rect 2610 2478 2644 2512
rect 2610 2406 2644 2440
rect 2610 2334 2644 2368
rect 2610 2262 2644 2296
rect 598 2215 632 2249
rect 382 2170 404 2183
rect 404 2170 416 2183
rect 454 2180 472 2183
rect 472 2180 488 2183
rect 382 2149 416 2170
rect 454 2149 488 2180
rect 526 2176 560 2210
rect 598 2142 632 2176
rect 382 2101 404 2110
rect 404 2101 416 2110
rect 382 2076 416 2101
rect 454 2076 488 2110
rect 526 2103 560 2137
rect 598 2069 632 2103
rect 382 2032 404 2037
rect 404 2032 416 2037
rect 382 2003 416 2032
rect 454 2006 488 2037
rect 526 2030 560 2064
rect 454 2003 472 2006
rect 472 2003 488 2006
rect 598 1996 632 2030
rect 382 1963 404 1964
rect 404 1963 416 1964
rect 382 1930 416 1963
rect 454 1937 488 1964
rect 526 1957 560 1991
rect 454 1930 472 1937
rect 472 1930 488 1937
rect 598 1923 632 1957
rect 382 1861 416 1891
rect 454 1868 488 1891
rect 526 1884 560 1918
rect 382 1857 404 1861
rect 404 1857 416 1861
rect 454 1857 472 1868
rect 472 1857 488 1868
rect 598 1850 632 1884
rect 382 1793 416 1818
rect 454 1799 488 1818
rect 526 1811 560 1845
rect 382 1784 404 1793
rect 404 1784 416 1793
rect 454 1784 472 1799
rect 472 1784 488 1799
rect 598 1777 632 1811
rect 382 1725 416 1745
rect 454 1730 488 1745
rect 526 1738 560 1772
rect 382 1711 404 1725
rect 404 1711 416 1725
rect 454 1711 472 1730
rect 472 1711 488 1730
rect 598 1704 632 1738
rect 382 1657 416 1672
rect 454 1661 488 1672
rect 526 1665 560 1699
rect 382 1638 404 1657
rect 404 1638 416 1657
rect 454 1638 472 1661
rect 472 1638 488 1661
rect 598 1631 632 1665
rect 382 1589 416 1599
rect 454 1592 488 1599
rect 526 1592 560 1626
rect 382 1565 404 1589
rect 404 1565 416 1589
rect 454 1565 472 1592
rect 472 1565 488 1592
rect 598 1558 632 1592
rect 382 1521 416 1526
rect 454 1523 488 1526
rect 382 1492 404 1521
rect 404 1492 416 1521
rect 454 1492 472 1523
rect 472 1492 488 1523
rect 526 1519 560 1553
rect 598 1485 632 1519
rect 382 1419 404 1453
rect 404 1419 416 1453
rect 454 1420 472 1453
rect 472 1420 488 1453
rect 526 1446 560 1480
rect 454 1419 488 1420
rect 598 1412 632 1446
rect 382 1351 404 1380
rect 404 1351 416 1380
rect 454 1351 472 1380
rect 472 1351 488 1380
rect 526 1373 560 1407
rect 382 1346 416 1351
rect 454 1346 488 1351
rect 598 1339 632 1373
rect 382 1283 416 1307
rect 454 1283 488 1307
rect 526 1300 560 1334
rect 382 1273 404 1283
rect 404 1273 416 1283
rect 454 1273 472 1283
rect 472 1273 488 1283
rect 598 1266 632 1300
rect 382 1212 416 1234
rect 454 1214 488 1234
rect 526 1227 560 1261
rect 382 1200 404 1212
rect 404 1200 416 1212
rect 454 1200 488 1214
rect 598 1193 632 1227
rect 526 1180 560 1188
rect 382 1141 416 1161
rect 382 1127 404 1141
rect 404 1127 416 1141
rect 454 1127 488 1161
rect 526 1154 540 1180
rect 540 1154 560 1180
rect 598 1120 632 1154
rect 526 1112 560 1115
rect 382 1070 416 1088
rect 382 1054 404 1070
rect 404 1054 416 1070
rect 454 1054 488 1088
rect 526 1081 540 1112
rect 540 1081 560 1112
rect 598 1047 632 1081
rect 382 999 416 1015
rect 382 981 404 999
rect 404 981 416 999
rect 454 981 488 1015
rect 526 1010 540 1042
rect 540 1010 560 1042
rect 526 1008 560 1010
rect 598 974 632 1008
rect 526 942 540 969
rect 540 942 560 969
rect 382 928 416 942
rect 382 908 404 928
rect 404 908 416 928
rect 454 908 488 942
rect 526 935 560 942
rect 598 901 632 935
rect 526 874 540 896
rect 540 874 560 896
rect 382 857 416 869
rect 382 835 404 857
rect 404 835 416 857
rect 454 835 488 869
rect 526 862 560 874
rect 598 828 632 862
rect 526 806 540 824
rect 540 806 560 824
rect 382 786 416 796
rect 382 762 404 786
rect 404 762 416 786
rect 454 762 488 796
rect 526 790 560 806
rect 598 755 632 789
rect 526 738 540 752
rect 540 738 560 752
rect 526 724 560 738
rect 382 715 416 723
rect 382 689 404 715
rect 404 689 416 715
rect 454 689 488 723
rect 526 718 540 724
rect 540 718 560 724
rect 798 2176 832 2210
rect 798 2103 832 2137
rect 798 2030 832 2064
rect 798 1958 832 1992
rect 798 1886 832 1920
rect 798 1814 832 1848
rect 798 1742 832 1776
rect 798 1670 832 1704
rect 798 1598 832 1632
rect 798 1526 832 1560
rect 798 1454 832 1488
rect 798 1382 832 1416
rect 798 1310 832 1344
rect 798 1238 832 1272
rect 798 1166 832 1200
rect 798 1094 832 1128
rect 798 1022 832 1056
rect 798 950 832 984
rect 798 878 832 912
rect 798 806 832 840
rect 798 734 832 768
rect 1110 2176 1144 2210
rect 1110 2103 1144 2137
rect 1110 2030 1144 2064
rect 1110 1958 1144 1992
rect 1110 1886 1144 1920
rect 1110 1814 1144 1848
rect 1110 1742 1144 1776
rect 1110 1670 1144 1704
rect 1110 1598 1144 1632
rect 1110 1526 1144 1560
rect 1110 1454 1144 1488
rect 1110 1382 1144 1416
rect 1110 1310 1144 1344
rect 1110 1238 1144 1272
rect 1110 1166 1144 1200
rect 1110 1094 1144 1128
rect 1110 1022 1144 1056
rect 1110 950 1144 984
rect 1110 878 1144 912
rect 1110 806 1144 840
rect 1110 734 1144 768
rect 1626 2176 1660 2210
rect 1626 2103 1660 2137
rect 1626 2030 1660 2064
rect 1626 1958 1660 1992
rect 1626 1886 1660 1920
rect 1626 1814 1660 1848
rect 1626 1742 1660 1776
rect 1626 1670 1660 1704
rect 1626 1598 1660 1632
rect 1626 1526 1660 1560
rect 1626 1454 1660 1488
rect 1626 1382 1660 1416
rect 1626 1310 1660 1344
rect 1626 1238 1660 1272
rect 1626 1166 1660 1200
rect 1626 1094 1660 1128
rect 1626 1022 1660 1056
rect 1626 950 1660 984
rect 1626 878 1660 912
rect 1626 806 1660 840
rect 598 682 632 716
rect 382 644 416 650
rect 382 616 404 644
rect 404 616 416 644
rect 454 616 488 650
rect 526 646 540 680
rect 540 646 560 680
rect 598 609 632 643
rect 688 642 703 676
rect 703 642 722 676
rect 764 642 774 676
rect 774 642 798 676
rect 840 642 845 676
rect 845 642 874 676
rect 916 642 917 676
rect 917 642 950 676
rect 992 642 1023 676
rect 1023 642 1026 676
rect 1068 642 1095 676
rect 1095 642 1102 676
rect 1144 642 1167 676
rect 1167 642 1178 676
rect 1221 642 1239 676
rect 1239 642 1255 676
rect 526 574 540 608
rect 540 574 560 608
rect 1626 734 1660 768
rect 1938 2176 1972 2210
rect 1938 2103 1972 2137
rect 1938 2030 1972 2064
rect 1938 1958 1972 1992
rect 1938 1886 1972 1920
rect 1938 1814 1972 1848
rect 1938 1742 1972 1776
rect 1938 1670 1972 1704
rect 1938 1598 1972 1632
rect 1938 1526 1972 1560
rect 1938 1454 1972 1488
rect 1938 1382 1972 1416
rect 1938 1310 1972 1344
rect 1938 1238 1972 1272
rect 1938 1166 1972 1200
rect 1938 1094 1972 1128
rect 1938 1022 1972 1056
rect 1938 950 1972 984
rect 1938 878 1972 912
rect 1938 806 1972 840
rect 1938 734 1972 768
rect 2454 2176 2488 2210
rect 2454 2103 2488 2137
rect 2454 2030 2488 2064
rect 2454 1958 2488 1992
rect 2454 1886 2488 1920
rect 2454 1814 2488 1848
rect 2454 1742 2488 1776
rect 2454 1670 2488 1704
rect 2454 1598 2488 1632
rect 2454 1526 2488 1560
rect 2454 1454 2488 1488
rect 2454 1382 2488 1416
rect 2454 1310 2488 1344
rect 2454 1238 2488 1272
rect 2454 1166 2488 1200
rect 2454 1094 2488 1128
rect 2454 1022 2488 1056
rect 2454 950 2488 984
rect 2454 878 2488 912
rect 2454 806 2488 840
rect 1516 642 1531 676
rect 1531 642 1550 676
rect 1592 642 1602 676
rect 1602 642 1626 676
rect 1668 642 1673 676
rect 1673 642 1702 676
rect 1744 642 1745 676
rect 1745 642 1778 676
rect 1820 642 1851 676
rect 1851 642 1854 676
rect 1896 642 1923 676
rect 1923 642 1930 676
rect 1972 642 1995 676
rect 1995 642 2006 676
rect 2049 642 2067 676
rect 2067 642 2083 676
rect 2454 734 2488 768
rect 2766 2176 2800 2210
rect 2766 2103 2800 2137
rect 2766 2030 2800 2064
rect 2766 1958 2800 1992
rect 2766 1886 2800 1920
rect 2766 1814 2800 1848
rect 2766 1742 2800 1776
rect 2766 1670 2800 1704
rect 2766 1598 2800 1632
rect 2766 1526 2800 1560
rect 2766 1454 2800 1488
rect 2766 1382 2800 1416
rect 2766 1310 2800 1344
rect 2766 1238 2800 1272
rect 2766 1166 2800 1200
rect 2766 1094 2800 1128
rect 2766 1022 2800 1056
rect 2766 950 2800 984
rect 2766 878 2800 912
rect 2766 806 2800 840
rect 2766 734 2800 768
rect 3171 3806 3205 3818
rect 3247 3806 3281 3818
rect 3323 3806 3357 3818
rect 3399 3806 3433 3818
rect 3475 3806 3509 3818
rect 3551 3806 3585 3818
rect 3628 3806 3662 3818
rect 3705 3806 3739 3818
rect 3171 3784 3187 3806
rect 3187 3784 3205 3806
rect 3247 3784 3258 3806
rect 3258 3784 3281 3806
rect 3323 3784 3329 3806
rect 3329 3784 3357 3806
rect 3399 3784 3401 3806
rect 3401 3784 3433 3806
rect 3475 3784 3507 3806
rect 3507 3784 3509 3806
rect 3551 3784 3579 3806
rect 3579 3784 3585 3806
rect 3628 3784 3651 3806
rect 3651 3784 3662 3806
rect 3705 3784 3723 3806
rect 3723 3784 3739 3806
rect 2952 3704 2986 3738
rect 3024 3704 3058 3738
rect 3096 3704 3130 3738
rect 2952 3631 2986 3665
rect 3024 3631 3058 3665
rect 3096 3631 3130 3665
rect 2952 2262 3130 3592
rect 2344 642 2359 676
rect 2359 642 2378 676
rect 2420 642 2430 676
rect 2430 642 2454 676
rect 2496 642 2501 676
rect 2501 642 2530 676
rect 2572 642 2573 676
rect 2573 642 2606 676
rect 2648 642 2679 676
rect 2679 642 2682 676
rect 2724 642 2751 676
rect 2751 642 2758 676
rect 2800 642 2823 676
rect 2823 642 2834 676
rect 2877 642 2895 676
rect 2895 642 2911 676
rect 3998 3806 4032 3818
rect 4074 3806 4108 3818
rect 4150 3806 4184 3818
rect 4226 3806 4260 3818
rect 4302 3806 4336 3818
rect 4379 3806 4413 3818
rect 4456 3806 4490 3818
rect 4533 3806 4567 3818
rect 3998 3784 4014 3806
rect 4014 3784 4032 3806
rect 4074 3784 4085 3806
rect 4085 3784 4108 3806
rect 4150 3784 4157 3806
rect 4157 3784 4184 3806
rect 4226 3784 4229 3806
rect 4229 3784 4260 3806
rect 4302 3784 4335 3806
rect 4335 3784 4336 3806
rect 4379 3784 4407 3806
rect 4407 3784 4413 3806
rect 4456 3784 4479 3806
rect 4479 3784 4490 3806
rect 4533 3784 4551 3806
rect 4551 3784 4567 3806
rect 5522 3856 5542 3890
rect 5542 3856 5556 3890
rect 5450 3821 5484 3855
rect 4827 3806 4861 3818
rect 4903 3806 4937 3818
rect 4979 3806 5013 3818
rect 5055 3806 5089 3818
rect 5131 3806 5165 3818
rect 5207 3806 5241 3818
rect 5284 3806 5318 3818
rect 5361 3806 5395 3818
rect 4827 3784 4843 3806
rect 4843 3784 4861 3806
rect 4903 3784 4914 3806
rect 4914 3784 4937 3806
rect 4979 3784 4985 3806
rect 4985 3784 5013 3806
rect 5055 3784 5057 3806
rect 5057 3784 5089 3806
rect 5131 3784 5163 3806
rect 5163 3784 5165 3806
rect 5207 3784 5235 3806
rect 5235 3784 5241 3806
rect 5284 3784 5307 3806
rect 5307 3784 5318 3806
rect 5361 3784 5379 3806
rect 5379 3784 5395 3806
rect 5450 3748 5484 3782
rect 3438 3704 3472 3738
rect 3438 3631 3472 3665
rect 3438 3558 3472 3592
rect 3438 3486 3472 3520
rect 3438 3414 3472 3448
rect 3438 3342 3472 3376
rect 3438 3270 3472 3304
rect 3438 3198 3472 3232
rect 3438 3126 3472 3160
rect 3438 3054 3472 3088
rect 3438 2982 3472 3016
rect 3438 2910 3472 2944
rect 3438 2838 3472 2872
rect 3438 2766 3472 2800
rect 3438 2694 3472 2728
rect 3438 2622 3472 2656
rect 3438 2550 3472 2584
rect 3438 2478 3472 2512
rect 3438 2406 3472 2440
rect 3438 2334 3472 2368
rect 3438 2262 3472 2296
rect 3781 3704 3815 3738
rect 3853 3704 3887 3738
rect 3925 3704 3959 3738
rect 3781 3631 3815 3665
rect 3853 3631 3887 3665
rect 3925 3631 3959 3665
rect 3781 2262 3959 3592
rect 4266 3704 4300 3738
rect 4266 3631 4300 3665
rect 4266 3558 4300 3592
rect 4266 3486 4300 3520
rect 4266 3414 4300 3448
rect 4266 3342 4300 3376
rect 4266 3270 4300 3304
rect 4266 3198 4300 3232
rect 4266 3126 4300 3160
rect 4266 3054 4300 3088
rect 4266 2982 4300 3016
rect 4266 2910 4300 2944
rect 4266 2838 4300 2872
rect 4266 2766 4300 2800
rect 4266 2694 4300 2728
rect 4266 2622 4300 2656
rect 4266 2550 4300 2584
rect 4266 2478 4300 2512
rect 4266 2406 4300 2440
rect 4266 2334 4300 2368
rect 4266 2262 4300 2296
rect 4608 3704 4642 3738
rect 4680 3704 4714 3738
rect 4752 3704 4786 3738
rect 4608 3631 4642 3665
rect 4680 3631 4714 3665
rect 4752 3631 4786 3665
rect 4608 2262 4786 3592
rect 5094 3704 5128 3738
rect 5094 3631 5128 3665
rect 5094 3558 5128 3592
rect 5094 3486 5128 3520
rect 5094 3414 5128 3448
rect 5094 3342 5128 3376
rect 5094 3270 5128 3304
rect 5094 3198 5128 3232
rect 5094 3126 5128 3160
rect 5094 3054 5128 3088
rect 5094 2982 5128 3016
rect 5094 2910 5128 2944
rect 5094 2838 5128 2872
rect 5094 2766 5128 2800
rect 5094 2694 5128 2728
rect 5094 2622 5128 2656
rect 5094 2550 5128 2584
rect 5094 2478 5128 2512
rect 5094 2406 5128 2440
rect 5094 2334 5128 2368
rect 5094 2262 5128 2296
rect 5450 3675 5484 3709
rect 5522 3692 5542 3850
rect 5542 3692 5700 3850
rect 5522 3658 5576 3692
rect 5576 3658 5700 3692
rect 5450 3602 5484 3636
rect 5522 3624 5542 3658
rect 5542 3624 5700 3658
rect 5522 3590 5576 3624
rect 5576 3590 5700 3624
rect 5522 3568 5542 3590
rect 5542 3568 5700 3590
rect 5450 3529 5484 3563
rect 5522 3522 5556 3529
rect 5522 3495 5542 3522
rect 5542 3495 5556 3522
rect 5450 3456 5484 3490
rect 5522 3454 5556 3456
rect 5522 3422 5542 3454
rect 5542 3422 5556 3454
rect 5450 3383 5484 3417
rect 5522 3352 5542 3383
rect 5542 3352 5556 3383
rect 5522 3349 5556 3352
rect 5450 3310 5484 3344
rect 5522 3284 5542 3310
rect 5542 3284 5556 3310
rect 5522 3276 5556 3284
rect 5450 3237 5484 3271
rect 5522 3216 5542 3237
rect 5542 3216 5556 3237
rect 5522 3203 5556 3216
rect 5450 3164 5484 3198
rect 5522 3148 5542 3164
rect 5542 3148 5556 3164
rect 5522 3130 5556 3148
rect 5450 3091 5484 3125
rect 5522 3080 5542 3091
rect 5542 3080 5556 3091
rect 5522 3057 5556 3080
rect 5450 3018 5484 3052
rect 5522 3012 5542 3018
rect 5542 3012 5556 3018
rect 5522 2984 5556 3012
rect 5450 2945 5484 2979
rect 5594 2952 5700 3568
rect 5522 2944 5542 2945
rect 5542 2944 5556 2945
rect 5522 2911 5556 2944
rect 5450 2872 5484 2906
rect 5594 2879 5628 2913
rect 5666 2879 5700 2913
rect 5522 2842 5556 2872
rect 5522 2838 5542 2842
rect 5542 2838 5556 2842
rect 5450 2799 5484 2833
rect 5594 2806 5628 2840
rect 5666 2806 5700 2840
rect 5522 2774 5556 2799
rect 5522 2765 5542 2774
rect 5542 2765 5556 2774
rect 5450 2726 5484 2760
rect 5594 2733 5628 2767
rect 5666 2733 5700 2767
rect 5522 2706 5556 2726
rect 5522 2692 5542 2706
rect 5542 2692 5556 2706
rect 5450 2653 5484 2687
rect 5594 2660 5628 2694
rect 5666 2660 5700 2694
rect 5522 2619 5556 2653
rect 5450 2580 5484 2614
rect 5594 2587 5610 2621
rect 5610 2587 5628 2621
rect 5666 2587 5700 2621
rect 5522 2546 5556 2580
rect 5450 2507 5484 2541
rect 5594 2535 5628 2548
rect 5666 2536 5678 2548
rect 5678 2536 5700 2548
rect 5594 2514 5610 2535
rect 5610 2514 5628 2535
rect 5666 2514 5700 2536
rect 5522 2473 5556 2507
rect 5450 2434 5484 2468
rect 5594 2466 5628 2475
rect 5666 2467 5678 2475
rect 5678 2467 5700 2475
rect 5594 2441 5610 2466
rect 5610 2441 5628 2466
rect 5666 2441 5700 2467
rect 5522 2400 5556 2434
rect 5594 2397 5628 2402
rect 5666 2398 5678 2402
rect 5678 2398 5700 2402
rect 5450 2361 5484 2395
rect 5594 2368 5610 2397
rect 5610 2368 5628 2397
rect 5666 2368 5700 2398
rect 5522 2327 5556 2361
rect 5594 2328 5628 2329
rect 5450 2288 5484 2322
rect 5594 2295 5610 2328
rect 5610 2295 5628 2328
rect 5666 2295 5700 2329
rect 5522 2254 5556 2288
rect 5450 2215 5484 2249
rect 5594 2225 5610 2256
rect 5610 2225 5628 2256
rect 5666 2225 5700 2256
rect 5594 2222 5628 2225
rect 5666 2222 5678 2225
rect 5678 2222 5700 2225
rect 3282 2176 3316 2210
rect 3282 2103 3316 2137
rect 3282 2030 3316 2064
rect 3282 1958 3316 1992
rect 3282 1886 3316 1920
rect 3282 1814 3316 1848
rect 3282 1742 3316 1776
rect 3282 1670 3316 1704
rect 3282 1598 3316 1632
rect 3282 1526 3316 1560
rect 3282 1454 3316 1488
rect 3282 1382 3316 1416
rect 3282 1310 3316 1344
rect 3282 1238 3316 1272
rect 3282 1166 3316 1200
rect 3282 1094 3316 1128
rect 3282 1022 3316 1056
rect 3282 950 3316 984
rect 3282 878 3316 912
rect 3282 806 3316 840
rect 3282 734 3316 768
rect 3594 2176 3628 2210
rect 3594 2103 3628 2137
rect 3594 2030 3628 2064
rect 3594 1958 3628 1992
rect 3594 1886 3628 1920
rect 3594 1814 3628 1848
rect 3594 1742 3628 1776
rect 3594 1670 3628 1704
rect 3594 1598 3628 1632
rect 3594 1526 3628 1560
rect 3594 1454 3628 1488
rect 3594 1382 3628 1416
rect 3594 1310 3628 1344
rect 3594 1238 3628 1272
rect 3594 1166 3628 1200
rect 3594 1094 3628 1128
rect 3594 1022 3628 1056
rect 3594 950 3628 984
rect 3594 878 3628 912
rect 3594 806 3628 840
rect 3594 734 3628 768
rect 4110 2176 4144 2210
rect 4110 2103 4144 2137
rect 4110 2030 4144 2064
rect 4110 1958 4144 1992
rect 4110 1886 4144 1920
rect 4110 1814 4144 1848
rect 4110 1742 4144 1776
rect 4110 1670 4144 1704
rect 4110 1598 4144 1632
rect 4110 1526 4144 1560
rect 4110 1454 4144 1488
rect 4110 1382 4144 1416
rect 4110 1310 4144 1344
rect 4110 1238 4144 1272
rect 4110 1166 4144 1200
rect 4110 1094 4144 1128
rect 4110 1022 4144 1056
rect 4110 950 4144 984
rect 4110 878 4144 912
rect 4110 806 4144 840
rect 3172 642 3187 676
rect 3187 642 3206 676
rect 3248 642 3258 676
rect 3258 642 3282 676
rect 3324 642 3329 676
rect 3329 642 3358 676
rect 3400 642 3401 676
rect 3401 642 3434 676
rect 3476 642 3507 676
rect 3507 642 3510 676
rect 3552 642 3579 676
rect 3579 642 3586 676
rect 3628 642 3651 676
rect 3651 642 3662 676
rect 3705 642 3723 676
rect 3723 642 3739 676
rect 4110 734 4144 768
rect 4422 2176 4456 2210
rect 4422 2103 4456 2137
rect 4422 2030 4456 2064
rect 4422 1958 4456 1992
rect 4422 1886 4456 1920
rect 4422 1814 4456 1848
rect 4422 1742 4456 1776
rect 4422 1670 4456 1704
rect 4422 1598 4456 1632
rect 4422 1526 4456 1560
rect 4422 1454 4456 1488
rect 4422 1382 4456 1416
rect 4422 1310 4456 1344
rect 4422 1238 4456 1272
rect 4422 1166 4456 1200
rect 4422 1094 4456 1128
rect 4422 1022 4456 1056
rect 4422 950 4456 984
rect 4422 878 4456 912
rect 4422 806 4456 840
rect 4422 734 4456 768
rect 4938 2176 4972 2210
rect 4938 2103 4972 2137
rect 4938 2030 4972 2064
rect 4938 1958 4972 1992
rect 4938 1886 4972 1920
rect 4938 1814 4972 1848
rect 4938 1742 4972 1776
rect 4938 1670 4972 1704
rect 4938 1598 4972 1632
rect 4938 1526 4972 1560
rect 4938 1454 4972 1488
rect 4938 1382 4972 1416
rect 4938 1310 4972 1344
rect 4938 1238 4972 1272
rect 4938 1166 4972 1200
rect 4938 1094 4972 1128
rect 4938 1022 4972 1056
rect 4938 950 4972 984
rect 4938 878 4972 912
rect 4938 806 4972 840
rect 4000 642 4015 676
rect 4015 642 4034 676
rect 4076 642 4086 676
rect 4086 642 4110 676
rect 4152 642 4157 676
rect 4157 642 4186 676
rect 4228 642 4229 676
rect 4229 642 4262 676
rect 4304 642 4335 676
rect 4335 642 4338 676
rect 4380 642 4407 676
rect 4407 642 4414 676
rect 4456 642 4479 676
rect 4479 642 4490 676
rect 4533 642 4551 676
rect 4551 642 4567 676
rect 4938 734 4972 768
rect 5250 2176 5284 2210
rect 5250 2103 5284 2137
rect 5250 2030 5284 2064
rect 5250 1958 5284 1992
rect 5250 1886 5284 1920
rect 5250 1814 5284 1848
rect 5250 1742 5284 1776
rect 5250 1670 5284 1704
rect 5250 1598 5284 1632
rect 5250 1526 5284 1560
rect 5250 1454 5284 1488
rect 5250 1382 5284 1416
rect 5250 1310 5284 1344
rect 5250 1238 5284 1272
rect 5250 1166 5284 1200
rect 5250 1094 5284 1128
rect 5250 1022 5284 1056
rect 5250 950 5284 984
rect 5250 878 5284 912
rect 5250 806 5284 840
rect 5250 734 5284 768
rect 5522 2181 5556 2215
rect 5450 2142 5484 2176
rect 5594 2156 5610 2183
rect 5610 2156 5628 2183
rect 5666 2156 5700 2183
rect 5594 2149 5628 2156
rect 5666 2149 5678 2156
rect 5678 2149 5700 2156
rect 5522 2108 5556 2142
rect 5450 2069 5484 2103
rect 5594 2087 5610 2110
rect 5610 2087 5628 2110
rect 5666 2087 5700 2110
rect 5594 2076 5628 2087
rect 5666 2076 5678 2087
rect 5678 2076 5700 2087
rect 5522 2035 5556 2069
rect 5450 1996 5484 2030
rect 5594 2018 5610 2037
rect 5610 2018 5628 2037
rect 5666 2018 5700 2037
rect 5594 2003 5628 2018
rect 5666 2003 5678 2018
rect 5678 2003 5700 2018
rect 5522 1962 5556 1996
rect 5450 1923 5484 1957
rect 5594 1949 5610 1964
rect 5610 1949 5628 1964
rect 5666 1949 5700 1964
rect 5594 1930 5628 1949
rect 5666 1930 5678 1949
rect 5678 1930 5700 1949
rect 5522 1889 5556 1923
rect 5450 1850 5484 1884
rect 5594 1880 5610 1891
rect 5610 1880 5628 1891
rect 5666 1880 5700 1891
rect 5594 1857 5628 1880
rect 5666 1857 5678 1880
rect 5678 1857 5700 1880
rect 5522 1816 5556 1850
rect 5594 1811 5610 1818
rect 5610 1811 5628 1818
rect 5666 1811 5700 1818
rect 5450 1777 5484 1811
rect 5594 1784 5628 1811
rect 5666 1784 5678 1811
rect 5678 1784 5700 1811
rect 5522 1743 5556 1777
rect 5594 1742 5610 1745
rect 5610 1742 5628 1745
rect 5666 1742 5700 1745
rect 5450 1704 5484 1738
rect 5594 1711 5628 1742
rect 5666 1711 5678 1742
rect 5678 1711 5700 1742
rect 5522 1670 5556 1704
rect 5450 1631 5484 1665
rect 5594 1638 5628 1672
rect 5666 1639 5678 1672
rect 5678 1639 5700 1672
rect 5666 1638 5700 1639
rect 5522 1597 5556 1631
rect 5450 1558 5484 1592
rect 5594 1569 5628 1599
rect 5666 1570 5678 1599
rect 5678 1570 5700 1599
rect 5594 1565 5610 1569
rect 5610 1565 5628 1569
rect 5666 1565 5700 1570
rect 5522 1524 5556 1558
rect 5450 1485 5484 1519
rect 5594 1500 5628 1526
rect 5666 1501 5678 1526
rect 5678 1501 5700 1526
rect 5594 1492 5610 1500
rect 5610 1492 5628 1500
rect 5666 1492 5700 1501
rect 5522 1451 5556 1485
rect 5450 1412 5484 1446
rect 5594 1431 5628 1453
rect 5666 1432 5678 1453
rect 5678 1432 5700 1453
rect 5594 1419 5610 1431
rect 5610 1419 5628 1431
rect 5666 1419 5700 1432
rect 5522 1378 5556 1412
rect 5450 1339 5484 1373
rect 5594 1362 5628 1380
rect 5666 1363 5678 1380
rect 5678 1363 5700 1380
rect 5594 1346 5610 1362
rect 5610 1346 5628 1362
rect 5666 1346 5700 1363
rect 5522 1305 5556 1339
rect 5450 1266 5484 1300
rect 5594 1293 5628 1307
rect 5666 1294 5678 1307
rect 5678 1294 5700 1307
rect 5594 1273 5610 1293
rect 5610 1273 5628 1293
rect 5666 1273 5700 1294
rect 5522 1232 5556 1266
rect 5450 1193 5484 1227
rect 5594 1224 5628 1234
rect 5666 1225 5678 1234
rect 5678 1225 5700 1234
rect 5594 1200 5610 1224
rect 5610 1200 5628 1224
rect 5666 1200 5700 1225
rect 5522 1159 5556 1193
rect 5594 1155 5628 1161
rect 5666 1156 5678 1161
rect 5678 1156 5700 1161
rect 5450 1120 5484 1154
rect 5594 1127 5610 1155
rect 5610 1127 5628 1155
rect 5666 1127 5700 1156
rect 5522 1086 5556 1120
rect 5594 1086 5628 1088
rect 5666 1087 5678 1088
rect 5678 1087 5700 1088
rect 5450 1047 5484 1081
rect 5594 1054 5610 1086
rect 5610 1054 5628 1086
rect 5666 1054 5700 1087
rect 5522 1013 5556 1047
rect 5450 974 5484 1008
rect 5594 983 5610 1015
rect 5610 983 5628 1015
rect 5666 983 5700 1015
rect 5594 981 5628 983
rect 5666 981 5678 983
rect 5678 981 5700 983
rect 5522 940 5556 974
rect 5450 901 5484 935
rect 5594 914 5610 942
rect 5610 914 5628 942
rect 5666 914 5700 942
rect 5594 908 5628 914
rect 5666 908 5678 914
rect 5678 908 5700 914
rect 5522 867 5556 901
rect 5450 828 5484 862
rect 5594 845 5610 869
rect 5610 845 5628 869
rect 5666 845 5700 869
rect 5594 835 5628 845
rect 5666 835 5678 845
rect 5678 835 5700 845
rect 5522 794 5556 828
rect 5450 755 5484 789
rect 5594 776 5610 796
rect 5610 776 5628 796
rect 5666 776 5700 796
rect 5594 762 5628 776
rect 5666 762 5678 776
rect 5678 762 5700 776
rect 5522 724 5556 755
rect 5522 721 5542 724
rect 5542 721 5556 724
rect 5450 682 5484 716
rect 5594 707 5610 723
rect 5610 707 5628 723
rect 5666 707 5700 723
rect 5594 689 5628 707
rect 5666 689 5678 707
rect 5678 689 5700 707
rect 4828 642 4843 676
rect 4843 642 4862 676
rect 4904 642 4914 676
rect 4914 642 4938 676
rect 4980 642 4985 676
rect 4985 642 5014 676
rect 5056 642 5057 676
rect 5057 642 5090 676
rect 5132 642 5163 676
rect 5163 642 5166 676
rect 5208 642 5235 676
rect 5235 642 5242 676
rect 5284 642 5307 676
rect 5307 642 5318 676
rect 5361 642 5379 676
rect 5379 642 5395 676
rect 5522 671 5556 682
rect 5522 648 5542 671
rect 5542 648 5556 671
rect 5450 609 5484 643
rect 5594 638 5610 650
rect 5610 638 5628 650
rect 5666 638 5700 650
rect 5594 616 5628 638
rect 5666 616 5678 638
rect 5678 616 5700 638
rect 5522 602 5556 609
rect 5522 575 5556 602
rect 598 568 609 570
rect 609 568 632 570
rect 671 568 678 570
rect 678 568 705 570
rect 744 568 747 570
rect 747 568 778 570
rect 598 536 632 568
rect 671 536 705 568
rect 744 536 778 568
rect 817 536 851 570
rect 890 536 924 570
rect 963 536 997 570
rect 1036 536 1070 570
rect 1109 536 1143 570
rect 1182 536 1216 570
rect 1255 536 1289 570
rect 1328 536 1362 570
rect 1401 536 1435 570
rect 1474 536 1508 570
rect 1547 536 1581 570
rect 1620 536 1654 570
rect 1693 536 1727 570
rect 1766 536 1800 570
rect 1839 536 1873 570
rect 1912 536 1946 570
rect 1985 536 2019 570
rect 2058 536 2092 570
rect 2131 536 2165 570
rect 2204 536 2238 570
rect 2277 536 2311 570
rect 2350 536 2384 570
rect 2423 536 2457 570
rect 2496 536 2530 570
rect 2569 536 2603 570
rect 564 466 598 498
rect 637 466 671 498
rect 710 466 714 498
rect 714 466 744 498
rect 564 464 576 466
rect 576 464 598 466
rect 637 464 645 466
rect 645 464 671 466
rect 710 464 744 466
rect 783 464 817 498
rect 856 464 890 498
rect 929 464 963 498
rect 1002 464 1036 498
rect 1075 464 1109 498
rect 1148 464 1182 498
rect 1221 464 1255 498
rect 1294 464 1328 498
rect 1367 464 1401 498
rect 1440 464 1474 498
rect 1513 464 1547 498
rect 1586 464 1620 498
rect 1659 464 1693 498
rect 1732 464 1766 498
rect 1805 464 1839 498
rect 1878 464 1912 498
rect 1951 464 1985 498
rect 2024 464 2058 498
rect 2097 464 2131 498
rect 2170 464 2204 498
rect 2243 464 2277 498
rect 2316 464 2350 498
rect 2388 464 2422 498
rect 2460 464 2494 498
rect 2532 464 2566 498
rect 2604 464 2638 498
rect 2642 464 5446 570
rect 5450 536 5484 570
rect 5522 502 5556 536
rect 5980 4218 6086 4548
rect 5980 4145 6014 4179
rect 6052 4146 6086 4180
rect 5980 4072 6014 4106
rect 6052 4074 6086 4108
rect 5980 3999 6014 4033
rect 6052 4002 6086 4036
rect 5980 3926 6014 3960
rect 6052 3930 6086 3964
rect 5980 3853 6014 3887
rect 6052 3858 6086 3892
rect 5980 3780 6014 3814
rect 6052 3786 6086 3820
rect 5980 3707 6014 3741
rect 6052 3714 6086 3748
rect 5980 3634 6014 3668
rect 6052 3642 6086 3676
rect 5980 3561 6014 3595
rect 6052 3570 6086 3604
rect 5980 3488 6014 3522
rect 6052 3498 6086 3532
rect 5980 3415 6014 3449
rect 6052 3426 6086 3460
rect 5980 3342 6014 3376
rect 6052 3354 6086 3388
rect 5980 3269 6014 3303
rect 6052 3282 6086 3316
rect 5980 3196 6014 3230
rect 6052 3210 6086 3244
rect 5980 3123 6014 3157
rect 6052 3138 6086 3172
rect 5980 3050 6014 3084
rect 6052 3066 6086 3100
rect 5980 2977 6014 3011
rect 6052 2994 6086 3028
rect 5980 2904 6014 2938
rect 6052 2922 6086 2956
rect 5980 2831 6014 2865
rect 6052 2850 6086 2884
rect 5980 2758 6014 2792
rect 6052 2778 6086 2812
rect 5980 2685 6014 2719
rect 6052 2706 6086 2740
rect 5980 2612 6014 2646
rect 6052 2634 6086 2668
rect 5980 2539 6014 2573
rect 6052 2562 6086 2596
rect 5980 2466 6014 2500
rect 6052 2490 6086 2524
rect 5980 2393 6014 2427
rect 6052 2418 6086 2452
rect 5980 2320 6014 2354
rect 6052 2346 6086 2380
rect 5980 2247 6014 2281
rect 6052 2274 6086 2308
rect 5980 2174 6014 2208
rect 6052 2202 6086 2236
rect 5980 2101 6014 2135
rect 6052 2130 6086 2164
rect 5980 2028 6014 2062
rect 6052 2058 6086 2092
rect 5980 1955 6014 1989
rect 6052 1986 6086 2020
rect 5980 1882 6014 1916
rect 6052 1914 6086 1948
rect 5980 1809 6014 1843
rect 6052 1842 6086 1876
rect 6052 1770 6086 1804
rect 5980 1736 6014 1770
rect 6052 1698 6086 1732
rect 5980 1663 6014 1697
rect 6052 1626 6086 1660
rect 5980 1590 6014 1624
rect 6052 1554 6086 1588
rect 5980 1517 6014 1551
rect 6052 1482 6086 1516
rect 5980 1444 6014 1478
rect 6052 1410 6086 1444
rect 5980 1371 6014 1405
rect 6052 1337 6086 1371
rect 5980 1298 6014 1332
rect 6052 1264 6086 1298
rect 5980 1225 6014 1259
rect 6052 1191 6086 1225
rect 5980 1152 6014 1186
rect 6052 1118 6086 1152
rect 5980 1079 6014 1113
rect 6052 1045 6086 1079
rect 5980 1006 6014 1040
rect 6052 972 6086 1006
rect 5980 933 6014 967
rect 6052 899 6086 933
rect 5980 860 6014 894
rect 6052 826 6086 860
rect 5980 787 6014 821
rect 6052 753 6086 787
rect 5980 714 6014 748
rect 6052 680 6086 714
rect 5980 641 6014 675
rect 6052 607 6086 641
rect 5980 568 6014 602
rect 6052 534 6086 568
rect 5980 495 6014 529
rect 6052 461 6086 495
rect 5980 422 6014 456
rect 6052 388 6086 422
rect 5980 349 6014 383
rect 6052 315 6086 349
rect 5980 276 6014 310
rect 6052 242 6086 276
rect 5980 203 6014 237
rect 6052 169 6086 203
rect 174 130 204 164
rect 204 130 208 164
rect 247 130 281 164
rect 320 130 354 164
rect 393 130 427 164
rect 466 130 500 164
rect 539 130 573 164
rect 612 130 646 164
rect 685 130 719 164
rect 758 130 792 164
rect 831 130 865 164
rect 904 130 938 164
rect 977 130 1011 164
rect 1050 130 1084 164
rect 1123 130 1157 164
rect 1196 130 1230 164
rect 1269 130 1303 164
rect 1342 130 1376 164
rect 1415 130 1449 164
rect 1488 130 1522 164
rect 1561 130 1595 164
rect 1634 130 1668 164
rect 1707 130 1741 164
rect 1780 130 1814 164
rect 1853 130 1887 164
rect 1926 130 1960 164
rect 1999 130 2033 164
rect 2072 130 2106 164
rect 2145 130 2179 164
rect 2218 130 2252 164
rect 2291 130 2325 164
rect 2364 130 2398 164
rect 2437 130 2471 164
rect 2510 130 2544 164
rect 2583 130 2617 164
rect 2656 130 2690 164
rect 2729 130 2763 164
rect 2802 130 2836 164
rect 2875 130 2909 164
rect 2948 130 2982 164
rect 3021 130 3055 164
rect 3094 130 3128 164
rect 3167 130 3201 164
rect 3240 130 3274 164
rect 3313 130 3347 164
rect 3386 130 3420 164
rect 3459 130 3493 164
rect 3532 128 5882 164
rect 5882 162 5948 164
rect 5948 162 5976 164
rect 5980 162 6014 164
rect 5882 128 5976 162
rect 5980 130 6014 162
rect 174 58 204 92
rect 204 58 208 92
rect 247 58 281 92
rect 320 58 354 92
rect 393 58 427 92
rect 466 58 500 92
rect 539 58 573 92
rect 612 58 646 92
rect 685 58 719 92
rect 758 58 792 92
rect 830 58 864 92
rect 902 58 936 92
rect 974 58 1008 92
rect 1046 58 1080 92
rect 1118 58 1152 92
rect 1190 58 1224 92
rect 1262 58 1296 92
rect 1334 58 1368 92
rect 1406 58 1440 92
rect 1478 58 1512 92
rect 1550 58 1584 92
rect 1622 58 1656 92
rect 1694 58 1728 92
rect 1766 58 1800 92
rect 1838 58 1872 92
rect 1910 58 1944 92
rect 1982 58 2016 92
rect 2054 58 2088 92
rect 2126 58 2160 92
rect 2198 58 2232 92
rect 2270 58 2304 92
rect 2342 58 2376 92
rect 2414 58 2448 92
rect 2486 58 2520 92
rect 2558 58 2592 92
rect 2630 58 2664 92
rect 2702 58 2736 92
rect 2774 58 2808 92
rect 2846 58 2880 92
rect 2918 58 2952 92
rect 2990 58 3024 92
rect 3062 58 3096 92
rect 3134 58 3168 92
rect 3206 58 3240 92
rect 3278 58 3312 92
rect 3350 58 3384 92
rect 3422 58 3456 92
rect 3494 58 3528 92
rect 3532 58 5950 128
rect 5950 58 5976 128
rect 6052 96 6086 130
<< metal1 >>
tri 21 4740 45 4764 se
rect 45 4740 234 4764
tri 234 4740 258 4764 sw
tri 5936 4740 5960 4764 se
rect 5960 4740 6117 4764
tri 15 4734 21 4740 se
rect 21 4734 6117 4740
rect 15 4700 209 4734
rect 243 4700 282 4734
rect 316 4700 355 4734
rect 389 4700 428 4734
rect 462 4700 501 4734
rect 535 4700 574 4734
rect 608 4700 647 4734
rect 681 4700 720 4734
rect 754 4700 793 4734
rect 827 4700 866 4734
rect 900 4700 939 4734
rect 973 4700 1012 4734
rect 1046 4700 1085 4734
rect 1119 4700 1158 4734
rect 1192 4700 1231 4734
rect 1265 4700 1304 4734
rect 1338 4700 1377 4734
rect 1411 4700 1450 4734
rect 1484 4700 1523 4734
rect 1557 4700 1596 4734
rect 1630 4700 1669 4734
rect 1703 4700 1742 4734
rect 1776 4700 1815 4734
rect 1849 4700 1888 4734
rect 1922 4700 1961 4734
rect 1995 4700 2034 4734
rect 2068 4700 2107 4734
rect 2141 4700 2180 4734
rect 2214 4700 2253 4734
rect 2287 4700 2326 4734
rect 2360 4700 2399 4734
rect 2433 4700 2472 4734
rect 2506 4700 2545 4734
rect 2579 4700 2618 4734
rect 2652 4700 2691 4734
rect 2725 4700 2764 4734
rect 2798 4700 2837 4734
rect 2871 4700 2910 4734
rect 2944 4700 2983 4734
rect 3017 4700 3056 4734
rect 3090 4700 3129 4734
rect 3163 4700 3202 4734
rect 3236 4700 3275 4734
rect 3309 4700 3348 4734
rect 3382 4700 3421 4734
rect 3455 4700 3494 4734
rect 3528 4700 3567 4734
rect 3601 4700 3640 4734
rect 3674 4700 3713 4734
rect 3747 4700 3786 4734
rect 3820 4700 3859 4734
rect 3893 4700 3932 4734
rect 3966 4700 4005 4734
rect 4039 4700 4078 4734
rect 4112 4700 4151 4734
rect 4185 4700 4224 4734
rect 4258 4700 4297 4734
rect 4331 4700 4370 4734
rect 4404 4700 4443 4734
rect 4477 4700 4516 4734
rect 4550 4700 4589 4734
rect 4623 4700 4662 4734
rect 4696 4700 4735 4734
rect 4769 4700 4808 4734
rect 4842 4700 4881 4734
rect 4915 4700 4954 4734
rect 15 4662 4954 4700
rect 15 4628 209 4662
rect 243 4628 282 4662
rect 316 4628 355 4662
rect 389 4628 428 4662
rect 462 4628 501 4662
rect 535 4628 574 4662
rect 608 4628 647 4662
rect 681 4628 720 4662
rect 754 4628 793 4662
rect 827 4628 866 4662
rect 900 4628 939 4662
rect 973 4628 1012 4662
rect 1046 4628 1085 4662
rect 1119 4628 1158 4662
rect 1192 4628 1231 4662
rect 1265 4628 1304 4662
rect 1338 4628 1377 4662
rect 1411 4628 1450 4662
rect 1484 4628 1523 4662
rect 1557 4628 1596 4662
rect 1630 4628 1669 4662
rect 1703 4628 1742 4662
rect 1776 4628 1815 4662
rect 1849 4628 1888 4662
rect 1922 4628 1961 4662
rect 1995 4628 2034 4662
rect 2068 4628 2107 4662
rect 2141 4628 2180 4662
rect 2214 4628 2253 4662
rect 2287 4628 2326 4662
rect 2360 4628 2399 4662
rect 2433 4628 2472 4662
rect 2506 4628 2545 4662
rect 2579 4628 2618 4662
rect 2652 4628 2691 4662
rect 2725 4628 2764 4662
rect 2798 4628 2837 4662
rect 2871 4628 2910 4662
rect 2944 4628 2983 4662
rect 3017 4628 3056 4662
rect 3090 4628 3129 4662
rect 3163 4628 3202 4662
rect 3236 4628 3275 4662
rect 3309 4628 3348 4662
rect 3382 4628 3421 4662
rect 3455 4628 3494 4662
rect 3528 4628 3567 4662
rect 3601 4628 3640 4662
rect 3674 4628 3713 4662
rect 3747 4628 3786 4662
rect 3820 4628 3859 4662
rect 3893 4628 3932 4662
rect 3966 4628 4005 4662
rect 4039 4628 4078 4662
rect 4112 4628 4151 4662
rect 4185 4628 4224 4662
rect 4258 4628 4297 4662
rect 4331 4628 4370 4662
rect 4404 4628 4443 4662
rect 4477 4628 4516 4662
rect 4550 4628 4589 4662
rect 4623 4628 4662 4662
rect 4696 4628 4735 4662
rect 4769 4628 4808 4662
rect 4842 4628 4881 4662
rect 4915 4628 4954 4662
rect 5924 4646 6117 4734
rect 5924 4628 6095 4646
rect 15 4624 6095 4628
tri 6095 4624 6117 4646 nw
rect 15 4622 6092 4624
rect 15 4612 208 4622
tri 208 4612 218 4622 nw
tri 5949 4612 5959 4622 ne
rect 5959 4612 6092 4622
tri 6092 4621 6095 4624 nw
rect 15 4603 199 4612
tri 199 4603 208 4612 nw
tri 5959 4603 5968 4612 ne
rect 5968 4603 5980 4612
tri 39 4597 45 4603 ne
rect 45 4597 193 4603
tri 193 4597 199 4603 nw
tri 5968 4597 5974 4603 ne
tri 45 4554 88 4597 ne
rect 88 4554 150 4597
tri 150 4554 193 4597 nw
rect 370 4288 5712 4294
rect 370 4254 382 4288
rect 416 4254 455 4288
rect 489 4254 528 4288
rect 562 4254 601 4288
rect 635 4254 674 4288
rect 708 4254 747 4288
rect 781 4254 820 4288
rect 854 4254 893 4288
rect 927 4254 966 4288
rect 1000 4254 1039 4288
rect 1073 4254 1112 4288
rect 1146 4254 1185 4288
rect 1219 4254 1258 4288
rect 1292 4254 1331 4288
rect 1365 4254 1404 4288
rect 1438 4254 1477 4288
rect 1511 4254 1550 4288
rect 1584 4254 1623 4288
rect 1657 4254 1696 4288
rect 1730 4254 1769 4288
rect 1803 4254 1842 4288
rect 1876 4254 1915 4288
rect 1949 4254 1988 4288
rect 2022 4254 2061 4288
rect 2095 4254 2134 4288
rect 2168 4254 2207 4288
rect 2241 4254 2280 4288
rect 2314 4254 2353 4288
rect 2387 4254 2426 4288
rect 370 4216 2426 4254
rect 370 4182 382 4216
rect 416 4182 455 4216
rect 489 4182 528 4216
rect 562 4182 601 4216
rect 635 4182 674 4216
rect 708 4182 747 4216
rect 781 4182 820 4216
rect 854 4182 893 4216
rect 927 4182 966 4216
rect 1000 4182 1039 4216
rect 1073 4182 1112 4216
rect 1146 4182 1185 4216
rect 1219 4182 1258 4216
rect 1292 4182 1331 4216
rect 1365 4182 1404 4216
rect 1438 4182 1477 4216
rect 1511 4182 1550 4216
rect 1584 4182 1623 4216
rect 1657 4182 1696 4216
rect 1730 4182 1769 4216
rect 1803 4182 1842 4216
rect 1876 4182 1915 4216
rect 1949 4182 1988 4216
rect 2022 4182 2061 4216
rect 2095 4182 2134 4216
rect 2168 4182 2207 4216
rect 2241 4182 2280 4216
rect 2314 4182 2353 4216
rect 2387 4182 2426 4216
rect 370 4144 2426 4182
rect 370 4110 382 4144
rect 416 4110 455 4144
rect 489 4110 528 4144
rect 562 4110 601 4144
rect 635 4110 674 4144
rect 708 4110 747 4144
rect 781 4110 820 4144
rect 854 4110 893 4144
rect 927 4110 966 4144
rect 1000 4110 1039 4144
rect 1073 4110 1112 4144
rect 1146 4110 1185 4144
rect 1219 4110 1258 4144
rect 1292 4110 1331 4144
rect 1365 4110 1404 4144
rect 1438 4110 1477 4144
rect 1511 4110 1550 4144
rect 1584 4110 1623 4144
rect 1657 4110 1696 4144
rect 1730 4110 1769 4144
rect 1803 4110 1842 4144
rect 1876 4110 1915 4144
rect 1949 4110 1988 4144
rect 2022 4110 2061 4144
rect 2095 4110 2134 4144
rect 2168 4110 2207 4144
rect 2241 4110 2280 4144
rect 2314 4110 2353 4144
rect 2387 4110 2426 4144
rect 370 4072 2426 4110
rect 370 4038 382 4072
rect 416 4038 455 4072
rect 489 4038 528 4072
rect 562 4038 601 4072
rect 635 4038 674 4072
rect 708 4038 747 4072
rect 781 4038 820 4072
rect 854 4038 893 4072
rect 927 4038 966 4072
rect 1000 4038 1039 4072
rect 1073 4038 1112 4072
rect 1146 4038 1185 4072
rect 1219 4038 1258 4072
rect 1292 4038 1331 4072
rect 1365 4038 1404 4072
rect 1438 4038 1477 4072
rect 1511 4038 1550 4072
rect 1584 4038 1623 4072
rect 1657 4038 1696 4072
rect 1730 4038 1769 4072
rect 1803 4038 1842 4072
rect 1876 4038 1915 4072
rect 1949 4038 1988 4072
rect 2022 4038 2061 4072
rect 2095 4038 2134 4072
rect 2168 4038 2207 4072
rect 2241 4038 2280 4072
rect 2314 4038 2353 4072
rect 2387 4038 2426 4072
rect 5700 4038 5712 4288
rect 370 4000 2426 4038
rect 370 3966 636 4000
rect 670 3966 708 4000
rect 742 3966 780 4000
rect 814 3966 852 4000
rect 886 3966 924 4000
rect 958 3966 996 4000
rect 1030 3966 1068 4000
rect 1102 3966 1140 4000
rect 1174 3966 1212 4000
rect 1246 3966 1284 4000
rect 1318 3966 1356 4000
rect 1390 3966 1428 4000
rect 1462 3966 1500 4000
rect 1534 3966 1572 4000
rect 1606 3966 1644 4000
rect 1678 3966 1716 4000
rect 1750 3966 1788 4000
rect 1822 3966 1860 4000
rect 1894 3966 1932 4000
rect 1966 3966 2004 4000
rect 2038 3966 2076 4000
rect 2110 3966 2148 4000
rect 2182 3966 2220 4000
rect 2254 3966 2292 4000
rect 2326 3966 2364 4000
rect 2398 3966 2426 4000
rect 3334 4000 5125 4038
rect 3334 3966 3373 4000
rect 3407 3966 3446 4000
rect 3480 3966 3519 4000
rect 3553 3966 3592 4000
rect 3626 3966 3665 4000
rect 3699 3966 3738 4000
rect 3772 3966 3811 4000
rect 3845 3966 3884 4000
rect 3918 3966 3957 4000
rect 3991 3966 4030 4000
rect 4064 3966 4103 4000
rect 4137 3966 4176 4000
rect 4210 3966 4249 4000
rect 4283 3966 4322 4000
rect 4356 3966 4395 4000
rect 4429 3966 4468 4000
rect 4502 3966 4541 4000
rect 4575 3966 4614 4000
rect 4648 3966 4687 4000
rect 4721 3966 4760 4000
rect 4794 3966 4833 4000
rect 4867 3966 4906 4000
rect 4940 3966 4979 4000
rect 5013 3966 5052 4000
rect 5086 3966 5125 4000
rect 370 3962 5125 3966
rect 370 3928 526 3962
rect 560 3928 5125 3962
rect 370 3894 598 3928
rect 632 3894 671 3928
rect 705 3894 744 3928
rect 778 3894 817 3928
rect 851 3894 890 3928
rect 924 3894 963 3928
rect 997 3894 1036 3928
rect 1070 3894 1109 3928
rect 1143 3894 1182 3928
rect 1216 3894 1255 3928
rect 1289 3894 1328 3928
rect 1362 3894 1401 3928
rect 1435 3894 1474 3928
rect 1508 3894 1547 3928
rect 1581 3894 1620 3928
rect 1654 3894 1693 3928
rect 1727 3894 1766 3928
rect 1800 3894 1839 3928
rect 1873 3894 1912 3928
rect 1946 3894 1985 3928
rect 2019 3894 2058 3928
rect 2092 3894 2131 3928
rect 2165 3894 2204 3928
rect 2238 3894 2277 3928
rect 2311 3894 2350 3928
rect 2384 3894 2423 3928
rect 2457 3894 2496 3928
rect 2530 3894 2569 3928
rect 2603 3894 2642 3928
rect 2676 3894 2715 3928
rect 2749 3894 2788 3928
rect 2822 3894 2861 3928
rect 2895 3894 2934 3928
rect 2968 3894 3007 3928
rect 3041 3894 3080 3928
rect 3114 3894 3153 3928
rect 3187 3894 3226 3928
rect 3260 3894 3299 3928
rect 3333 3894 3372 3928
rect 3406 3894 3445 3928
rect 3479 3894 3518 3928
rect 3552 3894 3591 3928
rect 3625 3894 3664 3928
rect 3698 3894 3737 3928
rect 3771 3894 3810 3928
rect 3844 3894 3883 3928
rect 3917 3894 3956 3928
rect 3990 3894 4029 3928
rect 4063 3894 4102 3928
rect 4136 3894 4175 3928
rect 4209 3894 4248 3928
rect 4282 3894 4321 3928
rect 4355 3894 4394 3928
rect 4428 3894 4467 3928
rect 4501 3894 4540 3928
rect 4574 3894 4613 3928
rect 4647 3894 4686 3928
rect 4720 3894 4759 3928
rect 4793 3894 4832 3928
rect 4866 3894 4905 3928
rect 4939 3894 4978 3928
rect 5012 3894 5051 3928
rect 5085 3894 5125 3928
rect 5231 4000 5712 4038
rect 5231 3966 5292 4000
rect 5326 3966 5388 4000
rect 5422 3966 5484 4000
rect 5518 3966 5712 4000
rect 5231 3928 5712 3966
rect 5231 3894 5281 3928
rect 5315 3894 5365 3928
rect 5399 3894 5450 3928
rect 5484 3894 5712 3928
rect 370 3890 5712 3894
rect 370 3889 5522 3890
rect 370 3855 526 3889
rect 560 3888 5522 3889
rect 560 3855 638 3888
tri 638 3863 663 3888 nw
tri 5419 3863 5444 3888 ne
rect 370 3850 598 3855
rect 370 2952 382 3850
rect 488 3821 598 3850
rect 632 3821 638 3855
rect 5444 3856 5522 3888
rect 5556 3856 5712 3890
rect 5444 3855 5712 3856
rect 488 3816 638 3821
rect 488 3782 526 3816
rect 560 3782 638 3816
rect 488 3748 598 3782
rect 632 3750 638 3782
rect 675 3818 5407 3830
rect 675 3784 687 3818
rect 721 3784 763 3818
rect 797 3784 839 3818
rect 873 3784 915 3818
rect 949 3784 991 3818
rect 1025 3784 1067 3818
rect 1101 3784 1144 3818
rect 1178 3784 1221 3818
rect 1255 3784 1515 3818
rect 1549 3784 1591 3818
rect 1625 3784 1667 3818
rect 1701 3784 1743 3818
rect 1777 3784 1819 3818
rect 1853 3784 1895 3818
rect 1929 3784 1972 3818
rect 2006 3784 2049 3818
rect 2083 3784 2343 3818
rect 2377 3784 2419 3818
rect 2453 3784 2495 3818
rect 2529 3784 2571 3818
rect 2605 3784 2647 3818
rect 2681 3784 2723 3818
rect 2757 3784 2800 3818
rect 2834 3784 2877 3818
rect 2911 3784 3171 3818
rect 3205 3784 3247 3818
rect 3281 3784 3323 3818
rect 3357 3784 3399 3818
rect 3433 3784 3475 3818
rect 3509 3784 3551 3818
rect 3585 3784 3628 3818
rect 3662 3784 3705 3818
rect 3739 3784 3998 3818
rect 4032 3784 4074 3818
rect 4108 3784 4150 3818
rect 4184 3784 4226 3818
rect 4260 3784 4302 3818
rect 4336 3784 4379 3818
rect 4413 3784 4456 3818
rect 4490 3784 4533 3818
rect 4567 3784 4827 3818
rect 4861 3784 4903 3818
rect 4937 3784 4979 3818
rect 5013 3784 5055 3818
rect 5089 3784 5131 3818
rect 5165 3784 5207 3818
rect 5241 3784 5284 3818
rect 5318 3784 5361 3818
rect 5395 3784 5407 3818
rect 675 3778 5407 3784
rect 5444 3821 5450 3855
rect 5484 3850 5712 3855
rect 5484 3821 5522 3850
rect 5444 3782 5522 3821
tri 638 3750 663 3775 sw
tri 5419 3750 5444 3775 se
rect 5444 3750 5450 3782
rect 632 3748 5450 3750
rect 5484 3748 5522 3782
rect 488 3743 5522 3748
rect 488 3709 526 3743
rect 560 3738 5522 3743
rect 560 3709 954 3738
rect 488 3675 598 3709
rect 632 3704 954 3709
rect 988 3704 1297 3738
rect 1331 3704 1369 3738
rect 1403 3704 1441 3738
rect 1475 3704 1782 3738
rect 1816 3704 2124 3738
rect 2158 3704 2196 3738
rect 2230 3704 2268 3738
rect 2302 3704 2610 3738
rect 2644 3704 2952 3738
rect 2986 3704 3024 3738
rect 3058 3704 3096 3738
rect 3130 3704 3438 3738
rect 3472 3704 3781 3738
rect 3815 3704 3853 3738
rect 3887 3704 3925 3738
rect 3959 3704 4266 3738
rect 4300 3704 4608 3738
rect 4642 3704 4680 3738
rect 4714 3704 4752 3738
rect 4786 3704 5094 3738
rect 5128 3709 5522 3738
rect 5128 3704 5450 3709
rect 632 3675 5450 3704
rect 5484 3675 5522 3709
rect 488 3670 5522 3675
rect 488 3636 526 3670
rect 560 3665 5522 3670
rect 560 3636 954 3665
rect 488 3602 598 3636
rect 632 3631 954 3636
rect 988 3631 1297 3665
rect 1331 3631 1369 3665
rect 1403 3631 1441 3665
rect 1475 3631 1782 3665
rect 1816 3631 2124 3665
rect 2158 3631 2196 3665
rect 2230 3631 2268 3665
rect 2302 3631 2610 3665
rect 2644 3631 2952 3665
rect 2986 3631 3024 3665
rect 3058 3631 3096 3665
rect 3130 3631 3438 3665
rect 3472 3631 3781 3665
rect 3815 3631 3853 3665
rect 3887 3631 3925 3665
rect 3959 3631 4266 3665
rect 4300 3631 4608 3665
rect 4642 3631 4680 3665
rect 4714 3631 4752 3665
rect 4786 3631 5094 3665
rect 5128 3636 5522 3665
rect 5128 3631 5450 3636
rect 632 3602 5450 3631
rect 5484 3602 5522 3636
rect 488 3597 5522 3602
rect 488 3563 526 3597
rect 560 3592 5522 3597
rect 560 3570 954 3592
rect 560 3563 651 3570
rect 488 3529 598 3563
rect 632 3558 651 3563
tri 651 3558 663 3570 nw
tri 923 3558 935 3570 ne
rect 935 3558 954 3570
rect 988 3570 1297 3592
rect 988 3558 994 3570
rect 632 3529 638 3558
tri 638 3545 651 3558 nw
tri 935 3545 948 3558 ne
rect 488 3524 638 3529
rect 488 3490 526 3524
rect 560 3490 638 3524
rect 948 3520 994 3558
tri 994 3545 1019 3570 nw
tri 1266 3545 1291 3570 ne
rect 488 3456 598 3490
rect 632 3486 638 3490
tri 638 3486 663 3511 sw
tri 923 3486 948 3511 se
rect 948 3486 954 3520
rect 988 3486 994 3520
tri 994 3486 1019 3511 sw
tri 1266 3486 1291 3511 se
rect 1291 3486 1297 3570
rect 632 3456 1297 3486
rect 488 3451 1297 3456
rect 488 3417 526 3451
rect 560 3448 1297 3451
rect 560 3417 954 3448
rect 488 3383 598 3417
rect 632 3414 954 3417
rect 988 3414 1297 3448
rect 632 3383 1297 3414
rect 488 3378 1297 3383
rect 488 3344 526 3378
rect 560 3376 1297 3378
rect 560 3344 954 3376
rect 488 3310 598 3344
rect 632 3342 954 3344
rect 988 3342 1297 3376
rect 632 3310 1297 3342
rect 488 3306 1297 3310
rect 488 3305 661 3306
rect 488 3271 526 3305
rect 560 3304 661 3305
tri 661 3304 663 3306 nw
tri 923 3304 925 3306 ne
rect 925 3304 994 3306
rect 560 3271 638 3304
tri 638 3281 661 3304 nw
tri 925 3281 948 3304 ne
rect 488 3237 598 3271
rect 632 3237 638 3271
rect 948 3270 954 3304
rect 988 3270 994 3304
tri 994 3281 1019 3306 nw
tri 1266 3281 1291 3306 ne
rect 488 3232 638 3237
tri 638 3232 653 3247 sw
tri 933 3232 948 3247 se
rect 948 3232 994 3270
rect 488 3198 526 3232
rect 560 3222 653 3232
tri 653 3222 663 3232 sw
tri 923 3222 933 3232 se
rect 933 3222 954 3232
rect 560 3198 954 3222
rect 988 3222 994 3232
tri 994 3222 1019 3247 sw
tri 1266 3222 1291 3247 se
rect 1291 3222 1297 3306
rect 988 3198 1297 3222
rect 488 3164 598 3198
rect 632 3164 1297 3198
rect 488 3160 1297 3164
rect 488 3159 954 3160
rect 488 3125 526 3159
rect 560 3126 954 3159
rect 988 3126 1297 3160
rect 560 3125 1297 3126
rect 488 3091 598 3125
rect 632 3091 1297 3125
rect 488 3088 1297 3091
rect 488 3086 954 3088
rect 488 3052 526 3086
rect 560 3054 954 3086
rect 988 3054 1297 3088
rect 560 3052 1297 3054
rect 488 3018 598 3052
rect 632 3042 1297 3052
rect 632 3018 638 3042
rect 488 3013 638 3018
tri 638 3017 663 3042 nw
tri 923 3017 948 3042 ne
rect 488 2979 526 3013
rect 560 2982 638 3013
rect 948 3016 994 3042
tri 994 3017 1019 3042 nw
tri 1266 3017 1291 3042 ne
tri 638 2982 639 2983 sw
tri 947 2982 948 2983 se
rect 948 2982 954 3016
rect 988 2982 994 3016
rect 560 2979 639 2982
rect 488 2952 598 2979
rect 370 2945 598 2952
rect 632 2958 639 2979
tri 639 2958 663 2982 sw
tri 923 2958 947 2982 se
rect 947 2958 994 2982
tri 994 2958 1019 2983 sw
tri 1266 2958 1291 2983 se
rect 1291 2958 1297 3042
rect 632 2945 1297 2958
rect 370 2944 1297 2945
rect 370 2940 954 2944
rect 370 2913 526 2940
rect 370 2879 382 2913
rect 416 2879 454 2913
rect 488 2906 526 2913
rect 560 2910 954 2940
rect 988 2910 1297 2944
rect 560 2906 1297 2910
rect 488 2879 598 2906
rect 370 2872 598 2879
rect 632 2872 1297 2906
rect 370 2867 954 2872
rect 370 2840 526 2867
rect 370 2806 382 2840
rect 416 2806 454 2840
rect 488 2833 526 2840
rect 560 2838 954 2867
rect 988 2838 1297 2872
rect 560 2833 1297 2838
rect 488 2806 598 2833
rect 370 2799 598 2806
rect 632 2800 1297 2833
rect 632 2799 954 2800
rect 370 2794 954 2799
rect 370 2767 526 2794
rect 370 2733 382 2767
rect 416 2733 454 2767
rect 488 2760 526 2767
rect 560 2778 954 2794
rect 560 2766 651 2778
tri 651 2766 663 2778 nw
tri 923 2766 935 2778 ne
rect 935 2766 954 2778
rect 988 2778 1297 2800
rect 988 2766 994 2778
rect 560 2760 638 2766
rect 488 2733 598 2760
rect 370 2726 598 2733
rect 632 2726 638 2760
tri 638 2753 651 2766 nw
tri 935 2753 948 2766 ne
rect 370 2721 638 2726
rect 370 2694 526 2721
rect 370 2660 382 2694
rect 416 2660 454 2694
rect 488 2687 526 2694
rect 560 2694 638 2721
rect 948 2728 994 2766
tri 994 2753 1019 2778 nw
tri 1266 2753 1291 2778 ne
tri 638 2694 663 2719 sw
tri 923 2694 948 2719 se
rect 948 2694 954 2728
rect 988 2694 994 2728
tri 994 2694 1019 2719 sw
tri 1266 2694 1291 2719 se
rect 1291 2694 1297 2778
rect 560 2687 1297 2694
rect 488 2660 598 2687
rect 370 2653 598 2660
rect 632 2656 1297 2687
rect 632 2653 954 2656
rect 370 2648 954 2653
rect 370 2621 526 2648
rect 370 2587 382 2621
rect 416 2587 454 2621
rect 488 2614 526 2621
rect 560 2622 954 2648
rect 988 2622 1297 2656
rect 560 2614 1297 2622
rect 488 2587 598 2614
rect 370 2580 598 2587
rect 632 2584 1297 2614
rect 632 2580 954 2584
rect 370 2575 954 2580
rect 370 2548 526 2575
rect 370 2514 382 2548
rect 416 2514 454 2548
rect 488 2541 526 2548
rect 560 2550 954 2575
rect 988 2550 1297 2584
rect 560 2541 1297 2550
rect 488 2514 598 2541
rect 370 2507 598 2514
rect 632 2514 1297 2541
rect 632 2512 661 2514
tri 661 2512 663 2514 nw
tri 923 2512 925 2514 ne
rect 925 2512 994 2514
rect 632 2507 638 2512
rect 370 2502 638 2507
rect 370 2475 526 2502
rect 370 2441 382 2475
rect 416 2441 454 2475
rect 488 2468 526 2475
rect 560 2468 638 2502
tri 638 2489 661 2512 nw
tri 925 2489 948 2512 ne
rect 488 2441 598 2468
rect 370 2434 598 2441
rect 632 2440 638 2468
rect 948 2478 954 2512
rect 988 2478 994 2512
tri 994 2489 1019 2514 nw
tri 1266 2489 1291 2514 ne
tri 638 2440 653 2455 sw
tri 933 2440 948 2455 se
rect 948 2440 994 2478
rect 632 2434 653 2440
rect 370 2430 653 2434
tri 653 2430 663 2440 sw
tri 923 2430 933 2440 se
rect 933 2430 954 2440
rect 370 2429 954 2430
rect 370 2402 526 2429
rect 370 2368 382 2402
rect 416 2368 454 2402
rect 488 2395 526 2402
rect 560 2406 954 2429
rect 988 2430 994 2440
tri 994 2430 1019 2455 sw
tri 1266 2430 1291 2455 se
rect 1291 2430 1297 2514
rect 988 2406 1297 2430
rect 560 2395 1297 2406
rect 488 2368 598 2395
rect 370 2361 598 2368
rect 632 2368 1297 2395
rect 632 2361 954 2368
rect 370 2356 954 2361
rect 370 2329 526 2356
rect 370 2295 382 2329
rect 416 2295 454 2329
rect 488 2322 526 2329
rect 560 2334 954 2356
rect 988 2334 1297 2368
rect 560 2322 1297 2334
rect 488 2295 598 2322
rect 370 2288 598 2295
rect 632 2296 1297 2322
rect 632 2288 954 2296
rect 370 2283 954 2288
rect 370 2256 526 2283
rect 370 2222 382 2256
rect 416 2222 454 2256
rect 488 2249 526 2256
rect 560 2262 954 2283
rect 988 2262 1297 2296
rect 1475 3570 1782 3592
rect 1475 3558 1494 3570
tri 1494 3558 1506 3570 nw
tri 1751 3558 1763 3570 ne
rect 1763 3558 1782 3570
rect 1816 3570 2124 3592
rect 1816 3558 1822 3570
rect 1475 3486 1481 3558
tri 1481 3545 1494 3558 nw
tri 1763 3545 1776 3558 ne
rect 1776 3520 1822 3558
tri 1822 3545 1847 3570 nw
tri 2093 3545 2118 3570 ne
tri 1481 3486 1506 3511 sw
tri 1751 3486 1776 3511 se
rect 1776 3486 1782 3520
rect 1816 3486 1822 3520
tri 1822 3486 1847 3511 sw
tri 2093 3486 2118 3511 se
rect 2118 3486 2124 3570
rect 1475 3448 2124 3486
rect 1475 3414 1782 3448
rect 1816 3414 2124 3448
rect 1475 3376 2124 3414
rect 1475 3342 1782 3376
rect 1816 3342 2124 3376
rect 1475 3306 2124 3342
rect 1475 3304 1504 3306
tri 1504 3304 1506 3306 nw
tri 1751 3304 1753 3306 ne
rect 1753 3304 1822 3306
rect 1475 3232 1481 3304
tri 1481 3281 1504 3304 nw
tri 1753 3281 1776 3304 ne
rect 1776 3270 1782 3304
rect 1816 3270 1822 3304
tri 1822 3281 1847 3306 nw
tri 2093 3281 2118 3306 ne
tri 1481 3232 1496 3247 sw
tri 1761 3232 1776 3247 se
rect 1776 3232 1822 3270
rect 1475 3222 1496 3232
tri 1496 3222 1506 3232 sw
tri 1751 3222 1761 3232 se
rect 1761 3222 1782 3232
rect 1475 3198 1782 3222
rect 1816 3222 1822 3232
tri 1822 3222 1847 3247 sw
tri 2093 3222 2118 3247 se
rect 2118 3222 2124 3306
rect 1816 3198 2124 3222
rect 1475 3160 2124 3198
rect 1475 3126 1782 3160
rect 1816 3126 2124 3160
rect 1475 3088 2124 3126
rect 1475 3054 1782 3088
rect 1816 3054 2124 3088
rect 1475 3042 2124 3054
rect 1475 2982 1481 3042
tri 1481 3017 1506 3042 nw
tri 1751 3017 1776 3042 ne
rect 1776 3016 1822 3042
tri 1822 3017 1847 3042 nw
tri 2093 3017 2118 3042 ne
tri 1481 2982 1482 2983 sw
tri 1775 2982 1776 2983 se
rect 1776 2982 1782 3016
rect 1816 2982 1822 3016
rect 1475 2958 1482 2982
tri 1482 2958 1506 2982 sw
tri 1751 2958 1775 2982 se
rect 1775 2958 1822 2982
tri 1822 2958 1847 2983 sw
tri 2093 2958 2118 2983 se
rect 2118 2958 2124 3042
rect 1475 2944 2124 2958
rect 1475 2910 1782 2944
rect 1816 2910 2124 2944
rect 1475 2872 2124 2910
rect 1475 2838 1782 2872
rect 1816 2838 2124 2872
rect 1475 2800 2124 2838
rect 1475 2778 1782 2800
rect 1475 2766 1494 2778
tri 1494 2766 1506 2778 nw
tri 1751 2766 1763 2778 ne
rect 1763 2766 1782 2778
rect 1816 2778 2124 2800
rect 1816 2766 1822 2778
rect 1475 2694 1481 2766
tri 1481 2753 1494 2766 nw
tri 1763 2753 1776 2766 ne
rect 1776 2728 1822 2766
tri 1822 2753 1847 2778 nw
tri 2093 2753 2118 2778 ne
tri 1481 2694 1506 2719 sw
tri 1751 2694 1776 2719 se
rect 1776 2694 1782 2728
rect 1816 2694 1822 2728
tri 1822 2694 1847 2719 sw
tri 2093 2694 2118 2719 se
rect 2118 2694 2124 2778
rect 1475 2656 2124 2694
rect 1475 2622 1782 2656
rect 1816 2622 2124 2656
rect 1475 2584 2124 2622
rect 1475 2550 1782 2584
rect 1816 2550 2124 2584
rect 1475 2514 2124 2550
rect 1475 2512 1504 2514
tri 1504 2512 1506 2514 nw
tri 1751 2512 1753 2514 ne
rect 1753 2512 1822 2514
rect 1475 2440 1481 2512
tri 1481 2489 1504 2512 nw
tri 1753 2489 1776 2512 ne
rect 1776 2478 1782 2512
rect 1816 2478 1822 2512
tri 1822 2489 1847 2514 nw
tri 2093 2489 2118 2514 ne
tri 1481 2440 1496 2455 sw
tri 1761 2440 1776 2455 se
rect 1776 2440 1822 2478
rect 1475 2430 1496 2440
tri 1496 2430 1506 2440 sw
tri 1751 2430 1761 2440 se
rect 1761 2430 1782 2440
rect 1475 2406 1782 2430
rect 1816 2430 1822 2440
tri 1822 2430 1847 2455 sw
tri 2093 2430 2118 2455 se
rect 2118 2430 2124 2514
rect 1816 2406 2124 2430
rect 1475 2368 2124 2406
rect 1475 2334 1782 2368
rect 1816 2334 2124 2368
rect 1475 2296 2124 2334
rect 1475 2262 1782 2296
rect 1816 2262 2124 2296
rect 2302 3570 2610 3592
rect 2302 3558 2321 3570
tri 2321 3558 2333 3570 nw
tri 2579 3558 2591 3570 ne
rect 2591 3558 2610 3570
rect 2644 3570 2952 3592
rect 2644 3558 2650 3570
rect 2302 3486 2308 3558
tri 2308 3545 2321 3558 nw
tri 2591 3545 2604 3558 ne
rect 2604 3520 2650 3558
tri 2650 3545 2675 3570 nw
tri 2921 3545 2946 3570 ne
tri 2308 3486 2333 3511 sw
tri 2579 3486 2604 3511 se
rect 2604 3486 2610 3520
rect 2644 3486 2650 3520
tri 2650 3486 2675 3511 sw
tri 2921 3486 2946 3511 se
rect 2946 3486 2952 3570
rect 2302 3448 2952 3486
rect 2302 3414 2610 3448
rect 2644 3414 2952 3448
rect 2302 3376 2952 3414
rect 2302 3342 2610 3376
rect 2644 3342 2952 3376
rect 2302 3306 2952 3342
rect 2302 3304 2331 3306
tri 2331 3304 2333 3306 nw
tri 2579 3304 2581 3306 ne
rect 2581 3304 2650 3306
rect 2302 3232 2308 3304
tri 2308 3281 2331 3304 nw
tri 2581 3281 2604 3304 ne
rect 2604 3270 2610 3304
rect 2644 3270 2650 3304
tri 2650 3281 2675 3306 nw
tri 2921 3281 2946 3306 ne
tri 2308 3232 2323 3247 sw
tri 2589 3232 2604 3247 se
rect 2604 3232 2650 3270
rect 2302 3222 2323 3232
tri 2323 3222 2333 3232 sw
tri 2579 3222 2589 3232 se
rect 2589 3222 2610 3232
rect 2302 3198 2610 3222
rect 2644 3222 2650 3232
tri 2650 3222 2675 3247 sw
tri 2921 3222 2946 3247 se
rect 2946 3222 2952 3306
rect 2644 3198 2952 3222
rect 2302 3160 2952 3198
rect 2302 3126 2610 3160
rect 2644 3126 2952 3160
rect 2302 3088 2952 3126
rect 2302 3054 2610 3088
rect 2644 3054 2952 3088
rect 2302 3042 2952 3054
rect 2302 2982 2308 3042
tri 2308 3017 2333 3042 nw
tri 2579 3017 2604 3042 ne
rect 2604 3016 2650 3042
tri 2650 3017 2675 3042 nw
tri 2921 3017 2946 3042 ne
tri 2308 2982 2309 2983 sw
tri 2603 2982 2604 2983 se
rect 2604 2982 2610 3016
rect 2644 2982 2650 3016
rect 2302 2958 2309 2982
tri 2309 2958 2333 2982 sw
tri 2579 2958 2603 2982 se
rect 2603 2958 2650 2982
tri 2650 2958 2675 2983 sw
tri 2921 2958 2946 2983 se
rect 2946 2958 2952 3042
rect 2302 2944 2952 2958
rect 2302 2910 2610 2944
rect 2644 2910 2952 2944
rect 2302 2872 2952 2910
rect 2302 2838 2610 2872
rect 2644 2838 2952 2872
rect 2302 2800 2952 2838
rect 2302 2778 2610 2800
rect 2302 2766 2321 2778
tri 2321 2766 2333 2778 nw
tri 2579 2766 2591 2778 ne
rect 2591 2766 2610 2778
rect 2644 2778 2952 2800
rect 2644 2766 2650 2778
rect 2302 2694 2308 2766
tri 2308 2753 2321 2766 nw
tri 2591 2753 2604 2766 ne
rect 2604 2728 2650 2766
tri 2650 2753 2675 2778 nw
tri 2921 2753 2946 2778 ne
tri 2308 2694 2333 2719 sw
tri 2579 2694 2604 2719 se
rect 2604 2694 2610 2728
rect 2644 2694 2650 2728
tri 2650 2694 2675 2719 sw
tri 2921 2694 2946 2719 se
rect 2946 2694 2952 2778
rect 2302 2656 2952 2694
rect 2302 2622 2610 2656
rect 2644 2622 2952 2656
rect 2302 2584 2952 2622
rect 2302 2550 2610 2584
rect 2644 2550 2952 2584
rect 2302 2514 2952 2550
rect 2302 2512 2331 2514
tri 2331 2512 2333 2514 nw
tri 2579 2512 2581 2514 ne
rect 2581 2512 2650 2514
rect 2302 2440 2308 2512
tri 2308 2489 2331 2512 nw
tri 2581 2489 2604 2512 ne
rect 2604 2478 2610 2512
rect 2644 2478 2650 2512
tri 2650 2489 2675 2514 nw
tri 2921 2489 2946 2514 ne
tri 2308 2440 2323 2455 sw
tri 2589 2440 2604 2455 se
rect 2604 2440 2650 2478
rect 2302 2430 2323 2440
tri 2323 2430 2333 2440 sw
tri 2579 2430 2589 2440 se
rect 2589 2430 2610 2440
rect 2302 2406 2610 2430
rect 2644 2430 2650 2440
tri 2650 2430 2675 2455 sw
tri 2921 2430 2946 2455 se
rect 2946 2430 2952 2514
rect 2644 2406 2952 2430
rect 2302 2368 2952 2406
rect 2302 2334 2610 2368
rect 2644 2334 2952 2368
rect 2302 2296 2952 2334
rect 2302 2262 2610 2296
rect 2644 2262 2952 2296
rect 3130 3570 3438 3592
rect 3130 3558 3149 3570
tri 3149 3558 3161 3570 nw
tri 3407 3558 3419 3570 ne
rect 3419 3558 3438 3570
rect 3472 3570 3781 3592
rect 3472 3558 3478 3570
rect 3130 3486 3136 3558
tri 3136 3545 3149 3558 nw
tri 3419 3545 3432 3558 ne
rect 3432 3520 3478 3558
tri 3478 3545 3503 3570 nw
tri 3750 3545 3775 3570 ne
tri 3136 3486 3161 3511 sw
tri 3407 3486 3432 3511 se
rect 3432 3486 3438 3520
rect 3472 3486 3478 3520
tri 3478 3486 3503 3511 sw
tri 3750 3486 3775 3511 se
rect 3775 3486 3781 3570
rect 3130 3448 3781 3486
rect 3130 3414 3438 3448
rect 3472 3414 3781 3448
rect 3130 3376 3781 3414
rect 3130 3342 3438 3376
rect 3472 3342 3781 3376
rect 3130 3306 3781 3342
rect 3130 3304 3159 3306
tri 3159 3304 3161 3306 nw
tri 3407 3304 3409 3306 ne
rect 3409 3304 3478 3306
rect 3130 3232 3136 3304
tri 3136 3281 3159 3304 nw
tri 3409 3281 3432 3304 ne
rect 3432 3270 3438 3304
rect 3472 3270 3478 3304
tri 3478 3281 3503 3306 nw
tri 3750 3281 3775 3306 ne
tri 3136 3232 3151 3247 sw
tri 3417 3232 3432 3247 se
rect 3432 3232 3478 3270
rect 3130 3222 3151 3232
tri 3151 3222 3161 3232 sw
tri 3407 3222 3417 3232 se
rect 3417 3222 3438 3232
rect 3130 3198 3438 3222
rect 3472 3222 3478 3232
tri 3478 3222 3503 3247 sw
tri 3750 3222 3775 3247 se
rect 3775 3222 3781 3306
rect 3472 3198 3781 3222
rect 3130 3160 3781 3198
rect 3130 3126 3438 3160
rect 3472 3126 3781 3160
rect 3130 3088 3781 3126
rect 3130 3054 3438 3088
rect 3472 3054 3781 3088
rect 3130 3042 3781 3054
rect 3130 2982 3136 3042
tri 3136 3017 3161 3042 nw
tri 3407 3017 3432 3042 ne
rect 3432 3016 3478 3042
tri 3478 3017 3503 3042 nw
tri 3750 3017 3775 3042 ne
tri 3136 2982 3137 2983 sw
tri 3431 2982 3432 2983 se
rect 3432 2982 3438 3016
rect 3472 2982 3478 3016
rect 3130 2958 3137 2982
tri 3137 2958 3161 2982 sw
tri 3407 2958 3431 2982 se
rect 3431 2958 3478 2982
tri 3478 2958 3503 2983 sw
tri 3750 2958 3775 2983 se
rect 3775 2958 3781 3042
rect 3130 2944 3781 2958
rect 3130 2910 3438 2944
rect 3472 2910 3781 2944
rect 3130 2872 3781 2910
rect 3130 2838 3438 2872
rect 3472 2838 3781 2872
rect 3130 2800 3781 2838
rect 3130 2778 3438 2800
rect 3130 2766 3149 2778
tri 3149 2766 3161 2778 nw
tri 3407 2766 3419 2778 ne
rect 3419 2766 3438 2778
rect 3472 2778 3781 2800
rect 3472 2766 3478 2778
rect 3130 2694 3136 2766
tri 3136 2753 3149 2766 nw
tri 3419 2753 3432 2766 ne
rect 3432 2728 3478 2766
tri 3478 2753 3503 2778 nw
tri 3750 2753 3775 2778 ne
tri 3136 2694 3161 2719 sw
tri 3407 2694 3432 2719 se
rect 3432 2694 3438 2728
rect 3472 2694 3478 2728
tri 3478 2694 3503 2719 sw
tri 3750 2694 3775 2719 se
rect 3775 2694 3781 2778
rect 3130 2656 3781 2694
rect 3130 2622 3438 2656
rect 3472 2622 3781 2656
rect 3130 2584 3781 2622
rect 3130 2550 3438 2584
rect 3472 2550 3781 2584
rect 3130 2514 3781 2550
rect 3130 2512 3159 2514
tri 3159 2512 3161 2514 nw
tri 3407 2512 3409 2514 ne
rect 3409 2512 3478 2514
rect 3130 2440 3136 2512
tri 3136 2489 3159 2512 nw
tri 3409 2489 3432 2512 ne
rect 3432 2478 3438 2512
rect 3472 2478 3478 2512
tri 3478 2489 3503 2514 nw
tri 3750 2489 3775 2514 ne
tri 3136 2440 3151 2455 sw
tri 3417 2440 3432 2455 se
rect 3432 2440 3478 2478
rect 3130 2430 3151 2440
tri 3151 2430 3161 2440 sw
tri 3407 2430 3417 2440 se
rect 3417 2430 3438 2440
rect 3130 2406 3438 2430
rect 3472 2430 3478 2440
tri 3478 2430 3503 2455 sw
tri 3750 2430 3775 2455 se
rect 3775 2430 3781 2514
rect 3472 2406 3781 2430
rect 3130 2368 3781 2406
rect 3130 2334 3438 2368
rect 3472 2334 3781 2368
rect 3130 2296 3781 2334
rect 3130 2262 3438 2296
rect 3472 2262 3781 2296
rect 3959 3570 4266 3592
rect 3959 3558 3978 3570
tri 3978 3558 3990 3570 nw
tri 4235 3558 4247 3570 ne
rect 4247 3558 4266 3570
rect 4300 3570 4608 3592
rect 4300 3558 4306 3570
rect 3959 3486 3965 3558
tri 3965 3545 3978 3558 nw
tri 4247 3545 4260 3558 ne
rect 4260 3520 4306 3558
tri 4306 3545 4331 3570 nw
tri 4577 3545 4602 3570 ne
tri 3965 3486 3990 3511 sw
tri 4235 3486 4260 3511 se
rect 4260 3486 4266 3520
rect 4300 3486 4306 3520
tri 4306 3486 4331 3511 sw
tri 4577 3486 4602 3511 se
rect 4602 3486 4608 3570
rect 3959 3448 4608 3486
rect 3959 3414 4266 3448
rect 4300 3414 4608 3448
rect 3959 3376 4608 3414
rect 3959 3342 4266 3376
rect 4300 3342 4608 3376
rect 3959 3306 4608 3342
rect 3959 3304 3988 3306
tri 3988 3304 3990 3306 nw
tri 4235 3304 4237 3306 ne
rect 4237 3304 4306 3306
rect 3959 3232 3965 3304
tri 3965 3281 3988 3304 nw
tri 4237 3281 4260 3304 ne
rect 4260 3270 4266 3304
rect 4300 3270 4306 3304
tri 4306 3281 4331 3306 nw
tri 4577 3281 4602 3306 ne
tri 3965 3232 3980 3247 sw
tri 4245 3232 4260 3247 se
rect 4260 3232 4306 3270
rect 3959 3222 3980 3232
tri 3980 3222 3990 3232 sw
tri 4235 3222 4245 3232 se
rect 4245 3222 4266 3232
rect 3959 3198 4266 3222
rect 4300 3222 4306 3232
tri 4306 3222 4331 3247 sw
tri 4577 3222 4602 3247 se
rect 4602 3222 4608 3306
rect 4300 3198 4608 3222
rect 3959 3160 4608 3198
rect 3959 3126 4266 3160
rect 4300 3126 4608 3160
rect 3959 3088 4608 3126
rect 3959 3054 4266 3088
rect 4300 3054 4608 3088
rect 3959 3042 4608 3054
rect 3959 2982 3965 3042
tri 3965 3017 3990 3042 nw
tri 4235 3017 4260 3042 ne
rect 4260 3016 4306 3042
tri 4306 3017 4331 3042 nw
tri 4577 3017 4602 3042 ne
tri 3965 2982 3966 2983 sw
tri 4259 2982 4260 2983 se
rect 4260 2982 4266 3016
rect 4300 2982 4306 3016
rect 3959 2958 3966 2982
tri 3966 2958 3990 2982 sw
tri 4235 2958 4259 2982 se
rect 4259 2958 4306 2982
tri 4306 2958 4331 2983 sw
tri 4577 2958 4602 2983 se
rect 4602 2958 4608 3042
rect 3959 2944 4608 2958
rect 3959 2910 4266 2944
rect 4300 2910 4608 2944
rect 3959 2872 4608 2910
rect 3959 2838 4266 2872
rect 4300 2838 4608 2872
rect 3959 2800 4608 2838
rect 3959 2778 4266 2800
rect 3959 2766 3978 2778
tri 3978 2766 3990 2778 nw
tri 4235 2766 4247 2778 ne
rect 4247 2766 4266 2778
rect 4300 2778 4608 2800
rect 4300 2766 4306 2778
rect 3959 2694 3965 2766
tri 3965 2753 3978 2766 nw
tri 4247 2753 4260 2766 ne
rect 4260 2728 4306 2766
tri 4306 2753 4331 2778 nw
tri 4577 2753 4602 2778 ne
tri 3965 2694 3990 2719 sw
tri 4235 2694 4260 2719 se
rect 4260 2694 4266 2728
rect 4300 2694 4306 2728
tri 4306 2694 4331 2719 sw
tri 4577 2694 4602 2719 se
rect 4602 2694 4608 2778
rect 3959 2656 4608 2694
rect 3959 2622 4266 2656
rect 4300 2622 4608 2656
rect 3959 2584 4608 2622
rect 3959 2550 4266 2584
rect 4300 2550 4608 2584
rect 3959 2514 4608 2550
rect 3959 2512 3988 2514
tri 3988 2512 3990 2514 nw
tri 4235 2512 4237 2514 ne
rect 4237 2512 4306 2514
rect 3959 2440 3965 2512
tri 3965 2489 3988 2512 nw
tri 4237 2489 4260 2512 ne
rect 4260 2478 4266 2512
rect 4300 2478 4306 2512
tri 4306 2489 4331 2514 nw
tri 4577 2489 4602 2514 ne
tri 3965 2440 3980 2455 sw
tri 4245 2440 4260 2455 se
rect 4260 2440 4306 2478
rect 3959 2430 3980 2440
tri 3980 2430 3990 2440 sw
tri 4235 2430 4245 2440 se
rect 4245 2430 4266 2440
rect 3959 2406 4266 2430
rect 4300 2430 4306 2440
tri 4306 2430 4331 2455 sw
tri 4577 2430 4602 2455 se
rect 4602 2430 4608 2514
rect 4300 2406 4608 2430
rect 3959 2368 4608 2406
rect 3959 2334 4266 2368
rect 4300 2334 4608 2368
rect 3959 2296 4608 2334
rect 3959 2262 4266 2296
rect 4300 2262 4608 2296
rect 4786 3570 5094 3592
rect 4786 3558 4805 3570
tri 4805 3558 4817 3570 nw
tri 5063 3558 5075 3570 ne
rect 5075 3558 5094 3570
rect 5128 3570 5522 3592
rect 5128 3568 5157 3570
tri 5157 3568 5159 3570 nw
tri 5419 3568 5421 3570 ne
rect 5421 3568 5522 3570
rect 5128 3563 5152 3568
tri 5152 3563 5157 3568 nw
tri 5421 3563 5426 3568 ne
rect 5426 3563 5594 3568
rect 5128 3558 5134 3563
rect 4786 3486 4792 3558
tri 4792 3545 4805 3558 nw
tri 5075 3545 5088 3558 ne
rect 5088 3520 5134 3558
tri 5134 3545 5152 3563 nw
tri 5426 3545 5444 3563 ne
tri 4792 3486 4817 3511 sw
tri 5063 3486 5088 3511 se
rect 5088 3486 5094 3520
rect 5128 3495 5134 3520
rect 5444 3529 5450 3563
rect 5484 3529 5594 3563
tri 5134 3495 5150 3511 sw
tri 5428 3495 5444 3511 se
rect 5444 3495 5522 3529
rect 5556 3495 5594 3529
rect 5128 3490 5150 3495
tri 5150 3490 5155 3495 sw
tri 5423 3490 5428 3495 se
rect 5428 3490 5594 3495
rect 5128 3486 5155 3490
tri 5155 3486 5159 3490 sw
tri 5419 3486 5423 3490 se
rect 5423 3486 5450 3490
rect 4786 3456 5450 3486
rect 5484 3456 5594 3490
rect 4786 3448 5522 3456
rect 4786 3414 5094 3448
rect 5128 3422 5522 3448
rect 5556 3422 5594 3456
rect 5128 3417 5594 3422
rect 5128 3414 5450 3417
rect 4786 3383 5450 3414
rect 5484 3383 5594 3417
rect 4786 3376 5522 3383
rect 4786 3342 5094 3376
rect 5128 3349 5522 3376
rect 5556 3349 5594 3383
rect 5128 3344 5594 3349
rect 5128 3342 5450 3344
rect 4786 3310 5450 3342
rect 5484 3310 5594 3344
rect 4786 3306 5522 3310
rect 4786 3304 4815 3306
tri 4815 3304 4817 3306 nw
tri 5063 3304 5065 3306 ne
rect 5065 3304 5134 3306
rect 4786 3237 4792 3304
tri 4792 3281 4815 3304 nw
tri 5065 3281 5088 3304 ne
rect 5088 3270 5094 3304
rect 5128 3270 5134 3304
tri 5134 3281 5159 3306 nw
tri 5419 3281 5444 3306 ne
tri 4792 3237 4802 3247 sw
tri 5078 3237 5088 3247 se
rect 5088 3237 5134 3270
rect 5444 3276 5522 3306
rect 5556 3276 5594 3310
rect 5444 3271 5594 3276
tri 5134 3237 5144 3247 sw
tri 5434 3237 5444 3247 se
rect 5444 3237 5450 3271
rect 5484 3237 5594 3271
rect 4786 3232 4802 3237
tri 4802 3232 4807 3237 sw
tri 5073 3232 5078 3237 se
rect 5078 3232 5144 3237
rect 4786 3222 4807 3232
tri 4807 3222 4817 3232 sw
tri 5063 3222 5073 3232 se
rect 5073 3222 5094 3232
rect 4786 3198 5094 3222
rect 5128 3222 5144 3232
tri 5144 3222 5159 3237 sw
tri 5419 3222 5434 3237 se
rect 5434 3222 5522 3237
rect 5128 3203 5522 3222
rect 5556 3203 5594 3237
rect 5128 3198 5594 3203
rect 4786 3164 5450 3198
rect 5484 3164 5594 3198
rect 4786 3160 5522 3164
rect 4786 3126 5094 3160
rect 5128 3130 5522 3160
rect 5556 3130 5594 3164
rect 5128 3126 5594 3130
rect 4786 3125 5594 3126
rect 4786 3091 5450 3125
rect 5484 3091 5594 3125
rect 4786 3088 5522 3091
rect 4786 3054 5094 3088
rect 5128 3057 5522 3088
rect 5556 3057 5594 3091
rect 5128 3054 5594 3057
rect 4786 3052 5594 3054
rect 4786 3042 5450 3052
rect 4786 3018 4793 3042
tri 4793 3018 4817 3042 nw
tri 5063 3018 5087 3042 ne
rect 5087 3018 5135 3042
tri 5135 3018 5159 3042 nw
tri 5419 3018 5443 3042 ne
rect 5443 3018 5450 3042
rect 5484 3018 5594 3052
rect 4786 2982 4792 3018
tri 4792 3017 4793 3018 nw
tri 5087 3017 5088 3018 ne
rect 5088 3016 5134 3018
tri 5134 3017 5135 3018 nw
tri 5443 3017 5444 3018 ne
tri 4792 2982 4793 2983 sw
tri 5087 2982 5088 2983 se
rect 5088 2982 5094 3016
rect 5128 2982 5134 3016
rect 5444 2984 5522 3018
rect 5556 2984 5594 3018
rect 4786 2979 4793 2982
tri 4793 2979 4796 2982 sw
tri 5084 2979 5087 2982 se
rect 5087 2979 5134 2982
tri 5134 2979 5138 2983 sw
tri 5440 2979 5444 2983 se
rect 5444 2979 5594 2984
rect 4786 2958 4796 2979
tri 4796 2958 4817 2979 sw
tri 5063 2958 5084 2979 se
rect 5084 2958 5138 2979
tri 5138 2958 5159 2979 sw
tri 5419 2958 5440 2979 se
rect 5440 2958 5450 2979
rect 4786 2945 5450 2958
rect 5484 2952 5594 2979
rect 5700 2952 5712 3850
rect 5484 2945 5712 2952
rect 4786 2944 5522 2945
rect 4786 2910 5094 2944
rect 5128 2911 5522 2944
rect 5556 2913 5712 2945
rect 5556 2911 5594 2913
rect 5128 2910 5594 2911
rect 4786 2906 5594 2910
rect 4786 2872 5450 2906
rect 5484 2879 5594 2906
rect 5628 2879 5666 2913
rect 5700 2879 5712 2913
rect 5484 2872 5712 2879
rect 4786 2838 5094 2872
rect 5128 2838 5522 2872
rect 5556 2840 5712 2872
rect 5556 2838 5594 2840
rect 4786 2833 5594 2838
rect 4786 2800 5450 2833
rect 4786 2778 5094 2800
rect 4786 2766 4805 2778
tri 4805 2766 4817 2778 nw
tri 5063 2766 5075 2778 ne
rect 5075 2766 5094 2778
rect 5128 2799 5450 2800
rect 5484 2806 5594 2833
rect 5628 2806 5666 2840
rect 5700 2806 5712 2840
rect 5484 2799 5712 2806
rect 5128 2778 5522 2799
rect 5128 2766 5146 2778
rect 4786 2765 4804 2766
tri 4804 2765 4805 2766 nw
tri 5075 2765 5076 2766 ne
rect 5076 2765 5146 2766
tri 5146 2765 5159 2778 nw
tri 5419 2765 5432 2778 ne
rect 5432 2765 5522 2778
rect 5556 2767 5712 2799
rect 5556 2765 5594 2767
rect 4786 2760 4799 2765
tri 4799 2760 4804 2765 nw
tri 5076 2760 5081 2765 ne
rect 5081 2760 5141 2765
tri 5141 2760 5146 2765 nw
tri 5432 2760 5437 2765 ne
rect 5437 2760 5594 2765
rect 4786 2694 4792 2760
tri 4792 2753 4799 2760 nw
tri 5081 2753 5088 2760 ne
rect 5088 2728 5134 2760
tri 5134 2753 5141 2760 nw
tri 5437 2753 5444 2760 ne
tri 4792 2694 4817 2719 sw
tri 5063 2694 5088 2719 se
rect 5088 2694 5094 2728
rect 5128 2694 5134 2728
rect 5444 2726 5450 2760
rect 5484 2733 5594 2760
rect 5628 2733 5666 2767
rect 5700 2733 5712 2767
rect 5484 2726 5712 2733
tri 5134 2694 5159 2719 sw
tri 5419 2694 5444 2719 se
rect 5444 2694 5522 2726
rect 4786 2692 5522 2694
rect 5556 2694 5712 2726
rect 5556 2692 5594 2694
rect 4786 2687 5594 2692
rect 4786 2656 5450 2687
rect 4786 2622 5094 2656
rect 5128 2653 5450 2656
rect 5484 2660 5594 2687
rect 5628 2660 5666 2694
rect 5700 2660 5712 2694
rect 5484 2653 5712 2660
rect 5128 2622 5522 2653
rect 4786 2619 5522 2622
rect 5556 2621 5712 2653
rect 5556 2619 5594 2621
rect 4786 2614 5594 2619
rect 4786 2584 5450 2614
rect 4786 2550 5094 2584
rect 5128 2580 5450 2584
rect 5484 2587 5594 2614
rect 5628 2587 5666 2621
rect 5700 2587 5712 2621
rect 5484 2580 5712 2587
rect 5128 2550 5522 2580
rect 4786 2546 5522 2550
rect 5556 2548 5712 2580
rect 5556 2546 5594 2548
rect 4786 2541 5594 2546
rect 4786 2514 5450 2541
rect 4786 2512 4815 2514
tri 4815 2512 4817 2514 nw
tri 5063 2512 5065 2514 ne
rect 5065 2512 5152 2514
rect 4786 2440 4792 2512
tri 4792 2489 4815 2512 nw
tri 5065 2489 5088 2512 ne
rect 5088 2478 5094 2512
rect 5128 2507 5152 2512
tri 5152 2507 5159 2514 nw
tri 5419 2507 5426 2514 ne
rect 5426 2507 5450 2514
rect 5484 2514 5594 2541
rect 5628 2514 5666 2548
rect 5700 2514 5712 2548
rect 5484 2507 5712 2514
rect 5128 2478 5134 2507
tri 5134 2489 5152 2507 nw
tri 5426 2489 5444 2507 ne
tri 4792 2440 4807 2455 sw
tri 5073 2440 5088 2455 se
rect 5088 2440 5134 2478
rect 5444 2473 5522 2507
rect 5556 2475 5712 2507
rect 5556 2473 5594 2475
rect 5444 2468 5594 2473
rect 4786 2430 4807 2440
tri 4807 2430 4817 2440 sw
tri 5063 2430 5073 2440 se
rect 5073 2430 5094 2440
rect 4786 2406 5094 2430
rect 5128 2434 5134 2440
tri 5134 2434 5155 2455 sw
tri 5423 2434 5444 2455 se
rect 5444 2434 5450 2468
rect 5484 2441 5594 2468
rect 5628 2441 5666 2475
rect 5700 2441 5712 2475
rect 5484 2434 5712 2441
rect 5128 2430 5155 2434
tri 5155 2430 5159 2434 sw
tri 5419 2430 5423 2434 se
rect 5423 2430 5522 2434
rect 5128 2406 5522 2430
rect 4786 2400 5522 2406
rect 5556 2402 5712 2434
rect 5556 2400 5594 2402
rect 4786 2395 5594 2400
rect 4786 2368 5450 2395
rect 4786 2334 5094 2368
rect 5128 2361 5450 2368
rect 5484 2368 5594 2395
rect 5628 2368 5666 2402
rect 5700 2368 5712 2402
rect 5484 2361 5712 2368
rect 5128 2334 5522 2361
rect 4786 2327 5522 2334
rect 5556 2329 5712 2361
rect 5556 2327 5594 2329
rect 4786 2322 5594 2327
rect 4786 2296 5450 2322
rect 4786 2262 5094 2296
rect 5128 2288 5450 2296
rect 5484 2295 5594 2322
rect 5628 2295 5666 2329
rect 5700 2295 5712 2329
rect 5484 2288 5712 2295
rect 5128 2262 5522 2288
rect 560 2254 5522 2262
rect 5556 2256 5712 2288
rect 5556 2254 5594 2256
rect 560 2250 5594 2254
rect 560 2249 662 2250
tri 662 2249 663 2250 nw
tri 5419 2249 5420 2250 ne
rect 5420 2249 5594 2250
rect 488 2222 598 2249
rect 370 2215 598 2222
rect 632 2215 638 2249
tri 638 2225 662 2249 nw
tri 5420 2225 5444 2249 ne
rect 370 2210 638 2215
rect 370 2183 526 2210
rect 370 2149 382 2183
rect 416 2149 454 2183
rect 488 2176 526 2183
rect 560 2176 638 2210
rect 488 2149 598 2176
rect 370 2142 598 2149
rect 632 2142 638 2176
rect 370 2137 638 2142
rect 370 2110 526 2137
rect 370 2076 382 2110
rect 416 2076 454 2110
rect 488 2103 526 2110
rect 560 2103 638 2137
rect 488 2076 598 2103
rect 370 2069 598 2076
rect 632 2069 638 2103
rect 370 2064 638 2069
rect 370 2037 526 2064
rect 370 2003 382 2037
rect 416 2003 454 2037
rect 488 2030 526 2037
rect 560 2030 638 2064
rect 488 2003 598 2030
rect 370 1996 598 2003
rect 632 1996 638 2030
rect 370 1991 638 1996
rect 370 1964 526 1991
rect 370 1930 382 1964
rect 416 1930 454 1964
rect 488 1957 526 1964
rect 560 1957 638 1991
rect 488 1930 598 1957
rect 370 1923 598 1930
rect 632 1923 638 1957
rect 370 1918 638 1923
rect 370 1891 526 1918
rect 370 1857 382 1891
rect 416 1857 454 1891
rect 488 1884 526 1891
rect 560 1884 638 1918
rect 488 1857 598 1884
rect 370 1850 598 1857
rect 632 1850 638 1884
rect 370 1845 638 1850
rect 370 1818 526 1845
rect 370 1784 382 1818
rect 416 1784 454 1818
rect 488 1811 526 1818
rect 560 1811 638 1845
rect 488 1784 598 1811
rect 370 1777 598 1784
rect 632 1777 638 1811
rect 370 1772 638 1777
rect 370 1745 526 1772
rect 370 1711 382 1745
rect 416 1711 454 1745
rect 488 1738 526 1745
rect 560 1738 638 1772
rect 488 1711 598 1738
rect 370 1704 598 1711
rect 632 1704 638 1738
rect 370 1699 638 1704
rect 370 1672 526 1699
rect 370 1638 382 1672
rect 416 1638 454 1672
rect 488 1665 526 1672
rect 560 1665 638 1699
rect 488 1638 598 1665
rect 370 1631 598 1638
rect 632 1631 638 1665
rect 370 1626 638 1631
rect 370 1599 526 1626
rect 370 1565 382 1599
rect 416 1565 454 1599
rect 488 1592 526 1599
rect 560 1592 638 1626
rect 488 1565 598 1592
rect 370 1558 598 1565
rect 632 1558 638 1592
rect 370 1553 638 1558
rect 370 1526 526 1553
rect 370 1492 382 1526
rect 416 1492 454 1526
rect 488 1519 526 1526
rect 560 1519 638 1553
rect 488 1492 598 1519
rect 370 1485 598 1492
rect 632 1485 638 1519
rect 370 1480 638 1485
rect 370 1453 526 1480
rect 370 1419 382 1453
rect 416 1419 454 1453
rect 488 1446 526 1453
rect 560 1446 638 1480
rect 488 1419 598 1446
rect 370 1412 598 1419
rect 632 1412 638 1446
rect 370 1407 638 1412
rect 370 1380 526 1407
rect 370 1346 382 1380
rect 416 1346 454 1380
rect 488 1373 526 1380
rect 560 1373 638 1407
rect 488 1346 598 1373
rect 370 1339 598 1346
rect 632 1339 638 1373
rect 370 1334 638 1339
rect 370 1307 526 1334
rect 370 1273 382 1307
rect 416 1273 454 1307
rect 488 1300 526 1307
rect 560 1300 638 1334
rect 488 1273 598 1300
rect 370 1266 598 1273
rect 632 1266 638 1300
rect 370 1261 638 1266
rect 370 1234 526 1261
rect 370 1200 382 1234
rect 416 1200 454 1234
rect 488 1227 526 1234
rect 560 1227 638 1261
rect 488 1200 598 1227
rect 370 1193 598 1200
rect 632 1193 638 1227
rect 370 1188 638 1193
rect 370 1161 526 1188
rect 370 1127 382 1161
rect 416 1127 454 1161
rect 488 1154 526 1161
rect 560 1154 638 1188
rect 488 1127 598 1154
rect 370 1120 598 1127
rect 632 1120 638 1154
rect 370 1115 638 1120
rect 370 1088 526 1115
rect 370 1054 382 1088
rect 416 1054 454 1088
rect 488 1081 526 1088
rect 560 1081 638 1115
rect 488 1054 598 1081
rect 370 1047 598 1054
rect 632 1047 638 1081
rect 370 1042 638 1047
rect 370 1015 526 1042
rect 370 981 382 1015
rect 416 981 454 1015
rect 488 1008 526 1015
rect 560 1008 638 1042
rect 488 981 598 1008
rect 370 974 598 981
rect 632 974 638 1008
rect 370 969 638 974
rect 370 942 526 969
rect 370 908 382 942
rect 416 908 454 942
rect 488 935 526 942
rect 560 935 638 969
rect 488 908 598 935
rect 370 901 598 908
rect 632 901 638 935
rect 370 896 638 901
rect 370 869 526 896
rect 370 835 382 869
rect 416 835 454 869
rect 488 862 526 869
rect 560 862 638 896
rect 488 835 598 862
rect 370 828 598 835
rect 632 828 638 862
rect 370 824 638 828
rect 370 796 526 824
rect 370 762 382 796
rect 416 762 454 796
rect 488 790 526 796
rect 560 790 638 824
rect 488 789 638 790
rect 488 762 598 789
rect 370 755 598 762
rect 632 755 638 789
rect 370 752 638 755
rect 370 723 526 752
rect 370 689 382 723
rect 416 689 454 723
rect 488 718 526 723
rect 560 718 638 752
rect 792 2210 5290 2222
rect 792 2176 798 2210
rect 832 2176 1110 2210
rect 1144 2176 1626 2210
rect 1660 2176 1938 2210
rect 1972 2176 2454 2210
rect 2488 2176 2766 2210
rect 2800 2176 3282 2210
rect 3316 2176 3594 2210
rect 3628 2176 4110 2210
rect 4144 2176 4422 2210
rect 4456 2176 4938 2210
rect 4972 2176 5250 2210
rect 5284 2176 5290 2210
rect 792 2137 5290 2176
rect 792 2103 798 2137
rect 832 2103 1110 2137
rect 1144 2103 1626 2137
rect 1660 2103 1938 2137
rect 1972 2103 2454 2137
rect 2488 2103 2766 2137
rect 2800 2103 3282 2137
rect 3316 2103 3594 2137
rect 3628 2103 4110 2137
rect 4144 2103 4422 2137
rect 4456 2103 4938 2137
rect 4972 2103 5250 2137
rect 5284 2103 5290 2137
rect 792 2064 5290 2103
rect 792 2030 798 2064
rect 832 2042 1110 2064
rect 832 2030 851 2042
tri 851 2030 863 2042 nw
tri 1079 2030 1091 2042 ne
rect 1091 2030 1110 2042
rect 1144 2042 1626 2064
rect 1144 2030 1163 2042
tri 1163 2030 1175 2042 nw
tri 1595 2030 1607 2042 ne
rect 1607 2030 1626 2042
rect 1660 2042 1938 2064
rect 1660 2030 1679 2042
tri 1679 2030 1691 2042 nw
tri 1907 2030 1919 2042 ne
rect 1919 2030 1938 2042
rect 1972 2042 2454 2064
rect 1972 2030 1991 2042
tri 1991 2030 2003 2042 nw
tri 2423 2030 2435 2042 ne
rect 2435 2030 2454 2042
rect 2488 2042 2766 2064
rect 2488 2030 2507 2042
tri 2507 2030 2519 2042 nw
tri 2735 2030 2747 2042 ne
rect 2747 2030 2766 2042
rect 2800 2042 3282 2064
rect 2800 2030 2819 2042
tri 2819 2030 2831 2042 nw
tri 3251 2030 3263 2042 ne
rect 3263 2030 3282 2042
rect 3316 2042 3594 2064
rect 3316 2030 3335 2042
tri 3335 2030 3347 2042 nw
tri 3563 2030 3575 2042 ne
rect 3575 2030 3594 2042
rect 3628 2042 4110 2064
rect 3628 2030 3647 2042
tri 3647 2030 3659 2042 nw
tri 4079 2030 4091 2042 ne
rect 4091 2030 4110 2042
rect 4144 2042 4422 2064
rect 4144 2030 4163 2042
tri 4163 2030 4175 2042 nw
tri 4391 2030 4403 2042 ne
rect 4403 2030 4422 2042
rect 4456 2042 4938 2064
rect 4456 2030 4475 2042
tri 4475 2030 4487 2042 nw
tri 4907 2030 4919 2042 ne
rect 4919 2030 4938 2042
rect 4972 2042 5250 2064
rect 4972 2030 4991 2042
tri 4991 2030 5003 2042 nw
tri 5219 2030 5231 2042 ne
rect 5231 2030 5250 2042
rect 5284 2030 5290 2064
rect 792 1992 838 2030
tri 838 2017 851 2030 nw
tri 1091 2017 1104 2030 ne
rect 792 1958 798 1992
rect 832 1958 838 1992
rect 1104 1992 1150 2030
tri 1150 2017 1163 2030 nw
tri 1607 2017 1620 2030 ne
tri 838 1958 863 1983 sw
tri 1079 1958 1104 1983 se
rect 1104 1958 1110 1992
rect 1144 1958 1150 1992
rect 1620 1992 1666 2030
tri 1666 2017 1679 2030 nw
tri 1919 2017 1932 2030 ne
tri 1150 1958 1175 1983 sw
tri 1595 1958 1620 1983 se
rect 1620 1958 1626 1992
rect 1660 1958 1666 1992
rect 1932 1992 1978 2030
tri 1978 2017 1991 2030 nw
tri 2435 2017 2448 2030 ne
tri 1666 1958 1691 1983 sw
tri 1907 1958 1932 1983 se
rect 1932 1958 1938 1992
rect 1972 1958 1978 1992
rect 2448 1992 2494 2030
tri 2494 2017 2507 2030 nw
tri 2747 2017 2760 2030 ne
tri 1978 1958 2003 1983 sw
tri 2423 1958 2448 1983 se
rect 2448 1958 2454 1992
rect 2488 1958 2494 1992
rect 2760 1992 2806 2030
tri 2806 2017 2819 2030 nw
tri 3263 2017 3276 2030 ne
tri 2494 1958 2519 1983 sw
tri 2735 1958 2760 1983 se
rect 2760 1958 2766 1992
rect 2800 1958 2806 1992
rect 3276 1992 3322 2030
tri 3322 2017 3335 2030 nw
tri 3575 2017 3588 2030 ne
tri 2806 1958 2831 1983 sw
tri 3251 1958 3276 1983 se
rect 3276 1958 3282 1992
rect 3316 1958 3322 1992
rect 3588 1992 3634 2030
tri 3634 2017 3647 2030 nw
tri 4091 2017 4104 2030 ne
tri 3322 1958 3347 1983 sw
tri 3563 1958 3588 1983 se
rect 3588 1958 3594 1992
rect 3628 1958 3634 1992
rect 4104 1992 4150 2030
tri 4150 2017 4163 2030 nw
tri 4403 2017 4416 2030 ne
tri 3634 1958 3659 1983 sw
tri 4079 1958 4104 1983 se
rect 4104 1958 4110 1992
rect 4144 1958 4150 1992
rect 4416 1992 4462 2030
tri 4462 2017 4475 2030 nw
tri 4919 2017 4932 2030 ne
tri 4150 1958 4175 1983 sw
tri 4391 1958 4416 1983 se
rect 4416 1958 4422 1992
rect 4456 1958 4462 1992
rect 4932 1992 4978 2030
tri 4978 2017 4991 2030 nw
tri 5231 2017 5244 2030 ne
tri 4462 1958 4487 1983 sw
tri 4907 1958 4932 1983 se
rect 4932 1958 4938 1992
rect 4972 1958 4978 1992
rect 5244 1992 5290 2030
tri 4978 1958 5003 1983 sw
tri 5219 1958 5244 1983 se
rect 5244 1958 5250 1992
rect 5284 1958 5290 1992
rect 792 1920 5290 1958
rect 792 1886 798 1920
rect 832 1886 1110 1920
rect 1144 1886 1626 1920
rect 1660 1886 1938 1920
rect 1972 1886 2454 1920
rect 2488 1886 2766 1920
rect 2800 1886 3282 1920
rect 3316 1886 3594 1920
rect 3628 1886 4110 1920
rect 4144 1886 4422 1920
rect 4456 1886 4938 1920
rect 4972 1886 5250 1920
rect 5284 1886 5290 1920
rect 792 1848 5290 1886
rect 792 1814 798 1848
rect 832 1814 1110 1848
rect 1144 1814 1626 1848
rect 1660 1814 1938 1848
rect 1972 1814 2454 1848
rect 2488 1814 2766 1848
rect 2800 1814 3282 1848
rect 3316 1814 3594 1848
rect 3628 1814 4110 1848
rect 4144 1814 4422 1848
rect 4456 1814 4938 1848
rect 4972 1814 5250 1848
rect 5284 1814 5290 1848
rect 792 1778 5290 1814
rect 792 1777 862 1778
tri 862 1777 863 1778 nw
tri 1079 1777 1080 1778 ne
rect 1080 1777 1174 1778
tri 1174 1777 1175 1778 nw
tri 1595 1777 1596 1778 ne
rect 1596 1777 1690 1778
tri 1690 1777 1691 1778 nw
tri 1907 1777 1908 1778 ne
rect 1908 1777 2002 1778
tri 2002 1777 2003 1778 nw
tri 2423 1777 2424 1778 ne
rect 2424 1777 2518 1778
tri 2518 1777 2519 1778 nw
tri 2735 1777 2736 1778 ne
rect 2736 1777 2830 1778
tri 2830 1777 2831 1778 nw
tri 3251 1777 3252 1778 ne
rect 3252 1777 3346 1778
tri 3346 1777 3347 1778 nw
tri 3563 1777 3564 1778 ne
rect 3564 1777 3658 1778
tri 3658 1777 3659 1778 nw
tri 4079 1777 4080 1778 ne
rect 4080 1777 4174 1778
tri 4174 1777 4175 1778 nw
tri 4391 1777 4392 1778 ne
rect 4392 1777 4486 1778
tri 4486 1777 4487 1778 nw
tri 4907 1777 4908 1778 ne
rect 4908 1777 5002 1778
tri 5002 1777 5003 1778 nw
tri 5219 1777 5220 1778 ne
rect 5220 1777 5290 1778
rect 792 1776 861 1777
tri 861 1776 862 1777 nw
tri 1080 1776 1081 1777 ne
rect 1081 1776 1173 1777
tri 1173 1776 1174 1777 nw
tri 1596 1776 1597 1777 ne
rect 1597 1776 1689 1777
tri 1689 1776 1690 1777 nw
tri 1908 1776 1909 1777 ne
rect 1909 1776 2001 1777
tri 2001 1776 2002 1777 nw
tri 2424 1776 2425 1777 ne
rect 2425 1776 2517 1777
tri 2517 1776 2518 1777 nw
tri 2736 1776 2737 1777 ne
rect 2737 1776 2829 1777
tri 2829 1776 2830 1777 nw
tri 3252 1776 3253 1777 ne
rect 3253 1776 3345 1777
tri 3345 1776 3346 1777 nw
tri 3564 1776 3565 1777 ne
rect 3565 1776 3657 1777
tri 3657 1776 3658 1777 nw
tri 4080 1776 4081 1777 ne
rect 4081 1776 4173 1777
tri 4173 1776 4174 1777 nw
tri 4392 1776 4393 1777 ne
rect 4393 1776 4485 1777
tri 4485 1776 4486 1777 nw
tri 4908 1776 4909 1777 ne
rect 4909 1776 5001 1777
tri 5001 1776 5002 1777 nw
tri 5220 1776 5221 1777 ne
rect 5221 1776 5290 1777
rect 792 1742 798 1776
rect 832 1742 838 1776
tri 838 1753 861 1776 nw
tri 1081 1753 1104 1776 ne
rect 792 1704 838 1742
rect 1104 1742 1110 1776
rect 1144 1742 1150 1776
tri 1150 1753 1173 1776 nw
tri 1597 1753 1620 1776 ne
tri 838 1704 853 1719 sw
tri 1089 1704 1104 1719 se
rect 1104 1704 1150 1742
rect 1620 1742 1626 1776
rect 1660 1742 1666 1776
tri 1666 1753 1689 1776 nw
tri 1909 1753 1932 1776 ne
tri 1150 1704 1165 1719 sw
tri 1605 1704 1620 1719 se
rect 1620 1704 1666 1742
rect 1932 1742 1938 1776
rect 1972 1742 1978 1776
tri 1978 1753 2001 1776 nw
tri 2425 1753 2448 1776 ne
tri 1666 1704 1681 1719 sw
tri 1917 1704 1932 1719 se
rect 1932 1704 1978 1742
rect 2448 1742 2454 1776
rect 2488 1742 2494 1776
tri 2494 1753 2517 1776 nw
tri 2737 1753 2760 1776 ne
tri 1978 1704 1993 1719 sw
tri 2433 1704 2448 1719 se
rect 2448 1704 2494 1742
rect 2760 1742 2766 1776
rect 2800 1742 2806 1776
tri 2806 1753 2829 1776 nw
tri 3253 1753 3276 1776 ne
tri 2494 1704 2509 1719 sw
tri 2745 1704 2760 1719 se
rect 2760 1704 2806 1742
rect 3276 1742 3282 1776
rect 3316 1742 3322 1776
tri 3322 1753 3345 1776 nw
tri 3565 1753 3588 1776 ne
tri 2806 1704 2821 1719 sw
tri 3261 1704 3276 1719 se
rect 3276 1704 3322 1742
rect 3588 1742 3594 1776
rect 3628 1742 3634 1776
tri 3634 1753 3657 1776 nw
tri 4081 1753 4104 1776 ne
tri 3322 1704 3337 1719 sw
tri 3573 1704 3588 1719 se
rect 3588 1704 3634 1742
rect 4104 1742 4110 1776
rect 4144 1742 4150 1776
tri 4150 1753 4173 1776 nw
tri 4393 1753 4416 1776 ne
tri 3634 1704 3649 1719 sw
tri 4089 1704 4104 1719 se
rect 4104 1704 4150 1742
rect 4416 1742 4422 1776
rect 4456 1742 4462 1776
tri 4462 1753 4485 1776 nw
tri 4909 1753 4932 1776 ne
tri 4150 1704 4165 1719 sw
tri 4401 1704 4416 1719 se
rect 4416 1704 4462 1742
rect 4932 1742 4938 1776
rect 4972 1742 4978 1776
tri 4978 1753 5001 1776 nw
tri 5221 1753 5244 1776 ne
tri 4462 1704 4477 1719 sw
tri 4917 1704 4932 1719 se
rect 4932 1704 4978 1742
rect 5244 1742 5250 1776
rect 5284 1742 5290 1776
tri 4978 1704 4993 1719 sw
tri 5229 1704 5244 1719 se
rect 5244 1704 5290 1742
rect 792 1670 798 1704
rect 832 1694 853 1704
tri 853 1694 863 1704 sw
tri 1079 1694 1089 1704 se
rect 1089 1694 1110 1704
rect 832 1670 1110 1694
rect 1144 1694 1165 1704
tri 1165 1694 1175 1704 sw
tri 1595 1694 1605 1704 se
rect 1605 1694 1626 1704
rect 1144 1670 1626 1694
rect 1660 1694 1681 1704
tri 1681 1694 1691 1704 sw
tri 1907 1694 1917 1704 se
rect 1917 1694 1938 1704
rect 1660 1670 1938 1694
rect 1972 1694 1993 1704
tri 1993 1694 2003 1704 sw
tri 2423 1694 2433 1704 se
rect 2433 1694 2454 1704
rect 1972 1670 2454 1694
rect 2488 1694 2509 1704
tri 2509 1694 2519 1704 sw
tri 2735 1694 2745 1704 se
rect 2745 1694 2766 1704
rect 2488 1670 2766 1694
rect 2800 1694 2821 1704
tri 2821 1694 2831 1704 sw
tri 3251 1694 3261 1704 se
rect 3261 1694 3282 1704
rect 2800 1670 3282 1694
rect 3316 1694 3337 1704
tri 3337 1694 3347 1704 sw
tri 3563 1694 3573 1704 se
rect 3573 1694 3594 1704
rect 3316 1670 3594 1694
rect 3628 1694 3649 1704
tri 3649 1694 3659 1704 sw
tri 4079 1694 4089 1704 se
rect 4089 1694 4110 1704
rect 3628 1670 4110 1694
rect 4144 1694 4165 1704
tri 4165 1694 4175 1704 sw
tri 4391 1694 4401 1704 se
rect 4401 1694 4422 1704
rect 4144 1670 4422 1694
rect 4456 1694 4477 1704
tri 4477 1694 4487 1704 sw
tri 4907 1694 4917 1704 se
rect 4917 1694 4938 1704
rect 4456 1670 4938 1694
rect 4972 1694 4993 1704
tri 4993 1694 5003 1704 sw
tri 5219 1694 5229 1704 se
rect 5229 1694 5250 1704
rect 4972 1670 5250 1694
rect 5284 1670 5290 1704
rect 792 1632 5290 1670
rect 792 1598 798 1632
rect 832 1598 1110 1632
rect 1144 1598 1626 1632
rect 1660 1598 1938 1632
rect 1972 1598 2454 1632
rect 2488 1598 2766 1632
rect 2800 1598 3282 1632
rect 3316 1598 3594 1632
rect 3628 1598 4110 1632
rect 4144 1598 4422 1632
rect 4456 1598 4938 1632
rect 4972 1598 5250 1632
rect 5284 1598 5290 1632
rect 792 1560 5290 1598
rect 792 1526 798 1560
rect 832 1526 1110 1560
rect 1144 1526 1626 1560
rect 1660 1526 1938 1560
rect 1972 1526 2454 1560
rect 2488 1526 2766 1560
rect 2800 1526 3282 1560
rect 3316 1526 3594 1560
rect 3628 1526 4110 1560
rect 4144 1526 4422 1560
rect 4456 1526 4938 1560
rect 4972 1526 5250 1560
rect 5284 1526 5290 1560
rect 792 1514 5290 1526
rect 792 1488 838 1514
tri 838 1489 863 1514 nw
tri 1079 1489 1104 1514 ne
rect 792 1454 798 1488
rect 832 1454 838 1488
rect 1104 1488 1150 1514
tri 1150 1489 1175 1514 nw
tri 1595 1489 1620 1514 ne
tri 838 1454 839 1455 sw
tri 1103 1454 1104 1455 se
rect 1104 1454 1110 1488
rect 1144 1454 1150 1488
rect 1620 1488 1666 1514
tri 1666 1489 1691 1514 nw
tri 1907 1489 1932 1514 ne
tri 1150 1454 1151 1455 sw
tri 1619 1454 1620 1455 se
rect 1620 1454 1626 1488
rect 1660 1454 1666 1488
rect 1932 1488 1978 1514
tri 1978 1489 2003 1514 nw
tri 2423 1489 2448 1514 ne
tri 1666 1454 1667 1455 sw
tri 1931 1454 1932 1455 se
rect 1932 1454 1938 1488
rect 1972 1454 1978 1488
rect 2448 1488 2494 1514
tri 2494 1489 2519 1514 nw
tri 2735 1489 2760 1514 ne
tri 1978 1454 1979 1455 sw
tri 2447 1454 2448 1455 se
rect 2448 1454 2454 1488
rect 2488 1454 2494 1488
rect 2760 1488 2806 1514
tri 2806 1489 2831 1514 nw
tri 3251 1489 3276 1514 ne
tri 2494 1454 2495 1455 sw
tri 2759 1454 2760 1455 se
rect 2760 1454 2766 1488
rect 2800 1454 2806 1488
rect 3276 1488 3322 1514
tri 3322 1489 3347 1514 nw
tri 3563 1489 3588 1514 ne
tri 2806 1454 2807 1455 sw
tri 3275 1454 3276 1455 se
rect 3276 1454 3282 1488
rect 3316 1454 3322 1488
rect 3588 1488 3634 1514
tri 3634 1489 3659 1514 nw
tri 4079 1489 4104 1514 ne
tri 3322 1454 3323 1455 sw
tri 3587 1454 3588 1455 se
rect 3588 1454 3594 1488
rect 3628 1454 3634 1488
rect 4104 1488 4150 1514
tri 4150 1489 4175 1514 nw
tri 4391 1489 4416 1514 ne
tri 3634 1454 3635 1455 sw
tri 4103 1454 4104 1455 se
rect 4104 1454 4110 1488
rect 4144 1454 4150 1488
rect 4416 1488 4462 1514
tri 4462 1489 4487 1514 nw
tri 4907 1489 4932 1514 ne
tri 4150 1454 4151 1455 sw
tri 4415 1454 4416 1455 se
rect 4416 1454 4422 1488
rect 4456 1454 4462 1488
rect 4932 1488 4978 1514
tri 4978 1489 5003 1514 nw
tri 5219 1489 5244 1514 ne
tri 4462 1454 4463 1455 sw
tri 4931 1454 4932 1455 se
rect 4932 1454 4938 1488
rect 4972 1454 4978 1488
rect 5244 1488 5290 1514
tri 4978 1454 4979 1455 sw
tri 5243 1454 5244 1455 se
rect 5244 1454 5250 1488
rect 5284 1454 5290 1488
rect 792 1451 839 1454
tri 839 1451 842 1454 sw
tri 1100 1451 1103 1454 se
rect 1103 1451 1151 1454
tri 1151 1451 1154 1454 sw
tri 1616 1451 1619 1454 se
rect 1619 1451 1667 1454
tri 1667 1451 1670 1454 sw
tri 1928 1451 1931 1454 se
rect 1931 1451 1979 1454
tri 1979 1451 1982 1454 sw
tri 2444 1451 2447 1454 se
rect 2447 1451 2495 1454
tri 2495 1451 2498 1454 sw
tri 2756 1451 2759 1454 se
rect 2759 1451 2807 1454
tri 2807 1451 2810 1454 sw
tri 3272 1451 3275 1454 se
rect 3275 1451 3323 1454
tri 3323 1451 3326 1454 sw
tri 3584 1451 3587 1454 se
rect 3587 1451 3635 1454
tri 3635 1451 3638 1454 sw
tri 4100 1451 4103 1454 se
rect 4103 1451 4151 1454
tri 4151 1451 4154 1454 sw
tri 4412 1451 4415 1454 se
rect 4415 1451 4463 1454
tri 4463 1451 4466 1454 sw
tri 4928 1451 4931 1454 se
rect 4931 1451 4979 1454
tri 4979 1451 4982 1454 sw
tri 5240 1451 5243 1454 se
rect 5243 1451 5290 1454
rect 792 1446 842 1451
tri 842 1446 847 1451 sw
tri 1095 1446 1100 1451 se
rect 1100 1446 1154 1451
tri 1154 1446 1159 1451 sw
tri 1611 1446 1616 1451 se
rect 1616 1446 1670 1451
tri 1670 1446 1675 1451 sw
tri 1923 1446 1928 1451 se
rect 1928 1446 1982 1451
tri 1982 1446 1987 1451 sw
tri 2439 1446 2444 1451 se
rect 2444 1446 2498 1451
tri 2498 1446 2503 1451 sw
tri 2751 1446 2756 1451 se
rect 2756 1446 2810 1451
tri 2810 1446 2815 1451 sw
tri 3267 1446 3272 1451 se
rect 3272 1446 3326 1451
tri 3326 1446 3331 1451 sw
tri 3579 1446 3584 1451 se
rect 3584 1446 3638 1451
tri 3638 1446 3643 1451 sw
tri 4095 1446 4100 1451 se
rect 4100 1446 4154 1451
tri 4154 1446 4159 1451 sw
tri 4407 1446 4412 1451 se
rect 4412 1446 4466 1451
tri 4466 1446 4471 1451 sw
tri 4923 1446 4928 1451 se
rect 4928 1446 4982 1451
tri 4982 1446 4987 1451 sw
tri 5235 1446 5240 1451 se
rect 5240 1446 5290 1451
rect 792 1430 847 1446
tri 847 1430 863 1446 sw
tri 1079 1430 1095 1446 se
rect 1095 1430 1159 1446
tri 1159 1430 1175 1446 sw
tri 1595 1430 1611 1446 se
rect 1611 1430 1675 1446
tri 1675 1430 1691 1446 sw
tri 1907 1430 1923 1446 se
rect 1923 1430 1987 1446
tri 1987 1430 2003 1446 sw
tri 2423 1430 2439 1446 se
rect 2439 1430 2503 1446
tri 2503 1430 2519 1446 sw
tri 2735 1430 2751 1446 se
rect 2751 1430 2815 1446
tri 2815 1430 2831 1446 sw
tri 3251 1430 3267 1446 se
rect 3267 1430 3331 1446
tri 3331 1430 3347 1446 sw
tri 3563 1430 3579 1446 se
rect 3579 1430 3643 1446
tri 3643 1430 3659 1446 sw
tri 4079 1430 4095 1446 se
rect 4095 1430 4159 1446
tri 4159 1430 4175 1446 sw
tri 4391 1430 4407 1446 se
rect 4407 1430 4471 1446
tri 4471 1430 4487 1446 sw
tri 4907 1430 4923 1446 se
rect 4923 1430 4987 1446
tri 4987 1430 5003 1446 sw
tri 5219 1430 5235 1446 se
rect 5235 1430 5290 1446
rect 792 1416 5290 1430
rect 792 1382 798 1416
rect 832 1382 1110 1416
rect 1144 1382 1626 1416
rect 1660 1382 1938 1416
rect 1972 1382 2454 1416
rect 2488 1382 2766 1416
rect 2800 1382 3282 1416
rect 3316 1382 3594 1416
rect 3628 1382 4110 1416
rect 4144 1382 4422 1416
rect 4456 1382 4938 1416
rect 4972 1382 5250 1416
rect 5284 1382 5290 1416
rect 792 1344 5290 1382
rect 792 1310 798 1344
rect 832 1310 1110 1344
rect 1144 1310 1626 1344
rect 1660 1310 1938 1344
rect 1972 1310 2454 1344
rect 2488 1310 2766 1344
rect 2800 1310 3282 1344
rect 3316 1310 3594 1344
rect 3628 1310 4110 1344
rect 4144 1310 4422 1344
rect 4456 1310 4938 1344
rect 4972 1310 5250 1344
rect 5284 1310 5290 1344
rect 792 1272 5290 1310
rect 792 1238 798 1272
rect 832 1250 1110 1272
rect 832 1238 851 1250
tri 851 1238 863 1250 nw
tri 1079 1238 1091 1250 ne
rect 1091 1238 1110 1250
rect 1144 1250 1626 1272
rect 1144 1238 1163 1250
tri 1163 1238 1175 1250 nw
tri 1595 1238 1607 1250 ne
rect 1607 1238 1626 1250
rect 1660 1250 1938 1272
rect 1660 1238 1679 1250
tri 1679 1238 1691 1250 nw
tri 1907 1238 1919 1250 ne
rect 1919 1238 1938 1250
rect 1972 1250 2454 1272
rect 1972 1238 1991 1250
tri 1991 1238 2003 1250 nw
tri 2423 1238 2435 1250 ne
rect 2435 1238 2454 1250
rect 2488 1250 2766 1272
rect 2488 1238 2507 1250
tri 2507 1238 2519 1250 nw
tri 2735 1238 2747 1250 ne
rect 2747 1238 2766 1250
rect 2800 1250 3282 1272
rect 2800 1238 2819 1250
tri 2819 1238 2831 1250 nw
tri 3251 1238 3263 1250 ne
rect 3263 1238 3282 1250
rect 3316 1250 3594 1272
rect 3316 1238 3335 1250
tri 3335 1238 3347 1250 nw
tri 3563 1238 3575 1250 ne
rect 3575 1238 3594 1250
rect 3628 1250 4110 1272
rect 3628 1238 3647 1250
tri 3647 1238 3659 1250 nw
tri 4079 1238 4091 1250 ne
rect 4091 1238 4110 1250
rect 4144 1250 4422 1272
rect 4144 1238 4163 1250
tri 4163 1238 4175 1250 nw
tri 4391 1238 4403 1250 ne
rect 4403 1238 4422 1250
rect 4456 1250 4938 1272
rect 4456 1238 4475 1250
tri 4475 1238 4487 1250 nw
tri 4907 1238 4919 1250 ne
rect 4919 1238 4938 1250
rect 4972 1250 5250 1272
rect 4972 1238 4991 1250
tri 4991 1238 5003 1250 nw
tri 5219 1238 5231 1250 ne
rect 5231 1238 5250 1250
rect 5284 1238 5290 1272
rect 792 1232 845 1238
tri 845 1232 851 1238 nw
tri 1091 1232 1097 1238 ne
rect 1097 1232 1157 1238
tri 1157 1232 1163 1238 nw
tri 1607 1232 1613 1238 ne
rect 1613 1232 1673 1238
tri 1673 1232 1679 1238 nw
tri 1919 1232 1925 1238 ne
rect 1925 1232 1985 1238
tri 1985 1232 1991 1238 nw
tri 2435 1232 2441 1238 ne
rect 2441 1232 2501 1238
tri 2501 1232 2507 1238 nw
tri 2747 1232 2753 1238 ne
rect 2753 1232 2813 1238
tri 2813 1232 2819 1238 nw
tri 3263 1232 3269 1238 ne
rect 3269 1232 3329 1238
tri 3329 1232 3335 1238 nw
tri 3575 1232 3581 1238 ne
rect 3581 1232 3641 1238
tri 3641 1232 3647 1238 nw
tri 4091 1232 4097 1238 ne
rect 4097 1232 4157 1238
tri 4157 1232 4163 1238 nw
tri 4403 1232 4409 1238 ne
rect 4409 1232 4469 1238
tri 4469 1232 4475 1238 nw
tri 4919 1232 4925 1238 ne
rect 4925 1232 4985 1238
tri 4985 1232 4991 1238 nw
tri 5231 1232 5237 1238 ne
rect 5237 1232 5290 1238
rect 792 1227 840 1232
tri 840 1227 845 1232 nw
tri 1097 1227 1102 1232 ne
rect 1102 1227 1152 1232
tri 1152 1227 1157 1232 nw
tri 1613 1227 1618 1232 ne
rect 1618 1227 1668 1232
tri 1668 1227 1673 1232 nw
tri 1925 1227 1930 1232 ne
rect 1930 1227 1980 1232
tri 1980 1227 1985 1232 nw
tri 2441 1227 2446 1232 ne
rect 2446 1227 2496 1232
tri 2496 1227 2501 1232 nw
tri 2753 1227 2758 1232 ne
rect 2758 1227 2808 1232
tri 2808 1227 2813 1232 nw
tri 3269 1227 3274 1232 ne
rect 3274 1227 3324 1232
tri 3324 1227 3329 1232 nw
tri 3581 1227 3586 1232 ne
rect 3586 1227 3636 1232
tri 3636 1227 3641 1232 nw
tri 4097 1227 4102 1232 ne
rect 4102 1227 4152 1232
tri 4152 1227 4157 1232 nw
tri 4409 1227 4414 1232 ne
rect 4414 1227 4464 1232
tri 4464 1227 4469 1232 nw
tri 4925 1227 4930 1232 ne
rect 4930 1227 4980 1232
tri 4980 1227 4985 1232 nw
tri 5237 1227 5242 1232 ne
rect 5242 1227 5290 1232
rect 792 1200 838 1227
tri 838 1225 840 1227 nw
tri 1102 1225 1104 1227 ne
rect 792 1166 798 1200
rect 832 1166 838 1200
rect 1104 1200 1150 1227
tri 1150 1225 1152 1227 nw
tri 1618 1225 1620 1227 ne
tri 838 1166 863 1191 sw
tri 1079 1166 1104 1191 se
rect 1104 1166 1110 1200
rect 1144 1166 1150 1200
rect 1620 1200 1666 1227
tri 1666 1225 1668 1227 nw
tri 1930 1225 1932 1227 ne
tri 1150 1166 1175 1191 sw
tri 1595 1166 1620 1191 se
rect 1620 1166 1626 1200
rect 1660 1166 1666 1200
rect 1932 1200 1978 1227
tri 1978 1225 1980 1227 nw
tri 2446 1225 2448 1227 ne
tri 1666 1166 1691 1191 sw
tri 1907 1166 1932 1191 se
rect 1932 1166 1938 1200
rect 1972 1166 1978 1200
rect 2448 1200 2494 1227
tri 2494 1225 2496 1227 nw
tri 2758 1225 2760 1227 ne
tri 1978 1166 2003 1191 sw
tri 2423 1166 2448 1191 se
rect 2448 1166 2454 1200
rect 2488 1166 2494 1200
rect 2760 1200 2806 1227
tri 2806 1225 2808 1227 nw
tri 3274 1225 3276 1227 ne
tri 2494 1166 2519 1191 sw
tri 2735 1166 2760 1191 se
rect 2760 1166 2766 1200
rect 2800 1166 2806 1200
rect 3276 1200 3322 1227
tri 3322 1225 3324 1227 nw
tri 3586 1225 3588 1227 ne
tri 2806 1166 2831 1191 sw
tri 3251 1166 3276 1191 se
rect 3276 1166 3282 1200
rect 3316 1166 3322 1200
rect 3588 1200 3634 1227
tri 3634 1225 3636 1227 nw
tri 4102 1225 4104 1227 ne
tri 3322 1166 3347 1191 sw
tri 3563 1166 3588 1191 se
rect 3588 1166 3594 1200
rect 3628 1166 3634 1200
rect 4104 1200 4150 1227
tri 4150 1225 4152 1227 nw
tri 4414 1225 4416 1227 ne
tri 3634 1166 3659 1191 sw
tri 4079 1166 4104 1191 se
rect 4104 1166 4110 1200
rect 4144 1166 4150 1200
rect 4416 1200 4462 1227
tri 4462 1225 4464 1227 nw
tri 4930 1225 4932 1227 ne
tri 4150 1166 4175 1191 sw
tri 4391 1166 4416 1191 se
rect 4416 1166 4422 1200
rect 4456 1166 4462 1200
rect 4932 1200 4978 1227
tri 4978 1225 4980 1227 nw
tri 5242 1225 5244 1227 ne
tri 4462 1166 4487 1191 sw
tri 4907 1166 4932 1191 se
rect 4932 1166 4938 1200
rect 4972 1166 4978 1200
rect 5244 1200 5290 1227
tri 4978 1166 5003 1191 sw
tri 5219 1166 5244 1191 se
rect 5244 1166 5250 1200
rect 5284 1166 5290 1200
rect 792 1128 5290 1166
rect 792 1094 798 1128
rect 832 1094 1110 1128
rect 1144 1094 1626 1128
rect 1660 1094 1938 1128
rect 1972 1094 2454 1128
rect 2488 1094 2766 1128
rect 2800 1094 3282 1128
rect 3316 1094 3594 1128
rect 3628 1094 4110 1128
rect 4144 1094 4422 1128
rect 4456 1094 4938 1128
rect 4972 1094 5250 1128
rect 5284 1094 5290 1128
rect 792 1056 5290 1094
rect 792 1022 798 1056
rect 832 1022 1110 1056
rect 1144 1022 1626 1056
rect 1660 1022 1938 1056
rect 1972 1022 2454 1056
rect 2488 1022 2766 1056
rect 2800 1022 3282 1056
rect 3316 1022 3594 1056
rect 3628 1022 4110 1056
rect 4144 1022 4422 1056
rect 4456 1022 4938 1056
rect 4972 1022 5250 1056
rect 5284 1022 5290 1056
rect 792 986 5290 1022
rect 792 984 861 986
tri 861 984 863 986 nw
tri 1079 984 1081 986 ne
rect 1081 984 1173 986
tri 1173 984 1175 986 nw
tri 1595 984 1597 986 ne
rect 1597 984 1689 986
tri 1689 984 1691 986 nw
tri 1907 984 1909 986 ne
rect 1909 984 2001 986
tri 2001 984 2003 986 nw
tri 2423 984 2425 986 ne
rect 2425 984 2517 986
tri 2517 984 2519 986 nw
tri 2735 984 2737 986 ne
rect 2737 984 2829 986
tri 2829 984 2831 986 nw
tri 3251 984 3253 986 ne
rect 3253 984 3345 986
tri 3345 984 3347 986 nw
tri 3563 984 3565 986 ne
rect 3565 984 3657 986
tri 3657 984 3659 986 nw
tri 4079 984 4081 986 ne
rect 4081 984 4173 986
tri 4173 984 4175 986 nw
tri 4391 984 4393 986 ne
rect 4393 984 4485 986
tri 4485 984 4487 986 nw
tri 4907 984 4909 986 ne
rect 4909 984 5001 986
tri 5001 984 5003 986 nw
tri 5219 984 5221 986 ne
rect 5221 984 5290 986
rect 792 950 798 984
rect 832 950 838 984
tri 838 961 861 984 nw
tri 1081 961 1104 984 ne
rect 792 912 838 950
rect 1104 950 1110 984
rect 1144 950 1150 984
tri 1150 961 1173 984 nw
tri 1597 961 1620 984 ne
tri 838 912 853 927 sw
tri 1089 912 1104 927 se
rect 1104 912 1150 950
rect 1620 950 1626 984
rect 1660 950 1666 984
tri 1666 961 1689 984 nw
tri 1909 961 1932 984 ne
tri 1150 912 1165 927 sw
tri 1605 912 1620 927 se
rect 1620 912 1666 950
rect 1932 950 1938 984
rect 1972 950 1978 984
tri 1978 961 2001 984 nw
tri 2425 961 2448 984 ne
tri 1666 912 1681 927 sw
tri 1917 912 1932 927 se
rect 1932 912 1978 950
rect 2448 950 2454 984
rect 2488 950 2494 984
tri 2494 961 2517 984 nw
tri 2737 961 2760 984 ne
tri 1978 912 1993 927 sw
tri 2433 912 2448 927 se
rect 2448 912 2494 950
rect 2760 950 2766 984
rect 2800 950 2806 984
tri 2806 961 2829 984 nw
tri 3253 961 3276 984 ne
tri 2494 912 2509 927 sw
tri 2745 912 2760 927 se
rect 2760 912 2806 950
rect 3276 950 3282 984
rect 3316 950 3322 984
tri 3322 961 3345 984 nw
tri 3565 961 3588 984 ne
tri 2806 912 2821 927 sw
tri 3261 912 3276 927 se
rect 3276 912 3322 950
rect 3588 950 3594 984
rect 3628 950 3634 984
tri 3634 961 3657 984 nw
tri 4081 961 4104 984 ne
tri 3322 912 3337 927 sw
tri 3573 912 3588 927 se
rect 3588 912 3634 950
rect 4104 950 4110 984
rect 4144 950 4150 984
tri 4150 961 4173 984 nw
tri 4393 961 4416 984 ne
tri 3634 912 3649 927 sw
tri 4089 912 4104 927 se
rect 4104 912 4150 950
rect 4416 950 4422 984
rect 4456 950 4462 984
tri 4462 961 4485 984 nw
tri 4909 961 4932 984 ne
tri 4150 912 4165 927 sw
tri 4401 912 4416 927 se
rect 4416 912 4462 950
rect 4932 950 4938 984
rect 4972 950 4978 984
tri 4978 961 5001 984 nw
tri 5221 961 5244 984 ne
tri 4462 912 4477 927 sw
tri 4917 912 4932 927 se
rect 4932 912 4978 950
rect 5244 950 5250 984
rect 5284 950 5290 984
tri 4978 912 4993 927 sw
tri 5229 912 5244 927 se
rect 5244 912 5290 950
rect 792 878 798 912
rect 832 902 853 912
tri 853 902 863 912 sw
tri 1079 902 1089 912 se
rect 1089 902 1110 912
rect 832 878 1110 902
rect 1144 902 1165 912
tri 1165 902 1175 912 sw
tri 1595 902 1605 912 se
rect 1605 902 1626 912
rect 1144 878 1626 902
rect 1660 902 1681 912
tri 1681 902 1691 912 sw
tri 1907 902 1917 912 se
rect 1917 902 1938 912
rect 1660 878 1938 902
rect 1972 902 1993 912
tri 1993 902 2003 912 sw
tri 2423 902 2433 912 se
rect 2433 902 2454 912
rect 1972 878 2454 902
rect 2488 902 2509 912
tri 2509 902 2519 912 sw
tri 2735 902 2745 912 se
rect 2745 902 2766 912
rect 2488 878 2766 902
rect 2800 902 2821 912
tri 2821 902 2831 912 sw
tri 3251 902 3261 912 se
rect 3261 902 3282 912
rect 2800 878 3282 902
rect 3316 902 3337 912
tri 3337 902 3347 912 sw
tri 3563 902 3573 912 se
rect 3573 902 3594 912
rect 3316 878 3594 902
rect 3628 902 3649 912
tri 3649 902 3659 912 sw
tri 4079 902 4089 912 se
rect 4089 902 4110 912
rect 3628 878 4110 902
rect 4144 902 4165 912
tri 4165 902 4175 912 sw
tri 4391 902 4401 912 se
rect 4401 902 4422 912
rect 4144 878 4422 902
rect 4456 902 4477 912
tri 4477 902 4487 912 sw
tri 4907 902 4917 912 se
rect 4917 902 4938 912
rect 4456 878 4938 902
rect 4972 902 4993 912
tri 4993 902 5003 912 sw
tri 5219 902 5229 912 se
rect 5229 902 5250 912
rect 4972 878 5250 902
rect 5284 878 5290 912
rect 792 840 5290 878
rect 792 806 798 840
rect 832 806 1110 840
rect 1144 806 1626 840
rect 1660 806 1938 840
rect 1972 806 2454 840
rect 2488 806 2766 840
rect 2800 806 3282 840
rect 3316 806 3594 840
rect 3628 806 4110 840
rect 4144 806 4422 840
rect 4456 806 4938 840
rect 4972 806 5250 840
rect 5284 806 5290 840
rect 792 768 5290 806
rect 792 734 798 768
rect 832 734 1110 768
rect 1144 734 1626 768
rect 1660 734 1938 768
rect 1972 734 2454 768
rect 2488 734 2766 768
rect 2800 734 3282 768
rect 3316 734 3594 768
rect 3628 734 4110 768
rect 4144 734 4422 768
rect 4456 734 4938 768
rect 4972 734 5250 768
rect 5284 734 5290 768
rect 792 722 5290 734
rect 5444 2215 5450 2249
rect 5484 2222 5594 2249
rect 5628 2222 5666 2256
rect 5700 2222 5712 2256
rect 5484 2215 5712 2222
rect 5444 2181 5522 2215
rect 5556 2183 5712 2215
rect 5556 2181 5594 2183
rect 5444 2176 5594 2181
rect 5444 2142 5450 2176
rect 5484 2149 5594 2176
rect 5628 2149 5666 2183
rect 5700 2149 5712 2183
rect 5484 2142 5712 2149
rect 5444 2108 5522 2142
rect 5556 2110 5712 2142
rect 5556 2108 5594 2110
rect 5444 2103 5594 2108
rect 5444 2069 5450 2103
rect 5484 2076 5594 2103
rect 5628 2076 5666 2110
rect 5700 2076 5712 2110
rect 5484 2069 5712 2076
rect 5444 2035 5522 2069
rect 5556 2037 5712 2069
rect 5556 2035 5594 2037
rect 5444 2030 5594 2035
rect 5444 1996 5450 2030
rect 5484 2003 5594 2030
rect 5628 2003 5666 2037
rect 5700 2003 5712 2037
rect 5484 1996 5712 2003
rect 5444 1962 5522 1996
rect 5556 1964 5712 1996
rect 5556 1962 5594 1964
rect 5444 1957 5594 1962
rect 5444 1923 5450 1957
rect 5484 1930 5594 1957
rect 5628 1930 5666 1964
rect 5700 1930 5712 1964
rect 5484 1923 5712 1930
rect 5444 1889 5522 1923
rect 5556 1891 5712 1923
rect 5556 1889 5594 1891
rect 5444 1884 5594 1889
rect 5444 1850 5450 1884
rect 5484 1857 5594 1884
rect 5628 1857 5666 1891
rect 5700 1857 5712 1891
rect 5484 1850 5712 1857
rect 5444 1816 5522 1850
rect 5556 1818 5712 1850
rect 5556 1816 5594 1818
rect 5444 1811 5594 1816
rect 5444 1777 5450 1811
rect 5484 1784 5594 1811
rect 5628 1784 5666 1818
rect 5700 1784 5712 1818
rect 5484 1777 5712 1784
rect 5444 1743 5522 1777
rect 5556 1745 5712 1777
rect 5556 1743 5594 1745
rect 5444 1738 5594 1743
rect 5444 1704 5450 1738
rect 5484 1711 5594 1738
rect 5628 1711 5666 1745
rect 5700 1711 5712 1745
rect 5484 1704 5712 1711
rect 5444 1670 5522 1704
rect 5556 1672 5712 1704
rect 5556 1670 5594 1672
rect 5444 1665 5594 1670
rect 5444 1631 5450 1665
rect 5484 1638 5594 1665
rect 5628 1638 5666 1672
rect 5700 1638 5712 1672
rect 5484 1631 5712 1638
rect 5444 1597 5522 1631
rect 5556 1599 5712 1631
rect 5556 1597 5594 1599
rect 5444 1592 5594 1597
rect 5444 1558 5450 1592
rect 5484 1565 5594 1592
rect 5628 1565 5666 1599
rect 5700 1565 5712 1599
rect 5484 1558 5712 1565
rect 5444 1524 5522 1558
rect 5556 1526 5712 1558
rect 5556 1524 5594 1526
rect 5444 1519 5594 1524
rect 5444 1485 5450 1519
rect 5484 1492 5594 1519
rect 5628 1492 5666 1526
rect 5700 1492 5712 1526
rect 5484 1485 5712 1492
rect 5444 1451 5522 1485
rect 5556 1453 5712 1485
rect 5556 1451 5594 1453
rect 5444 1446 5594 1451
rect 5444 1412 5450 1446
rect 5484 1419 5594 1446
rect 5628 1419 5666 1453
rect 5700 1419 5712 1453
rect 5484 1412 5712 1419
rect 5444 1378 5522 1412
rect 5556 1380 5712 1412
rect 5556 1378 5594 1380
rect 5444 1373 5594 1378
rect 5444 1339 5450 1373
rect 5484 1346 5594 1373
rect 5628 1346 5666 1380
rect 5700 1346 5712 1380
rect 5484 1339 5712 1346
rect 5444 1305 5522 1339
rect 5556 1307 5712 1339
rect 5556 1305 5594 1307
rect 5444 1300 5594 1305
rect 5444 1266 5450 1300
rect 5484 1273 5594 1300
rect 5628 1273 5666 1307
rect 5700 1273 5712 1307
rect 5484 1266 5712 1273
rect 5444 1232 5522 1266
rect 5556 1234 5712 1266
rect 5556 1232 5594 1234
rect 5444 1227 5594 1232
rect 5444 1193 5450 1227
rect 5484 1200 5594 1227
rect 5628 1200 5666 1234
rect 5700 1200 5712 1234
rect 5484 1193 5712 1200
rect 5444 1159 5522 1193
rect 5556 1161 5712 1193
rect 5556 1159 5594 1161
rect 5444 1154 5594 1159
rect 5444 1120 5450 1154
rect 5484 1127 5594 1154
rect 5628 1127 5666 1161
rect 5700 1127 5712 1161
rect 5484 1120 5712 1127
rect 5444 1086 5522 1120
rect 5556 1088 5712 1120
rect 5556 1086 5594 1088
rect 5444 1081 5594 1086
rect 5444 1047 5450 1081
rect 5484 1054 5594 1081
rect 5628 1054 5666 1088
rect 5700 1054 5712 1088
rect 5484 1047 5712 1054
rect 5444 1013 5522 1047
rect 5556 1015 5712 1047
rect 5556 1013 5594 1015
rect 5444 1008 5594 1013
rect 5444 974 5450 1008
rect 5484 981 5594 1008
rect 5628 981 5666 1015
rect 5700 981 5712 1015
rect 5484 974 5712 981
rect 5444 940 5522 974
rect 5556 942 5712 974
rect 5556 940 5594 942
rect 5444 935 5594 940
rect 5444 901 5450 935
rect 5484 908 5594 935
rect 5628 908 5666 942
rect 5700 908 5712 942
rect 5484 901 5712 908
rect 5444 867 5522 901
rect 5556 869 5712 901
rect 5556 867 5594 869
rect 5444 862 5594 867
rect 5444 828 5450 862
rect 5484 835 5594 862
rect 5628 835 5666 869
rect 5700 835 5712 869
rect 5484 828 5712 835
rect 5444 794 5522 828
rect 5556 796 5712 828
rect 5556 794 5594 796
rect 5444 789 5594 794
rect 5444 755 5450 789
rect 5484 762 5594 789
rect 5628 762 5666 796
rect 5700 762 5712 796
rect 5484 755 5712 762
rect 488 716 638 718
rect 488 689 598 716
rect 370 682 598 689
rect 632 682 638 716
rect 5444 721 5522 755
rect 5556 723 5712 755
rect 5556 721 5594 723
rect 5444 716 5594 721
rect 5444 682 5450 716
rect 5484 689 5594 716
rect 5628 689 5666 723
rect 5700 689 5712 723
rect 5484 682 5712 689
rect 370 680 638 682
rect 370 650 526 680
rect 370 616 382 650
rect 416 616 454 650
rect 488 646 526 650
rect 560 646 638 680
rect 488 643 638 646
rect 488 616 598 643
rect 370 609 598 616
rect 632 609 638 643
rect 676 676 5407 682
rect 676 642 688 676
rect 722 642 764 676
rect 798 642 840 676
rect 874 642 916 676
rect 950 642 992 676
rect 1026 642 1068 676
rect 1102 642 1144 676
rect 1178 642 1221 676
rect 1255 642 1516 676
rect 1550 642 1592 676
rect 1626 642 1668 676
rect 1702 642 1744 676
rect 1778 642 1820 676
rect 1854 642 1896 676
rect 1930 642 1972 676
rect 2006 642 2049 676
rect 2083 642 2344 676
rect 2378 642 2420 676
rect 2454 642 2496 676
rect 2530 642 2572 676
rect 2606 642 2648 676
rect 2682 642 2724 676
rect 2758 642 2800 676
rect 2834 642 2877 676
rect 2911 642 3172 676
rect 3206 642 3248 676
rect 3282 642 3324 676
rect 3358 642 3400 676
rect 3434 642 3476 676
rect 3510 642 3552 676
rect 3586 642 3628 676
rect 3662 642 3705 676
rect 3739 642 4000 676
rect 4034 642 4076 676
rect 4110 642 4152 676
rect 4186 642 4228 676
rect 4262 642 4304 676
rect 4338 642 4380 676
rect 4414 642 4456 676
rect 4490 642 4533 676
rect 4567 642 4828 676
rect 4862 642 4904 676
rect 4938 642 4980 676
rect 5014 642 5056 676
rect 5090 642 5132 676
rect 5166 642 5208 676
rect 5242 642 5284 676
rect 5318 642 5361 676
rect 5395 642 5407 676
rect 676 630 5407 642
rect 5444 648 5522 682
rect 5556 650 5712 682
rect 5556 648 5594 650
rect 5444 643 5594 648
rect 370 608 638 609
tri 370 604 374 608 ne
rect 374 604 526 608
tri 374 574 404 604 ne
rect 404 574 526 604
rect 560 576 638 608
rect 5444 609 5450 643
rect 5484 616 5594 643
rect 5628 616 5666 650
rect 5700 616 5712 650
rect 5484 609 5706 616
tri 5706 610 5712 616 nw
rect 5974 4218 5980 4603
rect 6086 4218 6092 4612
rect 5974 4180 6092 4218
rect 5974 4179 6052 4180
rect 5974 4145 5980 4179
rect 6014 4146 6052 4179
rect 6086 4146 6092 4180
rect 6014 4145 6092 4146
rect 5974 4108 6092 4145
rect 5974 4106 6052 4108
rect 5974 4072 5980 4106
rect 6014 4074 6052 4106
rect 6086 4074 6092 4108
rect 6014 4072 6092 4074
rect 5974 4036 6092 4072
rect 5974 4033 6052 4036
rect 5974 3999 5980 4033
rect 6014 4002 6052 4033
rect 6086 4002 6092 4036
rect 6014 3999 6092 4002
rect 5974 3964 6092 3999
rect 5974 3960 6052 3964
rect 5974 3926 5980 3960
rect 6014 3930 6052 3960
rect 6086 3930 6092 3964
rect 6014 3926 6092 3930
rect 5974 3892 6092 3926
rect 5974 3887 6052 3892
rect 5974 3853 5980 3887
rect 6014 3858 6052 3887
rect 6086 3858 6092 3892
rect 6014 3853 6092 3858
rect 5974 3820 6092 3853
rect 5974 3814 6052 3820
rect 5974 3780 5980 3814
rect 6014 3786 6052 3814
rect 6086 3786 6092 3820
rect 6014 3780 6092 3786
rect 5974 3748 6092 3780
rect 5974 3741 6052 3748
rect 5974 3707 5980 3741
rect 6014 3714 6052 3741
rect 6086 3714 6092 3748
rect 6014 3707 6092 3714
rect 5974 3676 6092 3707
rect 5974 3668 6052 3676
rect 5974 3634 5980 3668
rect 6014 3642 6052 3668
rect 6086 3642 6092 3676
rect 6014 3634 6092 3642
rect 5974 3604 6092 3634
rect 5974 3595 6052 3604
rect 5974 3561 5980 3595
rect 6014 3570 6052 3595
rect 6086 3570 6092 3604
rect 6014 3561 6092 3570
rect 5974 3532 6092 3561
rect 5974 3522 6052 3532
rect 5974 3488 5980 3522
rect 6014 3498 6052 3522
rect 6086 3498 6092 3532
rect 6014 3488 6092 3498
rect 5974 3460 6092 3488
rect 5974 3449 6052 3460
rect 5974 3415 5980 3449
rect 6014 3426 6052 3449
rect 6086 3426 6092 3460
rect 6014 3415 6092 3426
rect 5974 3388 6092 3415
rect 5974 3376 6052 3388
rect 5974 3342 5980 3376
rect 6014 3354 6052 3376
rect 6086 3354 6092 3388
rect 6014 3342 6092 3354
rect 5974 3316 6092 3342
rect 5974 3303 6052 3316
rect 5974 3269 5980 3303
rect 6014 3282 6052 3303
rect 6086 3282 6092 3316
rect 6014 3269 6092 3282
rect 5974 3244 6092 3269
rect 5974 3230 6052 3244
rect 5974 3196 5980 3230
rect 6014 3210 6052 3230
rect 6086 3210 6092 3244
rect 6014 3196 6092 3210
rect 5974 3172 6092 3196
rect 5974 3157 6052 3172
rect 5974 3123 5980 3157
rect 6014 3138 6052 3157
rect 6086 3138 6092 3172
rect 6014 3123 6092 3138
rect 5974 3100 6092 3123
rect 5974 3084 6052 3100
rect 5974 3050 5980 3084
rect 6014 3066 6052 3084
rect 6086 3066 6092 3100
rect 6014 3050 6092 3066
rect 5974 3028 6092 3050
rect 5974 3011 6052 3028
rect 5974 2977 5980 3011
rect 6014 2994 6052 3011
rect 6086 2994 6092 3028
rect 6014 2977 6092 2994
rect 5974 2956 6092 2977
rect 5974 2938 6052 2956
rect 5974 2904 5980 2938
rect 6014 2922 6052 2938
rect 6086 2922 6092 2956
rect 6014 2904 6092 2922
rect 5974 2884 6092 2904
rect 5974 2865 6052 2884
rect 5974 2831 5980 2865
rect 6014 2850 6052 2865
rect 6086 2850 6092 2884
rect 6014 2831 6092 2850
rect 5974 2812 6092 2831
rect 5974 2792 6052 2812
rect 5974 2758 5980 2792
rect 6014 2778 6052 2792
rect 6086 2778 6092 2812
rect 6014 2758 6092 2778
rect 5974 2740 6092 2758
rect 5974 2719 6052 2740
rect 5974 2685 5980 2719
rect 6014 2706 6052 2719
rect 6086 2706 6092 2740
rect 6014 2685 6092 2706
rect 5974 2668 6092 2685
rect 5974 2646 6052 2668
rect 5974 2612 5980 2646
rect 6014 2634 6052 2646
rect 6086 2634 6092 2668
rect 6014 2612 6092 2634
rect 5974 2596 6092 2612
rect 5974 2573 6052 2596
rect 5974 2539 5980 2573
rect 6014 2562 6052 2573
rect 6086 2562 6092 2596
rect 6014 2539 6092 2562
rect 5974 2524 6092 2539
rect 5974 2500 6052 2524
rect 5974 2466 5980 2500
rect 6014 2490 6052 2500
rect 6086 2490 6092 2524
rect 6014 2466 6092 2490
rect 5974 2452 6092 2466
rect 5974 2427 6052 2452
rect 5974 2393 5980 2427
rect 6014 2418 6052 2427
rect 6086 2418 6092 2452
rect 6014 2393 6092 2418
rect 5974 2380 6092 2393
rect 5974 2354 6052 2380
rect 5974 2320 5980 2354
rect 6014 2346 6052 2354
rect 6086 2346 6092 2380
rect 6014 2320 6092 2346
rect 5974 2308 6092 2320
rect 5974 2281 6052 2308
rect 5974 2247 5980 2281
rect 6014 2274 6052 2281
rect 6086 2274 6092 2308
rect 6014 2247 6092 2274
rect 5974 2236 6092 2247
rect 5974 2208 6052 2236
rect 5974 2174 5980 2208
rect 6014 2202 6052 2208
rect 6086 2202 6092 2236
rect 6014 2174 6092 2202
rect 5974 2164 6092 2174
rect 5974 2135 6052 2164
rect 5974 2101 5980 2135
rect 6014 2130 6052 2135
rect 6086 2130 6092 2164
rect 6014 2101 6092 2130
rect 5974 2092 6092 2101
rect 5974 2062 6052 2092
rect 5974 2028 5980 2062
rect 6014 2058 6052 2062
rect 6086 2058 6092 2092
rect 6014 2028 6092 2058
rect 5974 2020 6092 2028
rect 5974 1989 6052 2020
rect 5974 1955 5980 1989
rect 6014 1986 6052 1989
rect 6086 1986 6092 2020
rect 6014 1955 6092 1986
rect 5974 1948 6092 1955
rect 5974 1916 6052 1948
rect 5974 1882 5980 1916
rect 6014 1914 6052 1916
rect 6086 1914 6092 1948
rect 6014 1882 6092 1914
rect 5974 1876 6092 1882
rect 5974 1843 6052 1876
rect 5974 1809 5980 1843
rect 6014 1842 6052 1843
rect 6086 1842 6092 1876
rect 6014 1809 6092 1842
rect 5974 1804 6092 1809
rect 5974 1770 6052 1804
rect 6086 1770 6092 1804
rect 5974 1736 5980 1770
rect 6014 1736 6092 1770
rect 5974 1732 6092 1736
rect 5974 1698 6052 1732
rect 6086 1698 6092 1732
rect 5974 1697 6092 1698
rect 5974 1663 5980 1697
rect 6014 1663 6092 1697
rect 5974 1660 6092 1663
rect 5974 1626 6052 1660
rect 6086 1626 6092 1660
rect 5974 1624 6092 1626
rect 5974 1590 5980 1624
rect 6014 1590 6092 1624
rect 5974 1588 6092 1590
rect 5974 1554 6052 1588
rect 6086 1554 6092 1588
rect 5974 1551 6092 1554
rect 5974 1517 5980 1551
rect 6014 1517 6092 1551
rect 5974 1516 6092 1517
rect 5974 1482 6052 1516
rect 6086 1482 6092 1516
rect 5974 1478 6092 1482
rect 5974 1444 5980 1478
rect 6014 1444 6092 1478
rect 5974 1410 6052 1444
rect 6086 1410 6092 1444
rect 5974 1405 6092 1410
rect 5974 1371 5980 1405
rect 6014 1371 6092 1405
rect 5974 1337 6052 1371
rect 6086 1337 6092 1371
rect 5974 1332 6092 1337
rect 5974 1298 5980 1332
rect 6014 1298 6092 1332
rect 5974 1264 6052 1298
rect 6086 1264 6092 1298
rect 5974 1259 6092 1264
rect 5974 1225 5980 1259
rect 6014 1225 6092 1259
rect 5974 1191 6052 1225
rect 6086 1191 6092 1225
rect 5974 1186 6092 1191
rect 5974 1152 5980 1186
rect 6014 1152 6092 1186
rect 5974 1118 6052 1152
rect 6086 1118 6092 1152
rect 5974 1113 6092 1118
rect 5974 1079 5980 1113
rect 6014 1079 6092 1113
rect 5974 1045 6052 1079
rect 6086 1045 6092 1079
rect 5974 1040 6092 1045
rect 5974 1006 5980 1040
rect 6014 1006 6092 1040
rect 5974 972 6052 1006
rect 6086 972 6092 1006
rect 5974 967 6092 972
rect 5974 933 5980 967
rect 6014 933 6092 967
rect 5974 899 6052 933
rect 6086 899 6092 933
rect 5974 894 6092 899
rect 5974 860 5980 894
rect 6014 860 6092 894
rect 5974 826 6052 860
rect 6086 826 6092 860
rect 5974 821 6092 826
rect 5974 787 5980 821
rect 6014 787 6092 821
rect 5974 753 6052 787
rect 6086 753 6092 787
rect 5974 748 6092 753
rect 5974 714 5980 748
rect 6014 714 6092 748
rect 5974 680 6052 714
rect 6086 680 6092 714
rect 5974 675 6092 680
rect 5974 641 5980 675
rect 6014 641 6092 675
tri 638 576 663 601 sw
tri 5419 576 5444 601 se
rect 5444 576 5522 609
rect 560 575 5522 576
rect 5556 604 5706 609
rect 5974 607 6052 641
rect 6086 607 6092 641
rect 5556 602 5698 604
tri 5698 602 5700 604 nw
rect 5974 602 6092 607
rect 5556 575 5664 602
rect 560 574 5664 575
tri 404 570 408 574 ne
rect 408 570 5664 574
tri 408 536 442 570 ne
rect 442 536 598 570
rect 632 536 671 570
rect 705 536 744 570
rect 778 536 817 570
rect 851 536 890 570
rect 924 536 963 570
rect 997 536 1036 570
rect 1070 536 1109 570
rect 1143 536 1182 570
rect 1216 536 1255 570
rect 1289 536 1328 570
rect 1362 536 1401 570
rect 1435 536 1474 570
rect 1508 536 1547 570
rect 1581 536 1620 570
rect 1654 536 1693 570
rect 1727 536 1766 570
rect 1800 536 1839 570
rect 1873 536 1912 570
rect 1946 536 1985 570
rect 2019 536 2058 570
rect 2092 536 2131 570
rect 2165 536 2204 570
rect 2238 536 2277 570
rect 2311 536 2350 570
rect 2384 536 2423 570
rect 2457 536 2496 570
rect 2530 536 2569 570
rect 2603 536 2642 570
tri 442 498 480 536 ne
rect 480 498 2642 536
tri 480 464 514 498 ne
rect 514 464 564 498
rect 598 464 637 498
rect 671 464 710 498
rect 744 464 783 498
rect 817 464 856 498
rect 890 464 929 498
rect 963 464 1002 498
rect 1036 464 1075 498
rect 1109 464 1148 498
rect 1182 464 1221 498
rect 1255 464 1294 498
rect 1328 464 1367 498
rect 1401 464 1440 498
rect 1474 464 1513 498
rect 1547 464 1586 498
rect 1620 464 1659 498
rect 1693 464 1732 498
rect 1766 464 1805 498
rect 1839 464 1878 498
rect 1912 464 1951 498
rect 1985 464 2024 498
rect 2058 464 2097 498
rect 2131 464 2170 498
rect 2204 464 2243 498
rect 2277 464 2316 498
rect 2350 464 2388 498
rect 2422 464 2460 498
rect 2494 464 2532 498
rect 2566 464 2604 498
rect 2638 464 2642 498
rect 5446 536 5450 570
rect 5484 568 5664 570
tri 5664 568 5698 602 nw
rect 5974 568 5980 602
rect 6014 568 6092 602
rect 5484 536 5630 568
rect 5446 502 5522 536
rect 5556 534 5630 536
tri 5630 534 5664 568 nw
rect 5974 534 6052 568
rect 6086 534 6092 568
rect 5556 529 5625 534
tri 5625 529 5630 534 nw
rect 5974 529 6092 534
rect 5556 502 5591 529
rect 5446 495 5591 502
tri 5591 495 5625 529 nw
rect 5974 495 5980 529
rect 6014 495 6092 529
rect 5446 464 5562 495
tri 5562 466 5591 495 nw
tri 514 461 517 464 ne
rect 517 461 5562 464
tri 517 458 520 461 ne
rect 520 458 5562 461
rect 5974 461 6052 495
rect 6086 461 6092 495
rect 5974 456 6092 461
rect 5974 422 5980 456
rect 6014 422 6092 456
rect 5974 388 6052 422
rect 6086 388 6092 422
rect 5974 383 6092 388
rect 5974 349 5980 383
rect 6014 349 6092 383
rect 5974 315 6052 349
rect 6086 315 6092 349
rect 5974 310 6092 315
rect 5974 276 5980 310
rect 6014 276 6092 310
rect 5974 242 6052 276
rect 6086 242 6092 276
rect 5974 237 6092 242
rect 108 203 144 223
tri 144 203 164 223 sw
rect 5974 203 5980 237
rect 6014 203 6092 237
rect 108 170 164 203
tri 164 170 197 203 sw
tri 5949 170 5974 195 se
rect 5974 170 6052 203
rect 108 169 6052 170
rect 6086 169 6092 203
rect 108 164 6092 169
rect 108 130 174 164
rect 208 130 247 164
rect 281 130 320 164
rect 354 130 393 164
rect 427 130 466 164
rect 500 130 539 164
rect 573 130 612 164
rect 646 130 685 164
rect 719 130 758 164
rect 792 130 831 164
rect 865 130 904 164
rect 938 130 977 164
rect 1011 130 1050 164
rect 1084 130 1123 164
rect 1157 130 1196 164
rect 1230 130 1269 164
rect 1303 130 1342 164
rect 1376 130 1415 164
rect 1449 130 1488 164
rect 1522 130 1561 164
rect 1595 130 1634 164
rect 1668 130 1707 164
rect 1741 130 1780 164
rect 1814 130 1853 164
rect 1887 130 1926 164
rect 1960 130 1999 164
rect 2033 130 2072 164
rect 2106 130 2145 164
rect 2179 130 2218 164
rect 2252 130 2291 164
rect 2325 130 2364 164
rect 2398 130 2437 164
rect 2471 130 2510 164
rect 2544 130 2583 164
rect 2617 130 2656 164
rect 2690 130 2729 164
rect 2763 130 2802 164
rect 2836 130 2875 164
rect 2909 130 2948 164
rect 2982 130 3021 164
rect 3055 130 3094 164
rect 3128 130 3167 164
rect 3201 130 3240 164
rect 3274 130 3313 164
rect 3347 130 3386 164
rect 3420 130 3459 164
rect 3493 130 3532 164
rect 108 92 3532 130
rect 108 58 174 92
rect 208 58 247 92
rect 281 58 320 92
rect 354 58 393 92
rect 427 58 466 92
rect 500 58 539 92
rect 573 58 612 92
rect 646 58 685 92
rect 719 58 758 92
rect 792 58 830 92
rect 864 58 902 92
rect 936 58 974 92
rect 1008 58 1046 92
rect 1080 58 1118 92
rect 1152 58 1190 92
rect 1224 58 1262 92
rect 1296 58 1334 92
rect 1368 58 1406 92
rect 1440 58 1478 92
rect 1512 58 1550 92
rect 1584 58 1622 92
rect 1656 58 1694 92
rect 1728 58 1766 92
rect 1800 58 1838 92
rect 1872 58 1910 92
rect 1944 58 1982 92
rect 2016 58 2054 92
rect 2088 58 2126 92
rect 2160 58 2198 92
rect 2232 58 2270 92
rect 2304 58 2342 92
rect 2376 58 2414 92
rect 2448 58 2486 92
rect 2520 58 2558 92
rect 2592 58 2630 92
rect 2664 58 2702 92
rect 2736 58 2774 92
rect 2808 58 2846 92
rect 2880 58 2918 92
rect 2952 58 2990 92
rect 3024 58 3062 92
rect 3096 58 3134 92
rect 3168 58 3206 92
rect 3240 58 3278 92
rect 3312 58 3350 92
rect 3384 58 3422 92
rect 3456 58 3494 92
rect 3528 58 3532 92
rect 5976 130 5980 164
rect 6014 130 6092 164
rect 5976 96 6052 130
rect 6086 96 6092 130
rect 5976 58 6092 96
rect 108 52 6092 58
use pfet_CDNS_524688791851487  pfet_CDNS_524688791851487_0
timestamp 1707688321
transform 1 0 687 0 -1 3724
box -266 -66 894 3066
use pfet_CDNS_524688791851490  pfet_CDNS_524688791851490_0
timestamp 1707688321
transform 1 0 1515 0 -1 3724
box -326 -66 894 3066
use pfet_CDNS_524688791851490  pfet_CDNS_524688791851490_1
timestamp 1707688321
transform 1 0 3999 0 -1 3724
box -326 -66 894 3066
use pfet_CDNS_524688791851490  pfet_CDNS_524688791851490_2
timestamp 1707688321
transform 1 0 3171 0 -1 3724
box -326 -66 894 3066
use pfet_CDNS_524688791851490  pfet_CDNS_524688791851490_3
timestamp 1707688321
transform 1 0 2343 0 -1 3724
box -326 -66 894 3066
use pfet_CDNS_524688791851491  pfet_CDNS_524688791851491_0
timestamp 1707688321
transform 1 0 4827 0 -1 3724
box -326 -66 834 3066
<< labels >>
flabel comment s 2901 3020 2901 3020 0 FreeSans 5000 0 0 0 vpb_drvr
flabel metal1 s 4327 2045 5273 2218 0 FreeSans 800 0 0 0 vcc_io
port 1 nsew
flabel metal1 s 2965 631 3110 681 0 FreeSans 400 0 0 0 pswg_h
port 2 nsew
flabel metal1 s 514 2523 1451 2689 0 FreeSans 800 0 0 0 vpb_drvr
port 3 nsew
flabel metal1 s 514 2258 1451 2424 0 FreeSans 800 0 0 0 vpb_drvr
port 3 nsew
flabel metal1 s 514 2789 1451 2955 0 FreeSans 800 0 0 0 vpb_drvr
port 3 nsew
flabel metal1 s 514 3050 1451 3216 0 FreeSans 800 0 0 0 vpb_drvr
port 3 nsew
flabel metal1 s 514 3311 1451 3477 0 FreeSans 800 0 0 0 vpb_drvr
port 3 nsew
flabel metal1 s 514 3577 1451 3743 0 FreeSans 800 0 0 0 vpb_drvr
port 3 nsew
flabel metal1 s 4327 725 5273 898 0 FreeSans 800 0 0 0 vcc_io
port 1 nsew
flabel metal1 s 4327 989 5273 1162 0 FreeSans 800 0 0 0 vcc_io
port 1 nsew
flabel metal1 s 4327 1254 5273 1427 0 FreeSans 800 0 0 0 vcc_io
port 1 nsew
flabel metal1 s 4327 1520 5273 1693 0 FreeSans 800 0 0 0 vcc_io
port 1 nsew
flabel metal1 s 4327 1781 5273 1954 0 FreeSans 800 0 0 0 vcc_io
port 1 nsew
<< properties >>
string GDS_END 89691490
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 89393544
string path 10.500 105.900 142.075 105.900 
<< end >>
