magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -68 -26 3683 92
<< ndiff >>
rect -42 50 0 66
rect -42 16 -34 50
rect -42 0 0 16
rect 3615 50 3657 66
rect 3649 16 3657 50
rect 3615 0 3657 16
<< ndiffc >>
rect -34 16 0 50
rect 3615 16 3649 50
<< ndiffres >>
rect 0 0 3615 66
<< locali >>
rect -34 50 0 66
rect -34 0 0 16
rect 3615 50 3649 66
rect 3615 0 3649 16
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_0
timestamp 1707688321
transform -1 0 8 0 1 4
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_1
timestamp 1707688321
transform 1 0 3607 0 1 4
box 0 0 1 1
<< properties >>
string GDS_END 78443586
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 78443084
<< end >>
