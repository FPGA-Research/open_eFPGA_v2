magic
tech sky130B
timestamp 1707688321
<< metal1 >>
rect 0 0 3 58
rect 893 0 896 58
<< via1 >>
rect 3 0 893 58
<< metal2 >>
rect 0 0 3 58
rect 893 0 896 58
<< properties >>
string GDS_END 91727104
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 91723388
<< end >>
