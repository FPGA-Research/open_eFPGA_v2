magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< poly >>
rect 85 376 219 392
rect 85 342 101 376
rect 135 342 169 376
rect 203 342 219 376
rect 85 326 219 342
rect -58 268 76 284
rect -58 234 -42 268
rect -8 234 26 268
rect 60 234 76 268
rect -58 218 76 234
<< polycont >>
rect 101 342 135 376
rect 169 342 203 376
rect -42 234 -8 268
rect 26 234 60 268
<< locali >>
rect 74 556 108 594
rect 230 472 264 510
rect 135 342 143 376
rect 203 342 219 376
rect -58 234 -42 268
rect -8 234 26 268
rect 64 234 76 268
rect 53 112 87 150
rect -105 24 -67 58
<< viali >>
rect 74 594 108 628
rect 74 522 108 556
rect 230 510 264 544
rect 230 438 264 472
rect 71 342 101 376
rect 101 342 105 376
rect 143 342 169 376
rect 169 342 177 376
rect -42 234 -8 268
rect 30 234 60 268
rect 60 234 64 268
rect 53 150 87 184
rect 53 78 87 112
rect -139 24 -105 58
rect -67 24 -33 58
<< metal1 >>
rect 31 628 114 690
rect 31 594 74 628
rect 108 594 114 628
rect 31 590 114 594
tri 34 556 68 590 ne
rect 68 556 114 590
rect 68 522 74 556
rect 108 522 114 556
rect 68 510 114 522
rect 221 548 273 556
rect 221 484 273 496
rect 221 426 273 432
rect -54 376 189 382
rect -54 342 71 376
rect 105 342 143 376
rect 177 342 189 376
rect -54 270 189 342
rect -54 268 76 270
rect -54 234 -42 268
rect -8 234 30 268
rect 64 234 76 268
rect -54 228 76 234
rect 44 190 96 196
rect 44 126 96 138
rect 44 66 96 74
rect -244 58 -21 64
rect -244 24 -139 58
rect -105 24 -67 58
rect -33 24 -21 58
rect -244 0 -21 24
<< via1 >>
rect 221 544 273 548
rect 221 510 230 544
rect 230 510 264 544
rect 264 510 273 544
rect 221 496 273 510
rect 221 472 273 484
rect 221 438 230 472
rect 230 438 264 472
rect 264 438 273 472
rect 221 432 273 438
rect 44 184 96 190
rect 44 150 53 184
rect 53 150 87 184
rect 87 150 96 184
rect 44 138 96 150
rect 44 112 96 126
rect 44 78 53 112
rect 53 78 87 112
rect 87 78 96 112
rect 44 74 96 78
<< metal2 >>
rect 221 548 273 554
rect 221 484 273 496
tri 147 299 221 373 se
rect 221 351 273 432
tri 221 299 273 351 nw
tri 73 225 147 299 se
tri 147 225 221 299 nw
tri 44 196 73 225 se
rect 73 196 118 225
tri 118 196 147 225 nw
rect 44 190 96 196
tri 96 174 118 196 nw
rect 44 126 96 138
rect 44 68 96 74
use nfet_CDNS_52468879185814  nfet_CDNS_52468879185814_0
timestamp 1707688321
transform 1 0 -58 0 1 36
box -82 -32 182 182
use pfet_CDNS_52468879185725  pfet_CDNS_52468879185725_0
timestamp 1707688321
transform 1 0 119 0 -1 624
box -119 -66 219 266
<< properties >>
string GDS_END 25735924
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 25732910
string path 6.175 10.650 6.175 13.850 
<< end >>
