magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< metal1 >>
rect 62637 78584 62643 78636
rect 62695 78624 62701 78636
rect 62851 78624 62857 78636
rect 62695 78596 62857 78624
rect 62695 78584 62701 78596
rect 62851 78584 62857 78596
rect 62909 78584 62915 78636
rect 61683 78482 61689 78534
rect 61741 78522 61747 78534
rect 62513 78522 62519 78534
rect 61741 78494 62519 78522
rect 61741 78482 61747 78494
rect 62513 78482 62519 78494
rect 62571 78482 62577 78534
rect 62761 78482 62767 78534
rect 62819 78522 62825 78534
rect 64019 78522 64025 78534
rect 62819 78494 64025 78522
rect 62819 78482 62825 78494
rect 64019 78482 64025 78494
rect 64077 78482 64083 78534
rect 62761 77683 62767 77735
rect 62819 77683 62825 77735
rect 62637 76193 62643 76245
rect 62695 76193 62701 76245
rect 62513 74855 62519 74907
rect 62571 74855 62577 74907
<< via1 >>
rect 62643 78584 62695 78636
rect 62857 78584 62909 78636
rect 61689 78482 61741 78534
rect 62519 78482 62571 78534
rect 62767 78482 62819 78534
rect 64025 78482 64077 78534
rect 62767 77683 62819 77735
rect 62643 76193 62695 76245
rect 62519 74855 62571 74907
<< metal2 >>
rect 61701 78540 61729 79883
rect 62869 78642 62897 79883
rect 62643 78636 62695 78642
rect 62643 78578 62695 78584
rect 62857 78636 62909 78642
rect 62857 78578 62909 78584
rect 61689 78534 61741 78540
rect 61689 78476 61741 78482
rect 62519 78534 62571 78540
rect 62519 78476 62571 78482
rect 62531 74913 62559 78476
rect 62655 76251 62683 78578
rect 64037 78540 64065 79883
rect 62767 78534 62819 78540
rect 62767 78476 62819 78482
rect 64025 78534 64077 78540
rect 64025 78476 64077 78482
rect 62779 77741 62807 78476
rect 62767 77735 62819 77741
rect 62767 77677 62819 77683
rect 62643 76245 62695 76251
rect 62643 76187 62695 76193
rect 62519 74907 62571 74913
rect 62519 74849 62571 74855
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_0
timestamp 1707688321
transform 1 0 62851 0 1 78578
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_1
timestamp 1707688321
transform 1 0 62637 0 1 76187
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_2
timestamp 1707688321
transform 1 0 62637 0 1 78578
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_3
timestamp 1707688321
transform 1 0 64019 0 1 78476
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_4
timestamp 1707688321
transform 1 0 62761 0 1 77677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_5
timestamp 1707688321
transform 1 0 62761 0 1 78476
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_6
timestamp 1707688321
transform 1 0 61683 0 1 78476
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_7
timestamp 1707688321
transform 1 0 62513 0 1 74849
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_8
timestamp 1707688321
transform 1 0 62513 0 1 78476
box 0 0 1 1
<< properties >>
string FIXED_BBOX 61683 74849 64083 79883
string GDS_END 7023352
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_8x1024_8.gds
string GDS_START 7021786
<< end >>
