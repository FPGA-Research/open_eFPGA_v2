magic
tech sky130B
timestamp 1707688321
<< viali >>
rect 0 0 125 1889
<< metal1 >>
rect -6 1889 131 1892
rect -6 0 0 1889
rect 125 0 131 1889
rect -6 -3 131 0
<< properties >>
string GDS_END 98210024
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 98196324
<< end >>
