magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -26 -26 226 1026
<< ndiff >>
rect 0 930 60 1000
rect 0 896 11 930
rect 45 896 60 930
rect 0 862 60 896
rect 0 828 11 862
rect 45 828 60 862
rect 0 794 60 828
rect 0 760 11 794
rect 45 760 60 794
rect 0 726 60 760
rect 0 692 11 726
rect 45 692 60 726
rect 0 658 60 692
rect 0 624 11 658
rect 45 624 60 658
rect 0 590 60 624
rect 0 556 11 590
rect 45 556 60 590
rect 0 522 60 556
rect 0 488 11 522
rect 45 488 60 522
rect 0 454 60 488
rect 0 420 11 454
rect 45 420 60 454
rect 0 386 60 420
rect 0 352 11 386
rect 45 352 60 386
rect 0 318 60 352
rect 0 284 11 318
rect 45 284 60 318
rect 0 250 60 284
rect 0 216 11 250
rect 45 216 60 250
rect 0 182 60 216
rect 0 148 11 182
rect 45 148 60 182
rect 0 114 60 148
rect 0 80 11 114
rect 45 80 60 114
rect 0 46 60 80
rect 0 12 11 46
rect 45 12 60 46
rect 0 0 60 12
<< ndiffc >>
rect 11 896 45 930
rect 11 828 45 862
rect 11 760 45 794
rect 11 692 45 726
rect 11 624 45 658
rect 11 556 45 590
rect 11 488 45 522
rect 11 420 45 454
rect 11 352 45 386
rect 11 284 45 318
rect 11 216 45 250
rect 11 148 45 182
rect 11 80 45 114
rect 11 12 45 46
<< psubdiff >>
rect 60 942 200 1000
rect 60 908 79 942
rect 113 908 200 942
rect 60 874 200 908
rect 60 840 79 874
rect 113 840 200 874
rect 60 806 200 840
rect 60 772 79 806
rect 113 772 200 806
rect 60 738 200 772
rect 60 704 79 738
rect 113 704 200 738
rect 60 670 200 704
rect 60 636 79 670
rect 113 636 200 670
rect 60 602 200 636
rect 60 568 79 602
rect 113 568 200 602
rect 60 534 200 568
rect 60 500 79 534
rect 113 500 200 534
rect 60 466 200 500
rect 60 432 79 466
rect 113 432 200 466
rect 60 398 200 432
rect 60 364 79 398
rect 113 364 200 398
rect 60 330 200 364
rect 60 296 79 330
rect 113 296 200 330
rect 60 262 200 296
rect 60 228 79 262
rect 113 228 200 262
rect 60 194 200 228
rect 60 160 79 194
rect 113 160 200 194
rect 60 126 200 160
rect 60 92 79 126
rect 113 92 200 126
rect 60 58 200 92
rect 60 24 79 58
rect 113 24 200 58
rect 60 0 200 24
<< psubdiffcont >>
rect 79 908 113 942
rect 79 840 113 874
rect 79 772 113 806
rect 79 704 113 738
rect 79 636 113 670
rect 79 568 113 602
rect 79 500 113 534
rect 79 432 113 466
rect 79 364 113 398
rect 79 296 113 330
rect 79 228 113 262
rect 79 160 113 194
rect 79 92 113 126
rect 79 24 113 58
<< locali >>
rect 11 942 113 958
rect 11 930 79 942
rect 45 908 79 930
rect 45 896 113 908
rect 11 874 113 896
rect 11 862 79 874
rect 45 840 79 862
rect 45 828 113 840
rect 11 806 113 828
rect 11 794 79 806
rect 45 772 79 794
rect 45 760 113 772
rect 11 738 113 760
rect 11 726 79 738
rect 45 704 79 726
rect 45 692 113 704
rect 11 670 113 692
rect 11 658 79 670
rect 45 636 79 658
rect 45 624 113 636
rect 11 602 113 624
rect 11 590 79 602
rect 45 568 79 590
rect 45 556 113 568
rect 11 534 113 556
rect 11 522 79 534
rect 45 500 79 522
rect 45 488 113 500
rect 11 466 113 488
rect 11 454 79 466
rect 45 432 79 454
rect 45 420 113 432
rect 11 398 113 420
rect 11 386 79 398
rect 45 364 79 386
rect 45 352 113 364
rect 11 330 113 352
rect 11 318 79 330
rect 45 296 79 318
rect 45 284 113 296
rect 11 262 113 284
rect 11 250 79 262
rect 45 228 79 250
rect 45 216 113 228
rect 11 194 113 216
rect 11 182 79 194
rect 45 160 79 182
rect 45 148 113 160
rect 11 126 113 148
rect 11 114 79 126
rect 45 92 79 114
rect 45 80 113 92
rect 11 58 113 80
rect 11 46 79 58
rect 45 24 79 46
rect 45 12 113 24
rect 11 -4 113 12
<< properties >>
string GDS_END 13673102
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 13670922
<< end >>
