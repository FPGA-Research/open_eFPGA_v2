magic
tech sky130A
timestamp 1707688321
<< locali >>
rect 17 1344 36 1361
rect 53 1344 72 1361
rect 0 1313 89 1344
rect 17 1296 36 1313
rect 53 1296 72 1313
rect 0 1265 89 1296
rect 17 1248 36 1265
rect 53 1248 72 1265
rect 0 1217 89 1248
rect 17 1200 36 1217
rect 53 1200 72 1217
rect 0 1169 89 1200
rect 17 1152 36 1169
rect 53 1152 72 1169
rect 0 1121 89 1152
rect 17 1104 36 1121
rect 53 1104 72 1121
rect 0 1073 89 1104
rect 17 1056 36 1073
rect 53 1056 72 1073
rect 0 1025 89 1056
rect 17 1008 36 1025
rect 53 1008 72 1025
rect 0 977 89 1008
rect 17 960 36 977
rect 53 960 72 977
rect 0 929 89 960
rect 17 912 36 929
rect 53 912 72 929
rect 0 881 89 912
rect 17 864 36 881
rect 53 864 72 881
rect 0 833 89 864
rect 17 816 36 833
rect 53 816 72 833
rect 0 785 89 816
rect 17 768 36 785
rect 53 768 72 785
rect 0 737 89 768
rect 17 720 36 737
rect 53 720 72 737
rect 0 689 89 720
rect 17 672 36 689
rect 53 672 72 689
rect 0 641 89 672
rect 17 624 36 641
rect 53 624 72 641
rect 0 593 89 624
rect 17 576 36 593
rect 53 576 72 593
rect 0 545 89 576
rect 17 528 36 545
rect 53 528 72 545
rect 0 497 89 528
rect 17 480 36 497
rect 53 480 72 497
rect 0 449 89 480
rect 17 432 36 449
rect 53 432 72 449
rect 0 401 89 432
rect 17 384 36 401
rect 53 384 72 401
rect 0 353 89 384
rect 17 336 36 353
rect 53 336 72 353
rect 0 305 89 336
rect 17 288 36 305
rect 53 288 72 305
rect 0 257 89 288
rect 17 240 36 257
rect 53 240 72 257
rect 0 209 89 240
rect 17 192 36 209
rect 53 192 72 209
rect 0 161 89 192
rect 17 144 36 161
rect 53 144 72 161
rect 0 113 89 144
rect 17 96 36 113
rect 53 96 72 113
rect 0 65 89 96
rect 17 48 36 65
rect 53 48 72 65
rect 0 17 89 48
rect 17 0 36 17
rect 53 0 72 17
<< viali >>
rect 0 1344 17 1361
rect 36 1344 53 1361
rect 72 1344 89 1361
rect 0 1296 17 1313
rect 36 1296 53 1313
rect 72 1296 89 1313
rect 0 1248 17 1265
rect 36 1248 53 1265
rect 72 1248 89 1265
rect 0 1200 17 1217
rect 36 1200 53 1217
rect 72 1200 89 1217
rect 0 1152 17 1169
rect 36 1152 53 1169
rect 72 1152 89 1169
rect 0 1104 17 1121
rect 36 1104 53 1121
rect 72 1104 89 1121
rect 0 1056 17 1073
rect 36 1056 53 1073
rect 72 1056 89 1073
rect 0 1008 17 1025
rect 36 1008 53 1025
rect 72 1008 89 1025
rect 0 960 17 977
rect 36 960 53 977
rect 72 960 89 977
rect 0 912 17 929
rect 36 912 53 929
rect 72 912 89 929
rect 0 864 17 881
rect 36 864 53 881
rect 72 864 89 881
rect 0 816 17 833
rect 36 816 53 833
rect 72 816 89 833
rect 0 768 17 785
rect 36 768 53 785
rect 72 768 89 785
rect 0 720 17 737
rect 36 720 53 737
rect 72 720 89 737
rect 0 672 17 689
rect 36 672 53 689
rect 72 672 89 689
rect 0 624 17 641
rect 36 624 53 641
rect 72 624 89 641
rect 0 576 17 593
rect 36 576 53 593
rect 72 576 89 593
rect 0 528 17 545
rect 36 528 53 545
rect 72 528 89 545
rect 0 480 17 497
rect 36 480 53 497
rect 72 480 89 497
rect 0 432 17 449
rect 36 432 53 449
rect 72 432 89 449
rect 0 384 17 401
rect 36 384 53 401
rect 72 384 89 401
rect 0 336 17 353
rect 36 336 53 353
rect 72 336 89 353
rect 0 288 17 305
rect 36 288 53 305
rect 72 288 89 305
rect 0 240 17 257
rect 36 240 53 257
rect 72 240 89 257
rect 0 192 17 209
rect 36 192 53 209
rect 72 192 89 209
rect 0 144 17 161
rect 36 144 53 161
rect 72 144 89 161
rect 0 96 17 113
rect 36 96 53 113
rect 72 96 89 113
rect 0 48 17 65
rect 36 48 53 65
rect 72 48 89 65
rect 0 0 17 17
rect 36 0 53 17
rect 72 0 89 17
<< metal1 >>
rect -6 1361 95 1364
rect -6 1344 0 1361
rect 17 1344 36 1361
rect 53 1344 72 1361
rect 89 1344 95 1361
rect -6 1313 95 1344
rect -6 1296 0 1313
rect 17 1296 36 1313
rect 53 1296 72 1313
rect 89 1296 95 1313
rect -6 1265 95 1296
rect -6 1248 0 1265
rect 17 1248 36 1265
rect 53 1248 72 1265
rect 89 1248 95 1265
rect -6 1217 95 1248
rect -6 1200 0 1217
rect 17 1200 36 1217
rect 53 1200 72 1217
rect 89 1200 95 1217
rect -6 1169 95 1200
rect -6 1152 0 1169
rect 17 1152 36 1169
rect 53 1152 72 1169
rect 89 1152 95 1169
rect -6 1121 95 1152
rect -6 1104 0 1121
rect 17 1104 36 1121
rect 53 1104 72 1121
rect 89 1104 95 1121
rect -6 1073 95 1104
rect -6 1056 0 1073
rect 17 1056 36 1073
rect 53 1056 72 1073
rect 89 1056 95 1073
rect -6 1025 95 1056
rect -6 1008 0 1025
rect 17 1008 36 1025
rect 53 1008 72 1025
rect 89 1008 95 1025
rect -6 977 95 1008
rect -6 960 0 977
rect 17 960 36 977
rect 53 960 72 977
rect 89 960 95 977
rect -6 929 95 960
rect -6 912 0 929
rect 17 912 36 929
rect 53 912 72 929
rect 89 912 95 929
rect -6 881 95 912
rect -6 864 0 881
rect 17 864 36 881
rect 53 864 72 881
rect 89 864 95 881
rect -6 833 95 864
rect -6 816 0 833
rect 17 816 36 833
rect 53 816 72 833
rect 89 816 95 833
rect -6 785 95 816
rect -6 768 0 785
rect 17 768 36 785
rect 53 768 72 785
rect 89 768 95 785
rect -6 737 95 768
rect -6 720 0 737
rect 17 720 36 737
rect 53 720 72 737
rect 89 720 95 737
rect -6 689 95 720
rect -6 672 0 689
rect 17 672 36 689
rect 53 672 72 689
rect 89 672 95 689
rect -6 641 95 672
rect -6 624 0 641
rect 17 624 36 641
rect 53 624 72 641
rect 89 624 95 641
rect -6 593 95 624
rect -6 576 0 593
rect 17 576 36 593
rect 53 576 72 593
rect 89 576 95 593
rect -6 545 95 576
rect -6 528 0 545
rect 17 528 36 545
rect 53 528 72 545
rect 89 528 95 545
rect -6 497 95 528
rect -6 480 0 497
rect 17 480 36 497
rect 53 480 72 497
rect 89 480 95 497
rect -6 449 95 480
rect -6 432 0 449
rect 17 432 36 449
rect 53 432 72 449
rect 89 432 95 449
rect -6 401 95 432
rect -6 384 0 401
rect 17 384 36 401
rect 53 384 72 401
rect 89 384 95 401
rect -6 353 95 384
rect -6 336 0 353
rect 17 336 36 353
rect 53 336 72 353
rect 89 336 95 353
rect -6 305 95 336
rect -6 288 0 305
rect 17 288 36 305
rect 53 288 72 305
rect 89 288 95 305
rect -6 257 95 288
rect -6 240 0 257
rect 17 240 36 257
rect 53 240 72 257
rect 89 240 95 257
rect -6 209 95 240
rect -6 192 0 209
rect 17 192 36 209
rect 53 192 72 209
rect 89 192 95 209
rect -6 161 95 192
rect -6 144 0 161
rect 17 144 36 161
rect 53 144 72 161
rect 89 144 95 161
rect -6 113 95 144
rect -6 96 0 113
rect 17 96 36 113
rect 53 96 72 113
rect 89 96 95 113
rect -6 65 95 96
rect -6 48 0 65
rect 17 48 36 65
rect 53 48 72 65
rect 89 48 95 65
rect -6 17 95 48
rect -6 0 0 17
rect 17 0 36 17
rect 53 0 72 17
rect 89 0 95 17
rect -6 -3 95 0
<< properties >>
string GDS_END 42957968
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 42952268
<< end >>
