magic
tech sky130B
timestamp 1707688321
<< viali >>
rect 0 0 53 5417
<< metal1 >>
rect -6 5417 59 5420
rect -6 0 0 5417
rect 53 0 59 5417
rect -6 -3 59 0
<< properties >>
string GDS_END 92064410
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 92044950
<< end >>
