magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -89 -36 545 1036
<< pmoslvt >>
rect 0 0 200 1000
rect 256 0 456 1000
<< pdiff >>
rect -50 0 0 1000
rect 456 0 506 1000
<< poly >>
rect 0 1000 200 1026
rect 0 -26 200 0
rect 256 1000 456 1026
rect 256 -26 456 0
<< metal1 >>
rect -51 -16 -5 978
rect 205 -16 251 978
rect 461 -16 507 978
use DFM1sd2_CDNS_52468879185176  DFM1sd2_CDNS_52468879185176_0
timestamp 1707688321
transform 1 0 200 0 1 0
box -36 -36 92 1036
use DFM1sd_CDNS_52468879185574  DFM1sd_CDNS_52468879185574_0
timestamp 1707688321
transform -1 0 0 0 1 0
box -36 -36 89 1036
use DFM1sd_CDNS_52468879185574  DFM1sd_CDNS_52468879185574_1
timestamp 1707688321
transform 1 0 456 0 1 0
box -36 -36 89 1036
<< labels >>
flabel comment s -28 481 -28 481 0 FreeSans 300 0 0 0 S
flabel comment s 228 481 228 481 0 FreeSans 300 0 0 0 D
flabel comment s 484 481 484 481 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 86597460
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86596012
<< end >>
