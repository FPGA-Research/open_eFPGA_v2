magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< metal2 >>
rect 0 665 376 674
rect 56 609 80 665
rect 136 609 160 665
rect 216 609 240 665
rect 296 609 320 665
rect 0 465 376 609
rect 56 409 80 465
rect 136 409 160 465
rect 216 409 240 465
rect 296 409 320 465
rect 0 265 376 409
rect 56 209 80 265
rect 136 209 160 265
rect 216 209 240 265
rect 296 209 320 265
rect 0 65 376 209
rect 56 9 80 65
rect 136 9 160 65
rect 216 9 240 65
rect 296 9 320 65
rect 0 0 376 9
<< via2 >>
rect 0 609 56 665
rect 80 609 136 665
rect 160 609 216 665
rect 240 609 296 665
rect 320 609 376 665
rect 0 409 56 465
rect 80 409 136 465
rect 160 409 216 465
rect 240 409 296 465
rect 320 409 376 465
rect 0 209 56 265
rect 80 209 136 265
rect 160 209 216 265
rect 240 209 296 265
rect 320 209 376 265
rect 0 9 56 65
rect 80 9 136 65
rect 160 9 216 65
rect 240 9 296 65
rect 320 9 376 65
<< metal3 >>
rect -5 665 381 670
rect -5 609 0 665
rect 56 609 80 665
rect 136 609 160 665
rect 216 609 240 665
rect 296 609 320 665
rect 376 609 381 665
rect -5 465 381 609
rect -5 409 0 465
rect 56 409 80 465
rect 136 409 160 465
rect 216 409 240 465
rect 296 409 320 465
rect 376 409 381 465
rect -5 265 381 409
rect -5 209 0 265
rect 56 209 80 265
rect 136 209 160 265
rect 216 209 240 265
rect 296 209 320 265
rect 376 209 381 265
rect -5 65 381 209
rect -5 9 0 65
rect 56 9 80 65
rect 136 9 160 65
rect 216 9 240 65
rect 296 9 320 65
rect 376 9 381 65
rect -5 4 381 9
<< properties >>
string GDS_END 78399930
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 78398518
<< end >>
