magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< locali >>
rect 77 3096 111 3112
rect 1459 3096 1493 3112
rect 111 3062 1459 3096
rect 1493 3062 1942 3096
rect 77 3046 111 3062
rect 1459 3046 1493 3062
rect 3259 3023 3836 3057
rect 157 2984 191 3000
rect 1539 2984 1573 3000
rect 191 2950 1539 2984
rect 1573 2950 1832 2984
rect 157 2934 191 2950
rect 1539 2934 1573 2950
rect 237 2894 271 2910
rect 1619 2894 1653 2910
rect 271 2860 1619 2894
rect 1653 2860 1942 2894
rect 237 2844 271 2860
rect 1619 2844 1653 2860
rect 1603 2636 1619 2670
rect 1653 2636 1942 2670
rect 1523 2546 1539 2580
rect 1573 2546 1832 2580
rect 3259 2473 3836 2507
rect 1203 2434 1219 2468
rect 1253 2434 1942 2468
rect 1443 2272 1459 2306
rect 1493 2272 1942 2306
rect 3259 2233 3836 2267
rect 1283 2160 1299 2194
rect 1333 2160 1832 2194
rect 1603 2070 1619 2104
rect 1653 2070 1942 2104
rect 1603 1846 1619 1880
rect 1653 1846 1942 1880
rect 1283 1756 1299 1790
rect 1333 1756 1832 1790
rect 3259 1683 3836 1717
rect 1203 1644 1219 1678
rect 1253 1644 1942 1678
rect 1443 1482 1459 1516
rect 1493 1482 1942 1516
rect 3259 1443 3836 1477
rect 1523 1370 1539 1404
rect 1573 1370 1832 1404
rect 1363 1280 1379 1314
rect 1413 1280 1942 1314
rect 1363 1056 1379 1090
rect 1413 1056 1942 1090
rect 221 943 237 977
rect 271 943 494 977
rect 1523 966 1539 1000
rect 1573 966 1832 1000
rect 1125 927 1159 943
rect 3259 893 3836 927
rect 1125 877 1159 893
rect 1203 854 1219 888
rect 1253 854 1942 888
rect 1125 687 1159 703
rect 1443 692 1459 726
rect 1493 692 1942 726
rect 3259 653 3836 687
rect 1125 637 1159 653
rect 141 603 157 637
rect 191 603 494 637
rect 1283 580 1299 614
rect 1333 580 1832 614
rect 1363 490 1379 524
rect 1413 490 1942 524
rect 1363 266 1379 300
rect 1413 266 1942 300
rect 61 153 77 187
rect 111 153 494 187
rect 1283 176 1299 210
rect 1333 176 1832 210
rect 1125 137 1159 153
rect 3259 103 3836 137
rect 1125 87 1159 103
rect 1203 64 1219 98
rect 1253 64 1942 98
<< viali >>
rect 77 3062 111 3096
rect 1459 3062 1493 3096
rect 157 2950 191 2984
rect 1539 2950 1573 2984
rect 237 2860 271 2894
rect 1619 2860 1653 2894
rect 1619 2636 1653 2670
rect 1539 2546 1573 2580
rect 1219 2434 1253 2468
rect 1459 2272 1493 2306
rect 1299 2160 1333 2194
rect 1619 2070 1653 2104
rect 1619 1846 1653 1880
rect 1299 1756 1333 1790
rect 1219 1644 1253 1678
rect 1459 1482 1493 1516
rect 1539 1370 1573 1404
rect 1379 1280 1413 1314
rect 1379 1056 1413 1090
rect 237 943 271 977
rect 1539 966 1573 1000
rect 1125 893 1159 927
rect 1219 854 1253 888
rect 1459 692 1493 726
rect 1125 653 1159 687
rect 157 603 191 637
rect 1299 580 1333 614
rect 1379 490 1413 524
rect 1379 266 1413 300
rect 77 153 111 187
rect 1299 176 1333 210
rect 1125 103 1159 137
rect 1219 64 1253 98
<< metal1 >>
rect 1453 3102 1499 3108
rect 65 3096 123 3102
rect 65 3062 77 3096
rect 111 3062 123 3096
rect 1447 3096 1505 3102
rect 65 3056 123 3062
rect 80 199 108 3056
rect 160 2990 188 3080
rect 145 2984 203 2990
rect 145 2950 157 2984
rect 191 2950 203 2984
rect 145 2944 203 2950
rect 160 649 188 2944
rect 240 2900 268 3080
rect 225 2894 283 2900
rect 225 2860 237 2894
rect 271 2860 283 2894
rect 225 2854 283 2860
rect 240 989 268 2854
rect 1222 2480 1250 3080
rect 1213 2468 1259 2480
rect 1213 2434 1219 2468
rect 1253 2434 1259 2468
rect 1213 2422 1259 2434
rect 1222 1690 1250 2422
rect 1302 2206 1330 3080
rect 1293 2194 1339 2206
rect 1293 2160 1299 2194
rect 1333 2160 1339 2194
rect 1293 2148 1339 2160
rect 1302 1802 1330 2148
rect 1293 1790 1339 1802
rect 1293 1756 1299 1790
rect 1333 1756 1339 1790
rect 1293 1744 1339 1756
rect 1213 1678 1259 1690
rect 1213 1644 1219 1678
rect 1253 1644 1259 1678
rect 1213 1632 1259 1644
rect 231 977 277 989
rect 231 943 237 977
rect 271 943 277 977
rect 231 931 277 943
rect 151 637 197 649
rect 151 603 157 637
rect 191 603 197 637
rect 151 591 197 603
rect 71 187 117 199
rect 71 153 77 187
rect 111 153 117 187
rect 71 141 117 153
rect 80 80 108 141
rect 160 80 188 591
rect 240 80 268 931
rect 584 421 612 1185
rect 980 421 1008 1185
rect 1110 884 1116 936
rect 1168 884 1174 936
rect 1222 900 1250 1632
rect 1213 888 1259 900
rect 1213 854 1219 888
rect 1253 854 1259 888
rect 1213 842 1259 854
rect 1110 644 1116 696
rect 1168 644 1174 696
rect 566 369 572 421
rect 624 369 630 421
rect 962 369 968 421
rect 1020 369 1026 421
rect 584 80 612 369
rect 980 80 1008 369
rect 1222 343 1250 842
rect 1302 738 1330 1744
rect 1382 1326 1410 3080
rect 1447 3062 1459 3096
rect 1493 3062 1505 3096
rect 1447 3056 1505 3062
rect 1453 3050 1499 3056
rect 1462 2318 1490 3050
rect 1542 2996 1570 3080
rect 1533 2990 1579 2996
rect 1527 2984 1585 2990
rect 1527 2950 1539 2984
rect 1573 2950 1585 2984
rect 1527 2944 1585 2950
rect 1533 2938 1579 2944
rect 1542 2592 1570 2938
rect 1622 2906 1650 3080
rect 1613 2900 1659 2906
rect 1607 2894 1665 2900
rect 1607 2860 1619 2894
rect 1653 2860 1665 2894
rect 1607 2854 1665 2860
rect 1613 2848 1659 2854
rect 1622 2682 1650 2848
rect 2030 2814 2076 3204
rect 2454 2814 2502 3146
rect 2886 2814 2934 3146
rect 2021 2762 2027 2814
rect 2079 2762 2085 2814
rect 2446 2762 2452 2814
rect 2504 2762 2510 2814
rect 2878 2762 2884 2814
rect 2936 2762 2942 2814
rect 3278 2791 3306 3160
rect 3674 2791 3702 3160
rect 1613 2670 1659 2682
rect 1613 2636 1619 2670
rect 1653 2636 1659 2670
rect 1613 2624 1659 2636
rect 1533 2580 1579 2592
rect 1533 2546 1539 2580
rect 1573 2546 1579 2580
rect 1533 2534 1579 2546
rect 1453 2306 1499 2318
rect 1453 2272 1459 2306
rect 1493 2272 1499 2306
rect 1453 2260 1499 2272
rect 1462 1528 1490 2260
rect 1453 1516 1499 1528
rect 1453 1482 1459 1516
rect 1493 1482 1499 1516
rect 1453 1470 1499 1482
rect 1373 1314 1419 1326
rect 1373 1280 1379 1314
rect 1413 1280 1419 1314
rect 1373 1268 1419 1280
rect 1382 1133 1410 1268
rect 1370 1127 1422 1133
rect 1370 1069 1379 1075
rect 1373 1056 1379 1069
rect 1413 1069 1422 1075
rect 1413 1056 1419 1069
rect 1373 1044 1419 1056
rect 1290 732 1342 738
rect 1290 674 1342 680
rect 1302 626 1330 674
rect 1293 614 1339 626
rect 1293 580 1299 614
rect 1333 580 1339 614
rect 1293 568 1339 580
rect 1210 337 1262 343
rect 1210 279 1262 285
rect 1110 94 1116 146
rect 1168 94 1174 146
rect 1222 110 1250 279
rect 1302 222 1330 568
rect 1382 536 1410 1044
rect 1462 738 1490 1470
rect 1542 1416 1570 2534
rect 1622 2116 1650 2624
rect 1613 2104 1659 2116
rect 1613 2070 1619 2104
rect 1653 2070 1659 2104
rect 1613 2058 1659 2070
rect 1622 1892 1650 2058
rect 2030 2024 2076 2762
rect 2454 2024 2502 2762
rect 2886 2024 2934 2762
rect 3260 2739 3266 2791
rect 3318 2739 3324 2791
rect 3656 2739 3662 2791
rect 3714 2739 3720 2791
rect 2021 1972 2027 2024
rect 2079 1972 2085 2024
rect 2446 1972 2452 2024
rect 2504 1972 2510 2024
rect 2878 1972 2884 2024
rect 2936 1972 2942 2024
rect 3278 2001 3306 2739
rect 3674 2001 3702 2739
rect 1613 1880 1659 1892
rect 1613 1846 1619 1880
rect 1653 1846 1659 1880
rect 1613 1834 1659 1846
rect 1533 1404 1579 1416
rect 1533 1370 1539 1404
rect 1573 1370 1579 1404
rect 1533 1358 1579 1370
rect 1542 1012 1570 1358
rect 1533 1000 1579 1012
rect 1533 966 1539 1000
rect 1573 966 1579 1000
rect 1533 954 1579 966
rect 1453 726 1499 738
rect 1453 692 1459 726
rect 1493 692 1499 726
rect 1453 680 1499 692
rect 1373 524 1419 536
rect 1373 490 1379 524
rect 1413 490 1419 524
rect 1373 478 1419 490
rect 1382 312 1410 478
rect 1373 300 1419 312
rect 1373 266 1379 300
rect 1413 266 1419 300
rect 1373 254 1419 266
rect 1293 210 1339 222
rect 1293 176 1299 210
rect 1333 176 1339 210
rect 1293 164 1339 176
rect 1213 98 1259 110
rect 1213 64 1219 98
rect 1253 64 1259 98
rect 1302 80 1330 164
rect 1382 80 1410 254
rect 1462 80 1490 680
rect 1542 80 1570 954
rect 1622 80 1650 1834
rect 2030 1234 2076 1972
rect 2454 1234 2502 1972
rect 2886 1234 2934 1972
rect 3260 1949 3266 2001
rect 3318 1949 3324 2001
rect 3656 1949 3662 2001
rect 3714 1949 3720 2001
rect 2021 1182 2027 1234
rect 2079 1182 2085 1234
rect 2446 1182 2452 1234
rect 2504 1182 2510 1234
rect 2878 1182 2884 1234
rect 2936 1182 2942 1234
rect 3278 1211 3306 1949
rect 3674 1211 3702 1949
rect 2030 444 2076 1182
rect 2454 444 2502 1182
rect 2886 444 2934 1182
rect 3260 1159 3266 1211
rect 3318 1159 3324 1211
rect 3656 1159 3662 1211
rect 3714 1159 3720 1211
rect 2021 392 2027 444
rect 2079 392 2085 444
rect 2446 392 2452 444
rect 2504 392 2510 444
rect 2878 392 2884 444
rect 2936 392 2942 444
rect 3278 421 3306 1159
rect 3674 421 3702 1159
rect 2030 80 2076 392
rect 2454 80 2502 392
rect 2886 80 2934 392
rect 3260 369 3266 421
rect 3318 369 3324 421
rect 3656 369 3662 421
rect 3714 369 3720 421
rect 3278 80 3306 369
rect 3674 80 3702 369
rect 1213 52 1259 64
<< via1 >>
rect 1116 927 1168 936
rect 1116 893 1125 927
rect 1125 893 1159 927
rect 1159 893 1168 927
rect 1116 884 1168 893
rect 1116 687 1168 696
rect 1116 653 1125 687
rect 1125 653 1159 687
rect 1159 653 1168 687
rect 1116 644 1168 653
rect 572 369 624 421
rect 968 369 1020 421
rect 2027 2762 2079 2814
rect 2452 2762 2504 2814
rect 2884 2762 2936 2814
rect 1370 1090 1422 1127
rect 1370 1075 1379 1090
rect 1379 1075 1413 1090
rect 1413 1075 1422 1090
rect 1290 680 1342 732
rect 1210 285 1262 337
rect 1116 137 1168 146
rect 1116 103 1125 137
rect 1125 103 1159 137
rect 1159 103 1168 137
rect 1116 94 1168 103
rect 3266 2739 3318 2791
rect 3662 2739 3714 2791
rect 2027 1972 2079 2024
rect 2452 1972 2504 2024
rect 2884 1972 2936 2024
rect 3266 1949 3318 2001
rect 3662 1949 3714 2001
rect 2027 1182 2079 1234
rect 2452 1182 2504 1234
rect 2884 1182 2936 1234
rect 3266 1159 3318 1211
rect 3662 1159 3714 1211
rect 2027 392 2079 444
rect 2452 392 2504 444
rect 2884 392 2936 444
rect 3266 369 3318 421
rect 3662 369 3714 421
<< metal2 >>
rect 2025 2816 2081 2825
rect 2025 2751 2081 2760
rect 2450 2816 2506 2825
rect 2450 2751 2506 2760
rect 2882 2816 2938 2825
rect 2882 2751 2938 2760
rect 3264 2793 3320 2802
rect 3264 2728 3320 2737
rect 3660 2793 3716 2802
rect 3660 2728 3716 2737
rect 2025 2026 2081 2035
rect 2025 1961 2081 1970
rect 2450 2026 2506 2035
rect 2450 1961 2506 1970
rect 2882 2026 2938 2035
rect 2882 1961 2938 1970
rect 3264 2003 3320 2012
rect 3264 1938 3320 1947
rect 3660 2003 3716 2012
rect 3660 1938 3716 1947
rect 2025 1236 2081 1245
rect 2025 1171 2081 1180
rect 2450 1236 2506 1245
rect 2450 1171 2506 1180
rect 2882 1236 2938 1245
rect 2882 1171 2938 1180
rect 3264 1213 3320 1222
rect 3264 1148 3320 1157
rect 3660 1213 3716 1222
rect 3660 1148 3716 1157
rect 1364 1115 1370 1127
rect 1128 1087 1370 1115
rect 1128 942 1156 1087
rect 1364 1075 1370 1087
rect 1422 1075 1428 1127
rect 1116 936 1168 942
rect 1116 878 1168 884
rect 1284 720 1290 732
rect 1128 702 1290 720
rect 1116 696 1290 702
rect 1168 692 1290 696
rect 1284 680 1290 692
rect 1342 680 1348 732
rect 1116 638 1168 644
rect 2025 446 2081 455
rect 570 423 626 432
rect 570 358 626 367
rect 966 423 1022 432
rect 2025 381 2081 390
rect 2450 446 2506 455
rect 2450 381 2506 390
rect 2882 446 2938 455
rect 2882 381 2938 390
rect 3264 423 3320 432
rect 966 358 1022 367
rect 3264 358 3320 367
rect 3660 423 3716 432
rect 3660 358 3716 367
rect 1204 325 1210 337
rect 1128 297 1210 325
rect 1128 152 1156 297
rect 1204 285 1210 297
rect 1262 285 1268 337
rect 1116 146 1168 152
rect 1116 88 1168 94
<< via2 >>
rect 2025 2814 2081 2816
rect 2025 2762 2027 2814
rect 2027 2762 2079 2814
rect 2079 2762 2081 2814
rect 2025 2760 2081 2762
rect 2450 2814 2506 2816
rect 2450 2762 2452 2814
rect 2452 2762 2504 2814
rect 2504 2762 2506 2814
rect 2450 2760 2506 2762
rect 2882 2814 2938 2816
rect 2882 2762 2884 2814
rect 2884 2762 2936 2814
rect 2936 2762 2938 2814
rect 2882 2760 2938 2762
rect 3264 2791 3320 2793
rect 3264 2739 3266 2791
rect 3266 2739 3318 2791
rect 3318 2739 3320 2791
rect 3264 2737 3320 2739
rect 3660 2791 3716 2793
rect 3660 2739 3662 2791
rect 3662 2739 3714 2791
rect 3714 2739 3716 2791
rect 3660 2737 3716 2739
rect 2025 2024 2081 2026
rect 2025 1972 2027 2024
rect 2027 1972 2079 2024
rect 2079 1972 2081 2024
rect 2025 1970 2081 1972
rect 2450 2024 2506 2026
rect 2450 1972 2452 2024
rect 2452 1972 2504 2024
rect 2504 1972 2506 2024
rect 2450 1970 2506 1972
rect 2882 2024 2938 2026
rect 2882 1972 2884 2024
rect 2884 1972 2936 2024
rect 2936 1972 2938 2024
rect 2882 1970 2938 1972
rect 3264 2001 3320 2003
rect 3264 1949 3266 2001
rect 3266 1949 3318 2001
rect 3318 1949 3320 2001
rect 3264 1947 3320 1949
rect 3660 2001 3716 2003
rect 3660 1949 3662 2001
rect 3662 1949 3714 2001
rect 3714 1949 3716 2001
rect 3660 1947 3716 1949
rect 2025 1234 2081 1236
rect 2025 1182 2027 1234
rect 2027 1182 2079 1234
rect 2079 1182 2081 1234
rect 2025 1180 2081 1182
rect 2450 1234 2506 1236
rect 2450 1182 2452 1234
rect 2452 1182 2504 1234
rect 2504 1182 2506 1234
rect 2450 1180 2506 1182
rect 2882 1234 2938 1236
rect 2882 1182 2884 1234
rect 2884 1182 2936 1234
rect 2936 1182 2938 1234
rect 2882 1180 2938 1182
rect 3264 1211 3320 1213
rect 3264 1159 3266 1211
rect 3266 1159 3318 1211
rect 3318 1159 3320 1211
rect 3264 1157 3320 1159
rect 3660 1211 3716 1213
rect 3660 1159 3662 1211
rect 3662 1159 3714 1211
rect 3714 1159 3716 1211
rect 3660 1157 3716 1159
rect 2025 444 2081 446
rect 570 421 626 423
rect 570 369 572 421
rect 572 369 624 421
rect 624 369 626 421
rect 570 367 626 369
rect 966 421 1022 423
rect 966 369 968 421
rect 968 369 1020 421
rect 1020 369 1022 421
rect 2025 392 2027 444
rect 2027 392 2079 444
rect 2079 392 2081 444
rect 2025 390 2081 392
rect 2450 444 2506 446
rect 2450 392 2452 444
rect 2452 392 2504 444
rect 2504 392 2506 444
rect 2450 390 2506 392
rect 2882 444 2938 446
rect 2882 392 2884 444
rect 2884 392 2936 444
rect 2936 392 2938 444
rect 2882 390 2938 392
rect 3264 421 3320 423
rect 966 367 1022 369
rect 3264 369 3266 421
rect 3266 369 3318 421
rect 3318 369 3320 421
rect 3264 367 3320 369
rect 3660 421 3716 423
rect 3660 369 3662 421
rect 3662 369 3714 421
rect 3714 369 3716 421
rect 3660 367 3716 369
<< metal3 >>
rect 2004 2816 2102 2837
rect 2004 2760 2025 2816
rect 2081 2760 2102 2816
rect 2004 2739 2102 2760
rect 2429 2816 2527 2837
rect 2429 2760 2450 2816
rect 2506 2760 2527 2816
rect 2429 2739 2527 2760
rect 2861 2816 2959 2837
rect 2861 2760 2882 2816
rect 2938 2760 2959 2816
rect 2861 2739 2959 2760
rect 3243 2793 3341 2814
rect 3243 2737 3264 2793
rect 3320 2737 3341 2793
rect 3243 2716 3341 2737
rect 3639 2793 3737 2814
rect 3639 2737 3660 2793
rect 3716 2737 3737 2793
rect 3639 2716 3737 2737
rect 2004 2026 2102 2047
rect 2004 1970 2025 2026
rect 2081 1970 2102 2026
rect 2004 1949 2102 1970
rect 2429 2026 2527 2047
rect 2429 1970 2450 2026
rect 2506 1970 2527 2026
rect 2429 1949 2527 1970
rect 2861 2026 2959 2047
rect 2861 1970 2882 2026
rect 2938 1970 2959 2026
rect 2861 1949 2959 1970
rect 3243 2003 3341 2024
rect 3243 1947 3264 2003
rect 3320 1947 3341 2003
rect 3243 1926 3341 1947
rect 3639 2003 3737 2024
rect 3639 1947 3660 2003
rect 3716 1947 3737 2003
rect 3639 1926 3737 1947
rect 2004 1236 2102 1257
rect 2004 1180 2025 1236
rect 2081 1180 2102 1236
rect 2004 1159 2102 1180
rect 2429 1236 2527 1257
rect 2429 1180 2450 1236
rect 2506 1180 2527 1236
rect 2429 1159 2527 1180
rect 2861 1236 2959 1257
rect 2861 1180 2882 1236
rect 2938 1180 2959 1236
rect 2861 1159 2959 1180
rect 3243 1213 3341 1234
rect 3243 1157 3264 1213
rect 3320 1157 3341 1213
rect 3243 1136 3341 1157
rect 3639 1213 3737 1234
rect 3639 1157 3660 1213
rect 3716 1157 3737 1213
rect 3639 1136 3737 1157
rect 2004 446 2102 467
rect 549 423 647 444
rect 549 367 570 423
rect 626 367 647 423
rect 549 346 647 367
rect 945 423 1043 444
rect 945 367 966 423
rect 1022 367 1043 423
rect 2004 390 2025 446
rect 2081 390 2102 446
rect 2004 369 2102 390
rect 2429 446 2527 467
rect 2429 390 2450 446
rect 2506 390 2527 446
rect 2429 369 2527 390
rect 2861 446 2959 467
rect 2861 390 2882 446
rect 2938 390 2959 446
rect 2861 369 2959 390
rect 3243 423 3341 444
rect 945 346 1043 367
rect 3243 367 3264 423
rect 3320 367 3341 423
rect 3243 346 3341 367
rect 3639 423 3737 444
rect 3639 367 3660 423
rect 3716 367 3737 423
rect 3639 346 3737 367
use sky130_sram_2kbyte_1rw1r_32x512_8_and3_dec  sky130_sram_2kbyte_1rw1r_32x512_8_and3_dec_0
timestamp 1707688321
transform 1 0 1782 0 -1 3160
box 0 -60 2072 490
use sky130_sram_2kbyte_1rw1r_32x512_8_and3_dec  sky130_sram_2kbyte_1rw1r_32x512_8_and3_dec_1
timestamp 1707688321
transform 1 0 1782 0 1 2370
box 0 -60 2072 490
use sky130_sram_2kbyte_1rw1r_32x512_8_and3_dec  sky130_sram_2kbyte_1rw1r_32x512_8_and3_dec_2
timestamp 1707688321
transform 1 0 1782 0 -1 2370
box 0 -60 2072 490
use sky130_sram_2kbyte_1rw1r_32x512_8_and3_dec  sky130_sram_2kbyte_1rw1r_32x512_8_and3_dec_3
timestamp 1707688321
transform 1 0 1782 0 1 1580
box 0 -60 2072 490
use sky130_sram_2kbyte_1rw1r_32x512_8_and3_dec  sky130_sram_2kbyte_1rw1r_32x512_8_and3_dec_4
timestamp 1707688321
transform 1 0 1782 0 -1 1580
box 0 -60 2072 490
use sky130_sram_2kbyte_1rw1r_32x512_8_and3_dec  sky130_sram_2kbyte_1rw1r_32x512_8_and3_dec_5
timestamp 1707688321
transform 1 0 1782 0 1 790
box 0 -60 2072 490
use sky130_sram_2kbyte_1rw1r_32x512_8_and3_dec  sky130_sram_2kbyte_1rw1r_32x512_8_and3_dec_6
timestamp 1707688321
transform 1 0 1782 0 -1 790
box 0 -60 2072 490
use sky130_sram_2kbyte_1rw1r_32x512_8_and3_dec  sky130_sram_2kbyte_1rw1r_32x512_8_and3_dec_7
timestamp 1707688321
transform 1 0 1782 0 1 0
box 0 -60 2072 490
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_0
timestamp 1707688321
transform 1 0 2020 0 1 2751
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_1
timestamp 1707688321
transform 1 0 3259 0 1 2728
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_2
timestamp 1707688321
transform 1 0 2020 0 1 1961
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_3
timestamp 1707688321
transform 1 0 3259 0 1 1938
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_4
timestamp 1707688321
transform 1 0 2020 0 1 1171
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_5
timestamp 1707688321
transform 1 0 3259 0 1 1148
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_6
timestamp 1707688321
transform 1 0 2020 0 1 381
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_7
timestamp 1707688321
transform 1 0 3259 0 1 358
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_8
timestamp 1707688321
transform 1 0 565 0 1 358
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_9
timestamp 1707688321
transform 1 0 3655 0 1 2728
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_10
timestamp 1707688321
transform 1 0 2877 0 1 2751
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_11
timestamp 1707688321
transform 1 0 2445 0 1 2751
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_12
timestamp 1707688321
transform 1 0 3655 0 1 1938
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_13
timestamp 1707688321
transform 1 0 2877 0 1 1961
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_14
timestamp 1707688321
transform 1 0 2445 0 1 1961
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_15
timestamp 1707688321
transform 1 0 3655 0 1 1148
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_16
timestamp 1707688321
transform 1 0 2877 0 1 1171
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_17
timestamp 1707688321
transform 1 0 2445 0 1 1171
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_18
timestamp 1707688321
transform 1 0 3655 0 1 358
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_19
timestamp 1707688321
transform 1 0 2877 0 1 381
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_20
timestamp 1707688321
transform 1 0 2445 0 1 381
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_7  sky130_sram_2kbyte_1rw1r_32x512_8_contact_7_21
timestamp 1707688321
transform 1 0 961 0 1 358
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_0
timestamp 1707688321
transform 1 0 1607 0 1 2844
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_1
timestamp 1707688321
transform 1 0 225 0 1 2844
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_2
timestamp 1707688321
transform 1 0 1527 0 1 2934
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_3
timestamp 1707688321
transform 1 0 145 0 1 2934
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_4
timestamp 1707688321
transform 1 0 1447 0 1 3046
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_5
timestamp 1707688321
transform 1 0 65 0 1 3046
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_6
timestamp 1707688321
transform 1 0 1113 0 1 877
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_7
timestamp 1707688321
transform 1 0 1113 0 1 637
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_14  sky130_sram_2kbyte_1rw1r_32x512_8_contact_14_8
timestamp 1707688321
transform 1 0 1113 0 1 87
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_17  sky130_sram_2kbyte_1rw1r_32x512_8_contact_17_0
timestamp 1707688321
transform 1 0 1603 0 1 2848
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_17  sky130_sram_2kbyte_1rw1r_32x512_8_contact_17_1
timestamp 1707688321
transform 1 0 1523 0 1 2938
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_17  sky130_sram_2kbyte_1rw1r_32x512_8_contact_17_2
timestamp 1707688321
transform 1 0 1443 0 1 3050
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_17  sky130_sram_2kbyte_1rw1r_32x512_8_contact_17_3
timestamp 1707688321
transform 1 0 1603 0 1 2624
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_17  sky130_sram_2kbyte_1rw1r_32x512_8_contact_17_4
timestamp 1707688321
transform 1 0 1523 0 1 2534
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_17  sky130_sram_2kbyte_1rw1r_32x512_8_contact_17_5
timestamp 1707688321
transform 1 0 1203 0 1 2422
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_17  sky130_sram_2kbyte_1rw1r_32x512_8_contact_17_6
timestamp 1707688321
transform 1 0 1603 0 1 2058
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_17  sky130_sram_2kbyte_1rw1r_32x512_8_contact_17_7
timestamp 1707688321
transform 1 0 1283 0 1 2148
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_17  sky130_sram_2kbyte_1rw1r_32x512_8_contact_17_8
timestamp 1707688321
transform 1 0 1443 0 1 2260
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_17  sky130_sram_2kbyte_1rw1r_32x512_8_contact_17_9
timestamp 1707688321
transform 1 0 1603 0 1 1834
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_17  sky130_sram_2kbyte_1rw1r_32x512_8_contact_17_10
timestamp 1707688321
transform 1 0 1283 0 1 1744
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_17  sky130_sram_2kbyte_1rw1r_32x512_8_contact_17_11
timestamp 1707688321
transform 1 0 1203 0 1 1632
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_17  sky130_sram_2kbyte_1rw1r_32x512_8_contact_17_12
timestamp 1707688321
transform 1 0 1363 0 1 1268
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_17  sky130_sram_2kbyte_1rw1r_32x512_8_contact_17_13
timestamp 1707688321
transform 1 0 1523 0 1 1358
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_17  sky130_sram_2kbyte_1rw1r_32x512_8_contact_17_14
timestamp 1707688321
transform 1 0 1443 0 1 1470
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_17  sky130_sram_2kbyte_1rw1r_32x512_8_contact_17_15
timestamp 1707688321
transform 1 0 1363 0 1 1044
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_17  sky130_sram_2kbyte_1rw1r_32x512_8_contact_17_16
timestamp 1707688321
transform 1 0 1523 0 1 954
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_17  sky130_sram_2kbyte_1rw1r_32x512_8_contact_17_17
timestamp 1707688321
transform 1 0 1203 0 1 842
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_17  sky130_sram_2kbyte_1rw1r_32x512_8_contact_17_18
timestamp 1707688321
transform 1 0 1363 0 1 478
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_17  sky130_sram_2kbyte_1rw1r_32x512_8_contact_17_19
timestamp 1707688321
transform 1 0 1283 0 1 568
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_17  sky130_sram_2kbyte_1rw1r_32x512_8_contact_17_20
timestamp 1707688321
transform 1 0 1443 0 1 680
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_17  sky130_sram_2kbyte_1rw1r_32x512_8_contact_17_21
timestamp 1707688321
transform 1 0 1363 0 1 254
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_17  sky130_sram_2kbyte_1rw1r_32x512_8_contact_17_22
timestamp 1707688321
transform 1 0 1283 0 1 164
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_17  sky130_sram_2kbyte_1rw1r_32x512_8_contact_17_23
timestamp 1707688321
transform 1 0 1203 0 1 52
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_17  sky130_sram_2kbyte_1rw1r_32x512_8_contact_17_24
timestamp 1707688321
transform 1 0 221 0 1 931
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_17  sky130_sram_2kbyte_1rw1r_32x512_8_contact_17_25
timestamp 1707688321
transform 1 0 141 0 1 591
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_17  sky130_sram_2kbyte_1rw1r_32x512_8_contact_17_26
timestamp 1707688321
transform 1 0 61 0 1 141
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_0
timestamp 1707688321
transform 1 0 2021 0 1 2756
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_1
timestamp 1707688321
transform 1 0 3260 0 1 2733
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_2
timestamp 1707688321
transform 1 0 2021 0 1 1966
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_3
timestamp 1707688321
transform 1 0 3260 0 1 1943
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_4
timestamp 1707688321
transform 1 0 2021 0 1 1176
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_5
timestamp 1707688321
transform 1 0 3260 0 1 1153
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_6
timestamp 1707688321
transform 1 0 2021 0 1 386
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_7
timestamp 1707688321
transform 1 0 3260 0 1 363
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_8
timestamp 1707688321
transform 1 0 566 0 1 363
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_9
timestamp 1707688321
transform 1 0 3656 0 1 2733
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_10
timestamp 1707688321
transform 1 0 2878 0 1 2756
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_11
timestamp 1707688321
transform 1 0 2446 0 1 2756
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_12
timestamp 1707688321
transform 1 0 3656 0 1 1943
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_13
timestamp 1707688321
transform 1 0 2878 0 1 1966
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_14
timestamp 1707688321
transform 1 0 2446 0 1 1966
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_15
timestamp 1707688321
transform 1 0 3656 0 1 1153
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_16
timestamp 1707688321
transform 1 0 2878 0 1 1176
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_17
timestamp 1707688321
transform 1 0 2446 0 1 1176
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_18
timestamp 1707688321
transform 1 0 3656 0 1 363
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_19
timestamp 1707688321
transform 1 0 2878 0 1 386
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_20
timestamp 1707688321
transform 1 0 2446 0 1 386
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_21
timestamp 1707688321
transform 1 0 962 0 1 363
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_22
timestamp 1707688321
transform 1 0 1110 0 1 878
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_23
timestamp 1707688321
transform 1 0 1110 0 1 638
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_19  sky130_sram_2kbyte_1rw1r_32x512_8_contact_19_24
timestamp 1707688321
transform 1 0 1110 0 1 88
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_20  sky130_sram_2kbyte_1rw1r_32x512_8_contact_20_0
timestamp 1707688321
transform 1 0 1364 0 1 1069
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_20  sky130_sram_2kbyte_1rw1r_32x512_8_contact_20_1
timestamp 1707688321
transform 1 0 1284 0 1 674
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_20  sky130_sram_2kbyte_1rw1r_32x512_8_contact_20_2
timestamp 1707688321
transform 1 0 1204 0 1 279
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_pinv_dec  sky130_sram_2kbyte_1rw1r_32x512_8_pinv_dec_0
timestamp 1707688321
transform 1 0 400 0 1 790
box 44 0 760 490
use sky130_sram_2kbyte_1rw1r_32x512_8_pinv_dec  sky130_sram_2kbyte_1rw1r_32x512_8_pinv_dec_1
timestamp 1707688321
transform 1 0 400 0 -1 790
box 44 0 760 490
use sky130_sram_2kbyte_1rw1r_32x512_8_pinv_dec  sky130_sram_2kbyte_1rw1r_32x512_8_pinv_dec_2
timestamp 1707688321
transform 1 0 400 0 1 0
box 44 0 760 490
<< labels >>
rlabel metal3 s 945 346 1043 444 4 vdd
port 1 nsew
rlabel metal3 s 2861 369 2959 467 4 vdd
port 1 nsew
rlabel metal3 s 3639 346 3737 444 4 vdd
port 1 nsew
rlabel metal3 s 2429 1159 2527 1257 4 vdd
port 1 nsew
rlabel metal3 s 3639 2716 3737 2814 4 vdd
port 1 nsew
rlabel metal3 s 2861 1159 2959 1257 4 vdd
port 1 nsew
rlabel metal3 s 2429 369 2527 467 4 vdd
port 1 nsew
rlabel metal3 s 2861 1949 2959 2047 4 vdd
port 1 nsew
rlabel metal3 s 2861 2739 2959 2837 4 vdd
port 1 nsew
rlabel metal3 s 3639 1926 3737 2024 4 vdd
port 1 nsew
rlabel metal3 s 2429 1949 2527 2047 4 vdd
port 1 nsew
rlabel metal3 s 2429 2739 2527 2837 4 vdd
port 1 nsew
rlabel metal3 s 3639 1136 3737 1234 4 vdd
port 1 nsew
rlabel metal3 s 3243 2716 3341 2814 4 gnd
port 2 nsew
rlabel metal3 s 2004 1949 2102 2047 4 gnd
port 2 nsew
rlabel metal3 s 549 346 647 444 4 gnd
port 2 nsew
rlabel metal3 s 3243 1926 3341 2024 4 gnd
port 2 nsew
rlabel metal3 s 2004 369 2102 467 4 gnd
port 2 nsew
rlabel metal3 s 3243 1136 3341 1234 4 gnd
port 2 nsew
rlabel metal3 s 3243 346 3341 444 4 gnd
port 2 nsew
rlabel metal3 s 2004 1159 2102 1257 4 gnd
port 2 nsew
rlabel metal3 s 2004 2739 2102 2837 4 gnd
port 2 nsew
rlabel metal1 s 71 141 117 199 4 in_0
port 3 nsew
rlabel metal1 s 151 591 197 649 4 in_1
port 4 nsew
rlabel metal1 s 231 931 277 989 4 in_2
port 5 nsew
rlabel locali s 3547 120 3547 120 4 out_0
rlabel locali s 3547 670 3547 670 4 out_1
rlabel locali s 3547 910 3547 910 4 out_2
rlabel locali s 3547 1460 3547 1460 4 out_3
rlabel locali s 3547 1700 3547 1700 4 out_4
rlabel locali s 3547 2250 3547 2250 4 out_5
rlabel locali s 3547 2490 3547 2490 4 out_6
rlabel locali s 3547 3040 3547 3040 4 out_7
<< properties >>
string FIXED_BBOX 0 0 3836 3160
string GDS_END 212846
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_START 193464
<< end >>
