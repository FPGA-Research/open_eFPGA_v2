magic
tech sky130A
timestamp 1707688321
<< metal1 >>
rect 0 0 3 570
rect 253 0 256 570
<< via1 >>
rect 3 0 253 570
<< metal2 >>
rect 0 0 3 570
rect 253 0 256 570
<< properties >>
string GDS_END 88479722
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 88470374
<< end >>
