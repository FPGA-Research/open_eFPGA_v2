magic
tech sky130B
timestamp 1707688321
<< metal1 >>
rect 0 0 3 186
rect 381 0 384 186
<< via1 >>
rect 3 0 381 186
<< metal2 >>
rect 0 0 3 186
rect 381 0 384 186
<< properties >>
string GDS_END 94182640
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 94177900
<< end >>
