magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -122 -66 219 366
<< mvpmos >>
rect 0 0 100 300
<< mvpdiff >>
rect -56 250 0 300
rect -56 216 -45 250
rect -11 216 0 250
rect -56 182 0 216
rect -56 148 -45 182
rect -11 148 0 182
rect -56 114 0 148
rect -56 80 -45 114
rect -11 80 0 114
rect -56 46 0 80
rect -56 12 -45 46
rect -11 12 0 46
rect -56 0 0 12
rect 100 250 153 300
rect 100 216 111 250
rect 145 216 153 250
rect 100 182 153 216
rect 100 148 111 182
rect 145 148 153 182
rect 100 114 153 148
rect 100 80 111 114
rect 145 80 153 114
rect 100 46 153 80
rect 100 12 111 46
rect 145 12 153 46
rect 100 0 153 12
<< mvpdiffc >>
rect -45 216 -11 250
rect -45 148 -11 182
rect -45 80 -11 114
rect -45 12 -11 46
rect 111 216 145 250
rect 111 148 145 182
rect 111 80 145 114
rect 111 12 145 46
<< poly >>
rect 0 300 100 326
rect 0 -26 100 0
<< locali >>
rect -45 250 -11 266
rect -45 182 -11 216
rect -45 114 -11 148
rect -45 46 -11 80
rect -45 -4 -11 12
rect 111 250 145 266
rect 111 182 145 216
rect 111 114 145 148
rect 111 46 145 80
rect 111 -4 145 12
use hvDFL1sd2_CDNS_52468879185277  hvDFL1sd2_CDNS_52468879185277_0
timestamp 1707688321
transform -1 0 0 0 1 0
box 0 0 1 1
use hvDFL1sd_CDNS_52468879185669  hvDFL1sd_CDNS_52468879185669_0
timestamp 1707688321
transform 1 0 100 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 131 -28 131 0 FreeSans 300 0 0 0 S
flabel comment s 128 131 128 131 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 86353452
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86352432
<< end >>
