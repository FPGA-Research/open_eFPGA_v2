magic
tech sky130A
timestamp 1707688321
<< metal1 >>
rect 0 0 3 154
rect 381 0 384 154
<< via1 >>
rect 3 0 381 154
<< metal2 >>
rect 0 0 3 154
rect 381 0 384 154
<< properties >>
string GDS_END 91767086
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 91763114
<< end >>
