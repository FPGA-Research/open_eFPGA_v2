magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< pwell >>
rect 467 350 491 401
<< obsli1 >>
rect 0 0 876 918
<< obsm1 >>
rect 0 852 876 918
rect 0 66 66 852
rect 113 491 141 824
rect 169 519 197 852
rect 225 491 253 824
rect 281 519 309 852
rect 337 491 365 824
rect 411 491 465 824
rect 511 491 539 824
rect 567 519 595 852
rect 623 491 651 824
rect 679 519 707 852
rect 735 491 763 824
rect 113 427 763 491
rect 113 94 141 427
rect 169 66 197 399
rect 225 94 253 427
rect 281 66 309 399
rect 337 94 365 427
rect 411 94 465 427
rect 511 94 539 427
rect 567 66 595 399
rect 623 94 651 427
rect 679 66 707 399
rect 735 94 763 427
rect 810 66 876 852
rect 0 0 876 66
<< obsm2 >>
rect 0 852 383 918
rect 0 768 66 852
rect 411 824 465 918
rect 493 852 876 918
rect 94 796 782 824
rect 0 740 382 768
rect 0 656 66 740
rect 410 712 466 796
rect 810 768 876 852
rect 494 740 876 768
rect 94 684 782 712
rect 0 628 382 656
rect 0 544 66 628
rect 410 600 466 684
rect 810 656 876 740
rect 494 628 876 656
rect 94 572 782 600
rect 0 516 382 544
rect 0 514 66 516
rect 410 487 466 572
rect 810 544 876 628
rect 494 516 876 544
rect 810 514 876 516
rect 74 486 802 487
rect 0 432 876 486
rect 74 431 802 432
rect 0 402 66 404
rect 0 374 382 402
rect 0 290 66 374
rect 410 346 466 431
rect 810 402 876 404
rect 494 374 876 402
rect 94 318 782 346
rect 0 262 382 290
rect 0 178 66 262
rect 410 234 466 318
rect 810 290 876 374
rect 494 262 876 290
rect 94 206 782 234
rect 0 150 382 178
rect 0 66 66 150
rect 410 122 466 206
rect 810 178 876 262
rect 494 150 876 178
rect 94 94 782 122
rect 0 0 383 66
rect 411 0 465 94
rect 810 66 876 150
rect 493 0 876 66
<< metal3 >>
rect 0 852 876 918
rect 0 66 66 852
rect 126 492 186 792
rect 246 552 306 852
rect 405 492 471 792
rect 570 552 630 852
rect 690 492 750 792
rect 126 426 750 492
rect 126 126 186 426
rect 246 66 306 366
rect 405 126 471 426
rect 570 66 630 366
rect 690 126 750 426
rect 810 66 876 852
rect 0 0 876 66
<< labels >>
rlabel metal3 s 810 66 876 852 6 C0
port 1 nsew
rlabel metal3 s 570 552 630 852 6 C0
port 1 nsew
rlabel metal3 s 570 66 630 366 6 C0
port 1 nsew
rlabel metal3 s 246 552 306 852 6 C0
port 1 nsew
rlabel metal3 s 246 66 306 366 6 C0
port 1 nsew
rlabel metal3 s 0 852 876 918 6 C0
port 1 nsew
rlabel metal3 s 0 66 66 852 6 C0
port 1 nsew
rlabel metal3 s 0 0 876 66 6 C0
port 1 nsew
rlabel metal3 s 690 492 750 792 6 C1
port 2 nsew
rlabel metal3 s 690 126 750 426 6 C1
port 2 nsew
rlabel metal3 s 405 492 471 792 6 C1
port 2 nsew
rlabel metal3 s 405 126 471 426 6 C1
port 2 nsew
rlabel metal3 s 126 492 186 792 6 C1
port 2 nsew
rlabel metal3 s 126 426 750 492 6 C1
port 2 nsew
rlabel metal3 s 126 126 186 426 6 C1
port 2 nsew
rlabel pwell s 467 350 491 401 6 SUB
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 876 918
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 149780
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 135732
string device primitive
<< end >>
