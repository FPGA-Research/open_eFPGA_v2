magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -119 -66 1775 266
<< mvpmos >>
rect 0 0 800 200
rect 856 0 1656 200
<< mvpdiff >>
rect -53 182 0 200
rect -53 148 -45 182
rect -11 148 0 182
rect -53 114 0 148
rect -53 80 -45 114
rect -11 80 0 114
rect -53 46 0 80
rect -53 12 -45 46
rect -11 12 0 46
rect -53 0 0 12
rect 800 182 856 200
rect 800 148 811 182
rect 845 148 856 182
rect 800 114 856 148
rect 800 80 811 114
rect 845 80 856 114
rect 800 46 856 80
rect 800 12 811 46
rect 845 12 856 46
rect 800 0 856 12
rect 1656 182 1709 200
rect 1656 148 1667 182
rect 1701 148 1709 182
rect 1656 114 1709 148
rect 1656 80 1667 114
rect 1701 80 1709 114
rect 1656 46 1709 80
rect 1656 12 1667 46
rect 1701 12 1709 46
rect 1656 0 1709 12
<< mvpdiffc >>
rect -45 148 -11 182
rect -45 80 -11 114
rect -45 12 -11 46
rect 811 148 845 182
rect 811 80 845 114
rect 811 12 845 46
rect 1667 148 1701 182
rect 1667 80 1701 114
rect 1667 12 1701 46
<< poly >>
rect 0 200 800 226
rect 856 200 1656 226
rect 0 -26 800 0
rect 856 -26 1656 0
<< locali >>
rect -45 182 -11 198
rect -45 114 -11 148
rect -45 46 -11 80
rect -45 -4 -11 12
rect 811 182 845 198
rect 811 114 845 148
rect 811 46 845 80
rect 811 -4 845 12
rect 1667 182 1701 198
rect 1667 114 1701 148
rect 1667 46 1701 80
rect 1667 -4 1701 12
use hvDFL1sd2_CDNS_52468879185110  hvDFL1sd2_CDNS_52468879185110_0
timestamp 1707688321
transform 1 0 800 0 1 0
box 0 0 1 1
use hvDFL1sd_CDNS_5246887918589  hvDFL1sd_CDNS_5246887918589_0
timestamp 1707688321
transform -1 0 0 0 1 0
box 0 0 1 1
use hvDFL1sd_CDNS_5246887918589  hvDFL1sd_CDNS_5246887918589_1
timestamp 1707688321
transform 1 0 1656 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 97 -28 97 0 FreeSans 300 0 0 0 S
flabel comment s 828 97 828 97 0 FreeSans 300 0 0 0 D
flabel comment s 1684 97 1684 97 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 87859676
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87858158
<< end >>
