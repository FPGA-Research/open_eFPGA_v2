magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -76 -26 372 626
<< mvnmos >>
rect 0 0 120 600
rect 176 0 296 600
<< mvndiff >>
rect -50 0 0 600
rect 296 0 346 600
<< poly >>
rect 0 600 120 626
rect 0 -26 120 0
rect 176 600 296 626
rect 176 -26 296 0
<< metal1 >>
rect -51 -16 -5 546
rect 125 -16 171 546
rect 301 -16 347 546
use hvDFM1sd2_CDNS_52468879185154  hvDFM1sd2_CDNS_52468879185154_0
timestamp 1707688321
transform 1 0 120 0 1 0
box -26 -26 82 626
use hvDFM1sd_CDNS_52468879185149  hvDFM1sd_CDNS_52468879185149_0
timestamp 1707688321
transform -1 0 0 0 1 0
box -26 -26 79 626
use hvDFM1sd_CDNS_52468879185149  hvDFM1sd_CDNS_52468879185149_1
timestamp 1707688321
transform 1 0 296 0 1 0
box -26 -26 79 626
<< labels >>
flabel comment s -28 265 -28 265 0 FreeSans 300 0 0 0 S
flabel comment s 148 265 148 265 0 FreeSans 300 0 0 0 D
flabel comment s 324 265 324 265 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 85991986
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85990596
<< end >>
