magic
tech sky130B
timestamp 1707688321
<< metal1 >>
rect 0 0 3 282
rect 253 0 256 282
<< via1 >>
rect 3 0 253 282
<< metal2 >>
rect 0 0 3 282
rect 253 0 256 282
<< properties >>
string GDS_END 88470316
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 88465576
<< end >>
