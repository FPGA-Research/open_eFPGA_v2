magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect 0 2152 1591 2424
rect 0 272 272 2152
rect 1319 272 1591 2152
rect 0 0 1591 272
<< pwell >>
rect 332 332 1259 2092
<< mvnmosesd >>
tri 695 1712 735 1752 ne
tri 695 672 735 712 se
rect 735 672 855 1752
tri 855 1712 895 1752 nw
tri 855 672 895 712 sw
<< mvndiff >>
rect 594 1712 695 1752
tri 695 1712 735 1752 sw
rect 594 1635 735 1712
rect 594 1601 602 1635
rect 636 1601 735 1635
rect 594 1567 735 1601
rect 594 1533 602 1567
rect 636 1533 735 1567
rect 594 1499 735 1533
rect 594 1465 602 1499
rect 636 1465 735 1499
rect 594 1431 735 1465
rect 594 1397 602 1431
rect 636 1397 735 1431
rect 594 1363 735 1397
rect 594 1329 602 1363
rect 636 1329 735 1363
rect 594 1295 735 1329
rect 594 1261 602 1295
rect 636 1261 735 1295
rect 594 1227 735 1261
rect 594 1193 602 1227
rect 636 1193 735 1227
rect 594 1159 735 1193
rect 594 1125 602 1159
rect 636 1125 735 1159
rect 594 1091 735 1125
rect 594 1057 602 1091
rect 636 1057 735 1091
rect 594 1023 735 1057
rect 594 989 602 1023
rect 636 989 735 1023
rect 594 955 735 989
rect 594 921 602 955
rect 636 921 735 955
rect 594 887 735 921
rect 594 853 602 887
rect 636 853 735 887
rect 594 819 735 853
rect 594 785 602 819
rect 636 785 735 819
rect 594 751 735 785
rect 594 717 602 751
rect 636 717 735 751
rect 594 712 735 717
rect 594 672 695 712
tri 695 672 735 712 nw
tri 855 1712 895 1752 se
rect 895 1712 996 1752
rect 855 1635 996 1712
rect 855 1601 946 1635
rect 980 1601 996 1635
rect 855 1567 996 1601
rect 855 1533 946 1567
rect 980 1533 996 1567
rect 855 1499 996 1533
rect 855 1465 946 1499
rect 980 1465 996 1499
rect 855 1431 996 1465
rect 855 1397 946 1431
rect 980 1397 996 1431
rect 855 1363 996 1397
rect 855 1329 946 1363
rect 980 1329 996 1363
rect 855 1295 996 1329
rect 855 1261 946 1295
rect 980 1261 996 1295
rect 855 1227 996 1261
rect 855 1193 946 1227
rect 980 1193 996 1227
rect 855 1159 996 1193
rect 855 1125 946 1159
rect 980 1125 996 1159
rect 855 1091 996 1125
rect 855 1057 946 1091
rect 980 1057 996 1091
rect 855 1023 996 1057
rect 855 989 946 1023
rect 980 989 996 1023
rect 855 955 996 989
rect 855 921 946 955
rect 980 921 996 955
rect 855 887 996 921
rect 855 853 946 887
rect 980 853 996 887
rect 855 819 996 853
rect 855 785 946 819
rect 980 785 996 819
rect 855 751 996 785
rect 855 717 946 751
rect 980 717 996 751
rect 855 712 996 717
tri 855 672 895 712 ne
rect 895 672 996 712
<< mvndiffc >>
rect 602 1601 636 1635
rect 602 1533 636 1567
rect 602 1465 636 1499
rect 602 1397 636 1431
rect 602 1329 636 1363
rect 602 1261 636 1295
rect 602 1193 636 1227
rect 602 1125 636 1159
rect 602 1057 636 1091
rect 602 989 636 1023
rect 602 921 636 955
rect 602 853 636 887
rect 602 785 636 819
rect 602 717 636 751
rect 946 1601 980 1635
rect 946 1533 980 1567
rect 946 1465 980 1499
rect 946 1397 980 1431
rect 946 1329 980 1363
rect 946 1261 980 1295
rect 946 1193 980 1227
rect 946 1125 980 1159
rect 946 1057 980 1091
rect 946 989 980 1023
rect 946 921 980 955
rect 946 853 980 887
rect 946 785 980 819
rect 946 717 980 751
<< mvpsubdiff >>
rect 358 2013 1233 2066
rect 358 1979 473 2013
rect 507 1979 541 2013
rect 575 1979 609 2013
rect 643 1979 677 2013
rect 711 1979 745 2013
rect 779 1979 813 2013
rect 847 1979 881 2013
rect 915 1979 949 2013
rect 983 1979 1017 2013
rect 1051 1979 1085 2013
rect 1119 1979 1233 2013
rect 358 1926 1233 1979
rect 358 1791 462 1926
rect 358 1757 404 1791
rect 438 1757 462 1791
rect 358 1723 462 1757
rect 1129 1791 1233 1926
rect 1129 1757 1156 1791
rect 1190 1757 1233 1791
rect 358 1689 404 1723
rect 438 1689 462 1723
rect 358 1655 462 1689
rect 358 1621 404 1655
rect 438 1621 462 1655
rect 358 1587 462 1621
rect 358 1553 404 1587
rect 438 1553 462 1587
rect 358 1519 462 1553
rect 358 1485 404 1519
rect 438 1485 462 1519
rect 358 1451 462 1485
rect 358 1417 404 1451
rect 438 1417 462 1451
rect 358 1383 462 1417
rect 358 1349 404 1383
rect 438 1349 462 1383
rect 358 1315 462 1349
rect 358 1281 404 1315
rect 438 1281 462 1315
rect 358 1247 462 1281
rect 358 1213 404 1247
rect 438 1213 462 1247
rect 358 1179 462 1213
rect 358 1145 404 1179
rect 438 1145 462 1179
rect 358 1111 462 1145
rect 358 1077 404 1111
rect 438 1077 462 1111
rect 358 1043 462 1077
rect 358 1009 404 1043
rect 438 1009 462 1043
rect 358 975 462 1009
rect 358 941 404 975
rect 438 941 462 975
rect 358 907 462 941
rect 358 873 404 907
rect 438 873 462 907
rect 358 839 462 873
rect 358 805 404 839
rect 438 805 462 839
rect 358 771 462 805
rect 358 737 404 771
rect 438 737 462 771
rect 358 703 462 737
rect 358 669 404 703
rect 438 669 462 703
rect 1129 1723 1233 1757
rect 1129 1689 1156 1723
rect 1190 1689 1233 1723
rect 1129 1655 1233 1689
rect 1129 1621 1156 1655
rect 1190 1621 1233 1655
rect 1129 1587 1233 1621
rect 1129 1553 1156 1587
rect 1190 1553 1233 1587
rect 1129 1519 1233 1553
rect 1129 1485 1156 1519
rect 1190 1485 1233 1519
rect 1129 1451 1233 1485
rect 1129 1417 1156 1451
rect 1190 1417 1233 1451
rect 1129 1383 1233 1417
rect 1129 1349 1156 1383
rect 1190 1349 1233 1383
rect 1129 1315 1233 1349
rect 1129 1281 1156 1315
rect 1190 1281 1233 1315
rect 1129 1247 1233 1281
rect 1129 1213 1156 1247
rect 1190 1213 1233 1247
rect 1129 1179 1233 1213
rect 1129 1145 1156 1179
rect 1190 1145 1233 1179
rect 1129 1111 1233 1145
rect 1129 1077 1156 1111
rect 1190 1077 1233 1111
rect 1129 1043 1233 1077
rect 1129 1009 1156 1043
rect 1190 1009 1233 1043
rect 1129 975 1233 1009
rect 1129 941 1156 975
rect 1190 941 1233 975
rect 1129 907 1233 941
rect 1129 873 1156 907
rect 1190 873 1233 907
rect 1129 839 1233 873
rect 1129 805 1156 839
rect 1190 805 1233 839
rect 1129 771 1233 805
rect 1129 737 1156 771
rect 1190 737 1233 771
rect 1129 703 1233 737
rect 358 635 462 669
rect 358 601 404 635
rect 438 601 462 635
rect 358 567 462 601
rect 358 533 404 567
rect 438 533 462 567
rect 1129 669 1156 703
rect 1190 669 1233 703
rect 1129 635 1233 669
rect 1129 601 1156 635
rect 1190 601 1233 635
rect 1129 567 1233 601
rect 358 498 462 533
rect 1129 533 1156 567
rect 1190 533 1233 567
rect 1129 498 1233 533
rect 358 445 1233 498
rect 358 411 473 445
rect 507 411 541 445
rect 575 411 609 445
rect 643 411 677 445
rect 711 411 745 445
rect 779 411 813 445
rect 847 411 881 445
rect 915 411 949 445
rect 983 411 1017 445
rect 1051 411 1085 445
rect 1119 411 1233 445
rect 358 358 1233 411
<< mvnsubdiff >>
rect 66 2305 1525 2358
rect 66 2271 303 2305
rect 337 2271 371 2305
rect 405 2271 439 2305
rect 473 2271 507 2305
rect 541 2271 575 2305
rect 609 2271 643 2305
rect 677 2271 711 2305
rect 745 2271 779 2305
rect 813 2271 847 2305
rect 881 2271 915 2305
rect 949 2271 983 2305
rect 1017 2271 1051 2305
rect 1085 2271 1119 2305
rect 1153 2271 1187 2305
rect 1221 2271 1255 2305
rect 1289 2271 1525 2305
rect 66 2218 1525 2271
rect 66 2092 206 2218
rect 66 2058 119 2092
rect 153 2058 206 2092
rect 1385 2092 1525 2218
rect 66 2024 206 2058
rect 66 1990 119 2024
rect 153 1990 206 2024
rect 66 1956 206 1990
rect 66 1922 119 1956
rect 153 1922 206 1956
rect 66 1888 206 1922
rect 66 1854 119 1888
rect 153 1854 206 1888
rect 66 1820 206 1854
rect 66 1786 119 1820
rect 153 1786 206 1820
rect 66 1752 206 1786
rect 66 1718 119 1752
rect 153 1718 206 1752
rect 66 1684 206 1718
rect 66 1650 119 1684
rect 153 1650 206 1684
rect 66 1616 206 1650
rect 66 1582 119 1616
rect 153 1582 206 1616
rect 66 1548 206 1582
rect 66 1514 119 1548
rect 153 1514 206 1548
rect 66 1480 206 1514
rect 66 1446 119 1480
rect 153 1446 206 1480
rect 66 1412 206 1446
rect 66 1378 119 1412
rect 153 1378 206 1412
rect 66 1344 206 1378
rect 66 1310 119 1344
rect 153 1310 206 1344
rect 66 1276 206 1310
rect 66 1242 119 1276
rect 153 1242 206 1276
rect 66 1208 206 1242
rect 66 1174 119 1208
rect 153 1174 206 1208
rect 66 1140 206 1174
rect 66 1106 119 1140
rect 153 1106 206 1140
rect 66 1072 206 1106
rect 66 1038 119 1072
rect 153 1038 206 1072
rect 66 1004 206 1038
rect 66 970 119 1004
rect 153 970 206 1004
rect 66 936 206 970
rect 66 902 119 936
rect 153 902 206 936
rect 66 868 206 902
rect 66 834 119 868
rect 153 834 206 868
rect 66 800 206 834
rect 66 766 119 800
rect 153 766 206 800
rect 66 732 206 766
rect 66 698 119 732
rect 153 698 206 732
rect 66 664 206 698
rect 66 630 119 664
rect 153 630 206 664
rect 66 596 206 630
rect 66 562 119 596
rect 153 562 206 596
rect 66 528 206 562
rect 66 494 119 528
rect 153 494 206 528
rect 66 460 206 494
rect 66 426 119 460
rect 153 426 206 460
rect 66 392 206 426
rect 66 358 119 392
rect 153 358 206 392
rect 1385 2058 1438 2092
rect 1472 2058 1525 2092
rect 1385 2024 1525 2058
rect 1385 1990 1438 2024
rect 1472 1990 1525 2024
rect 1385 1956 1525 1990
rect 1385 1922 1438 1956
rect 1472 1922 1525 1956
rect 1385 1888 1525 1922
rect 1385 1854 1438 1888
rect 1472 1854 1525 1888
rect 1385 1820 1525 1854
rect 1385 1786 1438 1820
rect 1472 1786 1525 1820
rect 1385 1752 1525 1786
rect 1385 1718 1438 1752
rect 1472 1718 1525 1752
rect 1385 1684 1525 1718
rect 1385 1650 1438 1684
rect 1472 1650 1525 1684
rect 1385 1616 1525 1650
rect 1385 1582 1438 1616
rect 1472 1582 1525 1616
rect 1385 1548 1525 1582
rect 1385 1514 1438 1548
rect 1472 1514 1525 1548
rect 1385 1480 1525 1514
rect 1385 1446 1438 1480
rect 1472 1446 1525 1480
rect 1385 1412 1525 1446
rect 1385 1378 1438 1412
rect 1472 1378 1525 1412
rect 1385 1344 1525 1378
rect 1385 1310 1438 1344
rect 1472 1310 1525 1344
rect 1385 1276 1525 1310
rect 1385 1242 1438 1276
rect 1472 1242 1525 1276
rect 1385 1208 1525 1242
rect 1385 1174 1438 1208
rect 1472 1174 1525 1208
rect 1385 1140 1525 1174
rect 1385 1106 1438 1140
rect 1472 1106 1525 1140
rect 1385 1072 1525 1106
rect 1385 1038 1438 1072
rect 1472 1038 1525 1072
rect 1385 1004 1525 1038
rect 1385 970 1438 1004
rect 1472 970 1525 1004
rect 1385 936 1525 970
rect 1385 902 1438 936
rect 1472 902 1525 936
rect 1385 868 1525 902
rect 1385 834 1438 868
rect 1472 834 1525 868
rect 1385 800 1525 834
rect 1385 766 1438 800
rect 1472 766 1525 800
rect 1385 732 1525 766
rect 1385 698 1438 732
rect 1472 698 1525 732
rect 1385 664 1525 698
rect 1385 630 1438 664
rect 1472 630 1525 664
rect 1385 596 1525 630
rect 1385 562 1438 596
rect 1472 562 1525 596
rect 1385 528 1525 562
rect 1385 494 1438 528
rect 1472 494 1525 528
rect 1385 460 1525 494
rect 1385 426 1438 460
rect 1472 426 1525 460
rect 1385 392 1525 426
rect 1385 358 1438 392
rect 1472 358 1525 392
rect 66 324 206 358
rect 66 290 119 324
rect 153 290 206 324
rect 66 256 206 290
rect 66 222 119 256
rect 153 222 206 256
rect 66 206 206 222
rect 1385 324 1525 358
rect 1385 290 1438 324
rect 1472 290 1525 324
rect 1385 256 1525 290
rect 1385 222 1438 256
rect 1472 222 1525 256
rect 1385 206 1525 222
rect 66 153 1525 206
rect 66 119 303 153
rect 337 119 371 153
rect 405 119 439 153
rect 473 119 507 153
rect 541 119 575 153
rect 609 119 643 153
rect 677 119 711 153
rect 745 119 779 153
rect 813 119 847 153
rect 881 119 915 153
rect 949 119 983 153
rect 1017 119 1051 153
rect 1085 119 1119 153
rect 1153 119 1187 153
rect 1221 119 1255 153
rect 1289 119 1525 153
rect 66 66 1525 119
<< mvpsubdiffcont >>
rect 473 1979 507 2013
rect 541 1979 575 2013
rect 609 1979 643 2013
rect 677 1979 711 2013
rect 745 1979 779 2013
rect 813 1979 847 2013
rect 881 1979 915 2013
rect 949 1979 983 2013
rect 1017 1979 1051 2013
rect 1085 1979 1119 2013
rect 404 1757 438 1791
rect 1156 1757 1190 1791
rect 404 1689 438 1723
rect 404 1621 438 1655
rect 404 1553 438 1587
rect 404 1485 438 1519
rect 404 1417 438 1451
rect 404 1349 438 1383
rect 404 1281 438 1315
rect 404 1213 438 1247
rect 404 1145 438 1179
rect 404 1077 438 1111
rect 404 1009 438 1043
rect 404 941 438 975
rect 404 873 438 907
rect 404 805 438 839
rect 404 737 438 771
rect 404 669 438 703
rect 1156 1689 1190 1723
rect 1156 1621 1190 1655
rect 1156 1553 1190 1587
rect 1156 1485 1190 1519
rect 1156 1417 1190 1451
rect 1156 1349 1190 1383
rect 1156 1281 1190 1315
rect 1156 1213 1190 1247
rect 1156 1145 1190 1179
rect 1156 1077 1190 1111
rect 1156 1009 1190 1043
rect 1156 941 1190 975
rect 1156 873 1190 907
rect 1156 805 1190 839
rect 1156 737 1190 771
rect 404 601 438 635
rect 404 533 438 567
rect 1156 669 1190 703
rect 1156 601 1190 635
rect 1156 533 1190 567
rect 473 411 507 445
rect 541 411 575 445
rect 609 411 643 445
rect 677 411 711 445
rect 745 411 779 445
rect 813 411 847 445
rect 881 411 915 445
rect 949 411 983 445
rect 1017 411 1051 445
rect 1085 411 1119 445
<< mvnsubdiffcont >>
rect 303 2271 337 2305
rect 371 2271 405 2305
rect 439 2271 473 2305
rect 507 2271 541 2305
rect 575 2271 609 2305
rect 643 2271 677 2305
rect 711 2271 745 2305
rect 779 2271 813 2305
rect 847 2271 881 2305
rect 915 2271 949 2305
rect 983 2271 1017 2305
rect 1051 2271 1085 2305
rect 1119 2271 1153 2305
rect 1187 2271 1221 2305
rect 1255 2271 1289 2305
rect 119 2058 153 2092
rect 119 1990 153 2024
rect 119 1922 153 1956
rect 119 1854 153 1888
rect 119 1786 153 1820
rect 119 1718 153 1752
rect 119 1650 153 1684
rect 119 1582 153 1616
rect 119 1514 153 1548
rect 119 1446 153 1480
rect 119 1378 153 1412
rect 119 1310 153 1344
rect 119 1242 153 1276
rect 119 1174 153 1208
rect 119 1106 153 1140
rect 119 1038 153 1072
rect 119 970 153 1004
rect 119 902 153 936
rect 119 834 153 868
rect 119 766 153 800
rect 119 698 153 732
rect 119 630 153 664
rect 119 562 153 596
rect 119 494 153 528
rect 119 426 153 460
rect 119 358 153 392
rect 1438 2058 1472 2092
rect 1438 1990 1472 2024
rect 1438 1922 1472 1956
rect 1438 1854 1472 1888
rect 1438 1786 1472 1820
rect 1438 1718 1472 1752
rect 1438 1650 1472 1684
rect 1438 1582 1472 1616
rect 1438 1514 1472 1548
rect 1438 1446 1472 1480
rect 1438 1378 1472 1412
rect 1438 1310 1472 1344
rect 1438 1242 1472 1276
rect 1438 1174 1472 1208
rect 1438 1106 1472 1140
rect 1438 1038 1472 1072
rect 1438 970 1472 1004
rect 1438 902 1472 936
rect 1438 834 1472 868
rect 1438 766 1472 800
rect 1438 698 1472 732
rect 1438 630 1472 664
rect 1438 562 1472 596
rect 1438 494 1472 528
rect 1438 426 1472 460
rect 1438 358 1472 392
rect 119 290 153 324
rect 119 222 153 256
rect 1438 290 1472 324
rect 1438 222 1472 256
rect 303 119 337 153
rect 371 119 405 153
rect 439 119 473 153
rect 507 119 541 153
rect 575 119 609 153
rect 643 119 677 153
rect 711 119 745 153
rect 779 119 813 153
rect 847 119 881 153
rect 915 119 949 153
rect 983 119 1017 153
rect 1051 119 1085 153
rect 1119 119 1153 153
rect 1187 119 1221 153
rect 1255 119 1289 153
<< poly >>
rect 655 1846 935 1866
rect 655 1812 676 1846
rect 710 1812 744 1846
rect 778 1812 812 1846
rect 846 1812 880 1846
rect 914 1812 935 1846
rect 655 1792 935 1812
tri 655 1752 695 1792 ne
rect 695 1752 895 1792
tri 895 1752 935 1792 nw
tri 655 632 695 672 se
rect 695 632 895 672
tri 895 632 935 672 sw
rect 655 558 935 632
<< polycont >>
rect 676 1812 710 1846
rect 744 1812 778 1846
rect 812 1812 846 1846
rect 880 1812 914 1846
<< locali >>
rect 66 2305 1525 2358
rect 66 2271 303 2305
rect 341 2271 371 2305
rect 413 2271 439 2305
rect 485 2271 507 2305
rect 557 2271 575 2305
rect 629 2271 643 2305
rect 677 2271 711 2305
rect 745 2271 779 2305
rect 813 2271 847 2305
rect 881 2271 915 2305
rect 949 2271 959 2305
rect 1017 2271 1031 2305
rect 1085 2271 1103 2305
rect 1153 2271 1175 2305
rect 1221 2271 1247 2305
rect 1289 2271 1525 2305
rect 66 2218 1525 2271
rect 66 2092 206 2218
rect 66 2058 119 2092
rect 153 2058 206 2092
rect 1385 2092 1525 2218
rect 66 2035 206 2058
rect 66 1990 119 2035
rect 153 1990 206 2035
rect 66 1963 206 1990
rect 66 1922 119 1963
rect 153 1922 206 1963
rect 66 1891 206 1922
rect 66 1854 119 1891
rect 153 1854 206 1891
rect 66 1820 206 1854
rect 66 1785 119 1820
rect 153 1785 206 1820
rect 66 1752 206 1785
rect 66 1713 119 1752
rect 153 1713 206 1752
rect 66 1684 206 1713
rect 66 1641 119 1684
rect 153 1641 206 1684
rect 66 1616 206 1641
rect 66 1569 119 1616
rect 153 1569 206 1616
rect 66 1548 206 1569
rect 66 1497 119 1548
rect 153 1497 206 1548
rect 66 1480 206 1497
rect 66 1425 119 1480
rect 153 1425 206 1480
rect 66 1412 206 1425
rect 66 1353 119 1412
rect 153 1353 206 1412
rect 66 1344 206 1353
rect 66 1281 119 1344
rect 153 1281 206 1344
rect 66 1276 206 1281
rect 66 1209 119 1276
rect 153 1209 206 1276
rect 66 1208 206 1209
rect 66 1174 119 1208
rect 153 1174 206 1208
rect 66 1171 206 1174
rect 66 1106 119 1171
rect 153 1106 206 1171
rect 66 1099 206 1106
rect 66 1038 119 1099
rect 153 1038 206 1099
rect 66 1027 206 1038
rect 66 970 119 1027
rect 153 970 206 1027
rect 66 955 206 970
rect 66 902 119 955
rect 153 902 206 955
rect 66 883 206 902
rect 66 834 119 883
rect 153 834 206 883
rect 66 811 206 834
rect 66 766 119 811
rect 153 766 206 811
rect 66 739 206 766
rect 66 698 119 739
rect 153 698 206 739
rect 66 667 206 698
rect 66 630 119 667
rect 153 630 206 667
rect 66 596 206 630
rect 66 561 119 596
rect 153 561 206 596
rect 66 528 206 561
rect 66 489 119 528
rect 153 489 206 528
rect 66 460 206 489
rect 66 417 119 460
rect 153 417 206 460
rect 66 392 206 417
rect 66 345 119 392
rect 153 345 206 392
rect 358 2013 1233 2066
rect 358 2003 473 2013
rect 507 2003 541 2013
rect 575 2003 609 2013
rect 358 1969 454 2003
rect 507 1979 526 2003
rect 575 1979 598 2003
rect 643 1979 677 2013
rect 711 1979 745 2013
rect 779 1979 813 2013
rect 847 1979 881 2013
rect 915 2003 949 2013
rect 983 2003 1017 2013
rect 1051 2003 1085 2013
rect 915 1979 928 2003
rect 983 1979 1000 2003
rect 1051 1979 1072 2003
rect 1119 1979 1233 2013
rect 488 1969 526 1979
rect 560 1969 598 1979
rect 632 1969 928 1979
rect 962 1969 1000 1979
rect 1034 1969 1072 1979
rect 1106 1969 1233 1979
rect 358 1924 1233 1969
rect 358 1803 498 1924
rect 358 1769 395 1803
rect 429 1791 498 1803
rect 358 1757 404 1769
rect 438 1757 498 1791
rect 662 1847 927 1867
rect 662 1846 725 1847
rect 759 1846 797 1847
rect 831 1846 927 1847
rect 662 1812 676 1846
rect 710 1813 725 1846
rect 778 1813 797 1846
rect 710 1812 744 1813
rect 778 1812 812 1813
rect 846 1812 880 1846
rect 914 1812 927 1846
rect 662 1785 927 1812
rect 1093 1803 1233 1924
rect 358 1731 498 1757
rect 1093 1769 1146 1803
rect 1180 1791 1233 1803
rect 1093 1757 1156 1769
rect 1190 1757 1233 1791
rect 358 1697 395 1731
rect 429 1723 498 1731
rect 358 1689 404 1697
rect 438 1689 498 1723
rect 358 1659 498 1689
rect 358 1625 395 1659
rect 429 1655 498 1659
rect 358 1621 404 1625
rect 438 1621 498 1655
rect 358 1587 498 1621
rect 358 1553 395 1587
rect 438 1553 498 1587
rect 358 1519 498 1553
rect 358 1515 404 1519
rect 358 1481 395 1515
rect 438 1485 498 1519
rect 429 1481 498 1485
rect 358 1451 498 1481
rect 358 1443 404 1451
rect 358 1409 395 1443
rect 438 1417 498 1451
rect 429 1409 498 1417
rect 358 1383 498 1409
rect 358 1371 404 1383
rect 358 1337 395 1371
rect 438 1349 498 1383
rect 429 1337 498 1349
rect 358 1315 498 1337
rect 358 1299 404 1315
rect 358 1265 395 1299
rect 438 1281 498 1315
rect 429 1265 498 1281
rect 358 1247 498 1265
rect 358 1227 404 1247
rect 358 1193 395 1227
rect 438 1213 498 1247
rect 429 1193 498 1213
rect 358 1179 498 1193
rect 358 1155 404 1179
rect 358 1121 395 1155
rect 438 1145 498 1179
rect 429 1121 498 1145
rect 358 1111 498 1121
rect 358 1083 404 1111
rect 358 1049 395 1083
rect 438 1077 498 1111
rect 429 1049 498 1077
rect 358 1043 498 1049
rect 358 1011 404 1043
rect 358 977 395 1011
rect 438 1009 498 1043
rect 429 977 498 1009
rect 358 975 498 977
rect 358 941 404 975
rect 438 941 498 975
rect 358 939 498 941
rect 358 905 395 939
rect 429 907 498 939
rect 358 873 404 905
rect 438 873 498 907
rect 358 867 498 873
rect 358 833 395 867
rect 429 839 498 867
rect 358 805 404 833
rect 438 805 498 839
rect 358 795 498 805
rect 358 761 395 795
rect 429 771 498 795
rect 358 737 404 761
rect 438 737 498 771
rect 358 723 498 737
rect 358 689 395 723
rect 429 703 498 723
rect 358 669 404 689
rect 438 669 498 703
rect 593 1635 701 1751
rect 593 1601 602 1635
rect 636 1601 701 1635
rect 593 1583 701 1601
rect 593 1567 621 1583
rect 593 1533 602 1567
rect 655 1549 701 1583
rect 636 1533 701 1549
rect 593 1511 701 1533
rect 593 1499 621 1511
rect 593 1465 602 1499
rect 655 1477 701 1511
rect 636 1465 701 1477
rect 593 1439 701 1465
rect 593 1431 621 1439
rect 593 1397 602 1431
rect 655 1405 701 1439
rect 636 1397 701 1405
rect 593 1367 701 1397
rect 593 1363 621 1367
rect 593 1329 602 1363
rect 655 1333 701 1367
rect 636 1329 701 1333
rect 593 1295 701 1329
rect 593 1261 602 1295
rect 655 1261 701 1295
rect 593 1227 701 1261
rect 593 1193 602 1227
rect 636 1223 701 1227
rect 593 1189 621 1193
rect 655 1189 701 1223
rect 593 1159 701 1189
rect 593 1125 602 1159
rect 636 1151 701 1159
rect 593 1117 621 1125
rect 655 1117 701 1151
rect 593 1091 701 1117
rect 593 1057 602 1091
rect 636 1079 701 1091
rect 593 1045 621 1057
rect 655 1045 701 1079
rect 593 1023 701 1045
rect 593 989 602 1023
rect 636 1007 701 1023
rect 593 973 621 989
rect 655 973 701 1007
rect 593 955 701 973
rect 593 921 602 955
rect 636 935 701 955
rect 593 901 621 921
rect 655 901 701 935
rect 593 887 701 901
rect 593 853 602 887
rect 636 863 701 887
rect 593 829 621 853
rect 655 829 701 863
rect 593 819 701 829
rect 593 785 602 819
rect 636 791 701 819
rect 593 757 621 785
rect 655 757 701 791
rect 593 751 701 757
rect 593 717 602 751
rect 636 717 701 751
rect 593 672 701 717
rect 888 1635 996 1751
rect 888 1601 946 1635
rect 980 1601 996 1635
rect 888 1583 996 1601
rect 888 1549 915 1583
rect 949 1567 996 1583
rect 888 1533 946 1549
rect 980 1533 996 1567
rect 888 1511 996 1533
rect 888 1477 915 1511
rect 949 1499 996 1511
rect 888 1465 946 1477
rect 980 1465 996 1499
rect 888 1439 996 1465
rect 888 1405 915 1439
rect 949 1431 996 1439
rect 888 1397 946 1405
rect 980 1397 996 1431
rect 888 1367 996 1397
rect 888 1333 915 1367
rect 949 1363 996 1367
rect 888 1329 946 1333
rect 980 1329 996 1363
rect 888 1295 996 1329
rect 888 1261 915 1295
rect 980 1261 996 1295
rect 888 1227 996 1261
rect 888 1223 946 1227
rect 888 1189 915 1223
rect 980 1193 996 1227
rect 949 1189 996 1193
rect 888 1159 996 1189
rect 888 1151 946 1159
rect 888 1117 915 1151
rect 980 1125 996 1159
rect 949 1117 996 1125
rect 888 1091 996 1117
rect 888 1079 946 1091
rect 888 1045 915 1079
rect 980 1057 996 1091
rect 949 1045 996 1057
rect 888 1023 996 1045
rect 888 1007 946 1023
rect 888 973 915 1007
rect 980 989 996 1023
rect 949 973 996 989
rect 888 955 996 973
rect 888 935 946 955
rect 888 901 915 935
rect 980 921 996 955
rect 949 901 996 921
rect 888 887 996 901
rect 888 863 946 887
rect 888 829 915 863
rect 980 853 996 887
rect 949 829 996 853
rect 888 819 996 829
rect 888 791 946 819
rect 888 757 915 791
rect 980 785 996 819
rect 949 757 996 785
rect 888 751 996 757
rect 888 717 946 751
rect 980 717 996 751
rect 888 672 996 717
rect 1093 1731 1233 1757
rect 1093 1697 1146 1731
rect 1180 1723 1233 1731
rect 1093 1689 1156 1697
rect 1190 1689 1233 1723
rect 1093 1659 1233 1689
rect 1093 1625 1146 1659
rect 1180 1655 1233 1659
rect 1093 1621 1156 1625
rect 1190 1621 1233 1655
rect 1093 1587 1233 1621
rect 1093 1553 1146 1587
rect 1190 1553 1233 1587
rect 1093 1519 1233 1553
rect 1093 1515 1156 1519
rect 1093 1481 1146 1515
rect 1190 1485 1233 1519
rect 1180 1481 1233 1485
rect 1093 1451 1233 1481
rect 1093 1443 1156 1451
rect 1093 1409 1146 1443
rect 1190 1417 1233 1451
rect 1180 1409 1233 1417
rect 1093 1383 1233 1409
rect 1093 1371 1156 1383
rect 1093 1337 1146 1371
rect 1190 1349 1233 1383
rect 1180 1337 1233 1349
rect 1093 1315 1233 1337
rect 1093 1299 1156 1315
rect 1093 1265 1146 1299
rect 1190 1281 1233 1315
rect 1180 1265 1233 1281
rect 1093 1247 1233 1265
rect 1093 1227 1156 1247
rect 1093 1193 1146 1227
rect 1190 1213 1233 1247
rect 1180 1193 1233 1213
rect 1093 1179 1233 1193
rect 1093 1155 1156 1179
rect 1093 1121 1146 1155
rect 1190 1145 1233 1179
rect 1180 1121 1233 1145
rect 1093 1111 1233 1121
rect 1093 1083 1156 1111
rect 1093 1049 1146 1083
rect 1190 1077 1233 1111
rect 1180 1049 1233 1077
rect 1093 1043 1233 1049
rect 1093 1011 1156 1043
rect 1093 977 1146 1011
rect 1190 1009 1233 1043
rect 1180 977 1233 1009
rect 1093 975 1233 977
rect 1093 941 1156 975
rect 1190 941 1233 975
rect 1093 939 1233 941
rect 1093 905 1146 939
rect 1180 907 1233 939
rect 1093 873 1156 905
rect 1190 873 1233 907
rect 1093 867 1233 873
rect 1093 833 1146 867
rect 1180 839 1233 867
rect 1093 805 1156 833
rect 1190 805 1233 839
rect 1093 795 1233 805
rect 1093 761 1146 795
rect 1180 771 1233 795
rect 1093 737 1156 761
rect 1190 737 1233 771
rect 1093 723 1233 737
rect 1093 689 1146 723
rect 1180 703 1233 723
rect 358 651 498 669
rect 358 617 395 651
rect 429 635 498 651
rect 358 601 404 617
rect 438 601 498 635
rect 358 579 498 601
rect 358 545 395 579
rect 429 567 498 579
rect 358 533 404 545
rect 438 533 498 567
rect 358 507 498 533
rect 358 473 395 507
rect 429 498 498 507
rect 1093 669 1156 689
rect 1190 669 1233 703
rect 1093 651 1233 669
rect 1093 617 1146 651
rect 1180 635 1233 651
rect 1093 601 1156 617
rect 1190 601 1233 635
rect 1093 579 1233 601
rect 1093 545 1146 579
rect 1180 567 1233 579
rect 1093 533 1156 545
rect 1190 533 1233 567
rect 1093 507 1233 533
rect 1093 498 1146 507
rect 429 473 1146 498
rect 1180 473 1233 507
rect 358 445 1233 473
rect 358 435 473 445
rect 358 401 395 435
rect 429 411 473 435
rect 507 411 541 445
rect 575 411 609 445
rect 643 411 677 445
rect 711 411 745 445
rect 779 411 813 445
rect 847 411 881 445
rect 915 411 949 445
rect 983 411 1017 445
rect 1051 411 1085 445
rect 1119 435 1233 445
rect 1119 411 1146 435
rect 429 401 1146 411
rect 1180 401 1233 435
rect 358 358 1233 401
rect 1385 2058 1438 2092
rect 1472 2058 1525 2092
rect 1385 2035 1525 2058
rect 1385 1990 1438 2035
rect 1472 1990 1525 2035
rect 1385 1963 1525 1990
rect 1385 1922 1438 1963
rect 1472 1922 1525 1963
rect 1385 1891 1525 1922
rect 1385 1854 1438 1891
rect 1472 1854 1525 1891
rect 1385 1820 1525 1854
rect 1385 1785 1438 1820
rect 1472 1785 1525 1820
rect 1385 1752 1525 1785
rect 1385 1713 1438 1752
rect 1472 1713 1525 1752
rect 1385 1684 1525 1713
rect 1385 1641 1438 1684
rect 1472 1641 1525 1684
rect 1385 1616 1525 1641
rect 1385 1569 1438 1616
rect 1472 1569 1525 1616
rect 1385 1548 1525 1569
rect 1385 1497 1438 1548
rect 1472 1497 1525 1548
rect 1385 1480 1525 1497
rect 1385 1425 1438 1480
rect 1472 1425 1525 1480
rect 1385 1412 1525 1425
rect 1385 1353 1438 1412
rect 1472 1353 1525 1412
rect 1385 1344 1525 1353
rect 1385 1281 1438 1344
rect 1472 1281 1525 1344
rect 1385 1276 1525 1281
rect 1385 1209 1438 1276
rect 1472 1209 1525 1276
rect 1385 1208 1525 1209
rect 1385 1174 1438 1208
rect 1472 1174 1525 1208
rect 1385 1171 1525 1174
rect 1385 1106 1438 1171
rect 1472 1106 1525 1171
rect 1385 1099 1525 1106
rect 1385 1038 1438 1099
rect 1472 1038 1525 1099
rect 1385 1027 1525 1038
rect 1385 970 1438 1027
rect 1472 970 1525 1027
rect 1385 955 1525 970
rect 1385 902 1438 955
rect 1472 902 1525 955
rect 1385 883 1525 902
rect 1385 834 1438 883
rect 1472 834 1525 883
rect 1385 811 1525 834
rect 1385 766 1438 811
rect 1472 766 1525 811
rect 1385 739 1525 766
rect 1385 698 1438 739
rect 1472 698 1525 739
rect 1385 667 1525 698
rect 1385 630 1438 667
rect 1472 630 1525 667
rect 1385 596 1525 630
rect 1385 561 1438 596
rect 1472 561 1525 596
rect 1385 528 1525 561
rect 1385 489 1438 528
rect 1472 489 1525 528
rect 1385 460 1525 489
rect 1385 417 1438 460
rect 1472 417 1525 460
rect 1385 392 1525 417
rect 66 324 206 345
rect 66 273 119 324
rect 153 273 206 324
rect 66 256 206 273
rect 66 222 119 256
rect 153 222 206 256
rect 66 206 206 222
rect 1385 345 1438 392
rect 1472 345 1525 392
rect 1385 324 1525 345
rect 1385 273 1438 324
rect 1472 273 1525 324
rect 1385 256 1525 273
rect 1385 222 1438 256
rect 1472 222 1525 256
rect 1385 206 1525 222
rect 66 153 1525 206
rect 66 119 303 153
rect 337 119 371 153
rect 405 119 439 153
rect 473 119 507 153
rect 541 119 575 153
rect 609 119 643 153
rect 677 119 711 153
rect 745 119 779 153
rect 813 119 847 153
rect 881 119 915 153
rect 949 119 983 153
rect 1017 119 1051 153
rect 1085 142 1119 153
rect 1085 119 1118 142
rect 1153 119 1187 153
rect 1221 142 1255 153
rect 1289 142 1525 153
rect 1224 119 1255 142
rect 66 108 1118 119
rect 1152 108 1190 119
rect 1224 108 1262 119
rect 1296 108 1525 142
rect 66 66 1525 108
<< viali >>
rect 307 2271 337 2305
rect 337 2271 341 2305
rect 379 2271 405 2305
rect 405 2271 413 2305
rect 451 2271 473 2305
rect 473 2271 485 2305
rect 523 2271 541 2305
rect 541 2271 557 2305
rect 595 2271 609 2305
rect 609 2271 629 2305
rect 959 2271 983 2305
rect 983 2271 993 2305
rect 1031 2271 1051 2305
rect 1051 2271 1065 2305
rect 1103 2271 1119 2305
rect 1119 2271 1137 2305
rect 1175 2271 1187 2305
rect 1187 2271 1209 2305
rect 1247 2271 1255 2305
rect 1255 2271 1281 2305
rect 119 2024 153 2035
rect 119 2001 153 2024
rect 119 1956 153 1963
rect 119 1929 153 1956
rect 119 1888 153 1891
rect 119 1857 153 1888
rect 119 1786 153 1819
rect 119 1785 153 1786
rect 119 1718 153 1747
rect 119 1713 153 1718
rect 119 1650 153 1675
rect 119 1641 153 1650
rect 119 1582 153 1603
rect 119 1569 153 1582
rect 119 1514 153 1531
rect 119 1497 153 1514
rect 119 1446 153 1459
rect 119 1425 153 1446
rect 119 1378 153 1387
rect 119 1353 153 1378
rect 119 1310 153 1315
rect 119 1281 153 1310
rect 119 1242 153 1243
rect 119 1209 153 1242
rect 119 1140 153 1171
rect 119 1137 153 1140
rect 119 1072 153 1099
rect 119 1065 153 1072
rect 119 1004 153 1027
rect 119 993 153 1004
rect 119 936 153 955
rect 119 921 153 936
rect 119 868 153 883
rect 119 849 153 868
rect 119 800 153 811
rect 119 777 153 800
rect 119 732 153 739
rect 119 705 153 732
rect 119 664 153 667
rect 119 633 153 664
rect 119 562 153 595
rect 119 561 153 562
rect 119 494 153 523
rect 119 489 153 494
rect 119 426 153 451
rect 119 417 153 426
rect 119 358 153 379
rect 119 345 153 358
rect 454 1979 473 2003
rect 473 1979 488 2003
rect 526 1979 541 2003
rect 541 1979 560 2003
rect 598 1979 609 2003
rect 609 1979 632 2003
rect 928 1979 949 2003
rect 949 1979 962 2003
rect 1000 1979 1017 2003
rect 1017 1979 1034 2003
rect 1072 1979 1085 2003
rect 1085 1979 1106 2003
rect 454 1969 488 1979
rect 526 1969 560 1979
rect 598 1969 632 1979
rect 928 1969 962 1979
rect 1000 1969 1034 1979
rect 1072 1969 1106 1979
rect 395 1791 429 1803
rect 395 1769 404 1791
rect 404 1769 429 1791
rect 725 1846 759 1847
rect 797 1846 831 1847
rect 725 1813 744 1846
rect 744 1813 759 1846
rect 797 1813 812 1846
rect 812 1813 831 1846
rect 1146 1791 1180 1803
rect 1146 1769 1156 1791
rect 1156 1769 1180 1791
rect 395 1723 429 1731
rect 395 1697 404 1723
rect 404 1697 429 1723
rect 395 1655 429 1659
rect 395 1625 404 1655
rect 404 1625 429 1655
rect 395 1553 404 1587
rect 404 1553 429 1587
rect 395 1485 404 1515
rect 404 1485 429 1515
rect 395 1481 429 1485
rect 395 1417 404 1443
rect 404 1417 429 1443
rect 395 1409 429 1417
rect 395 1349 404 1371
rect 404 1349 429 1371
rect 395 1337 429 1349
rect 395 1281 404 1299
rect 404 1281 429 1299
rect 395 1265 429 1281
rect 395 1213 404 1227
rect 404 1213 429 1227
rect 395 1193 429 1213
rect 395 1145 404 1155
rect 404 1145 429 1155
rect 395 1121 429 1145
rect 395 1077 404 1083
rect 404 1077 429 1083
rect 395 1049 429 1077
rect 395 1009 404 1011
rect 404 1009 429 1011
rect 395 977 429 1009
rect 395 907 429 939
rect 395 905 404 907
rect 404 905 429 907
rect 395 839 429 867
rect 395 833 404 839
rect 404 833 429 839
rect 395 771 429 795
rect 395 761 404 771
rect 404 761 429 771
rect 395 703 429 723
rect 395 689 404 703
rect 404 689 429 703
rect 621 1567 655 1583
rect 621 1549 636 1567
rect 636 1549 655 1567
rect 621 1499 655 1511
rect 621 1477 636 1499
rect 636 1477 655 1499
rect 621 1431 655 1439
rect 621 1405 636 1431
rect 636 1405 655 1431
rect 621 1363 655 1367
rect 621 1333 636 1363
rect 636 1333 655 1363
rect 621 1261 636 1295
rect 636 1261 655 1295
rect 621 1193 636 1223
rect 636 1193 655 1223
rect 621 1189 655 1193
rect 621 1125 636 1151
rect 636 1125 655 1151
rect 621 1117 655 1125
rect 621 1057 636 1079
rect 636 1057 655 1079
rect 621 1045 655 1057
rect 621 989 636 1007
rect 636 989 655 1007
rect 621 973 655 989
rect 621 921 636 935
rect 636 921 655 935
rect 621 901 655 921
rect 621 853 636 863
rect 636 853 655 863
rect 621 829 655 853
rect 621 785 636 791
rect 636 785 655 791
rect 621 757 655 785
rect 915 1567 949 1583
rect 915 1549 946 1567
rect 946 1549 949 1567
rect 915 1499 949 1511
rect 915 1477 946 1499
rect 946 1477 949 1499
rect 915 1431 949 1439
rect 915 1405 946 1431
rect 946 1405 949 1431
rect 915 1363 949 1367
rect 915 1333 946 1363
rect 946 1333 949 1363
rect 915 1261 946 1295
rect 946 1261 949 1295
rect 915 1193 946 1223
rect 946 1193 949 1223
rect 915 1189 949 1193
rect 915 1125 946 1151
rect 946 1125 949 1151
rect 915 1117 949 1125
rect 915 1057 946 1079
rect 946 1057 949 1079
rect 915 1045 949 1057
rect 915 989 946 1007
rect 946 989 949 1007
rect 915 973 949 989
rect 915 921 946 935
rect 946 921 949 935
rect 915 901 949 921
rect 915 853 946 863
rect 946 853 949 863
rect 915 829 949 853
rect 915 785 946 791
rect 946 785 949 791
rect 915 757 949 785
rect 1146 1723 1180 1731
rect 1146 1697 1156 1723
rect 1156 1697 1180 1723
rect 1146 1655 1180 1659
rect 1146 1625 1156 1655
rect 1156 1625 1180 1655
rect 1146 1553 1156 1587
rect 1156 1553 1180 1587
rect 1146 1485 1156 1515
rect 1156 1485 1180 1515
rect 1146 1481 1180 1485
rect 1146 1417 1156 1443
rect 1156 1417 1180 1443
rect 1146 1409 1180 1417
rect 1146 1349 1156 1371
rect 1156 1349 1180 1371
rect 1146 1337 1180 1349
rect 1146 1281 1156 1299
rect 1156 1281 1180 1299
rect 1146 1265 1180 1281
rect 1146 1213 1156 1227
rect 1156 1213 1180 1227
rect 1146 1193 1180 1213
rect 1146 1145 1156 1155
rect 1156 1145 1180 1155
rect 1146 1121 1180 1145
rect 1146 1077 1156 1083
rect 1156 1077 1180 1083
rect 1146 1049 1180 1077
rect 1146 1009 1156 1011
rect 1156 1009 1180 1011
rect 1146 977 1180 1009
rect 1146 907 1180 939
rect 1146 905 1156 907
rect 1156 905 1180 907
rect 1146 839 1180 867
rect 1146 833 1156 839
rect 1156 833 1180 839
rect 1146 771 1180 795
rect 1146 761 1156 771
rect 1156 761 1180 771
rect 1146 703 1180 723
rect 1146 689 1156 703
rect 1156 689 1180 703
rect 395 635 429 651
rect 395 617 404 635
rect 404 617 429 635
rect 395 567 429 579
rect 395 545 404 567
rect 404 545 429 567
rect 395 473 429 507
rect 1146 635 1180 651
rect 1146 617 1156 635
rect 1156 617 1180 635
rect 1146 567 1180 579
rect 1146 545 1156 567
rect 1156 545 1180 567
rect 1146 473 1180 507
rect 395 401 429 435
rect 1146 401 1180 435
rect 1438 2024 1472 2035
rect 1438 2001 1472 2024
rect 1438 1956 1472 1963
rect 1438 1929 1472 1956
rect 1438 1888 1472 1891
rect 1438 1857 1472 1888
rect 1438 1786 1472 1819
rect 1438 1785 1472 1786
rect 1438 1718 1472 1747
rect 1438 1713 1472 1718
rect 1438 1650 1472 1675
rect 1438 1641 1472 1650
rect 1438 1582 1472 1603
rect 1438 1569 1472 1582
rect 1438 1514 1472 1531
rect 1438 1497 1472 1514
rect 1438 1446 1472 1459
rect 1438 1425 1472 1446
rect 1438 1378 1472 1387
rect 1438 1353 1472 1378
rect 1438 1310 1472 1315
rect 1438 1281 1472 1310
rect 1438 1242 1472 1243
rect 1438 1209 1472 1242
rect 1438 1140 1472 1171
rect 1438 1137 1472 1140
rect 1438 1072 1472 1099
rect 1438 1065 1472 1072
rect 1438 1004 1472 1027
rect 1438 993 1472 1004
rect 1438 936 1472 955
rect 1438 921 1472 936
rect 1438 868 1472 883
rect 1438 849 1472 868
rect 1438 800 1472 811
rect 1438 777 1472 800
rect 1438 732 1472 739
rect 1438 705 1472 732
rect 1438 664 1472 667
rect 1438 633 1472 664
rect 1438 562 1472 595
rect 1438 561 1472 562
rect 1438 494 1472 523
rect 1438 489 1472 494
rect 1438 426 1472 451
rect 1438 417 1472 426
rect 119 290 153 307
rect 119 273 153 290
rect 1438 358 1472 379
rect 1438 345 1472 358
rect 1438 290 1472 307
rect 1438 273 1472 290
rect 1118 119 1119 142
rect 1119 119 1152 142
rect 1190 119 1221 142
rect 1221 119 1224 142
rect 1262 119 1289 142
rect 1289 119 1296 142
rect 1118 108 1152 119
rect 1190 108 1224 119
rect 1262 108 1296 119
<< metal1 >>
tri 155 2305 208 2358 se
rect 208 2305 669 2358
tri 121 2271 155 2305 se
rect 155 2271 307 2305
rect 341 2271 379 2305
rect 413 2271 451 2305
rect 485 2271 523 2305
rect 557 2271 595 2305
rect 629 2271 669 2305
tri 66 2216 121 2271 se
rect 121 2218 669 2271
rect 121 2216 286 2218
tri 286 2216 288 2218 nw
rect 66 2035 206 2216
tri 206 2136 286 2216 nw
tri 393 2035 424 2066 se
rect 424 2035 669 2066
rect 66 2001 119 2035
rect 153 2001 206 2035
tri 361 2003 393 2035 se
rect 393 2003 669 2035
rect 66 1963 206 2001
rect 66 1929 119 1963
rect 153 1929 206 1963
rect 66 1891 206 1929
rect 66 1857 119 1891
rect 153 1857 206 1891
rect 66 1819 206 1857
rect 66 1785 119 1819
rect 153 1785 206 1819
rect 66 1747 206 1785
rect 66 1713 119 1747
rect 153 1713 206 1747
rect 66 1675 206 1713
rect 66 1641 119 1675
rect 153 1641 206 1675
rect 66 1603 206 1641
rect 66 1569 119 1603
rect 153 1569 206 1603
rect 66 1531 206 1569
rect 66 1497 119 1531
rect 153 1497 206 1531
rect 66 1459 206 1497
rect 66 1425 119 1459
rect 153 1425 206 1459
rect 66 1387 206 1425
rect 66 1353 119 1387
rect 153 1353 206 1387
rect 66 1315 206 1353
rect 66 1281 119 1315
rect 153 1281 206 1315
rect 66 1243 206 1281
rect 66 1209 119 1243
rect 153 1209 206 1243
rect 66 1171 206 1209
rect 66 1137 119 1171
rect 153 1137 206 1171
rect 66 1099 206 1137
rect 66 1065 119 1099
rect 153 1065 206 1099
rect 66 1027 206 1065
rect 66 993 119 1027
rect 153 993 206 1027
rect 66 955 206 993
rect 66 921 119 955
rect 153 921 206 955
rect 66 883 206 921
rect 66 849 119 883
rect 153 849 206 883
rect 66 811 206 849
rect 66 777 119 811
rect 153 777 206 811
rect 66 739 206 777
rect 66 705 119 739
rect 153 705 206 739
rect 66 667 206 705
rect 66 633 119 667
rect 153 633 206 667
rect 66 595 206 633
rect 66 561 119 595
rect 153 561 206 595
rect 66 523 206 561
rect 66 489 119 523
rect 153 489 206 523
rect 66 451 206 489
rect 66 417 119 451
rect 153 417 206 451
rect 66 379 206 417
rect 66 345 119 379
rect 153 345 206 379
rect 66 307 206 345
rect 66 273 119 307
rect 153 273 206 307
rect 66 69 206 273
rect 66 66 203 69
rect 204 67 205 68
tri 358 2000 361 2003 se
rect 361 2000 454 2003
rect 358 1969 454 2000
rect 488 1969 526 2003
rect 560 1969 598 2003
rect 632 1969 669 2003
rect 358 1901 669 1969
rect 358 1891 601 1901
tri 601 1891 611 1901 nw
rect 358 1857 567 1891
tri 567 1857 601 1891 nw
rect 358 1847 557 1857
tri 557 1847 567 1857 nw
rect 703 1847 852 2359
rect 886 2305 1383 2358
rect 886 2271 959 2305
rect 993 2271 1031 2305
rect 1065 2271 1103 2305
rect 1137 2271 1175 2305
rect 1209 2271 1247 2305
rect 1281 2271 1383 2305
rect 886 2218 1383 2271
tri 1289 2216 1291 2218 ne
rect 1291 2216 1383 2218
tri 1383 2216 1525 2358 sw
tri 1291 2124 1383 2216 ne
rect 1383 2124 1525 2216
tri 1383 2122 1385 2124 ne
rect 886 2035 1167 2066
tri 1167 2035 1198 2066 sw
rect 1385 2035 1525 2124
rect 886 2003 1198 2035
rect 886 1969 928 2003
rect 962 1969 1000 2003
rect 1034 1969 1072 2003
rect 1106 2001 1198 2003
tri 1198 2001 1232 2035 sw
rect 1385 2001 1438 2035
rect 1472 2001 1525 2035
rect 1106 2000 1232 2001
tri 1232 2000 1233 2001 sw
rect 1106 1969 1233 2000
rect 886 1901 1233 1969
tri 1012 1891 1022 1901 ne
rect 1022 1891 1233 1901
tri 1022 1857 1056 1891 ne
rect 1056 1857 1233 1891
rect 358 1803 536 1847
tri 536 1826 557 1847 nw
rect 358 1769 395 1803
rect 429 1769 536 1803
rect 703 1813 725 1847
rect 759 1813 797 1847
rect 831 1813 852 1847
tri 1056 1820 1093 1857 ne
rect 703 1791 852 1813
rect 1093 1803 1233 1857
rect 358 1731 536 1769
rect 1093 1769 1146 1803
rect 1180 1769 1233 1803
rect 358 1697 395 1731
rect 429 1697 536 1731
rect 358 1659 536 1697
rect 358 1625 395 1659
rect 429 1625 536 1659
rect 358 1587 536 1625
rect 358 1553 395 1587
rect 429 1553 536 1587
rect 358 1515 536 1553
rect 358 1481 395 1515
rect 429 1481 536 1515
rect 358 1443 536 1481
rect 358 1409 395 1443
rect 429 1409 536 1443
rect 358 1371 536 1409
rect 358 1337 395 1371
rect 429 1337 536 1371
rect 358 1299 536 1337
rect 358 1265 395 1299
rect 429 1265 536 1299
rect 358 1227 536 1265
rect 358 1193 395 1227
rect 429 1193 536 1227
rect 358 1155 536 1193
rect 358 1121 395 1155
rect 429 1121 536 1155
rect 358 1083 536 1121
rect 358 1049 395 1083
rect 429 1049 536 1083
rect 358 1011 536 1049
rect 358 977 395 1011
rect 429 977 536 1011
rect 358 939 536 977
rect 358 905 395 939
rect 429 905 536 939
rect 358 867 536 905
rect 358 833 395 867
rect 429 833 536 867
rect 358 795 536 833
rect 358 761 395 795
rect 429 761 536 795
rect 358 723 536 761
rect 358 689 395 723
rect 429 689 536 723
rect 358 651 536 689
rect 358 617 395 651
rect 429 617 536 651
rect 358 579 536 617
rect 358 545 395 579
rect 429 545 536 579
rect 358 507 536 545
rect 358 473 395 507
rect 429 473 536 507
rect 358 435 536 473
rect 358 401 395 435
rect 429 401 536 435
rect 358 69 536 401
rect 358 66 533 69
rect 534 67 535 68
rect 572 1583 772 1709
rect 572 1549 621 1583
rect 655 1549 772 1583
rect 572 1511 772 1549
rect 572 1477 621 1511
rect 655 1477 772 1511
rect 572 1439 772 1477
rect 572 1405 621 1439
rect 655 1405 772 1439
rect 572 1367 772 1405
rect 572 1333 621 1367
rect 655 1333 772 1367
rect 572 1295 772 1333
rect 572 1261 621 1295
rect 655 1261 772 1295
rect 572 1223 772 1261
rect 572 1189 621 1223
rect 655 1189 772 1223
rect 572 1151 772 1189
rect 572 1117 621 1151
rect 655 1117 772 1151
rect 572 1079 772 1117
rect 572 1045 621 1079
rect 655 1045 772 1079
rect 572 1007 772 1045
rect 572 973 621 1007
rect 655 973 772 1007
rect 572 935 772 973
rect 572 901 621 935
rect 655 901 772 935
rect 572 863 772 901
rect 572 829 621 863
rect 655 829 772 863
rect 572 791 772 829
rect 572 757 621 791
rect 655 757 772 791
rect 572 66 772 757
rect 831 1583 1031 1752
rect 831 1549 915 1583
rect 949 1549 1031 1583
rect 831 1511 1031 1549
rect 831 1477 915 1511
rect 949 1477 1031 1511
rect 831 1439 1031 1477
rect 831 1405 915 1439
rect 949 1405 1031 1439
rect 831 1367 1031 1405
rect 831 1333 915 1367
rect 949 1333 1031 1367
rect 831 1295 1031 1333
rect 831 1261 915 1295
rect 949 1261 1031 1295
rect 831 1223 1031 1261
rect 831 1189 915 1223
rect 949 1189 1031 1223
rect 831 1151 1031 1189
rect 831 1117 915 1151
rect 949 1117 1031 1151
rect 831 1079 1031 1117
rect 831 1045 915 1079
rect 949 1045 1031 1079
rect 831 1007 1031 1045
rect 831 973 915 1007
rect 949 973 1031 1007
rect 831 935 1031 973
rect 831 901 915 935
rect 949 901 1031 935
rect 831 863 1031 901
rect 831 829 915 863
rect 949 829 1031 863
rect 831 791 1031 829
rect 831 757 915 791
rect 949 757 1031 791
rect 831 66 1031 757
rect 1093 1731 1233 1769
rect 1093 1697 1146 1731
rect 1180 1697 1233 1731
rect 1093 1659 1233 1697
rect 1093 1625 1146 1659
rect 1180 1625 1233 1659
rect 1093 1587 1233 1625
rect 1093 1553 1146 1587
rect 1180 1553 1233 1587
rect 1093 1515 1233 1553
rect 1093 1481 1146 1515
rect 1180 1481 1233 1515
rect 1093 1443 1233 1481
rect 1093 1409 1146 1443
rect 1180 1409 1233 1443
rect 1093 1371 1233 1409
rect 1093 1337 1146 1371
rect 1180 1337 1233 1371
rect 1093 1299 1233 1337
rect 1093 1265 1146 1299
rect 1180 1265 1233 1299
rect 1093 1227 1233 1265
rect 1093 1193 1146 1227
rect 1180 1193 1233 1227
rect 1093 1155 1233 1193
rect 1093 1121 1146 1155
rect 1180 1121 1233 1155
rect 1093 1083 1233 1121
rect 1093 1049 1146 1083
rect 1180 1049 1233 1083
rect 1093 1011 1233 1049
rect 1093 977 1146 1011
rect 1180 977 1233 1011
rect 1093 939 1233 977
rect 1093 905 1146 939
rect 1180 905 1233 939
rect 1093 867 1233 905
rect 1093 833 1146 867
rect 1180 833 1233 867
rect 1093 795 1233 833
rect 1093 761 1146 795
rect 1180 761 1233 795
rect 1093 723 1233 761
rect 1093 689 1146 723
rect 1180 689 1233 723
rect 1093 651 1233 689
rect 1093 617 1146 651
rect 1180 617 1233 651
rect 1093 579 1233 617
rect 1093 545 1146 579
rect 1180 545 1233 579
rect 1093 507 1233 545
rect 1093 473 1146 507
rect 1180 473 1233 507
rect 1093 435 1233 473
rect 1093 401 1146 435
rect 1180 401 1233 435
rect 1093 358 1233 401
rect 1385 1963 1525 2001
rect 1385 1929 1438 1963
rect 1472 1929 1525 1963
rect 1385 1891 1525 1929
rect 1385 1857 1438 1891
rect 1472 1857 1525 1891
rect 1385 1819 1525 1857
rect 1385 1785 1438 1819
rect 1472 1785 1525 1819
rect 1385 1747 1525 1785
rect 1385 1713 1438 1747
rect 1472 1713 1525 1747
rect 1385 1675 1525 1713
rect 1385 1641 1438 1675
rect 1472 1641 1525 1675
rect 1385 1603 1525 1641
rect 1385 1569 1438 1603
rect 1472 1569 1525 1603
rect 1385 1531 1525 1569
rect 1385 1497 1438 1531
rect 1472 1497 1525 1531
rect 1385 1459 1525 1497
rect 1385 1425 1438 1459
rect 1472 1425 1525 1459
rect 1385 1387 1525 1425
rect 1385 1353 1438 1387
rect 1472 1353 1525 1387
rect 1385 1315 1525 1353
rect 1385 1281 1438 1315
rect 1472 1281 1525 1315
rect 1385 1243 1525 1281
rect 1385 1209 1438 1243
rect 1472 1209 1525 1243
rect 1385 1171 1525 1209
rect 1385 1137 1438 1171
rect 1472 1137 1525 1171
rect 1385 1099 1525 1137
rect 1385 1065 1438 1099
rect 1472 1065 1525 1099
rect 1385 1027 1525 1065
rect 1385 993 1438 1027
rect 1472 993 1525 1027
rect 1385 955 1525 993
rect 1385 921 1438 955
rect 1472 921 1525 955
rect 1385 883 1525 921
rect 1385 849 1438 883
rect 1472 849 1525 883
rect 1385 811 1525 849
rect 1385 777 1438 811
rect 1472 777 1525 811
rect 1385 739 1525 777
rect 1385 705 1438 739
rect 1472 705 1525 739
rect 1385 667 1525 705
rect 1385 633 1438 667
rect 1472 633 1525 667
rect 1385 595 1525 633
rect 1385 561 1438 595
rect 1472 561 1525 595
rect 1385 523 1525 561
rect 1385 489 1438 523
rect 1472 489 1525 523
rect 1385 451 1525 489
rect 1385 417 1438 451
rect 1472 417 1525 451
rect 1385 379 1525 417
rect 1385 345 1438 379
rect 1472 345 1525 379
rect 1385 307 1525 345
tri 1356 273 1385 302 se
rect 1385 273 1438 307
rect 1472 273 1525 307
tri 1289 206 1356 273 se
rect 1356 208 1525 273
rect 1356 206 1523 208
tri 1523 206 1525 208 nw
rect 1070 142 1383 206
rect 1070 108 1118 142
rect 1152 108 1190 142
rect 1224 108 1262 142
rect 1296 108 1383 142
rect 1070 66 1383 108
tri 1383 66 1523 206 nw
<< rmetal1 >>
rect 203 68 206 69
rect 203 67 204 68
rect 205 67 206 68
rect 203 66 206 67
rect 533 68 536 69
rect 533 67 534 68
rect 535 67 536 68
rect 533 66 536 67
use sky130_fd_pr__dfl1__example_55959141808158  sky130_fd_pr__dfl1__example_55959141808158_0
timestamp 1707688321
transform 1 0 938 0 1 705
box 0 0 1 1
use sky130_fd_pr__dfl1__example_55959141808158  sky130_fd_pr__dfl1__example_55959141808158_1
timestamp 1707688321
transform 1 0 594 0 1 705
box 0 0 1 1
use sky130_fd_pr__tpl1__example_55959141808148  sky130_fd_pr__tpl1__example_55959141808148_0
timestamp 1707688321
transform 1 0 279 0 1 95
box 0 0 1 1
use sky130_fd_pr__tpl1__example_55959141808148  sky130_fd_pr__tpl1__example_55959141808148_1
timestamp 1707688321
transform 1 0 279 0 1 2247
box 0 0 1 1
use sky130_fd_pr__tpl1__example_55959141808149  sky130_fd_pr__tpl1__example_55959141808149_0
timestamp 1707688321
transform 1 0 449 0 1 1955
box 0 0 1 1
use sky130_fd_pr__tpl1__example_55959141808149  sky130_fd_pr__tpl1__example_55959141808149_1
timestamp 1707688321
transform 1 0 449 0 1 387
box 0 0 1 1
use sky130_fd_pr__tpl1__example_55959141808150  sky130_fd_pr__tpl1__example_55959141808150_0
timestamp 1707688321
transform 1 0 380 0 1 509
box 0 0 1 1
use sky130_fd_pr__tpl1__example_55959141808150  sky130_fd_pr__tpl1__example_55959141808150_1
timestamp 1707688321
transform 1 0 1132 0 1 509
box 0 0 1 1
use sky130_fd_pr__tpl1__example_55959141808151  sky130_fd_pr__tpl1__example_55959141808151_0
timestamp 1707688321
transform 1 0 95 0 1 198
box 0 0 1 1
use sky130_fd_pr__tpl1__example_55959141808151  sky130_fd_pr__tpl1__example_55959141808151_1
timestamp 1707688321
transform 1 0 1414 0 1 198
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808152  sky130_fd_pr__via_l1m1__example_55959141808152_0
timestamp 1707688321
transform 1 0 1118 0 1 108
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808152  sky130_fd_pr__via_l1m1__example_55959141808152_1
timestamp 1707688321
transform 1 0 454 0 1 1969
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808152  sky130_fd_pr__via_l1m1__example_55959141808152_2
timestamp 1707688321
transform 1 0 928 0 1 1969
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808153  sky130_fd_pr__via_l1m1__example_55959141808153_0
timestamp 1707688321
transform 1 0 119 0 1 273
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808153  sky130_fd_pr__via_l1m1__example_55959141808153_1
timestamp 1707688321
transform 1 0 1438 0 1 273
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808154  sky130_fd_pr__via_l1m1__example_55959141808154_0
timestamp 1707688321
transform 1 0 1146 0 1 401
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808154  sky130_fd_pr__via_l1m1__example_55959141808154_1
timestamp 1707688321
transform 1 0 395 0 1 401
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808155  sky130_fd_pr__via_l1m1__example_55959141808155_0
timestamp 1707688321
transform 1 0 915 0 1 757
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808155  sky130_fd_pr__via_l1m1__example_55959141808155_1
timestamp 1707688321
transform 1 0 621 0 1 757
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808156  sky130_fd_pr__via_l1m1__example_55959141808156_0
timestamp 1707688321
transform 1 0 959 0 1 2271
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808156  sky130_fd_pr__via_l1m1__example_55959141808156_1
timestamp 1707688321
transform 1 0 307 0 1 2271
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808157  sky130_fd_pr__via_l1m1__example_55959141808157_0
timestamp 1707688321
transform 1 0 725 0 1 1813
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808147  sky130_fd_pr__via_pol1__example_55959141808147_0
timestamp 1707688321
transform 1 0 660 0 1 1796
box 0 0 1 1
<< labels >>
flabel comment s 1452 1103 1452 1103 0 FreeSans 500 270 0 0 DO NOT MERGE WITH PFET NWELL
flabel comment s 129 1085 129 1085 0 FreeSans 500 90 0 0 DO NOT MERGE WITH PFET NWELL
flabel comment s 783 2298 783 2298 0 FreeSans 500 0 0 0 DO NOT MERGE WITH PFET NWELL
flabel metal1 s 703 2259 852 2359 0 FreeSans 300 0 0 0 GATE
port 1 nsew
flabel metal1 s 68 77 204 117 0 FreeSans 200 0 0 0 NWELLRING
port 2 nsew
flabel metal1 s 628 78 721 118 0 FreeSans 200 0 0 0 VGND
port 3 nsew
flabel metal1 s 387 82 514 122 0 FreeSans 300 0 0 0 NBODY
port 4 nsew
flabel metal1 s 888 70 996 103 0 FreeSans 400 0 0 0 IN
port 5 nsew
<< properties >>
string GDS_END 16799308
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 16794544
<< end >>
