magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< dnwell >>
rect -336 1932 2037 4597
<< pwell >>
rect -88 4263 1789 4349
rect -88 2266 -2 4263
rect 1703 2266 1789 4263
rect -88 2180 1789 2266
<< psubdiff >>
rect -62 4289 29 4323
rect 63 4289 97 4323
rect 131 4289 165 4323
rect 199 4289 233 4323
rect 267 4289 301 4323
rect 335 4289 369 4323
rect 403 4289 437 4323
rect 471 4289 505 4323
rect 539 4289 573 4323
rect 607 4289 641 4323
rect 675 4289 709 4323
rect 743 4289 777 4323
rect 811 4289 845 4323
rect 879 4289 913 4323
rect 947 4289 981 4323
rect 1015 4289 1049 4323
rect 1083 4289 1117 4323
rect 1151 4289 1185 4323
rect 1219 4289 1253 4323
rect 1287 4289 1321 4323
rect 1355 4289 1389 4323
rect 1423 4289 1457 4323
rect 1491 4289 1525 4323
rect 1559 4289 1593 4323
rect 1627 4289 1661 4323
rect 1695 4289 1763 4323
rect -62 4255 -28 4289
rect -62 4187 -28 4221
rect 1729 4212 1763 4289
rect -62 4119 -28 4153
rect 1729 4144 1763 4178
rect -62 4051 -28 4085
rect -62 3983 -28 4017
rect -62 3915 -28 3949
rect -62 3847 -28 3881
rect 1729 4076 1763 4110
rect 1729 4008 1763 4042
rect 1729 3940 1763 3974
rect 1729 3872 1763 3906
rect -62 3779 -28 3813
rect 1729 3804 1763 3838
rect -62 3711 -28 3745
rect -62 3643 -28 3677
rect -62 3575 -28 3609
rect -62 3507 -28 3541
rect 1729 3736 1763 3770
rect 1729 3668 1763 3702
rect 1729 3600 1763 3634
rect 1729 3532 1763 3566
rect -62 3439 -28 3473
rect 1729 3464 1763 3498
rect -62 3371 -28 3405
rect -62 3303 -28 3337
rect -62 3235 -28 3269
rect -62 3167 -28 3201
rect -62 3099 -28 3133
rect -62 3031 -28 3065
rect 1729 3396 1763 3430
rect 1729 3328 1763 3362
rect 1729 3260 1763 3294
rect 1729 3192 1763 3226
rect 1729 3124 1763 3158
rect 1729 3056 1763 3090
rect -62 2963 -28 2997
rect 1729 2988 1763 3022
rect -62 2895 -28 2929
rect -62 2827 -28 2861
rect -62 2759 -28 2793
rect 1729 2920 1763 2954
rect 1729 2852 1763 2886
rect 1729 2784 1763 2818
rect -62 2691 -28 2725
rect 1729 2716 1763 2750
rect -62 2623 -28 2657
rect 1729 2648 1763 2682
rect -62 2555 -28 2589
rect -62 2487 -28 2521
rect -62 2419 -28 2453
rect -62 2351 -28 2385
rect -62 2240 -28 2317
rect 1729 2580 1763 2614
rect 1729 2512 1763 2546
rect 1729 2444 1763 2478
rect 1729 2376 1763 2410
rect 1729 2308 1763 2342
rect 1729 2240 1763 2274
rect -62 2206 6 2240
rect 40 2206 74 2240
rect 108 2206 142 2240
rect 176 2206 210 2240
rect 244 2206 278 2240
rect 312 2206 346 2240
rect 380 2206 414 2240
rect 448 2206 482 2240
rect 516 2206 550 2240
rect 584 2206 618 2240
rect 652 2206 686 2240
rect 720 2206 754 2240
rect 788 2206 822 2240
rect 856 2206 890 2240
rect 924 2206 1021 2240
rect 1055 2206 1089 2240
rect 1123 2206 1157 2240
rect 1191 2206 1225 2240
rect 1259 2206 1293 2240
rect 1327 2206 1361 2240
rect 1395 2206 1429 2240
rect 1463 2206 1497 2240
rect 1531 2206 1565 2240
rect 1599 2206 1633 2240
rect 1667 2206 1763 2240
<< psubdiffcont >>
rect 29 4289 63 4323
rect 97 4289 131 4323
rect 165 4289 199 4323
rect 233 4289 267 4323
rect 301 4289 335 4323
rect 369 4289 403 4323
rect 437 4289 471 4323
rect 505 4289 539 4323
rect 573 4289 607 4323
rect 641 4289 675 4323
rect 709 4289 743 4323
rect 777 4289 811 4323
rect 845 4289 879 4323
rect 913 4289 947 4323
rect 981 4289 1015 4323
rect 1049 4289 1083 4323
rect 1117 4289 1151 4323
rect 1185 4289 1219 4323
rect 1253 4289 1287 4323
rect 1321 4289 1355 4323
rect 1389 4289 1423 4323
rect 1457 4289 1491 4323
rect 1525 4289 1559 4323
rect 1593 4289 1627 4323
rect 1661 4289 1695 4323
rect -62 4221 -28 4255
rect -62 4153 -28 4187
rect 1729 4178 1763 4212
rect -62 4085 -28 4119
rect -62 4017 -28 4051
rect -62 3949 -28 3983
rect -62 3881 -28 3915
rect -62 3813 -28 3847
rect 1729 4110 1763 4144
rect 1729 4042 1763 4076
rect 1729 3974 1763 4008
rect 1729 3906 1763 3940
rect 1729 3838 1763 3872
rect -62 3745 -28 3779
rect 1729 3770 1763 3804
rect -62 3677 -28 3711
rect -62 3609 -28 3643
rect -62 3541 -28 3575
rect -62 3473 -28 3507
rect 1729 3702 1763 3736
rect 1729 3634 1763 3668
rect 1729 3566 1763 3600
rect 1729 3498 1763 3532
rect -62 3405 -28 3439
rect 1729 3430 1763 3464
rect -62 3337 -28 3371
rect -62 3269 -28 3303
rect -62 3201 -28 3235
rect -62 3133 -28 3167
rect -62 3065 -28 3099
rect 1729 3362 1763 3396
rect 1729 3294 1763 3328
rect 1729 3226 1763 3260
rect 1729 3158 1763 3192
rect 1729 3090 1763 3124
rect -62 2997 -28 3031
rect 1729 3022 1763 3056
rect -62 2929 -28 2963
rect -62 2861 -28 2895
rect -62 2793 -28 2827
rect -62 2725 -28 2759
rect 1729 2954 1763 2988
rect 1729 2886 1763 2920
rect 1729 2818 1763 2852
rect 1729 2750 1763 2784
rect -62 2657 -28 2691
rect -62 2589 -28 2623
rect 1729 2682 1763 2716
rect -62 2521 -28 2555
rect -62 2453 -28 2487
rect -62 2385 -28 2419
rect -62 2317 -28 2351
rect 1729 2614 1763 2648
rect 1729 2546 1763 2580
rect 1729 2478 1763 2512
rect 1729 2410 1763 2444
rect 1729 2342 1763 2376
rect 1729 2274 1763 2308
rect 6 2206 40 2240
rect 74 2206 108 2240
rect 142 2206 176 2240
rect 210 2206 244 2240
rect 278 2206 312 2240
rect 346 2206 380 2240
rect 414 2206 448 2240
rect 482 2206 516 2240
rect 550 2206 584 2240
rect 618 2206 652 2240
rect 686 2206 720 2240
rect 754 2206 788 2240
rect 822 2206 856 2240
rect 890 2206 924 2240
rect 1021 2206 1055 2240
rect 1089 2206 1123 2240
rect 1157 2206 1191 2240
rect 1225 2206 1259 2240
rect 1293 2206 1327 2240
rect 1361 2206 1395 2240
rect 1429 2206 1463 2240
rect 1497 2206 1531 2240
rect 1565 2206 1599 2240
rect 1633 2206 1667 2240
<< poly >>
rect 247 4194 535 4210
rect 247 4160 263 4194
rect 297 4160 337 4194
rect 371 4160 411 4194
rect 445 4160 485 4194
rect 519 4160 535 4194
rect 247 4144 535 4160
rect 1016 4194 1304 4210
rect 1016 4160 1032 4194
rect 1066 4160 1106 4194
rect 1140 4160 1180 4194
rect 1214 4160 1254 4194
rect 1288 4160 1304 4194
rect 1016 4144 1304 4160
rect 1134 3810 1562 3826
rect 1134 3776 1150 3810
rect 1184 3776 1222 3810
rect 1256 3776 1294 3810
rect 1328 3776 1366 3810
rect 1400 3776 1439 3810
rect 1473 3776 1512 3810
rect 1546 3776 1562 3810
rect 1134 3760 1562 3776
rect 141 3458 793 3474
rect 141 3424 157 3458
rect 191 3424 231 3458
rect 265 3424 305 3458
rect 339 3424 378 3458
rect 412 3424 451 3458
rect 485 3424 524 3458
rect 558 3424 597 3458
rect 631 3424 670 3458
rect 704 3424 743 3458
rect 777 3424 793 3458
rect 141 3408 793 3424
rect 257 3022 391 3038
rect 257 2988 273 3022
rect 307 2988 341 3022
rect 375 2988 391 3022
rect 257 2972 391 2988
rect 795 2722 929 2738
rect 795 2688 811 2722
rect 845 2688 879 2722
rect 913 2688 929 2722
rect 795 2672 929 2688
rect 1167 2672 1367 2688
rect 1167 2638 1183 2672
rect 1217 2638 1317 2672
rect 1351 2638 1367 2672
rect 1167 2622 1367 2638
rect 854 1883 988 1899
rect 854 1849 870 1883
rect 904 1849 938 1883
rect 972 1849 988 1883
rect 854 1833 988 1849
rect 1346 1750 1412 1766
rect 1346 1716 1362 1750
rect 1396 1716 1412 1750
rect 1346 1682 1412 1716
rect 1346 1648 1362 1682
rect 1396 1648 1412 1682
rect 1346 1632 1412 1648
rect 1346 1364 1412 1380
rect 1346 1330 1362 1364
rect 1396 1330 1412 1364
rect 1346 1296 1412 1330
rect 1346 1262 1362 1296
rect 1396 1262 1412 1296
rect 1346 1246 1412 1262
rect 447 1153 581 1169
rect 447 1119 463 1153
rect 497 1119 531 1153
rect 565 1119 581 1153
rect 447 1103 581 1119
<< polycont >>
rect 263 4160 297 4194
rect 337 4160 371 4194
rect 411 4160 445 4194
rect 485 4160 519 4194
rect 1032 4160 1066 4194
rect 1106 4160 1140 4194
rect 1180 4160 1214 4194
rect 1254 4160 1288 4194
rect 1150 3776 1184 3810
rect 1222 3776 1256 3810
rect 1294 3776 1328 3810
rect 1366 3776 1400 3810
rect 1439 3776 1473 3810
rect 1512 3776 1546 3810
rect 157 3424 191 3458
rect 231 3424 265 3458
rect 305 3424 339 3458
rect 378 3424 412 3458
rect 451 3424 485 3458
rect 524 3424 558 3458
rect 597 3424 631 3458
rect 670 3424 704 3458
rect 743 3424 777 3458
rect 273 2988 307 3022
rect 341 2988 375 3022
rect 811 2688 845 2722
rect 879 2688 913 2722
rect 1183 2638 1217 2672
rect 1317 2638 1351 2672
rect 870 1849 904 1883
rect 938 1849 972 1883
rect 1362 1716 1396 1750
rect 1362 1648 1396 1682
rect 1362 1330 1396 1364
rect 1362 1262 1396 1296
rect 463 1119 497 1153
rect 531 1119 565 1153
<< locali >>
rect -62 4289 29 4323
rect 63 4289 97 4323
rect 131 4289 165 4323
rect 199 4289 233 4323
rect 267 4289 301 4323
rect 335 4289 369 4323
rect 403 4289 437 4323
rect 471 4289 505 4323
rect 539 4289 573 4323
rect 607 4289 641 4323
rect 675 4289 709 4323
rect 743 4289 777 4323
rect 811 4289 845 4323
rect 879 4289 913 4323
rect 947 4289 981 4323
rect 1015 4289 1049 4323
rect 1083 4289 1117 4323
rect 1151 4289 1185 4323
rect 1219 4289 1253 4323
rect 1287 4289 1321 4323
rect 1355 4289 1389 4323
rect 1423 4289 1457 4323
rect 1491 4289 1525 4323
rect 1559 4289 1593 4323
rect 1627 4289 1661 4323
rect 1695 4289 1763 4323
rect -62 4255 -28 4289
rect -62 4187 -28 4221
rect 1729 4212 1763 4289
rect 247 4160 263 4194
rect 297 4160 326 4194
rect 371 4160 398 4194
rect 445 4160 485 4194
rect 519 4160 535 4194
rect 1016 4160 1032 4194
rect 1066 4160 1106 4194
rect 1158 4160 1180 4194
rect 1230 4160 1254 4194
rect 1288 4160 1304 4194
rect -62 4119 -28 4153
rect 1729 4144 1763 4178
rect -62 4051 -28 4076
rect -62 3983 -28 3992
rect -62 3942 -28 3949
rect 134 4076 168 4110
rect 202 4076 236 4110
rect 134 4026 236 4076
rect 134 3992 168 4026
rect 202 3992 236 4026
rect 134 3942 236 3992
rect 134 3908 168 3942
rect 202 3908 236 3942
rect -62 3847 -28 3881
rect -62 3779 -28 3813
rect 277 3798 333 4112
rect 374 4038 408 4076
rect 449 3798 505 4112
rect 546 4076 580 4110
rect 614 4076 648 4110
rect 546 4026 648 4076
rect 546 3992 580 4026
rect 614 3992 648 4026
rect 546 3942 648 3992
rect 546 3908 580 3942
rect 614 3908 648 3942
rect 903 4076 937 4110
rect 971 4076 1005 4110
rect 903 4026 1005 4076
rect 903 3992 937 4026
rect 971 3992 1005 4026
rect 1143 4042 1177 4080
rect 1315 4076 1349 4110
rect 1383 4076 1417 4110
rect 1315 4026 1417 4076
rect 903 3942 1005 3992
rect 1315 3992 1349 4026
rect 1383 3992 1417 4026
rect 903 3908 937 3942
rect 971 3908 1005 3942
rect 1057 3882 1091 3920
rect 1229 3882 1263 3920
rect 1315 3942 1417 3992
rect 1315 3908 1349 3942
rect 1383 3908 1417 3942
rect 1729 4026 1763 4042
rect 1729 3942 1763 3974
rect 1729 3872 1763 3906
rect -62 3711 -28 3745
rect -62 3643 -28 3677
rect -62 3575 -28 3609
rect -62 3507 -28 3541
rect 88 3748 613 3798
rect 1134 3776 1150 3810
rect 1184 3776 1222 3810
rect 1256 3776 1294 3810
rect 1328 3776 1366 3810
rect 1417 3776 1439 3810
rect 1489 3776 1512 3810
rect 1546 3776 1562 3810
rect 1729 3804 1763 3838
rect 88 3506 141 3748
rect 299 3579 405 3710
rect 333 3545 371 3579
rect 299 3508 405 3545
rect 557 3506 613 3748
rect 1729 3736 1763 3770
rect 768 3579 874 3710
rect 1729 3668 1763 3702
rect 802 3545 840 3579
rect 1089 3585 1123 3623
rect 1729 3600 1763 3634
rect 768 3508 874 3545
rect 1729 3532 1763 3566
rect -62 3439 -28 3473
rect 1729 3464 1763 3498
rect 141 3424 157 3458
rect 191 3424 231 3458
rect 265 3424 305 3458
rect 339 3424 378 3458
rect 412 3424 451 3458
rect 485 3424 523 3458
rect 558 3424 595 3458
rect 631 3424 670 3458
rect 704 3424 743 3458
rect 777 3424 793 3458
rect -62 3371 -28 3405
rect 1729 3396 1763 3430
rect -62 3303 -28 3337
rect -62 3235 -28 3269
rect -62 3167 -28 3201
rect 60 3340 231 3374
rect 60 3306 191 3340
rect 225 3306 231 3340
rect 60 3268 231 3306
rect 60 3234 191 3268
rect 225 3234 231 3268
rect 60 3172 231 3234
rect 299 3243 405 3374
rect 333 3209 371 3243
rect 299 3172 405 3209
rect 532 3346 638 3374
rect 566 3312 604 3346
rect 532 3172 638 3312
rect 768 3243 874 3374
rect 1729 3328 1763 3362
rect 1729 3260 1763 3294
rect 802 3209 840 3243
rect 768 3172 874 3209
rect 1397 3174 1431 3212
rect -62 3099 -28 3133
rect 1227 3120 1265 3154
rect 1573 3174 1607 3212
rect 1729 3192 1763 3226
rect 1729 3124 1763 3158
rect -62 3031 -28 3065
rect 1729 3056 1763 3090
rect 365 3022 403 3028
rect -62 2963 -28 2997
rect 257 2988 273 3022
rect 307 2994 331 3022
rect 375 2994 403 3022
rect 307 2988 341 2994
rect 375 2988 391 2994
rect 1729 2988 1763 3022
rect 1729 2940 1763 2954
rect -62 2895 -28 2906
rect 729 2856 767 2890
rect -62 2827 -28 2829
rect -62 2786 -28 2793
rect -62 2709 -28 2725
rect 935 2770 973 2804
rect 393 2726 427 2764
rect 1058 2752 1168 2924
rect 1344 2812 1378 2850
rect 1729 2863 1763 2886
rect 1729 2786 1763 2818
rect 1058 2734 1202 2752
rect 795 2688 807 2722
rect 845 2688 879 2722
rect 913 2688 929 2722
rect 1007 2710 1202 2734
rect 1729 2716 1763 2750
rect -62 2632 -28 2657
rect -62 2555 -28 2589
rect -62 2487 -28 2521
rect -62 2419 -28 2444
rect 217 2400 251 2438
rect 757 2400 791 2438
rect -62 2351 -28 2366
rect -62 2240 -28 2317
rect 858 2312 967 2638
rect 883 2278 921 2312
rect 955 2278 967 2312
rect 1007 2610 1129 2710
rect 1167 2638 1183 2672
rect 1217 2638 1253 2672
rect 1287 2638 1317 2672
rect 1359 2638 1367 2672
rect 1729 2648 1763 2675
rect 1007 2312 1082 2610
rect 1729 2580 1763 2598
rect 1361 2564 1653 2570
rect 1361 2530 1364 2564
rect 1398 2530 1436 2564
rect 1470 2558 1653 2564
rect 1470 2530 1613 2558
rect 1361 2524 1613 2530
rect 1647 2524 1653 2558
rect 1361 2486 1653 2524
rect 1122 2400 1156 2438
rect 1361 2452 1613 2486
rect 1647 2452 1653 2486
rect 1361 2436 1653 2452
rect 1729 2512 1763 2521
rect 1729 2400 1763 2410
rect 1007 2278 1019 2312
rect 1053 2278 1091 2312
rect 1729 2308 1763 2342
rect 1729 2240 1763 2274
rect -62 2206 6 2240
rect 40 2206 74 2240
rect 108 2206 142 2240
rect 176 2206 210 2240
rect 244 2206 278 2240
rect 312 2206 346 2240
rect 380 2206 414 2240
rect 448 2206 482 2240
rect 516 2206 550 2240
rect 584 2206 618 2240
rect 652 2206 686 2240
rect 720 2206 754 2240
rect 788 2206 822 2240
rect 856 2206 890 2240
rect 924 2206 1021 2240
rect 1055 2206 1089 2240
rect 1123 2206 1157 2240
rect 1191 2206 1225 2240
rect 1259 2206 1293 2240
rect 1327 2206 1361 2240
rect 1395 2206 1429 2240
rect 1463 2206 1497 2240
rect 1531 2206 1565 2240
rect 1599 2206 1633 2240
rect 1667 2206 1763 2240
rect 854 1849 870 1883
rect 904 1849 938 1883
rect 972 1849 1294 1883
rect 889 1793 1294 1849
rect 889 1775 1168 1793
rect 408 1658 442 1696
rect 686 1558 746 1751
rect 643 1524 709 1558
rect 743 1524 809 1558
rect 609 1474 843 1524
rect 643 1440 709 1474
rect 743 1440 809 1474
rect 686 1197 746 1440
rect 889 1390 950 1775
rect 1202 1759 1240 1793
rect 1274 1775 1294 1793
rect 1362 1750 1396 1766
rect 990 1658 1024 1696
rect 1362 1699 1396 1716
rect 1362 1682 1365 1699
rect 1399 1665 1449 1699
rect 1483 1665 1532 1699
rect 1362 1632 1396 1648
rect 1160 1524 1184 1535
rect 1218 1524 1256 1558
rect 1290 1524 1306 1535
rect 1160 1475 1306 1524
rect 1184 1474 1290 1475
rect 1218 1440 1256 1474
rect 889 1356 905 1390
rect 939 1356 950 1390
rect 889 1318 950 1356
rect 1362 1364 1396 1380
rect 889 1284 905 1318
rect 939 1284 950 1318
rect 1310 1300 1348 1334
rect 1382 1300 1396 1330
rect 889 1237 950 1284
rect 1362 1296 1396 1300
rect 1362 1246 1396 1262
rect 1160 1153 1294 1217
rect 447 1119 460 1153
rect 497 1119 531 1153
rect 566 1119 581 1153
rect 1160 1119 1168 1153
rect 1202 1119 1240 1153
rect 1274 1119 1294 1153
rect 1436 1153 1566 1665
rect 1436 1119 1448 1153
rect 1482 1119 1520 1153
rect 1554 1119 1566 1153
<< viali >>
rect 326 4160 337 4194
rect 337 4160 360 4194
rect 398 4160 411 4194
rect 411 4160 432 4194
rect 1124 4160 1140 4194
rect 1140 4160 1158 4194
rect 1196 4160 1214 4194
rect 1214 4160 1230 4194
rect -62 4085 -28 4110
rect -62 4076 -28 4085
rect -62 4017 -28 4026
rect -62 3992 -28 4017
rect -62 3915 -28 3942
rect -62 3908 -28 3915
rect 168 4076 202 4110
rect 168 3992 202 4026
rect 168 3908 202 3942
rect 374 4076 408 4110
rect 374 4004 408 4038
rect 580 4076 614 4110
rect 580 3992 614 4026
rect 580 3908 614 3942
rect 937 4076 971 4110
rect 937 3992 971 4026
rect 1143 4080 1177 4114
rect 1143 4008 1177 4042
rect 1349 4076 1383 4110
rect 1349 3992 1383 4026
rect 937 3908 971 3942
rect 1057 3920 1091 3954
rect 1057 3848 1091 3882
rect 1229 3920 1263 3954
rect 1349 3908 1383 3942
rect 1729 4076 1763 4110
rect 1729 4008 1763 4026
rect 1729 3992 1763 4008
rect 1729 3940 1763 3942
rect 1729 3908 1763 3940
rect 1229 3848 1263 3882
rect 1383 3776 1400 3810
rect 1400 3776 1417 3810
rect 1455 3776 1473 3810
rect 1473 3776 1489 3810
rect 299 3545 333 3579
rect 371 3545 405 3579
rect 768 3545 802 3579
rect 840 3545 874 3579
rect 1089 3623 1123 3657
rect 1089 3551 1123 3585
rect 523 3424 524 3458
rect 524 3424 557 3458
rect 595 3424 597 3458
rect 597 3424 629 3458
rect 191 3306 225 3340
rect 191 3234 225 3268
rect 299 3209 333 3243
rect 371 3209 405 3243
rect 532 3312 566 3346
rect 604 3312 638 3346
rect 768 3209 802 3243
rect 840 3209 874 3243
rect 1397 3212 1431 3246
rect 1193 3120 1227 3154
rect 1265 3120 1299 3154
rect 1397 3140 1431 3174
rect 1573 3212 1607 3246
rect 1573 3140 1607 3174
rect 331 3022 365 3028
rect 331 2994 341 3022
rect 341 2994 365 3022
rect 403 2994 437 3028
rect -62 2929 -28 2940
rect -62 2906 -28 2929
rect -62 2861 -28 2863
rect -62 2829 -28 2861
rect 695 2856 729 2890
rect 767 2856 801 2890
rect -62 2759 -28 2786
rect -62 2752 -28 2759
rect -62 2691 -28 2709
rect 393 2764 427 2798
rect 901 2770 935 2804
rect 973 2770 1007 2804
rect 1729 2920 1763 2940
rect 1729 2906 1763 2920
rect 1344 2850 1378 2884
rect 1344 2778 1378 2812
rect 1729 2852 1763 2863
rect 1729 2829 1763 2852
rect 1729 2784 1763 2786
rect 1729 2752 1763 2784
rect 393 2692 427 2726
rect -62 2675 -28 2691
rect 807 2688 811 2722
rect 811 2688 841 2722
rect 879 2688 913 2722
rect -62 2623 -28 2632
rect -62 2598 -28 2623
rect -62 2521 -28 2555
rect -62 2453 -28 2478
rect -62 2444 -28 2453
rect -62 2385 -28 2400
rect -62 2366 -28 2385
rect 217 2438 251 2472
rect 217 2366 251 2400
rect 757 2438 791 2472
rect 757 2366 791 2400
rect 849 2278 883 2312
rect 921 2278 955 2312
rect 1729 2682 1763 2709
rect 1729 2675 1763 2682
rect 1253 2638 1287 2672
rect 1325 2638 1351 2672
rect 1351 2638 1359 2672
rect 1729 2614 1763 2632
rect 1729 2598 1763 2614
rect 1364 2530 1398 2564
rect 1436 2530 1470 2564
rect 1613 2524 1647 2558
rect 1122 2438 1156 2472
rect 1613 2452 1647 2486
rect 1729 2546 1763 2555
rect 1729 2521 1763 2546
rect 1729 2444 1763 2478
rect 1122 2366 1156 2400
rect 1729 2376 1763 2400
rect 1729 2366 1763 2376
rect 1019 2278 1053 2312
rect 1091 2278 1125 2312
rect 408 1696 442 1730
rect 408 1624 442 1658
rect 609 1524 643 1558
rect 709 1524 743 1558
rect 809 1524 843 1558
rect 609 1440 643 1474
rect 709 1440 743 1474
rect 809 1440 843 1474
rect 1168 1759 1202 1793
rect 1240 1759 1274 1793
rect 990 1696 1024 1730
rect 990 1624 1024 1658
rect 1365 1682 1399 1699
rect 1365 1665 1396 1682
rect 1396 1665 1399 1682
rect 1449 1665 1483 1699
rect 1532 1665 1566 1699
rect 1184 1524 1218 1558
rect 1256 1524 1290 1558
rect 1184 1440 1218 1474
rect 1256 1440 1290 1474
rect 905 1356 939 1390
rect 905 1284 939 1318
rect 1276 1300 1310 1334
rect 1348 1330 1362 1334
rect 1362 1330 1382 1334
rect 1348 1300 1382 1330
rect 460 1119 463 1153
rect 463 1119 494 1153
rect 532 1119 565 1153
rect 565 1119 566 1153
rect 1168 1119 1202 1153
rect 1240 1119 1274 1153
rect 1448 1119 1482 1153
rect 1520 1119 1554 1153
<< metal1 >>
rect 314 4194 444 4200
rect 314 4160 326 4194
rect 360 4160 398 4194
rect 432 4160 444 4194
rect 314 4154 444 4160
rect 1112 4194 1242 4200
rect 1112 4160 1124 4194
rect 1158 4160 1196 4194
rect 1230 4160 1242 4194
rect 1112 4154 1242 4160
tri 1005 4122 1009 4126 se
rect 1009 4122 1015 4126
rect -68 4110 1015 4122
rect -68 4076 -62 4110
rect -28 4076 168 4110
rect 202 4076 374 4110
rect 408 4076 580 4110
rect 614 4076 937 4110
rect 971 4076 1015 4110
rect -68 4074 1015 4076
rect 1067 4074 1079 4126
rect 1131 4122 1183 4126
tri 1183 4122 1187 4126 sw
rect 1131 4114 1769 4122
rect 1131 4080 1143 4114
rect 1177 4110 1769 4114
rect 1177 4080 1349 4110
rect 1131 4076 1349 4080
rect 1383 4076 1729 4110
rect 1763 4076 1769 4110
rect 1131 4074 1769 4076
rect -68 4048 1769 4074
rect -68 4038 1015 4048
rect -68 4026 374 4038
rect -68 3992 -62 4026
rect -28 3992 168 4026
rect 202 4004 374 4026
rect 408 4026 1015 4038
rect 408 4004 580 4026
rect 202 3996 580 4004
rect 202 3992 279 3996
tri 279 3992 283 3996 nw
tri 364 3992 368 3996 ne
rect 368 3992 414 3996
tri 414 3992 418 3996 nw
tri 499 3992 503 3996 ne
rect 503 3992 580 3996
rect 614 3996 937 4026
rect 614 3992 691 3996
tri 691 3992 695 3996 nw
tri 856 3992 860 3996 ne
rect 860 3992 937 3996
rect 971 3996 1015 4026
rect 1067 3996 1079 4048
rect 1131 4042 1769 4048
rect 1131 4008 1143 4042
rect 1177 4026 1769 4042
rect 1177 4008 1349 4026
rect 1131 3996 1349 4008
rect 971 3992 1036 3996
tri 1036 3992 1040 3996 nw
tri 1280 3992 1284 3996 ne
rect 1284 3992 1349 3996
rect 1383 3996 1729 4026
rect 1383 3992 1460 3996
tri 1460 3992 1464 3996 nw
tri 1682 3992 1686 3996 ne
rect 1686 3992 1729 3996
rect 1763 3992 1769 4026
rect -68 3966 253 3992
tri 253 3966 279 3992 nw
tri 503 3966 529 3992 ne
rect 529 3966 665 3992
tri 665 3966 691 3992 nw
tri 860 3966 886 3992 ne
rect 886 3966 1011 3992
tri 1011 3967 1036 3992 nw
tri 1284 3967 1309 3992 ne
rect 1309 3966 1434 3992
tri 1434 3966 1460 3992 nw
tri 1686 3966 1712 3992 ne
rect 1712 3966 1769 3992
rect -68 3942 242 3966
tri 242 3955 253 3966 nw
tri 529 3955 540 3966 ne
rect -68 3908 -62 3942
rect -28 3908 168 3942
rect 202 3908 242 3942
rect -68 3896 242 3908
rect 540 3942 654 3966
tri 654 3955 665 3966 nw
tri 886 3955 897 3966 ne
rect 540 3908 580 3942
rect 614 3908 654 3942
rect 540 3896 654 3908
rect 897 3942 1011 3966
rect 897 3908 937 3942
rect 971 3908 1011 3942
rect 897 3896 1011 3908
rect 1051 3960 1269 3966
rect 1051 3954 1217 3960
rect 1051 3920 1057 3954
rect 1091 3920 1217 3954
rect 1051 3908 1217 3920
rect 1051 3896 1269 3908
rect 1309 3942 1423 3966
tri 1423 3955 1434 3966 nw
tri 1712 3955 1723 3966 ne
rect 1309 3908 1349 3942
rect 1383 3908 1423 3942
rect 1309 3896 1423 3908
rect 1723 3942 1769 3966
rect 1723 3908 1729 3942
rect 1763 3908 1769 3942
rect 1723 3896 1769 3908
rect 1051 3882 1217 3896
rect 1051 3848 1057 3882
rect 1091 3848 1217 3882
rect 1051 3844 1217 3848
rect 1051 3836 1269 3844
rect 1371 3810 1501 3816
rect 1371 3776 1383 3810
rect 1417 3776 1455 3810
rect 1489 3776 1501 3810
rect 1371 3770 1501 3776
rect 1083 3657 1129 3669
rect 1083 3623 1089 3657
rect 1123 3623 1129 3657
tri 1053 3585 1083 3615 se
rect 1083 3585 1129 3623
rect 287 3579 1089 3585
rect 287 3545 299 3579
rect 333 3545 371 3579
rect 405 3545 768 3579
rect 802 3545 840 3579
rect 874 3551 1089 3579
rect 1123 3551 1129 3585
rect 874 3545 1129 3551
rect 287 3539 1129 3545
rect 511 3458 641 3464
rect 511 3424 523 3458
rect 557 3424 595 3458
rect 629 3424 641 3458
rect 511 3418 641 3424
rect 185 3346 1227 3352
rect 185 3340 532 3346
rect 185 3306 191 3340
rect 225 3312 532 3340
rect 566 3312 604 3346
rect 638 3312 1227 3346
rect 225 3306 1227 3312
rect 185 3300 261 3306
tri 261 3300 267 3306 nw
tri 1215 3300 1221 3306 ne
rect 1221 3300 1227 3306
rect 1279 3300 1291 3352
rect 1343 3300 1349 3352
rect 185 3268 231 3300
tri 231 3270 261 3300 nw
rect 185 3234 191 3268
rect 225 3234 231 3268
tri 1382 3249 1391 3258 se
rect 1391 3249 1437 3258
rect 185 3222 231 3234
rect 287 3246 1437 3249
rect 287 3243 1397 3246
rect 287 3209 299 3243
rect 333 3209 371 3243
rect 405 3209 768 3243
rect 802 3209 840 3243
rect 874 3212 1397 3243
rect 1431 3212 1437 3246
rect 874 3209 1437 3212
rect 287 3203 1437 3209
tri 1355 3174 1384 3203 ne
rect 1384 3174 1437 3203
tri 1384 3167 1391 3174 ne
tri 1218 3160 1221 3163 se
rect 1221 3160 1227 3163
rect 1181 3154 1227 3160
rect 1279 3154 1291 3163
rect 1181 3120 1193 3154
rect 1181 3114 1227 3120
tri 1218 3111 1221 3114 ne
rect 1221 3111 1227 3114
rect 1279 3111 1291 3120
rect 1343 3111 1349 3163
rect 1391 3140 1397 3174
rect 1431 3140 1437 3174
rect 1391 3128 1437 3140
rect 1567 3256 1613 3258
tri 1613 3256 1615 3258 sw
rect 1567 3250 1656 3256
rect 1567 3246 1604 3250
rect 1567 3212 1573 3246
rect 1567 3198 1604 3212
rect 1567 3186 1656 3198
rect 1567 3174 1604 3186
rect 1567 3140 1573 3174
rect 1567 3134 1604 3140
rect 1567 3128 1656 3134
rect 319 3028 449 3034
rect 319 2994 331 3028
rect 365 2994 403 3028
rect 437 2994 449 3028
rect 319 2988 449 2994
rect -68 2940 1769 2952
rect -68 2906 -62 2940
rect -28 2906 1729 2940
rect 1763 2906 1769 2940
rect -68 2890 1769 2906
rect -68 2863 695 2890
rect -68 2829 -62 2863
rect -28 2856 695 2863
rect 729 2856 767 2890
rect 801 2884 1769 2890
rect 801 2856 1344 2884
rect -28 2850 1344 2856
rect 1378 2863 1769 2884
rect 1378 2850 1729 2863
rect -28 2829 192 2850
tri 192 2829 213 2850 nw
tri 1270 2829 1291 2850 ne
rect 1291 2829 1729 2850
rect 1763 2829 1769 2863
rect -68 2812 175 2829
tri 175 2812 192 2829 nw
tri 1291 2812 1308 2829 ne
rect 1308 2812 1769 2829
rect -68 2804 167 2812
tri 167 2804 175 2812 nw
tri 1308 2810 1310 2812 ne
rect 1310 2810 1344 2812
rect 387 2804 1019 2810
tri 1310 2808 1312 2810 ne
rect -68 2798 161 2804
tri 161 2798 167 2804 nw
rect 387 2798 901 2804
rect -68 2786 129 2798
rect -68 2752 -62 2786
rect -28 2766 129 2786
tri 129 2766 161 2798 nw
rect -28 2764 127 2766
tri 127 2764 129 2766 nw
rect 387 2764 393 2798
rect 427 2770 901 2798
rect 935 2770 973 2804
rect 1007 2770 1019 2804
rect 427 2764 1019 2770
rect 1312 2778 1344 2810
rect 1378 2786 1769 2812
rect 1378 2778 1729 2786
rect 1312 2766 1729 2778
tri 1670 2764 1672 2766 ne
rect 1672 2764 1729 2766
rect -28 2752 115 2764
tri 115 2752 127 2764 nw
rect 387 2752 456 2764
tri 456 2752 468 2764 nw
tri 932 2752 944 2764 ne
rect 944 2752 1013 2764
tri 1013 2758 1019 2764 nw
tri 1672 2758 1678 2764 ne
rect 1678 2758 1729 2764
tri 1678 2752 1684 2758 ne
rect 1684 2752 1729 2758
rect 1763 2752 1769 2786
rect -68 2709 95 2752
tri 95 2732 115 2752 nw
rect 387 2732 436 2752
tri 436 2732 456 2752 nw
tri 944 2732 964 2752 ne
rect 964 2732 1013 2752
rect -68 2675 -62 2709
rect -28 2675 95 2709
rect 387 2726 433 2732
tri 433 2729 436 2732 nw
tri 964 2729 967 2732 ne
rect 387 2692 393 2726
rect 427 2692 433 2726
rect 387 2680 433 2692
rect 795 2722 925 2728
rect 795 2688 807 2722
rect 841 2688 879 2722
rect 913 2688 925 2722
rect 795 2682 925 2688
rect 967 2713 1013 2732
tri 1684 2729 1707 2752 ne
rect 1707 2729 1769 2752
tri 1707 2718 1718 2729 ne
rect 1718 2718 1769 2729
tri 1013 2713 1018 2718 sw
tri 1718 2713 1723 2718 ne
rect 967 2709 1018 2713
tri 1018 2709 1022 2713 sw
rect 1723 2709 1769 2718
rect 967 2698 1022 2709
tri 967 2682 983 2698 ne
rect 983 2682 1022 2698
tri 1022 2682 1049 2709 sw
tri 802 2680 804 2682 ne
rect 804 2681 917 2682
tri 917 2681 918 2682 nw
tri 983 2681 984 2682 ne
rect 984 2681 1049 2682
tri 1049 2681 1050 2682 sw
rect 804 2680 911 2681
tri 804 2675 809 2680 ne
rect 809 2675 911 2680
tri 911 2675 917 2681 nw
tri 984 2678 987 2681 ne
rect 987 2678 1050 2681
tri 1050 2678 1053 2681 sw
tri 1218 2678 1221 2681 se
rect 1221 2678 1227 2681
tri 987 2675 990 2678 ne
rect 990 2675 1227 2678
rect -68 2632 95 2675
tri 809 2672 812 2675 ne
rect 812 2672 908 2675
tri 908 2672 911 2675 nw
tri 990 2672 993 2675 ne
rect 993 2672 1227 2675
rect 1279 2672 1291 2681
rect 1343 2678 1349 2681
tri 1349 2678 1352 2681 sw
rect 1343 2672 1371 2678
tri 812 2647 837 2672 ne
rect -68 2598 -62 2632
rect -28 2598 95 2632
tri 95 2598 99 2602 sw
rect 837 2598 883 2672
tri 883 2647 908 2672 nw
tri 993 2652 1013 2672 ne
rect 1013 2652 1227 2672
tri 1013 2647 1018 2652 ne
rect 1018 2647 1227 2652
tri 1018 2638 1027 2647 ne
rect 1027 2638 1227 2647
rect 1287 2638 1291 2672
rect 1359 2638 1371 2672
tri 1027 2632 1033 2638 ne
rect 1033 2632 1227 2638
tri 1218 2629 1221 2632 ne
rect 1221 2629 1227 2632
rect 1279 2629 1291 2638
rect 1343 2632 1371 2638
rect 1723 2675 1729 2709
rect 1763 2675 1769 2709
rect 1723 2632 1769 2675
rect 1343 2629 1349 2632
tri 1349 2629 1352 2632 nw
tri 883 2598 890 2605 sw
rect 1723 2598 1729 2632
rect 1763 2598 1769 2632
rect -68 2570 99 2598
tri 99 2570 127 2598 sw
rect 837 2570 890 2598
tri 890 2570 918 2598 sw
rect -68 2564 127 2570
tri 127 2564 133 2570 sw
rect 837 2564 1653 2570
rect -68 2555 133 2564
rect -68 2521 -62 2555
rect -28 2530 133 2555
tri 133 2530 167 2564 sw
rect 837 2530 1364 2564
rect 1398 2530 1436 2564
rect 1470 2560 1653 2564
rect 1470 2530 1601 2560
rect -28 2524 167 2530
tri 167 2524 173 2530 sw
rect 837 2524 1601 2530
rect -28 2521 173 2524
tri 173 2521 176 2524 sw
tri 1563 2521 1566 2524 ne
rect 1566 2521 1601 2524
rect -68 2486 176 2521
tri 176 2486 211 2521 sw
tri 1566 2486 1601 2521 ne
rect 1601 2496 1653 2508
rect -68 2484 211 2486
tri 211 2484 213 2486 sw
rect -68 2478 1015 2484
rect -68 2444 -62 2478
rect -28 2472 1015 2478
rect -28 2444 217 2472
rect -68 2438 217 2444
rect 251 2438 757 2472
rect 791 2438 1015 2472
rect -68 2432 1015 2438
rect 1067 2432 1079 2484
rect 1131 2472 1162 2484
rect 1156 2438 1162 2472
rect 1601 2438 1653 2444
rect 1723 2555 1769 2598
rect 1723 2521 1729 2555
rect 1763 2521 1769 2555
rect 1723 2478 1769 2521
rect 1723 2444 1729 2478
rect 1763 2444 1769 2478
rect 1131 2432 1162 2438
rect -68 2406 1162 2432
rect -68 2400 1015 2406
rect -68 2366 -62 2400
rect -28 2366 217 2400
rect 251 2366 757 2400
rect 791 2366 1015 2400
rect -68 2354 1015 2366
rect 1067 2354 1079 2406
rect 1131 2400 1162 2406
rect 1156 2366 1162 2400
rect 1131 2354 1162 2366
rect 1723 2400 1769 2444
rect 1723 2366 1729 2400
rect 1763 2366 1769 2400
rect 1723 2354 1769 2366
tri 837 2318 839 2320 se
rect 839 2318 845 2321
rect 837 2272 845 2318
tri 837 2270 839 2272 ne
rect 839 2269 845 2272
rect 897 2269 909 2321
rect 961 2269 967 2321
rect 1007 2269 1013 2321
rect 1065 2269 1077 2321
rect 1129 2318 1135 2321
tri 1135 2318 1137 2320 sw
rect 1129 2272 1137 2318
rect 1129 2269 1135 2272
tri 1135 2270 1137 2272 nw
tri 1218 1799 1221 1802 se
rect 1221 1799 1227 1802
rect 1156 1793 1227 1799
rect 866 1776 918 1782
rect 402 1730 448 1742
rect 402 1696 408 1730
rect 442 1700 448 1730
tri 857 1719 866 1728 se
rect 1156 1759 1168 1793
rect 1202 1759 1227 1793
rect 1156 1753 1227 1759
tri 1218 1750 1221 1753 ne
rect 1221 1750 1227 1753
rect 1279 1750 1291 1802
rect 1343 1750 1349 1802
rect 1600 1781 1652 1787
rect 866 1719 918 1724
tri 448 1700 467 1719 sw
tri 838 1700 857 1719 se
rect 857 1712 918 1719
rect 857 1700 866 1712
rect 442 1696 866 1700
rect 402 1660 866 1696
rect 402 1658 918 1660
rect 402 1624 408 1658
rect 442 1654 918 1658
rect 984 1736 1078 1742
rect 984 1730 1026 1736
rect 984 1696 990 1730
rect 1024 1696 1026 1730
rect 984 1684 1026 1696
tri 1565 1705 1600 1740 se
rect 1600 1717 1652 1729
rect 984 1672 1078 1684
rect 984 1658 1026 1672
rect 442 1624 448 1654
tri 448 1632 470 1654 nw
rect 402 1612 448 1624
rect 984 1624 990 1658
rect 1024 1624 1026 1658
rect 984 1620 1026 1624
rect 1353 1699 1600 1705
rect 1353 1665 1365 1699
rect 1399 1665 1449 1699
rect 1483 1665 1532 1699
rect 1566 1665 1600 1699
rect 1353 1659 1652 1665
rect 984 1614 1078 1620
rect 984 1612 1030 1614
tri 1030 1612 1032 1614 nw
rect 264 1558 1652 1564
rect 264 1524 609 1558
rect 643 1524 709 1558
rect 743 1524 809 1558
rect 843 1524 1184 1558
rect 1218 1524 1256 1558
rect 1290 1524 1652 1558
rect 264 1474 1652 1524
rect 264 1440 609 1474
rect 643 1440 709 1474
rect 743 1440 809 1474
rect 843 1440 1184 1474
rect 1218 1440 1256 1474
rect 1290 1440 1652 1474
rect 264 1434 1652 1440
rect 899 1390 945 1402
rect 899 1356 905 1390
rect 939 1356 945 1390
rect 899 1340 945 1356
tri 945 1340 970 1365 sw
rect 899 1334 1394 1340
rect 899 1318 1276 1334
rect 899 1284 905 1318
rect 939 1300 1276 1318
rect 1310 1300 1348 1334
rect 1382 1300 1394 1334
rect 939 1294 1394 1300
rect 939 1284 945 1294
rect 899 1272 945 1284
tri 945 1272 967 1294 nw
rect 448 1153 1566 1159
rect 448 1119 460 1153
rect 494 1119 532 1153
rect 566 1119 1168 1153
rect 1202 1119 1240 1153
rect 1274 1119 1448 1153
rect 1482 1119 1520 1153
rect 1554 1119 1566 1153
rect 448 1113 1566 1119
<< via1 >>
rect 1015 4074 1067 4126
rect 1079 4074 1131 4126
rect 1015 3996 1067 4048
rect 1079 3996 1131 4048
rect 1217 3954 1269 3960
rect 1217 3920 1229 3954
rect 1229 3920 1263 3954
rect 1263 3920 1269 3954
rect 1217 3908 1269 3920
rect 1217 3882 1269 3896
rect 1217 3848 1229 3882
rect 1229 3848 1263 3882
rect 1263 3848 1269 3882
rect 1217 3844 1269 3848
rect 1227 3300 1279 3352
rect 1291 3300 1343 3352
rect 1227 3154 1279 3163
rect 1291 3154 1343 3163
rect 1227 3120 1265 3154
rect 1265 3120 1279 3154
rect 1291 3120 1299 3154
rect 1299 3120 1343 3154
rect 1227 3111 1279 3120
rect 1291 3111 1343 3120
rect 1604 3246 1656 3250
rect 1604 3212 1607 3246
rect 1607 3212 1656 3246
rect 1604 3198 1656 3212
rect 1604 3174 1656 3186
rect 1604 3140 1607 3174
rect 1607 3140 1656 3174
rect 1604 3134 1656 3140
rect 1227 2672 1279 2681
rect 1291 2672 1343 2681
rect 1227 2638 1253 2672
rect 1253 2638 1279 2672
rect 1291 2638 1325 2672
rect 1325 2638 1343 2672
rect 1227 2629 1279 2638
rect 1291 2629 1343 2638
rect 1601 2558 1653 2560
rect 1601 2524 1613 2558
rect 1613 2524 1647 2558
rect 1647 2524 1653 2558
rect 1601 2508 1653 2524
rect 1601 2486 1653 2496
rect 1015 2432 1067 2484
rect 1079 2472 1131 2484
rect 1079 2438 1122 2472
rect 1122 2438 1131 2472
rect 1601 2452 1613 2486
rect 1613 2452 1647 2486
rect 1647 2452 1653 2486
rect 1601 2444 1653 2452
rect 1079 2432 1131 2438
rect 1015 2354 1067 2406
rect 1079 2400 1131 2406
rect 1079 2366 1122 2400
rect 1122 2366 1131 2400
rect 1079 2354 1131 2366
rect 845 2312 897 2321
rect 845 2278 849 2312
rect 849 2278 883 2312
rect 883 2278 897 2312
rect 845 2269 897 2278
rect 909 2312 961 2321
rect 909 2278 921 2312
rect 921 2278 955 2312
rect 955 2278 961 2312
rect 909 2269 961 2278
rect 1013 2312 1065 2321
rect 1013 2278 1019 2312
rect 1019 2278 1053 2312
rect 1053 2278 1065 2312
rect 1013 2269 1065 2278
rect 1077 2312 1129 2321
rect 1077 2278 1091 2312
rect 1091 2278 1125 2312
rect 1125 2278 1129 2312
rect 1077 2269 1129 2278
rect 1227 1793 1279 1802
rect 866 1724 918 1776
rect 1227 1759 1240 1793
rect 1240 1759 1274 1793
rect 1274 1759 1279 1793
rect 1227 1750 1279 1759
rect 1291 1750 1343 1802
rect 866 1660 918 1712
rect 1026 1684 1078 1736
rect 1600 1729 1652 1781
rect 1026 1620 1078 1672
rect 1600 1665 1652 1717
<< metal2 >>
rect 1009 4074 1015 4126
rect 1067 4074 1079 4126
rect 1131 4074 1137 4126
rect 1009 4048 1137 4074
rect 1009 3996 1015 4048
rect 1067 3996 1079 4048
rect 1131 3996 1137 4048
rect 1009 2484 1137 3996
rect 1217 3960 1269 3966
rect 1217 3896 1269 3908
rect 1217 3838 1269 3844
rect 1223 3352 1269 3838
rect 1221 3300 1227 3352
rect 1279 3300 1291 3352
rect 1343 3300 1349 3352
rect 1604 3250 1656 3256
rect 1604 3186 1656 3198
rect 1221 3111 1227 3163
rect 1279 3111 1291 3163
rect 1343 3111 1349 3163
rect 1604 3128 1656 3134
rect 1259 2681 1311 3111
rect 1221 2629 1227 2681
rect 1279 2629 1291 2681
rect 1343 2629 1349 2681
rect 1009 2432 1015 2484
rect 1067 2432 1079 2484
rect 1131 2432 1137 2484
rect 1009 2406 1137 2432
rect 1009 2354 1015 2406
rect 1067 2354 1079 2406
rect 1131 2354 1137 2406
rect 839 2269 845 2321
rect 897 2269 909 2321
rect 961 2269 967 2321
rect 1007 2269 1013 2321
rect 1065 2269 1077 2321
rect 1129 2269 1135 2321
rect 872 1782 918 2269
rect 866 1776 918 1782
rect 1054 1742 1100 2269
rect 1259 1802 1311 2629
rect 1607 2566 1653 3128
rect 1601 2560 1653 2566
rect 1601 2496 1653 2508
rect 1601 2438 1653 2444
rect 1221 1750 1227 1802
rect 1279 1750 1291 1802
rect 1343 1750 1349 1802
rect 1607 1787 1653 2438
rect 1600 1781 1653 1787
rect 866 1712 918 1724
rect 866 1654 918 1660
rect 1026 1736 1100 1742
rect 1078 1684 1100 1736
rect 1026 1672 1100 1684
rect 1078 1620 1100 1672
rect 1652 1729 1653 1781
rect 1600 1717 1653 1729
rect 1652 1685 1653 1717
rect 1600 1659 1652 1665
rect 1026 1614 1100 1620
use nfet_CDNS_52468879185512  nfet_CDNS_52468879185512_0
timestamp 1707688321
transform -1 0 1562 0 1 3128
box -79 -32 199 632
use nfet_CDNS_52468879185512  nfet_CDNS_52468879185512_1
timestamp 1707688321
transform -1 0 1254 0 1 3128
box -79 -32 199 632
use nfet_CDNS_52468879185512  nfet_CDNS_52468879185512_2
timestamp 1707688321
transform 1 0 262 0 1 2340
box -79 -32 199 632
use nfet_CDNS_52468879185793  nfet_CDNS_52468879185793_0
timestamp 1707688321
transform 1 0 141 0 -1 3706
box -79 -32 731 232
use nfet_CDNS_52468879185793  nfet_CDNS_52468879185793_1
timestamp 1707688321
transform 1 0 141 0 1 3176
box -79 -32 731 232
use nfet_CDNS_52468879185796  nfet_CDNS_52468879185796_0
timestamp 1707688321
transform 1 0 762 0 -1 2920
box -79 -32 279 182
use nfet_CDNS_52468879185796  nfet_CDNS_52468879185796_1
timestamp 1707688321
transform 1 0 1167 0 1 2440
box -79 -32 279 182
use nfet_CDNS_52468879185797  nfet_CDNS_52468879185797_0
timestamp 1707688321
transform -1 0 1333 0 -1 2920
box -79 -32 199 232
use nfet_CDNS_52468879185797  nfet_CDNS_52468879185797_1
timestamp 1707688321
transform 1 0 802 0 1 2440
box -79 -32 199 232
use nfet_CDNS_52468879185915  nfet_CDNS_52468879185915_0
timestamp 1707688321
transform 1 0 1016 0 1 3912
box -151 -32 439 232
use nfet_CDNS_52468879185915  nfet_CDNS_52468879185915_1
timestamp 1707688321
transform 1 0 247 0 1 3912
box -151 -32 439 232
use pfet_CDNS_52468879185911  pfet_CDNS_52468879185911_0
timestamp 1707688321
transform 0 1 1164 -1 0 1362
box -266 -66 219 216
use pfet_CDNS_52468879185911  pfet_CDNS_52468879185911_1
timestamp 1707688321
transform 0 1 1164 1 0 1648
box -266 -66 219 216
use pfet_CDNS_52468879185913  pfet_CDNS_52468879185913_0
timestamp 1707688321
transform -1 0 573 0 1 1201
box -266 -66 239 666
use pfet_CDNS_52468879185913  pfet_CDNS_52468879185913_1
timestamp 1707688321
transform 1 0 859 0 1 1201
box -266 -66 239 666
<< labels >>
flabel metal1 s 1409 3770 1477 3816 0 FreeSans 500 0 0 0 hld_h_n
port 2 nsew
flabel metal1 s 1152 4154 1211 4200 0 FreeSans 500 0 0 0 in
port 3 nsew
flabel metal1 s 359 4154 411 4200 0 FreeSans 500 0 0 0 in_n
port 4 nsew
flabel metal1 s 361 2988 418 3034 0 FreeSans 500 0 0 0 rst_h
port 5 nsew
flabel metal1 s 976 1435 1090 1563 0 FreeSans 500 0 0 0 vdda
port 6 nsew
flabel metal1 s 713 4016 820 4111 0 FreeSans 500 0 0 0 vssa
port 8 nsew
flabel metal1 s 553 3418 603 3464 0 FreeSans 500 0 0 0 vpwr
port 7 nsew
flabel metal2 s 1054 2178 1100 2231 0 FreeSans 500 90 0 0 out_h_n
port 9 nsew
flabel metal2 s 1281 2181 1281 2181 0 FreeSans 500 90 0 0 fbk
flabel metal2 s 1629 2180 1629 2180 0 FreeSans 500 90 0 0 fbk_n
flabel metal2 s 872 2174 918 2231 0 FreeSans 500 90 0 0 out_h
port 10 nsew
<< properties >>
string GDS_END 80698418
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 80661782
string path 31.075 95.950 31.075 99.150 
<< end >>
