magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< pwell >>
rect 1551 1747 1572 1796
<< obsli1 >>
rect 16 2216 2250 2250
rect 16 50 50 2216
rect 2216 50 2250 2216
rect 16 16 2250 50
<< obsm1 >>
rect 0 2200 2266 2266
rect 0 66 66 2200
rect 94 1164 122 2172
rect 150 1192 178 2200
rect 206 1164 234 2172
rect 262 1192 290 2200
rect 318 1164 346 2172
rect 374 1192 402 2200
rect 430 1164 458 2172
rect 486 1192 514 2200
rect 542 1164 570 2172
rect 598 1192 626 2200
rect 654 1164 682 2172
rect 710 1192 738 2200
rect 766 1164 794 2172
rect 822 1192 850 2200
rect 878 1164 906 2172
rect 934 1192 962 2200
rect 990 1164 1018 2172
rect 1046 1192 1074 2200
rect 1102 1164 1164 2172
rect 1192 1192 1220 2200
rect 1248 1164 1276 2172
rect 1304 1192 1332 2200
rect 1360 1164 1388 2172
rect 1416 1192 1444 2200
rect 1472 1164 1500 2172
rect 1528 1192 1556 2200
rect 1584 1164 1612 2172
rect 1640 1192 1668 2200
rect 1696 1164 1724 2172
rect 1752 1192 1780 2200
rect 1808 1164 1836 2172
rect 1864 1192 1892 2200
rect 1920 1164 1948 2172
rect 1976 1192 2004 2200
rect 2032 1164 2060 2172
rect 2088 1192 2116 2200
rect 2144 1164 2172 2172
rect 94 1102 2172 1164
rect 94 94 122 1102
rect 150 66 178 1074
rect 206 94 234 1102
rect 262 66 290 1074
rect 318 94 346 1102
rect 374 66 402 1074
rect 430 94 458 1102
rect 486 66 514 1074
rect 542 94 570 1102
rect 598 66 626 1074
rect 654 94 682 1102
rect 710 66 738 1074
rect 766 94 794 1102
rect 822 66 850 1074
rect 878 94 906 1102
rect 934 66 962 1074
rect 990 94 1018 1102
rect 1046 66 1074 1074
rect 1102 94 1164 1102
rect 1192 66 1220 1074
rect 1248 94 1276 1102
rect 1304 66 1332 1074
rect 1360 94 1388 1102
rect 1416 66 1444 1074
rect 1472 94 1500 1102
rect 1528 66 1556 1074
rect 1584 94 1612 1102
rect 1640 66 1668 1074
rect 1696 94 1724 1102
rect 1752 66 1780 1074
rect 1808 94 1836 1102
rect 1864 66 1892 1074
rect 1920 94 1948 1102
rect 1976 66 2004 1074
rect 2032 94 2060 1102
rect 2088 66 2116 1074
rect 2144 94 2172 1102
rect 2200 66 2266 2200
rect 0 0 2266 66
<< obsm2 >>
rect 0 2200 1074 2266
rect 1192 2200 2266 2266
rect 0 2116 66 2200
rect 1102 2172 1164 2200
rect 94 2144 2172 2172
rect 0 2088 1074 2116
rect 0 2004 66 2088
rect 1102 2060 1164 2144
rect 2200 2116 2266 2200
rect 1192 2088 2266 2116
rect 94 2032 2172 2060
rect 0 1976 1074 2004
rect 0 1892 66 1976
rect 1102 1948 1164 2032
rect 2200 2004 2266 2088
rect 1192 1976 2266 2004
rect 94 1920 2172 1948
rect 0 1864 1074 1892
rect 0 1780 66 1864
rect 1102 1836 1164 1920
rect 2200 1892 2266 1976
rect 1192 1864 2266 1892
rect 94 1808 2172 1836
rect 0 1752 1074 1780
rect 0 1668 66 1752
rect 1102 1724 1164 1808
rect 2200 1780 2266 1864
rect 1192 1752 2266 1780
rect 94 1696 2172 1724
rect 0 1640 1074 1668
rect 0 1556 66 1640
rect 1102 1612 1164 1696
rect 2200 1668 2266 1752
rect 1192 1640 2266 1668
rect 94 1584 2172 1612
rect 0 1528 1074 1556
rect 0 1444 66 1528
rect 1102 1500 1164 1584
rect 2200 1556 2266 1640
rect 1192 1528 2266 1556
rect 94 1472 2172 1500
rect 0 1416 1074 1444
rect 0 1332 66 1416
rect 1102 1388 1164 1472
rect 2200 1444 2266 1528
rect 1192 1416 2266 1444
rect 94 1360 2172 1388
rect 0 1304 1074 1332
rect 0 1220 66 1304
rect 1102 1276 1164 1360
rect 2200 1332 2266 1416
rect 1192 1304 2266 1332
rect 94 1248 2172 1276
rect 0 1192 1074 1220
rect 1102 1164 1164 1248
rect 2200 1220 2266 1304
rect 1192 1192 2266 1220
rect 66 1102 2200 1164
rect 0 1046 1074 1074
rect 0 962 66 1046
rect 1102 1018 1164 1102
rect 1192 1046 2266 1074
rect 94 990 2172 1018
rect 0 934 1074 962
rect 0 850 66 934
rect 1102 906 1164 990
rect 2200 962 2266 1046
rect 1192 934 2266 962
rect 94 878 2172 906
rect 0 822 1074 850
rect 0 738 66 822
rect 1102 794 1164 878
rect 2200 850 2266 934
rect 1192 822 2266 850
rect 94 766 2172 794
rect 0 710 1074 738
rect 0 626 66 710
rect 1102 682 1164 766
rect 2200 738 2266 822
rect 1192 710 2266 738
rect 94 654 2172 682
rect 0 598 1074 626
rect 0 514 66 598
rect 1102 570 1164 654
rect 2200 626 2266 710
rect 1192 598 2266 626
rect 94 542 2172 570
rect 0 486 1074 514
rect 0 402 66 486
rect 1102 458 1164 542
rect 2200 514 2266 598
rect 1192 486 2266 514
rect 94 430 2172 458
rect 0 374 1074 402
rect 0 290 66 374
rect 1102 346 1164 430
rect 2200 402 2266 486
rect 1192 374 2266 402
rect 94 318 2172 346
rect 0 262 1074 290
rect 0 178 66 262
rect 1102 234 1164 318
rect 2200 290 2266 374
rect 1192 262 2266 290
rect 94 206 2172 234
rect 0 150 1074 178
rect 0 66 66 150
rect 1102 122 1164 206
rect 2200 178 2266 262
rect 1192 150 2266 178
rect 94 94 2172 122
rect 1102 66 1164 94
rect 2200 66 2266 150
rect 0 0 1074 66
rect 1192 0 2266 66
<< obsm3 >>
rect 0 2200 1026 2266
rect 1240 2200 2266 2266
rect 0 1240 66 2200
rect 126 1180 186 2140
rect 246 1240 306 2200
rect 366 1180 426 2140
rect 486 1240 546 2200
rect 606 1180 666 2140
rect 726 1240 786 2200
rect 846 1180 906 2140
rect 966 1240 1026 2200
rect 1086 1180 1180 2200
rect 1240 1240 1300 2200
rect 1360 1180 1420 2140
rect 1480 1240 1540 2200
rect 1600 1180 1660 2140
rect 1720 1240 1780 2200
rect 1840 1180 1900 2140
rect 1960 1240 2020 2200
rect 2080 1180 2140 2140
rect 2200 1240 2266 2200
rect 66 1086 2200 1180
rect 0 66 66 1026
rect 126 126 186 1086
rect 246 66 306 1026
rect 366 126 426 1086
rect 486 66 546 1026
rect 606 126 666 1086
rect 726 66 786 1026
rect 846 126 906 1086
rect 966 66 1026 1026
rect 1086 66 1180 1086
rect 1240 66 1300 1026
rect 1360 126 1420 1086
rect 1480 66 1540 1026
rect 1600 126 1660 1086
rect 1720 66 1780 1026
rect 1840 126 1900 1086
rect 1960 66 2020 1026
rect 2080 126 2140 1086
rect 2200 66 2266 1026
rect 0 0 1026 66
rect 1240 0 2266 66
<< metal4 >>
rect 0 2200 2266 2266
rect 0 2020 66 2200
rect 126 2080 2140 2140
rect 0 1960 1026 2020
rect 0 1780 66 1960
rect 1086 1900 1180 2080
rect 2200 2020 2266 2200
rect 1240 1960 2266 2020
rect 126 1840 2140 1900
rect 0 1720 1026 1780
rect 0 1540 66 1720
rect 1086 1660 1180 1840
rect 2200 1780 2266 1960
rect 1240 1720 2266 1780
rect 126 1600 2140 1660
rect 0 1480 1026 1540
rect 0 1300 66 1480
rect 1086 1420 1180 1600
rect 2200 1540 2266 1720
rect 1240 1480 2266 1540
rect 126 1360 2140 1420
rect 0 1240 1026 1300
rect 0 1026 66 1240
rect 1086 1180 1180 1360
rect 2200 1300 2266 1480
rect 1240 1240 2266 1300
rect 126 1086 2140 1180
rect 0 966 1026 1026
rect 0 786 66 966
rect 1086 906 1180 1086
rect 2200 1026 2266 1240
rect 1240 966 2266 1026
rect 126 846 2140 906
rect 0 726 1026 786
rect 0 546 66 726
rect 1086 666 1180 846
rect 2200 786 2266 966
rect 1240 726 2266 786
rect 126 606 2140 666
rect 0 486 1026 546
rect 0 306 66 486
rect 1086 426 1180 606
rect 2200 546 2266 726
rect 1240 486 2266 546
rect 126 366 2140 426
rect 0 246 1026 306
rect 0 66 66 246
rect 1086 186 1180 366
rect 2200 306 2266 486
rect 1240 246 2266 306
rect 126 126 2140 186
rect 2200 66 2266 246
rect 0 0 2266 66
<< labels >>
rlabel metal4 s 2200 2020 2266 2200 6 C0
port 1 nsew
rlabel metal4 s 2200 1780 2266 1960 6 C0
port 1 nsew
rlabel metal4 s 2200 1540 2266 1720 6 C0
port 1 nsew
rlabel metal4 s 2200 1300 2266 1480 6 C0
port 1 nsew
rlabel metal4 s 2200 1026 2266 1240 6 C0
port 1 nsew
rlabel metal4 s 2200 786 2266 966 6 C0
port 1 nsew
rlabel metal4 s 2200 546 2266 726 6 C0
port 1 nsew
rlabel metal4 s 2200 306 2266 486 6 C0
port 1 nsew
rlabel metal4 s 2200 66 2266 246 6 C0
port 1 nsew
rlabel metal4 s 1240 1960 2266 2020 6 C0
port 1 nsew
rlabel metal4 s 1240 1720 2266 1780 6 C0
port 1 nsew
rlabel metal4 s 1240 1480 2266 1540 6 C0
port 1 nsew
rlabel metal4 s 1240 1240 2266 1300 6 C0
port 1 nsew
rlabel metal4 s 1240 966 2266 1026 6 C0
port 1 nsew
rlabel metal4 s 1240 726 2266 786 6 C0
port 1 nsew
rlabel metal4 s 1240 486 2266 546 6 C0
port 1 nsew
rlabel metal4 s 1240 246 2266 306 6 C0
port 1 nsew
rlabel metal4 s 0 2200 2266 2266 6 C0
port 1 nsew
rlabel metal4 s 0 2020 66 2200 6 C0
port 1 nsew
rlabel metal4 s 0 1960 1026 2020 6 C0
port 1 nsew
rlabel metal4 s 0 1780 66 1960 6 C0
port 1 nsew
rlabel metal4 s 0 1720 1026 1780 6 C0
port 1 nsew
rlabel metal4 s 0 1540 66 1720 6 C0
port 1 nsew
rlabel metal4 s 0 1480 1026 1540 6 C0
port 1 nsew
rlabel metal4 s 0 1300 66 1480 6 C0
port 1 nsew
rlabel metal4 s 0 1240 1026 1300 6 C0
port 1 nsew
rlabel metal4 s 0 1026 66 1240 6 C0
port 1 nsew
rlabel metal4 s 0 966 1026 1026 6 C0
port 1 nsew
rlabel metal4 s 0 786 66 966 6 C0
port 1 nsew
rlabel metal4 s 0 726 1026 786 6 C0
port 1 nsew
rlabel metal4 s 0 546 66 726 6 C0
port 1 nsew
rlabel metal4 s 0 486 1026 546 6 C0
port 1 nsew
rlabel metal4 s 0 306 66 486 6 C0
port 1 nsew
rlabel metal4 s 0 246 1026 306 6 C0
port 1 nsew
rlabel metal4 s 0 66 66 246 6 C0
port 1 nsew
rlabel metal4 s 0 0 2266 66 6 C0
port 1 nsew
rlabel metal4 s 1086 1900 1180 2080 6 C1
port 2 nsew
rlabel metal4 s 1086 1660 1180 1840 6 C1
port 2 nsew
rlabel metal4 s 1086 1420 1180 1600 6 C1
port 2 nsew
rlabel metal4 s 1086 1180 1180 1360 6 C1
port 2 nsew
rlabel metal4 s 1086 906 1180 1086 6 C1
port 2 nsew
rlabel metal4 s 1086 666 1180 846 6 C1
port 2 nsew
rlabel metal4 s 1086 426 1180 606 6 C1
port 2 nsew
rlabel metal4 s 1086 186 1180 366 6 C1
port 2 nsew
rlabel metal4 s 126 2080 2140 2140 6 C1
port 2 nsew
rlabel metal4 s 126 1840 2140 1900 6 C1
port 2 nsew
rlabel metal4 s 126 1600 2140 1660 6 C1
port 2 nsew
rlabel metal4 s 126 1360 2140 1420 6 C1
port 2 nsew
rlabel metal4 s 126 1086 2140 1180 6 C1
port 2 nsew
rlabel metal4 s 126 846 2140 906 6 C1
port 2 nsew
rlabel metal4 s 126 606 2140 666 6 C1
port 2 nsew
rlabel metal4 s 126 366 2140 426 6 C1
port 2 nsew
rlabel metal4 s 126 126 2140 186 6 C1
port 2 nsew
rlabel pwell s 1551 1747 1572 1796 6 SUB
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 2266 2266
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 479388
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 441852
string device primitive
<< end >>
