magic
tech sky130B
timestamp 1707688321
<< viali >>
rect 0 0 305 53
<< metal1 >>
rect -6 53 311 56
rect -6 0 0 53
rect 305 0 311 53
rect -6 -3 311 0
<< properties >>
string GDS_END 88002612
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 88001328
<< end >>
