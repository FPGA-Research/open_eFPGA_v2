magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< pwell >>
rect 74 -98 7067 -12
<< psubdiff >>
rect 100 -72 124 -38
rect 158 -72 192 -38
rect 226 -72 260 -38
rect 294 -72 328 -38
rect 362 -72 396 -38
rect 430 -72 464 -38
rect 498 -72 532 -38
rect 566 -72 600 -38
rect 634 -72 668 -38
rect 702 -72 736 -38
rect 770 -72 804 -38
rect 838 -72 872 -38
rect 906 -72 940 -38
rect 974 -72 1008 -38
rect 1042 -72 1076 -38
rect 1110 -72 1144 -38
rect 1178 -72 1212 -38
rect 1246 -72 1280 -38
rect 1314 -72 1348 -38
rect 1382 -72 1416 -38
rect 1450 -72 1484 -38
rect 1518 -72 1552 -38
rect 1586 -72 1620 -38
rect 1654 -72 1688 -38
rect 1722 -72 1756 -38
rect 1790 -72 1824 -38
rect 1858 -72 1892 -38
rect 1926 -72 1960 -38
rect 1994 -72 2028 -38
rect 2062 -72 2096 -38
rect 2130 -72 2164 -38
rect 2198 -72 2232 -38
rect 2266 -72 2300 -38
rect 2334 -72 2368 -38
rect 2402 -72 2436 -38
rect 2470 -72 2504 -38
rect 2538 -72 2572 -38
rect 2606 -72 2640 -38
rect 2674 -72 2708 -38
rect 2742 -72 2776 -38
rect 2810 -72 2844 -38
rect 2878 -72 2912 -38
rect 2946 -72 2980 -38
rect 3014 -72 3048 -38
rect 3082 -72 3116 -38
rect 3150 -72 3184 -38
rect 3218 -72 3252 -38
rect 3286 -72 3320 -38
rect 3354 -72 3388 -38
rect 3422 -72 3456 -38
rect 3490 -72 3524 -38
rect 3558 -72 3592 -38
rect 3626 -72 3660 -38
rect 3694 -72 3728 -38
rect 3762 -72 3796 -38
rect 3830 -72 3864 -38
rect 3898 -72 3932 -38
rect 3966 -72 4000 -38
rect 4034 -72 4068 -38
rect 4102 -72 4136 -38
rect 4170 -72 4204 -38
rect 4238 -72 4272 -38
rect 4306 -72 4340 -38
rect 4374 -72 4408 -38
rect 4442 -72 4476 -38
rect 4510 -72 4544 -38
rect 4578 -72 4612 -38
rect 4646 -72 4680 -38
rect 4714 -72 4748 -38
rect 4782 -72 4816 -38
rect 4850 -72 4884 -38
rect 4918 -72 4952 -38
rect 4986 -72 5020 -38
rect 5054 -72 5088 -38
rect 5122 -72 5156 -38
rect 5190 -72 5224 -38
rect 5258 -72 5292 -38
rect 5326 -72 5360 -38
rect 5394 -72 5428 -38
rect 5462 -72 5496 -38
rect 5530 -72 5564 -38
rect 5598 -72 5632 -38
rect 5666 -72 5700 -38
rect 5734 -72 5768 -38
rect 5802 -72 5836 -38
rect 5870 -72 5904 -38
rect 5938 -72 5972 -38
rect 6006 -72 6040 -38
rect 6074 -72 6108 -38
rect 6142 -72 6176 -38
rect 6210 -72 6244 -38
rect 6278 -72 6312 -38
rect 6346 -72 6380 -38
rect 6414 -72 6448 -38
rect 6482 -72 6516 -38
rect 6550 -72 6584 -38
rect 6618 -72 6652 -38
rect 6686 -72 6720 -38
rect 6754 -72 6788 -38
rect 6822 -72 6856 -38
rect 6890 -72 6924 -38
rect 6958 -72 7041 -38
<< psubdiffcont >>
rect 124 -72 158 -38
rect 192 -72 226 -38
rect 260 -72 294 -38
rect 328 -72 362 -38
rect 396 -72 430 -38
rect 464 -72 498 -38
rect 532 -72 566 -38
rect 600 -72 634 -38
rect 668 -72 702 -38
rect 736 -72 770 -38
rect 804 -72 838 -38
rect 872 -72 906 -38
rect 940 -72 974 -38
rect 1008 -72 1042 -38
rect 1076 -72 1110 -38
rect 1144 -72 1178 -38
rect 1212 -72 1246 -38
rect 1280 -72 1314 -38
rect 1348 -72 1382 -38
rect 1416 -72 1450 -38
rect 1484 -72 1518 -38
rect 1552 -72 1586 -38
rect 1620 -72 1654 -38
rect 1688 -72 1722 -38
rect 1756 -72 1790 -38
rect 1824 -72 1858 -38
rect 1892 -72 1926 -38
rect 1960 -72 1994 -38
rect 2028 -72 2062 -38
rect 2096 -72 2130 -38
rect 2164 -72 2198 -38
rect 2232 -72 2266 -38
rect 2300 -72 2334 -38
rect 2368 -72 2402 -38
rect 2436 -72 2470 -38
rect 2504 -72 2538 -38
rect 2572 -72 2606 -38
rect 2640 -72 2674 -38
rect 2708 -72 2742 -38
rect 2776 -72 2810 -38
rect 2844 -72 2878 -38
rect 2912 -72 2946 -38
rect 2980 -72 3014 -38
rect 3048 -72 3082 -38
rect 3116 -72 3150 -38
rect 3184 -72 3218 -38
rect 3252 -72 3286 -38
rect 3320 -72 3354 -38
rect 3388 -72 3422 -38
rect 3456 -72 3490 -38
rect 3524 -72 3558 -38
rect 3592 -72 3626 -38
rect 3660 -72 3694 -38
rect 3728 -72 3762 -38
rect 3796 -72 3830 -38
rect 3864 -72 3898 -38
rect 3932 -72 3966 -38
rect 4000 -72 4034 -38
rect 4068 -72 4102 -38
rect 4136 -72 4170 -38
rect 4204 -72 4238 -38
rect 4272 -72 4306 -38
rect 4340 -72 4374 -38
rect 4408 -72 4442 -38
rect 4476 -72 4510 -38
rect 4544 -72 4578 -38
rect 4612 -72 4646 -38
rect 4680 -72 4714 -38
rect 4748 -72 4782 -38
rect 4816 -72 4850 -38
rect 4884 -72 4918 -38
rect 4952 -72 4986 -38
rect 5020 -72 5054 -38
rect 5088 -72 5122 -38
rect 5156 -72 5190 -38
rect 5224 -72 5258 -38
rect 5292 -72 5326 -38
rect 5360 -72 5394 -38
rect 5428 -72 5462 -38
rect 5496 -72 5530 -38
rect 5564 -72 5598 -38
rect 5632 -72 5666 -38
rect 5700 -72 5734 -38
rect 5768 -72 5802 -38
rect 5836 -72 5870 -38
rect 5904 -72 5938 -38
rect 5972 -72 6006 -38
rect 6040 -72 6074 -38
rect 6108 -72 6142 -38
rect 6176 -72 6210 -38
rect 6244 -72 6278 -38
rect 6312 -72 6346 -38
rect 6380 -72 6414 -38
rect 6448 -72 6482 -38
rect 6516 -72 6550 -38
rect 6584 -72 6618 -38
rect 6652 -72 6686 -38
rect 6720 -72 6754 -38
rect 6788 -72 6822 -38
rect 6856 -72 6890 -38
rect 6924 -72 6958 -38
<< locali >>
rect 794 1613 847 1692
rect 1680 1620 1733 1686
rect 2566 1623 2619 1685
rect 3452 1613 3505 1698
rect 4338 1609 4391 1698
rect 5224 1618 5277 1700
rect 6110 1628 6163 1692
rect 6996 1625 7049 1684
rect 216 1517 254 1551
rect 182 324 288 1517
rect 1102 1517 1140 1551
rect 358 1431 396 1465
rect 324 324 430 1431
rect 539 1345 577 1379
rect 505 324 611 1345
rect 1068 324 1174 1517
rect 1988 1517 2026 1551
rect 1244 1431 1282 1465
rect 1210 324 1316 1431
rect 1425 1087 1463 1121
rect 1391 324 1497 1087
rect 1954 324 2060 1517
rect 2874 1517 2912 1551
rect 2311 1345 2349 1379
rect 2130 1173 2168 1207
rect 2096 324 2202 1173
rect 2277 324 2383 1345
rect 2840 324 2946 1517
rect 3902 1431 3940 1465
rect 3760 1259 3798 1293
rect 3016 1173 3054 1207
rect 2982 324 3088 1173
rect 3197 1087 3235 1121
rect 3163 324 3269 1087
rect 3726 324 3832 1259
rect 3868 324 3974 1431
rect 4788 1431 4826 1465
rect 4083 1345 4121 1379
rect 4049 324 4155 1345
rect 4646 1259 4684 1293
rect 4612 324 4718 1259
rect 4754 324 4860 1431
rect 5855 1345 5893 1379
rect 5532 1259 5570 1293
rect 4969 1087 5007 1121
rect 4935 324 5041 1087
rect 5498 324 5604 1259
rect 5674 1173 5712 1207
rect 5640 324 5746 1173
rect 5821 324 5927 1345
rect 6418 1259 6456 1293
rect 6384 324 6490 1259
rect 6560 1173 6598 1207
rect 6526 324 6632 1173
rect 6741 1087 6779 1121
rect 6707 324 6813 1087
rect 629 151 663 201
rect 629 67 663 117
rect 1515 151 1549 201
rect 1515 67 1549 117
rect 2401 151 2435 201
rect 2401 67 2435 117
rect 3287 151 3321 201
rect 3287 67 3321 117
rect 4173 151 4207 201
rect 4173 67 4207 117
rect 5059 151 5093 201
rect 5059 67 5093 117
rect 5945 151 5979 201
rect 5945 67 5979 117
rect 6831 151 6865 201
rect 6831 67 6865 117
rect 100 -72 112 -38
rect 158 -72 184 -38
rect 226 -72 256 -38
rect 294 -72 328 -38
rect 362 -72 396 -38
rect 434 -72 464 -38
rect 506 -72 532 -38
rect 578 -72 600 -38
rect 650 -72 668 -38
rect 722 -72 736 -38
rect 794 -72 804 -38
rect 866 -72 872 -38
rect 938 -72 940 -38
rect 974 -72 976 -38
rect 1042 -72 1048 -38
rect 1110 -72 1120 -38
rect 1178 -72 1192 -38
rect 1246 -72 1264 -38
rect 1314 -72 1336 -38
rect 1382 -72 1408 -38
rect 1450 -72 1480 -38
rect 1518 -72 1552 -38
rect 1586 -72 1620 -38
rect 1658 -72 1688 -38
rect 1730 -72 1756 -38
rect 1802 -72 1824 -38
rect 1874 -72 1892 -38
rect 1946 -72 1960 -38
rect 2018 -72 2028 -38
rect 2090 -72 2096 -38
rect 2162 -72 2164 -38
rect 2198 -72 2200 -38
rect 2266 -72 2272 -38
rect 2334 -72 2344 -38
rect 2402 -72 2416 -38
rect 2470 -72 2488 -38
rect 2538 -72 2560 -38
rect 2606 -72 2632 -38
rect 2674 -72 2704 -38
rect 2742 -72 2776 -38
rect 2810 -72 2844 -38
rect 2882 -72 2912 -38
rect 2954 -72 2980 -38
rect 3026 -72 3048 -38
rect 3099 -72 3116 -38
rect 3172 -72 3184 -38
rect 3245 -72 3252 -38
rect 3318 -72 3320 -38
rect 3354 -72 3357 -38
rect 3422 -72 3430 -38
rect 3490 -72 3503 -38
rect 3558 -72 3576 -38
rect 3626 -72 3649 -38
rect 3694 -72 3722 -38
rect 3762 -72 3795 -38
rect 3830 -72 3864 -38
rect 3902 -72 3932 -38
rect 3975 -72 4000 -38
rect 4048 -72 4068 -38
rect 4121 -72 4136 -38
rect 4194 -72 4204 -38
rect 4267 -72 4272 -38
rect 4374 -72 4379 -38
rect 4442 -72 4452 -38
rect 4510 -72 4525 -38
rect 4578 -72 4598 -38
rect 4646 -72 4671 -38
rect 4714 -72 4744 -38
rect 4782 -72 4816 -38
rect 4851 -72 4884 -38
rect 4924 -72 4952 -38
rect 4997 -72 5020 -38
rect 5070 -72 5088 -38
rect 5143 -72 5156 -38
rect 5216 -72 5224 -38
rect 5289 -72 5292 -38
rect 5326 -72 5328 -38
rect 5394 -72 5401 -38
rect 5462 -72 5474 -38
rect 5530 -72 5547 -38
rect 5598 -72 5620 -38
rect 5666 -72 5693 -38
rect 5734 -72 5766 -38
rect 5802 -72 5836 -38
rect 5873 -72 5904 -38
rect 5946 -72 5972 -38
rect 6019 -72 6040 -38
rect 6092 -72 6108 -38
rect 6165 -72 6176 -38
rect 6238 -72 6244 -38
rect 6311 -72 6312 -38
rect 6346 -72 6350 -38
rect 6414 -72 6423 -38
rect 6482 -72 6496 -38
rect 6550 -72 6569 -38
rect 6618 -72 6642 -38
rect 6686 -72 6715 -38
rect 6754 -72 6788 -38
rect 6822 -72 6856 -38
rect 6895 -72 6924 -38
rect 6968 -72 7007 -38
<< viali >>
rect 182 1517 216 1551
rect 254 1517 288 1551
rect 1068 1517 1102 1551
rect 1140 1517 1174 1551
rect 324 1431 358 1465
rect 396 1431 430 1465
rect 505 1345 539 1379
rect 577 1345 611 1379
rect 1954 1517 1988 1551
rect 2026 1517 2060 1551
rect 1210 1431 1244 1465
rect 1282 1431 1316 1465
rect 1391 1087 1425 1121
rect 1463 1087 1497 1121
rect 2840 1517 2874 1551
rect 2912 1517 2946 1551
rect 2277 1345 2311 1379
rect 2349 1345 2383 1379
rect 2096 1173 2130 1207
rect 2168 1173 2202 1207
rect 3868 1431 3902 1465
rect 3940 1431 3974 1465
rect 3726 1259 3760 1293
rect 3798 1259 3832 1293
rect 2982 1173 3016 1207
rect 3054 1173 3088 1207
rect 3163 1087 3197 1121
rect 3235 1087 3269 1121
rect 4754 1431 4788 1465
rect 4826 1431 4860 1465
rect 4049 1345 4083 1379
rect 4121 1345 4155 1379
rect 4612 1259 4646 1293
rect 4684 1259 4718 1293
rect 5821 1345 5855 1379
rect 5893 1345 5927 1379
rect 5498 1259 5532 1293
rect 5570 1259 5604 1293
rect 4935 1087 4969 1121
rect 5007 1087 5041 1121
rect 5640 1173 5674 1207
rect 5712 1173 5746 1207
rect 6384 1259 6418 1293
rect 6456 1259 6490 1293
rect 6526 1173 6560 1207
rect 6598 1173 6632 1207
rect 6707 1087 6741 1121
rect 6779 1087 6813 1121
rect 629 201 663 235
rect 629 117 663 151
rect 629 33 663 67
rect 1515 201 1549 235
rect 1515 117 1549 151
rect 1515 33 1549 67
rect 2401 201 2435 235
rect 2401 117 2435 151
rect 2401 33 2435 67
rect 3287 201 3321 235
rect 3287 117 3321 151
rect 3287 33 3321 67
rect 4173 201 4207 235
rect 4173 117 4207 151
rect 4173 33 4207 67
rect 5059 201 5093 235
rect 5059 117 5093 151
rect 5059 33 5093 67
rect 5945 201 5979 235
rect 5945 117 5979 151
rect 5945 33 5979 67
rect 6831 201 6865 235
rect 6831 117 6865 151
rect 6831 33 6865 67
rect 112 -72 124 -38
rect 124 -72 146 -38
rect 184 -72 192 -38
rect 192 -72 218 -38
rect 256 -72 260 -38
rect 260 -72 290 -38
rect 328 -72 362 -38
rect 400 -72 430 -38
rect 430 -72 434 -38
rect 472 -72 498 -38
rect 498 -72 506 -38
rect 544 -72 566 -38
rect 566 -72 578 -38
rect 616 -72 634 -38
rect 634 -72 650 -38
rect 688 -72 702 -38
rect 702 -72 722 -38
rect 760 -72 770 -38
rect 770 -72 794 -38
rect 832 -72 838 -38
rect 838 -72 866 -38
rect 904 -72 906 -38
rect 906 -72 938 -38
rect 976 -72 1008 -38
rect 1008 -72 1010 -38
rect 1048 -72 1076 -38
rect 1076 -72 1082 -38
rect 1120 -72 1144 -38
rect 1144 -72 1154 -38
rect 1192 -72 1212 -38
rect 1212 -72 1226 -38
rect 1264 -72 1280 -38
rect 1280 -72 1298 -38
rect 1336 -72 1348 -38
rect 1348 -72 1370 -38
rect 1408 -72 1416 -38
rect 1416 -72 1442 -38
rect 1480 -72 1484 -38
rect 1484 -72 1514 -38
rect 1552 -72 1586 -38
rect 1624 -72 1654 -38
rect 1654 -72 1658 -38
rect 1696 -72 1722 -38
rect 1722 -72 1730 -38
rect 1768 -72 1790 -38
rect 1790 -72 1802 -38
rect 1840 -72 1858 -38
rect 1858 -72 1874 -38
rect 1912 -72 1926 -38
rect 1926 -72 1946 -38
rect 1984 -72 1994 -38
rect 1994 -72 2018 -38
rect 2056 -72 2062 -38
rect 2062 -72 2090 -38
rect 2128 -72 2130 -38
rect 2130 -72 2162 -38
rect 2200 -72 2232 -38
rect 2232 -72 2234 -38
rect 2272 -72 2300 -38
rect 2300 -72 2306 -38
rect 2344 -72 2368 -38
rect 2368 -72 2378 -38
rect 2416 -72 2436 -38
rect 2436 -72 2450 -38
rect 2488 -72 2504 -38
rect 2504 -72 2522 -38
rect 2560 -72 2572 -38
rect 2572 -72 2594 -38
rect 2632 -72 2640 -38
rect 2640 -72 2666 -38
rect 2704 -72 2708 -38
rect 2708 -72 2738 -38
rect 2776 -72 2810 -38
rect 2848 -72 2878 -38
rect 2878 -72 2882 -38
rect 2920 -72 2946 -38
rect 2946 -72 2954 -38
rect 2992 -72 3014 -38
rect 3014 -72 3026 -38
rect 3065 -72 3082 -38
rect 3082 -72 3099 -38
rect 3138 -72 3150 -38
rect 3150 -72 3172 -38
rect 3211 -72 3218 -38
rect 3218 -72 3245 -38
rect 3284 -72 3286 -38
rect 3286 -72 3318 -38
rect 3357 -72 3388 -38
rect 3388 -72 3391 -38
rect 3430 -72 3456 -38
rect 3456 -72 3464 -38
rect 3503 -72 3524 -38
rect 3524 -72 3537 -38
rect 3576 -72 3592 -38
rect 3592 -72 3610 -38
rect 3649 -72 3660 -38
rect 3660 -72 3683 -38
rect 3722 -72 3728 -38
rect 3728 -72 3756 -38
rect 3795 -72 3796 -38
rect 3796 -72 3829 -38
rect 3868 -72 3898 -38
rect 3898 -72 3902 -38
rect 3941 -72 3966 -38
rect 3966 -72 3975 -38
rect 4014 -72 4034 -38
rect 4034 -72 4048 -38
rect 4087 -72 4102 -38
rect 4102 -72 4121 -38
rect 4160 -72 4170 -38
rect 4170 -72 4194 -38
rect 4233 -72 4238 -38
rect 4238 -72 4267 -38
rect 4306 -72 4340 -38
rect 4379 -72 4408 -38
rect 4408 -72 4413 -38
rect 4452 -72 4476 -38
rect 4476 -72 4486 -38
rect 4525 -72 4544 -38
rect 4544 -72 4559 -38
rect 4598 -72 4612 -38
rect 4612 -72 4632 -38
rect 4671 -72 4680 -38
rect 4680 -72 4705 -38
rect 4744 -72 4748 -38
rect 4748 -72 4778 -38
rect 4817 -72 4850 -38
rect 4850 -72 4851 -38
rect 4890 -72 4918 -38
rect 4918 -72 4924 -38
rect 4963 -72 4986 -38
rect 4986 -72 4997 -38
rect 5036 -72 5054 -38
rect 5054 -72 5070 -38
rect 5109 -72 5122 -38
rect 5122 -72 5143 -38
rect 5182 -72 5190 -38
rect 5190 -72 5216 -38
rect 5255 -72 5258 -38
rect 5258 -72 5289 -38
rect 5328 -72 5360 -38
rect 5360 -72 5362 -38
rect 5401 -72 5428 -38
rect 5428 -72 5435 -38
rect 5474 -72 5496 -38
rect 5496 -72 5508 -38
rect 5547 -72 5564 -38
rect 5564 -72 5581 -38
rect 5620 -72 5632 -38
rect 5632 -72 5654 -38
rect 5693 -72 5700 -38
rect 5700 -72 5727 -38
rect 5766 -72 5768 -38
rect 5768 -72 5800 -38
rect 5839 -72 5870 -38
rect 5870 -72 5873 -38
rect 5912 -72 5938 -38
rect 5938 -72 5946 -38
rect 5985 -72 6006 -38
rect 6006 -72 6019 -38
rect 6058 -72 6074 -38
rect 6074 -72 6092 -38
rect 6131 -72 6142 -38
rect 6142 -72 6165 -38
rect 6204 -72 6210 -38
rect 6210 -72 6238 -38
rect 6277 -72 6278 -38
rect 6278 -72 6311 -38
rect 6350 -72 6380 -38
rect 6380 -72 6384 -38
rect 6423 -72 6448 -38
rect 6448 -72 6457 -38
rect 6496 -72 6516 -38
rect 6516 -72 6530 -38
rect 6569 -72 6584 -38
rect 6584 -72 6603 -38
rect 6642 -72 6652 -38
rect 6652 -72 6676 -38
rect 6715 -72 6720 -38
rect 6720 -72 6749 -38
rect 6788 -72 6822 -38
rect 6861 -72 6890 -38
rect 6890 -72 6895 -38
rect 6934 -72 6958 -38
rect 6958 -72 6968 -38
rect 7007 -72 7041 -38
<< metal1 >>
rect 6720 1886 6808 1957
rect 35 1551 7100 1557
rect 35 1517 182 1551
rect 216 1517 254 1551
rect 288 1517 1068 1551
rect 1102 1517 1140 1551
rect 1174 1517 1954 1551
rect 1988 1517 2026 1551
rect 2060 1517 2840 1551
rect 2874 1517 2912 1551
rect 2946 1517 7100 1551
rect 35 1511 7100 1517
rect 35 1465 7100 1471
rect 35 1431 324 1465
rect 358 1431 396 1465
rect 430 1431 1210 1465
rect 1244 1431 1282 1465
rect 1316 1431 3868 1465
rect 3902 1431 3940 1465
rect 3974 1431 4754 1465
rect 4788 1431 4826 1465
rect 4860 1431 7100 1465
rect 35 1425 7100 1431
rect 35 1379 7100 1385
rect 35 1345 505 1379
rect 539 1345 577 1379
rect 611 1345 2277 1379
rect 2311 1345 2349 1379
rect 2383 1345 4049 1379
rect 4083 1345 4121 1379
rect 4155 1345 5821 1379
rect 5855 1345 5893 1379
rect 5927 1345 7100 1379
rect 35 1339 7100 1345
rect 35 1293 7100 1299
rect 35 1259 3726 1293
rect 3760 1259 3798 1293
rect 3832 1259 4612 1293
rect 4646 1259 4684 1293
rect 4718 1259 5498 1293
rect 5532 1259 5570 1293
rect 5604 1259 6384 1293
rect 6418 1259 6456 1293
rect 6490 1259 7100 1293
rect 35 1253 7100 1259
rect 35 1207 7100 1213
rect 35 1173 2096 1207
rect 2130 1173 2168 1207
rect 2202 1173 2982 1207
rect 3016 1173 3054 1207
rect 3088 1173 5640 1207
rect 5674 1173 5712 1207
rect 5746 1173 6526 1207
rect 6560 1173 6598 1207
rect 6632 1173 7100 1207
rect 35 1167 7100 1173
rect 35 1121 7100 1127
rect 35 1087 1391 1121
rect 1425 1087 1463 1121
rect 1497 1087 3163 1121
rect 3197 1087 3235 1121
rect 3269 1087 4935 1121
rect 4969 1087 5007 1121
rect 5041 1087 6707 1121
rect 6741 1087 6779 1121
rect 6813 1087 7100 1121
rect 35 1081 7100 1087
rect 27 235 7115 247
rect 27 201 629 235
rect 663 201 1515 235
rect 1549 201 2401 235
rect 2435 201 3287 235
rect 3321 201 4173 235
rect 4207 201 5059 235
rect 5093 201 5945 235
rect 5979 201 6831 235
rect 6865 201 7115 235
rect 27 151 7115 201
rect 27 117 629 151
rect 663 117 1515 151
rect 1549 117 2401 151
rect 2435 117 3287 151
rect 3321 117 4173 151
rect 4207 117 5059 151
rect 5093 117 5945 151
rect 5979 117 6831 151
rect 6865 117 7115 151
rect 27 67 7115 117
rect 27 33 629 67
rect 663 33 1515 67
rect 1549 33 2401 67
rect 2435 33 3287 67
rect 3321 33 4173 67
rect 4207 33 5059 67
rect 5093 33 5945 67
rect 5979 33 6831 67
rect 6865 33 7115 67
rect 27 21 7115 33
rect 100 -38 7053 21
rect 100 -72 112 -38
rect 146 -72 184 -38
rect 218 -72 256 -38
rect 290 -72 328 -38
rect 362 -72 400 -38
rect 434 -72 472 -38
rect 506 -72 544 -38
rect 578 -72 616 -38
rect 650 -72 688 -38
rect 722 -72 760 -38
rect 794 -72 832 -38
rect 866 -72 904 -38
rect 938 -72 976 -38
rect 1010 -72 1048 -38
rect 1082 -72 1120 -38
rect 1154 -72 1192 -38
rect 1226 -72 1264 -38
rect 1298 -72 1336 -38
rect 1370 -72 1408 -38
rect 1442 -72 1480 -38
rect 1514 -72 1552 -38
rect 1586 -72 1624 -38
rect 1658 -72 1696 -38
rect 1730 -72 1768 -38
rect 1802 -72 1840 -38
rect 1874 -72 1912 -38
rect 1946 -72 1984 -38
rect 2018 -72 2056 -38
rect 2090 -72 2128 -38
rect 2162 -72 2200 -38
rect 2234 -72 2272 -38
rect 2306 -72 2344 -38
rect 2378 -72 2416 -38
rect 2450 -72 2488 -38
rect 2522 -72 2560 -38
rect 2594 -72 2632 -38
rect 2666 -72 2704 -38
rect 2738 -72 2776 -38
rect 2810 -72 2848 -38
rect 2882 -72 2920 -38
rect 2954 -72 2992 -38
rect 3026 -72 3065 -38
rect 3099 -72 3138 -38
rect 3172 -72 3211 -38
rect 3245 -72 3284 -38
rect 3318 -72 3357 -38
rect 3391 -72 3430 -38
rect 3464 -72 3503 -38
rect 3537 -72 3576 -38
rect 3610 -72 3649 -38
rect 3683 -72 3722 -38
rect 3756 -72 3795 -38
rect 3829 -72 3868 -38
rect 3902 -72 3941 -38
rect 3975 -72 4014 -38
rect 4048 -72 4087 -38
rect 4121 -72 4160 -38
rect 4194 -72 4233 -38
rect 4267 -72 4306 -38
rect 4340 -72 4379 -38
rect 4413 -72 4452 -38
rect 4486 -72 4525 -38
rect 4559 -72 4598 -38
rect 4632 -72 4671 -38
rect 4705 -72 4744 -38
rect 4778 -72 4817 -38
rect 4851 -72 4890 -38
rect 4924 -72 4963 -38
rect 4997 -72 5036 -38
rect 5070 -72 5109 -38
rect 5143 -72 5182 -38
rect 5216 -72 5255 -38
rect 5289 -72 5328 -38
rect 5362 -72 5401 -38
rect 5435 -72 5474 -38
rect 5508 -72 5547 -38
rect 5581 -72 5620 -38
rect 5654 -72 5693 -38
rect 5727 -72 5766 -38
rect 5800 -72 5839 -38
rect 5873 -72 5912 -38
rect 5946 -72 5985 -38
rect 6019 -72 6058 -38
rect 6092 -72 6131 -38
rect 6165 -72 6204 -38
rect 6238 -72 6277 -38
rect 6311 -72 6350 -38
rect 6384 -72 6423 -38
rect 6457 -72 6496 -38
rect 6530 -72 6569 -38
rect 6603 -72 6642 -38
rect 6676 -72 6715 -38
rect 6749 -72 6788 -38
rect 6822 -72 6861 -38
rect 6895 -72 6934 -38
rect 6968 -72 7007 -38
rect 7041 -72 7053 -38
rect 100 -78 7053 -72
use sky130_fd_io__refgen_mux_and3  sky130_fd_io__refgen_mux_and3_0
timestamp 1707688321
transform 1 0 2685 0 1 -8
box 0 13 886 2173
use sky130_fd_io__refgen_mux_and3  sky130_fd_io__refgen_mux_and3_1
timestamp 1707688321
transform 1 0 27 0 1 -8
box 0 13 886 2173
use sky130_fd_io__refgen_mux_and3  sky130_fd_io__refgen_mux_and3_2
timestamp 1707688321
transform 1 0 4457 0 1 -8
box 0 13 886 2173
use sky130_fd_io__refgen_mux_and3  sky130_fd_io__refgen_mux_and3_3
timestamp 1707688321
transform 1 0 6229 0 1 -8
box 0 13 886 2173
use sky130_fd_io__refgen_mux_and3  sky130_fd_io__refgen_mux_and3_4
timestamp 1707688321
transform 1 0 3571 0 1 -8
box 0 13 886 2173
use sky130_fd_io__refgen_mux_and3  sky130_fd_io__refgen_mux_and3_5
timestamp 1707688321
transform 1 0 5343 0 1 -8
box 0 13 886 2173
use sky130_fd_io__refgen_mux_and3  sky130_fd_io__refgen_mux_and3_6
timestamp 1707688321
transform 1 0 913 0 1 -8
box 0 13 886 2173
use sky130_fd_io__refgen_mux_and3  sky130_fd_io__refgen_mux_and3_7
timestamp 1707688321
transform 1 0 1799 0 1 -8
box 0 13 886 2173
<< labels >>
flabel metal1 s 6187 1253 6257 1299 0 FreeSans 500 0 0 0 voh_sel_h<2>
port 3 nsew
flabel metal1 s 6187 1167 6257 1213 0 FreeSans 500 0 0 0 voh_sel_h<1>
port 5 nsew
flabel metal1 s 6187 1425 6257 1471 0 FreeSans 500 0 0 0 voh_sel_h_n<1>
port 4 nsew
flabel metal1 s 6187 1511 6257 1557 0 FreeSans 500 0 0 0 voh_sel_h_n<2>
port 8 nsew
flabel metal1 s 6187 1081 6257 1127 0 FreeSans 500 0 0 0 voh_sel_h<0>
port 1 nsew
flabel metal1 s 6720 1886 6808 1957 0 FreeSans 500 0 0 0 vddio
port 6 nsew
flabel metal1 s 6557 90 6641 179 0 FreeSans 500 0 0 0 vssio
port 7 nsew
flabel metal1 s 6187 1339 6257 1385 0 FreeSans 500 0 0 0 voh_sel_h_n<0>
port 2 nsew
flabel locali s 2566 1623 2619 1685 0 FreeSans 500 90 0 0 sel<2>
port 10 nsew
flabel locali s 3452 1613 3505 1698 0 FreeSans 500 90 0 0 sel<3>
port 11 nsew
flabel locali s 4338 1609 4391 1698 0 FreeSans 500 90 0 0 sel<4>
port 12 nsew
flabel locali s 6996 1625 7049 1684 0 FreeSans 500 90 0 0 sel<7>
port 13 nsew
flabel locali s 5224 1618 5277 1700 0 FreeSans 500 90 0 0 sel<5>
port 14 nsew
flabel locali s 6110 1628 6163 1692 0 FreeSans 500 90 0 0 sel<6>
port 15 nsew
flabel locali s 794 1613 847 1692 0 FreeSans 500 90 0 0 sel<0>
port 16 nsew
flabel locali s 1680 1620 1733 1686 0 FreeSans 500 90 0 0 sel<1>
port 17 nsew
<< properties >>
string GDS_END 80640712
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 80615068
string path 2.500 -1.375 176.025 -1.375 
<< end >>
