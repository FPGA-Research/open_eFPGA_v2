magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -82 -26 182 176
<< mvnmos >>
rect 0 0 100 150
<< mvndiff >>
rect -56 114 0 150
rect -56 80 -45 114
rect -11 80 0 114
rect -56 46 0 80
rect -56 12 -45 46
rect -11 12 0 46
rect -56 0 0 12
rect 100 114 156 150
rect 100 80 111 114
rect 145 80 156 114
rect 100 46 156 80
rect 100 12 111 46
rect 145 12 156 46
rect 100 0 156 12
<< mvndiffc >>
rect -45 80 -11 114
rect -45 12 -11 46
rect 111 80 145 114
rect 111 12 145 46
<< poly >>
rect 0 150 100 182
rect 0 -32 100 0
<< locali >>
rect -45 114 -11 130
rect -45 46 -11 68
rect 111 114 145 130
rect 111 46 145 68
<< viali >>
rect -45 80 -11 102
rect -45 68 -11 80
rect -45 12 -11 30
rect -45 -4 -11 12
rect 111 80 145 102
rect 111 68 145 80
rect 111 12 145 30
rect 111 -4 145 12
<< metal1 >>
rect -51 102 -5 114
rect -51 68 -45 102
rect -11 68 -5 102
rect -51 30 -5 68
rect -51 -4 -45 30
rect -11 -4 -5 30
rect -51 -16 -5 -4
rect 105 102 151 114
rect 105 68 111 102
rect 145 68 151 102
rect 105 30 151 68
rect 105 -4 111 30
rect 145 -4 151 30
rect 105 -16 151 -4
use hvDFM1sd2_CDNS_52468879185875  hvDFM1sd2_CDNS_52468879185875_0
timestamp 1707688321
transform -1 0 0 0 1 0
box 0 0 1 1
use hvDFM1sd2_CDNS_52468879185875  hvDFM1sd2_CDNS_52468879185875_1
timestamp 1707688321
transform 1 0 100 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 49 -28 49 0 FreeSans 300 0 0 0 S
flabel comment s 128 49 128 49 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 7609318
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7608424
<< end >>
