magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -116 -66 216 666
<< mvpmos >>
rect 0 0 100 600
<< mvpdiff >>
rect -50 0 0 600
rect 100 0 150 600
<< poly >>
rect 0 600 100 626
rect 0 -26 100 0
<< labels >>
flabel comment s -25 300 -25 300 0 FreeSans 300 0 0 0 S
flabel comment s 125 300 125 300 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 87874490
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87873722
<< end >>
