magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -38 261 1786 582
<< pwell >>
rect 704 157 886 201
rect 1194 157 1747 203
rect 1 21 1747 157
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 351 47 381 131
rect 463 47 493 119
rect 562 47 592 119
rect 661 47 691 131
rect 780 47 810 175
rect 881 47 911 119
rect 987 47 1017 119
rect 1082 47 1112 131
rect 1272 47 1302 177
rect 1356 47 1386 177
rect 1544 47 1574 131
rect 1639 47 1669 177
<< scpmoshvt >>
rect 79 363 109 491
rect 163 363 193 491
rect 351 413 381 497
rect 436 413 466 497
rect 531 413 561 497
rect 634 413 664 497
rect 766 347 796 497
rect 861 413 891 497
rect 945 413 975 497
rect 1059 413 1089 497
rect 1270 297 1300 497
rect 1354 297 1384 497
rect 1542 369 1572 497
rect 1639 297 1669 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 299 93 351 131
rect 299 59 307 93
rect 341 59 351 93
rect 299 47 351 59
rect 381 119 431 131
rect 730 131 780 175
rect 611 119 661 131
rect 381 107 463 119
rect 381 73 392 107
rect 426 73 463 107
rect 381 47 463 73
rect 493 107 562 119
rect 493 73 503 107
rect 537 73 562 107
rect 493 47 562 73
rect 592 47 661 119
rect 691 101 780 131
rect 691 67 702 101
rect 736 67 780 101
rect 691 47 780 67
rect 810 119 860 175
rect 1220 162 1272 177
rect 1032 119 1082 131
rect 810 107 881 119
rect 810 73 821 107
rect 855 73 881 107
rect 810 47 881 73
rect 911 107 987 119
rect 911 73 924 107
rect 958 73 987 107
rect 911 47 987 73
rect 1017 47 1082 119
rect 1112 107 1164 131
rect 1112 73 1122 107
rect 1156 73 1164 107
rect 1112 47 1164 73
rect 1220 128 1228 162
rect 1262 128 1272 162
rect 1220 94 1272 128
rect 1220 60 1228 94
rect 1262 60 1272 94
rect 1220 47 1272 60
rect 1302 123 1356 177
rect 1302 89 1312 123
rect 1346 89 1356 123
rect 1302 47 1356 89
rect 1386 164 1438 177
rect 1386 130 1396 164
rect 1430 130 1438 164
rect 1589 131 1639 177
rect 1386 96 1438 130
rect 1386 62 1396 96
rect 1430 62 1438 96
rect 1386 47 1438 62
rect 1492 119 1544 131
rect 1492 85 1500 119
rect 1534 85 1544 119
rect 1492 47 1544 85
rect 1574 93 1639 131
rect 1574 59 1595 93
rect 1629 59 1639 93
rect 1574 47 1639 59
rect 1669 131 1721 177
rect 1669 97 1679 131
rect 1713 97 1721 131
rect 1669 47 1721 97
<< pdiff >>
rect 27 477 79 491
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 363 79 375
rect 109 461 163 491
rect 109 427 119 461
rect 153 427 163 461
rect 109 363 163 427
rect 193 477 245 491
rect 193 443 203 477
rect 237 443 245 477
rect 193 409 245 443
rect 299 485 351 497
rect 299 451 307 485
rect 341 451 351 485
rect 299 413 351 451
rect 381 477 436 497
rect 381 443 391 477
rect 425 443 436 477
rect 381 413 436 443
rect 466 472 531 497
rect 466 438 483 472
rect 517 438 531 472
rect 466 413 531 438
rect 561 413 634 497
rect 664 485 766 497
rect 664 451 722 485
rect 756 451 766 485
rect 664 417 766 451
rect 664 413 722 417
rect 193 375 203 409
rect 237 375 245 409
rect 193 363 245 375
rect 679 383 722 413
rect 756 383 766 417
rect 679 347 766 383
rect 796 477 861 497
rect 796 443 806 477
rect 840 443 861 477
rect 796 413 861 443
rect 891 467 945 497
rect 891 433 901 467
rect 935 433 945 467
rect 891 413 945 433
rect 975 413 1059 497
rect 1089 477 1142 497
rect 1089 443 1100 477
rect 1134 443 1142 477
rect 1089 413 1142 443
rect 1216 485 1270 497
rect 1216 451 1224 485
rect 1258 451 1270 485
rect 1216 414 1270 451
rect 796 347 846 413
rect 1216 380 1224 414
rect 1258 380 1270 414
rect 1216 343 1270 380
rect 1216 309 1224 343
rect 1258 309 1270 343
rect 1216 297 1270 309
rect 1300 455 1354 497
rect 1300 421 1310 455
rect 1344 421 1354 455
rect 1300 375 1354 421
rect 1300 341 1310 375
rect 1344 341 1354 375
rect 1300 297 1354 341
rect 1384 479 1436 497
rect 1384 445 1394 479
rect 1428 445 1436 479
rect 1384 411 1436 445
rect 1384 377 1394 411
rect 1428 377 1436 411
rect 1384 343 1436 377
rect 1490 485 1542 497
rect 1490 451 1498 485
rect 1532 451 1542 485
rect 1490 417 1542 451
rect 1490 383 1498 417
rect 1532 383 1542 417
rect 1490 369 1542 383
rect 1572 485 1639 497
rect 1572 451 1595 485
rect 1629 451 1639 485
rect 1572 417 1639 451
rect 1572 383 1595 417
rect 1629 383 1639 417
rect 1572 369 1639 383
rect 1384 309 1394 343
rect 1428 309 1436 343
rect 1384 297 1436 309
rect 1587 349 1639 369
rect 1587 315 1595 349
rect 1629 315 1639 349
rect 1587 297 1639 315
rect 1669 485 1721 497
rect 1669 451 1679 485
rect 1713 451 1721 485
rect 1669 414 1721 451
rect 1669 380 1679 414
rect 1713 380 1721 414
rect 1669 343 1721 380
rect 1669 309 1679 343
rect 1713 309 1721 343
rect 1669 297 1721 309
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 307 59 341 93
rect 392 73 426 107
rect 503 73 537 107
rect 702 67 736 101
rect 821 73 855 107
rect 924 73 958 107
rect 1122 73 1156 107
rect 1228 128 1262 162
rect 1228 60 1262 94
rect 1312 89 1346 123
rect 1396 130 1430 164
rect 1396 62 1430 96
rect 1500 85 1534 119
rect 1595 59 1629 93
rect 1679 97 1713 131
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 427 153 461
rect 203 443 237 477
rect 307 451 341 485
rect 391 443 425 477
rect 483 438 517 472
rect 722 451 756 485
rect 203 375 237 409
rect 722 383 756 417
rect 806 443 840 477
rect 901 433 935 467
rect 1100 443 1134 477
rect 1224 451 1258 485
rect 1224 380 1258 414
rect 1224 309 1258 343
rect 1310 421 1344 455
rect 1310 341 1344 375
rect 1394 445 1428 479
rect 1394 377 1428 411
rect 1498 451 1532 485
rect 1498 383 1532 417
rect 1595 451 1629 485
rect 1595 383 1629 417
rect 1394 309 1428 343
rect 1595 315 1629 349
rect 1679 451 1713 485
rect 1679 380 1713 414
rect 1679 309 1713 343
<< poly >>
rect 79 491 109 517
rect 163 491 193 517
rect 351 497 381 523
rect 436 497 466 523
rect 531 497 561 523
rect 634 497 664 523
rect 766 497 796 523
rect 861 497 891 523
rect 945 497 975 523
rect 1059 497 1089 523
rect 1270 497 1300 523
rect 1354 497 1384 523
rect 1542 497 1572 523
rect 1639 497 1669 523
rect 79 348 109 363
rect 46 318 109 348
rect 46 265 76 318
rect 163 274 193 363
rect 351 333 381 413
rect 22 249 76 265
rect 22 215 32 249
rect 66 215 76 249
rect 118 264 193 274
rect 286 317 381 333
rect 286 283 296 317
rect 330 283 381 317
rect 436 297 466 413
rect 531 381 561 413
rect 531 365 592 381
rect 531 331 548 365
rect 582 331 592 365
rect 531 315 592 331
rect 286 267 381 283
rect 118 230 134 264
rect 168 230 193 264
rect 118 220 193 230
rect 22 199 76 215
rect 46 176 76 199
rect 46 146 109 176
rect 79 131 109 146
rect 163 131 193 220
rect 351 131 381 267
rect 423 287 489 297
rect 423 253 439 287
rect 473 273 489 287
rect 473 253 592 273
rect 423 243 592 253
rect 443 191 509 201
rect 443 157 459 191
rect 493 157 509 191
rect 443 147 509 157
rect 463 119 493 147
rect 562 119 592 243
rect 634 213 664 413
rect 766 309 796 347
rect 861 315 891 413
rect 945 375 975 413
rect 1059 381 1089 413
rect 944 365 1010 375
rect 944 331 960 365
rect 994 331 1010 365
rect 944 321 1010 331
rect 1059 365 1140 381
rect 1059 331 1096 365
rect 1130 331 1140 365
rect 1059 315 1140 331
rect 706 299 796 309
rect 706 265 722 299
rect 756 265 796 299
rect 706 255 796 265
rect 766 220 796 255
rect 848 299 902 315
rect 848 265 858 299
rect 892 279 902 299
rect 892 265 1017 279
rect 848 249 1017 265
rect 634 203 708 213
rect 634 169 658 203
rect 692 169 708 203
rect 766 190 810 220
rect 780 175 810 190
rect 881 191 945 207
rect 634 159 708 169
rect 661 131 691 159
rect 881 157 901 191
rect 935 157 945 191
rect 881 141 945 157
rect 881 119 911 141
rect 987 119 1017 249
rect 1082 131 1112 315
rect 1542 333 1572 369
rect 1533 303 1572 333
rect 1270 265 1300 297
rect 1354 265 1384 297
rect 1533 265 1563 303
rect 1639 265 1669 297
rect 1160 249 1302 265
rect 1160 215 1170 249
rect 1204 215 1302 249
rect 1160 199 1302 215
rect 1344 249 1563 265
rect 1344 215 1354 249
rect 1388 215 1563 249
rect 1344 199 1563 215
rect 1605 249 1669 265
rect 1605 215 1615 249
rect 1649 215 1669 249
rect 1605 199 1669 215
rect 1272 177 1302 199
rect 1356 177 1386 199
rect 1533 170 1563 199
rect 1639 177 1669 199
rect 1533 146 1574 170
rect 1544 131 1574 146
rect 79 21 109 47
rect 163 21 193 47
rect 351 21 381 47
rect 463 21 493 47
rect 562 21 592 47
rect 661 21 691 47
rect 780 21 810 47
rect 881 21 911 47
rect 987 21 1017 47
rect 1082 21 1112 47
rect 1272 21 1302 47
rect 1356 21 1386 47
rect 1544 21 1574 47
rect 1639 21 1669 47
<< polycont >>
rect 32 215 66 249
rect 296 283 330 317
rect 548 331 582 365
rect 134 230 168 264
rect 439 253 473 287
rect 459 157 493 191
rect 960 331 994 365
rect 1096 331 1130 365
rect 722 265 756 299
rect 858 265 892 299
rect 658 169 692 203
rect 901 157 935 191
rect 1170 215 1204 249
rect 1354 215 1388 249
rect 1615 215 1649 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 35 477 69 493
rect 35 409 69 443
rect 103 461 169 527
rect 103 427 119 461
rect 153 427 169 461
rect 203 477 240 493
rect 237 443 240 477
rect 203 409 240 443
rect 288 485 341 527
rect 288 451 307 485
rect 288 435 341 451
rect 375 477 425 493
rect 375 443 391 477
rect 722 485 756 527
rect 69 391 168 393
rect 69 375 126 391
rect 35 359 126 375
rect 122 357 126 359
rect 160 357 168 391
rect 18 249 88 325
rect 18 215 32 249
rect 66 215 88 249
rect 18 195 88 215
rect 122 264 168 357
rect 122 230 134 264
rect 122 161 168 230
rect 35 127 168 161
rect 237 375 240 409
rect 375 408 425 443
rect 467 438 483 472
rect 517 438 688 472
rect 203 323 240 375
rect 364 382 425 408
rect 514 391 620 404
rect 203 289 205 323
rect 239 289 240 323
rect 35 119 69 127
rect 203 119 240 289
rect 274 317 330 333
rect 274 283 296 317
rect 274 143 330 283
rect 364 161 398 382
rect 514 357 546 391
rect 580 365 620 391
rect 432 323 480 344
rect 432 289 443 323
rect 477 289 480 323
rect 432 287 480 289
rect 432 253 439 287
rect 473 253 480 287
rect 432 225 480 253
rect 514 191 548 357
rect 582 331 620 365
rect 654 315 688 438
rect 722 417 756 451
rect 722 367 756 383
rect 790 477 840 493
rect 790 443 806 477
rect 1098 477 1161 527
rect 790 427 840 443
rect 885 433 901 467
rect 935 433 1062 467
rect 654 299 756 315
rect 654 297 722 299
rect 364 135 409 161
rect 443 157 459 191
rect 493 157 548 191
rect 443 147 548 157
rect 582 265 722 297
rect 582 263 756 265
rect 35 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 237 85 240 119
rect 203 69 240 85
rect 291 93 341 109
rect 103 17 169 59
rect 291 59 307 93
rect 375 107 409 135
rect 582 107 616 263
rect 722 249 756 263
rect 658 213 698 219
rect 790 213 824 427
rect 858 391 896 393
rect 858 357 860 391
rect 894 357 896 391
rect 858 299 896 357
rect 892 265 896 299
rect 858 249 896 265
rect 930 365 994 399
rect 930 331 960 365
rect 930 323 994 331
rect 930 289 947 323
rect 981 289 994 323
rect 658 203 824 213
rect 930 207 994 289
rect 692 169 824 203
rect 658 153 824 169
rect 375 73 392 107
rect 426 73 442 107
rect 481 73 503 107
rect 537 73 616 107
rect 680 101 754 117
rect 291 17 341 59
rect 680 67 702 101
rect 736 67 754 101
rect 790 107 824 153
rect 901 191 994 207
rect 935 157 994 191
rect 901 141 994 157
rect 1028 265 1062 433
rect 1098 443 1100 477
rect 1134 443 1161 477
rect 1098 427 1161 443
rect 1208 485 1276 493
rect 1208 451 1224 485
rect 1258 451 1276 485
rect 1208 414 1276 451
rect 1208 381 1224 414
rect 1096 380 1224 381
rect 1258 380 1276 414
rect 1096 365 1276 380
rect 1130 343 1276 365
rect 1130 331 1224 343
rect 1096 309 1224 331
rect 1258 309 1276 343
rect 1310 455 1344 527
rect 1482 485 1548 489
rect 1310 375 1344 421
rect 1310 325 1344 341
rect 1378 479 1444 484
rect 1378 445 1394 479
rect 1428 445 1444 479
rect 1378 411 1444 445
rect 1378 377 1394 411
rect 1428 377 1444 411
rect 1378 343 1444 377
rect 1482 451 1498 485
rect 1532 451 1548 485
rect 1482 417 1548 451
rect 1482 383 1498 417
rect 1532 383 1548 417
rect 1482 343 1548 383
rect 1096 306 1276 309
rect 1238 265 1276 306
rect 1378 309 1394 343
rect 1428 315 1444 343
rect 1428 309 1460 315
rect 1378 299 1460 309
rect 1413 289 1460 299
rect 1028 249 1204 265
rect 1028 215 1170 249
rect 1028 199 1204 215
rect 1238 249 1388 265
rect 1238 215 1354 249
rect 1238 199 1388 215
rect 1028 107 1062 199
rect 1238 165 1278 199
rect 1422 173 1460 289
rect 1411 165 1460 173
rect 1212 162 1278 165
rect 1212 128 1228 162
rect 1262 128 1278 162
rect 1380 164 1460 165
rect 790 73 821 107
rect 855 73 871 107
rect 905 73 924 107
rect 958 73 1062 107
rect 1117 107 1159 123
rect 1117 73 1122 107
rect 1156 73 1159 107
rect 680 17 754 67
rect 1117 17 1159 73
rect 1212 94 1278 128
rect 1212 60 1228 94
rect 1262 60 1278 94
rect 1312 123 1346 139
rect 1312 17 1346 89
rect 1380 130 1396 164
rect 1430 148 1460 164
rect 1494 265 1548 343
rect 1586 485 1629 527
rect 1586 451 1595 485
rect 1586 417 1629 451
rect 1586 383 1595 417
rect 1586 349 1629 383
rect 1586 315 1595 349
rect 1586 299 1629 315
rect 1663 485 1730 493
rect 1663 451 1679 485
rect 1713 451 1730 485
rect 1663 414 1730 451
rect 1663 380 1679 414
rect 1713 380 1730 414
rect 1663 343 1730 380
rect 1663 309 1679 343
rect 1713 309 1730 343
rect 1663 296 1730 309
rect 1494 249 1649 265
rect 1494 215 1615 249
rect 1494 199 1649 215
rect 1430 130 1446 148
rect 1380 96 1446 130
rect 1494 123 1534 199
rect 1683 182 1730 296
rect 1380 62 1396 96
rect 1430 62 1446 96
rect 1484 119 1534 123
rect 1484 85 1500 119
rect 1679 131 1730 182
rect 1484 69 1534 85
rect 1581 93 1645 109
rect 1380 61 1446 62
rect 1581 59 1595 93
rect 1629 59 1645 93
rect 1581 17 1645 59
rect 1713 97 1730 131
rect 1679 51 1730 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 126 357 160 391
rect 205 289 239 323
rect 546 365 580 391
rect 546 357 548 365
rect 548 357 580 365
rect 443 289 477 323
rect 860 357 894 391
rect 947 289 981 323
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
<< metal1 >>
rect 0 561 1748 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 0 496 1748 527
rect 114 391 172 397
rect 114 357 126 391
rect 160 388 172 391
rect 534 391 592 397
rect 534 388 546 391
rect 160 360 546 388
rect 160 357 172 360
rect 114 351 172 357
rect 534 357 546 360
rect 580 388 592 391
rect 848 391 906 397
rect 848 388 860 391
rect 580 360 860 388
rect 580 357 592 360
rect 534 351 592 357
rect 848 357 860 360
rect 894 357 906 391
rect 848 351 906 357
rect 193 323 251 329
rect 193 289 205 323
rect 239 320 251 323
rect 431 323 489 329
rect 431 320 443 323
rect 239 292 443 320
rect 239 289 251 292
rect 193 283 251 289
rect 431 289 443 292
rect 477 320 489 323
rect 935 323 993 329
rect 935 320 947 323
rect 477 292 947 320
rect 477 289 489 292
rect 431 283 489 289
rect 935 289 947 292
rect 981 289 993 323
rect 935 283 993 289
rect 0 17 1748 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
rect 0 -48 1748 -17
<< labels >>
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel locali s 1685 304 1719 338 0 FreeSans 400 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 289 221 323 255 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 29 221 63 255 0 FreeSans 400 0 0 0 CLK
port 1 nsew clock input
flabel locali s 1390 85 1424 119 0 FreeSans 400 0 0 0 Q
port 7 nsew signal output
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
rlabel comment s 0 0 0 0 4 dfxbp_1
rlabel metal1 s 0 -48 1748 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1748 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1748 544
string GDS_END 2578756
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2564794
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 43.700 0.000 
<< end >>
