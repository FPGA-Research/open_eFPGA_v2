magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 1 21 459 203
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 177
rect 166 47 196 177
rect 267 47 297 177
rect 351 47 381 177
<< scpmoshvt >>
rect 79 297 109 497
rect 154 297 184 497
rect 277 297 307 497
rect 349 297 379 497
<< ndiff >>
rect 27 95 79 177
rect 27 61 35 95
rect 69 61 79 95
rect 27 47 79 61
rect 109 163 166 177
rect 109 129 119 163
rect 153 129 166 163
rect 109 47 166 129
rect 196 163 267 177
rect 196 129 219 163
rect 253 129 267 163
rect 196 95 267 129
rect 196 61 219 95
rect 253 61 267 95
rect 196 47 267 61
rect 297 89 351 177
rect 297 55 307 89
rect 341 55 351 89
rect 297 47 351 55
rect 381 163 433 177
rect 381 129 391 163
rect 425 129 433 163
rect 381 95 433 129
rect 381 61 391 95
rect 425 61 433 95
rect 381 47 433 61
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 297 79 451
rect 109 297 154 497
rect 184 477 277 497
rect 184 443 194 477
rect 228 443 277 477
rect 184 409 277 443
rect 184 375 194 409
rect 228 375 277 409
rect 184 297 277 375
rect 307 297 349 497
rect 379 481 433 497
rect 379 447 389 481
rect 423 447 433 481
rect 379 413 433 447
rect 379 379 389 413
rect 423 379 433 413
rect 379 345 433 379
rect 379 311 389 345
rect 423 311 433 345
rect 379 297 433 311
<< ndiffc >>
rect 35 61 69 95
rect 119 129 153 163
rect 219 129 253 163
rect 219 61 253 95
rect 307 55 341 89
rect 391 129 425 163
rect 391 61 425 95
<< pdiffc >>
rect 35 451 69 485
rect 194 443 228 477
rect 194 375 228 409
rect 389 447 423 481
rect 389 379 423 413
rect 389 311 423 345
<< poly >>
rect 79 497 109 523
rect 154 497 184 523
rect 277 497 307 523
rect 349 497 379 523
rect 79 265 109 297
rect 21 249 109 265
rect 21 215 31 249
rect 65 215 109 249
rect 21 199 109 215
rect 154 265 184 297
rect 277 265 307 297
rect 154 249 211 265
rect 154 215 167 249
rect 201 215 211 249
rect 154 199 211 215
rect 253 249 307 265
rect 253 215 263 249
rect 297 215 307 249
rect 253 199 307 215
rect 349 265 379 297
rect 349 249 415 265
rect 349 215 367 249
rect 401 215 415 249
rect 349 199 415 215
rect 79 177 109 199
rect 166 177 196 199
rect 267 177 297 199
rect 351 177 381 199
rect 79 21 109 47
rect 166 21 196 47
rect 267 21 297 47
rect 351 21 381 47
<< polycont >>
rect 31 215 65 249
rect 167 215 201 249
rect 263 215 297 249
rect 367 215 401 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 27 485 69 527
rect 27 451 35 485
rect 27 435 69 451
rect 167 477 267 493
rect 379 481 443 527
rect 167 443 194 477
rect 228 443 267 477
rect 167 409 267 443
rect 17 249 65 398
rect 17 215 31 249
rect 17 133 65 215
rect 99 375 194 409
rect 228 375 267 409
rect 99 367 267 375
rect 99 165 133 367
rect 167 283 247 333
rect 305 323 345 481
rect 281 289 345 323
rect 379 447 389 481
rect 423 447 443 481
rect 379 413 443 447
rect 379 379 389 413
rect 423 379 443 413
rect 379 345 443 379
rect 379 311 389 345
rect 423 311 443 345
rect 379 291 443 311
rect 167 249 201 283
rect 281 249 317 289
rect 244 215 263 249
rect 297 215 317 249
rect 351 249 443 255
rect 351 215 367 249
rect 401 215 443 249
rect 167 199 201 215
rect 237 165 443 173
rect 99 163 169 165
rect 99 129 119 163
rect 153 129 169 163
rect 203 163 443 165
rect 203 129 219 163
rect 253 139 391 163
rect 253 129 269 139
rect 203 95 269 129
rect 375 129 391 139
rect 425 129 443 163
rect 17 61 35 95
rect 69 61 219 95
rect 253 61 269 95
rect 17 59 269 61
rect 307 89 341 105
rect 375 95 443 129
rect 375 61 391 95
rect 425 61 443 95
rect 375 56 443 61
rect 307 17 341 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
flabel locali s 305 357 339 391 0 FreeSans 400 0 0 0 A2
port 2 nsew signal input
flabel locali s 29 153 63 187 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel locali s 213 425 247 459 0 FreeSans 400 0 0 0 Y
port 9 nsew signal output
flabel locali s 397 221 431 255 0 FreeSans 400 0 0 0 A1
port 1 nsew signal input
flabel locali s 213 289 247 323 0 FreeSans 400 0 0 0 B2
port 4 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 o22ai_1
rlabel metal1 s 0 -48 460 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 460 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 460 544
string GDS_END 1375324
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1370488
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 2.300 0.000 
<< end >>
