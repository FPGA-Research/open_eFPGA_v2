magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -38 261 590 582
<< pwell >>
rect 1 21 551 183
rect 29 -17 63 21
<< scnmos >>
rect 79 47 473 157
<< scpmoshvt >>
rect 79 323 473 497
<< ndiff >>
rect 27 112 79 157
rect 27 78 35 112
rect 69 78 79 112
rect 27 47 79 78
rect 473 112 525 157
rect 473 78 483 112
rect 517 78 525 112
rect 473 47 525 78
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 383 79 451
rect 27 349 35 383
rect 69 349 79 383
rect 27 323 79 349
rect 473 485 525 497
rect 473 451 483 485
rect 517 451 525 485
rect 473 383 525 451
rect 473 349 483 383
rect 517 349 525 383
rect 473 323 525 349
<< ndiffc >>
rect 35 78 69 112
rect 483 78 517 112
<< pdiffc >>
rect 35 451 69 485
rect 35 349 69 383
rect 483 451 517 485
rect 483 349 517 383
<< poly >>
rect 79 497 473 523
rect 79 297 473 323
rect 79 275 255 297
rect 79 241 95 275
rect 129 241 205 275
rect 239 241 255 275
rect 79 225 255 241
rect 297 239 473 255
rect 297 205 313 239
rect 347 205 423 239
rect 457 205 473 239
rect 297 183 473 205
rect 79 157 473 183
rect 79 21 473 47
<< polycont >>
rect 95 241 129 275
rect 205 241 239 275
rect 313 205 347 239
rect 423 205 457 239
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 17 485 535 527
rect 17 451 35 485
rect 69 451 483 485
rect 517 451 535 485
rect 17 383 535 451
rect 17 349 35 383
rect 69 349 483 383
rect 517 349 535 383
rect 17 309 535 349
rect 17 241 95 275
rect 129 241 205 275
rect 239 241 259 275
rect 17 171 259 241
rect 293 239 535 309
rect 293 205 313 239
rect 347 205 423 239
rect 457 205 535 239
rect 17 112 535 171
rect 17 78 35 112
rect 69 78 483 112
rect 517 78 535 112
rect 17 17 535 78
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 4 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 3 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 2 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 decap_6
rlabel metal1 s 0 -48 552 48 1 VGND
port 1 nsew ground bidirectional abutment
rlabel metal1 s 0 496 552 592 1 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 552 544
string GDS_END 3325654
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3322568
string LEFclass CORE SPACER
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 13.800 0.000 
<< end >>
