magic
tech sky130A
timestamp 1707688321
<< properties >>
string GDS_END 58599120
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 58597708
<< end >>
