magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< metal1 >>
rect 10137 2116 10143 2168
rect 10195 2156 10201 2168
rect 12498 2156 12526 2210
rect 10195 2128 12526 2156
rect 10195 2116 10201 2128
rect 15013 2048 15019 2100
rect 15071 2088 15077 2100
rect 15841 2088 15847 2100
rect 15071 2060 15847 2088
rect 15071 2048 15077 2060
rect 15841 2048 15847 2060
rect 15899 2048 15905 2100
rect 8297 1980 8303 2032
rect 8355 2020 8361 2032
rect 9033 2020 9039 2032
rect 8355 1992 9039 2020
rect 8355 1980 8361 1992
rect 9033 1980 9039 1992
rect 9091 1980 9097 2032
rect 12529 1980 12535 2032
rect 12587 2020 12593 2032
rect 15289 2020 15295 2032
rect 12587 1992 15295 2020
rect 12587 1980 12593 1992
rect 15289 1980 15295 1992
rect 15347 1980 15353 2032
rect 10689 1912 10695 1964
rect 10747 1952 10753 1964
rect 11977 1952 11983 1964
rect 10747 1924 11983 1952
rect 10747 1912 10753 1924
rect 11977 1912 11983 1924
rect 12035 1912 12041 1964
rect 13173 1912 13179 1964
rect 13231 1952 13237 1964
rect 15473 1952 15479 1964
rect 13231 1924 15479 1952
rect 13231 1912 13237 1924
rect 15473 1912 15479 1924
rect 15531 1912 15537 1964
rect 3973 1844 3979 1896
rect 4031 1884 4037 1896
rect 4433 1884 4439 1896
rect 4031 1856 4439 1884
rect 4031 1844 4037 1856
rect 4433 1844 4439 1856
rect 4491 1844 4497 1896
rect 9493 1844 9499 1896
rect 9551 1884 9557 1896
rect 9953 1884 9959 1896
rect 9551 1856 9959 1884
rect 9551 1844 9557 1856
rect 9953 1844 9959 1856
rect 10011 1844 10017 1896
rect 14369 1844 14375 1896
rect 14427 1884 14433 1896
rect 15749 1884 15755 1896
rect 14427 1856 15755 1884
rect 14427 1844 14433 1856
rect 15749 1844 15755 1856
rect 15807 1844 15813 1896
rect 1581 892 1587 944
rect 1639 932 1645 944
rect 2133 932 2139 944
rect 1639 904 2139 932
rect 1639 892 1645 904
rect 2133 892 2139 904
rect 2191 892 2197 944
rect 5169 892 5175 944
rect 5227 932 5233 944
rect 5721 932 5727 944
rect 5227 904 5727 932
rect 5227 892 5233 904
rect 5721 892 5727 904
rect 5779 892 5785 944
rect 11977 892 11983 944
rect 12035 932 12041 944
rect 13633 932 13639 944
rect 12035 904 13639 932
rect 12035 892 12041 904
rect 13633 892 13639 904
rect 13691 892 13697 944
rect 4525 824 4531 876
rect 4583 864 4589 876
rect 5353 864 5359 876
rect 4583 836 5359 864
rect 4583 824 4589 836
rect 5353 824 5359 836
rect 5411 824 5417 876
rect 11333 824 11339 876
rect 11391 864 11397 876
rect 13357 864 13363 876
rect 11391 836 13363 864
rect 11391 824 11397 836
rect 13357 824 13363 836
rect 13415 824 13421 876
<< via1 >>
rect 10143 2116 10195 2168
rect 15019 2048 15071 2100
rect 15847 2048 15899 2100
rect 8303 1980 8355 2032
rect 9039 1980 9091 2032
rect 12535 1980 12587 2032
rect 15295 1980 15347 2032
rect 10695 1912 10747 1964
rect 11983 1912 12035 1964
rect 13179 1912 13231 1964
rect 15479 1912 15531 1964
rect 3979 1844 4031 1896
rect 4439 1844 4491 1896
rect 9499 1844 9551 1896
rect 9959 1844 10011 1896
rect 14375 1844 14427 1896
rect 15755 1844 15807 1896
rect 1587 892 1639 944
rect 2139 892 2191 944
rect 5175 892 5227 944
rect 5727 892 5779 944
rect 11983 892 12035 944
rect 13639 892 13691 944
rect 4531 824 4583 876
rect 5359 824 5411 876
rect 11339 824 11391 876
rect 13363 824 13415 876
<< metal2 >>
rect 297 2128 353 2137
rect 297 2063 353 2072
rect 311 480 339 2063
rect 679 1162 707 2236
rect 1093 2114 1121 2236
rect 1093 2086 1167 2114
rect 1139 1434 1167 2086
rect 1231 1570 1259 2236
rect 2563 2114 2591 2236
rect 2563 2086 2731 2114
rect 1231 1542 1627 1570
rect 1139 1406 1535 1434
rect 679 1134 891 1162
rect 863 480 891 1134
rect 1507 480 1535 1406
rect 1599 950 1627 1542
rect 1587 944 1639 950
rect 1587 886 1639 892
rect 2139 944 2191 950
rect 2139 886 2191 892
rect 2151 480 2179 886
rect 2703 480 2731 2086
rect 3255 1162 3283 2236
rect 4451 2222 4497 2250
rect 5346 2222 5399 2250
rect 5724 2222 5767 2250
rect 6176 2222 6227 2250
rect 4451 1902 4479 2222
rect 3979 1896 4031 1902
rect 3979 1838 4031 1844
rect 4439 1896 4491 1902
rect 4439 1838 4491 1844
rect 3255 1134 3375 1162
rect 3347 480 3375 1134
rect 3991 480 4019 1838
rect 5175 944 5227 950
rect 5175 886 5227 892
rect 4531 876 4583 882
rect 4531 818 4583 824
rect 4543 480 4571 818
rect 5187 480 5215 886
rect 5371 882 5399 2222
rect 5739 950 5767 2222
rect 6199 1162 6227 2222
rect 5831 1134 6227 1162
rect 5727 944 5779 950
rect 5727 886 5779 892
rect 5359 876 5411 882
rect 5359 818 5411 824
rect 5831 480 5859 1134
rect 6383 480 6411 2236
rect 7119 1706 7147 2236
rect 7027 1678 7147 1706
rect 7027 480 7055 1678
rect 7671 480 7699 2236
rect 8853 2128 8909 2137
rect 8853 2063 8909 2072
rect 8303 2032 8355 2038
rect 8303 1974 8355 1980
rect 8315 480 8343 1974
rect 8867 480 8895 2063
rect 9051 2038 9079 2236
rect 9039 2032 9091 2038
rect 9039 1974 9091 1980
rect 9971 1902 9999 2236
rect 10143 2168 10195 2174
rect 10143 2110 10195 2116
rect 11981 2128 12037 2137
rect 9499 1896 9551 1902
rect 9499 1838 9551 1844
rect 9959 1896 10011 1902
rect 9959 1838 10011 1844
rect 9511 480 9539 1838
rect 10155 480 10183 2110
rect 11981 2063 12037 2072
rect 11995 1970 12023 2063
rect 12535 2032 12587 2038
rect 12535 1974 12587 1980
rect 10695 1964 10747 1970
rect 10695 1906 10747 1912
rect 11983 1964 12035 1970
rect 11983 1906 12035 1912
rect 10707 480 10735 1906
rect 11983 944 12035 950
rect 11983 886 12035 892
rect 11339 876 11391 882
rect 11339 818 11391 824
rect 11351 480 11379 818
rect 11995 480 12023 886
rect 12547 480 12575 1974
rect 13179 1964 13231 1970
rect 13179 1906 13231 1912
rect 13191 480 13219 1906
rect 13375 882 13403 2236
rect 13651 950 13679 2236
rect 15019 2100 15071 2106
rect 15019 2042 15071 2048
rect 13821 1992 13877 2001
rect 13821 1927 13877 1936
rect 13639 944 13691 950
rect 13639 886 13691 892
rect 13363 876 13415 882
rect 13363 818 13415 824
rect 13835 480 13863 1927
rect 14375 1896 14427 1902
rect 14375 1838 14427 1844
rect 14387 480 14415 1838
rect 15031 480 15059 2042
rect 15307 2038 15335 2236
rect 15534 2114 15562 2236
rect 15491 2086 15562 2114
rect 15295 2032 15347 2038
rect 15295 1974 15347 1980
rect 15491 1970 15519 2086
rect 15479 1964 15531 1970
rect 15479 1906 15531 1912
rect 15767 1902 15795 2236
rect 15845 2128 15901 2137
rect 15845 2063 15847 2072
rect 15899 2063 15901 2072
rect 15847 2042 15899 2048
rect 15755 1896 15807 1902
rect 15755 1838 15807 1844
rect 15951 1162 15979 2236
rect 15675 1134 15979 1162
rect 15675 480 15703 1134
rect 297 0 353 480
rect 849 0 905 480
rect 1493 0 1549 480
rect 2137 0 2193 480
rect 2689 0 2745 480
rect 3333 0 3389 480
rect 3977 0 4033 480
rect 4529 0 4585 480
rect 5173 0 5229 480
rect 5817 0 5873 480
rect 6369 0 6425 480
rect 7013 0 7069 480
rect 7657 0 7713 480
rect 8301 0 8357 480
rect 8853 0 8909 480
rect 9497 0 9553 480
rect 10141 0 10197 480
rect 10693 0 10749 480
rect 11337 0 11393 480
rect 11981 0 12037 480
rect 12533 0 12589 480
rect 13177 0 13233 480
rect 13821 0 13877 480
rect 14373 0 14429 480
rect 15017 0 15073 480
rect 15661 0 15717 480
<< via2 >>
rect 297 2072 353 2128
rect 8853 2072 8909 2128
rect 11981 2072 12037 2128
rect 13821 1936 13877 1992
rect 15845 2100 15901 2128
rect 15845 2072 15847 2100
rect 15847 2072 15899 2100
rect 15899 2072 15901 2100
<< metal3 >>
rect 62 2130 122 2236
rect 292 2130 358 2133
rect 62 2128 358 2130
rect 62 2072 297 2128
rect 353 2072 358 2128
rect 62 2070 358 2072
rect 292 2067 358 2070
rect 8848 2130 8914 2133
rect 9176 2130 9236 2236
rect 8848 2128 9236 2130
rect 8848 2072 8853 2128
rect 8909 2072 9236 2128
rect 8848 2070 9236 2072
rect 11976 2130 12042 2133
rect 12574 2130 12634 2236
rect 11976 2128 12634 2130
rect 11976 2072 11981 2128
rect 12037 2072 12634 2128
rect 11976 2070 12634 2072
rect 8848 2067 8914 2070
rect 11976 2067 12042 2070
rect 13816 1994 13882 1997
rect 15702 1994 15762 2236
rect 15851 2133 15911 2236
rect 15840 2128 15911 2133
rect 15840 2072 15845 2128
rect 15901 2072 15911 2128
rect 15840 2070 15911 2072
rect 15840 2067 15906 2070
rect 13816 1992 15762 1994
rect 13816 1936 13821 1992
rect 13877 1936 15762 1992
rect 13816 1934 15762 1936
rect 13816 1931 13882 1934
<< metal4 >>
rect 0 37350 254 42193
rect 15746 37350 16000 42193
rect 0 16200 254 21193
rect 15746 16200 16000 21193
rect 0 15010 254 15900
rect 15746 15010 16000 15900
rect 0 13840 254 14730
rect 15746 13840 16000 14730
rect 0 13474 522 13540
rect 9418 13474 16000 13540
rect 0 12818 7288 13414
rect 7752 12818 16000 13414
rect 0 12522 254 12758
rect 15746 12522 16000 12758
rect 0 11866 10429 12462
rect 10893 11866 16000 12462
rect 0 11740 522 11806
rect 9418 11740 16000 11806
rect 0 10510 254 11440
rect 15746 10510 16000 11440
rect 0 9540 254 10230
rect 15746 9540 16000 10230
rect 0 8570 254 9260
rect 15746 8570 16000 9260
rect 0 7360 254 8290
rect 15746 7360 16000 8290
rect 0 6150 254 7080
rect 15746 6150 16000 7080
rect 0 5180 193 5870
rect 15794 5180 16000 5870
rect 0 3970 254 4900
rect 15746 3970 16000 4900
rect 0 2600 254 3690
rect 15746 2600 16000 3690
<< metal5 >>
rect 2240 23105 14760 35595
rect 0 16200 254 21190
rect 15746 16200 16000 21190
rect 0 15030 254 15880
rect 15746 15030 16000 15880
rect 0 13860 254 14710
rect 15746 13860 16000 14710
rect 0 11740 254 13540
rect 15746 11740 16000 13540
rect 0 10530 254 11420
rect 15746 10530 16000 11420
rect 0 9561 254 10210
rect 15746 9561 16000 10210
rect 0 8590 254 9240
rect 15746 8590 16000 9240
rect 0 7380 254 8270
rect 15746 7380 16000 8270
rect 0 6170 254 7060
rect 15746 6170 16000 7060
rect 0 5200 193 5850
rect 15794 5200 16000 5850
rect 0 3990 254 4880
rect 15746 3990 16000 4880
rect 0 2620 254 3670
rect 15746 2620 16000 3670
use sky130_ef_io__gpiov2_pad  gpio
timestamp 1707688321
transform 1 0 0 0 1 2600
box -143 -506 16134 39593
<< labels >>
rlabel metal4 s 7752 12818 16000 13414 4 AMUXBUS_A
port 28 nsew
rlabel metal4 s 10893 11866 16000 12462 4 AMUXBUS_B
port 29 nsew
rlabel metal2 s 10141 0 10197 480 4 ANALOG_EN
port 22 nsew
rlabel metal2 s 8853 0 8909 480 4 ANALOG_POL
port 26 nsew
rlabel metal2 s 5817 0 5873 480 4 ANALOG_SEL
port 23 nsew
rlabel metal2 s 5173 0 5229 480 4 DM[2]
port 6 nsew
rlabel metal2 s 11337 0 11393 480 4 DM[1]
port 7 nsew
rlabel metal2 s 9497 0 9553 480 4 DM[0]
port 8 nsew
rlabel metal2 s 7013 0 7069 480 4 ENABLE_H
port 13 nsew
rlabel metal2 s 7657 0 7713 480 4 ENABLE_INP_H
port 15 nsew
rlabel metal2 s 2689 0 2745 480 4 ENABLE_VDDA_H
port 14 nsew
rlabel metal2 s 13821 0 13877 480 4 ENABLE_VDDIO
port 24 nsew
rlabel metal2 s 3333 0 3389 480 4 ENABLE_VSWITCH_H
port 25 nsew
rlabel metal2 s 6369 0 6425 480 4 HLD_H_N
port 9 nsew
rlabel metal2 s 4529 0 4585 480 4 HLD_OVR
port 21 nsew
rlabel metal2 s 1493 0 1549 480 4 IB_MODE_SEL
port 12 nsew
rlabel metal2 s 15017 0 15073 480 4 IN
port 10 nsew
rlabel metal2 s 297 0 353 480 4 IN_H
port 1 nsew
rlabel metal2 s 8301 0 8357 480 4 INP_DIS
port 11 nsew
rlabel metal2 s 849 0 905 480 4 OE_N
port 16 nsew
rlabel metal2 s 3977 0 4033 480 4 OUT
port 27 nsew
rlabel metal5 s 2240 23105 14760 35595 4 PAD
port 5 nsew
rlabel metal2 s 12533 0 12589 480 4 PAD_A_ESD_0_H
port 3 nsew
rlabel metal2 s 11981 0 12037 480 4 PAD_A_ESD_1_H
port 4 nsew
rlabel metal2 s 10693 0 10749 480 4 PAD_A_NOESD_H
port 2 nsew
rlabel metal2 s 13177 0 13233 480 4 SLOW
port 19 nsew
rlabel metal2 s 14373 0 14429 480 4 TIE_HI_ESD
port 17 nsew
rlabel metal2 s 15661 0 15717 480 4 TIE_LO_ESD
port 18 nsew
rlabel metal4 s 15746 3970 16000 4900 4 VCCD
port 36 nsew
rlabel metal4 s 15746 2600 16000 3690 4 VCCHIB
port 34 nsew
rlabel metal4 s 15794 5180 16000 5870 4 VDDA
port 31 nsew
rlabel metal4 s 15746 16200 16000 21193 4 VDDIO
port 35 nsew
rlabel metal4 s 15746 15010 16000 15900 4 VDDIO_Q
port 33 nsew
rlabel metal4 s 15746 9540 16000 10230 4 VSSA
port 30 nsew
rlabel metal4 s 15746 10510 16000 11440 4 VSSD
port 38 nsew
rlabel metal4 s 15746 7360 16000 8290 4 VSSIO
port 37 nsew
rlabel metal4 s 15746 13840 16000 14730 4 VSSIO_Q
port 39 nsew
rlabel metal4 s 15746 8570 16000 9260 4 VSWITCH
port 32 nsew
rlabel metal2 s 2137 0 2193 480 4 VTRIP_SEL
port 20 nsew
<< properties >>
string FIXED_BBOX 0 0 16000 42193
string GDS_END 23644
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__gpiov2_pad_wrapped.gds
string GDS_START 154
<< end >>
