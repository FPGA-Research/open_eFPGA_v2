magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< dnwell >>
rect -4856 80 15290 13020
<< nwell >>
rect -5020 12730 15370 13100
rect -5020 370 -4650 12730
rect 15000 370 15370 12730
rect -5020 0 15370 370
<< pwell >>
rect -4462 11634 14812 11856
rect -4462 666 -4240 11634
rect -4062 1109 14412 11359
rect 14590 666 14812 11634
rect -4462 444 14812 666
<< mvnmosesd >>
tri -3664 11313 -3644 11333 ne
tri -3664 1135 -3644 1155 se
rect -3644 1135 -3534 11333
tri -3534 11313 -3514 11333 nw
tri -2372 11313 -2352 11333 ne
tri -3534 1135 -3514 1155 sw
tri -2372 1135 -2352 1155 se
rect -2352 1135 -2242 11333
tri -2242 11313 -2222 11333 nw
tri -1860 11313 -1840 11333 ne
tri -2242 1135 -2222 1155 sw
tri -1860 1135 -1840 1155 se
rect -1840 1135 -1730 11333
tri -1730 11313 -1710 11333 nw
tri -568 11313 -548 11333 ne
tri -1730 1135 -1710 1155 sw
tri -568 1135 -548 1155 se
rect -548 1135 -438 11333
tri -438 11313 -418 11333 nw
tri -56 11313 -36 11333 ne
tri -438 1135 -418 1155 sw
tri -56 1135 -36 1155 se
rect -36 1135 74 11333
tri 74 11313 94 11333 nw
tri 1236 11313 1256 11333 ne
tri 74 1135 94 1155 sw
tri 1236 1135 1256 1155 se
rect 1256 1135 1366 11333
tri 1366 11313 1386 11333 nw
tri 1748 11313 1768 11333 ne
tri 1366 1135 1386 1155 sw
tri 1748 1135 1768 1155 se
rect 1768 1135 1878 11333
tri 1878 11313 1898 11333 nw
tri 3040 11313 3060 11333 ne
tri 1878 1135 1898 1155 sw
tri 3040 1135 3060 1155 se
rect 3060 1135 3170 11333
tri 3170 11313 3190 11333 nw
tri 3552 11313 3572 11333 ne
tri 3170 1135 3190 1155 sw
tri 3552 1135 3572 1155 se
rect 3572 1135 3682 11333
tri 3682 11313 3702 11333 nw
tri 4844 11313 4864 11333 ne
tri 3682 1135 3702 1155 sw
tri 4844 1135 4864 1155 se
rect 4864 1135 4974 11333
tri 4974 11313 4994 11333 nw
tri 5356 11313 5376 11333 ne
tri 4974 1135 4994 1155 sw
tri 5356 1135 5376 1155 se
rect 5376 1135 5486 11333
tri 5486 11313 5506 11333 nw
tri 6648 11313 6668 11333 ne
tri 5486 1135 5506 1155 sw
tri 6648 1135 6668 1155 se
rect 6668 1135 6778 11333
tri 6778 11313 6798 11333 nw
tri 7160 11313 7180 11333 ne
tri 6778 1135 6798 1155 sw
tri 7160 1135 7180 1155 se
rect 7180 1135 7290 11333
tri 7290 11313 7310 11333 nw
tri 8452 11313 8472 11333 ne
tri 7290 1135 7310 1155 sw
tri 8452 1135 8472 1155 se
rect 8472 1135 8582 11333
tri 8582 11313 8602 11333 nw
tri 8964 11313 8984 11333 ne
tri 8582 1135 8602 1155 sw
tri 8964 1135 8984 1155 se
rect 8984 1135 9094 11333
tri 9094 11313 9114 11333 nw
tri 10256 11313 10276 11333 ne
tri 9094 1135 9114 1155 sw
tri 10256 1135 10276 1155 se
rect 10276 1135 10386 11333
tri 10386 11313 10406 11333 nw
tri 10768 11313 10788 11333 ne
tri 10386 1135 10406 1155 sw
tri 10768 1135 10788 1155 se
rect 10788 1135 10898 11333
tri 10898 11313 10918 11333 nw
tri 12060 11313 12080 11333 ne
tri 10898 1135 10918 1155 sw
tri 12060 1135 12080 1155 se
rect 12080 1135 12190 11333
tri 12190 11313 12210 11333 nw
tri 12572 11313 12592 11333 ne
tri 12190 1135 12210 1155 sw
tri 12572 1135 12592 1155 se
rect 12592 1135 12702 11333
tri 12702 11313 12722 11333 nw
tri 13864 11313 13884 11333 ne
tri 12702 1135 12722 1155 sw
tri 13864 1135 13884 1155 se
rect 13884 1135 13994 11333
tri 13994 11313 14014 11333 nw
tri 13994 1135 14014 1155 sw
<< mvndiff >>
rect -4036 11313 -3664 11333
tri -3664 11313 -3644 11333 sw
rect -4036 11233 -3644 11313
rect -4036 3719 -3896 11233
rect -3794 3719 -3644 11233
rect -4036 3684 -3644 3719
rect -4036 3650 -3896 3684
rect -3862 3650 -3828 3684
rect -3794 3650 -3644 3684
rect -4036 3615 -3644 3650
rect -4036 3581 -3896 3615
rect -3862 3581 -3828 3615
rect -3794 3581 -3644 3615
rect -4036 3546 -3644 3581
rect -4036 3512 -3896 3546
rect -3862 3512 -3828 3546
rect -3794 3512 -3644 3546
rect -4036 3477 -3644 3512
rect -4036 3443 -3896 3477
rect -3862 3443 -3828 3477
rect -3794 3443 -3644 3477
rect -4036 3408 -3644 3443
rect -4036 3374 -3896 3408
rect -3862 3374 -3828 3408
rect -3794 3374 -3644 3408
rect -4036 3339 -3644 3374
rect -4036 3305 -3896 3339
rect -3862 3305 -3828 3339
rect -3794 3305 -3644 3339
rect -4036 3270 -3644 3305
rect -4036 3236 -3896 3270
rect -3862 3236 -3828 3270
rect -3794 3236 -3644 3270
rect -4036 3201 -3644 3236
rect -4036 3167 -3896 3201
rect -3862 3167 -3828 3201
rect -3794 3167 -3644 3201
rect -4036 3132 -3644 3167
rect -4036 3098 -3896 3132
rect -3862 3098 -3828 3132
rect -3794 3098 -3644 3132
rect -4036 3063 -3644 3098
rect -4036 3029 -3896 3063
rect -3862 3029 -3828 3063
rect -3794 3029 -3644 3063
rect -4036 2994 -3644 3029
rect -4036 2960 -3896 2994
rect -3862 2960 -3828 2994
rect -3794 2960 -3644 2994
rect -4036 2925 -3644 2960
rect -4036 2891 -3896 2925
rect -3862 2891 -3828 2925
rect -3794 2891 -3644 2925
rect -4036 2856 -3644 2891
rect -4036 2822 -3896 2856
rect -3862 2822 -3828 2856
rect -3794 2822 -3644 2856
rect -4036 2787 -3644 2822
rect -4036 2753 -3896 2787
rect -3862 2753 -3828 2787
rect -3794 2753 -3644 2787
rect -4036 2718 -3644 2753
rect -4036 2684 -3896 2718
rect -3862 2684 -3828 2718
rect -3794 2684 -3644 2718
rect -4036 2649 -3644 2684
rect -4036 2615 -3896 2649
rect -3862 2615 -3828 2649
rect -3794 2615 -3644 2649
rect -4036 2580 -3644 2615
rect -4036 2546 -3896 2580
rect -3862 2546 -3828 2580
rect -3794 2546 -3644 2580
rect -4036 2511 -3644 2546
rect -4036 2477 -3896 2511
rect -3862 2477 -3828 2511
rect -3794 2477 -3644 2511
rect -4036 2442 -3644 2477
rect -4036 2408 -3896 2442
rect -3862 2408 -3828 2442
rect -3794 2408 -3644 2442
rect -4036 2373 -3644 2408
rect -4036 2339 -3896 2373
rect -3862 2339 -3828 2373
rect -3794 2339 -3644 2373
rect -4036 2304 -3644 2339
rect -4036 2270 -3896 2304
rect -3862 2270 -3828 2304
rect -3794 2270 -3644 2304
rect -4036 2235 -3644 2270
rect -4036 2201 -3896 2235
rect -3862 2201 -3828 2235
rect -3794 2201 -3644 2235
rect -4036 2166 -3644 2201
rect -4036 2132 -3896 2166
rect -3862 2132 -3828 2166
rect -3794 2132 -3644 2166
rect -4036 2097 -3644 2132
rect -4036 2063 -3896 2097
rect -3862 2063 -3828 2097
rect -3794 2063 -3644 2097
rect -4036 2028 -3644 2063
rect -4036 1994 -3896 2028
rect -3862 1994 -3828 2028
rect -3794 1994 -3644 2028
rect -4036 1959 -3644 1994
rect -4036 1925 -3896 1959
rect -3862 1925 -3828 1959
rect -3794 1925 -3644 1959
rect -4036 1890 -3644 1925
rect -4036 1856 -3896 1890
rect -3862 1856 -3828 1890
rect -3794 1856 -3644 1890
rect -4036 1821 -3644 1856
rect -4036 1787 -3896 1821
rect -3862 1787 -3828 1821
rect -3794 1787 -3644 1821
rect -4036 1752 -3644 1787
rect -4036 1718 -3896 1752
rect -3862 1718 -3828 1752
rect -3794 1718 -3644 1752
rect -4036 1683 -3644 1718
rect -4036 1649 -3896 1683
rect -3862 1649 -3828 1683
rect -3794 1649 -3644 1683
rect -4036 1614 -3644 1649
rect -4036 1580 -3896 1614
rect -3862 1580 -3828 1614
rect -3794 1580 -3644 1614
rect -4036 1545 -3644 1580
rect -4036 1511 -3896 1545
rect -3862 1511 -3828 1545
rect -3794 1511 -3644 1545
rect -4036 1476 -3644 1511
rect -4036 1442 -3896 1476
rect -3862 1442 -3828 1476
rect -3794 1442 -3644 1476
rect -4036 1407 -3644 1442
rect -4036 1373 -3896 1407
rect -3862 1373 -3828 1407
rect -3794 1373 -3644 1407
rect -4036 1338 -3644 1373
rect -4036 1304 -3896 1338
rect -3862 1304 -3828 1338
rect -3794 1304 -3644 1338
rect -4036 1269 -3644 1304
rect -4036 1235 -3896 1269
rect -3862 1235 -3828 1269
rect -3794 1235 -3644 1269
rect -4036 1155 -3644 1235
rect -4036 1135 -3664 1155
tri -3664 1135 -3644 1155 nw
tri -3534 11313 -3514 11333 se
rect -3514 11313 -2372 11333
tri -2372 11313 -2352 11333 sw
rect -3534 11233 -2352 11313
rect -3534 3719 -2994 11233
rect -2892 3719 -2352 11233
rect -3534 3684 -2352 3719
rect -3534 3650 -2994 3684
rect -2960 3650 -2926 3684
rect -2892 3650 -2352 3684
rect -3534 3615 -2352 3650
rect -3534 3581 -2994 3615
rect -2960 3581 -2926 3615
rect -2892 3581 -2352 3615
rect -3534 3546 -2352 3581
rect -3534 3512 -2994 3546
rect -2960 3512 -2926 3546
rect -2892 3512 -2352 3546
rect -3534 3477 -2352 3512
rect -3534 3443 -2994 3477
rect -2960 3443 -2926 3477
rect -2892 3443 -2352 3477
rect -3534 3408 -2352 3443
rect -3534 3374 -2994 3408
rect -2960 3374 -2926 3408
rect -2892 3374 -2352 3408
rect -3534 3339 -2352 3374
rect -3534 3305 -2994 3339
rect -2960 3305 -2926 3339
rect -2892 3305 -2352 3339
rect -3534 3270 -2352 3305
rect -3534 3236 -2994 3270
rect -2960 3236 -2926 3270
rect -2892 3236 -2352 3270
rect -3534 3201 -2352 3236
rect -3534 3167 -2994 3201
rect -2960 3167 -2926 3201
rect -2892 3167 -2352 3201
rect -3534 3132 -2352 3167
rect -3534 3098 -2994 3132
rect -2960 3098 -2926 3132
rect -2892 3098 -2352 3132
rect -3534 3063 -2352 3098
rect -3534 3029 -2994 3063
rect -2960 3029 -2926 3063
rect -2892 3029 -2352 3063
rect -3534 2994 -2352 3029
rect -3534 2960 -2994 2994
rect -2960 2960 -2926 2994
rect -2892 2960 -2352 2994
rect -3534 2925 -2352 2960
rect -3534 2891 -2994 2925
rect -2960 2891 -2926 2925
rect -2892 2891 -2352 2925
rect -3534 2856 -2352 2891
rect -3534 2822 -2994 2856
rect -2960 2822 -2926 2856
rect -2892 2822 -2352 2856
rect -3534 2787 -2352 2822
rect -3534 2753 -2994 2787
rect -2960 2753 -2926 2787
rect -2892 2753 -2352 2787
rect -3534 2718 -2352 2753
rect -3534 2684 -2994 2718
rect -2960 2684 -2926 2718
rect -2892 2684 -2352 2718
rect -3534 2649 -2352 2684
rect -3534 2615 -2994 2649
rect -2960 2615 -2926 2649
rect -2892 2615 -2352 2649
rect -3534 2580 -2352 2615
rect -3534 2546 -2994 2580
rect -2960 2546 -2926 2580
rect -2892 2546 -2352 2580
rect -3534 2511 -2352 2546
rect -3534 2477 -2994 2511
rect -2960 2477 -2926 2511
rect -2892 2477 -2352 2511
rect -3534 2442 -2352 2477
rect -3534 2408 -2994 2442
rect -2960 2408 -2926 2442
rect -2892 2408 -2352 2442
rect -3534 2373 -2352 2408
rect -3534 2339 -2994 2373
rect -2960 2339 -2926 2373
rect -2892 2339 -2352 2373
rect -3534 2304 -2352 2339
rect -3534 2270 -2994 2304
rect -2960 2270 -2926 2304
rect -2892 2270 -2352 2304
rect -3534 2235 -2352 2270
rect -3534 2201 -2994 2235
rect -2960 2201 -2926 2235
rect -2892 2201 -2352 2235
rect -3534 2166 -2352 2201
rect -3534 2132 -2994 2166
rect -2960 2132 -2926 2166
rect -2892 2132 -2352 2166
rect -3534 2097 -2352 2132
rect -3534 2063 -2994 2097
rect -2960 2063 -2926 2097
rect -2892 2063 -2352 2097
rect -3534 2028 -2352 2063
rect -3534 1994 -2994 2028
rect -2960 1994 -2926 2028
rect -2892 1994 -2352 2028
rect -3534 1959 -2352 1994
rect -3534 1925 -2994 1959
rect -2960 1925 -2926 1959
rect -2892 1925 -2352 1959
rect -3534 1890 -2352 1925
rect -3534 1856 -2994 1890
rect -2960 1856 -2926 1890
rect -2892 1856 -2352 1890
rect -3534 1821 -2352 1856
rect -3534 1787 -2994 1821
rect -2960 1787 -2926 1821
rect -2892 1787 -2352 1821
rect -3534 1752 -2352 1787
rect -3534 1718 -2994 1752
rect -2960 1718 -2926 1752
rect -2892 1718 -2352 1752
rect -3534 1683 -2352 1718
rect -3534 1649 -2994 1683
rect -2960 1649 -2926 1683
rect -2892 1649 -2352 1683
rect -3534 1614 -2352 1649
rect -3534 1580 -2994 1614
rect -2960 1580 -2926 1614
rect -2892 1580 -2352 1614
rect -3534 1545 -2352 1580
rect -3534 1511 -2994 1545
rect -2960 1511 -2926 1545
rect -2892 1511 -2352 1545
rect -3534 1476 -2352 1511
rect -3534 1442 -2994 1476
rect -2960 1442 -2926 1476
rect -2892 1442 -2352 1476
rect -3534 1407 -2352 1442
rect -3534 1373 -2994 1407
rect -2960 1373 -2926 1407
rect -2892 1373 -2352 1407
rect -3534 1338 -2352 1373
rect -3534 1304 -2994 1338
rect -2960 1304 -2926 1338
rect -2892 1304 -2352 1338
rect -3534 1269 -2352 1304
rect -3534 1235 -2994 1269
rect -2960 1235 -2926 1269
rect -2892 1235 -2352 1269
rect -3534 1155 -2352 1235
tri -3534 1135 -3514 1155 ne
rect -3514 1135 -2372 1155
tri -2372 1135 -2352 1155 nw
tri -2242 11313 -2222 11333 se
rect -2222 11313 -1860 11333
tri -1860 11313 -1840 11333 sw
rect -2242 11233 -1840 11313
rect -2242 3719 -2092 11233
rect -1990 3719 -1840 11233
rect -2242 3684 -1840 3719
rect -2242 3650 -2092 3684
rect -2058 3650 -2024 3684
rect -1990 3650 -1840 3684
rect -2242 3615 -1840 3650
rect -2242 3581 -2092 3615
rect -2058 3581 -2024 3615
rect -1990 3581 -1840 3615
rect -2242 3546 -1840 3581
rect -2242 3512 -2092 3546
rect -2058 3512 -2024 3546
rect -1990 3512 -1840 3546
rect -2242 3477 -1840 3512
rect -2242 3443 -2092 3477
rect -2058 3443 -2024 3477
rect -1990 3443 -1840 3477
rect -2242 3408 -1840 3443
rect -2242 3374 -2092 3408
rect -2058 3374 -2024 3408
rect -1990 3374 -1840 3408
rect -2242 3339 -1840 3374
rect -2242 3305 -2092 3339
rect -2058 3305 -2024 3339
rect -1990 3305 -1840 3339
rect -2242 3270 -1840 3305
rect -2242 3236 -2092 3270
rect -2058 3236 -2024 3270
rect -1990 3236 -1840 3270
rect -2242 3201 -1840 3236
rect -2242 3167 -2092 3201
rect -2058 3167 -2024 3201
rect -1990 3167 -1840 3201
rect -2242 3132 -1840 3167
rect -2242 3098 -2092 3132
rect -2058 3098 -2024 3132
rect -1990 3098 -1840 3132
rect -2242 3063 -1840 3098
rect -2242 3029 -2092 3063
rect -2058 3029 -2024 3063
rect -1990 3029 -1840 3063
rect -2242 2994 -1840 3029
rect -2242 2960 -2092 2994
rect -2058 2960 -2024 2994
rect -1990 2960 -1840 2994
rect -2242 2925 -1840 2960
rect -2242 2891 -2092 2925
rect -2058 2891 -2024 2925
rect -1990 2891 -1840 2925
rect -2242 2856 -1840 2891
rect -2242 2822 -2092 2856
rect -2058 2822 -2024 2856
rect -1990 2822 -1840 2856
rect -2242 2787 -1840 2822
rect -2242 2753 -2092 2787
rect -2058 2753 -2024 2787
rect -1990 2753 -1840 2787
rect -2242 2718 -1840 2753
rect -2242 2684 -2092 2718
rect -2058 2684 -2024 2718
rect -1990 2684 -1840 2718
rect -2242 2649 -1840 2684
rect -2242 2615 -2092 2649
rect -2058 2615 -2024 2649
rect -1990 2615 -1840 2649
rect -2242 2580 -1840 2615
rect -2242 2546 -2092 2580
rect -2058 2546 -2024 2580
rect -1990 2546 -1840 2580
rect -2242 2511 -1840 2546
rect -2242 2477 -2092 2511
rect -2058 2477 -2024 2511
rect -1990 2477 -1840 2511
rect -2242 2442 -1840 2477
rect -2242 2408 -2092 2442
rect -2058 2408 -2024 2442
rect -1990 2408 -1840 2442
rect -2242 2373 -1840 2408
rect -2242 2339 -2092 2373
rect -2058 2339 -2024 2373
rect -1990 2339 -1840 2373
rect -2242 2304 -1840 2339
rect -2242 2270 -2092 2304
rect -2058 2270 -2024 2304
rect -1990 2270 -1840 2304
rect -2242 2235 -1840 2270
rect -2242 2201 -2092 2235
rect -2058 2201 -2024 2235
rect -1990 2201 -1840 2235
rect -2242 2166 -1840 2201
rect -2242 2132 -2092 2166
rect -2058 2132 -2024 2166
rect -1990 2132 -1840 2166
rect -2242 2097 -1840 2132
rect -2242 2063 -2092 2097
rect -2058 2063 -2024 2097
rect -1990 2063 -1840 2097
rect -2242 2028 -1840 2063
rect -2242 1994 -2092 2028
rect -2058 1994 -2024 2028
rect -1990 1994 -1840 2028
rect -2242 1959 -1840 1994
rect -2242 1925 -2092 1959
rect -2058 1925 -2024 1959
rect -1990 1925 -1840 1959
rect -2242 1890 -1840 1925
rect -2242 1856 -2092 1890
rect -2058 1856 -2024 1890
rect -1990 1856 -1840 1890
rect -2242 1821 -1840 1856
rect -2242 1787 -2092 1821
rect -2058 1787 -2024 1821
rect -1990 1787 -1840 1821
rect -2242 1752 -1840 1787
rect -2242 1718 -2092 1752
rect -2058 1718 -2024 1752
rect -1990 1718 -1840 1752
rect -2242 1683 -1840 1718
rect -2242 1649 -2092 1683
rect -2058 1649 -2024 1683
rect -1990 1649 -1840 1683
rect -2242 1614 -1840 1649
rect -2242 1580 -2092 1614
rect -2058 1580 -2024 1614
rect -1990 1580 -1840 1614
rect -2242 1545 -1840 1580
rect -2242 1511 -2092 1545
rect -2058 1511 -2024 1545
rect -1990 1511 -1840 1545
rect -2242 1476 -1840 1511
rect -2242 1442 -2092 1476
rect -2058 1442 -2024 1476
rect -1990 1442 -1840 1476
rect -2242 1407 -1840 1442
rect -2242 1373 -2092 1407
rect -2058 1373 -2024 1407
rect -1990 1373 -1840 1407
rect -2242 1338 -1840 1373
rect -2242 1304 -2092 1338
rect -2058 1304 -2024 1338
rect -1990 1304 -1840 1338
rect -2242 1269 -1840 1304
rect -2242 1235 -2092 1269
rect -2058 1235 -2024 1269
rect -1990 1235 -1840 1269
rect -2242 1155 -1840 1235
tri -2242 1135 -2222 1155 ne
rect -2222 1135 -1860 1155
tri -1860 1135 -1840 1155 nw
tri -1730 11313 -1710 11333 se
rect -1710 11313 -568 11333
tri -568 11313 -548 11333 sw
rect -1730 11233 -548 11313
rect -1730 3719 -1190 11233
rect -1088 3719 -548 11233
rect -1730 3684 -548 3719
rect -1730 3650 -1190 3684
rect -1156 3650 -1122 3684
rect -1088 3650 -548 3684
rect -1730 3615 -548 3650
rect -1730 3581 -1190 3615
rect -1156 3581 -1122 3615
rect -1088 3581 -548 3615
rect -1730 3546 -548 3581
rect -1730 3512 -1190 3546
rect -1156 3512 -1122 3546
rect -1088 3512 -548 3546
rect -1730 3477 -548 3512
rect -1730 3443 -1190 3477
rect -1156 3443 -1122 3477
rect -1088 3443 -548 3477
rect -1730 3408 -548 3443
rect -1730 3374 -1190 3408
rect -1156 3374 -1122 3408
rect -1088 3374 -548 3408
rect -1730 3339 -548 3374
rect -1730 3305 -1190 3339
rect -1156 3305 -1122 3339
rect -1088 3305 -548 3339
rect -1730 3270 -548 3305
rect -1730 3236 -1190 3270
rect -1156 3236 -1122 3270
rect -1088 3236 -548 3270
rect -1730 3201 -548 3236
rect -1730 3167 -1190 3201
rect -1156 3167 -1122 3201
rect -1088 3167 -548 3201
rect -1730 3132 -548 3167
rect -1730 3098 -1190 3132
rect -1156 3098 -1122 3132
rect -1088 3098 -548 3132
rect -1730 3063 -548 3098
rect -1730 3029 -1190 3063
rect -1156 3029 -1122 3063
rect -1088 3029 -548 3063
rect -1730 2994 -548 3029
rect -1730 2960 -1190 2994
rect -1156 2960 -1122 2994
rect -1088 2960 -548 2994
rect -1730 2925 -548 2960
rect -1730 2891 -1190 2925
rect -1156 2891 -1122 2925
rect -1088 2891 -548 2925
rect -1730 2856 -548 2891
rect -1730 2822 -1190 2856
rect -1156 2822 -1122 2856
rect -1088 2822 -548 2856
rect -1730 2787 -548 2822
rect -1730 2753 -1190 2787
rect -1156 2753 -1122 2787
rect -1088 2753 -548 2787
rect -1730 2718 -548 2753
rect -1730 2684 -1190 2718
rect -1156 2684 -1122 2718
rect -1088 2684 -548 2718
rect -1730 2649 -548 2684
rect -1730 2615 -1190 2649
rect -1156 2615 -1122 2649
rect -1088 2615 -548 2649
rect -1730 2580 -548 2615
rect -1730 2546 -1190 2580
rect -1156 2546 -1122 2580
rect -1088 2546 -548 2580
rect -1730 2511 -548 2546
rect -1730 2477 -1190 2511
rect -1156 2477 -1122 2511
rect -1088 2477 -548 2511
rect -1730 2442 -548 2477
rect -1730 2408 -1190 2442
rect -1156 2408 -1122 2442
rect -1088 2408 -548 2442
rect -1730 2373 -548 2408
rect -1730 2339 -1190 2373
rect -1156 2339 -1122 2373
rect -1088 2339 -548 2373
rect -1730 2304 -548 2339
rect -1730 2270 -1190 2304
rect -1156 2270 -1122 2304
rect -1088 2270 -548 2304
rect -1730 2235 -548 2270
rect -1730 2201 -1190 2235
rect -1156 2201 -1122 2235
rect -1088 2201 -548 2235
rect -1730 2166 -548 2201
rect -1730 2132 -1190 2166
rect -1156 2132 -1122 2166
rect -1088 2132 -548 2166
rect -1730 2097 -548 2132
rect -1730 2063 -1190 2097
rect -1156 2063 -1122 2097
rect -1088 2063 -548 2097
rect -1730 2028 -548 2063
rect -1730 1994 -1190 2028
rect -1156 1994 -1122 2028
rect -1088 1994 -548 2028
rect -1730 1959 -548 1994
rect -1730 1925 -1190 1959
rect -1156 1925 -1122 1959
rect -1088 1925 -548 1959
rect -1730 1890 -548 1925
rect -1730 1856 -1190 1890
rect -1156 1856 -1122 1890
rect -1088 1856 -548 1890
rect -1730 1821 -548 1856
rect -1730 1787 -1190 1821
rect -1156 1787 -1122 1821
rect -1088 1787 -548 1821
rect -1730 1752 -548 1787
rect -1730 1718 -1190 1752
rect -1156 1718 -1122 1752
rect -1088 1718 -548 1752
rect -1730 1683 -548 1718
rect -1730 1649 -1190 1683
rect -1156 1649 -1122 1683
rect -1088 1649 -548 1683
rect -1730 1614 -548 1649
rect -1730 1580 -1190 1614
rect -1156 1580 -1122 1614
rect -1088 1580 -548 1614
rect -1730 1545 -548 1580
rect -1730 1511 -1190 1545
rect -1156 1511 -1122 1545
rect -1088 1511 -548 1545
rect -1730 1476 -548 1511
rect -1730 1442 -1190 1476
rect -1156 1442 -1122 1476
rect -1088 1442 -548 1476
rect -1730 1407 -548 1442
rect -1730 1373 -1190 1407
rect -1156 1373 -1122 1407
rect -1088 1373 -548 1407
rect -1730 1338 -548 1373
rect -1730 1304 -1190 1338
rect -1156 1304 -1122 1338
rect -1088 1304 -548 1338
rect -1730 1269 -548 1304
rect -1730 1235 -1190 1269
rect -1156 1235 -1122 1269
rect -1088 1235 -548 1269
rect -1730 1155 -548 1235
tri -1730 1135 -1710 1155 ne
rect -1710 1135 -568 1155
tri -568 1135 -548 1155 nw
tri -438 11313 -418 11333 se
rect -418 11313 -56 11333
tri -56 11313 -36 11333 sw
rect -438 11233 -36 11313
rect -438 3719 -288 11233
rect -186 3719 -36 11233
rect -438 3684 -36 3719
rect -438 3650 -288 3684
rect -254 3650 -220 3684
rect -186 3650 -36 3684
rect -438 3615 -36 3650
rect -438 3581 -288 3615
rect -254 3581 -220 3615
rect -186 3581 -36 3615
rect -438 3546 -36 3581
rect -438 3512 -288 3546
rect -254 3512 -220 3546
rect -186 3512 -36 3546
rect -438 3477 -36 3512
rect -438 3443 -288 3477
rect -254 3443 -220 3477
rect -186 3443 -36 3477
rect -438 3408 -36 3443
rect -438 3374 -288 3408
rect -254 3374 -220 3408
rect -186 3374 -36 3408
rect -438 3339 -36 3374
rect -438 3305 -288 3339
rect -254 3305 -220 3339
rect -186 3305 -36 3339
rect -438 3270 -36 3305
rect -438 3236 -288 3270
rect -254 3236 -220 3270
rect -186 3236 -36 3270
rect -438 3201 -36 3236
rect -438 3167 -288 3201
rect -254 3167 -220 3201
rect -186 3167 -36 3201
rect -438 3132 -36 3167
rect -438 3098 -288 3132
rect -254 3098 -220 3132
rect -186 3098 -36 3132
rect -438 3063 -36 3098
rect -438 3029 -288 3063
rect -254 3029 -220 3063
rect -186 3029 -36 3063
rect -438 2994 -36 3029
rect -438 2960 -288 2994
rect -254 2960 -220 2994
rect -186 2960 -36 2994
rect -438 2925 -36 2960
rect -438 2891 -288 2925
rect -254 2891 -220 2925
rect -186 2891 -36 2925
rect -438 2856 -36 2891
rect -438 2822 -288 2856
rect -254 2822 -220 2856
rect -186 2822 -36 2856
rect -438 2787 -36 2822
rect -438 2753 -288 2787
rect -254 2753 -220 2787
rect -186 2753 -36 2787
rect -438 2718 -36 2753
rect -438 2684 -288 2718
rect -254 2684 -220 2718
rect -186 2684 -36 2718
rect -438 2649 -36 2684
rect -438 2615 -288 2649
rect -254 2615 -220 2649
rect -186 2615 -36 2649
rect -438 2580 -36 2615
rect -438 2546 -288 2580
rect -254 2546 -220 2580
rect -186 2546 -36 2580
rect -438 2511 -36 2546
rect -438 2477 -288 2511
rect -254 2477 -220 2511
rect -186 2477 -36 2511
rect -438 2442 -36 2477
rect -438 2408 -288 2442
rect -254 2408 -220 2442
rect -186 2408 -36 2442
rect -438 2373 -36 2408
rect -438 2339 -288 2373
rect -254 2339 -220 2373
rect -186 2339 -36 2373
rect -438 2304 -36 2339
rect -438 2270 -288 2304
rect -254 2270 -220 2304
rect -186 2270 -36 2304
rect -438 2235 -36 2270
rect -438 2201 -288 2235
rect -254 2201 -220 2235
rect -186 2201 -36 2235
rect -438 2166 -36 2201
rect -438 2132 -288 2166
rect -254 2132 -220 2166
rect -186 2132 -36 2166
rect -438 2097 -36 2132
rect -438 2063 -288 2097
rect -254 2063 -220 2097
rect -186 2063 -36 2097
rect -438 2028 -36 2063
rect -438 1994 -288 2028
rect -254 1994 -220 2028
rect -186 1994 -36 2028
rect -438 1959 -36 1994
rect -438 1925 -288 1959
rect -254 1925 -220 1959
rect -186 1925 -36 1959
rect -438 1890 -36 1925
rect -438 1856 -288 1890
rect -254 1856 -220 1890
rect -186 1856 -36 1890
rect -438 1821 -36 1856
rect -438 1787 -288 1821
rect -254 1787 -220 1821
rect -186 1787 -36 1821
rect -438 1752 -36 1787
rect -438 1718 -288 1752
rect -254 1718 -220 1752
rect -186 1718 -36 1752
rect -438 1683 -36 1718
rect -438 1649 -288 1683
rect -254 1649 -220 1683
rect -186 1649 -36 1683
rect -438 1614 -36 1649
rect -438 1580 -288 1614
rect -254 1580 -220 1614
rect -186 1580 -36 1614
rect -438 1545 -36 1580
rect -438 1511 -288 1545
rect -254 1511 -220 1545
rect -186 1511 -36 1545
rect -438 1476 -36 1511
rect -438 1442 -288 1476
rect -254 1442 -220 1476
rect -186 1442 -36 1476
rect -438 1407 -36 1442
rect -438 1373 -288 1407
rect -254 1373 -220 1407
rect -186 1373 -36 1407
rect -438 1338 -36 1373
rect -438 1304 -288 1338
rect -254 1304 -220 1338
rect -186 1304 -36 1338
rect -438 1269 -36 1304
rect -438 1235 -288 1269
rect -254 1235 -220 1269
rect -186 1235 -36 1269
rect -438 1155 -36 1235
tri -438 1135 -418 1155 ne
rect -418 1135 -56 1155
tri -56 1135 -36 1155 nw
tri 74 11313 94 11333 se
rect 94 11313 1236 11333
tri 1236 11313 1256 11333 sw
rect 74 11233 1256 11313
rect 74 3719 614 11233
rect 716 3719 1256 11233
rect 74 3684 1256 3719
rect 74 3650 614 3684
rect 648 3650 682 3684
rect 716 3650 1256 3684
rect 74 3615 1256 3650
rect 74 3581 614 3615
rect 648 3581 682 3615
rect 716 3581 1256 3615
rect 74 3546 1256 3581
rect 74 3512 614 3546
rect 648 3512 682 3546
rect 716 3512 1256 3546
rect 74 3477 1256 3512
rect 74 3443 614 3477
rect 648 3443 682 3477
rect 716 3443 1256 3477
rect 74 3408 1256 3443
rect 74 3374 614 3408
rect 648 3374 682 3408
rect 716 3374 1256 3408
rect 74 3339 1256 3374
rect 74 3305 614 3339
rect 648 3305 682 3339
rect 716 3305 1256 3339
rect 74 3270 1256 3305
rect 74 3236 614 3270
rect 648 3236 682 3270
rect 716 3236 1256 3270
rect 74 3201 1256 3236
rect 74 3167 614 3201
rect 648 3167 682 3201
rect 716 3167 1256 3201
rect 74 3132 1256 3167
rect 74 3098 614 3132
rect 648 3098 682 3132
rect 716 3098 1256 3132
rect 74 3063 1256 3098
rect 74 3029 614 3063
rect 648 3029 682 3063
rect 716 3029 1256 3063
rect 74 2994 1256 3029
rect 74 2960 614 2994
rect 648 2960 682 2994
rect 716 2960 1256 2994
rect 74 2925 1256 2960
rect 74 2891 614 2925
rect 648 2891 682 2925
rect 716 2891 1256 2925
rect 74 2856 1256 2891
rect 74 2822 614 2856
rect 648 2822 682 2856
rect 716 2822 1256 2856
rect 74 2787 1256 2822
rect 74 2753 614 2787
rect 648 2753 682 2787
rect 716 2753 1256 2787
rect 74 2718 1256 2753
rect 74 2684 614 2718
rect 648 2684 682 2718
rect 716 2684 1256 2718
rect 74 2649 1256 2684
rect 74 2615 614 2649
rect 648 2615 682 2649
rect 716 2615 1256 2649
rect 74 2580 1256 2615
rect 74 2546 614 2580
rect 648 2546 682 2580
rect 716 2546 1256 2580
rect 74 2511 1256 2546
rect 74 2477 614 2511
rect 648 2477 682 2511
rect 716 2477 1256 2511
rect 74 2442 1256 2477
rect 74 2408 614 2442
rect 648 2408 682 2442
rect 716 2408 1256 2442
rect 74 2373 1256 2408
rect 74 2339 614 2373
rect 648 2339 682 2373
rect 716 2339 1256 2373
rect 74 2304 1256 2339
rect 74 2270 614 2304
rect 648 2270 682 2304
rect 716 2270 1256 2304
rect 74 2235 1256 2270
rect 74 2201 614 2235
rect 648 2201 682 2235
rect 716 2201 1256 2235
rect 74 2166 1256 2201
rect 74 2132 614 2166
rect 648 2132 682 2166
rect 716 2132 1256 2166
rect 74 2097 1256 2132
rect 74 2063 614 2097
rect 648 2063 682 2097
rect 716 2063 1256 2097
rect 74 2028 1256 2063
rect 74 1994 614 2028
rect 648 1994 682 2028
rect 716 1994 1256 2028
rect 74 1959 1256 1994
rect 74 1925 614 1959
rect 648 1925 682 1959
rect 716 1925 1256 1959
rect 74 1890 1256 1925
rect 74 1856 614 1890
rect 648 1856 682 1890
rect 716 1856 1256 1890
rect 74 1821 1256 1856
rect 74 1787 614 1821
rect 648 1787 682 1821
rect 716 1787 1256 1821
rect 74 1752 1256 1787
rect 74 1718 614 1752
rect 648 1718 682 1752
rect 716 1718 1256 1752
rect 74 1683 1256 1718
rect 74 1649 614 1683
rect 648 1649 682 1683
rect 716 1649 1256 1683
rect 74 1614 1256 1649
rect 74 1580 614 1614
rect 648 1580 682 1614
rect 716 1580 1256 1614
rect 74 1545 1256 1580
rect 74 1511 614 1545
rect 648 1511 682 1545
rect 716 1511 1256 1545
rect 74 1476 1256 1511
rect 74 1442 614 1476
rect 648 1442 682 1476
rect 716 1442 1256 1476
rect 74 1407 1256 1442
rect 74 1373 614 1407
rect 648 1373 682 1407
rect 716 1373 1256 1407
rect 74 1338 1256 1373
rect 74 1304 614 1338
rect 648 1304 682 1338
rect 716 1304 1256 1338
rect 74 1269 1256 1304
rect 74 1235 614 1269
rect 648 1235 682 1269
rect 716 1235 1256 1269
rect 74 1155 1256 1235
tri 74 1135 94 1155 ne
rect 94 1135 1236 1155
tri 1236 1135 1256 1155 nw
tri 1366 11313 1386 11333 se
rect 1386 11313 1748 11333
tri 1748 11313 1768 11333 sw
rect 1366 11233 1768 11313
rect 1366 3719 1516 11233
rect 1618 3719 1768 11233
rect 1366 3684 1768 3719
rect 1366 3650 1516 3684
rect 1550 3650 1584 3684
rect 1618 3650 1768 3684
rect 1366 3615 1768 3650
rect 1366 3581 1516 3615
rect 1550 3581 1584 3615
rect 1618 3581 1768 3615
rect 1366 3546 1768 3581
rect 1366 3512 1516 3546
rect 1550 3512 1584 3546
rect 1618 3512 1768 3546
rect 1366 3477 1768 3512
rect 1366 3443 1516 3477
rect 1550 3443 1584 3477
rect 1618 3443 1768 3477
rect 1366 3408 1768 3443
rect 1366 3374 1516 3408
rect 1550 3374 1584 3408
rect 1618 3374 1768 3408
rect 1366 3339 1768 3374
rect 1366 3305 1516 3339
rect 1550 3305 1584 3339
rect 1618 3305 1768 3339
rect 1366 3270 1768 3305
rect 1366 3236 1516 3270
rect 1550 3236 1584 3270
rect 1618 3236 1768 3270
rect 1366 3201 1768 3236
rect 1366 3167 1516 3201
rect 1550 3167 1584 3201
rect 1618 3167 1768 3201
rect 1366 3132 1768 3167
rect 1366 3098 1516 3132
rect 1550 3098 1584 3132
rect 1618 3098 1768 3132
rect 1366 3063 1768 3098
rect 1366 3029 1516 3063
rect 1550 3029 1584 3063
rect 1618 3029 1768 3063
rect 1366 2994 1768 3029
rect 1366 2960 1516 2994
rect 1550 2960 1584 2994
rect 1618 2960 1768 2994
rect 1366 2925 1768 2960
rect 1366 2891 1516 2925
rect 1550 2891 1584 2925
rect 1618 2891 1768 2925
rect 1366 2856 1768 2891
rect 1366 2822 1516 2856
rect 1550 2822 1584 2856
rect 1618 2822 1768 2856
rect 1366 2787 1768 2822
rect 1366 2753 1516 2787
rect 1550 2753 1584 2787
rect 1618 2753 1768 2787
rect 1366 2718 1768 2753
rect 1366 2684 1516 2718
rect 1550 2684 1584 2718
rect 1618 2684 1768 2718
rect 1366 2649 1768 2684
rect 1366 2615 1516 2649
rect 1550 2615 1584 2649
rect 1618 2615 1768 2649
rect 1366 2580 1768 2615
rect 1366 2546 1516 2580
rect 1550 2546 1584 2580
rect 1618 2546 1768 2580
rect 1366 2511 1768 2546
rect 1366 2477 1516 2511
rect 1550 2477 1584 2511
rect 1618 2477 1768 2511
rect 1366 2442 1768 2477
rect 1366 2408 1516 2442
rect 1550 2408 1584 2442
rect 1618 2408 1768 2442
rect 1366 2373 1768 2408
rect 1366 2339 1516 2373
rect 1550 2339 1584 2373
rect 1618 2339 1768 2373
rect 1366 2304 1768 2339
rect 1366 2270 1516 2304
rect 1550 2270 1584 2304
rect 1618 2270 1768 2304
rect 1366 2235 1768 2270
rect 1366 2201 1516 2235
rect 1550 2201 1584 2235
rect 1618 2201 1768 2235
rect 1366 2166 1768 2201
rect 1366 2132 1516 2166
rect 1550 2132 1584 2166
rect 1618 2132 1768 2166
rect 1366 2097 1768 2132
rect 1366 2063 1516 2097
rect 1550 2063 1584 2097
rect 1618 2063 1768 2097
rect 1366 2028 1768 2063
rect 1366 1994 1516 2028
rect 1550 1994 1584 2028
rect 1618 1994 1768 2028
rect 1366 1959 1768 1994
rect 1366 1925 1516 1959
rect 1550 1925 1584 1959
rect 1618 1925 1768 1959
rect 1366 1890 1768 1925
rect 1366 1856 1516 1890
rect 1550 1856 1584 1890
rect 1618 1856 1768 1890
rect 1366 1821 1768 1856
rect 1366 1787 1516 1821
rect 1550 1787 1584 1821
rect 1618 1787 1768 1821
rect 1366 1752 1768 1787
rect 1366 1718 1516 1752
rect 1550 1718 1584 1752
rect 1618 1718 1768 1752
rect 1366 1683 1768 1718
rect 1366 1649 1516 1683
rect 1550 1649 1584 1683
rect 1618 1649 1768 1683
rect 1366 1614 1768 1649
rect 1366 1580 1516 1614
rect 1550 1580 1584 1614
rect 1618 1580 1768 1614
rect 1366 1545 1768 1580
rect 1366 1511 1516 1545
rect 1550 1511 1584 1545
rect 1618 1511 1768 1545
rect 1366 1476 1768 1511
rect 1366 1442 1516 1476
rect 1550 1442 1584 1476
rect 1618 1442 1768 1476
rect 1366 1407 1768 1442
rect 1366 1373 1516 1407
rect 1550 1373 1584 1407
rect 1618 1373 1768 1407
rect 1366 1338 1768 1373
rect 1366 1304 1516 1338
rect 1550 1304 1584 1338
rect 1618 1304 1768 1338
rect 1366 1269 1768 1304
rect 1366 1235 1516 1269
rect 1550 1235 1584 1269
rect 1618 1235 1768 1269
rect 1366 1155 1768 1235
tri 1366 1135 1386 1155 ne
rect 1386 1135 1748 1155
tri 1748 1135 1768 1155 nw
tri 1878 11313 1898 11333 se
rect 1898 11313 3040 11333
tri 3040 11313 3060 11333 sw
rect 1878 11233 3060 11313
rect 1878 3719 2418 11233
rect 2520 3719 3060 11233
rect 1878 3684 3060 3719
rect 1878 3650 2418 3684
rect 2452 3650 2486 3684
rect 2520 3650 3060 3684
rect 1878 3615 3060 3650
rect 1878 3581 2418 3615
rect 2452 3581 2486 3615
rect 2520 3581 3060 3615
rect 1878 3546 3060 3581
rect 1878 3512 2418 3546
rect 2452 3512 2486 3546
rect 2520 3512 3060 3546
rect 1878 3477 3060 3512
rect 1878 3443 2418 3477
rect 2452 3443 2486 3477
rect 2520 3443 3060 3477
rect 1878 3408 3060 3443
rect 1878 3374 2418 3408
rect 2452 3374 2486 3408
rect 2520 3374 3060 3408
rect 1878 3339 3060 3374
rect 1878 3305 2418 3339
rect 2452 3305 2486 3339
rect 2520 3305 3060 3339
rect 1878 3270 3060 3305
rect 1878 3236 2418 3270
rect 2452 3236 2486 3270
rect 2520 3236 3060 3270
rect 1878 3201 3060 3236
rect 1878 3167 2418 3201
rect 2452 3167 2486 3201
rect 2520 3167 3060 3201
rect 1878 3132 3060 3167
rect 1878 3098 2418 3132
rect 2452 3098 2486 3132
rect 2520 3098 3060 3132
rect 1878 3063 3060 3098
rect 1878 3029 2418 3063
rect 2452 3029 2486 3063
rect 2520 3029 3060 3063
rect 1878 2994 3060 3029
rect 1878 2960 2418 2994
rect 2452 2960 2486 2994
rect 2520 2960 3060 2994
rect 1878 2925 3060 2960
rect 1878 2891 2418 2925
rect 2452 2891 2486 2925
rect 2520 2891 3060 2925
rect 1878 2856 3060 2891
rect 1878 2822 2418 2856
rect 2452 2822 2486 2856
rect 2520 2822 3060 2856
rect 1878 2787 3060 2822
rect 1878 2753 2418 2787
rect 2452 2753 2486 2787
rect 2520 2753 3060 2787
rect 1878 2718 3060 2753
rect 1878 2684 2418 2718
rect 2452 2684 2486 2718
rect 2520 2684 3060 2718
rect 1878 2649 3060 2684
rect 1878 2615 2418 2649
rect 2452 2615 2486 2649
rect 2520 2615 3060 2649
rect 1878 2580 3060 2615
rect 1878 2546 2418 2580
rect 2452 2546 2486 2580
rect 2520 2546 3060 2580
rect 1878 2511 3060 2546
rect 1878 2477 2418 2511
rect 2452 2477 2486 2511
rect 2520 2477 3060 2511
rect 1878 2442 3060 2477
rect 1878 2408 2418 2442
rect 2452 2408 2486 2442
rect 2520 2408 3060 2442
rect 1878 2373 3060 2408
rect 1878 2339 2418 2373
rect 2452 2339 2486 2373
rect 2520 2339 3060 2373
rect 1878 2304 3060 2339
rect 1878 2270 2418 2304
rect 2452 2270 2486 2304
rect 2520 2270 3060 2304
rect 1878 2235 3060 2270
rect 1878 2201 2418 2235
rect 2452 2201 2486 2235
rect 2520 2201 3060 2235
rect 1878 2166 3060 2201
rect 1878 2132 2418 2166
rect 2452 2132 2486 2166
rect 2520 2132 3060 2166
rect 1878 2097 3060 2132
rect 1878 2063 2418 2097
rect 2452 2063 2486 2097
rect 2520 2063 3060 2097
rect 1878 2028 3060 2063
rect 1878 1994 2418 2028
rect 2452 1994 2486 2028
rect 2520 1994 3060 2028
rect 1878 1959 3060 1994
rect 1878 1925 2418 1959
rect 2452 1925 2486 1959
rect 2520 1925 3060 1959
rect 1878 1890 3060 1925
rect 1878 1856 2418 1890
rect 2452 1856 2486 1890
rect 2520 1856 3060 1890
rect 1878 1821 3060 1856
rect 1878 1787 2418 1821
rect 2452 1787 2486 1821
rect 2520 1787 3060 1821
rect 1878 1752 3060 1787
rect 1878 1718 2418 1752
rect 2452 1718 2486 1752
rect 2520 1718 3060 1752
rect 1878 1683 3060 1718
rect 1878 1649 2418 1683
rect 2452 1649 2486 1683
rect 2520 1649 3060 1683
rect 1878 1614 3060 1649
rect 1878 1580 2418 1614
rect 2452 1580 2486 1614
rect 2520 1580 3060 1614
rect 1878 1545 3060 1580
rect 1878 1511 2418 1545
rect 2452 1511 2486 1545
rect 2520 1511 3060 1545
rect 1878 1476 3060 1511
rect 1878 1442 2418 1476
rect 2452 1442 2486 1476
rect 2520 1442 3060 1476
rect 1878 1407 3060 1442
rect 1878 1373 2418 1407
rect 2452 1373 2486 1407
rect 2520 1373 3060 1407
rect 1878 1338 3060 1373
rect 1878 1304 2418 1338
rect 2452 1304 2486 1338
rect 2520 1304 3060 1338
rect 1878 1269 3060 1304
rect 1878 1235 2418 1269
rect 2452 1235 2486 1269
rect 2520 1235 3060 1269
rect 1878 1155 3060 1235
tri 1878 1135 1898 1155 ne
rect 1898 1135 3040 1155
tri 3040 1135 3060 1155 nw
tri 3170 11313 3190 11333 se
rect 3190 11313 3552 11333
tri 3552 11313 3572 11333 sw
rect 3170 11233 3572 11313
rect 3170 3719 3320 11233
rect 3422 3719 3572 11233
rect 3170 3684 3572 3719
rect 3170 3650 3320 3684
rect 3354 3650 3388 3684
rect 3422 3650 3572 3684
rect 3170 3615 3572 3650
rect 3170 3581 3320 3615
rect 3354 3581 3388 3615
rect 3422 3581 3572 3615
rect 3170 3546 3572 3581
rect 3170 3512 3320 3546
rect 3354 3512 3388 3546
rect 3422 3512 3572 3546
rect 3170 3477 3572 3512
rect 3170 3443 3320 3477
rect 3354 3443 3388 3477
rect 3422 3443 3572 3477
rect 3170 3408 3572 3443
rect 3170 3374 3320 3408
rect 3354 3374 3388 3408
rect 3422 3374 3572 3408
rect 3170 3339 3572 3374
rect 3170 3305 3320 3339
rect 3354 3305 3388 3339
rect 3422 3305 3572 3339
rect 3170 3270 3572 3305
rect 3170 3236 3320 3270
rect 3354 3236 3388 3270
rect 3422 3236 3572 3270
rect 3170 3201 3572 3236
rect 3170 3167 3320 3201
rect 3354 3167 3388 3201
rect 3422 3167 3572 3201
rect 3170 3132 3572 3167
rect 3170 3098 3320 3132
rect 3354 3098 3388 3132
rect 3422 3098 3572 3132
rect 3170 3063 3572 3098
rect 3170 3029 3320 3063
rect 3354 3029 3388 3063
rect 3422 3029 3572 3063
rect 3170 2994 3572 3029
rect 3170 2960 3320 2994
rect 3354 2960 3388 2994
rect 3422 2960 3572 2994
rect 3170 2925 3572 2960
rect 3170 2891 3320 2925
rect 3354 2891 3388 2925
rect 3422 2891 3572 2925
rect 3170 2856 3572 2891
rect 3170 2822 3320 2856
rect 3354 2822 3388 2856
rect 3422 2822 3572 2856
rect 3170 2787 3572 2822
rect 3170 2753 3320 2787
rect 3354 2753 3388 2787
rect 3422 2753 3572 2787
rect 3170 2718 3572 2753
rect 3170 2684 3320 2718
rect 3354 2684 3388 2718
rect 3422 2684 3572 2718
rect 3170 2649 3572 2684
rect 3170 2615 3320 2649
rect 3354 2615 3388 2649
rect 3422 2615 3572 2649
rect 3170 2580 3572 2615
rect 3170 2546 3320 2580
rect 3354 2546 3388 2580
rect 3422 2546 3572 2580
rect 3170 2511 3572 2546
rect 3170 2477 3320 2511
rect 3354 2477 3388 2511
rect 3422 2477 3572 2511
rect 3170 2442 3572 2477
rect 3170 2408 3320 2442
rect 3354 2408 3388 2442
rect 3422 2408 3572 2442
rect 3170 2373 3572 2408
rect 3170 2339 3320 2373
rect 3354 2339 3388 2373
rect 3422 2339 3572 2373
rect 3170 2304 3572 2339
rect 3170 2270 3320 2304
rect 3354 2270 3388 2304
rect 3422 2270 3572 2304
rect 3170 2235 3572 2270
rect 3170 2201 3320 2235
rect 3354 2201 3388 2235
rect 3422 2201 3572 2235
rect 3170 2166 3572 2201
rect 3170 2132 3320 2166
rect 3354 2132 3388 2166
rect 3422 2132 3572 2166
rect 3170 2097 3572 2132
rect 3170 2063 3320 2097
rect 3354 2063 3388 2097
rect 3422 2063 3572 2097
rect 3170 2028 3572 2063
rect 3170 1994 3320 2028
rect 3354 1994 3388 2028
rect 3422 1994 3572 2028
rect 3170 1959 3572 1994
rect 3170 1925 3320 1959
rect 3354 1925 3388 1959
rect 3422 1925 3572 1959
rect 3170 1890 3572 1925
rect 3170 1856 3320 1890
rect 3354 1856 3388 1890
rect 3422 1856 3572 1890
rect 3170 1821 3572 1856
rect 3170 1787 3320 1821
rect 3354 1787 3388 1821
rect 3422 1787 3572 1821
rect 3170 1752 3572 1787
rect 3170 1718 3320 1752
rect 3354 1718 3388 1752
rect 3422 1718 3572 1752
rect 3170 1683 3572 1718
rect 3170 1649 3320 1683
rect 3354 1649 3388 1683
rect 3422 1649 3572 1683
rect 3170 1614 3572 1649
rect 3170 1580 3320 1614
rect 3354 1580 3388 1614
rect 3422 1580 3572 1614
rect 3170 1545 3572 1580
rect 3170 1511 3320 1545
rect 3354 1511 3388 1545
rect 3422 1511 3572 1545
rect 3170 1476 3572 1511
rect 3170 1442 3320 1476
rect 3354 1442 3388 1476
rect 3422 1442 3572 1476
rect 3170 1407 3572 1442
rect 3170 1373 3320 1407
rect 3354 1373 3388 1407
rect 3422 1373 3572 1407
rect 3170 1338 3572 1373
rect 3170 1304 3320 1338
rect 3354 1304 3388 1338
rect 3422 1304 3572 1338
rect 3170 1269 3572 1304
rect 3170 1235 3320 1269
rect 3354 1235 3388 1269
rect 3422 1235 3572 1269
rect 3170 1155 3572 1235
tri 3170 1135 3190 1155 ne
rect 3190 1135 3552 1155
tri 3552 1135 3572 1155 nw
tri 3682 11313 3702 11333 se
rect 3702 11313 4844 11333
tri 4844 11313 4864 11333 sw
rect 3682 11233 4864 11313
rect 3682 3719 4222 11233
rect 4324 3719 4864 11233
rect 3682 3684 4864 3719
rect 3682 3650 4222 3684
rect 4256 3650 4290 3684
rect 4324 3650 4864 3684
rect 3682 3615 4864 3650
rect 3682 3581 4222 3615
rect 4256 3581 4290 3615
rect 4324 3581 4864 3615
rect 3682 3546 4864 3581
rect 3682 3512 4222 3546
rect 4256 3512 4290 3546
rect 4324 3512 4864 3546
rect 3682 3477 4864 3512
rect 3682 3443 4222 3477
rect 4256 3443 4290 3477
rect 4324 3443 4864 3477
rect 3682 3408 4864 3443
rect 3682 3374 4222 3408
rect 4256 3374 4290 3408
rect 4324 3374 4864 3408
rect 3682 3339 4864 3374
rect 3682 3305 4222 3339
rect 4256 3305 4290 3339
rect 4324 3305 4864 3339
rect 3682 3270 4864 3305
rect 3682 3236 4222 3270
rect 4256 3236 4290 3270
rect 4324 3236 4864 3270
rect 3682 3201 4864 3236
rect 3682 3167 4222 3201
rect 4256 3167 4290 3201
rect 4324 3167 4864 3201
rect 3682 3132 4864 3167
rect 3682 3098 4222 3132
rect 4256 3098 4290 3132
rect 4324 3098 4864 3132
rect 3682 3063 4864 3098
rect 3682 3029 4222 3063
rect 4256 3029 4290 3063
rect 4324 3029 4864 3063
rect 3682 2994 4864 3029
rect 3682 2960 4222 2994
rect 4256 2960 4290 2994
rect 4324 2960 4864 2994
rect 3682 2925 4864 2960
rect 3682 2891 4222 2925
rect 4256 2891 4290 2925
rect 4324 2891 4864 2925
rect 3682 2856 4864 2891
rect 3682 2822 4222 2856
rect 4256 2822 4290 2856
rect 4324 2822 4864 2856
rect 3682 2787 4864 2822
rect 3682 2753 4222 2787
rect 4256 2753 4290 2787
rect 4324 2753 4864 2787
rect 3682 2718 4864 2753
rect 3682 2684 4222 2718
rect 4256 2684 4290 2718
rect 4324 2684 4864 2718
rect 3682 2649 4864 2684
rect 3682 2615 4222 2649
rect 4256 2615 4290 2649
rect 4324 2615 4864 2649
rect 3682 2580 4864 2615
rect 3682 2546 4222 2580
rect 4256 2546 4290 2580
rect 4324 2546 4864 2580
rect 3682 2511 4864 2546
rect 3682 2477 4222 2511
rect 4256 2477 4290 2511
rect 4324 2477 4864 2511
rect 3682 2442 4864 2477
rect 3682 2408 4222 2442
rect 4256 2408 4290 2442
rect 4324 2408 4864 2442
rect 3682 2373 4864 2408
rect 3682 2339 4222 2373
rect 4256 2339 4290 2373
rect 4324 2339 4864 2373
rect 3682 2304 4864 2339
rect 3682 2270 4222 2304
rect 4256 2270 4290 2304
rect 4324 2270 4864 2304
rect 3682 2235 4864 2270
rect 3682 2201 4222 2235
rect 4256 2201 4290 2235
rect 4324 2201 4864 2235
rect 3682 2166 4864 2201
rect 3682 2132 4222 2166
rect 4256 2132 4290 2166
rect 4324 2132 4864 2166
rect 3682 2097 4864 2132
rect 3682 2063 4222 2097
rect 4256 2063 4290 2097
rect 4324 2063 4864 2097
rect 3682 2028 4864 2063
rect 3682 1994 4222 2028
rect 4256 1994 4290 2028
rect 4324 1994 4864 2028
rect 3682 1959 4864 1994
rect 3682 1925 4222 1959
rect 4256 1925 4290 1959
rect 4324 1925 4864 1959
rect 3682 1890 4864 1925
rect 3682 1856 4222 1890
rect 4256 1856 4290 1890
rect 4324 1856 4864 1890
rect 3682 1821 4864 1856
rect 3682 1787 4222 1821
rect 4256 1787 4290 1821
rect 4324 1787 4864 1821
rect 3682 1752 4864 1787
rect 3682 1718 4222 1752
rect 4256 1718 4290 1752
rect 4324 1718 4864 1752
rect 3682 1683 4864 1718
rect 3682 1649 4222 1683
rect 4256 1649 4290 1683
rect 4324 1649 4864 1683
rect 3682 1614 4864 1649
rect 3682 1580 4222 1614
rect 4256 1580 4290 1614
rect 4324 1580 4864 1614
rect 3682 1545 4864 1580
rect 3682 1511 4222 1545
rect 4256 1511 4290 1545
rect 4324 1511 4864 1545
rect 3682 1476 4864 1511
rect 3682 1442 4222 1476
rect 4256 1442 4290 1476
rect 4324 1442 4864 1476
rect 3682 1407 4864 1442
rect 3682 1373 4222 1407
rect 4256 1373 4290 1407
rect 4324 1373 4864 1407
rect 3682 1338 4864 1373
rect 3682 1304 4222 1338
rect 4256 1304 4290 1338
rect 4324 1304 4864 1338
rect 3682 1269 4864 1304
rect 3682 1235 4222 1269
rect 4256 1235 4290 1269
rect 4324 1235 4864 1269
rect 3682 1155 4864 1235
tri 3682 1135 3702 1155 ne
rect 3702 1135 4844 1155
tri 4844 1135 4864 1155 nw
tri 4974 11313 4994 11333 se
rect 4994 11313 5356 11333
tri 5356 11313 5376 11333 sw
rect 4974 11233 5376 11313
rect 4974 3719 5124 11233
rect 5226 3719 5376 11233
rect 4974 3684 5376 3719
rect 4974 3650 5124 3684
rect 5158 3650 5192 3684
rect 5226 3650 5376 3684
rect 4974 3615 5376 3650
rect 4974 3581 5124 3615
rect 5158 3581 5192 3615
rect 5226 3581 5376 3615
rect 4974 3546 5376 3581
rect 4974 3512 5124 3546
rect 5158 3512 5192 3546
rect 5226 3512 5376 3546
rect 4974 3477 5376 3512
rect 4974 3443 5124 3477
rect 5158 3443 5192 3477
rect 5226 3443 5376 3477
rect 4974 3408 5376 3443
rect 4974 3374 5124 3408
rect 5158 3374 5192 3408
rect 5226 3374 5376 3408
rect 4974 3339 5376 3374
rect 4974 3305 5124 3339
rect 5158 3305 5192 3339
rect 5226 3305 5376 3339
rect 4974 3270 5376 3305
rect 4974 3236 5124 3270
rect 5158 3236 5192 3270
rect 5226 3236 5376 3270
rect 4974 3201 5376 3236
rect 4974 3167 5124 3201
rect 5158 3167 5192 3201
rect 5226 3167 5376 3201
rect 4974 3132 5376 3167
rect 4974 3098 5124 3132
rect 5158 3098 5192 3132
rect 5226 3098 5376 3132
rect 4974 3063 5376 3098
rect 4974 3029 5124 3063
rect 5158 3029 5192 3063
rect 5226 3029 5376 3063
rect 4974 2994 5376 3029
rect 4974 2960 5124 2994
rect 5158 2960 5192 2994
rect 5226 2960 5376 2994
rect 4974 2925 5376 2960
rect 4974 2891 5124 2925
rect 5158 2891 5192 2925
rect 5226 2891 5376 2925
rect 4974 2856 5376 2891
rect 4974 2822 5124 2856
rect 5158 2822 5192 2856
rect 5226 2822 5376 2856
rect 4974 2787 5376 2822
rect 4974 2753 5124 2787
rect 5158 2753 5192 2787
rect 5226 2753 5376 2787
rect 4974 2718 5376 2753
rect 4974 2684 5124 2718
rect 5158 2684 5192 2718
rect 5226 2684 5376 2718
rect 4974 2649 5376 2684
rect 4974 2615 5124 2649
rect 5158 2615 5192 2649
rect 5226 2615 5376 2649
rect 4974 2580 5376 2615
rect 4974 2546 5124 2580
rect 5158 2546 5192 2580
rect 5226 2546 5376 2580
rect 4974 2511 5376 2546
rect 4974 2477 5124 2511
rect 5158 2477 5192 2511
rect 5226 2477 5376 2511
rect 4974 2442 5376 2477
rect 4974 2408 5124 2442
rect 5158 2408 5192 2442
rect 5226 2408 5376 2442
rect 4974 2373 5376 2408
rect 4974 2339 5124 2373
rect 5158 2339 5192 2373
rect 5226 2339 5376 2373
rect 4974 2304 5376 2339
rect 4974 2270 5124 2304
rect 5158 2270 5192 2304
rect 5226 2270 5376 2304
rect 4974 2235 5376 2270
rect 4974 2201 5124 2235
rect 5158 2201 5192 2235
rect 5226 2201 5376 2235
rect 4974 2166 5376 2201
rect 4974 2132 5124 2166
rect 5158 2132 5192 2166
rect 5226 2132 5376 2166
rect 4974 2097 5376 2132
rect 4974 2063 5124 2097
rect 5158 2063 5192 2097
rect 5226 2063 5376 2097
rect 4974 2028 5376 2063
rect 4974 1994 5124 2028
rect 5158 1994 5192 2028
rect 5226 1994 5376 2028
rect 4974 1959 5376 1994
rect 4974 1925 5124 1959
rect 5158 1925 5192 1959
rect 5226 1925 5376 1959
rect 4974 1890 5376 1925
rect 4974 1856 5124 1890
rect 5158 1856 5192 1890
rect 5226 1856 5376 1890
rect 4974 1821 5376 1856
rect 4974 1787 5124 1821
rect 5158 1787 5192 1821
rect 5226 1787 5376 1821
rect 4974 1752 5376 1787
rect 4974 1718 5124 1752
rect 5158 1718 5192 1752
rect 5226 1718 5376 1752
rect 4974 1683 5376 1718
rect 4974 1649 5124 1683
rect 5158 1649 5192 1683
rect 5226 1649 5376 1683
rect 4974 1614 5376 1649
rect 4974 1580 5124 1614
rect 5158 1580 5192 1614
rect 5226 1580 5376 1614
rect 4974 1545 5376 1580
rect 4974 1511 5124 1545
rect 5158 1511 5192 1545
rect 5226 1511 5376 1545
rect 4974 1476 5376 1511
rect 4974 1442 5124 1476
rect 5158 1442 5192 1476
rect 5226 1442 5376 1476
rect 4974 1407 5376 1442
rect 4974 1373 5124 1407
rect 5158 1373 5192 1407
rect 5226 1373 5376 1407
rect 4974 1338 5376 1373
rect 4974 1304 5124 1338
rect 5158 1304 5192 1338
rect 5226 1304 5376 1338
rect 4974 1269 5376 1304
rect 4974 1235 5124 1269
rect 5158 1235 5192 1269
rect 5226 1235 5376 1269
rect 4974 1155 5376 1235
tri 4974 1135 4994 1155 ne
rect 4994 1135 5356 1155
tri 5356 1135 5376 1155 nw
tri 5486 11313 5506 11333 se
rect 5506 11313 6648 11333
tri 6648 11313 6668 11333 sw
rect 5486 11233 6668 11313
rect 5486 3719 6026 11233
rect 6128 3719 6668 11233
rect 5486 3684 6668 3719
rect 5486 3650 6026 3684
rect 6060 3650 6094 3684
rect 6128 3650 6668 3684
rect 5486 3615 6668 3650
rect 5486 3581 6026 3615
rect 6060 3581 6094 3615
rect 6128 3581 6668 3615
rect 5486 3546 6668 3581
rect 5486 3512 6026 3546
rect 6060 3512 6094 3546
rect 6128 3512 6668 3546
rect 5486 3477 6668 3512
rect 5486 3443 6026 3477
rect 6060 3443 6094 3477
rect 6128 3443 6668 3477
rect 5486 3408 6668 3443
rect 5486 3374 6026 3408
rect 6060 3374 6094 3408
rect 6128 3374 6668 3408
rect 5486 3339 6668 3374
rect 5486 3305 6026 3339
rect 6060 3305 6094 3339
rect 6128 3305 6668 3339
rect 5486 3270 6668 3305
rect 5486 3236 6026 3270
rect 6060 3236 6094 3270
rect 6128 3236 6668 3270
rect 5486 3201 6668 3236
rect 5486 3167 6026 3201
rect 6060 3167 6094 3201
rect 6128 3167 6668 3201
rect 5486 3132 6668 3167
rect 5486 3098 6026 3132
rect 6060 3098 6094 3132
rect 6128 3098 6668 3132
rect 5486 3063 6668 3098
rect 5486 3029 6026 3063
rect 6060 3029 6094 3063
rect 6128 3029 6668 3063
rect 5486 2994 6668 3029
rect 5486 2960 6026 2994
rect 6060 2960 6094 2994
rect 6128 2960 6668 2994
rect 5486 2925 6668 2960
rect 5486 2891 6026 2925
rect 6060 2891 6094 2925
rect 6128 2891 6668 2925
rect 5486 2856 6668 2891
rect 5486 2822 6026 2856
rect 6060 2822 6094 2856
rect 6128 2822 6668 2856
rect 5486 2787 6668 2822
rect 5486 2753 6026 2787
rect 6060 2753 6094 2787
rect 6128 2753 6668 2787
rect 5486 2718 6668 2753
rect 5486 2684 6026 2718
rect 6060 2684 6094 2718
rect 6128 2684 6668 2718
rect 5486 2649 6668 2684
rect 5486 2615 6026 2649
rect 6060 2615 6094 2649
rect 6128 2615 6668 2649
rect 5486 2580 6668 2615
rect 5486 2546 6026 2580
rect 6060 2546 6094 2580
rect 6128 2546 6668 2580
rect 5486 2511 6668 2546
rect 5486 2477 6026 2511
rect 6060 2477 6094 2511
rect 6128 2477 6668 2511
rect 5486 2442 6668 2477
rect 5486 2408 6026 2442
rect 6060 2408 6094 2442
rect 6128 2408 6668 2442
rect 5486 2373 6668 2408
rect 5486 2339 6026 2373
rect 6060 2339 6094 2373
rect 6128 2339 6668 2373
rect 5486 2304 6668 2339
rect 5486 2270 6026 2304
rect 6060 2270 6094 2304
rect 6128 2270 6668 2304
rect 5486 2235 6668 2270
rect 5486 2201 6026 2235
rect 6060 2201 6094 2235
rect 6128 2201 6668 2235
rect 5486 2166 6668 2201
rect 5486 2132 6026 2166
rect 6060 2132 6094 2166
rect 6128 2132 6668 2166
rect 5486 2097 6668 2132
rect 5486 2063 6026 2097
rect 6060 2063 6094 2097
rect 6128 2063 6668 2097
rect 5486 2028 6668 2063
rect 5486 1994 6026 2028
rect 6060 1994 6094 2028
rect 6128 1994 6668 2028
rect 5486 1959 6668 1994
rect 5486 1925 6026 1959
rect 6060 1925 6094 1959
rect 6128 1925 6668 1959
rect 5486 1890 6668 1925
rect 5486 1856 6026 1890
rect 6060 1856 6094 1890
rect 6128 1856 6668 1890
rect 5486 1821 6668 1856
rect 5486 1787 6026 1821
rect 6060 1787 6094 1821
rect 6128 1787 6668 1821
rect 5486 1752 6668 1787
rect 5486 1718 6026 1752
rect 6060 1718 6094 1752
rect 6128 1718 6668 1752
rect 5486 1683 6668 1718
rect 5486 1649 6026 1683
rect 6060 1649 6094 1683
rect 6128 1649 6668 1683
rect 5486 1614 6668 1649
rect 5486 1580 6026 1614
rect 6060 1580 6094 1614
rect 6128 1580 6668 1614
rect 5486 1545 6668 1580
rect 5486 1511 6026 1545
rect 6060 1511 6094 1545
rect 6128 1511 6668 1545
rect 5486 1476 6668 1511
rect 5486 1442 6026 1476
rect 6060 1442 6094 1476
rect 6128 1442 6668 1476
rect 5486 1407 6668 1442
rect 5486 1373 6026 1407
rect 6060 1373 6094 1407
rect 6128 1373 6668 1407
rect 5486 1338 6668 1373
rect 5486 1304 6026 1338
rect 6060 1304 6094 1338
rect 6128 1304 6668 1338
rect 5486 1269 6668 1304
rect 5486 1235 6026 1269
rect 6060 1235 6094 1269
rect 6128 1235 6668 1269
rect 5486 1155 6668 1235
tri 5486 1135 5506 1155 ne
rect 5506 1135 6648 1155
tri 6648 1135 6668 1155 nw
tri 6778 11313 6798 11333 se
rect 6798 11313 7160 11333
tri 7160 11313 7180 11333 sw
rect 6778 11233 7180 11313
rect 6778 3719 6928 11233
rect 7030 3719 7180 11233
rect 6778 3684 7180 3719
rect 6778 3650 6928 3684
rect 6962 3650 6996 3684
rect 7030 3650 7180 3684
rect 6778 3615 7180 3650
rect 6778 3581 6928 3615
rect 6962 3581 6996 3615
rect 7030 3581 7180 3615
rect 6778 3546 7180 3581
rect 6778 3512 6928 3546
rect 6962 3512 6996 3546
rect 7030 3512 7180 3546
rect 6778 3477 7180 3512
rect 6778 3443 6928 3477
rect 6962 3443 6996 3477
rect 7030 3443 7180 3477
rect 6778 3408 7180 3443
rect 6778 3374 6928 3408
rect 6962 3374 6996 3408
rect 7030 3374 7180 3408
rect 6778 3339 7180 3374
rect 6778 3305 6928 3339
rect 6962 3305 6996 3339
rect 7030 3305 7180 3339
rect 6778 3270 7180 3305
rect 6778 3236 6928 3270
rect 6962 3236 6996 3270
rect 7030 3236 7180 3270
rect 6778 3201 7180 3236
rect 6778 3167 6928 3201
rect 6962 3167 6996 3201
rect 7030 3167 7180 3201
rect 6778 3132 7180 3167
rect 6778 3098 6928 3132
rect 6962 3098 6996 3132
rect 7030 3098 7180 3132
rect 6778 3063 7180 3098
rect 6778 3029 6928 3063
rect 6962 3029 6996 3063
rect 7030 3029 7180 3063
rect 6778 2994 7180 3029
rect 6778 2960 6928 2994
rect 6962 2960 6996 2994
rect 7030 2960 7180 2994
rect 6778 2925 7180 2960
rect 6778 2891 6928 2925
rect 6962 2891 6996 2925
rect 7030 2891 7180 2925
rect 6778 2856 7180 2891
rect 6778 2822 6928 2856
rect 6962 2822 6996 2856
rect 7030 2822 7180 2856
rect 6778 2787 7180 2822
rect 6778 2753 6928 2787
rect 6962 2753 6996 2787
rect 7030 2753 7180 2787
rect 6778 2718 7180 2753
rect 6778 2684 6928 2718
rect 6962 2684 6996 2718
rect 7030 2684 7180 2718
rect 6778 2649 7180 2684
rect 6778 2615 6928 2649
rect 6962 2615 6996 2649
rect 7030 2615 7180 2649
rect 6778 2580 7180 2615
rect 6778 2546 6928 2580
rect 6962 2546 6996 2580
rect 7030 2546 7180 2580
rect 6778 2511 7180 2546
rect 6778 2477 6928 2511
rect 6962 2477 6996 2511
rect 7030 2477 7180 2511
rect 6778 2442 7180 2477
rect 6778 2408 6928 2442
rect 6962 2408 6996 2442
rect 7030 2408 7180 2442
rect 6778 2373 7180 2408
rect 6778 2339 6928 2373
rect 6962 2339 6996 2373
rect 7030 2339 7180 2373
rect 6778 2304 7180 2339
rect 6778 2270 6928 2304
rect 6962 2270 6996 2304
rect 7030 2270 7180 2304
rect 6778 2235 7180 2270
rect 6778 2201 6928 2235
rect 6962 2201 6996 2235
rect 7030 2201 7180 2235
rect 6778 2166 7180 2201
rect 6778 2132 6928 2166
rect 6962 2132 6996 2166
rect 7030 2132 7180 2166
rect 6778 2097 7180 2132
rect 6778 2063 6928 2097
rect 6962 2063 6996 2097
rect 7030 2063 7180 2097
rect 6778 2028 7180 2063
rect 6778 1994 6928 2028
rect 6962 1994 6996 2028
rect 7030 1994 7180 2028
rect 6778 1959 7180 1994
rect 6778 1925 6928 1959
rect 6962 1925 6996 1959
rect 7030 1925 7180 1959
rect 6778 1890 7180 1925
rect 6778 1856 6928 1890
rect 6962 1856 6996 1890
rect 7030 1856 7180 1890
rect 6778 1821 7180 1856
rect 6778 1787 6928 1821
rect 6962 1787 6996 1821
rect 7030 1787 7180 1821
rect 6778 1752 7180 1787
rect 6778 1718 6928 1752
rect 6962 1718 6996 1752
rect 7030 1718 7180 1752
rect 6778 1683 7180 1718
rect 6778 1649 6928 1683
rect 6962 1649 6996 1683
rect 7030 1649 7180 1683
rect 6778 1614 7180 1649
rect 6778 1580 6928 1614
rect 6962 1580 6996 1614
rect 7030 1580 7180 1614
rect 6778 1545 7180 1580
rect 6778 1511 6928 1545
rect 6962 1511 6996 1545
rect 7030 1511 7180 1545
rect 6778 1476 7180 1511
rect 6778 1442 6928 1476
rect 6962 1442 6996 1476
rect 7030 1442 7180 1476
rect 6778 1407 7180 1442
rect 6778 1373 6928 1407
rect 6962 1373 6996 1407
rect 7030 1373 7180 1407
rect 6778 1338 7180 1373
rect 6778 1304 6928 1338
rect 6962 1304 6996 1338
rect 7030 1304 7180 1338
rect 6778 1269 7180 1304
rect 6778 1235 6928 1269
rect 6962 1235 6996 1269
rect 7030 1235 7180 1269
rect 6778 1155 7180 1235
tri 6778 1135 6798 1155 ne
rect 6798 1135 7160 1155
tri 7160 1135 7180 1155 nw
tri 7290 11313 7310 11333 se
rect 7310 11313 8452 11333
tri 8452 11313 8472 11333 sw
rect 7290 11233 8472 11313
rect 7290 3719 7830 11233
rect 7932 3719 8472 11233
rect 7290 3684 8472 3719
rect 7290 3650 7830 3684
rect 7864 3650 7898 3684
rect 7932 3650 8472 3684
rect 7290 3615 8472 3650
rect 7290 3581 7830 3615
rect 7864 3581 7898 3615
rect 7932 3581 8472 3615
rect 7290 3546 8472 3581
rect 7290 3512 7830 3546
rect 7864 3512 7898 3546
rect 7932 3512 8472 3546
rect 7290 3477 8472 3512
rect 7290 3443 7830 3477
rect 7864 3443 7898 3477
rect 7932 3443 8472 3477
rect 7290 3408 8472 3443
rect 7290 3374 7830 3408
rect 7864 3374 7898 3408
rect 7932 3374 8472 3408
rect 7290 3339 8472 3374
rect 7290 3305 7830 3339
rect 7864 3305 7898 3339
rect 7932 3305 8472 3339
rect 7290 3270 8472 3305
rect 7290 3236 7830 3270
rect 7864 3236 7898 3270
rect 7932 3236 8472 3270
rect 7290 3201 8472 3236
rect 7290 3167 7830 3201
rect 7864 3167 7898 3201
rect 7932 3167 8472 3201
rect 7290 3132 8472 3167
rect 7290 3098 7830 3132
rect 7864 3098 7898 3132
rect 7932 3098 8472 3132
rect 7290 3063 8472 3098
rect 7290 3029 7830 3063
rect 7864 3029 7898 3063
rect 7932 3029 8472 3063
rect 7290 2994 8472 3029
rect 7290 2960 7830 2994
rect 7864 2960 7898 2994
rect 7932 2960 8472 2994
rect 7290 2925 8472 2960
rect 7290 2891 7830 2925
rect 7864 2891 7898 2925
rect 7932 2891 8472 2925
rect 7290 2856 8472 2891
rect 7290 2822 7830 2856
rect 7864 2822 7898 2856
rect 7932 2822 8472 2856
rect 7290 2787 8472 2822
rect 7290 2753 7830 2787
rect 7864 2753 7898 2787
rect 7932 2753 8472 2787
rect 7290 2718 8472 2753
rect 7290 2684 7830 2718
rect 7864 2684 7898 2718
rect 7932 2684 8472 2718
rect 7290 2649 8472 2684
rect 7290 2615 7830 2649
rect 7864 2615 7898 2649
rect 7932 2615 8472 2649
rect 7290 2580 8472 2615
rect 7290 2546 7830 2580
rect 7864 2546 7898 2580
rect 7932 2546 8472 2580
rect 7290 2511 8472 2546
rect 7290 2477 7830 2511
rect 7864 2477 7898 2511
rect 7932 2477 8472 2511
rect 7290 2442 8472 2477
rect 7290 2408 7830 2442
rect 7864 2408 7898 2442
rect 7932 2408 8472 2442
rect 7290 2373 8472 2408
rect 7290 2339 7830 2373
rect 7864 2339 7898 2373
rect 7932 2339 8472 2373
rect 7290 2304 8472 2339
rect 7290 2270 7830 2304
rect 7864 2270 7898 2304
rect 7932 2270 8472 2304
rect 7290 2235 8472 2270
rect 7290 2201 7830 2235
rect 7864 2201 7898 2235
rect 7932 2201 8472 2235
rect 7290 2166 8472 2201
rect 7290 2132 7830 2166
rect 7864 2132 7898 2166
rect 7932 2132 8472 2166
rect 7290 2097 8472 2132
rect 7290 2063 7830 2097
rect 7864 2063 7898 2097
rect 7932 2063 8472 2097
rect 7290 2028 8472 2063
rect 7290 1994 7830 2028
rect 7864 1994 7898 2028
rect 7932 1994 8472 2028
rect 7290 1959 8472 1994
rect 7290 1925 7830 1959
rect 7864 1925 7898 1959
rect 7932 1925 8472 1959
rect 7290 1890 8472 1925
rect 7290 1856 7830 1890
rect 7864 1856 7898 1890
rect 7932 1856 8472 1890
rect 7290 1821 8472 1856
rect 7290 1787 7830 1821
rect 7864 1787 7898 1821
rect 7932 1787 8472 1821
rect 7290 1752 8472 1787
rect 7290 1718 7830 1752
rect 7864 1718 7898 1752
rect 7932 1718 8472 1752
rect 7290 1683 8472 1718
rect 7290 1649 7830 1683
rect 7864 1649 7898 1683
rect 7932 1649 8472 1683
rect 7290 1614 8472 1649
rect 7290 1580 7830 1614
rect 7864 1580 7898 1614
rect 7932 1580 8472 1614
rect 7290 1545 8472 1580
rect 7290 1511 7830 1545
rect 7864 1511 7898 1545
rect 7932 1511 8472 1545
rect 7290 1476 8472 1511
rect 7290 1442 7830 1476
rect 7864 1442 7898 1476
rect 7932 1442 8472 1476
rect 7290 1407 8472 1442
rect 7290 1373 7830 1407
rect 7864 1373 7898 1407
rect 7932 1373 8472 1407
rect 7290 1338 8472 1373
rect 7290 1304 7830 1338
rect 7864 1304 7898 1338
rect 7932 1304 8472 1338
rect 7290 1269 8472 1304
rect 7290 1235 7830 1269
rect 7864 1235 7898 1269
rect 7932 1235 8472 1269
rect 7290 1155 8472 1235
tri 7290 1135 7310 1155 ne
rect 7310 1135 8452 1155
tri 8452 1135 8472 1155 nw
tri 8582 11313 8602 11333 se
rect 8602 11313 8964 11333
tri 8964 11313 8984 11333 sw
rect 8582 11233 8984 11313
rect 8582 3719 8732 11233
rect 8834 3719 8984 11233
rect 8582 3684 8984 3719
rect 8582 3650 8732 3684
rect 8766 3650 8800 3684
rect 8834 3650 8984 3684
rect 8582 3615 8984 3650
rect 8582 3581 8732 3615
rect 8766 3581 8800 3615
rect 8834 3581 8984 3615
rect 8582 3546 8984 3581
rect 8582 3512 8732 3546
rect 8766 3512 8800 3546
rect 8834 3512 8984 3546
rect 8582 3477 8984 3512
rect 8582 3443 8732 3477
rect 8766 3443 8800 3477
rect 8834 3443 8984 3477
rect 8582 3408 8984 3443
rect 8582 3374 8732 3408
rect 8766 3374 8800 3408
rect 8834 3374 8984 3408
rect 8582 3339 8984 3374
rect 8582 3305 8732 3339
rect 8766 3305 8800 3339
rect 8834 3305 8984 3339
rect 8582 3270 8984 3305
rect 8582 3236 8732 3270
rect 8766 3236 8800 3270
rect 8834 3236 8984 3270
rect 8582 3201 8984 3236
rect 8582 3167 8732 3201
rect 8766 3167 8800 3201
rect 8834 3167 8984 3201
rect 8582 3132 8984 3167
rect 8582 3098 8732 3132
rect 8766 3098 8800 3132
rect 8834 3098 8984 3132
rect 8582 3063 8984 3098
rect 8582 3029 8732 3063
rect 8766 3029 8800 3063
rect 8834 3029 8984 3063
rect 8582 2994 8984 3029
rect 8582 2960 8732 2994
rect 8766 2960 8800 2994
rect 8834 2960 8984 2994
rect 8582 2925 8984 2960
rect 8582 2891 8732 2925
rect 8766 2891 8800 2925
rect 8834 2891 8984 2925
rect 8582 2856 8984 2891
rect 8582 2822 8732 2856
rect 8766 2822 8800 2856
rect 8834 2822 8984 2856
rect 8582 2787 8984 2822
rect 8582 2753 8732 2787
rect 8766 2753 8800 2787
rect 8834 2753 8984 2787
rect 8582 2718 8984 2753
rect 8582 2684 8732 2718
rect 8766 2684 8800 2718
rect 8834 2684 8984 2718
rect 8582 2649 8984 2684
rect 8582 2615 8732 2649
rect 8766 2615 8800 2649
rect 8834 2615 8984 2649
rect 8582 2580 8984 2615
rect 8582 2546 8732 2580
rect 8766 2546 8800 2580
rect 8834 2546 8984 2580
rect 8582 2511 8984 2546
rect 8582 2477 8732 2511
rect 8766 2477 8800 2511
rect 8834 2477 8984 2511
rect 8582 2442 8984 2477
rect 8582 2408 8732 2442
rect 8766 2408 8800 2442
rect 8834 2408 8984 2442
rect 8582 2373 8984 2408
rect 8582 2339 8732 2373
rect 8766 2339 8800 2373
rect 8834 2339 8984 2373
rect 8582 2304 8984 2339
rect 8582 2270 8732 2304
rect 8766 2270 8800 2304
rect 8834 2270 8984 2304
rect 8582 2235 8984 2270
rect 8582 2201 8732 2235
rect 8766 2201 8800 2235
rect 8834 2201 8984 2235
rect 8582 2166 8984 2201
rect 8582 2132 8732 2166
rect 8766 2132 8800 2166
rect 8834 2132 8984 2166
rect 8582 2097 8984 2132
rect 8582 2063 8732 2097
rect 8766 2063 8800 2097
rect 8834 2063 8984 2097
rect 8582 2028 8984 2063
rect 8582 1994 8732 2028
rect 8766 1994 8800 2028
rect 8834 1994 8984 2028
rect 8582 1959 8984 1994
rect 8582 1925 8732 1959
rect 8766 1925 8800 1959
rect 8834 1925 8984 1959
rect 8582 1890 8984 1925
rect 8582 1856 8732 1890
rect 8766 1856 8800 1890
rect 8834 1856 8984 1890
rect 8582 1821 8984 1856
rect 8582 1787 8732 1821
rect 8766 1787 8800 1821
rect 8834 1787 8984 1821
rect 8582 1752 8984 1787
rect 8582 1718 8732 1752
rect 8766 1718 8800 1752
rect 8834 1718 8984 1752
rect 8582 1683 8984 1718
rect 8582 1649 8732 1683
rect 8766 1649 8800 1683
rect 8834 1649 8984 1683
rect 8582 1614 8984 1649
rect 8582 1580 8732 1614
rect 8766 1580 8800 1614
rect 8834 1580 8984 1614
rect 8582 1545 8984 1580
rect 8582 1511 8732 1545
rect 8766 1511 8800 1545
rect 8834 1511 8984 1545
rect 8582 1476 8984 1511
rect 8582 1442 8732 1476
rect 8766 1442 8800 1476
rect 8834 1442 8984 1476
rect 8582 1407 8984 1442
rect 8582 1373 8732 1407
rect 8766 1373 8800 1407
rect 8834 1373 8984 1407
rect 8582 1338 8984 1373
rect 8582 1304 8732 1338
rect 8766 1304 8800 1338
rect 8834 1304 8984 1338
rect 8582 1269 8984 1304
rect 8582 1235 8732 1269
rect 8766 1235 8800 1269
rect 8834 1235 8984 1269
rect 8582 1155 8984 1235
tri 8582 1135 8602 1155 ne
rect 8602 1135 8964 1155
tri 8964 1135 8984 1155 nw
tri 9094 11313 9114 11333 se
rect 9114 11313 10256 11333
tri 10256 11313 10276 11333 sw
rect 9094 11233 10276 11313
rect 9094 3719 9634 11233
rect 9736 3719 10276 11233
rect 9094 3684 10276 3719
rect 9094 3650 9634 3684
rect 9668 3650 9702 3684
rect 9736 3650 10276 3684
rect 9094 3615 10276 3650
rect 9094 3581 9634 3615
rect 9668 3581 9702 3615
rect 9736 3581 10276 3615
rect 9094 3546 10276 3581
rect 9094 3512 9634 3546
rect 9668 3512 9702 3546
rect 9736 3512 10276 3546
rect 9094 3477 10276 3512
rect 9094 3443 9634 3477
rect 9668 3443 9702 3477
rect 9736 3443 10276 3477
rect 9094 3408 10276 3443
rect 9094 3374 9634 3408
rect 9668 3374 9702 3408
rect 9736 3374 10276 3408
rect 9094 3339 10276 3374
rect 9094 3305 9634 3339
rect 9668 3305 9702 3339
rect 9736 3305 10276 3339
rect 9094 3270 10276 3305
rect 9094 3236 9634 3270
rect 9668 3236 9702 3270
rect 9736 3236 10276 3270
rect 9094 3201 10276 3236
rect 9094 3167 9634 3201
rect 9668 3167 9702 3201
rect 9736 3167 10276 3201
rect 9094 3132 10276 3167
rect 9094 3098 9634 3132
rect 9668 3098 9702 3132
rect 9736 3098 10276 3132
rect 9094 3063 10276 3098
rect 9094 3029 9634 3063
rect 9668 3029 9702 3063
rect 9736 3029 10276 3063
rect 9094 2994 10276 3029
rect 9094 2960 9634 2994
rect 9668 2960 9702 2994
rect 9736 2960 10276 2994
rect 9094 2925 10276 2960
rect 9094 2891 9634 2925
rect 9668 2891 9702 2925
rect 9736 2891 10276 2925
rect 9094 2856 10276 2891
rect 9094 2822 9634 2856
rect 9668 2822 9702 2856
rect 9736 2822 10276 2856
rect 9094 2787 10276 2822
rect 9094 2753 9634 2787
rect 9668 2753 9702 2787
rect 9736 2753 10276 2787
rect 9094 2718 10276 2753
rect 9094 2684 9634 2718
rect 9668 2684 9702 2718
rect 9736 2684 10276 2718
rect 9094 2649 10276 2684
rect 9094 2615 9634 2649
rect 9668 2615 9702 2649
rect 9736 2615 10276 2649
rect 9094 2580 10276 2615
rect 9094 2546 9634 2580
rect 9668 2546 9702 2580
rect 9736 2546 10276 2580
rect 9094 2511 10276 2546
rect 9094 2477 9634 2511
rect 9668 2477 9702 2511
rect 9736 2477 10276 2511
rect 9094 2442 10276 2477
rect 9094 2408 9634 2442
rect 9668 2408 9702 2442
rect 9736 2408 10276 2442
rect 9094 2373 10276 2408
rect 9094 2339 9634 2373
rect 9668 2339 9702 2373
rect 9736 2339 10276 2373
rect 9094 2304 10276 2339
rect 9094 2270 9634 2304
rect 9668 2270 9702 2304
rect 9736 2270 10276 2304
rect 9094 2235 10276 2270
rect 9094 2201 9634 2235
rect 9668 2201 9702 2235
rect 9736 2201 10276 2235
rect 9094 2166 10276 2201
rect 9094 2132 9634 2166
rect 9668 2132 9702 2166
rect 9736 2132 10276 2166
rect 9094 2097 10276 2132
rect 9094 2063 9634 2097
rect 9668 2063 9702 2097
rect 9736 2063 10276 2097
rect 9094 2028 10276 2063
rect 9094 1994 9634 2028
rect 9668 1994 9702 2028
rect 9736 1994 10276 2028
rect 9094 1959 10276 1994
rect 9094 1925 9634 1959
rect 9668 1925 9702 1959
rect 9736 1925 10276 1959
rect 9094 1890 10276 1925
rect 9094 1856 9634 1890
rect 9668 1856 9702 1890
rect 9736 1856 10276 1890
rect 9094 1821 10276 1856
rect 9094 1787 9634 1821
rect 9668 1787 9702 1821
rect 9736 1787 10276 1821
rect 9094 1752 10276 1787
rect 9094 1718 9634 1752
rect 9668 1718 9702 1752
rect 9736 1718 10276 1752
rect 9094 1683 10276 1718
rect 9094 1649 9634 1683
rect 9668 1649 9702 1683
rect 9736 1649 10276 1683
rect 9094 1614 10276 1649
rect 9094 1580 9634 1614
rect 9668 1580 9702 1614
rect 9736 1580 10276 1614
rect 9094 1545 10276 1580
rect 9094 1511 9634 1545
rect 9668 1511 9702 1545
rect 9736 1511 10276 1545
rect 9094 1476 10276 1511
rect 9094 1442 9634 1476
rect 9668 1442 9702 1476
rect 9736 1442 10276 1476
rect 9094 1407 10276 1442
rect 9094 1373 9634 1407
rect 9668 1373 9702 1407
rect 9736 1373 10276 1407
rect 9094 1338 10276 1373
rect 9094 1304 9634 1338
rect 9668 1304 9702 1338
rect 9736 1304 10276 1338
rect 9094 1269 10276 1304
rect 9094 1235 9634 1269
rect 9668 1235 9702 1269
rect 9736 1235 10276 1269
rect 9094 1155 10276 1235
tri 9094 1135 9114 1155 ne
rect 9114 1135 10256 1155
tri 10256 1135 10276 1155 nw
tri 10386 11313 10406 11333 se
rect 10406 11313 10768 11333
tri 10768 11313 10788 11333 sw
rect 10386 11233 10788 11313
rect 10386 3719 10536 11233
rect 10638 3719 10788 11233
rect 10386 3684 10788 3719
rect 10386 3650 10536 3684
rect 10570 3650 10604 3684
rect 10638 3650 10788 3684
rect 10386 3615 10788 3650
rect 10386 3581 10536 3615
rect 10570 3581 10604 3615
rect 10638 3581 10788 3615
rect 10386 3546 10788 3581
rect 10386 3512 10536 3546
rect 10570 3512 10604 3546
rect 10638 3512 10788 3546
rect 10386 3477 10788 3512
rect 10386 3443 10536 3477
rect 10570 3443 10604 3477
rect 10638 3443 10788 3477
rect 10386 3408 10788 3443
rect 10386 3374 10536 3408
rect 10570 3374 10604 3408
rect 10638 3374 10788 3408
rect 10386 3339 10788 3374
rect 10386 3305 10536 3339
rect 10570 3305 10604 3339
rect 10638 3305 10788 3339
rect 10386 3270 10788 3305
rect 10386 3236 10536 3270
rect 10570 3236 10604 3270
rect 10638 3236 10788 3270
rect 10386 3201 10788 3236
rect 10386 3167 10536 3201
rect 10570 3167 10604 3201
rect 10638 3167 10788 3201
rect 10386 3132 10788 3167
rect 10386 3098 10536 3132
rect 10570 3098 10604 3132
rect 10638 3098 10788 3132
rect 10386 3063 10788 3098
rect 10386 3029 10536 3063
rect 10570 3029 10604 3063
rect 10638 3029 10788 3063
rect 10386 2994 10788 3029
rect 10386 2960 10536 2994
rect 10570 2960 10604 2994
rect 10638 2960 10788 2994
rect 10386 2925 10788 2960
rect 10386 2891 10536 2925
rect 10570 2891 10604 2925
rect 10638 2891 10788 2925
rect 10386 2856 10788 2891
rect 10386 2822 10536 2856
rect 10570 2822 10604 2856
rect 10638 2822 10788 2856
rect 10386 2787 10788 2822
rect 10386 2753 10536 2787
rect 10570 2753 10604 2787
rect 10638 2753 10788 2787
rect 10386 2718 10788 2753
rect 10386 2684 10536 2718
rect 10570 2684 10604 2718
rect 10638 2684 10788 2718
rect 10386 2649 10788 2684
rect 10386 2615 10536 2649
rect 10570 2615 10604 2649
rect 10638 2615 10788 2649
rect 10386 2580 10788 2615
rect 10386 2546 10536 2580
rect 10570 2546 10604 2580
rect 10638 2546 10788 2580
rect 10386 2511 10788 2546
rect 10386 2477 10536 2511
rect 10570 2477 10604 2511
rect 10638 2477 10788 2511
rect 10386 2442 10788 2477
rect 10386 2408 10536 2442
rect 10570 2408 10604 2442
rect 10638 2408 10788 2442
rect 10386 2373 10788 2408
rect 10386 2339 10536 2373
rect 10570 2339 10604 2373
rect 10638 2339 10788 2373
rect 10386 2304 10788 2339
rect 10386 2270 10536 2304
rect 10570 2270 10604 2304
rect 10638 2270 10788 2304
rect 10386 2235 10788 2270
rect 10386 2201 10536 2235
rect 10570 2201 10604 2235
rect 10638 2201 10788 2235
rect 10386 2166 10788 2201
rect 10386 2132 10536 2166
rect 10570 2132 10604 2166
rect 10638 2132 10788 2166
rect 10386 2097 10788 2132
rect 10386 2063 10536 2097
rect 10570 2063 10604 2097
rect 10638 2063 10788 2097
rect 10386 2028 10788 2063
rect 10386 1994 10536 2028
rect 10570 1994 10604 2028
rect 10638 1994 10788 2028
rect 10386 1959 10788 1994
rect 10386 1925 10536 1959
rect 10570 1925 10604 1959
rect 10638 1925 10788 1959
rect 10386 1890 10788 1925
rect 10386 1856 10536 1890
rect 10570 1856 10604 1890
rect 10638 1856 10788 1890
rect 10386 1821 10788 1856
rect 10386 1787 10536 1821
rect 10570 1787 10604 1821
rect 10638 1787 10788 1821
rect 10386 1752 10788 1787
rect 10386 1718 10536 1752
rect 10570 1718 10604 1752
rect 10638 1718 10788 1752
rect 10386 1683 10788 1718
rect 10386 1649 10536 1683
rect 10570 1649 10604 1683
rect 10638 1649 10788 1683
rect 10386 1614 10788 1649
rect 10386 1580 10536 1614
rect 10570 1580 10604 1614
rect 10638 1580 10788 1614
rect 10386 1545 10788 1580
rect 10386 1511 10536 1545
rect 10570 1511 10604 1545
rect 10638 1511 10788 1545
rect 10386 1476 10788 1511
rect 10386 1442 10536 1476
rect 10570 1442 10604 1476
rect 10638 1442 10788 1476
rect 10386 1407 10788 1442
rect 10386 1373 10536 1407
rect 10570 1373 10604 1407
rect 10638 1373 10788 1407
rect 10386 1338 10788 1373
rect 10386 1304 10536 1338
rect 10570 1304 10604 1338
rect 10638 1304 10788 1338
rect 10386 1269 10788 1304
rect 10386 1235 10536 1269
rect 10570 1235 10604 1269
rect 10638 1235 10788 1269
rect 10386 1155 10788 1235
tri 10386 1135 10406 1155 ne
rect 10406 1135 10768 1155
tri 10768 1135 10788 1155 nw
tri 10898 11313 10918 11333 se
rect 10918 11313 12060 11333
tri 12060 11313 12080 11333 sw
rect 10898 11233 12080 11313
rect 10898 3719 11438 11233
rect 11540 3719 12080 11233
rect 10898 3684 12080 3719
rect 10898 3650 11438 3684
rect 11472 3650 11506 3684
rect 11540 3650 12080 3684
rect 10898 3615 12080 3650
rect 10898 3581 11438 3615
rect 11472 3581 11506 3615
rect 11540 3581 12080 3615
rect 10898 3546 12080 3581
rect 10898 3512 11438 3546
rect 11472 3512 11506 3546
rect 11540 3512 12080 3546
rect 10898 3477 12080 3512
rect 10898 3443 11438 3477
rect 11472 3443 11506 3477
rect 11540 3443 12080 3477
rect 10898 3408 12080 3443
rect 10898 3374 11438 3408
rect 11472 3374 11506 3408
rect 11540 3374 12080 3408
rect 10898 3339 12080 3374
rect 10898 3305 11438 3339
rect 11472 3305 11506 3339
rect 11540 3305 12080 3339
rect 10898 3270 12080 3305
rect 10898 3236 11438 3270
rect 11472 3236 11506 3270
rect 11540 3236 12080 3270
rect 10898 3201 12080 3236
rect 10898 3167 11438 3201
rect 11472 3167 11506 3201
rect 11540 3167 12080 3201
rect 10898 3132 12080 3167
rect 10898 3098 11438 3132
rect 11472 3098 11506 3132
rect 11540 3098 12080 3132
rect 10898 3063 12080 3098
rect 10898 3029 11438 3063
rect 11472 3029 11506 3063
rect 11540 3029 12080 3063
rect 10898 2994 12080 3029
rect 10898 2960 11438 2994
rect 11472 2960 11506 2994
rect 11540 2960 12080 2994
rect 10898 2925 12080 2960
rect 10898 2891 11438 2925
rect 11472 2891 11506 2925
rect 11540 2891 12080 2925
rect 10898 2856 12080 2891
rect 10898 2822 11438 2856
rect 11472 2822 11506 2856
rect 11540 2822 12080 2856
rect 10898 2787 12080 2822
rect 10898 2753 11438 2787
rect 11472 2753 11506 2787
rect 11540 2753 12080 2787
rect 10898 2718 12080 2753
rect 10898 2684 11438 2718
rect 11472 2684 11506 2718
rect 11540 2684 12080 2718
rect 10898 2649 12080 2684
rect 10898 2615 11438 2649
rect 11472 2615 11506 2649
rect 11540 2615 12080 2649
rect 10898 2580 12080 2615
rect 10898 2546 11438 2580
rect 11472 2546 11506 2580
rect 11540 2546 12080 2580
rect 10898 2511 12080 2546
rect 10898 2477 11438 2511
rect 11472 2477 11506 2511
rect 11540 2477 12080 2511
rect 10898 2442 12080 2477
rect 10898 2408 11438 2442
rect 11472 2408 11506 2442
rect 11540 2408 12080 2442
rect 10898 2373 12080 2408
rect 10898 2339 11438 2373
rect 11472 2339 11506 2373
rect 11540 2339 12080 2373
rect 10898 2304 12080 2339
rect 10898 2270 11438 2304
rect 11472 2270 11506 2304
rect 11540 2270 12080 2304
rect 10898 2235 12080 2270
rect 10898 2201 11438 2235
rect 11472 2201 11506 2235
rect 11540 2201 12080 2235
rect 10898 2166 12080 2201
rect 10898 2132 11438 2166
rect 11472 2132 11506 2166
rect 11540 2132 12080 2166
rect 10898 2097 12080 2132
rect 10898 2063 11438 2097
rect 11472 2063 11506 2097
rect 11540 2063 12080 2097
rect 10898 2028 12080 2063
rect 10898 1994 11438 2028
rect 11472 1994 11506 2028
rect 11540 1994 12080 2028
rect 10898 1959 12080 1994
rect 10898 1925 11438 1959
rect 11472 1925 11506 1959
rect 11540 1925 12080 1959
rect 10898 1890 12080 1925
rect 10898 1856 11438 1890
rect 11472 1856 11506 1890
rect 11540 1856 12080 1890
rect 10898 1821 12080 1856
rect 10898 1787 11438 1821
rect 11472 1787 11506 1821
rect 11540 1787 12080 1821
rect 10898 1752 12080 1787
rect 10898 1718 11438 1752
rect 11472 1718 11506 1752
rect 11540 1718 12080 1752
rect 10898 1683 12080 1718
rect 10898 1649 11438 1683
rect 11472 1649 11506 1683
rect 11540 1649 12080 1683
rect 10898 1614 12080 1649
rect 10898 1580 11438 1614
rect 11472 1580 11506 1614
rect 11540 1580 12080 1614
rect 10898 1545 12080 1580
rect 10898 1511 11438 1545
rect 11472 1511 11506 1545
rect 11540 1511 12080 1545
rect 10898 1476 12080 1511
rect 10898 1442 11438 1476
rect 11472 1442 11506 1476
rect 11540 1442 12080 1476
rect 10898 1407 12080 1442
rect 10898 1373 11438 1407
rect 11472 1373 11506 1407
rect 11540 1373 12080 1407
rect 10898 1338 12080 1373
rect 10898 1304 11438 1338
rect 11472 1304 11506 1338
rect 11540 1304 12080 1338
rect 10898 1269 12080 1304
rect 10898 1235 11438 1269
rect 11472 1235 11506 1269
rect 11540 1235 12080 1269
rect 10898 1155 12080 1235
tri 10898 1135 10918 1155 ne
rect 10918 1135 12060 1155
tri 12060 1135 12080 1155 nw
tri 12190 11313 12210 11333 se
rect 12210 11313 12572 11333
tri 12572 11313 12592 11333 sw
rect 12190 11233 12592 11313
rect 12190 3719 12340 11233
rect 12442 3719 12592 11233
rect 12190 3684 12592 3719
rect 12190 3650 12340 3684
rect 12374 3650 12408 3684
rect 12442 3650 12592 3684
rect 12190 3615 12592 3650
rect 12190 3581 12340 3615
rect 12374 3581 12408 3615
rect 12442 3581 12592 3615
rect 12190 3546 12592 3581
rect 12190 3512 12340 3546
rect 12374 3512 12408 3546
rect 12442 3512 12592 3546
rect 12190 3477 12592 3512
rect 12190 3443 12340 3477
rect 12374 3443 12408 3477
rect 12442 3443 12592 3477
rect 12190 3408 12592 3443
rect 12190 3374 12340 3408
rect 12374 3374 12408 3408
rect 12442 3374 12592 3408
rect 12190 3339 12592 3374
rect 12190 3305 12340 3339
rect 12374 3305 12408 3339
rect 12442 3305 12592 3339
rect 12190 3270 12592 3305
rect 12190 3236 12340 3270
rect 12374 3236 12408 3270
rect 12442 3236 12592 3270
rect 12190 3201 12592 3236
rect 12190 3167 12340 3201
rect 12374 3167 12408 3201
rect 12442 3167 12592 3201
rect 12190 3132 12592 3167
rect 12190 3098 12340 3132
rect 12374 3098 12408 3132
rect 12442 3098 12592 3132
rect 12190 3063 12592 3098
rect 12190 3029 12340 3063
rect 12374 3029 12408 3063
rect 12442 3029 12592 3063
rect 12190 2994 12592 3029
rect 12190 2960 12340 2994
rect 12374 2960 12408 2994
rect 12442 2960 12592 2994
rect 12190 2925 12592 2960
rect 12190 2891 12340 2925
rect 12374 2891 12408 2925
rect 12442 2891 12592 2925
rect 12190 2856 12592 2891
rect 12190 2822 12340 2856
rect 12374 2822 12408 2856
rect 12442 2822 12592 2856
rect 12190 2787 12592 2822
rect 12190 2753 12340 2787
rect 12374 2753 12408 2787
rect 12442 2753 12592 2787
rect 12190 2718 12592 2753
rect 12190 2684 12340 2718
rect 12374 2684 12408 2718
rect 12442 2684 12592 2718
rect 12190 2649 12592 2684
rect 12190 2615 12340 2649
rect 12374 2615 12408 2649
rect 12442 2615 12592 2649
rect 12190 2580 12592 2615
rect 12190 2546 12340 2580
rect 12374 2546 12408 2580
rect 12442 2546 12592 2580
rect 12190 2511 12592 2546
rect 12190 2477 12340 2511
rect 12374 2477 12408 2511
rect 12442 2477 12592 2511
rect 12190 2442 12592 2477
rect 12190 2408 12340 2442
rect 12374 2408 12408 2442
rect 12442 2408 12592 2442
rect 12190 2373 12592 2408
rect 12190 2339 12340 2373
rect 12374 2339 12408 2373
rect 12442 2339 12592 2373
rect 12190 2304 12592 2339
rect 12190 2270 12340 2304
rect 12374 2270 12408 2304
rect 12442 2270 12592 2304
rect 12190 2235 12592 2270
rect 12190 2201 12340 2235
rect 12374 2201 12408 2235
rect 12442 2201 12592 2235
rect 12190 2166 12592 2201
rect 12190 2132 12340 2166
rect 12374 2132 12408 2166
rect 12442 2132 12592 2166
rect 12190 2097 12592 2132
rect 12190 2063 12340 2097
rect 12374 2063 12408 2097
rect 12442 2063 12592 2097
rect 12190 2028 12592 2063
rect 12190 1994 12340 2028
rect 12374 1994 12408 2028
rect 12442 1994 12592 2028
rect 12190 1959 12592 1994
rect 12190 1925 12340 1959
rect 12374 1925 12408 1959
rect 12442 1925 12592 1959
rect 12190 1890 12592 1925
rect 12190 1856 12340 1890
rect 12374 1856 12408 1890
rect 12442 1856 12592 1890
rect 12190 1821 12592 1856
rect 12190 1787 12340 1821
rect 12374 1787 12408 1821
rect 12442 1787 12592 1821
rect 12190 1752 12592 1787
rect 12190 1718 12340 1752
rect 12374 1718 12408 1752
rect 12442 1718 12592 1752
rect 12190 1683 12592 1718
rect 12190 1649 12340 1683
rect 12374 1649 12408 1683
rect 12442 1649 12592 1683
rect 12190 1614 12592 1649
rect 12190 1580 12340 1614
rect 12374 1580 12408 1614
rect 12442 1580 12592 1614
rect 12190 1545 12592 1580
rect 12190 1511 12340 1545
rect 12374 1511 12408 1545
rect 12442 1511 12592 1545
rect 12190 1476 12592 1511
rect 12190 1442 12340 1476
rect 12374 1442 12408 1476
rect 12442 1442 12592 1476
rect 12190 1407 12592 1442
rect 12190 1373 12340 1407
rect 12374 1373 12408 1407
rect 12442 1373 12592 1407
rect 12190 1338 12592 1373
rect 12190 1304 12340 1338
rect 12374 1304 12408 1338
rect 12442 1304 12592 1338
rect 12190 1269 12592 1304
rect 12190 1235 12340 1269
rect 12374 1235 12408 1269
rect 12442 1235 12592 1269
rect 12190 1155 12592 1235
tri 12190 1135 12210 1155 ne
rect 12210 1135 12572 1155
tri 12572 1135 12592 1155 nw
tri 12702 11313 12722 11333 se
rect 12722 11313 13864 11333
tri 13864 11313 13884 11333 sw
rect 12702 11233 13884 11313
rect 12702 3719 13242 11233
rect 13344 3719 13884 11233
rect 12702 3684 13884 3719
rect 12702 3650 13242 3684
rect 13276 3650 13310 3684
rect 13344 3650 13884 3684
rect 12702 3615 13884 3650
rect 12702 3581 13242 3615
rect 13276 3581 13310 3615
rect 13344 3581 13884 3615
rect 12702 3546 13884 3581
rect 12702 3512 13242 3546
rect 13276 3512 13310 3546
rect 13344 3512 13884 3546
rect 12702 3477 13884 3512
rect 12702 3443 13242 3477
rect 13276 3443 13310 3477
rect 13344 3443 13884 3477
rect 12702 3408 13884 3443
rect 12702 3374 13242 3408
rect 13276 3374 13310 3408
rect 13344 3374 13884 3408
rect 12702 3339 13884 3374
rect 12702 3305 13242 3339
rect 13276 3305 13310 3339
rect 13344 3305 13884 3339
rect 12702 3270 13884 3305
rect 12702 3236 13242 3270
rect 13276 3236 13310 3270
rect 13344 3236 13884 3270
rect 12702 3201 13884 3236
rect 12702 3167 13242 3201
rect 13276 3167 13310 3201
rect 13344 3167 13884 3201
rect 12702 3132 13884 3167
rect 12702 3098 13242 3132
rect 13276 3098 13310 3132
rect 13344 3098 13884 3132
rect 12702 3063 13884 3098
rect 12702 3029 13242 3063
rect 13276 3029 13310 3063
rect 13344 3029 13884 3063
rect 12702 2994 13884 3029
rect 12702 2960 13242 2994
rect 13276 2960 13310 2994
rect 13344 2960 13884 2994
rect 12702 2925 13884 2960
rect 12702 2891 13242 2925
rect 13276 2891 13310 2925
rect 13344 2891 13884 2925
rect 12702 2856 13884 2891
rect 12702 2822 13242 2856
rect 13276 2822 13310 2856
rect 13344 2822 13884 2856
rect 12702 2787 13884 2822
rect 12702 2753 13242 2787
rect 13276 2753 13310 2787
rect 13344 2753 13884 2787
rect 12702 2718 13884 2753
rect 12702 2684 13242 2718
rect 13276 2684 13310 2718
rect 13344 2684 13884 2718
rect 12702 2649 13884 2684
rect 12702 2615 13242 2649
rect 13276 2615 13310 2649
rect 13344 2615 13884 2649
rect 12702 2580 13884 2615
rect 12702 2546 13242 2580
rect 13276 2546 13310 2580
rect 13344 2546 13884 2580
rect 12702 2511 13884 2546
rect 12702 2477 13242 2511
rect 13276 2477 13310 2511
rect 13344 2477 13884 2511
rect 12702 2442 13884 2477
rect 12702 2408 13242 2442
rect 13276 2408 13310 2442
rect 13344 2408 13884 2442
rect 12702 2373 13884 2408
rect 12702 2339 13242 2373
rect 13276 2339 13310 2373
rect 13344 2339 13884 2373
rect 12702 2304 13884 2339
rect 12702 2270 13242 2304
rect 13276 2270 13310 2304
rect 13344 2270 13884 2304
rect 12702 2235 13884 2270
rect 12702 2201 13242 2235
rect 13276 2201 13310 2235
rect 13344 2201 13884 2235
rect 12702 2166 13884 2201
rect 12702 2132 13242 2166
rect 13276 2132 13310 2166
rect 13344 2132 13884 2166
rect 12702 2097 13884 2132
rect 12702 2063 13242 2097
rect 13276 2063 13310 2097
rect 13344 2063 13884 2097
rect 12702 2028 13884 2063
rect 12702 1994 13242 2028
rect 13276 1994 13310 2028
rect 13344 1994 13884 2028
rect 12702 1959 13884 1994
rect 12702 1925 13242 1959
rect 13276 1925 13310 1959
rect 13344 1925 13884 1959
rect 12702 1890 13884 1925
rect 12702 1856 13242 1890
rect 13276 1856 13310 1890
rect 13344 1856 13884 1890
rect 12702 1821 13884 1856
rect 12702 1787 13242 1821
rect 13276 1787 13310 1821
rect 13344 1787 13884 1821
rect 12702 1752 13884 1787
rect 12702 1718 13242 1752
rect 13276 1718 13310 1752
rect 13344 1718 13884 1752
rect 12702 1683 13884 1718
rect 12702 1649 13242 1683
rect 13276 1649 13310 1683
rect 13344 1649 13884 1683
rect 12702 1614 13884 1649
rect 12702 1580 13242 1614
rect 13276 1580 13310 1614
rect 13344 1580 13884 1614
rect 12702 1545 13884 1580
rect 12702 1511 13242 1545
rect 13276 1511 13310 1545
rect 13344 1511 13884 1545
rect 12702 1476 13884 1511
rect 12702 1442 13242 1476
rect 13276 1442 13310 1476
rect 13344 1442 13884 1476
rect 12702 1407 13884 1442
rect 12702 1373 13242 1407
rect 13276 1373 13310 1407
rect 13344 1373 13884 1407
rect 12702 1338 13884 1373
rect 12702 1304 13242 1338
rect 13276 1304 13310 1338
rect 13344 1304 13884 1338
rect 12702 1269 13884 1304
rect 12702 1235 13242 1269
rect 13276 1235 13310 1269
rect 13344 1235 13884 1269
rect 12702 1155 13884 1235
tri 12702 1135 12722 1155 ne
rect 12722 1135 13864 1155
tri 13864 1135 13884 1155 nw
tri 13994 11313 14014 11333 se
rect 14014 11313 14386 11333
rect 13994 11233 14386 11313
rect 13994 3719 14144 11233
rect 14246 3719 14386 11233
rect 13994 3684 14386 3719
rect 13994 3650 14144 3684
rect 14178 3650 14212 3684
rect 14246 3650 14386 3684
rect 13994 3615 14386 3650
rect 13994 3581 14144 3615
rect 14178 3581 14212 3615
rect 14246 3581 14386 3615
rect 13994 3546 14386 3581
rect 13994 3512 14144 3546
rect 14178 3512 14212 3546
rect 14246 3512 14386 3546
rect 13994 3477 14386 3512
rect 13994 3443 14144 3477
rect 14178 3443 14212 3477
rect 14246 3443 14386 3477
rect 13994 3408 14386 3443
rect 13994 3374 14144 3408
rect 14178 3374 14212 3408
rect 14246 3374 14386 3408
rect 13994 3339 14386 3374
rect 13994 3305 14144 3339
rect 14178 3305 14212 3339
rect 14246 3305 14386 3339
rect 13994 3270 14386 3305
rect 13994 3236 14144 3270
rect 14178 3236 14212 3270
rect 14246 3236 14386 3270
rect 13994 3201 14386 3236
rect 13994 3167 14144 3201
rect 14178 3167 14212 3201
rect 14246 3167 14386 3201
rect 13994 3132 14386 3167
rect 13994 3098 14144 3132
rect 14178 3098 14212 3132
rect 14246 3098 14386 3132
rect 13994 3063 14386 3098
rect 13994 3029 14144 3063
rect 14178 3029 14212 3063
rect 14246 3029 14386 3063
rect 13994 2994 14386 3029
rect 13994 2960 14144 2994
rect 14178 2960 14212 2994
rect 14246 2960 14386 2994
rect 13994 2925 14386 2960
rect 13994 2891 14144 2925
rect 14178 2891 14212 2925
rect 14246 2891 14386 2925
rect 13994 2856 14386 2891
rect 13994 2822 14144 2856
rect 14178 2822 14212 2856
rect 14246 2822 14386 2856
rect 13994 2787 14386 2822
rect 13994 2753 14144 2787
rect 14178 2753 14212 2787
rect 14246 2753 14386 2787
rect 13994 2718 14386 2753
rect 13994 2684 14144 2718
rect 14178 2684 14212 2718
rect 14246 2684 14386 2718
rect 13994 2649 14386 2684
rect 13994 2615 14144 2649
rect 14178 2615 14212 2649
rect 14246 2615 14386 2649
rect 13994 2580 14386 2615
rect 13994 2546 14144 2580
rect 14178 2546 14212 2580
rect 14246 2546 14386 2580
rect 13994 2511 14386 2546
rect 13994 2477 14144 2511
rect 14178 2477 14212 2511
rect 14246 2477 14386 2511
rect 13994 2442 14386 2477
rect 13994 2408 14144 2442
rect 14178 2408 14212 2442
rect 14246 2408 14386 2442
rect 13994 2373 14386 2408
rect 13994 2339 14144 2373
rect 14178 2339 14212 2373
rect 14246 2339 14386 2373
rect 13994 2304 14386 2339
rect 13994 2270 14144 2304
rect 14178 2270 14212 2304
rect 14246 2270 14386 2304
rect 13994 2235 14386 2270
rect 13994 2201 14144 2235
rect 14178 2201 14212 2235
rect 14246 2201 14386 2235
rect 13994 2166 14386 2201
rect 13994 2132 14144 2166
rect 14178 2132 14212 2166
rect 14246 2132 14386 2166
rect 13994 2097 14386 2132
rect 13994 2063 14144 2097
rect 14178 2063 14212 2097
rect 14246 2063 14386 2097
rect 13994 2028 14386 2063
rect 13994 1994 14144 2028
rect 14178 1994 14212 2028
rect 14246 1994 14386 2028
rect 13994 1959 14386 1994
rect 13994 1925 14144 1959
rect 14178 1925 14212 1959
rect 14246 1925 14386 1959
rect 13994 1890 14386 1925
rect 13994 1856 14144 1890
rect 14178 1856 14212 1890
rect 14246 1856 14386 1890
rect 13994 1821 14386 1856
rect 13994 1787 14144 1821
rect 14178 1787 14212 1821
rect 14246 1787 14386 1821
rect 13994 1752 14386 1787
rect 13994 1718 14144 1752
rect 14178 1718 14212 1752
rect 14246 1718 14386 1752
rect 13994 1683 14386 1718
rect 13994 1649 14144 1683
rect 14178 1649 14212 1683
rect 14246 1649 14386 1683
rect 13994 1614 14386 1649
rect 13994 1580 14144 1614
rect 14178 1580 14212 1614
rect 14246 1580 14386 1614
rect 13994 1545 14386 1580
rect 13994 1511 14144 1545
rect 14178 1511 14212 1545
rect 14246 1511 14386 1545
rect 13994 1476 14386 1511
rect 13994 1442 14144 1476
rect 14178 1442 14212 1476
rect 14246 1442 14386 1476
rect 13994 1407 14386 1442
rect 13994 1373 14144 1407
rect 14178 1373 14212 1407
rect 14246 1373 14386 1407
rect 13994 1338 14386 1373
rect 13994 1304 14144 1338
rect 14178 1304 14212 1338
rect 14246 1304 14386 1338
rect 13994 1269 14386 1304
rect 13994 1235 14144 1269
rect 14178 1235 14212 1269
rect 14246 1235 14386 1269
rect 13994 1155 14386 1235
tri 13994 1135 14014 1155 ne
rect 14014 1135 14386 1155
<< mvndiffc >>
rect -3896 3719 -3794 11233
rect -3896 3650 -3862 3684
rect -3828 3650 -3794 3684
rect -3896 3581 -3862 3615
rect -3828 3581 -3794 3615
rect -3896 3512 -3862 3546
rect -3828 3512 -3794 3546
rect -3896 3443 -3862 3477
rect -3828 3443 -3794 3477
rect -3896 3374 -3862 3408
rect -3828 3374 -3794 3408
rect -3896 3305 -3862 3339
rect -3828 3305 -3794 3339
rect -3896 3236 -3862 3270
rect -3828 3236 -3794 3270
rect -3896 3167 -3862 3201
rect -3828 3167 -3794 3201
rect -3896 3098 -3862 3132
rect -3828 3098 -3794 3132
rect -3896 3029 -3862 3063
rect -3828 3029 -3794 3063
rect -3896 2960 -3862 2994
rect -3828 2960 -3794 2994
rect -3896 2891 -3862 2925
rect -3828 2891 -3794 2925
rect -3896 2822 -3862 2856
rect -3828 2822 -3794 2856
rect -3896 2753 -3862 2787
rect -3828 2753 -3794 2787
rect -3896 2684 -3862 2718
rect -3828 2684 -3794 2718
rect -3896 2615 -3862 2649
rect -3828 2615 -3794 2649
rect -3896 2546 -3862 2580
rect -3828 2546 -3794 2580
rect -3896 2477 -3862 2511
rect -3828 2477 -3794 2511
rect -3896 2408 -3862 2442
rect -3828 2408 -3794 2442
rect -3896 2339 -3862 2373
rect -3828 2339 -3794 2373
rect -3896 2270 -3862 2304
rect -3828 2270 -3794 2304
rect -3896 2201 -3862 2235
rect -3828 2201 -3794 2235
rect -3896 2132 -3862 2166
rect -3828 2132 -3794 2166
rect -3896 2063 -3862 2097
rect -3828 2063 -3794 2097
rect -3896 1994 -3862 2028
rect -3828 1994 -3794 2028
rect -3896 1925 -3862 1959
rect -3828 1925 -3794 1959
rect -3896 1856 -3862 1890
rect -3828 1856 -3794 1890
rect -3896 1787 -3862 1821
rect -3828 1787 -3794 1821
rect -3896 1718 -3862 1752
rect -3828 1718 -3794 1752
rect -3896 1649 -3862 1683
rect -3828 1649 -3794 1683
rect -3896 1580 -3862 1614
rect -3828 1580 -3794 1614
rect -3896 1511 -3862 1545
rect -3828 1511 -3794 1545
rect -3896 1442 -3862 1476
rect -3828 1442 -3794 1476
rect -3896 1373 -3862 1407
rect -3828 1373 -3794 1407
rect -3896 1304 -3862 1338
rect -3828 1304 -3794 1338
rect -3896 1235 -3862 1269
rect -3828 1235 -3794 1269
rect -2994 3719 -2892 11233
rect -2994 3650 -2960 3684
rect -2926 3650 -2892 3684
rect -2994 3581 -2960 3615
rect -2926 3581 -2892 3615
rect -2994 3512 -2960 3546
rect -2926 3512 -2892 3546
rect -2994 3443 -2960 3477
rect -2926 3443 -2892 3477
rect -2994 3374 -2960 3408
rect -2926 3374 -2892 3408
rect -2994 3305 -2960 3339
rect -2926 3305 -2892 3339
rect -2994 3236 -2960 3270
rect -2926 3236 -2892 3270
rect -2994 3167 -2960 3201
rect -2926 3167 -2892 3201
rect -2994 3098 -2960 3132
rect -2926 3098 -2892 3132
rect -2994 3029 -2960 3063
rect -2926 3029 -2892 3063
rect -2994 2960 -2960 2994
rect -2926 2960 -2892 2994
rect -2994 2891 -2960 2925
rect -2926 2891 -2892 2925
rect -2994 2822 -2960 2856
rect -2926 2822 -2892 2856
rect -2994 2753 -2960 2787
rect -2926 2753 -2892 2787
rect -2994 2684 -2960 2718
rect -2926 2684 -2892 2718
rect -2994 2615 -2960 2649
rect -2926 2615 -2892 2649
rect -2994 2546 -2960 2580
rect -2926 2546 -2892 2580
rect -2994 2477 -2960 2511
rect -2926 2477 -2892 2511
rect -2994 2408 -2960 2442
rect -2926 2408 -2892 2442
rect -2994 2339 -2960 2373
rect -2926 2339 -2892 2373
rect -2994 2270 -2960 2304
rect -2926 2270 -2892 2304
rect -2994 2201 -2960 2235
rect -2926 2201 -2892 2235
rect -2994 2132 -2960 2166
rect -2926 2132 -2892 2166
rect -2994 2063 -2960 2097
rect -2926 2063 -2892 2097
rect -2994 1994 -2960 2028
rect -2926 1994 -2892 2028
rect -2994 1925 -2960 1959
rect -2926 1925 -2892 1959
rect -2994 1856 -2960 1890
rect -2926 1856 -2892 1890
rect -2994 1787 -2960 1821
rect -2926 1787 -2892 1821
rect -2994 1718 -2960 1752
rect -2926 1718 -2892 1752
rect -2994 1649 -2960 1683
rect -2926 1649 -2892 1683
rect -2994 1580 -2960 1614
rect -2926 1580 -2892 1614
rect -2994 1511 -2960 1545
rect -2926 1511 -2892 1545
rect -2994 1442 -2960 1476
rect -2926 1442 -2892 1476
rect -2994 1373 -2960 1407
rect -2926 1373 -2892 1407
rect -2994 1304 -2960 1338
rect -2926 1304 -2892 1338
rect -2994 1235 -2960 1269
rect -2926 1235 -2892 1269
rect -2092 3719 -1990 11233
rect -2092 3650 -2058 3684
rect -2024 3650 -1990 3684
rect -2092 3581 -2058 3615
rect -2024 3581 -1990 3615
rect -2092 3512 -2058 3546
rect -2024 3512 -1990 3546
rect -2092 3443 -2058 3477
rect -2024 3443 -1990 3477
rect -2092 3374 -2058 3408
rect -2024 3374 -1990 3408
rect -2092 3305 -2058 3339
rect -2024 3305 -1990 3339
rect -2092 3236 -2058 3270
rect -2024 3236 -1990 3270
rect -2092 3167 -2058 3201
rect -2024 3167 -1990 3201
rect -2092 3098 -2058 3132
rect -2024 3098 -1990 3132
rect -2092 3029 -2058 3063
rect -2024 3029 -1990 3063
rect -2092 2960 -2058 2994
rect -2024 2960 -1990 2994
rect -2092 2891 -2058 2925
rect -2024 2891 -1990 2925
rect -2092 2822 -2058 2856
rect -2024 2822 -1990 2856
rect -2092 2753 -2058 2787
rect -2024 2753 -1990 2787
rect -2092 2684 -2058 2718
rect -2024 2684 -1990 2718
rect -2092 2615 -2058 2649
rect -2024 2615 -1990 2649
rect -2092 2546 -2058 2580
rect -2024 2546 -1990 2580
rect -2092 2477 -2058 2511
rect -2024 2477 -1990 2511
rect -2092 2408 -2058 2442
rect -2024 2408 -1990 2442
rect -2092 2339 -2058 2373
rect -2024 2339 -1990 2373
rect -2092 2270 -2058 2304
rect -2024 2270 -1990 2304
rect -2092 2201 -2058 2235
rect -2024 2201 -1990 2235
rect -2092 2132 -2058 2166
rect -2024 2132 -1990 2166
rect -2092 2063 -2058 2097
rect -2024 2063 -1990 2097
rect -2092 1994 -2058 2028
rect -2024 1994 -1990 2028
rect -2092 1925 -2058 1959
rect -2024 1925 -1990 1959
rect -2092 1856 -2058 1890
rect -2024 1856 -1990 1890
rect -2092 1787 -2058 1821
rect -2024 1787 -1990 1821
rect -2092 1718 -2058 1752
rect -2024 1718 -1990 1752
rect -2092 1649 -2058 1683
rect -2024 1649 -1990 1683
rect -2092 1580 -2058 1614
rect -2024 1580 -1990 1614
rect -2092 1511 -2058 1545
rect -2024 1511 -1990 1545
rect -2092 1442 -2058 1476
rect -2024 1442 -1990 1476
rect -2092 1373 -2058 1407
rect -2024 1373 -1990 1407
rect -2092 1304 -2058 1338
rect -2024 1304 -1990 1338
rect -2092 1235 -2058 1269
rect -2024 1235 -1990 1269
rect -1190 3719 -1088 11233
rect -1190 3650 -1156 3684
rect -1122 3650 -1088 3684
rect -1190 3581 -1156 3615
rect -1122 3581 -1088 3615
rect -1190 3512 -1156 3546
rect -1122 3512 -1088 3546
rect -1190 3443 -1156 3477
rect -1122 3443 -1088 3477
rect -1190 3374 -1156 3408
rect -1122 3374 -1088 3408
rect -1190 3305 -1156 3339
rect -1122 3305 -1088 3339
rect -1190 3236 -1156 3270
rect -1122 3236 -1088 3270
rect -1190 3167 -1156 3201
rect -1122 3167 -1088 3201
rect -1190 3098 -1156 3132
rect -1122 3098 -1088 3132
rect -1190 3029 -1156 3063
rect -1122 3029 -1088 3063
rect -1190 2960 -1156 2994
rect -1122 2960 -1088 2994
rect -1190 2891 -1156 2925
rect -1122 2891 -1088 2925
rect -1190 2822 -1156 2856
rect -1122 2822 -1088 2856
rect -1190 2753 -1156 2787
rect -1122 2753 -1088 2787
rect -1190 2684 -1156 2718
rect -1122 2684 -1088 2718
rect -1190 2615 -1156 2649
rect -1122 2615 -1088 2649
rect -1190 2546 -1156 2580
rect -1122 2546 -1088 2580
rect -1190 2477 -1156 2511
rect -1122 2477 -1088 2511
rect -1190 2408 -1156 2442
rect -1122 2408 -1088 2442
rect -1190 2339 -1156 2373
rect -1122 2339 -1088 2373
rect -1190 2270 -1156 2304
rect -1122 2270 -1088 2304
rect -1190 2201 -1156 2235
rect -1122 2201 -1088 2235
rect -1190 2132 -1156 2166
rect -1122 2132 -1088 2166
rect -1190 2063 -1156 2097
rect -1122 2063 -1088 2097
rect -1190 1994 -1156 2028
rect -1122 1994 -1088 2028
rect -1190 1925 -1156 1959
rect -1122 1925 -1088 1959
rect -1190 1856 -1156 1890
rect -1122 1856 -1088 1890
rect -1190 1787 -1156 1821
rect -1122 1787 -1088 1821
rect -1190 1718 -1156 1752
rect -1122 1718 -1088 1752
rect -1190 1649 -1156 1683
rect -1122 1649 -1088 1683
rect -1190 1580 -1156 1614
rect -1122 1580 -1088 1614
rect -1190 1511 -1156 1545
rect -1122 1511 -1088 1545
rect -1190 1442 -1156 1476
rect -1122 1442 -1088 1476
rect -1190 1373 -1156 1407
rect -1122 1373 -1088 1407
rect -1190 1304 -1156 1338
rect -1122 1304 -1088 1338
rect -1190 1235 -1156 1269
rect -1122 1235 -1088 1269
rect -288 3719 -186 11233
rect -288 3650 -254 3684
rect -220 3650 -186 3684
rect -288 3581 -254 3615
rect -220 3581 -186 3615
rect -288 3512 -254 3546
rect -220 3512 -186 3546
rect -288 3443 -254 3477
rect -220 3443 -186 3477
rect -288 3374 -254 3408
rect -220 3374 -186 3408
rect -288 3305 -254 3339
rect -220 3305 -186 3339
rect -288 3236 -254 3270
rect -220 3236 -186 3270
rect -288 3167 -254 3201
rect -220 3167 -186 3201
rect -288 3098 -254 3132
rect -220 3098 -186 3132
rect -288 3029 -254 3063
rect -220 3029 -186 3063
rect -288 2960 -254 2994
rect -220 2960 -186 2994
rect -288 2891 -254 2925
rect -220 2891 -186 2925
rect -288 2822 -254 2856
rect -220 2822 -186 2856
rect -288 2753 -254 2787
rect -220 2753 -186 2787
rect -288 2684 -254 2718
rect -220 2684 -186 2718
rect -288 2615 -254 2649
rect -220 2615 -186 2649
rect -288 2546 -254 2580
rect -220 2546 -186 2580
rect -288 2477 -254 2511
rect -220 2477 -186 2511
rect -288 2408 -254 2442
rect -220 2408 -186 2442
rect -288 2339 -254 2373
rect -220 2339 -186 2373
rect -288 2270 -254 2304
rect -220 2270 -186 2304
rect -288 2201 -254 2235
rect -220 2201 -186 2235
rect -288 2132 -254 2166
rect -220 2132 -186 2166
rect -288 2063 -254 2097
rect -220 2063 -186 2097
rect -288 1994 -254 2028
rect -220 1994 -186 2028
rect -288 1925 -254 1959
rect -220 1925 -186 1959
rect -288 1856 -254 1890
rect -220 1856 -186 1890
rect -288 1787 -254 1821
rect -220 1787 -186 1821
rect -288 1718 -254 1752
rect -220 1718 -186 1752
rect -288 1649 -254 1683
rect -220 1649 -186 1683
rect -288 1580 -254 1614
rect -220 1580 -186 1614
rect -288 1511 -254 1545
rect -220 1511 -186 1545
rect -288 1442 -254 1476
rect -220 1442 -186 1476
rect -288 1373 -254 1407
rect -220 1373 -186 1407
rect -288 1304 -254 1338
rect -220 1304 -186 1338
rect -288 1235 -254 1269
rect -220 1235 -186 1269
rect 614 3719 716 11233
rect 614 3650 648 3684
rect 682 3650 716 3684
rect 614 3581 648 3615
rect 682 3581 716 3615
rect 614 3512 648 3546
rect 682 3512 716 3546
rect 614 3443 648 3477
rect 682 3443 716 3477
rect 614 3374 648 3408
rect 682 3374 716 3408
rect 614 3305 648 3339
rect 682 3305 716 3339
rect 614 3236 648 3270
rect 682 3236 716 3270
rect 614 3167 648 3201
rect 682 3167 716 3201
rect 614 3098 648 3132
rect 682 3098 716 3132
rect 614 3029 648 3063
rect 682 3029 716 3063
rect 614 2960 648 2994
rect 682 2960 716 2994
rect 614 2891 648 2925
rect 682 2891 716 2925
rect 614 2822 648 2856
rect 682 2822 716 2856
rect 614 2753 648 2787
rect 682 2753 716 2787
rect 614 2684 648 2718
rect 682 2684 716 2718
rect 614 2615 648 2649
rect 682 2615 716 2649
rect 614 2546 648 2580
rect 682 2546 716 2580
rect 614 2477 648 2511
rect 682 2477 716 2511
rect 614 2408 648 2442
rect 682 2408 716 2442
rect 614 2339 648 2373
rect 682 2339 716 2373
rect 614 2270 648 2304
rect 682 2270 716 2304
rect 614 2201 648 2235
rect 682 2201 716 2235
rect 614 2132 648 2166
rect 682 2132 716 2166
rect 614 2063 648 2097
rect 682 2063 716 2097
rect 614 1994 648 2028
rect 682 1994 716 2028
rect 614 1925 648 1959
rect 682 1925 716 1959
rect 614 1856 648 1890
rect 682 1856 716 1890
rect 614 1787 648 1821
rect 682 1787 716 1821
rect 614 1718 648 1752
rect 682 1718 716 1752
rect 614 1649 648 1683
rect 682 1649 716 1683
rect 614 1580 648 1614
rect 682 1580 716 1614
rect 614 1511 648 1545
rect 682 1511 716 1545
rect 614 1442 648 1476
rect 682 1442 716 1476
rect 614 1373 648 1407
rect 682 1373 716 1407
rect 614 1304 648 1338
rect 682 1304 716 1338
rect 614 1235 648 1269
rect 682 1235 716 1269
rect 1516 3719 1618 11233
rect 1516 3650 1550 3684
rect 1584 3650 1618 3684
rect 1516 3581 1550 3615
rect 1584 3581 1618 3615
rect 1516 3512 1550 3546
rect 1584 3512 1618 3546
rect 1516 3443 1550 3477
rect 1584 3443 1618 3477
rect 1516 3374 1550 3408
rect 1584 3374 1618 3408
rect 1516 3305 1550 3339
rect 1584 3305 1618 3339
rect 1516 3236 1550 3270
rect 1584 3236 1618 3270
rect 1516 3167 1550 3201
rect 1584 3167 1618 3201
rect 1516 3098 1550 3132
rect 1584 3098 1618 3132
rect 1516 3029 1550 3063
rect 1584 3029 1618 3063
rect 1516 2960 1550 2994
rect 1584 2960 1618 2994
rect 1516 2891 1550 2925
rect 1584 2891 1618 2925
rect 1516 2822 1550 2856
rect 1584 2822 1618 2856
rect 1516 2753 1550 2787
rect 1584 2753 1618 2787
rect 1516 2684 1550 2718
rect 1584 2684 1618 2718
rect 1516 2615 1550 2649
rect 1584 2615 1618 2649
rect 1516 2546 1550 2580
rect 1584 2546 1618 2580
rect 1516 2477 1550 2511
rect 1584 2477 1618 2511
rect 1516 2408 1550 2442
rect 1584 2408 1618 2442
rect 1516 2339 1550 2373
rect 1584 2339 1618 2373
rect 1516 2270 1550 2304
rect 1584 2270 1618 2304
rect 1516 2201 1550 2235
rect 1584 2201 1618 2235
rect 1516 2132 1550 2166
rect 1584 2132 1618 2166
rect 1516 2063 1550 2097
rect 1584 2063 1618 2097
rect 1516 1994 1550 2028
rect 1584 1994 1618 2028
rect 1516 1925 1550 1959
rect 1584 1925 1618 1959
rect 1516 1856 1550 1890
rect 1584 1856 1618 1890
rect 1516 1787 1550 1821
rect 1584 1787 1618 1821
rect 1516 1718 1550 1752
rect 1584 1718 1618 1752
rect 1516 1649 1550 1683
rect 1584 1649 1618 1683
rect 1516 1580 1550 1614
rect 1584 1580 1618 1614
rect 1516 1511 1550 1545
rect 1584 1511 1618 1545
rect 1516 1442 1550 1476
rect 1584 1442 1618 1476
rect 1516 1373 1550 1407
rect 1584 1373 1618 1407
rect 1516 1304 1550 1338
rect 1584 1304 1618 1338
rect 1516 1235 1550 1269
rect 1584 1235 1618 1269
rect 2418 3719 2520 11233
rect 2418 3650 2452 3684
rect 2486 3650 2520 3684
rect 2418 3581 2452 3615
rect 2486 3581 2520 3615
rect 2418 3512 2452 3546
rect 2486 3512 2520 3546
rect 2418 3443 2452 3477
rect 2486 3443 2520 3477
rect 2418 3374 2452 3408
rect 2486 3374 2520 3408
rect 2418 3305 2452 3339
rect 2486 3305 2520 3339
rect 2418 3236 2452 3270
rect 2486 3236 2520 3270
rect 2418 3167 2452 3201
rect 2486 3167 2520 3201
rect 2418 3098 2452 3132
rect 2486 3098 2520 3132
rect 2418 3029 2452 3063
rect 2486 3029 2520 3063
rect 2418 2960 2452 2994
rect 2486 2960 2520 2994
rect 2418 2891 2452 2925
rect 2486 2891 2520 2925
rect 2418 2822 2452 2856
rect 2486 2822 2520 2856
rect 2418 2753 2452 2787
rect 2486 2753 2520 2787
rect 2418 2684 2452 2718
rect 2486 2684 2520 2718
rect 2418 2615 2452 2649
rect 2486 2615 2520 2649
rect 2418 2546 2452 2580
rect 2486 2546 2520 2580
rect 2418 2477 2452 2511
rect 2486 2477 2520 2511
rect 2418 2408 2452 2442
rect 2486 2408 2520 2442
rect 2418 2339 2452 2373
rect 2486 2339 2520 2373
rect 2418 2270 2452 2304
rect 2486 2270 2520 2304
rect 2418 2201 2452 2235
rect 2486 2201 2520 2235
rect 2418 2132 2452 2166
rect 2486 2132 2520 2166
rect 2418 2063 2452 2097
rect 2486 2063 2520 2097
rect 2418 1994 2452 2028
rect 2486 1994 2520 2028
rect 2418 1925 2452 1959
rect 2486 1925 2520 1959
rect 2418 1856 2452 1890
rect 2486 1856 2520 1890
rect 2418 1787 2452 1821
rect 2486 1787 2520 1821
rect 2418 1718 2452 1752
rect 2486 1718 2520 1752
rect 2418 1649 2452 1683
rect 2486 1649 2520 1683
rect 2418 1580 2452 1614
rect 2486 1580 2520 1614
rect 2418 1511 2452 1545
rect 2486 1511 2520 1545
rect 2418 1442 2452 1476
rect 2486 1442 2520 1476
rect 2418 1373 2452 1407
rect 2486 1373 2520 1407
rect 2418 1304 2452 1338
rect 2486 1304 2520 1338
rect 2418 1235 2452 1269
rect 2486 1235 2520 1269
rect 3320 3719 3422 11233
rect 3320 3650 3354 3684
rect 3388 3650 3422 3684
rect 3320 3581 3354 3615
rect 3388 3581 3422 3615
rect 3320 3512 3354 3546
rect 3388 3512 3422 3546
rect 3320 3443 3354 3477
rect 3388 3443 3422 3477
rect 3320 3374 3354 3408
rect 3388 3374 3422 3408
rect 3320 3305 3354 3339
rect 3388 3305 3422 3339
rect 3320 3236 3354 3270
rect 3388 3236 3422 3270
rect 3320 3167 3354 3201
rect 3388 3167 3422 3201
rect 3320 3098 3354 3132
rect 3388 3098 3422 3132
rect 3320 3029 3354 3063
rect 3388 3029 3422 3063
rect 3320 2960 3354 2994
rect 3388 2960 3422 2994
rect 3320 2891 3354 2925
rect 3388 2891 3422 2925
rect 3320 2822 3354 2856
rect 3388 2822 3422 2856
rect 3320 2753 3354 2787
rect 3388 2753 3422 2787
rect 3320 2684 3354 2718
rect 3388 2684 3422 2718
rect 3320 2615 3354 2649
rect 3388 2615 3422 2649
rect 3320 2546 3354 2580
rect 3388 2546 3422 2580
rect 3320 2477 3354 2511
rect 3388 2477 3422 2511
rect 3320 2408 3354 2442
rect 3388 2408 3422 2442
rect 3320 2339 3354 2373
rect 3388 2339 3422 2373
rect 3320 2270 3354 2304
rect 3388 2270 3422 2304
rect 3320 2201 3354 2235
rect 3388 2201 3422 2235
rect 3320 2132 3354 2166
rect 3388 2132 3422 2166
rect 3320 2063 3354 2097
rect 3388 2063 3422 2097
rect 3320 1994 3354 2028
rect 3388 1994 3422 2028
rect 3320 1925 3354 1959
rect 3388 1925 3422 1959
rect 3320 1856 3354 1890
rect 3388 1856 3422 1890
rect 3320 1787 3354 1821
rect 3388 1787 3422 1821
rect 3320 1718 3354 1752
rect 3388 1718 3422 1752
rect 3320 1649 3354 1683
rect 3388 1649 3422 1683
rect 3320 1580 3354 1614
rect 3388 1580 3422 1614
rect 3320 1511 3354 1545
rect 3388 1511 3422 1545
rect 3320 1442 3354 1476
rect 3388 1442 3422 1476
rect 3320 1373 3354 1407
rect 3388 1373 3422 1407
rect 3320 1304 3354 1338
rect 3388 1304 3422 1338
rect 3320 1235 3354 1269
rect 3388 1235 3422 1269
rect 4222 3719 4324 11233
rect 4222 3650 4256 3684
rect 4290 3650 4324 3684
rect 4222 3581 4256 3615
rect 4290 3581 4324 3615
rect 4222 3512 4256 3546
rect 4290 3512 4324 3546
rect 4222 3443 4256 3477
rect 4290 3443 4324 3477
rect 4222 3374 4256 3408
rect 4290 3374 4324 3408
rect 4222 3305 4256 3339
rect 4290 3305 4324 3339
rect 4222 3236 4256 3270
rect 4290 3236 4324 3270
rect 4222 3167 4256 3201
rect 4290 3167 4324 3201
rect 4222 3098 4256 3132
rect 4290 3098 4324 3132
rect 4222 3029 4256 3063
rect 4290 3029 4324 3063
rect 4222 2960 4256 2994
rect 4290 2960 4324 2994
rect 4222 2891 4256 2925
rect 4290 2891 4324 2925
rect 4222 2822 4256 2856
rect 4290 2822 4324 2856
rect 4222 2753 4256 2787
rect 4290 2753 4324 2787
rect 4222 2684 4256 2718
rect 4290 2684 4324 2718
rect 4222 2615 4256 2649
rect 4290 2615 4324 2649
rect 4222 2546 4256 2580
rect 4290 2546 4324 2580
rect 4222 2477 4256 2511
rect 4290 2477 4324 2511
rect 4222 2408 4256 2442
rect 4290 2408 4324 2442
rect 4222 2339 4256 2373
rect 4290 2339 4324 2373
rect 4222 2270 4256 2304
rect 4290 2270 4324 2304
rect 4222 2201 4256 2235
rect 4290 2201 4324 2235
rect 4222 2132 4256 2166
rect 4290 2132 4324 2166
rect 4222 2063 4256 2097
rect 4290 2063 4324 2097
rect 4222 1994 4256 2028
rect 4290 1994 4324 2028
rect 4222 1925 4256 1959
rect 4290 1925 4324 1959
rect 4222 1856 4256 1890
rect 4290 1856 4324 1890
rect 4222 1787 4256 1821
rect 4290 1787 4324 1821
rect 4222 1718 4256 1752
rect 4290 1718 4324 1752
rect 4222 1649 4256 1683
rect 4290 1649 4324 1683
rect 4222 1580 4256 1614
rect 4290 1580 4324 1614
rect 4222 1511 4256 1545
rect 4290 1511 4324 1545
rect 4222 1442 4256 1476
rect 4290 1442 4324 1476
rect 4222 1373 4256 1407
rect 4290 1373 4324 1407
rect 4222 1304 4256 1338
rect 4290 1304 4324 1338
rect 4222 1235 4256 1269
rect 4290 1235 4324 1269
rect 5124 3719 5226 11233
rect 5124 3650 5158 3684
rect 5192 3650 5226 3684
rect 5124 3581 5158 3615
rect 5192 3581 5226 3615
rect 5124 3512 5158 3546
rect 5192 3512 5226 3546
rect 5124 3443 5158 3477
rect 5192 3443 5226 3477
rect 5124 3374 5158 3408
rect 5192 3374 5226 3408
rect 5124 3305 5158 3339
rect 5192 3305 5226 3339
rect 5124 3236 5158 3270
rect 5192 3236 5226 3270
rect 5124 3167 5158 3201
rect 5192 3167 5226 3201
rect 5124 3098 5158 3132
rect 5192 3098 5226 3132
rect 5124 3029 5158 3063
rect 5192 3029 5226 3063
rect 5124 2960 5158 2994
rect 5192 2960 5226 2994
rect 5124 2891 5158 2925
rect 5192 2891 5226 2925
rect 5124 2822 5158 2856
rect 5192 2822 5226 2856
rect 5124 2753 5158 2787
rect 5192 2753 5226 2787
rect 5124 2684 5158 2718
rect 5192 2684 5226 2718
rect 5124 2615 5158 2649
rect 5192 2615 5226 2649
rect 5124 2546 5158 2580
rect 5192 2546 5226 2580
rect 5124 2477 5158 2511
rect 5192 2477 5226 2511
rect 5124 2408 5158 2442
rect 5192 2408 5226 2442
rect 5124 2339 5158 2373
rect 5192 2339 5226 2373
rect 5124 2270 5158 2304
rect 5192 2270 5226 2304
rect 5124 2201 5158 2235
rect 5192 2201 5226 2235
rect 5124 2132 5158 2166
rect 5192 2132 5226 2166
rect 5124 2063 5158 2097
rect 5192 2063 5226 2097
rect 5124 1994 5158 2028
rect 5192 1994 5226 2028
rect 5124 1925 5158 1959
rect 5192 1925 5226 1959
rect 5124 1856 5158 1890
rect 5192 1856 5226 1890
rect 5124 1787 5158 1821
rect 5192 1787 5226 1821
rect 5124 1718 5158 1752
rect 5192 1718 5226 1752
rect 5124 1649 5158 1683
rect 5192 1649 5226 1683
rect 5124 1580 5158 1614
rect 5192 1580 5226 1614
rect 5124 1511 5158 1545
rect 5192 1511 5226 1545
rect 5124 1442 5158 1476
rect 5192 1442 5226 1476
rect 5124 1373 5158 1407
rect 5192 1373 5226 1407
rect 5124 1304 5158 1338
rect 5192 1304 5226 1338
rect 5124 1235 5158 1269
rect 5192 1235 5226 1269
rect 6026 3719 6128 11233
rect 6026 3650 6060 3684
rect 6094 3650 6128 3684
rect 6026 3581 6060 3615
rect 6094 3581 6128 3615
rect 6026 3512 6060 3546
rect 6094 3512 6128 3546
rect 6026 3443 6060 3477
rect 6094 3443 6128 3477
rect 6026 3374 6060 3408
rect 6094 3374 6128 3408
rect 6026 3305 6060 3339
rect 6094 3305 6128 3339
rect 6026 3236 6060 3270
rect 6094 3236 6128 3270
rect 6026 3167 6060 3201
rect 6094 3167 6128 3201
rect 6026 3098 6060 3132
rect 6094 3098 6128 3132
rect 6026 3029 6060 3063
rect 6094 3029 6128 3063
rect 6026 2960 6060 2994
rect 6094 2960 6128 2994
rect 6026 2891 6060 2925
rect 6094 2891 6128 2925
rect 6026 2822 6060 2856
rect 6094 2822 6128 2856
rect 6026 2753 6060 2787
rect 6094 2753 6128 2787
rect 6026 2684 6060 2718
rect 6094 2684 6128 2718
rect 6026 2615 6060 2649
rect 6094 2615 6128 2649
rect 6026 2546 6060 2580
rect 6094 2546 6128 2580
rect 6026 2477 6060 2511
rect 6094 2477 6128 2511
rect 6026 2408 6060 2442
rect 6094 2408 6128 2442
rect 6026 2339 6060 2373
rect 6094 2339 6128 2373
rect 6026 2270 6060 2304
rect 6094 2270 6128 2304
rect 6026 2201 6060 2235
rect 6094 2201 6128 2235
rect 6026 2132 6060 2166
rect 6094 2132 6128 2166
rect 6026 2063 6060 2097
rect 6094 2063 6128 2097
rect 6026 1994 6060 2028
rect 6094 1994 6128 2028
rect 6026 1925 6060 1959
rect 6094 1925 6128 1959
rect 6026 1856 6060 1890
rect 6094 1856 6128 1890
rect 6026 1787 6060 1821
rect 6094 1787 6128 1821
rect 6026 1718 6060 1752
rect 6094 1718 6128 1752
rect 6026 1649 6060 1683
rect 6094 1649 6128 1683
rect 6026 1580 6060 1614
rect 6094 1580 6128 1614
rect 6026 1511 6060 1545
rect 6094 1511 6128 1545
rect 6026 1442 6060 1476
rect 6094 1442 6128 1476
rect 6026 1373 6060 1407
rect 6094 1373 6128 1407
rect 6026 1304 6060 1338
rect 6094 1304 6128 1338
rect 6026 1235 6060 1269
rect 6094 1235 6128 1269
rect 6928 3719 7030 11233
rect 6928 3650 6962 3684
rect 6996 3650 7030 3684
rect 6928 3581 6962 3615
rect 6996 3581 7030 3615
rect 6928 3512 6962 3546
rect 6996 3512 7030 3546
rect 6928 3443 6962 3477
rect 6996 3443 7030 3477
rect 6928 3374 6962 3408
rect 6996 3374 7030 3408
rect 6928 3305 6962 3339
rect 6996 3305 7030 3339
rect 6928 3236 6962 3270
rect 6996 3236 7030 3270
rect 6928 3167 6962 3201
rect 6996 3167 7030 3201
rect 6928 3098 6962 3132
rect 6996 3098 7030 3132
rect 6928 3029 6962 3063
rect 6996 3029 7030 3063
rect 6928 2960 6962 2994
rect 6996 2960 7030 2994
rect 6928 2891 6962 2925
rect 6996 2891 7030 2925
rect 6928 2822 6962 2856
rect 6996 2822 7030 2856
rect 6928 2753 6962 2787
rect 6996 2753 7030 2787
rect 6928 2684 6962 2718
rect 6996 2684 7030 2718
rect 6928 2615 6962 2649
rect 6996 2615 7030 2649
rect 6928 2546 6962 2580
rect 6996 2546 7030 2580
rect 6928 2477 6962 2511
rect 6996 2477 7030 2511
rect 6928 2408 6962 2442
rect 6996 2408 7030 2442
rect 6928 2339 6962 2373
rect 6996 2339 7030 2373
rect 6928 2270 6962 2304
rect 6996 2270 7030 2304
rect 6928 2201 6962 2235
rect 6996 2201 7030 2235
rect 6928 2132 6962 2166
rect 6996 2132 7030 2166
rect 6928 2063 6962 2097
rect 6996 2063 7030 2097
rect 6928 1994 6962 2028
rect 6996 1994 7030 2028
rect 6928 1925 6962 1959
rect 6996 1925 7030 1959
rect 6928 1856 6962 1890
rect 6996 1856 7030 1890
rect 6928 1787 6962 1821
rect 6996 1787 7030 1821
rect 6928 1718 6962 1752
rect 6996 1718 7030 1752
rect 6928 1649 6962 1683
rect 6996 1649 7030 1683
rect 6928 1580 6962 1614
rect 6996 1580 7030 1614
rect 6928 1511 6962 1545
rect 6996 1511 7030 1545
rect 6928 1442 6962 1476
rect 6996 1442 7030 1476
rect 6928 1373 6962 1407
rect 6996 1373 7030 1407
rect 6928 1304 6962 1338
rect 6996 1304 7030 1338
rect 6928 1235 6962 1269
rect 6996 1235 7030 1269
rect 7830 3719 7932 11233
rect 7830 3650 7864 3684
rect 7898 3650 7932 3684
rect 7830 3581 7864 3615
rect 7898 3581 7932 3615
rect 7830 3512 7864 3546
rect 7898 3512 7932 3546
rect 7830 3443 7864 3477
rect 7898 3443 7932 3477
rect 7830 3374 7864 3408
rect 7898 3374 7932 3408
rect 7830 3305 7864 3339
rect 7898 3305 7932 3339
rect 7830 3236 7864 3270
rect 7898 3236 7932 3270
rect 7830 3167 7864 3201
rect 7898 3167 7932 3201
rect 7830 3098 7864 3132
rect 7898 3098 7932 3132
rect 7830 3029 7864 3063
rect 7898 3029 7932 3063
rect 7830 2960 7864 2994
rect 7898 2960 7932 2994
rect 7830 2891 7864 2925
rect 7898 2891 7932 2925
rect 7830 2822 7864 2856
rect 7898 2822 7932 2856
rect 7830 2753 7864 2787
rect 7898 2753 7932 2787
rect 7830 2684 7864 2718
rect 7898 2684 7932 2718
rect 7830 2615 7864 2649
rect 7898 2615 7932 2649
rect 7830 2546 7864 2580
rect 7898 2546 7932 2580
rect 7830 2477 7864 2511
rect 7898 2477 7932 2511
rect 7830 2408 7864 2442
rect 7898 2408 7932 2442
rect 7830 2339 7864 2373
rect 7898 2339 7932 2373
rect 7830 2270 7864 2304
rect 7898 2270 7932 2304
rect 7830 2201 7864 2235
rect 7898 2201 7932 2235
rect 7830 2132 7864 2166
rect 7898 2132 7932 2166
rect 7830 2063 7864 2097
rect 7898 2063 7932 2097
rect 7830 1994 7864 2028
rect 7898 1994 7932 2028
rect 7830 1925 7864 1959
rect 7898 1925 7932 1959
rect 7830 1856 7864 1890
rect 7898 1856 7932 1890
rect 7830 1787 7864 1821
rect 7898 1787 7932 1821
rect 7830 1718 7864 1752
rect 7898 1718 7932 1752
rect 7830 1649 7864 1683
rect 7898 1649 7932 1683
rect 7830 1580 7864 1614
rect 7898 1580 7932 1614
rect 7830 1511 7864 1545
rect 7898 1511 7932 1545
rect 7830 1442 7864 1476
rect 7898 1442 7932 1476
rect 7830 1373 7864 1407
rect 7898 1373 7932 1407
rect 7830 1304 7864 1338
rect 7898 1304 7932 1338
rect 7830 1235 7864 1269
rect 7898 1235 7932 1269
rect 8732 3719 8834 11233
rect 8732 3650 8766 3684
rect 8800 3650 8834 3684
rect 8732 3581 8766 3615
rect 8800 3581 8834 3615
rect 8732 3512 8766 3546
rect 8800 3512 8834 3546
rect 8732 3443 8766 3477
rect 8800 3443 8834 3477
rect 8732 3374 8766 3408
rect 8800 3374 8834 3408
rect 8732 3305 8766 3339
rect 8800 3305 8834 3339
rect 8732 3236 8766 3270
rect 8800 3236 8834 3270
rect 8732 3167 8766 3201
rect 8800 3167 8834 3201
rect 8732 3098 8766 3132
rect 8800 3098 8834 3132
rect 8732 3029 8766 3063
rect 8800 3029 8834 3063
rect 8732 2960 8766 2994
rect 8800 2960 8834 2994
rect 8732 2891 8766 2925
rect 8800 2891 8834 2925
rect 8732 2822 8766 2856
rect 8800 2822 8834 2856
rect 8732 2753 8766 2787
rect 8800 2753 8834 2787
rect 8732 2684 8766 2718
rect 8800 2684 8834 2718
rect 8732 2615 8766 2649
rect 8800 2615 8834 2649
rect 8732 2546 8766 2580
rect 8800 2546 8834 2580
rect 8732 2477 8766 2511
rect 8800 2477 8834 2511
rect 8732 2408 8766 2442
rect 8800 2408 8834 2442
rect 8732 2339 8766 2373
rect 8800 2339 8834 2373
rect 8732 2270 8766 2304
rect 8800 2270 8834 2304
rect 8732 2201 8766 2235
rect 8800 2201 8834 2235
rect 8732 2132 8766 2166
rect 8800 2132 8834 2166
rect 8732 2063 8766 2097
rect 8800 2063 8834 2097
rect 8732 1994 8766 2028
rect 8800 1994 8834 2028
rect 8732 1925 8766 1959
rect 8800 1925 8834 1959
rect 8732 1856 8766 1890
rect 8800 1856 8834 1890
rect 8732 1787 8766 1821
rect 8800 1787 8834 1821
rect 8732 1718 8766 1752
rect 8800 1718 8834 1752
rect 8732 1649 8766 1683
rect 8800 1649 8834 1683
rect 8732 1580 8766 1614
rect 8800 1580 8834 1614
rect 8732 1511 8766 1545
rect 8800 1511 8834 1545
rect 8732 1442 8766 1476
rect 8800 1442 8834 1476
rect 8732 1373 8766 1407
rect 8800 1373 8834 1407
rect 8732 1304 8766 1338
rect 8800 1304 8834 1338
rect 8732 1235 8766 1269
rect 8800 1235 8834 1269
rect 9634 3719 9736 11233
rect 9634 3650 9668 3684
rect 9702 3650 9736 3684
rect 9634 3581 9668 3615
rect 9702 3581 9736 3615
rect 9634 3512 9668 3546
rect 9702 3512 9736 3546
rect 9634 3443 9668 3477
rect 9702 3443 9736 3477
rect 9634 3374 9668 3408
rect 9702 3374 9736 3408
rect 9634 3305 9668 3339
rect 9702 3305 9736 3339
rect 9634 3236 9668 3270
rect 9702 3236 9736 3270
rect 9634 3167 9668 3201
rect 9702 3167 9736 3201
rect 9634 3098 9668 3132
rect 9702 3098 9736 3132
rect 9634 3029 9668 3063
rect 9702 3029 9736 3063
rect 9634 2960 9668 2994
rect 9702 2960 9736 2994
rect 9634 2891 9668 2925
rect 9702 2891 9736 2925
rect 9634 2822 9668 2856
rect 9702 2822 9736 2856
rect 9634 2753 9668 2787
rect 9702 2753 9736 2787
rect 9634 2684 9668 2718
rect 9702 2684 9736 2718
rect 9634 2615 9668 2649
rect 9702 2615 9736 2649
rect 9634 2546 9668 2580
rect 9702 2546 9736 2580
rect 9634 2477 9668 2511
rect 9702 2477 9736 2511
rect 9634 2408 9668 2442
rect 9702 2408 9736 2442
rect 9634 2339 9668 2373
rect 9702 2339 9736 2373
rect 9634 2270 9668 2304
rect 9702 2270 9736 2304
rect 9634 2201 9668 2235
rect 9702 2201 9736 2235
rect 9634 2132 9668 2166
rect 9702 2132 9736 2166
rect 9634 2063 9668 2097
rect 9702 2063 9736 2097
rect 9634 1994 9668 2028
rect 9702 1994 9736 2028
rect 9634 1925 9668 1959
rect 9702 1925 9736 1959
rect 9634 1856 9668 1890
rect 9702 1856 9736 1890
rect 9634 1787 9668 1821
rect 9702 1787 9736 1821
rect 9634 1718 9668 1752
rect 9702 1718 9736 1752
rect 9634 1649 9668 1683
rect 9702 1649 9736 1683
rect 9634 1580 9668 1614
rect 9702 1580 9736 1614
rect 9634 1511 9668 1545
rect 9702 1511 9736 1545
rect 9634 1442 9668 1476
rect 9702 1442 9736 1476
rect 9634 1373 9668 1407
rect 9702 1373 9736 1407
rect 9634 1304 9668 1338
rect 9702 1304 9736 1338
rect 9634 1235 9668 1269
rect 9702 1235 9736 1269
rect 10536 3719 10638 11233
rect 10536 3650 10570 3684
rect 10604 3650 10638 3684
rect 10536 3581 10570 3615
rect 10604 3581 10638 3615
rect 10536 3512 10570 3546
rect 10604 3512 10638 3546
rect 10536 3443 10570 3477
rect 10604 3443 10638 3477
rect 10536 3374 10570 3408
rect 10604 3374 10638 3408
rect 10536 3305 10570 3339
rect 10604 3305 10638 3339
rect 10536 3236 10570 3270
rect 10604 3236 10638 3270
rect 10536 3167 10570 3201
rect 10604 3167 10638 3201
rect 10536 3098 10570 3132
rect 10604 3098 10638 3132
rect 10536 3029 10570 3063
rect 10604 3029 10638 3063
rect 10536 2960 10570 2994
rect 10604 2960 10638 2994
rect 10536 2891 10570 2925
rect 10604 2891 10638 2925
rect 10536 2822 10570 2856
rect 10604 2822 10638 2856
rect 10536 2753 10570 2787
rect 10604 2753 10638 2787
rect 10536 2684 10570 2718
rect 10604 2684 10638 2718
rect 10536 2615 10570 2649
rect 10604 2615 10638 2649
rect 10536 2546 10570 2580
rect 10604 2546 10638 2580
rect 10536 2477 10570 2511
rect 10604 2477 10638 2511
rect 10536 2408 10570 2442
rect 10604 2408 10638 2442
rect 10536 2339 10570 2373
rect 10604 2339 10638 2373
rect 10536 2270 10570 2304
rect 10604 2270 10638 2304
rect 10536 2201 10570 2235
rect 10604 2201 10638 2235
rect 10536 2132 10570 2166
rect 10604 2132 10638 2166
rect 10536 2063 10570 2097
rect 10604 2063 10638 2097
rect 10536 1994 10570 2028
rect 10604 1994 10638 2028
rect 10536 1925 10570 1959
rect 10604 1925 10638 1959
rect 10536 1856 10570 1890
rect 10604 1856 10638 1890
rect 10536 1787 10570 1821
rect 10604 1787 10638 1821
rect 10536 1718 10570 1752
rect 10604 1718 10638 1752
rect 10536 1649 10570 1683
rect 10604 1649 10638 1683
rect 10536 1580 10570 1614
rect 10604 1580 10638 1614
rect 10536 1511 10570 1545
rect 10604 1511 10638 1545
rect 10536 1442 10570 1476
rect 10604 1442 10638 1476
rect 10536 1373 10570 1407
rect 10604 1373 10638 1407
rect 10536 1304 10570 1338
rect 10604 1304 10638 1338
rect 10536 1235 10570 1269
rect 10604 1235 10638 1269
rect 11438 3719 11540 11233
rect 11438 3650 11472 3684
rect 11506 3650 11540 3684
rect 11438 3581 11472 3615
rect 11506 3581 11540 3615
rect 11438 3512 11472 3546
rect 11506 3512 11540 3546
rect 11438 3443 11472 3477
rect 11506 3443 11540 3477
rect 11438 3374 11472 3408
rect 11506 3374 11540 3408
rect 11438 3305 11472 3339
rect 11506 3305 11540 3339
rect 11438 3236 11472 3270
rect 11506 3236 11540 3270
rect 11438 3167 11472 3201
rect 11506 3167 11540 3201
rect 11438 3098 11472 3132
rect 11506 3098 11540 3132
rect 11438 3029 11472 3063
rect 11506 3029 11540 3063
rect 11438 2960 11472 2994
rect 11506 2960 11540 2994
rect 11438 2891 11472 2925
rect 11506 2891 11540 2925
rect 11438 2822 11472 2856
rect 11506 2822 11540 2856
rect 11438 2753 11472 2787
rect 11506 2753 11540 2787
rect 11438 2684 11472 2718
rect 11506 2684 11540 2718
rect 11438 2615 11472 2649
rect 11506 2615 11540 2649
rect 11438 2546 11472 2580
rect 11506 2546 11540 2580
rect 11438 2477 11472 2511
rect 11506 2477 11540 2511
rect 11438 2408 11472 2442
rect 11506 2408 11540 2442
rect 11438 2339 11472 2373
rect 11506 2339 11540 2373
rect 11438 2270 11472 2304
rect 11506 2270 11540 2304
rect 11438 2201 11472 2235
rect 11506 2201 11540 2235
rect 11438 2132 11472 2166
rect 11506 2132 11540 2166
rect 11438 2063 11472 2097
rect 11506 2063 11540 2097
rect 11438 1994 11472 2028
rect 11506 1994 11540 2028
rect 11438 1925 11472 1959
rect 11506 1925 11540 1959
rect 11438 1856 11472 1890
rect 11506 1856 11540 1890
rect 11438 1787 11472 1821
rect 11506 1787 11540 1821
rect 11438 1718 11472 1752
rect 11506 1718 11540 1752
rect 11438 1649 11472 1683
rect 11506 1649 11540 1683
rect 11438 1580 11472 1614
rect 11506 1580 11540 1614
rect 11438 1511 11472 1545
rect 11506 1511 11540 1545
rect 11438 1442 11472 1476
rect 11506 1442 11540 1476
rect 11438 1373 11472 1407
rect 11506 1373 11540 1407
rect 11438 1304 11472 1338
rect 11506 1304 11540 1338
rect 11438 1235 11472 1269
rect 11506 1235 11540 1269
rect 12340 3719 12442 11233
rect 12340 3650 12374 3684
rect 12408 3650 12442 3684
rect 12340 3581 12374 3615
rect 12408 3581 12442 3615
rect 12340 3512 12374 3546
rect 12408 3512 12442 3546
rect 12340 3443 12374 3477
rect 12408 3443 12442 3477
rect 12340 3374 12374 3408
rect 12408 3374 12442 3408
rect 12340 3305 12374 3339
rect 12408 3305 12442 3339
rect 12340 3236 12374 3270
rect 12408 3236 12442 3270
rect 12340 3167 12374 3201
rect 12408 3167 12442 3201
rect 12340 3098 12374 3132
rect 12408 3098 12442 3132
rect 12340 3029 12374 3063
rect 12408 3029 12442 3063
rect 12340 2960 12374 2994
rect 12408 2960 12442 2994
rect 12340 2891 12374 2925
rect 12408 2891 12442 2925
rect 12340 2822 12374 2856
rect 12408 2822 12442 2856
rect 12340 2753 12374 2787
rect 12408 2753 12442 2787
rect 12340 2684 12374 2718
rect 12408 2684 12442 2718
rect 12340 2615 12374 2649
rect 12408 2615 12442 2649
rect 12340 2546 12374 2580
rect 12408 2546 12442 2580
rect 12340 2477 12374 2511
rect 12408 2477 12442 2511
rect 12340 2408 12374 2442
rect 12408 2408 12442 2442
rect 12340 2339 12374 2373
rect 12408 2339 12442 2373
rect 12340 2270 12374 2304
rect 12408 2270 12442 2304
rect 12340 2201 12374 2235
rect 12408 2201 12442 2235
rect 12340 2132 12374 2166
rect 12408 2132 12442 2166
rect 12340 2063 12374 2097
rect 12408 2063 12442 2097
rect 12340 1994 12374 2028
rect 12408 1994 12442 2028
rect 12340 1925 12374 1959
rect 12408 1925 12442 1959
rect 12340 1856 12374 1890
rect 12408 1856 12442 1890
rect 12340 1787 12374 1821
rect 12408 1787 12442 1821
rect 12340 1718 12374 1752
rect 12408 1718 12442 1752
rect 12340 1649 12374 1683
rect 12408 1649 12442 1683
rect 12340 1580 12374 1614
rect 12408 1580 12442 1614
rect 12340 1511 12374 1545
rect 12408 1511 12442 1545
rect 12340 1442 12374 1476
rect 12408 1442 12442 1476
rect 12340 1373 12374 1407
rect 12408 1373 12442 1407
rect 12340 1304 12374 1338
rect 12408 1304 12442 1338
rect 12340 1235 12374 1269
rect 12408 1235 12442 1269
rect 13242 3719 13344 11233
rect 13242 3650 13276 3684
rect 13310 3650 13344 3684
rect 13242 3581 13276 3615
rect 13310 3581 13344 3615
rect 13242 3512 13276 3546
rect 13310 3512 13344 3546
rect 13242 3443 13276 3477
rect 13310 3443 13344 3477
rect 13242 3374 13276 3408
rect 13310 3374 13344 3408
rect 13242 3305 13276 3339
rect 13310 3305 13344 3339
rect 13242 3236 13276 3270
rect 13310 3236 13344 3270
rect 13242 3167 13276 3201
rect 13310 3167 13344 3201
rect 13242 3098 13276 3132
rect 13310 3098 13344 3132
rect 13242 3029 13276 3063
rect 13310 3029 13344 3063
rect 13242 2960 13276 2994
rect 13310 2960 13344 2994
rect 13242 2891 13276 2925
rect 13310 2891 13344 2925
rect 13242 2822 13276 2856
rect 13310 2822 13344 2856
rect 13242 2753 13276 2787
rect 13310 2753 13344 2787
rect 13242 2684 13276 2718
rect 13310 2684 13344 2718
rect 13242 2615 13276 2649
rect 13310 2615 13344 2649
rect 13242 2546 13276 2580
rect 13310 2546 13344 2580
rect 13242 2477 13276 2511
rect 13310 2477 13344 2511
rect 13242 2408 13276 2442
rect 13310 2408 13344 2442
rect 13242 2339 13276 2373
rect 13310 2339 13344 2373
rect 13242 2270 13276 2304
rect 13310 2270 13344 2304
rect 13242 2201 13276 2235
rect 13310 2201 13344 2235
rect 13242 2132 13276 2166
rect 13310 2132 13344 2166
rect 13242 2063 13276 2097
rect 13310 2063 13344 2097
rect 13242 1994 13276 2028
rect 13310 1994 13344 2028
rect 13242 1925 13276 1959
rect 13310 1925 13344 1959
rect 13242 1856 13276 1890
rect 13310 1856 13344 1890
rect 13242 1787 13276 1821
rect 13310 1787 13344 1821
rect 13242 1718 13276 1752
rect 13310 1718 13344 1752
rect 13242 1649 13276 1683
rect 13310 1649 13344 1683
rect 13242 1580 13276 1614
rect 13310 1580 13344 1614
rect 13242 1511 13276 1545
rect 13310 1511 13344 1545
rect 13242 1442 13276 1476
rect 13310 1442 13344 1476
rect 13242 1373 13276 1407
rect 13310 1373 13344 1407
rect 13242 1304 13276 1338
rect 13310 1304 13344 1338
rect 13242 1235 13276 1269
rect 13310 1235 13344 1269
rect 14144 3719 14246 11233
rect 14144 3650 14178 3684
rect 14212 3650 14246 3684
rect 14144 3581 14178 3615
rect 14212 3581 14246 3615
rect 14144 3512 14178 3546
rect 14212 3512 14246 3546
rect 14144 3443 14178 3477
rect 14212 3443 14246 3477
rect 14144 3374 14178 3408
rect 14212 3374 14246 3408
rect 14144 3305 14178 3339
rect 14212 3305 14246 3339
rect 14144 3236 14178 3270
rect 14212 3236 14246 3270
rect 14144 3167 14178 3201
rect 14212 3167 14246 3201
rect 14144 3098 14178 3132
rect 14212 3098 14246 3132
rect 14144 3029 14178 3063
rect 14212 3029 14246 3063
rect 14144 2960 14178 2994
rect 14212 2960 14246 2994
rect 14144 2891 14178 2925
rect 14212 2891 14246 2925
rect 14144 2822 14178 2856
rect 14212 2822 14246 2856
rect 14144 2753 14178 2787
rect 14212 2753 14246 2787
rect 14144 2684 14178 2718
rect 14212 2684 14246 2718
rect 14144 2615 14178 2649
rect 14212 2615 14246 2649
rect 14144 2546 14178 2580
rect 14212 2546 14246 2580
rect 14144 2477 14178 2511
rect 14212 2477 14246 2511
rect 14144 2408 14178 2442
rect 14212 2408 14246 2442
rect 14144 2339 14178 2373
rect 14212 2339 14246 2373
rect 14144 2270 14178 2304
rect 14212 2270 14246 2304
rect 14144 2201 14178 2235
rect 14212 2201 14246 2235
rect 14144 2132 14178 2166
rect 14212 2132 14246 2166
rect 14144 2063 14178 2097
rect 14212 2063 14246 2097
rect 14144 1994 14178 2028
rect 14212 1994 14246 2028
rect 14144 1925 14178 1959
rect 14212 1925 14246 1959
rect 14144 1856 14178 1890
rect 14212 1856 14246 1890
rect 14144 1787 14178 1821
rect 14212 1787 14246 1821
rect 14144 1718 14178 1752
rect 14212 1718 14246 1752
rect 14144 1649 14178 1683
rect 14212 1649 14246 1683
rect 14144 1580 14178 1614
rect 14212 1580 14246 1614
rect 14144 1511 14178 1545
rect 14212 1511 14246 1545
rect 14144 1442 14178 1476
rect 14212 1442 14246 1476
rect 14144 1373 14178 1407
rect 14212 1373 14246 1407
rect 14144 1304 14178 1338
rect 14212 1304 14246 1338
rect 14144 1235 14178 1269
rect 14212 1235 14246 1269
<< mvpsubdiff >>
rect -4436 11796 -4368 11830
rect -4334 11796 -4299 11830
rect -4265 11796 -4227 11830
rect -4193 11796 -4158 11830
rect -4124 11796 -4089 11830
rect -4055 11796 -4020 11830
rect -3986 11796 -3933 11830
rect -3899 11796 -3864 11830
rect -3830 11796 -3795 11830
rect -3761 11796 -3726 11830
rect -3692 11796 -3657 11830
rect -3623 11796 -3588 11830
rect -3554 11796 -3519 11830
rect -3485 11796 -3450 11830
rect -3416 11796 -3381 11830
rect -3347 11796 -3312 11830
rect -3278 11796 -3243 11830
rect -3209 11796 -3174 11830
rect -3140 11796 -3105 11830
rect -3071 11796 -3036 11830
rect -3002 11796 -2967 11830
rect -2933 11796 -2898 11830
rect -2864 11796 -2829 11830
rect -2795 11796 -2760 11830
rect -2726 11796 -2691 11830
rect -2657 11796 -2622 11830
rect -2588 11796 -2553 11830
rect -2519 11796 -2484 11830
rect -2450 11796 -2415 11830
rect -2381 11796 -2346 11830
rect -2312 11796 -2277 11830
rect -2243 11796 -2208 11830
rect -2174 11796 -2139 11830
rect -2105 11796 -2070 11830
rect -2036 11796 -2001 11830
rect -1967 11796 -1932 11830
rect -1898 11796 -1863 11830
rect -1829 11796 -1794 11830
rect -4436 11762 -1794 11796
rect -4436 11728 -4368 11762
rect -4334 11728 -4299 11762
rect -4265 11728 -4227 11762
rect -4193 11728 -4158 11762
rect -4124 11728 -4089 11762
rect -4055 11728 -4020 11762
rect -3986 11728 -3933 11762
rect -3899 11728 -3864 11762
rect -3830 11728 -3795 11762
rect -3761 11728 -3726 11762
rect -3692 11728 -3657 11762
rect -3623 11728 -3588 11762
rect -3554 11728 -3519 11762
rect -3485 11728 -3450 11762
rect -3416 11728 -3381 11762
rect -3347 11728 -3312 11762
rect -3278 11728 -3243 11762
rect -3209 11728 -3174 11762
rect -3140 11728 -3105 11762
rect -3071 11728 -3036 11762
rect -3002 11728 -2967 11762
rect -2933 11728 -2898 11762
rect -2864 11728 -2829 11762
rect -2795 11728 -2760 11762
rect -2726 11728 -2691 11762
rect -2657 11728 -2622 11762
rect -2588 11728 -2553 11762
rect -2519 11728 -2484 11762
rect -2450 11728 -2415 11762
rect -2381 11728 -2346 11762
rect -2312 11728 -2277 11762
rect -2243 11728 -2208 11762
rect -2174 11728 -2139 11762
rect -2105 11728 -2070 11762
rect -2036 11728 -2001 11762
rect -1967 11728 -1932 11762
rect -1898 11728 -1863 11762
rect -1829 11728 -1794 11762
rect -4436 11694 -1794 11728
rect -4436 11660 -4368 11694
rect -4334 11660 -4299 11694
rect -4265 11660 -4227 11694
rect -4193 11660 -4158 11694
rect -4124 11660 -4089 11694
rect -4055 11660 -4020 11694
rect -3986 11660 -3933 11694
rect -3899 11660 -3864 11694
rect -3830 11660 -3795 11694
rect -3761 11660 -3726 11694
rect -3692 11660 -3657 11694
rect -3623 11660 -3588 11694
rect -3554 11660 -3519 11694
rect -3485 11660 -3450 11694
rect -3416 11660 -3381 11694
rect -3347 11660 -3312 11694
rect -3278 11660 -3243 11694
rect -3209 11660 -3174 11694
rect -3140 11660 -3105 11694
rect -3071 11660 -3036 11694
rect -3002 11660 -2967 11694
rect -2933 11660 -2898 11694
rect -2864 11660 -2829 11694
rect -2795 11660 -2760 11694
rect -2726 11660 -2691 11694
rect -2657 11660 -2622 11694
rect -2588 11660 -2553 11694
rect -2519 11660 -2484 11694
rect -2450 11660 -2415 11694
rect -2381 11660 -2346 11694
rect -2312 11660 -2277 11694
rect -2243 11660 -2208 11694
rect -2174 11660 -2139 11694
rect -2105 11660 -2070 11694
rect -2036 11660 -2001 11694
rect -1967 11660 -1932 11694
rect -1898 11660 -1863 11694
rect -1829 11660 -1794 11694
rect 824 11796 859 11830
rect 893 11796 928 11830
rect 962 11796 997 11830
rect 1031 11796 1066 11830
rect 1100 11796 1135 11830
rect 1169 11796 1204 11830
rect 1238 11796 1273 11830
rect 1307 11796 1342 11830
rect 1376 11796 1411 11830
rect 1445 11796 1480 11830
rect 1514 11796 1549 11830
rect 1583 11796 1618 11830
rect 1652 11796 1687 11830
rect 1721 11796 1756 11830
rect 1790 11796 1825 11830
rect 1859 11796 1894 11830
rect 1928 11796 1963 11830
rect 1997 11796 2032 11830
rect 2066 11796 2101 11830
rect 2135 11796 2170 11830
rect 2204 11796 2239 11830
rect 2273 11796 2308 11830
rect 824 11762 2308 11796
rect 824 11728 859 11762
rect 893 11728 928 11762
rect 962 11728 997 11762
rect 1031 11728 1066 11762
rect 1100 11728 1135 11762
rect 1169 11728 1204 11762
rect 1238 11728 1273 11762
rect 1307 11728 1342 11762
rect 1376 11728 1411 11762
rect 1445 11728 1480 11762
rect 1514 11728 1549 11762
rect 1583 11728 1618 11762
rect 1652 11728 1687 11762
rect 1721 11728 1756 11762
rect 1790 11728 1825 11762
rect 1859 11728 1894 11762
rect 1928 11728 1963 11762
rect 1997 11728 2032 11762
rect 2066 11728 2101 11762
rect 2135 11728 2170 11762
rect 2204 11728 2239 11762
rect 2273 11728 2308 11762
rect 824 11694 2308 11728
rect 824 11660 859 11694
rect 893 11660 928 11694
rect 962 11660 997 11694
rect 1031 11660 1066 11694
rect 1100 11660 1135 11694
rect 1169 11660 1204 11694
rect 1238 11660 1273 11694
rect 1307 11660 1342 11694
rect 1376 11660 1411 11694
rect 1445 11660 1480 11694
rect 1514 11660 1549 11694
rect 1583 11660 1618 11694
rect 1652 11660 1687 11694
rect 1721 11660 1756 11694
rect 1790 11660 1825 11694
rect 1859 11660 1894 11694
rect 1928 11660 1963 11694
rect 1997 11660 2032 11694
rect 2066 11660 2101 11694
rect 2135 11660 2170 11694
rect 2204 11660 2239 11694
rect 2273 11660 2308 11694
rect 14718 11660 14786 11830
rect -4436 11617 -4266 11660
rect -4402 11583 -4368 11617
rect -4334 11583 -4300 11617
rect -4436 11502 -4266 11583
rect 14616 11617 14786 11660
rect 14650 11583 14684 11617
rect 14718 11583 14752 11617
rect 14616 11502 14786 11583
rect -4436 1777 -4266 1812
rect -4402 1743 -4368 1777
rect -4334 1743 -4300 1777
rect -4436 1708 -4266 1743
rect -4402 1674 -4368 1708
rect -4334 1674 -4300 1708
rect -4436 1639 -4266 1674
rect -4402 1605 -4368 1639
rect -4334 1605 -4300 1639
rect -4436 1570 -4266 1605
rect -4402 1536 -4368 1570
rect -4334 1536 -4300 1570
rect -4436 1501 -4266 1536
rect -4402 1467 -4368 1501
rect -4334 1467 -4300 1501
rect -4436 1432 -4266 1467
rect -4402 1398 -4368 1432
rect -4334 1398 -4300 1432
rect -4436 1363 -4266 1398
rect -4402 1329 -4368 1363
rect -4334 1329 -4300 1363
rect -4436 1294 -4266 1329
rect -4402 1260 -4368 1294
rect -4334 1260 -4300 1294
rect -4436 1225 -4266 1260
rect -4402 1191 -4368 1225
rect -4334 1191 -4300 1225
rect -4436 1156 -4266 1191
rect -4402 1122 -4368 1156
rect -4334 1122 -4300 1156
rect 14616 1777 14786 1812
rect 14650 1743 14684 1777
rect 14718 1743 14752 1777
rect 14616 1708 14786 1743
rect 14650 1674 14684 1708
rect 14718 1674 14752 1708
rect 14616 1639 14786 1674
rect 14650 1605 14684 1639
rect 14718 1605 14752 1639
rect 14616 1570 14786 1605
rect 14650 1536 14684 1570
rect 14718 1536 14752 1570
rect 14616 1501 14786 1536
rect 14650 1467 14684 1501
rect 14718 1467 14752 1501
rect 14616 1432 14786 1467
rect 14650 1398 14684 1432
rect 14718 1398 14752 1432
rect 14616 1363 14786 1398
rect 14650 1329 14684 1363
rect 14718 1329 14752 1363
rect 14616 1294 14786 1329
rect 14650 1260 14684 1294
rect 14718 1260 14752 1294
rect 14616 1225 14786 1260
rect 14650 1191 14684 1225
rect 14718 1191 14752 1225
rect 14616 1156 14786 1191
rect -4436 1087 -4266 1122
rect -4402 1053 -4368 1087
rect -4334 1053 -4300 1087
rect -4436 1018 -4266 1053
rect -4402 984 -4368 1018
rect -4334 984 -4300 1018
rect 14650 1122 14684 1156
rect 14718 1122 14752 1156
rect 14616 1087 14786 1122
rect 14650 1053 14684 1087
rect 14718 1053 14752 1087
rect 14616 1018 14786 1053
rect -4436 949 -4266 984
rect -4402 915 -4368 949
rect -4334 915 -4300 949
rect -4436 880 -4266 915
rect -4402 846 -4368 880
rect -4334 846 -4300 880
rect -4436 811 -4266 846
rect -4402 777 -4368 811
rect -4334 777 -4300 811
rect -4436 742 -4266 777
rect -4402 708 -4368 742
rect -4334 708 -4300 742
rect -4436 640 -4266 708
rect 14650 984 14684 1018
rect 14718 984 14752 1018
rect 14616 949 14786 984
rect 14650 915 14684 949
rect 14718 915 14752 949
rect 14616 880 14786 915
rect 14650 846 14684 880
rect 14718 846 14752 880
rect 14616 811 14786 846
rect 14650 777 14684 811
rect 14718 777 14752 811
rect 14616 742 14786 777
rect 14650 708 14684 742
rect 14718 708 14752 742
rect 14616 640 14786 708
rect -4436 606 -4368 640
rect -4334 606 -4299 640
rect -4265 606 -4230 640
rect -4196 606 -4158 640
rect -4124 606 -4089 640
rect -4055 606 -4020 640
rect -3986 606 -3933 640
rect -3899 606 -3864 640
rect -3830 606 -3795 640
rect -3761 606 -3726 640
rect -3692 606 -3657 640
rect -3623 606 -3588 640
rect -3554 606 -3519 640
rect -3485 606 -3450 640
rect -3416 606 -3381 640
rect -3347 606 -3312 640
rect -3278 606 -3243 640
rect -3209 606 -3174 640
rect -3140 606 -3105 640
rect -3071 606 -3036 640
rect -3002 606 -2967 640
rect -2933 606 -2898 640
rect -2864 606 -2829 640
rect -2795 606 -2760 640
rect -2726 606 -2691 640
rect -2657 606 -2622 640
rect -2588 606 -2553 640
rect -2519 606 -2484 640
rect -2450 606 -2415 640
rect -2381 606 -2346 640
rect -2312 606 -2277 640
rect -2243 606 -2208 640
rect -2174 606 -2139 640
rect -2105 606 -2070 640
rect -2036 606 -2001 640
rect -1967 606 -1932 640
rect -1898 606 -1863 640
rect -1829 606 -1794 640
rect -4436 572 -1794 606
rect -4436 538 -4368 572
rect -4334 538 -4299 572
rect -4265 538 -4230 572
rect -4196 538 -4158 572
rect -4124 538 -4089 572
rect -4055 538 -4020 572
rect -3986 538 -3933 572
rect -3899 538 -3864 572
rect -3830 538 -3795 572
rect -3761 538 -3726 572
rect -3692 538 -3657 572
rect -3623 538 -3588 572
rect -3554 538 -3519 572
rect -3485 538 -3450 572
rect -3416 538 -3381 572
rect -3347 538 -3312 572
rect -3278 538 -3243 572
rect -3209 538 -3174 572
rect -3140 538 -3105 572
rect -3071 538 -3036 572
rect -3002 538 -2967 572
rect -2933 538 -2898 572
rect -2864 538 -2829 572
rect -2795 538 -2760 572
rect -2726 538 -2691 572
rect -2657 538 -2622 572
rect -2588 538 -2553 572
rect -2519 538 -2484 572
rect -2450 538 -2415 572
rect -2381 538 -2346 572
rect -2312 538 -2277 572
rect -2243 538 -2208 572
rect -2174 538 -2139 572
rect -2105 538 -2070 572
rect -2036 538 -2001 572
rect -1967 538 -1932 572
rect -1898 538 -1863 572
rect -1829 538 -1794 572
rect -4436 504 -1794 538
rect -4436 470 -4368 504
rect -4334 470 -4299 504
rect -4265 470 -4230 504
rect -4196 470 -4158 504
rect -4124 470 -4089 504
rect -4055 470 -4020 504
rect -3986 470 -3933 504
rect -3899 470 -3864 504
rect -3830 470 -3795 504
rect -3761 470 -3726 504
rect -3692 470 -3657 504
rect -3623 470 -3588 504
rect -3554 470 -3519 504
rect -3485 470 -3450 504
rect -3416 470 -3381 504
rect -3347 470 -3312 504
rect -3278 470 -3243 504
rect -3209 470 -3174 504
rect -3140 470 -3105 504
rect -3071 470 -3036 504
rect -3002 470 -2967 504
rect -2933 470 -2898 504
rect -2864 470 -2829 504
rect -2795 470 -2760 504
rect -2726 470 -2691 504
rect -2657 470 -2622 504
rect -2588 470 -2553 504
rect -2519 470 -2484 504
rect -2450 470 -2415 504
rect -2381 470 -2346 504
rect -2312 470 -2277 504
rect -2243 470 -2208 504
rect -2174 470 -2139 504
rect -2105 470 -2070 504
rect -2036 470 -2001 504
rect -1967 470 -1932 504
rect -1898 470 -1863 504
rect -1829 470 -1794 504
rect 824 606 859 640
rect 893 606 928 640
rect 962 606 997 640
rect 1031 606 1066 640
rect 1100 606 1135 640
rect 1169 606 1204 640
rect 1238 606 1273 640
rect 1307 606 1342 640
rect 1376 606 1411 640
rect 1445 606 1480 640
rect 1514 606 1549 640
rect 1583 606 1618 640
rect 1652 606 1687 640
rect 1721 606 1756 640
rect 1790 606 1825 640
rect 1859 606 1894 640
rect 1928 606 1963 640
rect 1997 606 2032 640
rect 2066 606 2101 640
rect 2135 606 2170 640
rect 2204 606 2239 640
rect 2273 606 2308 640
rect 824 572 2308 606
rect 824 538 859 572
rect 893 538 928 572
rect 962 538 997 572
rect 1031 538 1066 572
rect 1100 538 1135 572
rect 1169 538 1204 572
rect 1238 538 1273 572
rect 1307 538 1342 572
rect 1376 538 1411 572
rect 1445 538 1480 572
rect 1514 538 1549 572
rect 1583 538 1618 572
rect 1652 538 1687 572
rect 1721 538 1756 572
rect 1790 538 1825 572
rect 1859 538 1894 572
rect 1928 538 1963 572
rect 1997 538 2032 572
rect 2066 538 2101 572
rect 2135 538 2170 572
rect 2204 538 2239 572
rect 2273 538 2308 572
rect 824 504 2308 538
rect 824 470 859 504
rect 893 470 928 504
rect 962 470 997 504
rect 1031 470 1066 504
rect 1100 470 1135 504
rect 1169 470 1204 504
rect 1238 470 1273 504
rect 1307 470 1342 504
rect 1376 470 1411 504
rect 1445 470 1480 504
rect 1514 470 1549 504
rect 1583 470 1618 504
rect 1652 470 1687 504
rect 1721 470 1756 504
rect 1790 470 1825 504
rect 1859 470 1894 504
rect 1928 470 1963 504
rect 1997 470 2032 504
rect 2066 470 2101 504
rect 2135 470 2170 504
rect 2204 470 2239 504
rect 2273 470 2308 504
rect 14718 470 14786 640
<< mvnsubdiff >>
rect -4920 12966 -4852 13000
rect -4818 12966 -4783 13000
rect -4749 12966 -4703 13000
rect -4669 12966 -4634 13000
rect -4600 12966 -4565 13000
rect -4531 12966 -4496 13000
rect -4462 12966 -4427 13000
rect -4393 12966 -4358 13000
rect -4324 12966 -4289 13000
rect -4255 12966 -4220 13000
rect -4186 12966 -4151 13000
rect -4117 12966 -4082 13000
rect -4048 12966 -4013 13000
rect -3979 12966 -3944 13000
rect -3910 12966 -3875 13000
rect -3841 12966 -3806 13000
rect -3772 12966 -3737 13000
rect -3703 12966 -3668 13000
rect -3634 12966 -3599 13000
rect -3565 12966 -3530 13000
rect -3496 12966 -3461 13000
rect -3427 12966 -3392 13000
rect -3358 12966 -3323 13000
rect -3289 12966 -3254 13000
rect -3220 12966 -3185 13000
rect -3151 12966 -3116 13000
rect -3082 12966 -3029 13000
rect -2995 12966 -2960 13000
rect -2926 12966 -2891 13000
rect -2857 12966 -2822 13000
rect -4920 12932 -2822 12966
rect -4920 12898 -4852 12932
rect -4818 12898 -4783 12932
rect -4749 12898 -4703 12932
rect -4669 12898 -4634 12932
rect -4600 12898 -4565 12932
rect -4531 12898 -4496 12932
rect -4462 12898 -4427 12932
rect -4393 12898 -4358 12932
rect -4324 12898 -4289 12932
rect -4255 12898 -4220 12932
rect -4186 12898 -4151 12932
rect -4117 12898 -4082 12932
rect -4048 12898 -4013 12932
rect -3979 12898 -3944 12932
rect -3910 12898 -3875 12932
rect -3841 12898 -3806 12932
rect -3772 12898 -3737 12932
rect -3703 12898 -3668 12932
rect -3634 12898 -3599 12932
rect -3565 12898 -3530 12932
rect -3496 12898 -3461 12932
rect -3427 12898 -3392 12932
rect -3358 12898 -3323 12932
rect -3289 12898 -3254 12932
rect -3220 12898 -3185 12932
rect -3151 12898 -3116 12932
rect -3082 12898 -3029 12932
rect -2995 12898 -2960 12932
rect -2926 12898 -2891 12932
rect -2857 12898 -2822 12932
rect -4920 12864 -2822 12898
rect -4920 12830 -4852 12864
rect -4818 12830 -4783 12864
rect -4749 12830 -4703 12864
rect -4669 12830 -4634 12864
rect -4600 12830 -4565 12864
rect -4531 12830 -4496 12864
rect -4462 12830 -4427 12864
rect -4393 12830 -4358 12864
rect -4324 12830 -4289 12864
rect -4255 12830 -4220 12864
rect -4186 12830 -4151 12864
rect -4117 12830 -4082 12864
rect -4048 12830 -4013 12864
rect -3979 12830 -3944 12864
rect -3910 12830 -3875 12864
rect -3841 12830 -3806 12864
rect -3772 12830 -3737 12864
rect -3703 12830 -3668 12864
rect -3634 12830 -3599 12864
rect -3565 12830 -3530 12864
rect -3496 12830 -3461 12864
rect -3427 12830 -3392 12864
rect -3358 12830 -3323 12864
rect -3289 12830 -3254 12864
rect -3220 12830 -3185 12864
rect -3151 12830 -3116 12864
rect -3082 12830 -3029 12864
rect -2995 12830 -2960 12864
rect -2926 12830 -2891 12864
rect -2857 12830 -2822 12864
rect 340 12966 375 13000
rect 409 12966 444 13000
rect 478 12966 513 13000
rect 547 12966 582 13000
rect 616 12966 651 13000
rect 685 12966 720 13000
rect 754 12966 789 13000
rect 823 12966 858 13000
rect 892 12966 927 13000
rect 961 12966 996 13000
rect 1030 12966 1065 13000
rect 1099 12966 1134 13000
rect 1168 12966 1203 13000
rect 1237 12966 1272 13000
rect 340 12932 1272 12966
rect 340 12898 375 12932
rect 409 12898 444 12932
rect 478 12898 513 12932
rect 547 12898 582 12932
rect 616 12898 651 12932
rect 685 12898 720 12932
rect 754 12898 789 12932
rect 823 12898 858 12932
rect 892 12898 927 12932
rect 961 12898 996 12932
rect 1030 12898 1065 12932
rect 1099 12898 1134 12932
rect 1168 12898 1203 12932
rect 1237 12898 1272 12932
rect 340 12864 1272 12898
rect 340 12830 375 12864
rect 409 12830 444 12864
rect 478 12830 513 12864
rect 547 12830 582 12864
rect 616 12830 651 12864
rect 685 12830 720 12864
rect 754 12830 789 12864
rect 823 12830 858 12864
rect 892 12830 927 12864
rect 961 12830 996 12864
rect 1030 12830 1065 12864
rect 1099 12830 1134 12864
rect 1168 12830 1203 12864
rect 1237 12830 1272 12864
rect 14974 12830 15032 13000
rect 15202 12830 15270 13000
rect -4920 12726 -4750 12830
rect -4886 12692 -4852 12726
rect -4818 12692 -4784 12726
rect -4920 12650 -4750 12692
rect -4886 12616 -4852 12650
rect -4818 12616 -4784 12650
rect -4920 12574 -4750 12616
rect 15100 12726 15270 12830
rect 15134 12692 15168 12726
rect 15202 12692 15236 12726
rect 15100 12650 15270 12692
rect 15134 12616 15168 12650
rect 15202 12616 15236 12650
rect 15100 12574 15270 12616
rect -4920 11543 -4750 11588
rect -4886 11509 -4852 11543
rect -4818 11509 -4784 11543
rect -4920 11464 -4750 11509
rect -4920 855 -4750 890
rect -4886 821 -4852 855
rect -4818 821 -4784 855
rect -4920 786 -4750 821
rect -4886 752 -4852 786
rect -4818 752 -4784 786
rect -4920 717 -4750 752
rect -4886 683 -4852 717
rect -4818 683 -4784 717
rect -4920 648 -4750 683
rect -4886 614 -4852 648
rect -4818 614 -4784 648
rect -4920 579 -4750 614
rect -4886 545 -4852 579
rect -4818 545 -4784 579
rect -4920 510 -4750 545
rect -4886 476 -4852 510
rect -4818 476 -4784 510
rect -4920 441 -4750 476
rect 15100 11543 15270 11588
rect 15134 11509 15168 11543
rect 15202 11509 15236 11543
rect 15100 11464 15270 11509
rect 15100 855 15270 890
rect 15134 821 15168 855
rect 15202 821 15236 855
rect 15100 786 15270 821
rect 15134 752 15168 786
rect 15202 752 15236 786
rect 15100 717 15270 752
rect 15134 683 15168 717
rect 15202 683 15236 717
rect 15100 648 15270 683
rect 15134 614 15168 648
rect 15202 614 15236 648
rect 15100 579 15270 614
rect 15134 545 15168 579
rect 15202 545 15236 579
rect 15100 510 15270 545
rect 15134 476 15168 510
rect 15202 476 15236 510
rect -4886 407 -4852 441
rect -4818 407 -4784 441
rect -4920 372 -4750 407
rect -4886 338 -4852 372
rect -4818 338 -4784 372
rect -4920 270 -4750 338
rect 15100 441 15270 476
rect 15134 407 15168 441
rect 15202 407 15236 441
rect 15100 372 15270 407
rect 15134 338 15168 372
rect 15202 338 15236 372
rect 15100 270 15270 338
rect -4920 236 -4852 270
rect -4818 236 -4783 270
rect -4749 236 -4703 270
rect -4669 236 -4634 270
rect -4600 236 -4565 270
rect -4531 236 -4496 270
rect -4462 236 -4427 270
rect -4393 236 -4358 270
rect -4324 236 -4289 270
rect -4255 236 -4220 270
rect -4186 236 -4151 270
rect -4117 236 -4082 270
rect -4048 236 -4013 270
rect -3979 236 -3913 270
rect -4920 202 -3913 236
rect -4920 168 -4852 202
rect -4818 168 -4783 202
rect -4749 168 -4703 202
rect -4669 168 -4634 202
rect -4600 168 -4565 202
rect -4531 168 -4496 202
rect -4462 168 -4427 202
rect -4393 168 -4358 202
rect -4324 168 -4289 202
rect -4255 168 -4220 202
rect -4186 168 -4151 202
rect -4117 168 -4082 202
rect -4048 168 -4013 202
rect -3979 168 -3913 202
rect -4920 134 -3913 168
rect -4920 100 -4852 134
rect -4818 100 -4783 134
rect -4749 100 -4703 134
rect -4669 100 -4634 134
rect -4600 100 -4565 134
rect -4531 100 -4496 134
rect -4462 100 -4427 134
rect -4393 100 -4358 134
rect -4324 100 -4289 134
rect -4255 100 -4220 134
rect -4186 100 -4151 134
rect -4117 100 -4082 134
rect -4048 100 -4013 134
rect -3979 100 -3913 134
rect -2995 236 -2960 270
rect -2926 236 -2891 270
rect -2857 236 -2822 270
rect -2995 202 -2822 236
rect -2995 168 -2960 202
rect -2926 168 -2891 202
rect -2857 168 -2822 202
rect -2995 134 -2822 168
rect -2995 100 -2960 134
rect -2926 100 -2891 134
rect -2857 100 -2822 134
rect 340 236 375 270
rect 409 236 444 270
rect 478 236 513 270
rect 547 236 582 270
rect 616 236 651 270
rect 685 236 720 270
rect 754 236 789 270
rect 823 236 858 270
rect 892 236 927 270
rect 961 236 996 270
rect 1030 236 1065 270
rect 1099 236 1134 270
rect 1168 236 1203 270
rect 1237 236 1272 270
rect 340 202 1272 236
rect 340 168 375 202
rect 409 168 444 202
rect 478 168 513 202
rect 547 168 582 202
rect 616 168 651 202
rect 685 168 720 202
rect 754 168 789 202
rect 823 168 858 202
rect 892 168 927 202
rect 961 168 996 202
rect 1030 168 1065 202
rect 1099 168 1134 202
rect 1168 168 1203 202
rect 1237 168 1272 202
rect 340 134 1272 168
rect 340 100 375 134
rect 409 100 444 134
rect 478 100 513 134
rect 547 100 582 134
rect 616 100 651 134
rect 685 100 720 134
rect 754 100 789 134
rect 823 100 858 134
rect 892 100 927 134
rect 961 100 996 134
rect 1030 100 1065 134
rect 1099 100 1134 134
rect 1168 100 1203 134
rect 1237 100 1272 134
rect 14974 100 15032 270
rect 15202 100 15270 270
<< mvpsubdiffcont >>
rect -4368 11796 -4334 11830
rect -4299 11796 -4265 11830
rect -4227 11796 -4193 11830
rect -4158 11796 -4124 11830
rect -4089 11796 -4055 11830
rect -4020 11796 -3986 11830
rect -3933 11796 -3899 11830
rect -3864 11796 -3830 11830
rect -3795 11796 -3761 11830
rect -3726 11796 -3692 11830
rect -3657 11796 -3623 11830
rect -3588 11796 -3554 11830
rect -3519 11796 -3485 11830
rect -3450 11796 -3416 11830
rect -3381 11796 -3347 11830
rect -3312 11796 -3278 11830
rect -3243 11796 -3209 11830
rect -3174 11796 -3140 11830
rect -3105 11796 -3071 11830
rect -3036 11796 -3002 11830
rect -2967 11796 -2933 11830
rect -2898 11796 -2864 11830
rect -2829 11796 -2795 11830
rect -2760 11796 -2726 11830
rect -2691 11796 -2657 11830
rect -2622 11796 -2588 11830
rect -2553 11796 -2519 11830
rect -2484 11796 -2450 11830
rect -2415 11796 -2381 11830
rect -2346 11796 -2312 11830
rect -2277 11796 -2243 11830
rect -2208 11796 -2174 11830
rect -2139 11796 -2105 11830
rect -2070 11796 -2036 11830
rect -2001 11796 -1967 11830
rect -1932 11796 -1898 11830
rect -1863 11796 -1829 11830
rect -4368 11728 -4334 11762
rect -4299 11728 -4265 11762
rect -4227 11728 -4193 11762
rect -4158 11728 -4124 11762
rect -4089 11728 -4055 11762
rect -4020 11728 -3986 11762
rect -3933 11728 -3899 11762
rect -3864 11728 -3830 11762
rect -3795 11728 -3761 11762
rect -3726 11728 -3692 11762
rect -3657 11728 -3623 11762
rect -3588 11728 -3554 11762
rect -3519 11728 -3485 11762
rect -3450 11728 -3416 11762
rect -3381 11728 -3347 11762
rect -3312 11728 -3278 11762
rect -3243 11728 -3209 11762
rect -3174 11728 -3140 11762
rect -3105 11728 -3071 11762
rect -3036 11728 -3002 11762
rect -2967 11728 -2933 11762
rect -2898 11728 -2864 11762
rect -2829 11728 -2795 11762
rect -2760 11728 -2726 11762
rect -2691 11728 -2657 11762
rect -2622 11728 -2588 11762
rect -2553 11728 -2519 11762
rect -2484 11728 -2450 11762
rect -2415 11728 -2381 11762
rect -2346 11728 -2312 11762
rect -2277 11728 -2243 11762
rect -2208 11728 -2174 11762
rect -2139 11728 -2105 11762
rect -2070 11728 -2036 11762
rect -2001 11728 -1967 11762
rect -1932 11728 -1898 11762
rect -1863 11728 -1829 11762
rect -4368 11660 -4334 11694
rect -4299 11660 -4265 11694
rect -4227 11660 -4193 11694
rect -4158 11660 -4124 11694
rect -4089 11660 -4055 11694
rect -4020 11660 -3986 11694
rect -3933 11660 -3899 11694
rect -3864 11660 -3830 11694
rect -3795 11660 -3761 11694
rect -3726 11660 -3692 11694
rect -3657 11660 -3623 11694
rect -3588 11660 -3554 11694
rect -3519 11660 -3485 11694
rect -3450 11660 -3416 11694
rect -3381 11660 -3347 11694
rect -3312 11660 -3278 11694
rect -3243 11660 -3209 11694
rect -3174 11660 -3140 11694
rect -3105 11660 -3071 11694
rect -3036 11660 -3002 11694
rect -2967 11660 -2933 11694
rect -2898 11660 -2864 11694
rect -2829 11660 -2795 11694
rect -2760 11660 -2726 11694
rect -2691 11660 -2657 11694
rect -2622 11660 -2588 11694
rect -2553 11660 -2519 11694
rect -2484 11660 -2450 11694
rect -2415 11660 -2381 11694
rect -2346 11660 -2312 11694
rect -2277 11660 -2243 11694
rect -2208 11660 -2174 11694
rect -2139 11660 -2105 11694
rect -2070 11660 -2036 11694
rect -2001 11660 -1967 11694
rect -1932 11660 -1898 11694
rect -1863 11660 -1829 11694
rect -1794 11660 824 11830
rect 859 11796 893 11830
rect 928 11796 962 11830
rect 997 11796 1031 11830
rect 1066 11796 1100 11830
rect 1135 11796 1169 11830
rect 1204 11796 1238 11830
rect 1273 11796 1307 11830
rect 1342 11796 1376 11830
rect 1411 11796 1445 11830
rect 1480 11796 1514 11830
rect 1549 11796 1583 11830
rect 1618 11796 1652 11830
rect 1687 11796 1721 11830
rect 1756 11796 1790 11830
rect 1825 11796 1859 11830
rect 1894 11796 1928 11830
rect 1963 11796 1997 11830
rect 2032 11796 2066 11830
rect 2101 11796 2135 11830
rect 2170 11796 2204 11830
rect 2239 11796 2273 11830
rect 859 11728 893 11762
rect 928 11728 962 11762
rect 997 11728 1031 11762
rect 1066 11728 1100 11762
rect 1135 11728 1169 11762
rect 1204 11728 1238 11762
rect 1273 11728 1307 11762
rect 1342 11728 1376 11762
rect 1411 11728 1445 11762
rect 1480 11728 1514 11762
rect 1549 11728 1583 11762
rect 1618 11728 1652 11762
rect 1687 11728 1721 11762
rect 1756 11728 1790 11762
rect 1825 11728 1859 11762
rect 1894 11728 1928 11762
rect 1963 11728 1997 11762
rect 2032 11728 2066 11762
rect 2101 11728 2135 11762
rect 2170 11728 2204 11762
rect 2239 11728 2273 11762
rect 859 11660 893 11694
rect 928 11660 962 11694
rect 997 11660 1031 11694
rect 1066 11660 1100 11694
rect 1135 11660 1169 11694
rect 1204 11660 1238 11694
rect 1273 11660 1307 11694
rect 1342 11660 1376 11694
rect 1411 11660 1445 11694
rect 1480 11660 1514 11694
rect 1549 11660 1583 11694
rect 1618 11660 1652 11694
rect 1687 11660 1721 11694
rect 1756 11660 1790 11694
rect 1825 11660 1859 11694
rect 1894 11660 1928 11694
rect 1963 11660 1997 11694
rect 2032 11660 2066 11694
rect 2101 11660 2135 11694
rect 2170 11660 2204 11694
rect 2239 11660 2273 11694
rect 2308 11660 14718 11830
rect -4436 11583 -4402 11617
rect -4368 11583 -4334 11617
rect -4300 11583 -4266 11617
rect -4436 1812 -4266 11502
rect 14616 11583 14650 11617
rect 14684 11583 14718 11617
rect 14752 11583 14786 11617
rect -4436 1743 -4402 1777
rect -4368 1743 -4334 1777
rect -4300 1743 -4266 1777
rect -4436 1674 -4402 1708
rect -4368 1674 -4334 1708
rect -4300 1674 -4266 1708
rect -4436 1605 -4402 1639
rect -4368 1605 -4334 1639
rect -4300 1605 -4266 1639
rect -4436 1536 -4402 1570
rect -4368 1536 -4334 1570
rect -4300 1536 -4266 1570
rect -4436 1467 -4402 1501
rect -4368 1467 -4334 1501
rect -4300 1467 -4266 1501
rect -4436 1398 -4402 1432
rect -4368 1398 -4334 1432
rect -4300 1398 -4266 1432
rect -4436 1329 -4402 1363
rect -4368 1329 -4334 1363
rect -4300 1329 -4266 1363
rect -4436 1260 -4402 1294
rect -4368 1260 -4334 1294
rect -4300 1260 -4266 1294
rect -4436 1191 -4402 1225
rect -4368 1191 -4334 1225
rect -4300 1191 -4266 1225
rect -4436 1122 -4402 1156
rect -4368 1122 -4334 1156
rect -4300 1122 -4266 1156
rect 14616 1812 14786 11502
rect 14616 1743 14650 1777
rect 14684 1743 14718 1777
rect 14752 1743 14786 1777
rect 14616 1674 14650 1708
rect 14684 1674 14718 1708
rect 14752 1674 14786 1708
rect 14616 1605 14650 1639
rect 14684 1605 14718 1639
rect 14752 1605 14786 1639
rect 14616 1536 14650 1570
rect 14684 1536 14718 1570
rect 14752 1536 14786 1570
rect 14616 1467 14650 1501
rect 14684 1467 14718 1501
rect 14752 1467 14786 1501
rect 14616 1398 14650 1432
rect 14684 1398 14718 1432
rect 14752 1398 14786 1432
rect 14616 1329 14650 1363
rect 14684 1329 14718 1363
rect 14752 1329 14786 1363
rect 14616 1260 14650 1294
rect 14684 1260 14718 1294
rect 14752 1260 14786 1294
rect 14616 1191 14650 1225
rect 14684 1191 14718 1225
rect 14752 1191 14786 1225
rect -4436 1053 -4402 1087
rect -4368 1053 -4334 1087
rect -4300 1053 -4266 1087
rect -4436 984 -4402 1018
rect -4368 984 -4334 1018
rect -4300 984 -4266 1018
rect 14616 1122 14650 1156
rect 14684 1122 14718 1156
rect 14752 1122 14786 1156
rect 14616 1053 14650 1087
rect 14684 1053 14718 1087
rect 14752 1053 14786 1087
rect -4436 915 -4402 949
rect -4368 915 -4334 949
rect -4300 915 -4266 949
rect -4436 846 -4402 880
rect -4368 846 -4334 880
rect -4300 846 -4266 880
rect -4436 777 -4402 811
rect -4368 777 -4334 811
rect -4300 777 -4266 811
rect -4436 708 -4402 742
rect -4368 708 -4334 742
rect -4300 708 -4266 742
rect 14616 984 14650 1018
rect 14684 984 14718 1018
rect 14752 984 14786 1018
rect 14616 915 14650 949
rect 14684 915 14718 949
rect 14752 915 14786 949
rect 14616 846 14650 880
rect 14684 846 14718 880
rect 14752 846 14786 880
rect 14616 777 14650 811
rect 14684 777 14718 811
rect 14752 777 14786 811
rect 14616 708 14650 742
rect 14684 708 14718 742
rect 14752 708 14786 742
rect -4368 606 -4334 640
rect -4299 606 -4265 640
rect -4230 606 -4196 640
rect -4158 606 -4124 640
rect -4089 606 -4055 640
rect -4020 606 -3986 640
rect -3933 606 -3899 640
rect -3864 606 -3830 640
rect -3795 606 -3761 640
rect -3726 606 -3692 640
rect -3657 606 -3623 640
rect -3588 606 -3554 640
rect -3519 606 -3485 640
rect -3450 606 -3416 640
rect -3381 606 -3347 640
rect -3312 606 -3278 640
rect -3243 606 -3209 640
rect -3174 606 -3140 640
rect -3105 606 -3071 640
rect -3036 606 -3002 640
rect -2967 606 -2933 640
rect -2898 606 -2864 640
rect -2829 606 -2795 640
rect -2760 606 -2726 640
rect -2691 606 -2657 640
rect -2622 606 -2588 640
rect -2553 606 -2519 640
rect -2484 606 -2450 640
rect -2415 606 -2381 640
rect -2346 606 -2312 640
rect -2277 606 -2243 640
rect -2208 606 -2174 640
rect -2139 606 -2105 640
rect -2070 606 -2036 640
rect -2001 606 -1967 640
rect -1932 606 -1898 640
rect -1863 606 -1829 640
rect -4368 538 -4334 572
rect -4299 538 -4265 572
rect -4230 538 -4196 572
rect -4158 538 -4124 572
rect -4089 538 -4055 572
rect -4020 538 -3986 572
rect -3933 538 -3899 572
rect -3864 538 -3830 572
rect -3795 538 -3761 572
rect -3726 538 -3692 572
rect -3657 538 -3623 572
rect -3588 538 -3554 572
rect -3519 538 -3485 572
rect -3450 538 -3416 572
rect -3381 538 -3347 572
rect -3312 538 -3278 572
rect -3243 538 -3209 572
rect -3174 538 -3140 572
rect -3105 538 -3071 572
rect -3036 538 -3002 572
rect -2967 538 -2933 572
rect -2898 538 -2864 572
rect -2829 538 -2795 572
rect -2760 538 -2726 572
rect -2691 538 -2657 572
rect -2622 538 -2588 572
rect -2553 538 -2519 572
rect -2484 538 -2450 572
rect -2415 538 -2381 572
rect -2346 538 -2312 572
rect -2277 538 -2243 572
rect -2208 538 -2174 572
rect -2139 538 -2105 572
rect -2070 538 -2036 572
rect -2001 538 -1967 572
rect -1932 538 -1898 572
rect -1863 538 -1829 572
rect -4368 470 -4334 504
rect -4299 470 -4265 504
rect -4230 470 -4196 504
rect -4158 470 -4124 504
rect -4089 470 -4055 504
rect -4020 470 -3986 504
rect -3933 470 -3899 504
rect -3864 470 -3830 504
rect -3795 470 -3761 504
rect -3726 470 -3692 504
rect -3657 470 -3623 504
rect -3588 470 -3554 504
rect -3519 470 -3485 504
rect -3450 470 -3416 504
rect -3381 470 -3347 504
rect -3312 470 -3278 504
rect -3243 470 -3209 504
rect -3174 470 -3140 504
rect -3105 470 -3071 504
rect -3036 470 -3002 504
rect -2967 470 -2933 504
rect -2898 470 -2864 504
rect -2829 470 -2795 504
rect -2760 470 -2726 504
rect -2691 470 -2657 504
rect -2622 470 -2588 504
rect -2553 470 -2519 504
rect -2484 470 -2450 504
rect -2415 470 -2381 504
rect -2346 470 -2312 504
rect -2277 470 -2243 504
rect -2208 470 -2174 504
rect -2139 470 -2105 504
rect -2070 470 -2036 504
rect -2001 470 -1967 504
rect -1932 470 -1898 504
rect -1863 470 -1829 504
rect -1794 470 824 640
rect 859 606 893 640
rect 928 606 962 640
rect 997 606 1031 640
rect 1066 606 1100 640
rect 1135 606 1169 640
rect 1204 606 1238 640
rect 1273 606 1307 640
rect 1342 606 1376 640
rect 1411 606 1445 640
rect 1480 606 1514 640
rect 1549 606 1583 640
rect 1618 606 1652 640
rect 1687 606 1721 640
rect 1756 606 1790 640
rect 1825 606 1859 640
rect 1894 606 1928 640
rect 1963 606 1997 640
rect 2032 606 2066 640
rect 2101 606 2135 640
rect 2170 606 2204 640
rect 2239 606 2273 640
rect 859 538 893 572
rect 928 538 962 572
rect 997 538 1031 572
rect 1066 538 1100 572
rect 1135 538 1169 572
rect 1204 538 1238 572
rect 1273 538 1307 572
rect 1342 538 1376 572
rect 1411 538 1445 572
rect 1480 538 1514 572
rect 1549 538 1583 572
rect 1618 538 1652 572
rect 1687 538 1721 572
rect 1756 538 1790 572
rect 1825 538 1859 572
rect 1894 538 1928 572
rect 1963 538 1997 572
rect 2032 538 2066 572
rect 2101 538 2135 572
rect 2170 538 2204 572
rect 2239 538 2273 572
rect 859 470 893 504
rect 928 470 962 504
rect 997 470 1031 504
rect 1066 470 1100 504
rect 1135 470 1169 504
rect 1204 470 1238 504
rect 1273 470 1307 504
rect 1342 470 1376 504
rect 1411 470 1445 504
rect 1480 470 1514 504
rect 1549 470 1583 504
rect 1618 470 1652 504
rect 1687 470 1721 504
rect 1756 470 1790 504
rect 1825 470 1859 504
rect 1894 470 1928 504
rect 1963 470 1997 504
rect 2032 470 2066 504
rect 2101 470 2135 504
rect 2170 470 2204 504
rect 2239 470 2273 504
rect 2308 470 14718 640
<< mvnsubdiffcont >>
rect -4852 12966 -4818 13000
rect -4783 12966 -4749 13000
rect -4703 12966 -4669 13000
rect -4634 12966 -4600 13000
rect -4565 12966 -4531 13000
rect -4496 12966 -4462 13000
rect -4427 12966 -4393 13000
rect -4358 12966 -4324 13000
rect -4289 12966 -4255 13000
rect -4220 12966 -4186 13000
rect -4151 12966 -4117 13000
rect -4082 12966 -4048 13000
rect -4013 12966 -3979 13000
rect -3944 12966 -3910 13000
rect -3875 12966 -3841 13000
rect -3806 12966 -3772 13000
rect -3737 12966 -3703 13000
rect -3668 12966 -3634 13000
rect -3599 12966 -3565 13000
rect -3530 12966 -3496 13000
rect -3461 12966 -3427 13000
rect -3392 12966 -3358 13000
rect -3323 12966 -3289 13000
rect -3254 12966 -3220 13000
rect -3185 12966 -3151 13000
rect -3116 12966 -3082 13000
rect -3029 12966 -2995 13000
rect -2960 12966 -2926 13000
rect -2891 12966 -2857 13000
rect -4852 12898 -4818 12932
rect -4783 12898 -4749 12932
rect -4703 12898 -4669 12932
rect -4634 12898 -4600 12932
rect -4565 12898 -4531 12932
rect -4496 12898 -4462 12932
rect -4427 12898 -4393 12932
rect -4358 12898 -4324 12932
rect -4289 12898 -4255 12932
rect -4220 12898 -4186 12932
rect -4151 12898 -4117 12932
rect -4082 12898 -4048 12932
rect -4013 12898 -3979 12932
rect -3944 12898 -3910 12932
rect -3875 12898 -3841 12932
rect -3806 12898 -3772 12932
rect -3737 12898 -3703 12932
rect -3668 12898 -3634 12932
rect -3599 12898 -3565 12932
rect -3530 12898 -3496 12932
rect -3461 12898 -3427 12932
rect -3392 12898 -3358 12932
rect -3323 12898 -3289 12932
rect -3254 12898 -3220 12932
rect -3185 12898 -3151 12932
rect -3116 12898 -3082 12932
rect -3029 12898 -2995 12932
rect -2960 12898 -2926 12932
rect -2891 12898 -2857 12932
rect -4852 12830 -4818 12864
rect -4783 12830 -4749 12864
rect -4703 12830 -4669 12864
rect -4634 12830 -4600 12864
rect -4565 12830 -4531 12864
rect -4496 12830 -4462 12864
rect -4427 12830 -4393 12864
rect -4358 12830 -4324 12864
rect -4289 12830 -4255 12864
rect -4220 12830 -4186 12864
rect -4151 12830 -4117 12864
rect -4082 12830 -4048 12864
rect -4013 12830 -3979 12864
rect -3944 12830 -3910 12864
rect -3875 12830 -3841 12864
rect -3806 12830 -3772 12864
rect -3737 12830 -3703 12864
rect -3668 12830 -3634 12864
rect -3599 12830 -3565 12864
rect -3530 12830 -3496 12864
rect -3461 12830 -3427 12864
rect -3392 12830 -3358 12864
rect -3323 12830 -3289 12864
rect -3254 12830 -3220 12864
rect -3185 12830 -3151 12864
rect -3116 12830 -3082 12864
rect -3029 12830 -2995 12864
rect -2960 12830 -2926 12864
rect -2891 12830 -2857 12864
rect -2822 12830 340 13000
rect 375 12966 409 13000
rect 444 12966 478 13000
rect 513 12966 547 13000
rect 582 12966 616 13000
rect 651 12966 685 13000
rect 720 12966 754 13000
rect 789 12966 823 13000
rect 858 12966 892 13000
rect 927 12966 961 13000
rect 996 12966 1030 13000
rect 1065 12966 1099 13000
rect 1134 12966 1168 13000
rect 1203 12966 1237 13000
rect 375 12898 409 12932
rect 444 12898 478 12932
rect 513 12898 547 12932
rect 582 12898 616 12932
rect 651 12898 685 12932
rect 720 12898 754 12932
rect 789 12898 823 12932
rect 858 12898 892 12932
rect 927 12898 961 12932
rect 996 12898 1030 12932
rect 1065 12898 1099 12932
rect 1134 12898 1168 12932
rect 1203 12898 1237 12932
rect 375 12830 409 12864
rect 444 12830 478 12864
rect 513 12830 547 12864
rect 582 12830 616 12864
rect 651 12830 685 12864
rect 720 12830 754 12864
rect 789 12830 823 12864
rect 858 12830 892 12864
rect 927 12830 961 12864
rect 996 12830 1030 12864
rect 1065 12830 1099 12864
rect 1134 12830 1168 12864
rect 1203 12830 1237 12864
rect 1272 12830 14974 13000
rect 15032 12830 15202 13000
rect -4920 12692 -4886 12726
rect -4852 12692 -4818 12726
rect -4784 12692 -4750 12726
rect -4920 12616 -4886 12650
rect -4852 12616 -4818 12650
rect -4784 12616 -4750 12650
rect -4920 11588 -4750 12574
rect 15100 12692 15134 12726
rect 15168 12692 15202 12726
rect 15236 12692 15270 12726
rect 15100 12616 15134 12650
rect 15168 12616 15202 12650
rect 15236 12616 15270 12650
rect -4920 11509 -4886 11543
rect -4852 11509 -4818 11543
rect -4784 11509 -4750 11543
rect -4920 890 -4750 11464
rect -4920 821 -4886 855
rect -4852 821 -4818 855
rect -4784 821 -4750 855
rect -4920 752 -4886 786
rect -4852 752 -4818 786
rect -4784 752 -4750 786
rect -4920 683 -4886 717
rect -4852 683 -4818 717
rect -4784 683 -4750 717
rect -4920 614 -4886 648
rect -4852 614 -4818 648
rect -4784 614 -4750 648
rect -4920 545 -4886 579
rect -4852 545 -4818 579
rect -4784 545 -4750 579
rect -4920 476 -4886 510
rect -4852 476 -4818 510
rect -4784 476 -4750 510
rect 15100 11588 15270 12574
rect 15100 11509 15134 11543
rect 15168 11509 15202 11543
rect 15236 11509 15270 11543
rect 15100 890 15270 11464
rect 15100 821 15134 855
rect 15168 821 15202 855
rect 15236 821 15270 855
rect 15100 752 15134 786
rect 15168 752 15202 786
rect 15236 752 15270 786
rect 15100 683 15134 717
rect 15168 683 15202 717
rect 15236 683 15270 717
rect 15100 614 15134 648
rect 15168 614 15202 648
rect 15236 614 15270 648
rect 15100 545 15134 579
rect 15168 545 15202 579
rect 15236 545 15270 579
rect 15100 476 15134 510
rect 15168 476 15202 510
rect 15236 476 15270 510
rect -4920 407 -4886 441
rect -4852 407 -4818 441
rect -4784 407 -4750 441
rect -4920 338 -4886 372
rect -4852 338 -4818 372
rect -4784 338 -4750 372
rect 15100 407 15134 441
rect 15168 407 15202 441
rect 15236 407 15270 441
rect 15100 338 15134 372
rect 15168 338 15202 372
rect 15236 338 15270 372
rect -4852 236 -4818 270
rect -4783 236 -4749 270
rect -4703 236 -4669 270
rect -4634 236 -4600 270
rect -4565 236 -4531 270
rect -4496 236 -4462 270
rect -4427 236 -4393 270
rect -4358 236 -4324 270
rect -4289 236 -4255 270
rect -4220 236 -4186 270
rect -4151 236 -4117 270
rect -4082 236 -4048 270
rect -4013 236 -3979 270
rect -4852 168 -4818 202
rect -4783 168 -4749 202
rect -4703 168 -4669 202
rect -4634 168 -4600 202
rect -4565 168 -4531 202
rect -4496 168 -4462 202
rect -4427 168 -4393 202
rect -4358 168 -4324 202
rect -4289 168 -4255 202
rect -4220 168 -4186 202
rect -4151 168 -4117 202
rect -4082 168 -4048 202
rect -4013 168 -3979 202
rect -4852 100 -4818 134
rect -4783 100 -4749 134
rect -4703 100 -4669 134
rect -4634 100 -4600 134
rect -4565 100 -4531 134
rect -4496 100 -4462 134
rect -4427 100 -4393 134
rect -4358 100 -4324 134
rect -4289 100 -4255 134
rect -4220 100 -4186 134
rect -4151 100 -4117 134
rect -4082 100 -4048 134
rect -4013 100 -3979 134
rect -3913 100 -2995 270
rect -2960 236 -2926 270
rect -2891 236 -2857 270
rect -2960 168 -2926 202
rect -2891 168 -2857 202
rect -2960 100 -2926 134
rect -2891 100 -2857 134
rect -2822 100 340 270
rect 375 236 409 270
rect 444 236 478 270
rect 513 236 547 270
rect 582 236 616 270
rect 651 236 685 270
rect 720 236 754 270
rect 789 236 823 270
rect 858 236 892 270
rect 927 236 961 270
rect 996 236 1030 270
rect 1065 236 1099 270
rect 1134 236 1168 270
rect 1203 236 1237 270
rect 375 168 409 202
rect 444 168 478 202
rect 513 168 547 202
rect 582 168 616 202
rect 651 168 685 202
rect 720 168 754 202
rect 789 168 823 202
rect 858 168 892 202
rect 927 168 961 202
rect 996 168 1030 202
rect 1065 168 1099 202
rect 1134 168 1168 202
rect 1203 168 1237 202
rect 375 100 409 134
rect 444 100 478 134
rect 513 100 547 134
rect 582 100 616 134
rect 651 100 685 134
rect 720 100 754 134
rect 789 100 823 134
rect 858 100 892 134
rect 927 100 961 134
rect 996 100 1030 134
rect 1065 100 1099 134
rect 1134 100 1168 134
rect 1203 100 1237 134
rect 1272 100 14974 270
rect 15032 100 15202 270
<< poly >>
rect -3684 11353 -3494 11476
tri -3684 11333 -3664 11353 ne
rect -3664 11333 -3514 11353
tri -3514 11333 -3494 11353 nw
rect -2392 11353 -2202 11476
tri -2392 11333 -2372 11353 ne
rect -2372 11333 -2222 11353
tri -2222 11333 -2202 11353 nw
rect -1880 11353 -1690 11476
tri -1880 11333 -1860 11353 ne
rect -1860 11333 -1710 11353
tri -1710 11333 -1690 11353 nw
rect -588 11353 -398 11476
tri -588 11333 -568 11353 ne
rect -568 11333 -418 11353
tri -418 11333 -398 11353 nw
rect -76 11353 114 11476
tri -76 11333 -56 11353 ne
rect -56 11333 94 11353
tri 94 11333 114 11353 nw
rect 1216 11353 1406 11476
tri 1216 11333 1236 11353 ne
rect 1236 11333 1386 11353
tri 1386 11333 1406 11353 nw
rect 1728 11353 1918 11476
tri 1728 11333 1748 11353 ne
rect 1748 11333 1898 11353
tri 1898 11333 1918 11353 nw
rect 3020 11353 3210 11476
tri 3020 11333 3040 11353 ne
rect 3040 11333 3190 11353
tri 3190 11333 3210 11353 nw
rect 3532 11353 3722 11476
tri 3532 11333 3552 11353 ne
rect 3552 11333 3702 11353
tri 3702 11333 3722 11353 nw
rect 4824 11353 5014 11476
tri 4824 11333 4844 11353 ne
rect 4844 11333 4994 11353
tri 4994 11333 5014 11353 nw
rect 5336 11353 5526 11476
tri 5336 11333 5356 11353 ne
rect 5356 11333 5506 11353
tri 5506 11333 5526 11353 nw
rect 6628 11353 6818 11476
tri 6628 11333 6648 11353 ne
rect 6648 11333 6798 11353
tri 6798 11333 6818 11353 nw
rect 7140 11353 7330 11476
tri 7140 11333 7160 11353 ne
rect 7160 11333 7310 11353
tri 7310 11333 7330 11353 nw
rect 8432 11353 8622 11476
tri 8432 11333 8452 11353 ne
rect 8452 11333 8602 11353
tri 8602 11333 8622 11353 nw
rect 8944 11353 9134 11476
tri 8944 11333 8964 11353 ne
rect 8964 11333 9114 11353
tri 9114 11333 9134 11353 nw
rect 10236 11353 10426 11476
tri 10236 11333 10256 11353 ne
rect 10256 11333 10406 11353
tri 10406 11333 10426 11353 nw
rect 10748 11353 10938 11476
tri 10748 11333 10768 11353 ne
rect 10768 11333 10918 11353
tri 10918 11333 10938 11353 nw
rect 12040 11353 12230 11476
tri 12040 11333 12060 11353 ne
rect 12060 11333 12210 11353
tri 12210 11333 12230 11353 nw
rect 12552 11353 12742 11476
tri 12552 11333 12572 11353 ne
rect 12572 11333 12722 11353
tri 12722 11333 12742 11353 nw
rect 13844 11353 14034 11476
tri 13844 11333 13864 11353 ne
rect 13864 11333 14014 11353
tri 14014 11333 14034 11353 nw
tri -3684 1115 -3664 1135 se
rect -3664 1115 -3514 1135
tri -3514 1115 -3494 1135 sw
rect -3684 1042 -3494 1115
rect -3684 1008 -3642 1042
rect -3608 1008 -3574 1042
rect -3540 1008 -3494 1042
rect -3684 992 -3494 1008
tri -2392 1115 -2372 1135 se
rect -2372 1115 -2222 1135
tri -2222 1115 -2202 1135 sw
rect -2392 1042 -2202 1115
rect -2392 1008 -2350 1042
rect -2316 1008 -2282 1042
rect -2248 1008 -2202 1042
rect -2392 992 -2202 1008
tri -1880 1115 -1860 1135 se
rect -1860 1115 -1710 1135
tri -1710 1115 -1690 1135 sw
rect -1880 1042 -1690 1115
rect -1880 1008 -1838 1042
rect -1804 1008 -1770 1042
rect -1736 1008 -1690 1042
rect -1880 992 -1690 1008
tri -588 1115 -568 1135 se
rect -568 1115 -418 1135
tri -418 1115 -398 1135 sw
rect -588 1042 -398 1115
rect -588 1008 -546 1042
rect -512 1008 -478 1042
rect -444 1008 -398 1042
rect -588 992 -398 1008
tri -76 1115 -56 1135 se
rect -56 1115 94 1135
tri 94 1115 114 1135 sw
rect -76 1042 114 1115
rect -76 1008 -34 1042
rect 0 1008 34 1042
rect 68 1008 114 1042
rect -76 992 114 1008
tri 1216 1115 1236 1135 se
rect 1236 1115 1386 1135
tri 1386 1115 1406 1135 sw
rect 1216 1042 1406 1115
rect 1216 1008 1258 1042
rect 1292 1008 1326 1042
rect 1360 1008 1406 1042
rect 1216 992 1406 1008
tri 1728 1115 1748 1135 se
rect 1748 1115 1898 1135
tri 1898 1115 1918 1135 sw
rect 1728 1042 1918 1115
rect 1728 1008 1770 1042
rect 1804 1008 1838 1042
rect 1872 1008 1918 1042
rect 1728 992 1918 1008
tri 3020 1115 3040 1135 se
rect 3040 1115 3190 1135
tri 3190 1115 3210 1135 sw
rect 3020 1042 3210 1115
rect 3020 1008 3062 1042
rect 3096 1008 3130 1042
rect 3164 1008 3210 1042
rect 3020 992 3210 1008
tri 3532 1115 3552 1135 se
rect 3552 1115 3702 1135
tri 3702 1115 3722 1135 sw
rect 3532 1042 3722 1115
rect 3532 1008 3574 1042
rect 3608 1008 3642 1042
rect 3676 1008 3722 1042
rect 3532 992 3722 1008
tri 4824 1115 4844 1135 se
rect 4844 1115 4994 1135
tri 4994 1115 5014 1135 sw
rect 4824 1042 5014 1115
rect 4824 1008 4866 1042
rect 4900 1008 4934 1042
rect 4968 1008 5014 1042
rect 4824 992 5014 1008
tri 5336 1115 5356 1135 se
rect 5356 1115 5506 1135
tri 5506 1115 5526 1135 sw
rect 5336 1042 5526 1115
rect 5336 1008 5378 1042
rect 5412 1008 5446 1042
rect 5480 1008 5526 1042
rect 5336 992 5526 1008
tri 6628 1115 6648 1135 se
rect 6648 1115 6798 1135
tri 6798 1115 6818 1135 sw
rect 6628 1042 6818 1115
rect 6628 1008 6670 1042
rect 6704 1008 6738 1042
rect 6772 1008 6818 1042
rect 6628 992 6818 1008
tri 7140 1115 7160 1135 se
rect 7160 1115 7310 1135
tri 7310 1115 7330 1135 sw
rect 7140 1042 7330 1115
rect 7140 1008 7182 1042
rect 7216 1008 7250 1042
rect 7284 1008 7330 1042
rect 7140 992 7330 1008
tri 8432 1115 8452 1135 se
rect 8452 1115 8602 1135
tri 8602 1115 8622 1135 sw
rect 8432 1042 8622 1115
rect 8432 1008 8474 1042
rect 8508 1008 8542 1042
rect 8576 1008 8622 1042
rect 8432 992 8622 1008
tri 8944 1115 8964 1135 se
rect 8964 1115 9114 1135
tri 9114 1115 9134 1135 sw
rect 8944 1042 9134 1115
rect 8944 1008 8986 1042
rect 9020 1008 9054 1042
rect 9088 1008 9134 1042
rect 8944 992 9134 1008
tri 10236 1115 10256 1135 se
rect 10256 1115 10406 1135
tri 10406 1115 10426 1135 sw
rect 10236 1042 10426 1115
rect 10236 1008 10278 1042
rect 10312 1008 10346 1042
rect 10380 1008 10426 1042
rect 10236 992 10426 1008
tri 10748 1115 10768 1135 se
rect 10768 1115 10918 1135
tri 10918 1115 10938 1135 sw
rect 10748 1042 10938 1115
rect 10748 1008 10790 1042
rect 10824 1008 10858 1042
rect 10892 1008 10938 1042
rect 10748 992 10938 1008
tri 12040 1115 12060 1135 se
rect 12060 1115 12210 1135
tri 12210 1115 12230 1135 sw
rect 12040 1042 12230 1115
rect 12040 1008 12082 1042
rect 12116 1008 12150 1042
rect 12184 1008 12230 1042
rect 12040 992 12230 1008
tri 12552 1115 12572 1135 se
rect 12572 1115 12722 1135
tri 12722 1115 12742 1135 sw
rect 12552 1042 12742 1115
rect 12552 1008 12594 1042
rect 12628 1008 12662 1042
rect 12696 1008 12742 1042
rect 12552 992 12742 1008
tri 13844 1115 13864 1135 se
rect 13864 1115 14014 1135
tri 14014 1115 14034 1135 sw
rect 13844 1042 14034 1115
rect 13844 1008 13886 1042
rect 13920 1008 13954 1042
rect 13988 1008 14034 1042
rect 13844 992 14034 1008
<< polycont >>
rect -3642 1008 -3608 1042
rect -3574 1008 -3540 1042
rect -2350 1008 -2316 1042
rect -2282 1008 -2248 1042
rect -1838 1008 -1804 1042
rect -1770 1008 -1736 1042
rect -546 1008 -512 1042
rect -478 1008 -444 1042
rect -34 1008 0 1042
rect 34 1008 68 1042
rect 1258 1008 1292 1042
rect 1326 1008 1360 1042
rect 1770 1008 1804 1042
rect 1838 1008 1872 1042
rect 3062 1008 3096 1042
rect 3130 1008 3164 1042
rect 3574 1008 3608 1042
rect 3642 1008 3676 1042
rect 4866 1008 4900 1042
rect 4934 1008 4968 1042
rect 5378 1008 5412 1042
rect 5446 1008 5480 1042
rect 6670 1008 6704 1042
rect 6738 1008 6772 1042
rect 7182 1008 7216 1042
rect 7250 1008 7284 1042
rect 8474 1008 8508 1042
rect 8542 1008 8576 1042
rect 8986 1008 9020 1042
rect 9054 1008 9088 1042
rect 10278 1008 10312 1042
rect 10346 1008 10380 1042
rect 10790 1008 10824 1042
rect 10858 1008 10892 1042
rect 12082 1008 12116 1042
rect 12150 1008 12184 1042
rect 12594 1008 12628 1042
rect 12662 1008 12696 1042
rect 13886 1008 13920 1042
rect 13954 1008 13988 1042
<< locali >>
rect -4920 12966 -4852 13000
rect -4818 12966 -4783 13000
rect -4749 12966 -4703 13000
rect -4669 12966 -4634 13000
rect -4600 12966 -4565 13000
rect -4531 12966 -4496 13000
rect -4462 12966 -4427 13000
rect -4393 12966 -4358 13000
rect -4324 12966 -4289 13000
rect -4255 12966 -4220 13000
rect -4186 12966 -4151 13000
rect -4117 12966 -4082 13000
rect -4048 12966 -4013 13000
rect -3979 12966 -3944 13000
rect -3910 12966 -3875 13000
rect -3841 12966 -3806 13000
rect -3772 12966 -3737 13000
rect -3703 12966 -3668 13000
rect -3634 12966 -3599 13000
rect -3565 12966 -3530 13000
rect -3496 12966 -3461 13000
rect -3427 12966 -3392 13000
rect -3358 12966 -3323 13000
rect -3289 12966 -3254 13000
rect -3220 12966 -3185 13000
rect -3151 12966 -3116 13000
rect -3082 12966 -3029 13000
rect -2995 12966 -2960 13000
rect -2926 12966 -2891 13000
rect -2857 12966 -2822 13000
rect -4920 12932 -2822 12966
rect -4920 12898 -4852 12932
rect -4818 12898 -4783 12932
rect -4749 12898 -4703 12932
rect -4669 12898 -4634 12932
rect -4600 12898 -4565 12932
rect -4531 12898 -4496 12932
rect -4462 12898 -4427 12932
rect -4393 12898 -4358 12932
rect -4324 12898 -4289 12932
rect -4255 12898 -4220 12932
rect -4186 12898 -4151 12932
rect -4117 12898 -4082 12932
rect -4048 12898 -4013 12932
rect -3979 12898 -3944 12932
rect -3910 12898 -3875 12932
rect -3841 12898 -3806 12932
rect -3772 12898 -3737 12932
rect -3703 12898 -3668 12932
rect -3634 12898 -3599 12932
rect -3565 12898 -3530 12932
rect -3496 12898 -3461 12932
rect -3427 12898 -3392 12932
rect -3358 12898 -3323 12932
rect -3289 12898 -3254 12932
rect -3220 12898 -3185 12932
rect -3151 12898 -3116 12932
rect -3082 12898 -3029 12932
rect -2995 12898 -2960 12932
rect -2926 12898 -2891 12932
rect -2857 12898 -2822 12932
rect -4920 12864 -2822 12898
rect -4920 12830 -4852 12864
rect -4818 12830 -4783 12864
rect -4749 12830 -4703 12864
rect -4669 12830 -4634 12864
rect -4600 12830 -4565 12864
rect -4531 12830 -4496 12864
rect -4462 12830 -4427 12864
rect -4393 12830 -4358 12864
rect -4324 12830 -4289 12864
rect -4255 12830 -4220 12864
rect -4186 12830 -4151 12864
rect -4117 12830 -4082 12864
rect -4048 12830 -4013 12864
rect -3979 12830 -3944 12864
rect -3910 12830 -3875 12864
rect -3841 12830 -3806 12864
rect -3772 12830 -3737 12864
rect -3703 12830 -3668 12864
rect -3634 12830 -3599 12864
rect -3565 12830 -3530 12864
rect -3496 12830 -3461 12864
rect -3427 12830 -3392 12864
rect -3358 12830 -3323 12864
rect -3289 12830 -3254 12864
rect -3220 12830 -3185 12864
rect -3151 12830 -3116 12864
rect -3082 12830 -3029 12864
rect -2995 12830 -2960 12864
rect -2926 12830 -2891 12864
rect -2857 12830 -2822 12864
rect 340 12966 375 13000
rect 409 12966 444 13000
rect 478 12966 513 13000
rect 547 12966 582 13000
rect 616 12966 651 13000
rect 685 12966 720 13000
rect 754 12966 789 13000
rect 823 12966 858 13000
rect 892 12966 927 13000
rect 961 12966 996 13000
rect 1030 12966 1065 13000
rect 1099 12966 1134 13000
rect 1168 12966 1203 13000
rect 1237 12966 1272 13000
rect 340 12932 1272 12966
rect 340 12898 375 12932
rect 409 12898 444 12932
rect 478 12898 513 12932
rect 547 12898 582 12932
rect 616 12898 651 12932
rect 685 12898 720 12932
rect 754 12898 789 12932
rect 823 12898 858 12932
rect 892 12898 927 12932
rect 961 12898 996 12932
rect 1030 12898 1065 12932
rect 1099 12898 1134 12932
rect 1168 12898 1203 12932
rect 1237 12898 1272 12932
rect 340 12864 1272 12898
rect 340 12830 375 12864
rect 409 12830 444 12864
rect 478 12830 513 12864
rect 547 12830 582 12864
rect 616 12830 651 12864
rect 685 12830 720 12864
rect 754 12830 789 12864
rect 823 12830 858 12864
rect 892 12830 927 12864
rect 961 12830 996 12864
rect 1030 12830 1065 12864
rect 1099 12830 1134 12864
rect 1168 12830 1203 12864
rect 1237 12830 1272 12864
rect 14974 12830 15032 13000
rect 15202 12830 15270 13000
rect -4920 12757 -4750 12830
rect -4920 12726 -4888 12757
rect -4782 12726 -4750 12757
rect -4920 12650 -4888 12692
rect -4782 12650 -4750 12692
rect -4920 12574 -4888 12616
rect -4782 12574 -4750 12616
rect 15100 12757 15270 12830
rect 15100 12726 15132 12757
rect 15238 12726 15270 12757
rect 15100 12650 15132 12692
rect 15238 12650 15270 12692
rect 15100 12574 15132 12616
rect 15238 12574 15270 12616
rect -4920 11562 -4750 11588
rect -4920 11543 -4888 11562
rect -4854 11543 -4816 11562
rect -4782 11543 -4750 11562
rect -4854 11528 -4852 11543
rect -4886 11509 -4852 11528
rect -4818 11528 -4816 11543
rect -4818 11509 -4784 11528
rect -4920 11483 -4750 11509
rect -4920 11464 -4888 11483
rect -4782 11464 -4750 11483
rect -4920 878 -4888 890
rect -4854 878 -4816 890
rect -4782 878 -4750 890
rect -4920 855 -4750 878
rect -4886 839 -4852 855
rect -4854 821 -4852 839
rect -4818 839 -4784 855
rect -4818 821 -4816 839
rect -4920 805 -4888 821
rect -4854 805 -4816 821
rect -4782 805 -4750 821
rect -4920 786 -4750 805
rect -4886 766 -4852 786
rect -4854 752 -4852 766
rect -4818 766 -4784 786
rect -4818 752 -4816 766
rect -4920 732 -4888 752
rect -4854 732 -4816 752
rect -4782 732 -4750 752
rect -4920 717 -4750 732
rect -4886 693 -4852 717
rect -4854 683 -4852 693
rect -4818 693 -4784 717
rect -4818 683 -4816 693
rect -4920 659 -4888 683
rect -4854 659 -4816 683
rect -4782 659 -4750 683
rect -4920 648 -4750 659
rect -4886 620 -4852 648
rect -4854 614 -4852 620
rect -4818 620 -4784 648
rect -4818 614 -4816 620
rect -4920 586 -4888 614
rect -4854 586 -4816 614
rect -4782 586 -4750 614
rect -4920 579 -4750 586
rect -4886 547 -4852 579
rect -4854 545 -4852 547
rect -4818 547 -4784 579
rect -4818 545 -4816 547
rect -4920 513 -4888 545
rect -4854 513 -4816 545
rect -4782 513 -4750 545
rect -4920 510 -4750 513
rect -4886 476 -4852 510
rect -4818 476 -4784 510
rect -4920 474 -4750 476
rect -4920 441 -4888 474
rect -4854 441 -4816 474
rect -4782 441 -4750 474
rect -4436 11796 -4368 11830
rect -4334 11796 -4299 11830
rect -4265 11796 -4227 11830
rect -4193 11796 -4158 11830
rect -4124 11796 -4089 11830
rect -4055 11796 -4020 11830
rect -3986 11796 -3933 11830
rect -3899 11796 -3864 11830
rect -3830 11796 -3795 11830
rect -3761 11796 -3726 11830
rect -3692 11796 -3657 11830
rect -3623 11796 -3588 11830
rect -3554 11796 -3519 11830
rect -3485 11796 -3450 11830
rect -3416 11796 -3381 11830
rect -3347 11796 -3312 11830
rect -3278 11796 -3243 11830
rect -3209 11796 -3174 11830
rect -3140 11796 -3105 11830
rect -3071 11796 -3036 11830
rect -3002 11796 -2967 11830
rect -2933 11796 -2898 11830
rect -2864 11796 -2829 11830
rect -2795 11796 -2760 11830
rect -2726 11796 -2691 11830
rect -2657 11796 -2622 11830
rect -2588 11796 -2553 11830
rect -2519 11796 -2484 11830
rect -2450 11796 -2415 11830
rect -2381 11796 -2346 11830
rect -2312 11796 -2277 11830
rect -2243 11796 -2208 11830
rect -2174 11796 -2139 11830
rect -2105 11796 -2070 11830
rect -2036 11796 -2001 11830
rect -1967 11796 -1932 11830
rect -1898 11796 -1863 11830
rect -1829 11796 -1794 11830
rect -4436 11762 -1794 11796
rect -4436 11728 -4368 11762
rect -4334 11728 -4299 11762
rect -4265 11728 -4227 11762
rect -4193 11728 -4158 11762
rect -4124 11728 -4089 11762
rect -4055 11728 -4020 11762
rect -3986 11728 -3933 11762
rect -3899 11728 -3864 11762
rect -3830 11728 -3795 11762
rect -3761 11728 -3726 11762
rect -3692 11728 -3657 11762
rect -3623 11728 -3588 11762
rect -3554 11728 -3519 11762
rect -3485 11728 -3450 11762
rect -3416 11728 -3381 11762
rect -3347 11728 -3312 11762
rect -3278 11728 -3243 11762
rect -3209 11728 -3174 11762
rect -3140 11728 -3105 11762
rect -3071 11728 -3036 11762
rect -3002 11728 -2967 11762
rect -2933 11728 -2898 11762
rect -2864 11728 -2829 11762
rect -2795 11728 -2760 11762
rect -2726 11728 -2691 11762
rect -2657 11728 -2622 11762
rect -2588 11728 -2553 11762
rect -2519 11728 -2484 11762
rect -2450 11728 -2415 11762
rect -2381 11728 -2346 11762
rect -2312 11728 -2277 11762
rect -2243 11728 -2208 11762
rect -2174 11728 -2139 11762
rect -2105 11728 -2070 11762
rect -2036 11728 -2001 11762
rect -1967 11728 -1932 11762
rect -1898 11728 -1863 11762
rect -1829 11728 -1794 11762
rect -4436 11694 -1794 11728
rect -4436 11660 -4368 11694
rect -4334 11660 -4299 11694
rect -4265 11660 -4227 11694
rect -4193 11660 -4158 11694
rect -4124 11660 -4089 11694
rect -4055 11660 -4020 11694
rect -3986 11660 -3933 11694
rect -3899 11660 -3864 11694
rect -3830 11660 -3795 11694
rect -3761 11660 -3726 11694
rect -3692 11660 -3657 11694
rect -3623 11660 -3588 11694
rect -3554 11660 -3519 11694
rect -3485 11660 -3450 11694
rect -3416 11660 -3381 11694
rect -3347 11660 -3312 11694
rect -3278 11660 -3243 11694
rect -3209 11660 -3174 11694
rect -3140 11660 -3105 11694
rect -3071 11660 -3036 11694
rect -3002 11660 -2967 11694
rect -2933 11660 -2898 11694
rect -2864 11660 -2829 11694
rect -2795 11660 -2760 11694
rect -2726 11660 -2691 11694
rect -2657 11660 -2622 11694
rect -2588 11660 -2553 11694
rect -2519 11660 -2484 11694
rect -2450 11660 -2415 11694
rect -2381 11660 -2346 11694
rect -2312 11660 -2277 11694
rect -2243 11660 -2208 11694
rect -2174 11660 -2139 11694
rect -2105 11660 -2070 11694
rect -2036 11660 -2001 11694
rect -1967 11660 -1932 11694
rect -1898 11660 -1863 11694
rect -1829 11660 -1794 11694
rect 824 11796 859 11830
rect 893 11796 928 11830
rect 962 11796 997 11830
rect 1031 11796 1066 11830
rect 1100 11796 1135 11830
rect 1169 11796 1204 11830
rect 1238 11796 1273 11830
rect 1307 11796 1342 11830
rect 1376 11796 1411 11830
rect 1445 11796 1480 11830
rect 1514 11796 1549 11830
rect 1583 11796 1618 11830
rect 1652 11796 1687 11830
rect 1721 11796 1756 11830
rect 1790 11796 1825 11830
rect 1859 11796 1894 11830
rect 1928 11796 1963 11830
rect 1997 11796 2032 11830
rect 2066 11796 2101 11830
rect 2135 11796 2170 11830
rect 2204 11796 2239 11830
rect 2273 11796 2308 11830
rect 824 11762 2308 11796
rect 824 11728 859 11762
rect 893 11728 928 11762
rect 962 11728 997 11762
rect 1031 11728 1066 11762
rect 1100 11728 1135 11762
rect 1169 11728 1204 11762
rect 1238 11728 1273 11762
rect 1307 11728 1342 11762
rect 1376 11728 1411 11762
rect 1445 11728 1480 11762
rect 1514 11728 1549 11762
rect 1583 11728 1618 11762
rect 1652 11728 1687 11762
rect 1721 11728 1756 11762
rect 1790 11728 1825 11762
rect 1859 11728 1894 11762
rect 1928 11728 1963 11762
rect 1997 11728 2032 11762
rect 2066 11728 2101 11762
rect 2135 11728 2170 11762
rect 2204 11728 2239 11762
rect 2273 11728 2308 11762
rect 824 11694 2308 11728
rect 824 11660 859 11694
rect 893 11660 928 11694
rect 962 11660 997 11694
rect 1031 11660 1066 11694
rect 1100 11660 1135 11694
rect 1169 11660 1204 11694
rect 1238 11660 1273 11694
rect 1307 11660 1342 11694
rect 1376 11660 1411 11694
rect 1445 11660 1480 11694
rect 1514 11660 1549 11694
rect 1583 11660 1618 11694
rect 1652 11660 1687 11694
rect 1721 11660 1756 11694
rect 1790 11660 1825 11694
rect 1859 11660 1894 11694
rect 1928 11660 1963 11694
rect 1997 11660 2032 11694
rect 2066 11660 2101 11694
rect 2135 11660 2170 11694
rect 2204 11660 2239 11694
rect 2273 11660 2308 11694
rect 14718 11660 14786 11830
rect -4436 11617 -4266 11660
rect -4402 11583 -4368 11617
rect -4334 11583 -4300 11617
rect -4436 11502 -4266 11583
rect 14616 11617 14786 11660
rect 14650 11583 14684 11617
rect 14718 11583 14752 11617
rect 14616 11502 14786 11583
rect -4436 1777 -4266 1812
rect -4402 1743 -4368 1777
rect -4334 1743 -4300 1777
rect -4436 1708 -4266 1743
rect -4402 1674 -4368 1708
rect -4334 1674 -4300 1708
rect -4436 1639 -4266 1674
rect -4402 1605 -4368 1639
rect -4334 1605 -4300 1639
rect -4436 1570 -4266 1605
rect -4402 1536 -4368 1570
rect -4334 1536 -4300 1570
rect -4436 1501 -4266 1536
rect -4402 1467 -4368 1501
rect -4334 1467 -4300 1501
rect -4436 1432 -4266 1467
rect -4402 1398 -4368 1432
rect -4334 1398 -4300 1432
rect -4436 1363 -4266 1398
rect -4402 1329 -4368 1363
rect -4334 1329 -4300 1363
rect -4436 1294 -4266 1329
rect -4402 1260 -4368 1294
rect -4334 1260 -4300 1294
rect -4436 1225 -4266 1260
rect -4402 1191 -4368 1225
rect -4334 1191 -4300 1225
rect -4436 1156 -4266 1191
rect -4402 1122 -4368 1156
rect -4334 1122 -4300 1156
rect -4145 11233 -3545 11333
rect -4145 3279 -3898 11233
rect -3792 3279 -3545 11233
rect -4145 3270 -3545 3279
rect -4145 3240 -3896 3270
rect -4145 3206 -3898 3240
rect -3862 3236 -3828 3270
rect -3794 3240 -3545 3270
rect -3864 3206 -3826 3236
rect -3792 3206 -3545 3240
rect -4145 3201 -3545 3206
rect -4145 3167 -3896 3201
rect -3862 3167 -3828 3201
rect -3794 3167 -3545 3201
rect -4145 3133 -3898 3167
rect -3864 3133 -3826 3167
rect -3792 3133 -3545 3167
rect -4145 3132 -3545 3133
rect -4145 3098 -3896 3132
rect -3862 3098 -3828 3132
rect -3794 3098 -3545 3132
rect -4145 3094 -3545 3098
rect -4145 3060 -3898 3094
rect -3864 3063 -3826 3094
rect -4145 3029 -3896 3060
rect -3862 3029 -3828 3063
rect -3792 3060 -3545 3094
rect -3794 3029 -3545 3060
rect -4145 3021 -3545 3029
rect -4145 2987 -3898 3021
rect -3864 2994 -3826 3021
rect -4145 2960 -3896 2987
rect -3862 2960 -3828 2994
rect -3792 2987 -3545 3021
rect -3794 2960 -3545 2987
rect -4145 2948 -3545 2960
rect -4145 2914 -3898 2948
rect -3864 2925 -3826 2948
rect -4145 2891 -3896 2914
rect -3862 2891 -3828 2925
rect -3792 2914 -3545 2948
rect -3794 2891 -3545 2914
rect -4145 2875 -3545 2891
rect -4145 2841 -3898 2875
rect -3864 2856 -3826 2875
rect -4145 2822 -3896 2841
rect -3862 2822 -3828 2856
rect -3792 2841 -3545 2875
rect -3794 2822 -3545 2841
rect -4145 2802 -3545 2822
rect -4145 2768 -3898 2802
rect -3864 2787 -3826 2802
rect -4145 2753 -3896 2768
rect -3862 2753 -3828 2787
rect -3792 2768 -3545 2802
rect -3794 2753 -3545 2768
rect -4145 2729 -3545 2753
rect -4145 2695 -3898 2729
rect -3864 2718 -3826 2729
rect -4145 2684 -3896 2695
rect -3862 2684 -3828 2718
rect -3792 2695 -3545 2729
rect -3794 2684 -3545 2695
rect -4145 2656 -3545 2684
rect -4145 2622 -3898 2656
rect -3864 2649 -3826 2656
rect -4145 2615 -3896 2622
rect -3862 2615 -3828 2649
rect -3792 2622 -3545 2656
rect -3794 2615 -3545 2622
rect -4145 2583 -3545 2615
rect -4145 2549 -3898 2583
rect -3864 2580 -3826 2583
rect -4145 2546 -3896 2549
rect -3862 2546 -3828 2580
rect -3792 2549 -3545 2583
rect -3794 2546 -3545 2549
rect -4145 2511 -3545 2546
rect -4145 2510 -3896 2511
rect -4145 2476 -3898 2510
rect -3862 2477 -3828 2511
rect -3794 2510 -3545 2511
rect -3864 2476 -3826 2477
rect -3792 2476 -3545 2510
rect -4145 2442 -3545 2476
rect -4145 2437 -3896 2442
rect -4145 2403 -3898 2437
rect -3862 2408 -3828 2442
rect -3794 2437 -3545 2442
rect -3864 2403 -3826 2408
rect -3792 2403 -3545 2437
rect -4145 2373 -3545 2403
rect -4145 2364 -3896 2373
rect -4145 2330 -3898 2364
rect -3862 2339 -3828 2373
rect -3794 2364 -3545 2373
rect -3864 2330 -3826 2339
rect -3792 2330 -3545 2364
rect -4145 2304 -3545 2330
rect -4145 2291 -3896 2304
rect -4145 2257 -3898 2291
rect -3862 2270 -3828 2304
rect -3794 2291 -3545 2304
rect -3864 2257 -3826 2270
rect -3792 2257 -3545 2291
rect -4145 2235 -3545 2257
rect -4145 2218 -3896 2235
rect -4145 2184 -3898 2218
rect -3862 2201 -3828 2235
rect -3794 2218 -3545 2235
rect -3864 2184 -3826 2201
rect -3792 2184 -3545 2218
rect -4145 2166 -3545 2184
rect -4145 2145 -3896 2166
rect -4145 2111 -3898 2145
rect -3862 2132 -3828 2166
rect -3794 2145 -3545 2166
rect -3864 2111 -3826 2132
rect -3792 2111 -3545 2145
rect -4145 2097 -3545 2111
rect -4145 2072 -3896 2097
rect -4145 2038 -3898 2072
rect -3862 2063 -3828 2097
rect -3794 2072 -3545 2097
rect -3864 2038 -3826 2063
rect -3792 2038 -3545 2072
rect -4145 2028 -3545 2038
rect -4145 1999 -3896 2028
rect -4145 1965 -3898 1999
rect -3862 1994 -3828 2028
rect -3794 1999 -3545 2028
rect -3864 1965 -3826 1994
rect -3792 1965 -3545 1999
rect -4145 1959 -3545 1965
rect -4145 1926 -3896 1959
rect -4145 1892 -3898 1926
rect -3862 1925 -3828 1959
rect -3794 1926 -3545 1959
rect -3864 1892 -3826 1925
rect -3792 1892 -3545 1926
rect -4145 1890 -3545 1892
rect -4145 1856 -3896 1890
rect -3862 1856 -3828 1890
rect -3794 1856 -3545 1890
rect -4145 1853 -3545 1856
rect -4145 1819 -3898 1853
rect -3864 1821 -3826 1853
rect -4145 1787 -3896 1819
rect -3862 1787 -3828 1821
rect -3792 1819 -3545 1853
rect -3794 1787 -3545 1819
rect -4145 1780 -3545 1787
rect -4145 1746 -3898 1780
rect -3864 1752 -3826 1780
rect -4145 1718 -3896 1746
rect -3862 1718 -3828 1752
rect -3792 1746 -3545 1780
rect -3794 1718 -3545 1746
rect -4145 1707 -3545 1718
rect -4145 1673 -3898 1707
rect -3864 1683 -3826 1707
rect -4145 1649 -3896 1673
rect -3862 1649 -3828 1683
rect -3792 1673 -3545 1707
rect -3794 1649 -3545 1673
rect -4145 1634 -3545 1649
rect -4145 1600 -3898 1634
rect -3864 1614 -3826 1634
rect -4145 1580 -3896 1600
rect -3862 1580 -3828 1614
rect -3792 1600 -3545 1634
rect -3794 1580 -3545 1600
rect -4145 1561 -3545 1580
rect -4145 1527 -3898 1561
rect -3864 1545 -3826 1561
rect -4145 1511 -3896 1527
rect -3862 1511 -3828 1545
rect -3792 1527 -3545 1561
rect -3794 1511 -3545 1527
rect -4145 1488 -3545 1511
rect -4145 1454 -3898 1488
rect -3864 1476 -3826 1488
rect -4145 1442 -3896 1454
rect -3862 1442 -3828 1476
rect -3792 1454 -3545 1488
rect -3794 1442 -3545 1454
rect -4145 1415 -3545 1442
rect -4145 1381 -3898 1415
rect -3864 1407 -3826 1415
rect -4145 1373 -3896 1381
rect -3862 1373 -3828 1407
rect -3792 1381 -3545 1415
rect -3794 1373 -3545 1381
rect -4145 1342 -3545 1373
rect -4145 1308 -3898 1342
rect -3864 1338 -3826 1342
rect -4145 1304 -3896 1308
rect -3862 1304 -3828 1338
rect -3792 1308 -3545 1342
rect -3794 1304 -3545 1308
rect -4145 1269 -3545 1304
rect -4145 1235 -3898 1269
rect -3862 1235 -3828 1269
rect -3792 1235 -3545 1269
rect -4145 1135 -3545 1235
rect -3243 11233 -2643 11333
rect -3243 3279 -2996 11233
rect -2890 3279 -2643 11233
rect -3243 3270 -2643 3279
rect -3243 3240 -2994 3270
rect -3243 3206 -2996 3240
rect -2960 3236 -2926 3270
rect -2892 3240 -2643 3270
rect -2962 3206 -2924 3236
rect -2890 3206 -2643 3240
rect -3243 3201 -2643 3206
rect -3243 3167 -2994 3201
rect -2960 3167 -2926 3201
rect -2892 3167 -2643 3201
rect -3243 3133 -2996 3167
rect -2962 3133 -2924 3167
rect -2890 3133 -2643 3167
rect -3243 3132 -2643 3133
rect -3243 3098 -2994 3132
rect -2960 3098 -2926 3132
rect -2892 3098 -2643 3132
rect -3243 3094 -2643 3098
rect -3243 3060 -2996 3094
rect -2962 3063 -2924 3094
rect -3243 3029 -2994 3060
rect -2960 3029 -2926 3063
rect -2890 3060 -2643 3094
rect -2892 3029 -2643 3060
rect -3243 3021 -2643 3029
rect -3243 2987 -2996 3021
rect -2962 2994 -2924 3021
rect -3243 2960 -2994 2987
rect -2960 2960 -2926 2994
rect -2890 2987 -2643 3021
rect -2892 2960 -2643 2987
rect -3243 2948 -2643 2960
rect -3243 2914 -2996 2948
rect -2962 2925 -2924 2948
rect -3243 2891 -2994 2914
rect -2960 2891 -2926 2925
rect -2890 2914 -2643 2948
rect -2892 2891 -2643 2914
rect -3243 2875 -2643 2891
rect -3243 2841 -2996 2875
rect -2962 2856 -2924 2875
rect -3243 2822 -2994 2841
rect -2960 2822 -2926 2856
rect -2890 2841 -2643 2875
rect -2892 2822 -2643 2841
rect -3243 2802 -2643 2822
rect -3243 2768 -2996 2802
rect -2962 2787 -2924 2802
rect -3243 2753 -2994 2768
rect -2960 2753 -2926 2787
rect -2890 2768 -2643 2802
rect -2892 2753 -2643 2768
rect -3243 2729 -2643 2753
rect -3243 2695 -2996 2729
rect -2962 2718 -2924 2729
rect -3243 2684 -2994 2695
rect -2960 2684 -2926 2718
rect -2890 2695 -2643 2729
rect -2892 2684 -2643 2695
rect -3243 2656 -2643 2684
rect -3243 2622 -2996 2656
rect -2962 2649 -2924 2656
rect -3243 2615 -2994 2622
rect -2960 2615 -2926 2649
rect -2890 2622 -2643 2656
rect -2892 2615 -2643 2622
rect -3243 2583 -2643 2615
rect -3243 2549 -2996 2583
rect -2962 2580 -2924 2583
rect -3243 2546 -2994 2549
rect -2960 2546 -2926 2580
rect -2890 2549 -2643 2583
rect -2892 2546 -2643 2549
rect -3243 2511 -2643 2546
rect -3243 2510 -2994 2511
rect -3243 2476 -2996 2510
rect -2960 2477 -2926 2511
rect -2892 2510 -2643 2511
rect -2962 2476 -2924 2477
rect -2890 2476 -2643 2510
rect -3243 2442 -2643 2476
rect -3243 2437 -2994 2442
rect -3243 2403 -2996 2437
rect -2960 2408 -2926 2442
rect -2892 2437 -2643 2442
rect -2962 2403 -2924 2408
rect -2890 2403 -2643 2437
rect -3243 2373 -2643 2403
rect -3243 2364 -2994 2373
rect -3243 2330 -2996 2364
rect -2960 2339 -2926 2373
rect -2892 2364 -2643 2373
rect -2962 2330 -2924 2339
rect -2890 2330 -2643 2364
rect -3243 2304 -2643 2330
rect -3243 2291 -2994 2304
rect -3243 2257 -2996 2291
rect -2960 2270 -2926 2304
rect -2892 2291 -2643 2304
rect -2962 2257 -2924 2270
rect -2890 2257 -2643 2291
rect -3243 2235 -2643 2257
rect -3243 2218 -2994 2235
rect -3243 2184 -2996 2218
rect -2960 2201 -2926 2235
rect -2892 2218 -2643 2235
rect -2962 2184 -2924 2201
rect -2890 2184 -2643 2218
rect -3243 2166 -2643 2184
rect -3243 2145 -2994 2166
rect -3243 2111 -2996 2145
rect -2960 2132 -2926 2166
rect -2892 2145 -2643 2166
rect -2962 2111 -2924 2132
rect -2890 2111 -2643 2145
rect -3243 2097 -2643 2111
rect -3243 2072 -2994 2097
rect -3243 2038 -2996 2072
rect -2960 2063 -2926 2097
rect -2892 2072 -2643 2097
rect -2962 2038 -2924 2063
rect -2890 2038 -2643 2072
rect -3243 2028 -2643 2038
rect -3243 1999 -2994 2028
rect -3243 1965 -2996 1999
rect -2960 1994 -2926 2028
rect -2892 1999 -2643 2028
rect -2962 1965 -2924 1994
rect -2890 1965 -2643 1999
rect -3243 1959 -2643 1965
rect -3243 1926 -2994 1959
rect -3243 1892 -2996 1926
rect -2960 1925 -2926 1959
rect -2892 1926 -2643 1959
rect -2962 1892 -2924 1925
rect -2890 1892 -2643 1926
rect -3243 1890 -2643 1892
rect -3243 1856 -2994 1890
rect -2960 1856 -2926 1890
rect -2892 1856 -2643 1890
rect -3243 1853 -2643 1856
rect -3243 1819 -2996 1853
rect -2962 1821 -2924 1853
rect -3243 1787 -2994 1819
rect -2960 1787 -2926 1821
rect -2890 1819 -2643 1853
rect -2892 1787 -2643 1819
rect -3243 1780 -2643 1787
rect -3243 1746 -2996 1780
rect -2962 1752 -2924 1780
rect -3243 1718 -2994 1746
rect -2960 1718 -2926 1752
rect -2890 1746 -2643 1780
rect -2892 1718 -2643 1746
rect -3243 1707 -2643 1718
rect -3243 1673 -2996 1707
rect -2962 1683 -2924 1707
rect -3243 1649 -2994 1673
rect -2960 1649 -2926 1683
rect -2890 1673 -2643 1707
rect -2892 1649 -2643 1673
rect -3243 1634 -2643 1649
rect -3243 1600 -2996 1634
rect -2962 1614 -2924 1634
rect -3243 1580 -2994 1600
rect -2960 1580 -2926 1614
rect -2890 1600 -2643 1634
rect -2892 1580 -2643 1600
rect -3243 1561 -2643 1580
rect -3243 1527 -2996 1561
rect -2962 1545 -2924 1561
rect -3243 1511 -2994 1527
rect -2960 1511 -2926 1545
rect -2890 1527 -2643 1561
rect -2892 1511 -2643 1527
rect -3243 1488 -2643 1511
rect -3243 1454 -2996 1488
rect -2962 1476 -2924 1488
rect -3243 1442 -2994 1454
rect -2960 1442 -2926 1476
rect -2890 1454 -2643 1488
rect -2892 1442 -2643 1454
rect -3243 1415 -2643 1442
rect -3243 1381 -2996 1415
rect -2962 1407 -2924 1415
rect -3243 1373 -2994 1381
rect -2960 1373 -2926 1407
rect -2890 1381 -2643 1415
rect -2892 1373 -2643 1381
rect -3243 1342 -2643 1373
rect -3243 1308 -2996 1342
rect -2962 1338 -2924 1342
rect -3243 1304 -2994 1308
rect -2960 1304 -2926 1338
rect -2890 1308 -2643 1342
rect -2892 1304 -2643 1308
rect -3243 1269 -2643 1304
rect -3243 1235 -2996 1269
rect -2960 1235 -2926 1269
rect -2890 1235 -2643 1269
rect -3243 1135 -2643 1235
rect -2341 11233 -1741 11333
rect -2341 3279 -2094 11233
rect -1988 3279 -1741 11233
rect -2341 3270 -1741 3279
rect -2341 3240 -2092 3270
rect -2341 3206 -2094 3240
rect -2058 3236 -2024 3270
rect -1990 3240 -1741 3270
rect -2060 3206 -2022 3236
rect -1988 3206 -1741 3240
rect -2341 3201 -1741 3206
rect -2341 3167 -2092 3201
rect -2058 3167 -2024 3201
rect -1990 3167 -1741 3201
rect -2341 3133 -2094 3167
rect -2060 3133 -2022 3167
rect -1988 3133 -1741 3167
rect -2341 3132 -1741 3133
rect -2341 3098 -2092 3132
rect -2058 3098 -2024 3132
rect -1990 3098 -1741 3132
rect -2341 3094 -1741 3098
rect -2341 3060 -2094 3094
rect -2060 3063 -2022 3094
rect -2341 3029 -2092 3060
rect -2058 3029 -2024 3063
rect -1988 3060 -1741 3094
rect -1990 3029 -1741 3060
rect -2341 3021 -1741 3029
rect -2341 2987 -2094 3021
rect -2060 2994 -2022 3021
rect -2341 2960 -2092 2987
rect -2058 2960 -2024 2994
rect -1988 2987 -1741 3021
rect -1990 2960 -1741 2987
rect -2341 2948 -1741 2960
rect -2341 2914 -2094 2948
rect -2060 2925 -2022 2948
rect -2341 2891 -2092 2914
rect -2058 2891 -2024 2925
rect -1988 2914 -1741 2948
rect -1990 2891 -1741 2914
rect -2341 2875 -1741 2891
rect -2341 2841 -2094 2875
rect -2060 2856 -2022 2875
rect -2341 2822 -2092 2841
rect -2058 2822 -2024 2856
rect -1988 2841 -1741 2875
rect -1990 2822 -1741 2841
rect -2341 2802 -1741 2822
rect -2341 2768 -2094 2802
rect -2060 2787 -2022 2802
rect -2341 2753 -2092 2768
rect -2058 2753 -2024 2787
rect -1988 2768 -1741 2802
rect -1990 2753 -1741 2768
rect -2341 2729 -1741 2753
rect -2341 2695 -2094 2729
rect -2060 2718 -2022 2729
rect -2341 2684 -2092 2695
rect -2058 2684 -2024 2718
rect -1988 2695 -1741 2729
rect -1990 2684 -1741 2695
rect -2341 2656 -1741 2684
rect -2341 2622 -2094 2656
rect -2060 2649 -2022 2656
rect -2341 2615 -2092 2622
rect -2058 2615 -2024 2649
rect -1988 2622 -1741 2656
rect -1990 2615 -1741 2622
rect -2341 2583 -1741 2615
rect -2341 2549 -2094 2583
rect -2060 2580 -2022 2583
rect -2341 2546 -2092 2549
rect -2058 2546 -2024 2580
rect -1988 2549 -1741 2583
rect -1990 2546 -1741 2549
rect -2341 2511 -1741 2546
rect -2341 2510 -2092 2511
rect -2341 2476 -2094 2510
rect -2058 2477 -2024 2511
rect -1990 2510 -1741 2511
rect -2060 2476 -2022 2477
rect -1988 2476 -1741 2510
rect -2341 2442 -1741 2476
rect -2341 2437 -2092 2442
rect -2341 2403 -2094 2437
rect -2058 2408 -2024 2442
rect -1990 2437 -1741 2442
rect -2060 2403 -2022 2408
rect -1988 2403 -1741 2437
rect -2341 2373 -1741 2403
rect -2341 2364 -2092 2373
rect -2341 2330 -2094 2364
rect -2058 2339 -2024 2373
rect -1990 2364 -1741 2373
rect -2060 2330 -2022 2339
rect -1988 2330 -1741 2364
rect -2341 2304 -1741 2330
rect -2341 2291 -2092 2304
rect -2341 2257 -2094 2291
rect -2058 2270 -2024 2304
rect -1990 2291 -1741 2304
rect -2060 2257 -2022 2270
rect -1988 2257 -1741 2291
rect -2341 2235 -1741 2257
rect -2341 2218 -2092 2235
rect -2341 2184 -2094 2218
rect -2058 2201 -2024 2235
rect -1990 2218 -1741 2235
rect -2060 2184 -2022 2201
rect -1988 2184 -1741 2218
rect -2341 2166 -1741 2184
rect -2341 2145 -2092 2166
rect -2341 2111 -2094 2145
rect -2058 2132 -2024 2166
rect -1990 2145 -1741 2166
rect -2060 2111 -2022 2132
rect -1988 2111 -1741 2145
rect -2341 2097 -1741 2111
rect -2341 2072 -2092 2097
rect -2341 2038 -2094 2072
rect -2058 2063 -2024 2097
rect -1990 2072 -1741 2097
rect -2060 2038 -2022 2063
rect -1988 2038 -1741 2072
rect -2341 2028 -1741 2038
rect -2341 1999 -2092 2028
rect -2341 1965 -2094 1999
rect -2058 1994 -2024 2028
rect -1990 1999 -1741 2028
rect -2060 1965 -2022 1994
rect -1988 1965 -1741 1999
rect -2341 1959 -1741 1965
rect -2341 1926 -2092 1959
rect -2341 1892 -2094 1926
rect -2058 1925 -2024 1959
rect -1990 1926 -1741 1959
rect -2060 1892 -2022 1925
rect -1988 1892 -1741 1926
rect -2341 1890 -1741 1892
rect -2341 1856 -2092 1890
rect -2058 1856 -2024 1890
rect -1990 1856 -1741 1890
rect -2341 1853 -1741 1856
rect -2341 1819 -2094 1853
rect -2060 1821 -2022 1853
rect -2341 1787 -2092 1819
rect -2058 1787 -2024 1821
rect -1988 1819 -1741 1853
rect -1990 1787 -1741 1819
rect -2341 1780 -1741 1787
rect -2341 1746 -2094 1780
rect -2060 1752 -2022 1780
rect -2341 1718 -2092 1746
rect -2058 1718 -2024 1752
rect -1988 1746 -1741 1780
rect -1990 1718 -1741 1746
rect -2341 1707 -1741 1718
rect -2341 1673 -2094 1707
rect -2060 1683 -2022 1707
rect -2341 1649 -2092 1673
rect -2058 1649 -2024 1683
rect -1988 1673 -1741 1707
rect -1990 1649 -1741 1673
rect -2341 1634 -1741 1649
rect -2341 1600 -2094 1634
rect -2060 1614 -2022 1634
rect -2341 1580 -2092 1600
rect -2058 1580 -2024 1614
rect -1988 1600 -1741 1634
rect -1990 1580 -1741 1600
rect -2341 1561 -1741 1580
rect -2341 1527 -2094 1561
rect -2060 1545 -2022 1561
rect -2341 1511 -2092 1527
rect -2058 1511 -2024 1545
rect -1988 1527 -1741 1561
rect -1990 1511 -1741 1527
rect -2341 1488 -1741 1511
rect -2341 1454 -2094 1488
rect -2060 1476 -2022 1488
rect -2341 1442 -2092 1454
rect -2058 1442 -2024 1476
rect -1988 1454 -1741 1488
rect -1990 1442 -1741 1454
rect -2341 1415 -1741 1442
rect -2341 1381 -2094 1415
rect -2060 1407 -2022 1415
rect -2341 1373 -2092 1381
rect -2058 1373 -2024 1407
rect -1988 1381 -1741 1415
rect -1990 1373 -1741 1381
rect -2341 1342 -1741 1373
rect -2341 1308 -2094 1342
rect -2060 1338 -2022 1342
rect -2341 1304 -2092 1308
rect -2058 1304 -2024 1338
rect -1988 1308 -1741 1342
rect -1990 1304 -1741 1308
rect -2341 1269 -1741 1304
rect -2341 1235 -2094 1269
rect -2058 1235 -2024 1269
rect -1988 1235 -1741 1269
rect -2341 1135 -1741 1235
rect -1439 11233 -839 11333
rect -1439 3279 -1192 11233
rect -1086 3279 -839 11233
rect -1439 3270 -839 3279
rect -1439 3240 -1190 3270
rect -1439 3206 -1192 3240
rect -1156 3236 -1122 3270
rect -1088 3240 -839 3270
rect -1158 3206 -1120 3236
rect -1086 3206 -839 3240
rect -1439 3201 -839 3206
rect -1439 3167 -1190 3201
rect -1156 3167 -1122 3201
rect -1088 3167 -839 3201
rect -1439 3133 -1192 3167
rect -1158 3133 -1120 3167
rect -1086 3133 -839 3167
rect -1439 3132 -839 3133
rect -1439 3098 -1190 3132
rect -1156 3098 -1122 3132
rect -1088 3098 -839 3132
rect -1439 3094 -839 3098
rect -1439 3060 -1192 3094
rect -1158 3063 -1120 3094
rect -1439 3029 -1190 3060
rect -1156 3029 -1122 3063
rect -1086 3060 -839 3094
rect -1088 3029 -839 3060
rect -1439 3021 -839 3029
rect -1439 2987 -1192 3021
rect -1158 2994 -1120 3021
rect -1439 2960 -1190 2987
rect -1156 2960 -1122 2994
rect -1086 2987 -839 3021
rect -1088 2960 -839 2987
rect -1439 2948 -839 2960
rect -1439 2914 -1192 2948
rect -1158 2925 -1120 2948
rect -1439 2891 -1190 2914
rect -1156 2891 -1122 2925
rect -1086 2914 -839 2948
rect -1088 2891 -839 2914
rect -1439 2875 -839 2891
rect -1439 2841 -1192 2875
rect -1158 2856 -1120 2875
rect -1439 2822 -1190 2841
rect -1156 2822 -1122 2856
rect -1086 2841 -839 2875
rect -1088 2822 -839 2841
rect -1439 2802 -839 2822
rect -1439 2768 -1192 2802
rect -1158 2787 -1120 2802
rect -1439 2753 -1190 2768
rect -1156 2753 -1122 2787
rect -1086 2768 -839 2802
rect -1088 2753 -839 2768
rect -1439 2729 -839 2753
rect -1439 2695 -1192 2729
rect -1158 2718 -1120 2729
rect -1439 2684 -1190 2695
rect -1156 2684 -1122 2718
rect -1086 2695 -839 2729
rect -1088 2684 -839 2695
rect -1439 2656 -839 2684
rect -1439 2622 -1192 2656
rect -1158 2649 -1120 2656
rect -1439 2615 -1190 2622
rect -1156 2615 -1122 2649
rect -1086 2622 -839 2656
rect -1088 2615 -839 2622
rect -1439 2583 -839 2615
rect -1439 2549 -1192 2583
rect -1158 2580 -1120 2583
rect -1439 2546 -1190 2549
rect -1156 2546 -1122 2580
rect -1086 2549 -839 2583
rect -1088 2546 -839 2549
rect -1439 2511 -839 2546
rect -1439 2510 -1190 2511
rect -1439 2476 -1192 2510
rect -1156 2477 -1122 2511
rect -1088 2510 -839 2511
rect -1158 2476 -1120 2477
rect -1086 2476 -839 2510
rect -1439 2442 -839 2476
rect -1439 2437 -1190 2442
rect -1439 2403 -1192 2437
rect -1156 2408 -1122 2442
rect -1088 2437 -839 2442
rect -1158 2403 -1120 2408
rect -1086 2403 -839 2437
rect -1439 2373 -839 2403
rect -1439 2364 -1190 2373
rect -1439 2330 -1192 2364
rect -1156 2339 -1122 2373
rect -1088 2364 -839 2373
rect -1158 2330 -1120 2339
rect -1086 2330 -839 2364
rect -1439 2304 -839 2330
rect -1439 2291 -1190 2304
rect -1439 2257 -1192 2291
rect -1156 2270 -1122 2304
rect -1088 2291 -839 2304
rect -1158 2257 -1120 2270
rect -1086 2257 -839 2291
rect -1439 2235 -839 2257
rect -1439 2218 -1190 2235
rect -1439 2184 -1192 2218
rect -1156 2201 -1122 2235
rect -1088 2218 -839 2235
rect -1158 2184 -1120 2201
rect -1086 2184 -839 2218
rect -1439 2166 -839 2184
rect -1439 2145 -1190 2166
rect -1439 2111 -1192 2145
rect -1156 2132 -1122 2166
rect -1088 2145 -839 2166
rect -1158 2111 -1120 2132
rect -1086 2111 -839 2145
rect -1439 2097 -839 2111
rect -1439 2072 -1190 2097
rect -1439 2038 -1192 2072
rect -1156 2063 -1122 2097
rect -1088 2072 -839 2097
rect -1158 2038 -1120 2063
rect -1086 2038 -839 2072
rect -1439 2028 -839 2038
rect -1439 1999 -1190 2028
rect -1439 1965 -1192 1999
rect -1156 1994 -1122 2028
rect -1088 1999 -839 2028
rect -1158 1965 -1120 1994
rect -1086 1965 -839 1999
rect -1439 1959 -839 1965
rect -1439 1926 -1190 1959
rect -1439 1892 -1192 1926
rect -1156 1925 -1122 1959
rect -1088 1926 -839 1959
rect -1158 1892 -1120 1925
rect -1086 1892 -839 1926
rect -1439 1890 -839 1892
rect -1439 1856 -1190 1890
rect -1156 1856 -1122 1890
rect -1088 1856 -839 1890
rect -1439 1853 -839 1856
rect -1439 1819 -1192 1853
rect -1158 1821 -1120 1853
rect -1439 1787 -1190 1819
rect -1156 1787 -1122 1821
rect -1086 1819 -839 1853
rect -1088 1787 -839 1819
rect -1439 1780 -839 1787
rect -1439 1746 -1192 1780
rect -1158 1752 -1120 1780
rect -1439 1718 -1190 1746
rect -1156 1718 -1122 1752
rect -1086 1746 -839 1780
rect -1088 1718 -839 1746
rect -1439 1707 -839 1718
rect -1439 1673 -1192 1707
rect -1158 1683 -1120 1707
rect -1439 1649 -1190 1673
rect -1156 1649 -1122 1683
rect -1086 1673 -839 1707
rect -1088 1649 -839 1673
rect -1439 1634 -839 1649
rect -1439 1600 -1192 1634
rect -1158 1614 -1120 1634
rect -1439 1580 -1190 1600
rect -1156 1580 -1122 1614
rect -1086 1600 -839 1634
rect -1088 1580 -839 1600
rect -1439 1561 -839 1580
rect -1439 1527 -1192 1561
rect -1158 1545 -1120 1561
rect -1439 1511 -1190 1527
rect -1156 1511 -1122 1545
rect -1086 1527 -839 1561
rect -1088 1511 -839 1527
rect -1439 1488 -839 1511
rect -1439 1454 -1192 1488
rect -1158 1476 -1120 1488
rect -1439 1442 -1190 1454
rect -1156 1442 -1122 1476
rect -1086 1454 -839 1488
rect -1088 1442 -839 1454
rect -1439 1415 -839 1442
rect -1439 1381 -1192 1415
rect -1158 1407 -1120 1415
rect -1439 1373 -1190 1381
rect -1156 1373 -1122 1407
rect -1086 1381 -839 1415
rect -1088 1373 -839 1381
rect -1439 1342 -839 1373
rect -1439 1308 -1192 1342
rect -1158 1338 -1120 1342
rect -1439 1304 -1190 1308
rect -1156 1304 -1122 1338
rect -1086 1308 -839 1342
rect -1088 1304 -839 1308
rect -1439 1269 -839 1304
rect -1439 1235 -1192 1269
rect -1156 1235 -1122 1269
rect -1086 1235 -839 1269
rect -1439 1135 -839 1235
rect -537 11233 63 11333
rect -537 3279 -290 11233
rect -184 3279 63 11233
rect -537 3270 63 3279
rect -537 3240 -288 3270
rect -537 3206 -290 3240
rect -254 3236 -220 3270
rect -186 3240 63 3270
rect -256 3206 -218 3236
rect -184 3206 63 3240
rect -537 3201 63 3206
rect -537 3167 -288 3201
rect -254 3167 -220 3201
rect -186 3167 63 3201
rect -537 3133 -290 3167
rect -256 3133 -218 3167
rect -184 3133 63 3167
rect -537 3132 63 3133
rect -537 3098 -288 3132
rect -254 3098 -220 3132
rect -186 3098 63 3132
rect -537 3094 63 3098
rect -537 3060 -290 3094
rect -256 3063 -218 3094
rect -537 3029 -288 3060
rect -254 3029 -220 3063
rect -184 3060 63 3094
rect -186 3029 63 3060
rect -537 3021 63 3029
rect -537 2987 -290 3021
rect -256 2994 -218 3021
rect -537 2960 -288 2987
rect -254 2960 -220 2994
rect -184 2987 63 3021
rect -186 2960 63 2987
rect -537 2948 63 2960
rect -537 2914 -290 2948
rect -256 2925 -218 2948
rect -537 2891 -288 2914
rect -254 2891 -220 2925
rect -184 2914 63 2948
rect -186 2891 63 2914
rect -537 2875 63 2891
rect -537 2841 -290 2875
rect -256 2856 -218 2875
rect -537 2822 -288 2841
rect -254 2822 -220 2856
rect -184 2841 63 2875
rect -186 2822 63 2841
rect -537 2802 63 2822
rect -537 2768 -290 2802
rect -256 2787 -218 2802
rect -537 2753 -288 2768
rect -254 2753 -220 2787
rect -184 2768 63 2802
rect -186 2753 63 2768
rect -537 2729 63 2753
rect -537 2695 -290 2729
rect -256 2718 -218 2729
rect -537 2684 -288 2695
rect -254 2684 -220 2718
rect -184 2695 63 2729
rect -186 2684 63 2695
rect -537 2656 63 2684
rect -537 2622 -290 2656
rect -256 2649 -218 2656
rect -537 2615 -288 2622
rect -254 2615 -220 2649
rect -184 2622 63 2656
rect -186 2615 63 2622
rect -537 2583 63 2615
rect -537 2549 -290 2583
rect -256 2580 -218 2583
rect -537 2546 -288 2549
rect -254 2546 -220 2580
rect -184 2549 63 2583
rect -186 2546 63 2549
rect -537 2511 63 2546
rect -537 2510 -288 2511
rect -537 2476 -290 2510
rect -254 2477 -220 2511
rect -186 2510 63 2511
rect -256 2476 -218 2477
rect -184 2476 63 2510
rect -537 2442 63 2476
rect -537 2437 -288 2442
rect -537 2403 -290 2437
rect -254 2408 -220 2442
rect -186 2437 63 2442
rect -256 2403 -218 2408
rect -184 2403 63 2437
rect -537 2373 63 2403
rect -537 2364 -288 2373
rect -537 2330 -290 2364
rect -254 2339 -220 2373
rect -186 2364 63 2373
rect -256 2330 -218 2339
rect -184 2330 63 2364
rect -537 2304 63 2330
rect -537 2291 -288 2304
rect -537 2257 -290 2291
rect -254 2270 -220 2304
rect -186 2291 63 2304
rect -256 2257 -218 2270
rect -184 2257 63 2291
rect -537 2235 63 2257
rect -537 2218 -288 2235
rect -537 2184 -290 2218
rect -254 2201 -220 2235
rect -186 2218 63 2235
rect -256 2184 -218 2201
rect -184 2184 63 2218
rect -537 2166 63 2184
rect -537 2145 -288 2166
rect -537 2111 -290 2145
rect -254 2132 -220 2166
rect -186 2145 63 2166
rect -256 2111 -218 2132
rect -184 2111 63 2145
rect -537 2097 63 2111
rect -537 2072 -288 2097
rect -537 2038 -290 2072
rect -254 2063 -220 2097
rect -186 2072 63 2097
rect -256 2038 -218 2063
rect -184 2038 63 2072
rect -537 2028 63 2038
rect -537 1999 -288 2028
rect -537 1965 -290 1999
rect -254 1994 -220 2028
rect -186 1999 63 2028
rect -256 1965 -218 1994
rect -184 1965 63 1999
rect -537 1959 63 1965
rect -537 1926 -288 1959
rect -537 1892 -290 1926
rect -254 1925 -220 1959
rect -186 1926 63 1959
rect -256 1892 -218 1925
rect -184 1892 63 1926
rect -537 1890 63 1892
rect -537 1856 -288 1890
rect -254 1856 -220 1890
rect -186 1856 63 1890
rect -537 1853 63 1856
rect -537 1819 -290 1853
rect -256 1821 -218 1853
rect -537 1787 -288 1819
rect -254 1787 -220 1821
rect -184 1819 63 1853
rect -186 1787 63 1819
rect -537 1780 63 1787
rect -537 1746 -290 1780
rect -256 1752 -218 1780
rect -537 1718 -288 1746
rect -254 1718 -220 1752
rect -184 1746 63 1780
rect -186 1718 63 1746
rect -537 1707 63 1718
rect -537 1673 -290 1707
rect -256 1683 -218 1707
rect -537 1649 -288 1673
rect -254 1649 -220 1683
rect -184 1673 63 1707
rect -186 1649 63 1673
rect -537 1634 63 1649
rect -537 1600 -290 1634
rect -256 1614 -218 1634
rect -537 1580 -288 1600
rect -254 1580 -220 1614
rect -184 1600 63 1634
rect -186 1580 63 1600
rect -537 1561 63 1580
rect -537 1527 -290 1561
rect -256 1545 -218 1561
rect -537 1511 -288 1527
rect -254 1511 -220 1545
rect -184 1527 63 1561
rect -186 1511 63 1527
rect -537 1488 63 1511
rect -537 1454 -290 1488
rect -256 1476 -218 1488
rect -537 1442 -288 1454
rect -254 1442 -220 1476
rect -184 1454 63 1488
rect -186 1442 63 1454
rect -537 1415 63 1442
rect -537 1381 -290 1415
rect -256 1407 -218 1415
rect -537 1373 -288 1381
rect -254 1373 -220 1407
rect -184 1381 63 1415
rect -186 1373 63 1381
rect -537 1342 63 1373
rect -537 1308 -290 1342
rect -256 1338 -218 1342
rect -537 1304 -288 1308
rect -254 1304 -220 1338
rect -184 1308 63 1342
rect -186 1304 63 1308
rect -537 1269 63 1304
rect -537 1235 -290 1269
rect -254 1235 -220 1269
rect -184 1235 63 1269
rect -537 1135 63 1235
rect 365 11233 965 11333
rect 365 3279 612 11233
rect 718 3279 965 11233
rect 365 3270 965 3279
rect 365 3240 614 3270
rect 365 3206 612 3240
rect 648 3236 682 3270
rect 716 3240 965 3270
rect 646 3206 684 3236
rect 718 3206 965 3240
rect 365 3201 965 3206
rect 365 3167 614 3201
rect 648 3167 682 3201
rect 716 3167 965 3201
rect 365 3133 612 3167
rect 646 3133 684 3167
rect 718 3133 965 3167
rect 365 3132 965 3133
rect 365 3098 614 3132
rect 648 3098 682 3132
rect 716 3098 965 3132
rect 365 3094 965 3098
rect 365 3060 612 3094
rect 646 3063 684 3094
rect 365 3029 614 3060
rect 648 3029 682 3063
rect 718 3060 965 3094
rect 716 3029 965 3060
rect 365 3021 965 3029
rect 365 2987 612 3021
rect 646 2994 684 3021
rect 365 2960 614 2987
rect 648 2960 682 2994
rect 718 2987 965 3021
rect 716 2960 965 2987
rect 365 2948 965 2960
rect 365 2914 612 2948
rect 646 2925 684 2948
rect 365 2891 614 2914
rect 648 2891 682 2925
rect 718 2914 965 2948
rect 716 2891 965 2914
rect 365 2875 965 2891
rect 365 2841 612 2875
rect 646 2856 684 2875
rect 365 2822 614 2841
rect 648 2822 682 2856
rect 718 2841 965 2875
rect 716 2822 965 2841
rect 365 2802 965 2822
rect 365 2768 612 2802
rect 646 2787 684 2802
rect 365 2753 614 2768
rect 648 2753 682 2787
rect 718 2768 965 2802
rect 716 2753 965 2768
rect 365 2729 965 2753
rect 365 2695 612 2729
rect 646 2718 684 2729
rect 365 2684 614 2695
rect 648 2684 682 2718
rect 718 2695 965 2729
rect 716 2684 965 2695
rect 365 2656 965 2684
rect 365 2622 612 2656
rect 646 2649 684 2656
rect 365 2615 614 2622
rect 648 2615 682 2649
rect 718 2622 965 2656
rect 716 2615 965 2622
rect 365 2583 965 2615
rect 365 2549 612 2583
rect 646 2580 684 2583
rect 365 2546 614 2549
rect 648 2546 682 2580
rect 718 2549 965 2583
rect 716 2546 965 2549
rect 365 2511 965 2546
rect 365 2510 614 2511
rect 365 2476 612 2510
rect 648 2477 682 2511
rect 716 2510 965 2511
rect 646 2476 684 2477
rect 718 2476 965 2510
rect 365 2442 965 2476
rect 365 2437 614 2442
rect 365 2403 612 2437
rect 648 2408 682 2442
rect 716 2437 965 2442
rect 646 2403 684 2408
rect 718 2403 965 2437
rect 365 2373 965 2403
rect 365 2364 614 2373
rect 365 2330 612 2364
rect 648 2339 682 2373
rect 716 2364 965 2373
rect 646 2330 684 2339
rect 718 2330 965 2364
rect 365 2304 965 2330
rect 365 2291 614 2304
rect 365 2257 612 2291
rect 648 2270 682 2304
rect 716 2291 965 2304
rect 646 2257 684 2270
rect 718 2257 965 2291
rect 365 2235 965 2257
rect 365 2218 614 2235
rect 365 2184 612 2218
rect 648 2201 682 2235
rect 716 2218 965 2235
rect 646 2184 684 2201
rect 718 2184 965 2218
rect 365 2166 965 2184
rect 365 2145 614 2166
rect 365 2111 612 2145
rect 648 2132 682 2166
rect 716 2145 965 2166
rect 646 2111 684 2132
rect 718 2111 965 2145
rect 365 2097 965 2111
rect 365 2072 614 2097
rect 365 2038 612 2072
rect 648 2063 682 2097
rect 716 2072 965 2097
rect 646 2038 684 2063
rect 718 2038 965 2072
rect 365 2028 965 2038
rect 365 1999 614 2028
rect 365 1965 612 1999
rect 648 1994 682 2028
rect 716 1999 965 2028
rect 646 1965 684 1994
rect 718 1965 965 1999
rect 365 1959 965 1965
rect 365 1926 614 1959
rect 365 1892 612 1926
rect 648 1925 682 1959
rect 716 1926 965 1959
rect 646 1892 684 1925
rect 718 1892 965 1926
rect 365 1890 965 1892
rect 365 1856 614 1890
rect 648 1856 682 1890
rect 716 1856 965 1890
rect 365 1853 965 1856
rect 365 1819 612 1853
rect 646 1821 684 1853
rect 365 1787 614 1819
rect 648 1787 682 1821
rect 718 1819 965 1853
rect 716 1787 965 1819
rect 365 1780 965 1787
rect 365 1746 612 1780
rect 646 1752 684 1780
rect 365 1718 614 1746
rect 648 1718 682 1752
rect 718 1746 965 1780
rect 716 1718 965 1746
rect 365 1707 965 1718
rect 365 1673 612 1707
rect 646 1683 684 1707
rect 365 1649 614 1673
rect 648 1649 682 1683
rect 718 1673 965 1707
rect 716 1649 965 1673
rect 365 1634 965 1649
rect 365 1600 612 1634
rect 646 1614 684 1634
rect 365 1580 614 1600
rect 648 1580 682 1614
rect 718 1600 965 1634
rect 716 1580 965 1600
rect 365 1561 965 1580
rect 365 1527 612 1561
rect 646 1545 684 1561
rect 365 1511 614 1527
rect 648 1511 682 1545
rect 718 1527 965 1561
rect 716 1511 965 1527
rect 365 1488 965 1511
rect 365 1454 612 1488
rect 646 1476 684 1488
rect 365 1442 614 1454
rect 648 1442 682 1476
rect 718 1454 965 1488
rect 716 1442 965 1454
rect 365 1415 965 1442
rect 365 1381 612 1415
rect 646 1407 684 1415
rect 365 1373 614 1381
rect 648 1373 682 1407
rect 718 1381 965 1415
rect 716 1373 965 1381
rect 365 1342 965 1373
rect 365 1308 612 1342
rect 646 1338 684 1342
rect 365 1304 614 1308
rect 648 1304 682 1338
rect 718 1308 965 1342
rect 716 1304 965 1308
rect 365 1269 965 1304
rect 365 1235 612 1269
rect 648 1235 682 1269
rect 718 1235 965 1269
rect 365 1135 965 1235
rect 1267 11233 1867 11333
rect 1267 3279 1514 11233
rect 1620 3279 1867 11233
rect 1267 3270 1867 3279
rect 1267 3240 1516 3270
rect 1267 3206 1514 3240
rect 1550 3236 1584 3270
rect 1618 3240 1867 3270
rect 1548 3206 1586 3236
rect 1620 3206 1867 3240
rect 1267 3201 1867 3206
rect 1267 3167 1516 3201
rect 1550 3167 1584 3201
rect 1618 3167 1867 3201
rect 1267 3133 1514 3167
rect 1548 3133 1586 3167
rect 1620 3133 1867 3167
rect 1267 3132 1867 3133
rect 1267 3098 1516 3132
rect 1550 3098 1584 3132
rect 1618 3098 1867 3132
rect 1267 3094 1867 3098
rect 1267 3060 1514 3094
rect 1548 3063 1586 3094
rect 1267 3029 1516 3060
rect 1550 3029 1584 3063
rect 1620 3060 1867 3094
rect 1618 3029 1867 3060
rect 1267 3021 1867 3029
rect 1267 2987 1514 3021
rect 1548 2994 1586 3021
rect 1267 2960 1516 2987
rect 1550 2960 1584 2994
rect 1620 2987 1867 3021
rect 1618 2960 1867 2987
rect 1267 2948 1867 2960
rect 1267 2914 1514 2948
rect 1548 2925 1586 2948
rect 1267 2891 1516 2914
rect 1550 2891 1584 2925
rect 1620 2914 1867 2948
rect 1618 2891 1867 2914
rect 1267 2875 1867 2891
rect 1267 2841 1514 2875
rect 1548 2856 1586 2875
rect 1267 2822 1516 2841
rect 1550 2822 1584 2856
rect 1620 2841 1867 2875
rect 1618 2822 1867 2841
rect 1267 2802 1867 2822
rect 1267 2768 1514 2802
rect 1548 2787 1586 2802
rect 1267 2753 1516 2768
rect 1550 2753 1584 2787
rect 1620 2768 1867 2802
rect 1618 2753 1867 2768
rect 1267 2729 1867 2753
rect 1267 2695 1514 2729
rect 1548 2718 1586 2729
rect 1267 2684 1516 2695
rect 1550 2684 1584 2718
rect 1620 2695 1867 2729
rect 1618 2684 1867 2695
rect 1267 2656 1867 2684
rect 1267 2622 1514 2656
rect 1548 2649 1586 2656
rect 1267 2615 1516 2622
rect 1550 2615 1584 2649
rect 1620 2622 1867 2656
rect 1618 2615 1867 2622
rect 1267 2583 1867 2615
rect 1267 2549 1514 2583
rect 1548 2580 1586 2583
rect 1267 2546 1516 2549
rect 1550 2546 1584 2580
rect 1620 2549 1867 2583
rect 1618 2546 1867 2549
rect 1267 2511 1867 2546
rect 1267 2510 1516 2511
rect 1267 2476 1514 2510
rect 1550 2477 1584 2511
rect 1618 2510 1867 2511
rect 1548 2476 1586 2477
rect 1620 2476 1867 2510
rect 1267 2442 1867 2476
rect 1267 2437 1516 2442
rect 1267 2403 1514 2437
rect 1550 2408 1584 2442
rect 1618 2437 1867 2442
rect 1548 2403 1586 2408
rect 1620 2403 1867 2437
rect 1267 2373 1867 2403
rect 1267 2364 1516 2373
rect 1267 2330 1514 2364
rect 1550 2339 1584 2373
rect 1618 2364 1867 2373
rect 1548 2330 1586 2339
rect 1620 2330 1867 2364
rect 1267 2304 1867 2330
rect 1267 2291 1516 2304
rect 1267 2257 1514 2291
rect 1550 2270 1584 2304
rect 1618 2291 1867 2304
rect 1548 2257 1586 2270
rect 1620 2257 1867 2291
rect 1267 2235 1867 2257
rect 1267 2218 1516 2235
rect 1267 2184 1514 2218
rect 1550 2201 1584 2235
rect 1618 2218 1867 2235
rect 1548 2184 1586 2201
rect 1620 2184 1867 2218
rect 1267 2166 1867 2184
rect 1267 2145 1516 2166
rect 1267 2111 1514 2145
rect 1550 2132 1584 2166
rect 1618 2145 1867 2166
rect 1548 2111 1586 2132
rect 1620 2111 1867 2145
rect 1267 2097 1867 2111
rect 1267 2072 1516 2097
rect 1267 2038 1514 2072
rect 1550 2063 1584 2097
rect 1618 2072 1867 2097
rect 1548 2038 1586 2063
rect 1620 2038 1867 2072
rect 1267 2028 1867 2038
rect 1267 1999 1516 2028
rect 1267 1965 1514 1999
rect 1550 1994 1584 2028
rect 1618 1999 1867 2028
rect 1548 1965 1586 1994
rect 1620 1965 1867 1999
rect 1267 1959 1867 1965
rect 1267 1926 1516 1959
rect 1267 1892 1514 1926
rect 1550 1925 1584 1959
rect 1618 1926 1867 1959
rect 1548 1892 1586 1925
rect 1620 1892 1867 1926
rect 1267 1890 1867 1892
rect 1267 1856 1516 1890
rect 1550 1856 1584 1890
rect 1618 1856 1867 1890
rect 1267 1853 1867 1856
rect 1267 1819 1514 1853
rect 1548 1821 1586 1853
rect 1267 1787 1516 1819
rect 1550 1787 1584 1821
rect 1620 1819 1867 1853
rect 1618 1787 1867 1819
rect 1267 1780 1867 1787
rect 1267 1746 1514 1780
rect 1548 1752 1586 1780
rect 1267 1718 1516 1746
rect 1550 1718 1584 1752
rect 1620 1746 1867 1780
rect 1618 1718 1867 1746
rect 1267 1707 1867 1718
rect 1267 1673 1514 1707
rect 1548 1683 1586 1707
rect 1267 1649 1516 1673
rect 1550 1649 1584 1683
rect 1620 1673 1867 1707
rect 1618 1649 1867 1673
rect 1267 1634 1867 1649
rect 1267 1600 1514 1634
rect 1548 1614 1586 1634
rect 1267 1580 1516 1600
rect 1550 1580 1584 1614
rect 1620 1600 1867 1634
rect 1618 1580 1867 1600
rect 1267 1561 1867 1580
rect 1267 1527 1514 1561
rect 1548 1545 1586 1561
rect 1267 1511 1516 1527
rect 1550 1511 1584 1545
rect 1620 1527 1867 1561
rect 1618 1511 1867 1527
rect 1267 1488 1867 1511
rect 1267 1454 1514 1488
rect 1548 1476 1586 1488
rect 1267 1442 1516 1454
rect 1550 1442 1584 1476
rect 1620 1454 1867 1488
rect 1618 1442 1867 1454
rect 1267 1415 1867 1442
rect 1267 1381 1514 1415
rect 1548 1407 1586 1415
rect 1267 1373 1516 1381
rect 1550 1373 1584 1407
rect 1620 1381 1867 1415
rect 1618 1373 1867 1381
rect 1267 1342 1867 1373
rect 1267 1308 1514 1342
rect 1548 1338 1586 1342
rect 1267 1304 1516 1308
rect 1550 1304 1584 1338
rect 1620 1308 1867 1342
rect 1618 1304 1867 1308
rect 1267 1269 1867 1304
rect 1267 1235 1514 1269
rect 1550 1235 1584 1269
rect 1620 1235 1867 1269
rect 1267 1135 1867 1235
rect 2169 11233 2769 11333
rect 2169 3279 2416 11233
rect 2522 3279 2769 11233
rect 2169 3270 2769 3279
rect 2169 3240 2418 3270
rect 2169 3206 2416 3240
rect 2452 3236 2486 3270
rect 2520 3240 2769 3270
rect 2450 3206 2488 3236
rect 2522 3206 2769 3240
rect 2169 3201 2769 3206
rect 2169 3167 2418 3201
rect 2452 3167 2486 3201
rect 2520 3167 2769 3201
rect 2169 3133 2416 3167
rect 2450 3133 2488 3167
rect 2522 3133 2769 3167
rect 2169 3132 2769 3133
rect 2169 3098 2418 3132
rect 2452 3098 2486 3132
rect 2520 3098 2769 3132
rect 2169 3094 2769 3098
rect 2169 3060 2416 3094
rect 2450 3063 2488 3094
rect 2169 3029 2418 3060
rect 2452 3029 2486 3063
rect 2522 3060 2769 3094
rect 2520 3029 2769 3060
rect 2169 3021 2769 3029
rect 2169 2987 2416 3021
rect 2450 2994 2488 3021
rect 2169 2960 2418 2987
rect 2452 2960 2486 2994
rect 2522 2987 2769 3021
rect 2520 2960 2769 2987
rect 2169 2948 2769 2960
rect 2169 2914 2416 2948
rect 2450 2925 2488 2948
rect 2169 2891 2418 2914
rect 2452 2891 2486 2925
rect 2522 2914 2769 2948
rect 2520 2891 2769 2914
rect 2169 2875 2769 2891
rect 2169 2841 2416 2875
rect 2450 2856 2488 2875
rect 2169 2822 2418 2841
rect 2452 2822 2486 2856
rect 2522 2841 2769 2875
rect 2520 2822 2769 2841
rect 2169 2802 2769 2822
rect 2169 2768 2416 2802
rect 2450 2787 2488 2802
rect 2169 2753 2418 2768
rect 2452 2753 2486 2787
rect 2522 2768 2769 2802
rect 2520 2753 2769 2768
rect 2169 2729 2769 2753
rect 2169 2695 2416 2729
rect 2450 2718 2488 2729
rect 2169 2684 2418 2695
rect 2452 2684 2486 2718
rect 2522 2695 2769 2729
rect 2520 2684 2769 2695
rect 2169 2656 2769 2684
rect 2169 2622 2416 2656
rect 2450 2649 2488 2656
rect 2169 2615 2418 2622
rect 2452 2615 2486 2649
rect 2522 2622 2769 2656
rect 2520 2615 2769 2622
rect 2169 2583 2769 2615
rect 2169 2549 2416 2583
rect 2450 2580 2488 2583
rect 2169 2546 2418 2549
rect 2452 2546 2486 2580
rect 2522 2549 2769 2583
rect 2520 2546 2769 2549
rect 2169 2511 2769 2546
rect 2169 2510 2418 2511
rect 2169 2476 2416 2510
rect 2452 2477 2486 2511
rect 2520 2510 2769 2511
rect 2450 2476 2488 2477
rect 2522 2476 2769 2510
rect 2169 2442 2769 2476
rect 2169 2437 2418 2442
rect 2169 2403 2416 2437
rect 2452 2408 2486 2442
rect 2520 2437 2769 2442
rect 2450 2403 2488 2408
rect 2522 2403 2769 2437
rect 2169 2373 2769 2403
rect 2169 2364 2418 2373
rect 2169 2330 2416 2364
rect 2452 2339 2486 2373
rect 2520 2364 2769 2373
rect 2450 2330 2488 2339
rect 2522 2330 2769 2364
rect 2169 2304 2769 2330
rect 2169 2291 2418 2304
rect 2169 2257 2416 2291
rect 2452 2270 2486 2304
rect 2520 2291 2769 2304
rect 2450 2257 2488 2270
rect 2522 2257 2769 2291
rect 2169 2235 2769 2257
rect 2169 2218 2418 2235
rect 2169 2184 2416 2218
rect 2452 2201 2486 2235
rect 2520 2218 2769 2235
rect 2450 2184 2488 2201
rect 2522 2184 2769 2218
rect 2169 2166 2769 2184
rect 2169 2145 2418 2166
rect 2169 2111 2416 2145
rect 2452 2132 2486 2166
rect 2520 2145 2769 2166
rect 2450 2111 2488 2132
rect 2522 2111 2769 2145
rect 2169 2097 2769 2111
rect 2169 2072 2418 2097
rect 2169 2038 2416 2072
rect 2452 2063 2486 2097
rect 2520 2072 2769 2097
rect 2450 2038 2488 2063
rect 2522 2038 2769 2072
rect 2169 2028 2769 2038
rect 2169 1999 2418 2028
rect 2169 1965 2416 1999
rect 2452 1994 2486 2028
rect 2520 1999 2769 2028
rect 2450 1965 2488 1994
rect 2522 1965 2769 1999
rect 2169 1959 2769 1965
rect 2169 1926 2418 1959
rect 2169 1892 2416 1926
rect 2452 1925 2486 1959
rect 2520 1926 2769 1959
rect 2450 1892 2488 1925
rect 2522 1892 2769 1926
rect 2169 1890 2769 1892
rect 2169 1856 2418 1890
rect 2452 1856 2486 1890
rect 2520 1856 2769 1890
rect 2169 1853 2769 1856
rect 2169 1819 2416 1853
rect 2450 1821 2488 1853
rect 2169 1787 2418 1819
rect 2452 1787 2486 1821
rect 2522 1819 2769 1853
rect 2520 1787 2769 1819
rect 2169 1780 2769 1787
rect 2169 1746 2416 1780
rect 2450 1752 2488 1780
rect 2169 1718 2418 1746
rect 2452 1718 2486 1752
rect 2522 1746 2769 1780
rect 2520 1718 2769 1746
rect 2169 1707 2769 1718
rect 2169 1673 2416 1707
rect 2450 1683 2488 1707
rect 2169 1649 2418 1673
rect 2452 1649 2486 1683
rect 2522 1673 2769 1707
rect 2520 1649 2769 1673
rect 2169 1634 2769 1649
rect 2169 1600 2416 1634
rect 2450 1614 2488 1634
rect 2169 1580 2418 1600
rect 2452 1580 2486 1614
rect 2522 1600 2769 1634
rect 2520 1580 2769 1600
rect 2169 1561 2769 1580
rect 2169 1527 2416 1561
rect 2450 1545 2488 1561
rect 2169 1511 2418 1527
rect 2452 1511 2486 1545
rect 2522 1527 2769 1561
rect 2520 1511 2769 1527
rect 2169 1488 2769 1511
rect 2169 1454 2416 1488
rect 2450 1476 2488 1488
rect 2169 1442 2418 1454
rect 2452 1442 2486 1476
rect 2522 1454 2769 1488
rect 2520 1442 2769 1454
rect 2169 1415 2769 1442
rect 2169 1381 2416 1415
rect 2450 1407 2488 1415
rect 2169 1373 2418 1381
rect 2452 1373 2486 1407
rect 2522 1381 2769 1415
rect 2520 1373 2769 1381
rect 2169 1342 2769 1373
rect 2169 1308 2416 1342
rect 2450 1338 2488 1342
rect 2169 1304 2418 1308
rect 2452 1304 2486 1338
rect 2522 1308 2769 1342
rect 2520 1304 2769 1308
rect 2169 1269 2769 1304
rect 2169 1235 2416 1269
rect 2452 1235 2486 1269
rect 2522 1235 2769 1269
rect 2169 1135 2769 1235
rect 3071 11233 3671 11333
rect 3071 3279 3318 11233
rect 3424 3279 3671 11233
rect 3071 3270 3671 3279
rect 3071 3240 3320 3270
rect 3071 3206 3318 3240
rect 3354 3236 3388 3270
rect 3422 3240 3671 3270
rect 3352 3206 3390 3236
rect 3424 3206 3671 3240
rect 3071 3201 3671 3206
rect 3071 3167 3320 3201
rect 3354 3167 3388 3201
rect 3422 3167 3671 3201
rect 3071 3133 3318 3167
rect 3352 3133 3390 3167
rect 3424 3133 3671 3167
rect 3071 3132 3671 3133
rect 3071 3098 3320 3132
rect 3354 3098 3388 3132
rect 3422 3098 3671 3132
rect 3071 3094 3671 3098
rect 3071 3060 3318 3094
rect 3352 3063 3390 3094
rect 3071 3029 3320 3060
rect 3354 3029 3388 3063
rect 3424 3060 3671 3094
rect 3422 3029 3671 3060
rect 3071 3021 3671 3029
rect 3071 2987 3318 3021
rect 3352 2994 3390 3021
rect 3071 2960 3320 2987
rect 3354 2960 3388 2994
rect 3424 2987 3671 3021
rect 3422 2960 3671 2987
rect 3071 2948 3671 2960
rect 3071 2914 3318 2948
rect 3352 2925 3390 2948
rect 3071 2891 3320 2914
rect 3354 2891 3388 2925
rect 3424 2914 3671 2948
rect 3422 2891 3671 2914
rect 3071 2875 3671 2891
rect 3071 2841 3318 2875
rect 3352 2856 3390 2875
rect 3071 2822 3320 2841
rect 3354 2822 3388 2856
rect 3424 2841 3671 2875
rect 3422 2822 3671 2841
rect 3071 2802 3671 2822
rect 3071 2768 3318 2802
rect 3352 2787 3390 2802
rect 3071 2753 3320 2768
rect 3354 2753 3388 2787
rect 3424 2768 3671 2802
rect 3422 2753 3671 2768
rect 3071 2729 3671 2753
rect 3071 2695 3318 2729
rect 3352 2718 3390 2729
rect 3071 2684 3320 2695
rect 3354 2684 3388 2718
rect 3424 2695 3671 2729
rect 3422 2684 3671 2695
rect 3071 2656 3671 2684
rect 3071 2622 3318 2656
rect 3352 2649 3390 2656
rect 3071 2615 3320 2622
rect 3354 2615 3388 2649
rect 3424 2622 3671 2656
rect 3422 2615 3671 2622
rect 3071 2583 3671 2615
rect 3071 2549 3318 2583
rect 3352 2580 3390 2583
rect 3071 2546 3320 2549
rect 3354 2546 3388 2580
rect 3424 2549 3671 2583
rect 3422 2546 3671 2549
rect 3071 2511 3671 2546
rect 3071 2510 3320 2511
rect 3071 2476 3318 2510
rect 3354 2477 3388 2511
rect 3422 2510 3671 2511
rect 3352 2476 3390 2477
rect 3424 2476 3671 2510
rect 3071 2442 3671 2476
rect 3071 2437 3320 2442
rect 3071 2403 3318 2437
rect 3354 2408 3388 2442
rect 3422 2437 3671 2442
rect 3352 2403 3390 2408
rect 3424 2403 3671 2437
rect 3071 2373 3671 2403
rect 3071 2364 3320 2373
rect 3071 2330 3318 2364
rect 3354 2339 3388 2373
rect 3422 2364 3671 2373
rect 3352 2330 3390 2339
rect 3424 2330 3671 2364
rect 3071 2304 3671 2330
rect 3071 2291 3320 2304
rect 3071 2257 3318 2291
rect 3354 2270 3388 2304
rect 3422 2291 3671 2304
rect 3352 2257 3390 2270
rect 3424 2257 3671 2291
rect 3071 2235 3671 2257
rect 3071 2218 3320 2235
rect 3071 2184 3318 2218
rect 3354 2201 3388 2235
rect 3422 2218 3671 2235
rect 3352 2184 3390 2201
rect 3424 2184 3671 2218
rect 3071 2166 3671 2184
rect 3071 2145 3320 2166
rect 3071 2111 3318 2145
rect 3354 2132 3388 2166
rect 3422 2145 3671 2166
rect 3352 2111 3390 2132
rect 3424 2111 3671 2145
rect 3071 2097 3671 2111
rect 3071 2072 3320 2097
rect 3071 2038 3318 2072
rect 3354 2063 3388 2097
rect 3422 2072 3671 2097
rect 3352 2038 3390 2063
rect 3424 2038 3671 2072
rect 3071 2028 3671 2038
rect 3071 1999 3320 2028
rect 3071 1965 3318 1999
rect 3354 1994 3388 2028
rect 3422 1999 3671 2028
rect 3352 1965 3390 1994
rect 3424 1965 3671 1999
rect 3071 1959 3671 1965
rect 3071 1926 3320 1959
rect 3071 1892 3318 1926
rect 3354 1925 3388 1959
rect 3422 1926 3671 1959
rect 3352 1892 3390 1925
rect 3424 1892 3671 1926
rect 3071 1890 3671 1892
rect 3071 1856 3320 1890
rect 3354 1856 3388 1890
rect 3422 1856 3671 1890
rect 3071 1853 3671 1856
rect 3071 1819 3318 1853
rect 3352 1821 3390 1853
rect 3071 1787 3320 1819
rect 3354 1787 3388 1821
rect 3424 1819 3671 1853
rect 3422 1787 3671 1819
rect 3071 1780 3671 1787
rect 3071 1746 3318 1780
rect 3352 1752 3390 1780
rect 3071 1718 3320 1746
rect 3354 1718 3388 1752
rect 3424 1746 3671 1780
rect 3422 1718 3671 1746
rect 3071 1707 3671 1718
rect 3071 1673 3318 1707
rect 3352 1683 3390 1707
rect 3071 1649 3320 1673
rect 3354 1649 3388 1683
rect 3424 1673 3671 1707
rect 3422 1649 3671 1673
rect 3071 1634 3671 1649
rect 3071 1600 3318 1634
rect 3352 1614 3390 1634
rect 3071 1580 3320 1600
rect 3354 1580 3388 1614
rect 3424 1600 3671 1634
rect 3422 1580 3671 1600
rect 3071 1561 3671 1580
rect 3071 1527 3318 1561
rect 3352 1545 3390 1561
rect 3071 1511 3320 1527
rect 3354 1511 3388 1545
rect 3424 1527 3671 1561
rect 3422 1511 3671 1527
rect 3071 1488 3671 1511
rect 3071 1454 3318 1488
rect 3352 1476 3390 1488
rect 3071 1442 3320 1454
rect 3354 1442 3388 1476
rect 3424 1454 3671 1488
rect 3422 1442 3671 1454
rect 3071 1415 3671 1442
rect 3071 1381 3318 1415
rect 3352 1407 3390 1415
rect 3071 1373 3320 1381
rect 3354 1373 3388 1407
rect 3424 1381 3671 1415
rect 3422 1373 3671 1381
rect 3071 1342 3671 1373
rect 3071 1308 3318 1342
rect 3352 1338 3390 1342
rect 3071 1304 3320 1308
rect 3354 1304 3388 1338
rect 3424 1308 3671 1342
rect 3422 1304 3671 1308
rect 3071 1269 3671 1304
rect 3071 1235 3318 1269
rect 3354 1235 3388 1269
rect 3424 1235 3671 1269
rect 3071 1135 3671 1235
rect 3973 11233 4573 11333
rect 3973 3279 4220 11233
rect 4326 3279 4573 11233
rect 3973 3270 4573 3279
rect 3973 3240 4222 3270
rect 3973 3206 4220 3240
rect 4256 3236 4290 3270
rect 4324 3240 4573 3270
rect 4254 3206 4292 3236
rect 4326 3206 4573 3240
rect 3973 3201 4573 3206
rect 3973 3167 4222 3201
rect 4256 3167 4290 3201
rect 4324 3167 4573 3201
rect 3973 3133 4220 3167
rect 4254 3133 4292 3167
rect 4326 3133 4573 3167
rect 3973 3132 4573 3133
rect 3973 3098 4222 3132
rect 4256 3098 4290 3132
rect 4324 3098 4573 3132
rect 3973 3094 4573 3098
rect 3973 3060 4220 3094
rect 4254 3063 4292 3094
rect 3973 3029 4222 3060
rect 4256 3029 4290 3063
rect 4326 3060 4573 3094
rect 4324 3029 4573 3060
rect 3973 3021 4573 3029
rect 3973 2987 4220 3021
rect 4254 2994 4292 3021
rect 3973 2960 4222 2987
rect 4256 2960 4290 2994
rect 4326 2987 4573 3021
rect 4324 2960 4573 2987
rect 3973 2948 4573 2960
rect 3973 2914 4220 2948
rect 4254 2925 4292 2948
rect 3973 2891 4222 2914
rect 4256 2891 4290 2925
rect 4326 2914 4573 2948
rect 4324 2891 4573 2914
rect 3973 2875 4573 2891
rect 3973 2841 4220 2875
rect 4254 2856 4292 2875
rect 3973 2822 4222 2841
rect 4256 2822 4290 2856
rect 4326 2841 4573 2875
rect 4324 2822 4573 2841
rect 3973 2802 4573 2822
rect 3973 2768 4220 2802
rect 4254 2787 4292 2802
rect 3973 2753 4222 2768
rect 4256 2753 4290 2787
rect 4326 2768 4573 2802
rect 4324 2753 4573 2768
rect 3973 2729 4573 2753
rect 3973 2695 4220 2729
rect 4254 2718 4292 2729
rect 3973 2684 4222 2695
rect 4256 2684 4290 2718
rect 4326 2695 4573 2729
rect 4324 2684 4573 2695
rect 3973 2656 4573 2684
rect 3973 2622 4220 2656
rect 4254 2649 4292 2656
rect 3973 2615 4222 2622
rect 4256 2615 4290 2649
rect 4326 2622 4573 2656
rect 4324 2615 4573 2622
rect 3973 2583 4573 2615
rect 3973 2549 4220 2583
rect 4254 2580 4292 2583
rect 3973 2546 4222 2549
rect 4256 2546 4290 2580
rect 4326 2549 4573 2583
rect 4324 2546 4573 2549
rect 3973 2511 4573 2546
rect 3973 2510 4222 2511
rect 3973 2476 4220 2510
rect 4256 2477 4290 2511
rect 4324 2510 4573 2511
rect 4254 2476 4292 2477
rect 4326 2476 4573 2510
rect 3973 2442 4573 2476
rect 3973 2437 4222 2442
rect 3973 2403 4220 2437
rect 4256 2408 4290 2442
rect 4324 2437 4573 2442
rect 4254 2403 4292 2408
rect 4326 2403 4573 2437
rect 3973 2373 4573 2403
rect 3973 2364 4222 2373
rect 3973 2330 4220 2364
rect 4256 2339 4290 2373
rect 4324 2364 4573 2373
rect 4254 2330 4292 2339
rect 4326 2330 4573 2364
rect 3973 2304 4573 2330
rect 3973 2291 4222 2304
rect 3973 2257 4220 2291
rect 4256 2270 4290 2304
rect 4324 2291 4573 2304
rect 4254 2257 4292 2270
rect 4326 2257 4573 2291
rect 3973 2235 4573 2257
rect 3973 2218 4222 2235
rect 3973 2184 4220 2218
rect 4256 2201 4290 2235
rect 4324 2218 4573 2235
rect 4254 2184 4292 2201
rect 4326 2184 4573 2218
rect 3973 2166 4573 2184
rect 3973 2145 4222 2166
rect 3973 2111 4220 2145
rect 4256 2132 4290 2166
rect 4324 2145 4573 2166
rect 4254 2111 4292 2132
rect 4326 2111 4573 2145
rect 3973 2097 4573 2111
rect 3973 2072 4222 2097
rect 3973 2038 4220 2072
rect 4256 2063 4290 2097
rect 4324 2072 4573 2097
rect 4254 2038 4292 2063
rect 4326 2038 4573 2072
rect 3973 2028 4573 2038
rect 3973 1999 4222 2028
rect 3973 1965 4220 1999
rect 4256 1994 4290 2028
rect 4324 1999 4573 2028
rect 4254 1965 4292 1994
rect 4326 1965 4573 1999
rect 3973 1959 4573 1965
rect 3973 1926 4222 1959
rect 3973 1892 4220 1926
rect 4256 1925 4290 1959
rect 4324 1926 4573 1959
rect 4254 1892 4292 1925
rect 4326 1892 4573 1926
rect 3973 1890 4573 1892
rect 3973 1856 4222 1890
rect 4256 1856 4290 1890
rect 4324 1856 4573 1890
rect 3973 1853 4573 1856
rect 3973 1819 4220 1853
rect 4254 1821 4292 1853
rect 3973 1787 4222 1819
rect 4256 1787 4290 1821
rect 4326 1819 4573 1853
rect 4324 1787 4573 1819
rect 3973 1780 4573 1787
rect 3973 1746 4220 1780
rect 4254 1752 4292 1780
rect 3973 1718 4222 1746
rect 4256 1718 4290 1752
rect 4326 1746 4573 1780
rect 4324 1718 4573 1746
rect 3973 1707 4573 1718
rect 3973 1673 4220 1707
rect 4254 1683 4292 1707
rect 3973 1649 4222 1673
rect 4256 1649 4290 1683
rect 4326 1673 4573 1707
rect 4324 1649 4573 1673
rect 3973 1634 4573 1649
rect 3973 1600 4220 1634
rect 4254 1614 4292 1634
rect 3973 1580 4222 1600
rect 4256 1580 4290 1614
rect 4326 1600 4573 1634
rect 4324 1580 4573 1600
rect 3973 1561 4573 1580
rect 3973 1527 4220 1561
rect 4254 1545 4292 1561
rect 3973 1511 4222 1527
rect 4256 1511 4290 1545
rect 4326 1527 4573 1561
rect 4324 1511 4573 1527
rect 3973 1488 4573 1511
rect 3973 1454 4220 1488
rect 4254 1476 4292 1488
rect 3973 1442 4222 1454
rect 4256 1442 4290 1476
rect 4326 1454 4573 1488
rect 4324 1442 4573 1454
rect 3973 1415 4573 1442
rect 3973 1381 4220 1415
rect 4254 1407 4292 1415
rect 3973 1373 4222 1381
rect 4256 1373 4290 1407
rect 4326 1381 4573 1415
rect 4324 1373 4573 1381
rect 3973 1342 4573 1373
rect 3973 1308 4220 1342
rect 4254 1338 4292 1342
rect 3973 1304 4222 1308
rect 4256 1304 4290 1338
rect 4326 1308 4573 1342
rect 4324 1304 4573 1308
rect 3973 1269 4573 1304
rect 3973 1235 4220 1269
rect 4256 1235 4290 1269
rect 4326 1235 4573 1269
rect 3973 1135 4573 1235
rect 4875 11233 5475 11333
rect 4875 3279 5122 11233
rect 5228 3279 5475 11233
rect 4875 3270 5475 3279
rect 4875 3240 5124 3270
rect 4875 3206 5122 3240
rect 5158 3236 5192 3270
rect 5226 3240 5475 3270
rect 5156 3206 5194 3236
rect 5228 3206 5475 3240
rect 4875 3201 5475 3206
rect 4875 3167 5124 3201
rect 5158 3167 5192 3201
rect 5226 3167 5475 3201
rect 4875 3133 5122 3167
rect 5156 3133 5194 3167
rect 5228 3133 5475 3167
rect 4875 3132 5475 3133
rect 4875 3098 5124 3132
rect 5158 3098 5192 3132
rect 5226 3098 5475 3132
rect 4875 3094 5475 3098
rect 4875 3060 5122 3094
rect 5156 3063 5194 3094
rect 4875 3029 5124 3060
rect 5158 3029 5192 3063
rect 5228 3060 5475 3094
rect 5226 3029 5475 3060
rect 4875 3021 5475 3029
rect 4875 2987 5122 3021
rect 5156 2994 5194 3021
rect 4875 2960 5124 2987
rect 5158 2960 5192 2994
rect 5228 2987 5475 3021
rect 5226 2960 5475 2987
rect 4875 2948 5475 2960
rect 4875 2914 5122 2948
rect 5156 2925 5194 2948
rect 4875 2891 5124 2914
rect 5158 2891 5192 2925
rect 5228 2914 5475 2948
rect 5226 2891 5475 2914
rect 4875 2875 5475 2891
rect 4875 2841 5122 2875
rect 5156 2856 5194 2875
rect 4875 2822 5124 2841
rect 5158 2822 5192 2856
rect 5228 2841 5475 2875
rect 5226 2822 5475 2841
rect 4875 2802 5475 2822
rect 4875 2768 5122 2802
rect 5156 2787 5194 2802
rect 4875 2753 5124 2768
rect 5158 2753 5192 2787
rect 5228 2768 5475 2802
rect 5226 2753 5475 2768
rect 4875 2729 5475 2753
rect 4875 2695 5122 2729
rect 5156 2718 5194 2729
rect 4875 2684 5124 2695
rect 5158 2684 5192 2718
rect 5228 2695 5475 2729
rect 5226 2684 5475 2695
rect 4875 2656 5475 2684
rect 4875 2622 5122 2656
rect 5156 2649 5194 2656
rect 4875 2615 5124 2622
rect 5158 2615 5192 2649
rect 5228 2622 5475 2656
rect 5226 2615 5475 2622
rect 4875 2583 5475 2615
rect 4875 2549 5122 2583
rect 5156 2580 5194 2583
rect 4875 2546 5124 2549
rect 5158 2546 5192 2580
rect 5228 2549 5475 2583
rect 5226 2546 5475 2549
rect 4875 2511 5475 2546
rect 4875 2510 5124 2511
rect 4875 2476 5122 2510
rect 5158 2477 5192 2511
rect 5226 2510 5475 2511
rect 5156 2476 5194 2477
rect 5228 2476 5475 2510
rect 4875 2442 5475 2476
rect 4875 2437 5124 2442
rect 4875 2403 5122 2437
rect 5158 2408 5192 2442
rect 5226 2437 5475 2442
rect 5156 2403 5194 2408
rect 5228 2403 5475 2437
rect 4875 2373 5475 2403
rect 4875 2364 5124 2373
rect 4875 2330 5122 2364
rect 5158 2339 5192 2373
rect 5226 2364 5475 2373
rect 5156 2330 5194 2339
rect 5228 2330 5475 2364
rect 4875 2304 5475 2330
rect 4875 2291 5124 2304
rect 4875 2257 5122 2291
rect 5158 2270 5192 2304
rect 5226 2291 5475 2304
rect 5156 2257 5194 2270
rect 5228 2257 5475 2291
rect 4875 2235 5475 2257
rect 4875 2218 5124 2235
rect 4875 2184 5122 2218
rect 5158 2201 5192 2235
rect 5226 2218 5475 2235
rect 5156 2184 5194 2201
rect 5228 2184 5475 2218
rect 4875 2166 5475 2184
rect 4875 2145 5124 2166
rect 4875 2111 5122 2145
rect 5158 2132 5192 2166
rect 5226 2145 5475 2166
rect 5156 2111 5194 2132
rect 5228 2111 5475 2145
rect 4875 2097 5475 2111
rect 4875 2072 5124 2097
rect 4875 2038 5122 2072
rect 5158 2063 5192 2097
rect 5226 2072 5475 2097
rect 5156 2038 5194 2063
rect 5228 2038 5475 2072
rect 4875 2028 5475 2038
rect 4875 1999 5124 2028
rect 4875 1965 5122 1999
rect 5158 1994 5192 2028
rect 5226 1999 5475 2028
rect 5156 1965 5194 1994
rect 5228 1965 5475 1999
rect 4875 1959 5475 1965
rect 4875 1926 5124 1959
rect 4875 1892 5122 1926
rect 5158 1925 5192 1959
rect 5226 1926 5475 1959
rect 5156 1892 5194 1925
rect 5228 1892 5475 1926
rect 4875 1890 5475 1892
rect 4875 1856 5124 1890
rect 5158 1856 5192 1890
rect 5226 1856 5475 1890
rect 4875 1853 5475 1856
rect 4875 1819 5122 1853
rect 5156 1821 5194 1853
rect 4875 1787 5124 1819
rect 5158 1787 5192 1821
rect 5228 1819 5475 1853
rect 5226 1787 5475 1819
rect 4875 1780 5475 1787
rect 4875 1746 5122 1780
rect 5156 1752 5194 1780
rect 4875 1718 5124 1746
rect 5158 1718 5192 1752
rect 5228 1746 5475 1780
rect 5226 1718 5475 1746
rect 4875 1707 5475 1718
rect 4875 1673 5122 1707
rect 5156 1683 5194 1707
rect 4875 1649 5124 1673
rect 5158 1649 5192 1683
rect 5228 1673 5475 1707
rect 5226 1649 5475 1673
rect 4875 1634 5475 1649
rect 4875 1600 5122 1634
rect 5156 1614 5194 1634
rect 4875 1580 5124 1600
rect 5158 1580 5192 1614
rect 5228 1600 5475 1634
rect 5226 1580 5475 1600
rect 4875 1561 5475 1580
rect 4875 1527 5122 1561
rect 5156 1545 5194 1561
rect 4875 1511 5124 1527
rect 5158 1511 5192 1545
rect 5228 1527 5475 1561
rect 5226 1511 5475 1527
rect 4875 1488 5475 1511
rect 4875 1454 5122 1488
rect 5156 1476 5194 1488
rect 4875 1442 5124 1454
rect 5158 1442 5192 1476
rect 5228 1454 5475 1488
rect 5226 1442 5475 1454
rect 4875 1415 5475 1442
rect 4875 1381 5122 1415
rect 5156 1407 5194 1415
rect 4875 1373 5124 1381
rect 5158 1373 5192 1407
rect 5228 1381 5475 1415
rect 5226 1373 5475 1381
rect 4875 1342 5475 1373
rect 4875 1308 5122 1342
rect 5156 1338 5194 1342
rect 4875 1304 5124 1308
rect 5158 1304 5192 1338
rect 5228 1308 5475 1342
rect 5226 1304 5475 1308
rect 4875 1269 5475 1304
rect 4875 1235 5122 1269
rect 5158 1235 5192 1269
rect 5228 1235 5475 1269
rect 4875 1135 5475 1235
rect 5777 11233 6377 11333
rect 5777 3279 6024 11233
rect 6130 3279 6377 11233
rect 5777 3270 6377 3279
rect 5777 3240 6026 3270
rect 5777 3206 6024 3240
rect 6060 3236 6094 3270
rect 6128 3240 6377 3270
rect 6058 3206 6096 3236
rect 6130 3206 6377 3240
rect 5777 3201 6377 3206
rect 5777 3167 6026 3201
rect 6060 3167 6094 3201
rect 6128 3167 6377 3201
rect 5777 3133 6024 3167
rect 6058 3133 6096 3167
rect 6130 3133 6377 3167
rect 5777 3132 6377 3133
rect 5777 3098 6026 3132
rect 6060 3098 6094 3132
rect 6128 3098 6377 3132
rect 5777 3094 6377 3098
rect 5777 3060 6024 3094
rect 6058 3063 6096 3094
rect 5777 3029 6026 3060
rect 6060 3029 6094 3063
rect 6130 3060 6377 3094
rect 6128 3029 6377 3060
rect 5777 3021 6377 3029
rect 5777 2987 6024 3021
rect 6058 2994 6096 3021
rect 5777 2960 6026 2987
rect 6060 2960 6094 2994
rect 6130 2987 6377 3021
rect 6128 2960 6377 2987
rect 5777 2948 6377 2960
rect 5777 2914 6024 2948
rect 6058 2925 6096 2948
rect 5777 2891 6026 2914
rect 6060 2891 6094 2925
rect 6130 2914 6377 2948
rect 6128 2891 6377 2914
rect 5777 2875 6377 2891
rect 5777 2841 6024 2875
rect 6058 2856 6096 2875
rect 5777 2822 6026 2841
rect 6060 2822 6094 2856
rect 6130 2841 6377 2875
rect 6128 2822 6377 2841
rect 5777 2802 6377 2822
rect 5777 2768 6024 2802
rect 6058 2787 6096 2802
rect 5777 2753 6026 2768
rect 6060 2753 6094 2787
rect 6130 2768 6377 2802
rect 6128 2753 6377 2768
rect 5777 2729 6377 2753
rect 5777 2695 6024 2729
rect 6058 2718 6096 2729
rect 5777 2684 6026 2695
rect 6060 2684 6094 2718
rect 6130 2695 6377 2729
rect 6128 2684 6377 2695
rect 5777 2656 6377 2684
rect 5777 2622 6024 2656
rect 6058 2649 6096 2656
rect 5777 2615 6026 2622
rect 6060 2615 6094 2649
rect 6130 2622 6377 2656
rect 6128 2615 6377 2622
rect 5777 2583 6377 2615
rect 5777 2549 6024 2583
rect 6058 2580 6096 2583
rect 5777 2546 6026 2549
rect 6060 2546 6094 2580
rect 6130 2549 6377 2583
rect 6128 2546 6377 2549
rect 5777 2511 6377 2546
rect 5777 2510 6026 2511
rect 5777 2476 6024 2510
rect 6060 2477 6094 2511
rect 6128 2510 6377 2511
rect 6058 2476 6096 2477
rect 6130 2476 6377 2510
rect 5777 2442 6377 2476
rect 5777 2437 6026 2442
rect 5777 2403 6024 2437
rect 6060 2408 6094 2442
rect 6128 2437 6377 2442
rect 6058 2403 6096 2408
rect 6130 2403 6377 2437
rect 5777 2373 6377 2403
rect 5777 2364 6026 2373
rect 5777 2330 6024 2364
rect 6060 2339 6094 2373
rect 6128 2364 6377 2373
rect 6058 2330 6096 2339
rect 6130 2330 6377 2364
rect 5777 2304 6377 2330
rect 5777 2291 6026 2304
rect 5777 2257 6024 2291
rect 6060 2270 6094 2304
rect 6128 2291 6377 2304
rect 6058 2257 6096 2270
rect 6130 2257 6377 2291
rect 5777 2235 6377 2257
rect 5777 2218 6026 2235
rect 5777 2184 6024 2218
rect 6060 2201 6094 2235
rect 6128 2218 6377 2235
rect 6058 2184 6096 2201
rect 6130 2184 6377 2218
rect 5777 2166 6377 2184
rect 5777 2145 6026 2166
rect 5777 2111 6024 2145
rect 6060 2132 6094 2166
rect 6128 2145 6377 2166
rect 6058 2111 6096 2132
rect 6130 2111 6377 2145
rect 5777 2097 6377 2111
rect 5777 2072 6026 2097
rect 5777 2038 6024 2072
rect 6060 2063 6094 2097
rect 6128 2072 6377 2097
rect 6058 2038 6096 2063
rect 6130 2038 6377 2072
rect 5777 2028 6377 2038
rect 5777 1999 6026 2028
rect 5777 1965 6024 1999
rect 6060 1994 6094 2028
rect 6128 1999 6377 2028
rect 6058 1965 6096 1994
rect 6130 1965 6377 1999
rect 5777 1959 6377 1965
rect 5777 1926 6026 1959
rect 5777 1892 6024 1926
rect 6060 1925 6094 1959
rect 6128 1926 6377 1959
rect 6058 1892 6096 1925
rect 6130 1892 6377 1926
rect 5777 1890 6377 1892
rect 5777 1856 6026 1890
rect 6060 1856 6094 1890
rect 6128 1856 6377 1890
rect 5777 1853 6377 1856
rect 5777 1819 6024 1853
rect 6058 1821 6096 1853
rect 5777 1787 6026 1819
rect 6060 1787 6094 1821
rect 6130 1819 6377 1853
rect 6128 1787 6377 1819
rect 5777 1780 6377 1787
rect 5777 1746 6024 1780
rect 6058 1752 6096 1780
rect 5777 1718 6026 1746
rect 6060 1718 6094 1752
rect 6130 1746 6377 1780
rect 6128 1718 6377 1746
rect 5777 1707 6377 1718
rect 5777 1673 6024 1707
rect 6058 1683 6096 1707
rect 5777 1649 6026 1673
rect 6060 1649 6094 1683
rect 6130 1673 6377 1707
rect 6128 1649 6377 1673
rect 5777 1634 6377 1649
rect 5777 1600 6024 1634
rect 6058 1614 6096 1634
rect 5777 1580 6026 1600
rect 6060 1580 6094 1614
rect 6130 1600 6377 1634
rect 6128 1580 6377 1600
rect 5777 1561 6377 1580
rect 5777 1527 6024 1561
rect 6058 1545 6096 1561
rect 5777 1511 6026 1527
rect 6060 1511 6094 1545
rect 6130 1527 6377 1561
rect 6128 1511 6377 1527
rect 5777 1488 6377 1511
rect 5777 1454 6024 1488
rect 6058 1476 6096 1488
rect 5777 1442 6026 1454
rect 6060 1442 6094 1476
rect 6130 1454 6377 1488
rect 6128 1442 6377 1454
rect 5777 1415 6377 1442
rect 5777 1381 6024 1415
rect 6058 1407 6096 1415
rect 5777 1373 6026 1381
rect 6060 1373 6094 1407
rect 6130 1381 6377 1415
rect 6128 1373 6377 1381
rect 5777 1342 6377 1373
rect 5777 1308 6024 1342
rect 6058 1338 6096 1342
rect 5777 1304 6026 1308
rect 6060 1304 6094 1338
rect 6130 1308 6377 1342
rect 6128 1304 6377 1308
rect 5777 1269 6377 1304
rect 5777 1235 6024 1269
rect 6060 1235 6094 1269
rect 6130 1235 6377 1269
rect 5777 1135 6377 1235
rect 6679 11233 7279 11333
rect 6679 3279 6926 11233
rect 7032 3279 7279 11233
rect 6679 3270 7279 3279
rect 6679 3240 6928 3270
rect 6679 3206 6926 3240
rect 6962 3236 6996 3270
rect 7030 3240 7279 3270
rect 6960 3206 6998 3236
rect 7032 3206 7279 3240
rect 6679 3201 7279 3206
rect 6679 3167 6928 3201
rect 6962 3167 6996 3201
rect 7030 3167 7279 3201
rect 6679 3133 6926 3167
rect 6960 3133 6998 3167
rect 7032 3133 7279 3167
rect 6679 3132 7279 3133
rect 6679 3098 6928 3132
rect 6962 3098 6996 3132
rect 7030 3098 7279 3132
rect 6679 3094 7279 3098
rect 6679 3060 6926 3094
rect 6960 3063 6998 3094
rect 6679 3029 6928 3060
rect 6962 3029 6996 3063
rect 7032 3060 7279 3094
rect 7030 3029 7279 3060
rect 6679 3021 7279 3029
rect 6679 2987 6926 3021
rect 6960 2994 6998 3021
rect 6679 2960 6928 2987
rect 6962 2960 6996 2994
rect 7032 2987 7279 3021
rect 7030 2960 7279 2987
rect 6679 2948 7279 2960
rect 6679 2914 6926 2948
rect 6960 2925 6998 2948
rect 6679 2891 6928 2914
rect 6962 2891 6996 2925
rect 7032 2914 7279 2948
rect 7030 2891 7279 2914
rect 6679 2875 7279 2891
rect 6679 2841 6926 2875
rect 6960 2856 6998 2875
rect 6679 2822 6928 2841
rect 6962 2822 6996 2856
rect 7032 2841 7279 2875
rect 7030 2822 7279 2841
rect 6679 2802 7279 2822
rect 6679 2768 6926 2802
rect 6960 2787 6998 2802
rect 6679 2753 6928 2768
rect 6962 2753 6996 2787
rect 7032 2768 7279 2802
rect 7030 2753 7279 2768
rect 6679 2729 7279 2753
rect 6679 2695 6926 2729
rect 6960 2718 6998 2729
rect 6679 2684 6928 2695
rect 6962 2684 6996 2718
rect 7032 2695 7279 2729
rect 7030 2684 7279 2695
rect 6679 2656 7279 2684
rect 6679 2622 6926 2656
rect 6960 2649 6998 2656
rect 6679 2615 6928 2622
rect 6962 2615 6996 2649
rect 7032 2622 7279 2656
rect 7030 2615 7279 2622
rect 6679 2583 7279 2615
rect 6679 2549 6926 2583
rect 6960 2580 6998 2583
rect 6679 2546 6928 2549
rect 6962 2546 6996 2580
rect 7032 2549 7279 2583
rect 7030 2546 7279 2549
rect 6679 2511 7279 2546
rect 6679 2510 6928 2511
rect 6679 2476 6926 2510
rect 6962 2477 6996 2511
rect 7030 2510 7279 2511
rect 6960 2476 6998 2477
rect 7032 2476 7279 2510
rect 6679 2442 7279 2476
rect 6679 2437 6928 2442
rect 6679 2403 6926 2437
rect 6962 2408 6996 2442
rect 7030 2437 7279 2442
rect 6960 2403 6998 2408
rect 7032 2403 7279 2437
rect 6679 2373 7279 2403
rect 6679 2364 6928 2373
rect 6679 2330 6926 2364
rect 6962 2339 6996 2373
rect 7030 2364 7279 2373
rect 6960 2330 6998 2339
rect 7032 2330 7279 2364
rect 6679 2304 7279 2330
rect 6679 2291 6928 2304
rect 6679 2257 6926 2291
rect 6962 2270 6996 2304
rect 7030 2291 7279 2304
rect 6960 2257 6998 2270
rect 7032 2257 7279 2291
rect 6679 2235 7279 2257
rect 6679 2218 6928 2235
rect 6679 2184 6926 2218
rect 6962 2201 6996 2235
rect 7030 2218 7279 2235
rect 6960 2184 6998 2201
rect 7032 2184 7279 2218
rect 6679 2166 7279 2184
rect 6679 2145 6928 2166
rect 6679 2111 6926 2145
rect 6962 2132 6996 2166
rect 7030 2145 7279 2166
rect 6960 2111 6998 2132
rect 7032 2111 7279 2145
rect 6679 2097 7279 2111
rect 6679 2072 6928 2097
rect 6679 2038 6926 2072
rect 6962 2063 6996 2097
rect 7030 2072 7279 2097
rect 6960 2038 6998 2063
rect 7032 2038 7279 2072
rect 6679 2028 7279 2038
rect 6679 1999 6928 2028
rect 6679 1965 6926 1999
rect 6962 1994 6996 2028
rect 7030 1999 7279 2028
rect 6960 1965 6998 1994
rect 7032 1965 7279 1999
rect 6679 1959 7279 1965
rect 6679 1926 6928 1959
rect 6679 1892 6926 1926
rect 6962 1925 6996 1959
rect 7030 1926 7279 1959
rect 6960 1892 6998 1925
rect 7032 1892 7279 1926
rect 6679 1890 7279 1892
rect 6679 1856 6928 1890
rect 6962 1856 6996 1890
rect 7030 1856 7279 1890
rect 6679 1853 7279 1856
rect 6679 1819 6926 1853
rect 6960 1821 6998 1853
rect 6679 1787 6928 1819
rect 6962 1787 6996 1821
rect 7032 1819 7279 1853
rect 7030 1787 7279 1819
rect 6679 1780 7279 1787
rect 6679 1746 6926 1780
rect 6960 1752 6998 1780
rect 6679 1718 6928 1746
rect 6962 1718 6996 1752
rect 7032 1746 7279 1780
rect 7030 1718 7279 1746
rect 6679 1707 7279 1718
rect 6679 1673 6926 1707
rect 6960 1683 6998 1707
rect 6679 1649 6928 1673
rect 6962 1649 6996 1683
rect 7032 1673 7279 1707
rect 7030 1649 7279 1673
rect 6679 1634 7279 1649
rect 6679 1600 6926 1634
rect 6960 1614 6998 1634
rect 6679 1580 6928 1600
rect 6962 1580 6996 1614
rect 7032 1600 7279 1634
rect 7030 1580 7279 1600
rect 6679 1561 7279 1580
rect 6679 1527 6926 1561
rect 6960 1545 6998 1561
rect 6679 1511 6928 1527
rect 6962 1511 6996 1545
rect 7032 1527 7279 1561
rect 7030 1511 7279 1527
rect 6679 1488 7279 1511
rect 6679 1454 6926 1488
rect 6960 1476 6998 1488
rect 6679 1442 6928 1454
rect 6962 1442 6996 1476
rect 7032 1454 7279 1488
rect 7030 1442 7279 1454
rect 6679 1415 7279 1442
rect 6679 1381 6926 1415
rect 6960 1407 6998 1415
rect 6679 1373 6928 1381
rect 6962 1373 6996 1407
rect 7032 1381 7279 1415
rect 7030 1373 7279 1381
rect 6679 1342 7279 1373
rect 6679 1308 6926 1342
rect 6960 1338 6998 1342
rect 6679 1304 6928 1308
rect 6962 1304 6996 1338
rect 7032 1308 7279 1342
rect 7030 1304 7279 1308
rect 6679 1269 7279 1304
rect 6679 1235 6926 1269
rect 6962 1235 6996 1269
rect 7032 1235 7279 1269
rect 6679 1135 7279 1235
rect 7581 11233 8181 11333
rect 7581 3279 7828 11233
rect 7934 3279 8181 11233
rect 7581 3270 8181 3279
rect 7581 3240 7830 3270
rect 7581 3206 7828 3240
rect 7864 3236 7898 3270
rect 7932 3240 8181 3270
rect 7862 3206 7900 3236
rect 7934 3206 8181 3240
rect 7581 3201 8181 3206
rect 7581 3167 7830 3201
rect 7864 3167 7898 3201
rect 7932 3167 8181 3201
rect 7581 3133 7828 3167
rect 7862 3133 7900 3167
rect 7934 3133 8181 3167
rect 7581 3132 8181 3133
rect 7581 3098 7830 3132
rect 7864 3098 7898 3132
rect 7932 3098 8181 3132
rect 7581 3094 8181 3098
rect 7581 3060 7828 3094
rect 7862 3063 7900 3094
rect 7581 3029 7830 3060
rect 7864 3029 7898 3063
rect 7934 3060 8181 3094
rect 7932 3029 8181 3060
rect 7581 3021 8181 3029
rect 7581 2987 7828 3021
rect 7862 2994 7900 3021
rect 7581 2960 7830 2987
rect 7864 2960 7898 2994
rect 7934 2987 8181 3021
rect 7932 2960 8181 2987
rect 7581 2948 8181 2960
rect 7581 2914 7828 2948
rect 7862 2925 7900 2948
rect 7581 2891 7830 2914
rect 7864 2891 7898 2925
rect 7934 2914 8181 2948
rect 7932 2891 8181 2914
rect 7581 2875 8181 2891
rect 7581 2841 7828 2875
rect 7862 2856 7900 2875
rect 7581 2822 7830 2841
rect 7864 2822 7898 2856
rect 7934 2841 8181 2875
rect 7932 2822 8181 2841
rect 7581 2802 8181 2822
rect 7581 2768 7828 2802
rect 7862 2787 7900 2802
rect 7581 2753 7830 2768
rect 7864 2753 7898 2787
rect 7934 2768 8181 2802
rect 7932 2753 8181 2768
rect 7581 2729 8181 2753
rect 7581 2695 7828 2729
rect 7862 2718 7900 2729
rect 7581 2684 7830 2695
rect 7864 2684 7898 2718
rect 7934 2695 8181 2729
rect 7932 2684 8181 2695
rect 7581 2656 8181 2684
rect 7581 2622 7828 2656
rect 7862 2649 7900 2656
rect 7581 2615 7830 2622
rect 7864 2615 7898 2649
rect 7934 2622 8181 2656
rect 7932 2615 8181 2622
rect 7581 2583 8181 2615
rect 7581 2549 7828 2583
rect 7862 2580 7900 2583
rect 7581 2546 7830 2549
rect 7864 2546 7898 2580
rect 7934 2549 8181 2583
rect 7932 2546 8181 2549
rect 7581 2511 8181 2546
rect 7581 2510 7830 2511
rect 7581 2476 7828 2510
rect 7864 2477 7898 2511
rect 7932 2510 8181 2511
rect 7862 2476 7900 2477
rect 7934 2476 8181 2510
rect 7581 2442 8181 2476
rect 7581 2437 7830 2442
rect 7581 2403 7828 2437
rect 7864 2408 7898 2442
rect 7932 2437 8181 2442
rect 7862 2403 7900 2408
rect 7934 2403 8181 2437
rect 7581 2373 8181 2403
rect 7581 2364 7830 2373
rect 7581 2330 7828 2364
rect 7864 2339 7898 2373
rect 7932 2364 8181 2373
rect 7862 2330 7900 2339
rect 7934 2330 8181 2364
rect 7581 2304 8181 2330
rect 7581 2291 7830 2304
rect 7581 2257 7828 2291
rect 7864 2270 7898 2304
rect 7932 2291 8181 2304
rect 7862 2257 7900 2270
rect 7934 2257 8181 2291
rect 7581 2235 8181 2257
rect 7581 2218 7830 2235
rect 7581 2184 7828 2218
rect 7864 2201 7898 2235
rect 7932 2218 8181 2235
rect 7862 2184 7900 2201
rect 7934 2184 8181 2218
rect 7581 2166 8181 2184
rect 7581 2145 7830 2166
rect 7581 2111 7828 2145
rect 7864 2132 7898 2166
rect 7932 2145 8181 2166
rect 7862 2111 7900 2132
rect 7934 2111 8181 2145
rect 7581 2097 8181 2111
rect 7581 2072 7830 2097
rect 7581 2038 7828 2072
rect 7864 2063 7898 2097
rect 7932 2072 8181 2097
rect 7862 2038 7900 2063
rect 7934 2038 8181 2072
rect 7581 2028 8181 2038
rect 7581 1999 7830 2028
rect 7581 1965 7828 1999
rect 7864 1994 7898 2028
rect 7932 1999 8181 2028
rect 7862 1965 7900 1994
rect 7934 1965 8181 1999
rect 7581 1959 8181 1965
rect 7581 1926 7830 1959
rect 7581 1892 7828 1926
rect 7864 1925 7898 1959
rect 7932 1926 8181 1959
rect 7862 1892 7900 1925
rect 7934 1892 8181 1926
rect 7581 1890 8181 1892
rect 7581 1856 7830 1890
rect 7864 1856 7898 1890
rect 7932 1856 8181 1890
rect 7581 1853 8181 1856
rect 7581 1819 7828 1853
rect 7862 1821 7900 1853
rect 7581 1787 7830 1819
rect 7864 1787 7898 1821
rect 7934 1819 8181 1853
rect 7932 1787 8181 1819
rect 7581 1780 8181 1787
rect 7581 1746 7828 1780
rect 7862 1752 7900 1780
rect 7581 1718 7830 1746
rect 7864 1718 7898 1752
rect 7934 1746 8181 1780
rect 7932 1718 8181 1746
rect 7581 1707 8181 1718
rect 7581 1673 7828 1707
rect 7862 1683 7900 1707
rect 7581 1649 7830 1673
rect 7864 1649 7898 1683
rect 7934 1673 8181 1707
rect 7932 1649 8181 1673
rect 7581 1634 8181 1649
rect 7581 1600 7828 1634
rect 7862 1614 7900 1634
rect 7581 1580 7830 1600
rect 7864 1580 7898 1614
rect 7934 1600 8181 1634
rect 7932 1580 8181 1600
rect 7581 1561 8181 1580
rect 7581 1527 7828 1561
rect 7862 1545 7900 1561
rect 7581 1511 7830 1527
rect 7864 1511 7898 1545
rect 7934 1527 8181 1561
rect 7932 1511 8181 1527
rect 7581 1488 8181 1511
rect 7581 1454 7828 1488
rect 7862 1476 7900 1488
rect 7581 1442 7830 1454
rect 7864 1442 7898 1476
rect 7934 1454 8181 1488
rect 7932 1442 8181 1454
rect 7581 1415 8181 1442
rect 7581 1381 7828 1415
rect 7862 1407 7900 1415
rect 7581 1373 7830 1381
rect 7864 1373 7898 1407
rect 7934 1381 8181 1415
rect 7932 1373 8181 1381
rect 7581 1342 8181 1373
rect 7581 1308 7828 1342
rect 7862 1338 7900 1342
rect 7581 1304 7830 1308
rect 7864 1304 7898 1338
rect 7934 1308 8181 1342
rect 7932 1304 8181 1308
rect 7581 1269 8181 1304
rect 7581 1235 7828 1269
rect 7864 1235 7898 1269
rect 7934 1235 8181 1269
rect 7581 1135 8181 1235
rect 8483 11233 9083 11333
rect 8483 3279 8730 11233
rect 8836 3279 9083 11233
rect 8483 3270 9083 3279
rect 8483 3240 8732 3270
rect 8483 3206 8730 3240
rect 8766 3236 8800 3270
rect 8834 3240 9083 3270
rect 8764 3206 8802 3236
rect 8836 3206 9083 3240
rect 8483 3201 9083 3206
rect 8483 3167 8732 3201
rect 8766 3167 8800 3201
rect 8834 3167 9083 3201
rect 8483 3133 8730 3167
rect 8764 3133 8802 3167
rect 8836 3133 9083 3167
rect 8483 3132 9083 3133
rect 8483 3098 8732 3132
rect 8766 3098 8800 3132
rect 8834 3098 9083 3132
rect 8483 3094 9083 3098
rect 8483 3060 8730 3094
rect 8764 3063 8802 3094
rect 8483 3029 8732 3060
rect 8766 3029 8800 3063
rect 8836 3060 9083 3094
rect 8834 3029 9083 3060
rect 8483 3021 9083 3029
rect 8483 2987 8730 3021
rect 8764 2994 8802 3021
rect 8483 2960 8732 2987
rect 8766 2960 8800 2994
rect 8836 2987 9083 3021
rect 8834 2960 9083 2987
rect 8483 2948 9083 2960
rect 8483 2914 8730 2948
rect 8764 2925 8802 2948
rect 8483 2891 8732 2914
rect 8766 2891 8800 2925
rect 8836 2914 9083 2948
rect 8834 2891 9083 2914
rect 8483 2875 9083 2891
rect 8483 2841 8730 2875
rect 8764 2856 8802 2875
rect 8483 2822 8732 2841
rect 8766 2822 8800 2856
rect 8836 2841 9083 2875
rect 8834 2822 9083 2841
rect 8483 2802 9083 2822
rect 8483 2768 8730 2802
rect 8764 2787 8802 2802
rect 8483 2753 8732 2768
rect 8766 2753 8800 2787
rect 8836 2768 9083 2802
rect 8834 2753 9083 2768
rect 8483 2729 9083 2753
rect 8483 2695 8730 2729
rect 8764 2718 8802 2729
rect 8483 2684 8732 2695
rect 8766 2684 8800 2718
rect 8836 2695 9083 2729
rect 8834 2684 9083 2695
rect 8483 2656 9083 2684
rect 8483 2622 8730 2656
rect 8764 2649 8802 2656
rect 8483 2615 8732 2622
rect 8766 2615 8800 2649
rect 8836 2622 9083 2656
rect 8834 2615 9083 2622
rect 8483 2583 9083 2615
rect 8483 2549 8730 2583
rect 8764 2580 8802 2583
rect 8483 2546 8732 2549
rect 8766 2546 8800 2580
rect 8836 2549 9083 2583
rect 8834 2546 9083 2549
rect 8483 2511 9083 2546
rect 8483 2510 8732 2511
rect 8483 2476 8730 2510
rect 8766 2477 8800 2511
rect 8834 2510 9083 2511
rect 8764 2476 8802 2477
rect 8836 2476 9083 2510
rect 8483 2442 9083 2476
rect 8483 2437 8732 2442
rect 8483 2403 8730 2437
rect 8766 2408 8800 2442
rect 8834 2437 9083 2442
rect 8764 2403 8802 2408
rect 8836 2403 9083 2437
rect 8483 2373 9083 2403
rect 8483 2364 8732 2373
rect 8483 2330 8730 2364
rect 8766 2339 8800 2373
rect 8834 2364 9083 2373
rect 8764 2330 8802 2339
rect 8836 2330 9083 2364
rect 8483 2304 9083 2330
rect 8483 2291 8732 2304
rect 8483 2257 8730 2291
rect 8766 2270 8800 2304
rect 8834 2291 9083 2304
rect 8764 2257 8802 2270
rect 8836 2257 9083 2291
rect 8483 2235 9083 2257
rect 8483 2218 8732 2235
rect 8483 2184 8730 2218
rect 8766 2201 8800 2235
rect 8834 2218 9083 2235
rect 8764 2184 8802 2201
rect 8836 2184 9083 2218
rect 8483 2166 9083 2184
rect 8483 2145 8732 2166
rect 8483 2111 8730 2145
rect 8766 2132 8800 2166
rect 8834 2145 9083 2166
rect 8764 2111 8802 2132
rect 8836 2111 9083 2145
rect 8483 2097 9083 2111
rect 8483 2072 8732 2097
rect 8483 2038 8730 2072
rect 8766 2063 8800 2097
rect 8834 2072 9083 2097
rect 8764 2038 8802 2063
rect 8836 2038 9083 2072
rect 8483 2028 9083 2038
rect 8483 1999 8732 2028
rect 8483 1965 8730 1999
rect 8766 1994 8800 2028
rect 8834 1999 9083 2028
rect 8764 1965 8802 1994
rect 8836 1965 9083 1999
rect 8483 1959 9083 1965
rect 8483 1926 8732 1959
rect 8483 1892 8730 1926
rect 8766 1925 8800 1959
rect 8834 1926 9083 1959
rect 8764 1892 8802 1925
rect 8836 1892 9083 1926
rect 8483 1890 9083 1892
rect 8483 1856 8732 1890
rect 8766 1856 8800 1890
rect 8834 1856 9083 1890
rect 8483 1853 9083 1856
rect 8483 1819 8730 1853
rect 8764 1821 8802 1853
rect 8483 1787 8732 1819
rect 8766 1787 8800 1821
rect 8836 1819 9083 1853
rect 8834 1787 9083 1819
rect 8483 1780 9083 1787
rect 8483 1746 8730 1780
rect 8764 1752 8802 1780
rect 8483 1718 8732 1746
rect 8766 1718 8800 1752
rect 8836 1746 9083 1780
rect 8834 1718 9083 1746
rect 8483 1707 9083 1718
rect 8483 1673 8730 1707
rect 8764 1683 8802 1707
rect 8483 1649 8732 1673
rect 8766 1649 8800 1683
rect 8836 1673 9083 1707
rect 8834 1649 9083 1673
rect 8483 1634 9083 1649
rect 8483 1600 8730 1634
rect 8764 1614 8802 1634
rect 8483 1580 8732 1600
rect 8766 1580 8800 1614
rect 8836 1600 9083 1634
rect 8834 1580 9083 1600
rect 8483 1561 9083 1580
rect 8483 1527 8730 1561
rect 8764 1545 8802 1561
rect 8483 1511 8732 1527
rect 8766 1511 8800 1545
rect 8836 1527 9083 1561
rect 8834 1511 9083 1527
rect 8483 1488 9083 1511
rect 8483 1454 8730 1488
rect 8764 1476 8802 1488
rect 8483 1442 8732 1454
rect 8766 1442 8800 1476
rect 8836 1454 9083 1488
rect 8834 1442 9083 1454
rect 8483 1415 9083 1442
rect 8483 1381 8730 1415
rect 8764 1407 8802 1415
rect 8483 1373 8732 1381
rect 8766 1373 8800 1407
rect 8836 1381 9083 1415
rect 8834 1373 9083 1381
rect 8483 1342 9083 1373
rect 8483 1308 8730 1342
rect 8764 1338 8802 1342
rect 8483 1304 8732 1308
rect 8766 1304 8800 1338
rect 8836 1308 9083 1342
rect 8834 1304 9083 1308
rect 8483 1269 9083 1304
rect 8483 1235 8730 1269
rect 8766 1235 8800 1269
rect 8836 1235 9083 1269
rect 8483 1135 9083 1235
rect 9385 11233 9985 11333
rect 9385 3279 9632 11233
rect 9738 3279 9985 11233
rect 9385 3270 9985 3279
rect 9385 3240 9634 3270
rect 9385 3206 9632 3240
rect 9668 3236 9702 3270
rect 9736 3240 9985 3270
rect 9666 3206 9704 3236
rect 9738 3206 9985 3240
rect 9385 3201 9985 3206
rect 9385 3167 9634 3201
rect 9668 3167 9702 3201
rect 9736 3167 9985 3201
rect 9385 3133 9632 3167
rect 9666 3133 9704 3167
rect 9738 3133 9985 3167
rect 9385 3132 9985 3133
rect 9385 3098 9634 3132
rect 9668 3098 9702 3132
rect 9736 3098 9985 3132
rect 9385 3094 9985 3098
rect 9385 3060 9632 3094
rect 9666 3063 9704 3094
rect 9385 3029 9634 3060
rect 9668 3029 9702 3063
rect 9738 3060 9985 3094
rect 9736 3029 9985 3060
rect 9385 3021 9985 3029
rect 9385 2987 9632 3021
rect 9666 2994 9704 3021
rect 9385 2960 9634 2987
rect 9668 2960 9702 2994
rect 9738 2987 9985 3021
rect 9736 2960 9985 2987
rect 9385 2948 9985 2960
rect 9385 2914 9632 2948
rect 9666 2925 9704 2948
rect 9385 2891 9634 2914
rect 9668 2891 9702 2925
rect 9738 2914 9985 2948
rect 9736 2891 9985 2914
rect 9385 2875 9985 2891
rect 9385 2841 9632 2875
rect 9666 2856 9704 2875
rect 9385 2822 9634 2841
rect 9668 2822 9702 2856
rect 9738 2841 9985 2875
rect 9736 2822 9985 2841
rect 9385 2802 9985 2822
rect 9385 2768 9632 2802
rect 9666 2787 9704 2802
rect 9385 2753 9634 2768
rect 9668 2753 9702 2787
rect 9738 2768 9985 2802
rect 9736 2753 9985 2768
rect 9385 2729 9985 2753
rect 9385 2695 9632 2729
rect 9666 2718 9704 2729
rect 9385 2684 9634 2695
rect 9668 2684 9702 2718
rect 9738 2695 9985 2729
rect 9736 2684 9985 2695
rect 9385 2656 9985 2684
rect 9385 2622 9632 2656
rect 9666 2649 9704 2656
rect 9385 2615 9634 2622
rect 9668 2615 9702 2649
rect 9738 2622 9985 2656
rect 9736 2615 9985 2622
rect 9385 2583 9985 2615
rect 9385 2549 9632 2583
rect 9666 2580 9704 2583
rect 9385 2546 9634 2549
rect 9668 2546 9702 2580
rect 9738 2549 9985 2583
rect 9736 2546 9985 2549
rect 9385 2511 9985 2546
rect 9385 2510 9634 2511
rect 9385 2476 9632 2510
rect 9668 2477 9702 2511
rect 9736 2510 9985 2511
rect 9666 2476 9704 2477
rect 9738 2476 9985 2510
rect 9385 2442 9985 2476
rect 9385 2437 9634 2442
rect 9385 2403 9632 2437
rect 9668 2408 9702 2442
rect 9736 2437 9985 2442
rect 9666 2403 9704 2408
rect 9738 2403 9985 2437
rect 9385 2373 9985 2403
rect 9385 2364 9634 2373
rect 9385 2330 9632 2364
rect 9668 2339 9702 2373
rect 9736 2364 9985 2373
rect 9666 2330 9704 2339
rect 9738 2330 9985 2364
rect 9385 2304 9985 2330
rect 9385 2291 9634 2304
rect 9385 2257 9632 2291
rect 9668 2270 9702 2304
rect 9736 2291 9985 2304
rect 9666 2257 9704 2270
rect 9738 2257 9985 2291
rect 9385 2235 9985 2257
rect 9385 2218 9634 2235
rect 9385 2184 9632 2218
rect 9668 2201 9702 2235
rect 9736 2218 9985 2235
rect 9666 2184 9704 2201
rect 9738 2184 9985 2218
rect 9385 2166 9985 2184
rect 9385 2145 9634 2166
rect 9385 2111 9632 2145
rect 9668 2132 9702 2166
rect 9736 2145 9985 2166
rect 9666 2111 9704 2132
rect 9738 2111 9985 2145
rect 9385 2097 9985 2111
rect 9385 2072 9634 2097
rect 9385 2038 9632 2072
rect 9668 2063 9702 2097
rect 9736 2072 9985 2097
rect 9666 2038 9704 2063
rect 9738 2038 9985 2072
rect 9385 2028 9985 2038
rect 9385 1999 9634 2028
rect 9385 1965 9632 1999
rect 9668 1994 9702 2028
rect 9736 1999 9985 2028
rect 9666 1965 9704 1994
rect 9738 1965 9985 1999
rect 9385 1959 9985 1965
rect 9385 1926 9634 1959
rect 9385 1892 9632 1926
rect 9668 1925 9702 1959
rect 9736 1926 9985 1959
rect 9666 1892 9704 1925
rect 9738 1892 9985 1926
rect 9385 1890 9985 1892
rect 9385 1856 9634 1890
rect 9668 1856 9702 1890
rect 9736 1856 9985 1890
rect 9385 1853 9985 1856
rect 9385 1819 9632 1853
rect 9666 1821 9704 1853
rect 9385 1787 9634 1819
rect 9668 1787 9702 1821
rect 9738 1819 9985 1853
rect 9736 1787 9985 1819
rect 9385 1780 9985 1787
rect 9385 1746 9632 1780
rect 9666 1752 9704 1780
rect 9385 1718 9634 1746
rect 9668 1718 9702 1752
rect 9738 1746 9985 1780
rect 9736 1718 9985 1746
rect 9385 1707 9985 1718
rect 9385 1673 9632 1707
rect 9666 1683 9704 1707
rect 9385 1649 9634 1673
rect 9668 1649 9702 1683
rect 9738 1673 9985 1707
rect 9736 1649 9985 1673
rect 9385 1634 9985 1649
rect 9385 1600 9632 1634
rect 9666 1614 9704 1634
rect 9385 1580 9634 1600
rect 9668 1580 9702 1614
rect 9738 1600 9985 1634
rect 9736 1580 9985 1600
rect 9385 1561 9985 1580
rect 9385 1527 9632 1561
rect 9666 1545 9704 1561
rect 9385 1511 9634 1527
rect 9668 1511 9702 1545
rect 9738 1527 9985 1561
rect 9736 1511 9985 1527
rect 9385 1488 9985 1511
rect 9385 1454 9632 1488
rect 9666 1476 9704 1488
rect 9385 1442 9634 1454
rect 9668 1442 9702 1476
rect 9738 1454 9985 1488
rect 9736 1442 9985 1454
rect 9385 1415 9985 1442
rect 9385 1381 9632 1415
rect 9666 1407 9704 1415
rect 9385 1373 9634 1381
rect 9668 1373 9702 1407
rect 9738 1381 9985 1415
rect 9736 1373 9985 1381
rect 9385 1342 9985 1373
rect 9385 1308 9632 1342
rect 9666 1338 9704 1342
rect 9385 1304 9634 1308
rect 9668 1304 9702 1338
rect 9738 1308 9985 1342
rect 9736 1304 9985 1308
rect 9385 1269 9985 1304
rect 9385 1235 9632 1269
rect 9668 1235 9702 1269
rect 9738 1235 9985 1269
rect 9385 1135 9985 1235
rect 10287 11233 10887 11333
rect 10287 3279 10534 11233
rect 10640 3279 10887 11233
rect 10287 3270 10887 3279
rect 10287 3240 10536 3270
rect 10287 3206 10534 3240
rect 10570 3236 10604 3270
rect 10638 3240 10887 3270
rect 10568 3206 10606 3236
rect 10640 3206 10887 3240
rect 10287 3201 10887 3206
rect 10287 3167 10536 3201
rect 10570 3167 10604 3201
rect 10638 3167 10887 3201
rect 10287 3133 10534 3167
rect 10568 3133 10606 3167
rect 10640 3133 10887 3167
rect 10287 3132 10887 3133
rect 10287 3098 10536 3132
rect 10570 3098 10604 3132
rect 10638 3098 10887 3132
rect 10287 3094 10887 3098
rect 10287 3060 10534 3094
rect 10568 3063 10606 3094
rect 10287 3029 10536 3060
rect 10570 3029 10604 3063
rect 10640 3060 10887 3094
rect 10638 3029 10887 3060
rect 10287 3021 10887 3029
rect 10287 2987 10534 3021
rect 10568 2994 10606 3021
rect 10287 2960 10536 2987
rect 10570 2960 10604 2994
rect 10640 2987 10887 3021
rect 10638 2960 10887 2987
rect 10287 2948 10887 2960
rect 10287 2914 10534 2948
rect 10568 2925 10606 2948
rect 10287 2891 10536 2914
rect 10570 2891 10604 2925
rect 10640 2914 10887 2948
rect 10638 2891 10887 2914
rect 10287 2875 10887 2891
rect 10287 2841 10534 2875
rect 10568 2856 10606 2875
rect 10287 2822 10536 2841
rect 10570 2822 10604 2856
rect 10640 2841 10887 2875
rect 10638 2822 10887 2841
rect 10287 2802 10887 2822
rect 10287 2768 10534 2802
rect 10568 2787 10606 2802
rect 10287 2753 10536 2768
rect 10570 2753 10604 2787
rect 10640 2768 10887 2802
rect 10638 2753 10887 2768
rect 10287 2729 10887 2753
rect 10287 2695 10534 2729
rect 10568 2718 10606 2729
rect 10287 2684 10536 2695
rect 10570 2684 10604 2718
rect 10640 2695 10887 2729
rect 10638 2684 10887 2695
rect 10287 2656 10887 2684
rect 10287 2622 10534 2656
rect 10568 2649 10606 2656
rect 10287 2615 10536 2622
rect 10570 2615 10604 2649
rect 10640 2622 10887 2656
rect 10638 2615 10887 2622
rect 10287 2583 10887 2615
rect 10287 2549 10534 2583
rect 10568 2580 10606 2583
rect 10287 2546 10536 2549
rect 10570 2546 10604 2580
rect 10640 2549 10887 2583
rect 10638 2546 10887 2549
rect 10287 2511 10887 2546
rect 10287 2510 10536 2511
rect 10287 2476 10534 2510
rect 10570 2477 10604 2511
rect 10638 2510 10887 2511
rect 10568 2476 10606 2477
rect 10640 2476 10887 2510
rect 10287 2442 10887 2476
rect 10287 2437 10536 2442
rect 10287 2403 10534 2437
rect 10570 2408 10604 2442
rect 10638 2437 10887 2442
rect 10568 2403 10606 2408
rect 10640 2403 10887 2437
rect 10287 2373 10887 2403
rect 10287 2364 10536 2373
rect 10287 2330 10534 2364
rect 10570 2339 10604 2373
rect 10638 2364 10887 2373
rect 10568 2330 10606 2339
rect 10640 2330 10887 2364
rect 10287 2304 10887 2330
rect 10287 2291 10536 2304
rect 10287 2257 10534 2291
rect 10570 2270 10604 2304
rect 10638 2291 10887 2304
rect 10568 2257 10606 2270
rect 10640 2257 10887 2291
rect 10287 2235 10887 2257
rect 10287 2218 10536 2235
rect 10287 2184 10534 2218
rect 10570 2201 10604 2235
rect 10638 2218 10887 2235
rect 10568 2184 10606 2201
rect 10640 2184 10887 2218
rect 10287 2166 10887 2184
rect 10287 2145 10536 2166
rect 10287 2111 10534 2145
rect 10570 2132 10604 2166
rect 10638 2145 10887 2166
rect 10568 2111 10606 2132
rect 10640 2111 10887 2145
rect 10287 2097 10887 2111
rect 10287 2072 10536 2097
rect 10287 2038 10534 2072
rect 10570 2063 10604 2097
rect 10638 2072 10887 2097
rect 10568 2038 10606 2063
rect 10640 2038 10887 2072
rect 10287 2028 10887 2038
rect 10287 1999 10536 2028
rect 10287 1965 10534 1999
rect 10570 1994 10604 2028
rect 10638 1999 10887 2028
rect 10568 1965 10606 1994
rect 10640 1965 10887 1999
rect 10287 1959 10887 1965
rect 10287 1926 10536 1959
rect 10287 1892 10534 1926
rect 10570 1925 10604 1959
rect 10638 1926 10887 1959
rect 10568 1892 10606 1925
rect 10640 1892 10887 1926
rect 10287 1890 10887 1892
rect 10287 1856 10536 1890
rect 10570 1856 10604 1890
rect 10638 1856 10887 1890
rect 10287 1853 10887 1856
rect 10287 1819 10534 1853
rect 10568 1821 10606 1853
rect 10287 1787 10536 1819
rect 10570 1787 10604 1821
rect 10640 1819 10887 1853
rect 10638 1787 10887 1819
rect 10287 1780 10887 1787
rect 10287 1746 10534 1780
rect 10568 1752 10606 1780
rect 10287 1718 10536 1746
rect 10570 1718 10604 1752
rect 10640 1746 10887 1780
rect 10638 1718 10887 1746
rect 10287 1707 10887 1718
rect 10287 1673 10534 1707
rect 10568 1683 10606 1707
rect 10287 1649 10536 1673
rect 10570 1649 10604 1683
rect 10640 1673 10887 1707
rect 10638 1649 10887 1673
rect 10287 1634 10887 1649
rect 10287 1600 10534 1634
rect 10568 1614 10606 1634
rect 10287 1580 10536 1600
rect 10570 1580 10604 1614
rect 10640 1600 10887 1634
rect 10638 1580 10887 1600
rect 10287 1561 10887 1580
rect 10287 1527 10534 1561
rect 10568 1545 10606 1561
rect 10287 1511 10536 1527
rect 10570 1511 10604 1545
rect 10640 1527 10887 1561
rect 10638 1511 10887 1527
rect 10287 1488 10887 1511
rect 10287 1454 10534 1488
rect 10568 1476 10606 1488
rect 10287 1442 10536 1454
rect 10570 1442 10604 1476
rect 10640 1454 10887 1488
rect 10638 1442 10887 1454
rect 10287 1415 10887 1442
rect 10287 1381 10534 1415
rect 10568 1407 10606 1415
rect 10287 1373 10536 1381
rect 10570 1373 10604 1407
rect 10640 1381 10887 1415
rect 10638 1373 10887 1381
rect 10287 1342 10887 1373
rect 10287 1308 10534 1342
rect 10568 1338 10606 1342
rect 10287 1304 10536 1308
rect 10570 1304 10604 1338
rect 10640 1308 10887 1342
rect 10638 1304 10887 1308
rect 10287 1269 10887 1304
rect 10287 1235 10534 1269
rect 10570 1235 10604 1269
rect 10640 1235 10887 1269
rect 10287 1135 10887 1235
rect 11189 11233 11789 11333
rect 11189 3279 11436 11233
rect 11542 3279 11789 11233
rect 11189 3270 11789 3279
rect 11189 3240 11438 3270
rect 11189 3206 11436 3240
rect 11472 3236 11506 3270
rect 11540 3240 11789 3270
rect 11470 3206 11508 3236
rect 11542 3206 11789 3240
rect 11189 3201 11789 3206
rect 11189 3167 11438 3201
rect 11472 3167 11506 3201
rect 11540 3167 11789 3201
rect 11189 3133 11436 3167
rect 11470 3133 11508 3167
rect 11542 3133 11789 3167
rect 11189 3132 11789 3133
rect 11189 3098 11438 3132
rect 11472 3098 11506 3132
rect 11540 3098 11789 3132
rect 11189 3094 11789 3098
rect 11189 3060 11436 3094
rect 11470 3063 11508 3094
rect 11189 3029 11438 3060
rect 11472 3029 11506 3063
rect 11542 3060 11789 3094
rect 11540 3029 11789 3060
rect 11189 3021 11789 3029
rect 11189 2987 11436 3021
rect 11470 2994 11508 3021
rect 11189 2960 11438 2987
rect 11472 2960 11506 2994
rect 11542 2987 11789 3021
rect 11540 2960 11789 2987
rect 11189 2948 11789 2960
rect 11189 2914 11436 2948
rect 11470 2925 11508 2948
rect 11189 2891 11438 2914
rect 11472 2891 11506 2925
rect 11542 2914 11789 2948
rect 11540 2891 11789 2914
rect 11189 2875 11789 2891
rect 11189 2841 11436 2875
rect 11470 2856 11508 2875
rect 11189 2822 11438 2841
rect 11472 2822 11506 2856
rect 11542 2841 11789 2875
rect 11540 2822 11789 2841
rect 11189 2802 11789 2822
rect 11189 2768 11436 2802
rect 11470 2787 11508 2802
rect 11189 2753 11438 2768
rect 11472 2753 11506 2787
rect 11542 2768 11789 2802
rect 11540 2753 11789 2768
rect 11189 2729 11789 2753
rect 11189 2695 11436 2729
rect 11470 2718 11508 2729
rect 11189 2684 11438 2695
rect 11472 2684 11506 2718
rect 11542 2695 11789 2729
rect 11540 2684 11789 2695
rect 11189 2656 11789 2684
rect 11189 2622 11436 2656
rect 11470 2649 11508 2656
rect 11189 2615 11438 2622
rect 11472 2615 11506 2649
rect 11542 2622 11789 2656
rect 11540 2615 11789 2622
rect 11189 2583 11789 2615
rect 11189 2549 11436 2583
rect 11470 2580 11508 2583
rect 11189 2546 11438 2549
rect 11472 2546 11506 2580
rect 11542 2549 11789 2583
rect 11540 2546 11789 2549
rect 11189 2511 11789 2546
rect 11189 2510 11438 2511
rect 11189 2476 11436 2510
rect 11472 2477 11506 2511
rect 11540 2510 11789 2511
rect 11470 2476 11508 2477
rect 11542 2476 11789 2510
rect 11189 2442 11789 2476
rect 11189 2437 11438 2442
rect 11189 2403 11436 2437
rect 11472 2408 11506 2442
rect 11540 2437 11789 2442
rect 11470 2403 11508 2408
rect 11542 2403 11789 2437
rect 11189 2373 11789 2403
rect 11189 2364 11438 2373
rect 11189 2330 11436 2364
rect 11472 2339 11506 2373
rect 11540 2364 11789 2373
rect 11470 2330 11508 2339
rect 11542 2330 11789 2364
rect 11189 2304 11789 2330
rect 11189 2291 11438 2304
rect 11189 2257 11436 2291
rect 11472 2270 11506 2304
rect 11540 2291 11789 2304
rect 11470 2257 11508 2270
rect 11542 2257 11789 2291
rect 11189 2235 11789 2257
rect 11189 2218 11438 2235
rect 11189 2184 11436 2218
rect 11472 2201 11506 2235
rect 11540 2218 11789 2235
rect 11470 2184 11508 2201
rect 11542 2184 11789 2218
rect 11189 2166 11789 2184
rect 11189 2145 11438 2166
rect 11189 2111 11436 2145
rect 11472 2132 11506 2166
rect 11540 2145 11789 2166
rect 11470 2111 11508 2132
rect 11542 2111 11789 2145
rect 11189 2097 11789 2111
rect 11189 2072 11438 2097
rect 11189 2038 11436 2072
rect 11472 2063 11506 2097
rect 11540 2072 11789 2097
rect 11470 2038 11508 2063
rect 11542 2038 11789 2072
rect 11189 2028 11789 2038
rect 11189 1999 11438 2028
rect 11189 1965 11436 1999
rect 11472 1994 11506 2028
rect 11540 1999 11789 2028
rect 11470 1965 11508 1994
rect 11542 1965 11789 1999
rect 11189 1959 11789 1965
rect 11189 1926 11438 1959
rect 11189 1892 11436 1926
rect 11472 1925 11506 1959
rect 11540 1926 11789 1959
rect 11470 1892 11508 1925
rect 11542 1892 11789 1926
rect 11189 1890 11789 1892
rect 11189 1856 11438 1890
rect 11472 1856 11506 1890
rect 11540 1856 11789 1890
rect 11189 1853 11789 1856
rect 11189 1819 11436 1853
rect 11470 1821 11508 1853
rect 11189 1787 11438 1819
rect 11472 1787 11506 1821
rect 11542 1819 11789 1853
rect 11540 1787 11789 1819
rect 11189 1780 11789 1787
rect 11189 1746 11436 1780
rect 11470 1752 11508 1780
rect 11189 1718 11438 1746
rect 11472 1718 11506 1752
rect 11542 1746 11789 1780
rect 11540 1718 11789 1746
rect 11189 1707 11789 1718
rect 11189 1673 11436 1707
rect 11470 1683 11508 1707
rect 11189 1649 11438 1673
rect 11472 1649 11506 1683
rect 11542 1673 11789 1707
rect 11540 1649 11789 1673
rect 11189 1634 11789 1649
rect 11189 1600 11436 1634
rect 11470 1614 11508 1634
rect 11189 1580 11438 1600
rect 11472 1580 11506 1614
rect 11542 1600 11789 1634
rect 11540 1580 11789 1600
rect 11189 1561 11789 1580
rect 11189 1527 11436 1561
rect 11470 1545 11508 1561
rect 11189 1511 11438 1527
rect 11472 1511 11506 1545
rect 11542 1527 11789 1561
rect 11540 1511 11789 1527
rect 11189 1488 11789 1511
rect 11189 1454 11436 1488
rect 11470 1476 11508 1488
rect 11189 1442 11438 1454
rect 11472 1442 11506 1476
rect 11542 1454 11789 1488
rect 11540 1442 11789 1454
rect 11189 1415 11789 1442
rect 11189 1381 11436 1415
rect 11470 1407 11508 1415
rect 11189 1373 11438 1381
rect 11472 1373 11506 1407
rect 11542 1381 11789 1415
rect 11540 1373 11789 1381
rect 11189 1342 11789 1373
rect 11189 1308 11436 1342
rect 11470 1338 11508 1342
rect 11189 1304 11438 1308
rect 11472 1304 11506 1338
rect 11542 1308 11789 1342
rect 11540 1304 11789 1308
rect 11189 1269 11789 1304
rect 11189 1235 11436 1269
rect 11472 1235 11506 1269
rect 11542 1235 11789 1269
rect 11189 1135 11789 1235
rect 12091 11233 12691 11333
rect 12091 3279 12338 11233
rect 12444 3279 12691 11233
rect 12091 3270 12691 3279
rect 12091 3240 12340 3270
rect 12091 3206 12338 3240
rect 12374 3236 12408 3270
rect 12442 3240 12691 3270
rect 12372 3206 12410 3236
rect 12444 3206 12691 3240
rect 12091 3201 12691 3206
rect 12091 3167 12340 3201
rect 12374 3167 12408 3201
rect 12442 3167 12691 3201
rect 12091 3133 12338 3167
rect 12372 3133 12410 3167
rect 12444 3133 12691 3167
rect 12091 3132 12691 3133
rect 12091 3098 12340 3132
rect 12374 3098 12408 3132
rect 12442 3098 12691 3132
rect 12091 3094 12691 3098
rect 12091 3060 12338 3094
rect 12372 3063 12410 3094
rect 12091 3029 12340 3060
rect 12374 3029 12408 3063
rect 12444 3060 12691 3094
rect 12442 3029 12691 3060
rect 12091 3021 12691 3029
rect 12091 2987 12338 3021
rect 12372 2994 12410 3021
rect 12091 2960 12340 2987
rect 12374 2960 12408 2994
rect 12444 2987 12691 3021
rect 12442 2960 12691 2987
rect 12091 2948 12691 2960
rect 12091 2914 12338 2948
rect 12372 2925 12410 2948
rect 12091 2891 12340 2914
rect 12374 2891 12408 2925
rect 12444 2914 12691 2948
rect 12442 2891 12691 2914
rect 12091 2875 12691 2891
rect 12091 2841 12338 2875
rect 12372 2856 12410 2875
rect 12091 2822 12340 2841
rect 12374 2822 12408 2856
rect 12444 2841 12691 2875
rect 12442 2822 12691 2841
rect 12091 2802 12691 2822
rect 12091 2768 12338 2802
rect 12372 2787 12410 2802
rect 12091 2753 12340 2768
rect 12374 2753 12408 2787
rect 12444 2768 12691 2802
rect 12442 2753 12691 2768
rect 12091 2729 12691 2753
rect 12091 2695 12338 2729
rect 12372 2718 12410 2729
rect 12091 2684 12340 2695
rect 12374 2684 12408 2718
rect 12444 2695 12691 2729
rect 12442 2684 12691 2695
rect 12091 2656 12691 2684
rect 12091 2622 12338 2656
rect 12372 2649 12410 2656
rect 12091 2615 12340 2622
rect 12374 2615 12408 2649
rect 12444 2622 12691 2656
rect 12442 2615 12691 2622
rect 12091 2583 12691 2615
rect 12091 2549 12338 2583
rect 12372 2580 12410 2583
rect 12091 2546 12340 2549
rect 12374 2546 12408 2580
rect 12444 2549 12691 2583
rect 12442 2546 12691 2549
rect 12091 2511 12691 2546
rect 12091 2510 12340 2511
rect 12091 2476 12338 2510
rect 12374 2477 12408 2511
rect 12442 2510 12691 2511
rect 12372 2476 12410 2477
rect 12444 2476 12691 2510
rect 12091 2442 12691 2476
rect 12091 2437 12340 2442
rect 12091 2403 12338 2437
rect 12374 2408 12408 2442
rect 12442 2437 12691 2442
rect 12372 2403 12410 2408
rect 12444 2403 12691 2437
rect 12091 2373 12691 2403
rect 12091 2364 12340 2373
rect 12091 2330 12338 2364
rect 12374 2339 12408 2373
rect 12442 2364 12691 2373
rect 12372 2330 12410 2339
rect 12444 2330 12691 2364
rect 12091 2304 12691 2330
rect 12091 2291 12340 2304
rect 12091 2257 12338 2291
rect 12374 2270 12408 2304
rect 12442 2291 12691 2304
rect 12372 2257 12410 2270
rect 12444 2257 12691 2291
rect 12091 2235 12691 2257
rect 12091 2218 12340 2235
rect 12091 2184 12338 2218
rect 12374 2201 12408 2235
rect 12442 2218 12691 2235
rect 12372 2184 12410 2201
rect 12444 2184 12691 2218
rect 12091 2166 12691 2184
rect 12091 2145 12340 2166
rect 12091 2111 12338 2145
rect 12374 2132 12408 2166
rect 12442 2145 12691 2166
rect 12372 2111 12410 2132
rect 12444 2111 12691 2145
rect 12091 2097 12691 2111
rect 12091 2072 12340 2097
rect 12091 2038 12338 2072
rect 12374 2063 12408 2097
rect 12442 2072 12691 2097
rect 12372 2038 12410 2063
rect 12444 2038 12691 2072
rect 12091 2028 12691 2038
rect 12091 1999 12340 2028
rect 12091 1965 12338 1999
rect 12374 1994 12408 2028
rect 12442 1999 12691 2028
rect 12372 1965 12410 1994
rect 12444 1965 12691 1999
rect 12091 1959 12691 1965
rect 12091 1926 12340 1959
rect 12091 1892 12338 1926
rect 12374 1925 12408 1959
rect 12442 1926 12691 1959
rect 12372 1892 12410 1925
rect 12444 1892 12691 1926
rect 12091 1890 12691 1892
rect 12091 1856 12340 1890
rect 12374 1856 12408 1890
rect 12442 1856 12691 1890
rect 12091 1853 12691 1856
rect 12091 1819 12338 1853
rect 12372 1821 12410 1853
rect 12091 1787 12340 1819
rect 12374 1787 12408 1821
rect 12444 1819 12691 1853
rect 12442 1787 12691 1819
rect 12091 1780 12691 1787
rect 12091 1746 12338 1780
rect 12372 1752 12410 1780
rect 12091 1718 12340 1746
rect 12374 1718 12408 1752
rect 12444 1746 12691 1780
rect 12442 1718 12691 1746
rect 12091 1707 12691 1718
rect 12091 1673 12338 1707
rect 12372 1683 12410 1707
rect 12091 1649 12340 1673
rect 12374 1649 12408 1683
rect 12444 1673 12691 1707
rect 12442 1649 12691 1673
rect 12091 1634 12691 1649
rect 12091 1600 12338 1634
rect 12372 1614 12410 1634
rect 12091 1580 12340 1600
rect 12374 1580 12408 1614
rect 12444 1600 12691 1634
rect 12442 1580 12691 1600
rect 12091 1561 12691 1580
rect 12091 1527 12338 1561
rect 12372 1545 12410 1561
rect 12091 1511 12340 1527
rect 12374 1511 12408 1545
rect 12444 1527 12691 1561
rect 12442 1511 12691 1527
rect 12091 1488 12691 1511
rect 12091 1454 12338 1488
rect 12372 1476 12410 1488
rect 12091 1442 12340 1454
rect 12374 1442 12408 1476
rect 12444 1454 12691 1488
rect 12442 1442 12691 1454
rect 12091 1415 12691 1442
rect 12091 1381 12338 1415
rect 12372 1407 12410 1415
rect 12091 1373 12340 1381
rect 12374 1373 12408 1407
rect 12444 1381 12691 1415
rect 12442 1373 12691 1381
rect 12091 1342 12691 1373
rect 12091 1308 12338 1342
rect 12372 1338 12410 1342
rect 12091 1304 12340 1308
rect 12374 1304 12408 1338
rect 12444 1308 12691 1342
rect 12442 1304 12691 1308
rect 12091 1269 12691 1304
rect 12091 1235 12338 1269
rect 12374 1235 12408 1269
rect 12444 1235 12691 1269
rect 12091 1135 12691 1235
rect 12993 11233 13593 11333
rect 12993 3279 13240 11233
rect 13346 3279 13593 11233
rect 12993 3270 13593 3279
rect 12993 3240 13242 3270
rect 12993 3206 13240 3240
rect 13276 3236 13310 3270
rect 13344 3240 13593 3270
rect 13274 3206 13312 3236
rect 13346 3206 13593 3240
rect 12993 3201 13593 3206
rect 12993 3167 13242 3201
rect 13276 3167 13310 3201
rect 13344 3167 13593 3201
rect 12993 3133 13240 3167
rect 13274 3133 13312 3167
rect 13346 3133 13593 3167
rect 12993 3132 13593 3133
rect 12993 3098 13242 3132
rect 13276 3098 13310 3132
rect 13344 3098 13593 3132
rect 12993 3094 13593 3098
rect 12993 3060 13240 3094
rect 13274 3063 13312 3094
rect 12993 3029 13242 3060
rect 13276 3029 13310 3063
rect 13346 3060 13593 3094
rect 13344 3029 13593 3060
rect 12993 3021 13593 3029
rect 12993 2987 13240 3021
rect 13274 2994 13312 3021
rect 12993 2960 13242 2987
rect 13276 2960 13310 2994
rect 13346 2987 13593 3021
rect 13344 2960 13593 2987
rect 12993 2948 13593 2960
rect 12993 2914 13240 2948
rect 13274 2925 13312 2948
rect 12993 2891 13242 2914
rect 13276 2891 13310 2925
rect 13346 2914 13593 2948
rect 13344 2891 13593 2914
rect 12993 2875 13593 2891
rect 12993 2841 13240 2875
rect 13274 2856 13312 2875
rect 12993 2822 13242 2841
rect 13276 2822 13310 2856
rect 13346 2841 13593 2875
rect 13344 2822 13593 2841
rect 12993 2802 13593 2822
rect 12993 2768 13240 2802
rect 13274 2787 13312 2802
rect 12993 2753 13242 2768
rect 13276 2753 13310 2787
rect 13346 2768 13593 2802
rect 13344 2753 13593 2768
rect 12993 2729 13593 2753
rect 12993 2695 13240 2729
rect 13274 2718 13312 2729
rect 12993 2684 13242 2695
rect 13276 2684 13310 2718
rect 13346 2695 13593 2729
rect 13344 2684 13593 2695
rect 12993 2656 13593 2684
rect 12993 2622 13240 2656
rect 13274 2649 13312 2656
rect 12993 2615 13242 2622
rect 13276 2615 13310 2649
rect 13346 2622 13593 2656
rect 13344 2615 13593 2622
rect 12993 2583 13593 2615
rect 12993 2549 13240 2583
rect 13274 2580 13312 2583
rect 12993 2546 13242 2549
rect 13276 2546 13310 2580
rect 13346 2549 13593 2583
rect 13344 2546 13593 2549
rect 12993 2511 13593 2546
rect 12993 2510 13242 2511
rect 12993 2476 13240 2510
rect 13276 2477 13310 2511
rect 13344 2510 13593 2511
rect 13274 2476 13312 2477
rect 13346 2476 13593 2510
rect 12993 2442 13593 2476
rect 12993 2437 13242 2442
rect 12993 2403 13240 2437
rect 13276 2408 13310 2442
rect 13344 2437 13593 2442
rect 13274 2403 13312 2408
rect 13346 2403 13593 2437
rect 12993 2373 13593 2403
rect 12993 2364 13242 2373
rect 12993 2330 13240 2364
rect 13276 2339 13310 2373
rect 13344 2364 13593 2373
rect 13274 2330 13312 2339
rect 13346 2330 13593 2364
rect 12993 2304 13593 2330
rect 12993 2291 13242 2304
rect 12993 2257 13240 2291
rect 13276 2270 13310 2304
rect 13344 2291 13593 2304
rect 13274 2257 13312 2270
rect 13346 2257 13593 2291
rect 12993 2235 13593 2257
rect 12993 2218 13242 2235
rect 12993 2184 13240 2218
rect 13276 2201 13310 2235
rect 13344 2218 13593 2235
rect 13274 2184 13312 2201
rect 13346 2184 13593 2218
rect 12993 2166 13593 2184
rect 12993 2145 13242 2166
rect 12993 2111 13240 2145
rect 13276 2132 13310 2166
rect 13344 2145 13593 2166
rect 13274 2111 13312 2132
rect 13346 2111 13593 2145
rect 12993 2097 13593 2111
rect 12993 2072 13242 2097
rect 12993 2038 13240 2072
rect 13276 2063 13310 2097
rect 13344 2072 13593 2097
rect 13274 2038 13312 2063
rect 13346 2038 13593 2072
rect 12993 2028 13593 2038
rect 12993 1999 13242 2028
rect 12993 1965 13240 1999
rect 13276 1994 13310 2028
rect 13344 1999 13593 2028
rect 13274 1965 13312 1994
rect 13346 1965 13593 1999
rect 12993 1959 13593 1965
rect 12993 1926 13242 1959
rect 12993 1892 13240 1926
rect 13276 1925 13310 1959
rect 13344 1926 13593 1959
rect 13274 1892 13312 1925
rect 13346 1892 13593 1926
rect 12993 1890 13593 1892
rect 12993 1856 13242 1890
rect 13276 1856 13310 1890
rect 13344 1856 13593 1890
rect 12993 1853 13593 1856
rect 12993 1819 13240 1853
rect 13274 1821 13312 1853
rect 12993 1787 13242 1819
rect 13276 1787 13310 1821
rect 13346 1819 13593 1853
rect 13344 1787 13593 1819
rect 12993 1780 13593 1787
rect 12993 1746 13240 1780
rect 13274 1752 13312 1780
rect 12993 1718 13242 1746
rect 13276 1718 13310 1752
rect 13346 1746 13593 1780
rect 13344 1718 13593 1746
rect 12993 1707 13593 1718
rect 12993 1673 13240 1707
rect 13274 1683 13312 1707
rect 12993 1649 13242 1673
rect 13276 1649 13310 1683
rect 13346 1673 13593 1707
rect 13344 1649 13593 1673
rect 12993 1634 13593 1649
rect 12993 1600 13240 1634
rect 13274 1614 13312 1634
rect 12993 1580 13242 1600
rect 13276 1580 13310 1614
rect 13346 1600 13593 1634
rect 13344 1580 13593 1600
rect 12993 1561 13593 1580
rect 12993 1527 13240 1561
rect 13274 1545 13312 1561
rect 12993 1511 13242 1527
rect 13276 1511 13310 1545
rect 13346 1527 13593 1561
rect 13344 1511 13593 1527
rect 12993 1488 13593 1511
rect 12993 1454 13240 1488
rect 13274 1476 13312 1488
rect 12993 1442 13242 1454
rect 13276 1442 13310 1476
rect 13346 1454 13593 1488
rect 13344 1442 13593 1454
rect 12993 1415 13593 1442
rect 12993 1381 13240 1415
rect 13274 1407 13312 1415
rect 12993 1373 13242 1381
rect 13276 1373 13310 1407
rect 13346 1381 13593 1415
rect 13344 1373 13593 1381
rect 12993 1342 13593 1373
rect 12993 1308 13240 1342
rect 13274 1338 13312 1342
rect 12993 1304 13242 1308
rect 13276 1304 13310 1338
rect 13346 1308 13593 1342
rect 13344 1304 13593 1308
rect 12993 1269 13593 1304
rect 12993 1235 13240 1269
rect 13276 1235 13310 1269
rect 13346 1235 13593 1269
rect 12993 1135 13593 1235
rect 13895 11233 14495 11333
rect 13895 3279 14142 11233
rect 14248 3279 14495 11233
rect 13895 3270 14495 3279
rect 13895 3240 14144 3270
rect 13895 3206 14142 3240
rect 14178 3236 14212 3270
rect 14246 3240 14495 3270
rect 14176 3206 14214 3236
rect 14248 3206 14495 3240
rect 13895 3201 14495 3206
rect 13895 3167 14144 3201
rect 14178 3167 14212 3201
rect 14246 3167 14495 3201
rect 13895 3133 14142 3167
rect 14176 3133 14214 3167
rect 14248 3133 14495 3167
rect 13895 3132 14495 3133
rect 13895 3098 14144 3132
rect 14178 3098 14212 3132
rect 14246 3098 14495 3132
rect 13895 3094 14495 3098
rect 13895 3060 14142 3094
rect 14176 3063 14214 3094
rect 13895 3029 14144 3060
rect 14178 3029 14212 3063
rect 14248 3060 14495 3094
rect 14246 3029 14495 3060
rect 13895 3021 14495 3029
rect 13895 2987 14142 3021
rect 14176 2994 14214 3021
rect 13895 2960 14144 2987
rect 14178 2960 14212 2994
rect 14248 2987 14495 3021
rect 14246 2960 14495 2987
rect 13895 2948 14495 2960
rect 13895 2914 14142 2948
rect 14176 2925 14214 2948
rect 13895 2891 14144 2914
rect 14178 2891 14212 2925
rect 14248 2914 14495 2948
rect 14246 2891 14495 2914
rect 13895 2875 14495 2891
rect 13895 2841 14142 2875
rect 14176 2856 14214 2875
rect 13895 2822 14144 2841
rect 14178 2822 14212 2856
rect 14248 2841 14495 2875
rect 14246 2822 14495 2841
rect 13895 2802 14495 2822
rect 13895 2768 14142 2802
rect 14176 2787 14214 2802
rect 13895 2753 14144 2768
rect 14178 2753 14212 2787
rect 14248 2768 14495 2802
rect 14246 2753 14495 2768
rect 13895 2729 14495 2753
rect 13895 2695 14142 2729
rect 14176 2718 14214 2729
rect 13895 2684 14144 2695
rect 14178 2684 14212 2718
rect 14248 2695 14495 2729
rect 14246 2684 14495 2695
rect 13895 2656 14495 2684
rect 13895 2622 14142 2656
rect 14176 2649 14214 2656
rect 13895 2615 14144 2622
rect 14178 2615 14212 2649
rect 14248 2622 14495 2656
rect 14246 2615 14495 2622
rect 13895 2583 14495 2615
rect 13895 2549 14142 2583
rect 14176 2580 14214 2583
rect 13895 2546 14144 2549
rect 14178 2546 14212 2580
rect 14248 2549 14495 2583
rect 14246 2546 14495 2549
rect 13895 2511 14495 2546
rect 13895 2510 14144 2511
rect 13895 2476 14142 2510
rect 14178 2477 14212 2511
rect 14246 2510 14495 2511
rect 14176 2476 14214 2477
rect 14248 2476 14495 2510
rect 13895 2442 14495 2476
rect 13895 2437 14144 2442
rect 13895 2403 14142 2437
rect 14178 2408 14212 2442
rect 14246 2437 14495 2442
rect 14176 2403 14214 2408
rect 14248 2403 14495 2437
rect 13895 2373 14495 2403
rect 13895 2364 14144 2373
rect 13895 2330 14142 2364
rect 14178 2339 14212 2373
rect 14246 2364 14495 2373
rect 14176 2330 14214 2339
rect 14248 2330 14495 2364
rect 13895 2304 14495 2330
rect 13895 2291 14144 2304
rect 13895 2257 14142 2291
rect 14178 2270 14212 2304
rect 14246 2291 14495 2304
rect 14176 2257 14214 2270
rect 14248 2257 14495 2291
rect 13895 2235 14495 2257
rect 13895 2218 14144 2235
rect 13895 2184 14142 2218
rect 14178 2201 14212 2235
rect 14246 2218 14495 2235
rect 14176 2184 14214 2201
rect 14248 2184 14495 2218
rect 13895 2166 14495 2184
rect 13895 2145 14144 2166
rect 13895 2111 14142 2145
rect 14178 2132 14212 2166
rect 14246 2145 14495 2166
rect 14176 2111 14214 2132
rect 14248 2111 14495 2145
rect 13895 2097 14495 2111
rect 13895 2072 14144 2097
rect 13895 2038 14142 2072
rect 14178 2063 14212 2097
rect 14246 2072 14495 2097
rect 14176 2038 14214 2063
rect 14248 2038 14495 2072
rect 13895 2028 14495 2038
rect 13895 1999 14144 2028
rect 13895 1965 14142 1999
rect 14178 1994 14212 2028
rect 14246 1999 14495 2028
rect 14176 1965 14214 1994
rect 14248 1965 14495 1999
rect 13895 1959 14495 1965
rect 13895 1926 14144 1959
rect 13895 1892 14142 1926
rect 14178 1925 14212 1959
rect 14246 1926 14495 1959
rect 14176 1892 14214 1925
rect 14248 1892 14495 1926
rect 13895 1890 14495 1892
rect 13895 1856 14144 1890
rect 14178 1856 14212 1890
rect 14246 1856 14495 1890
rect 13895 1853 14495 1856
rect 13895 1819 14142 1853
rect 14176 1821 14214 1853
rect 13895 1787 14144 1819
rect 14178 1787 14212 1821
rect 14248 1819 14495 1853
rect 14246 1787 14495 1819
rect 13895 1780 14495 1787
rect 13895 1746 14142 1780
rect 14176 1752 14214 1780
rect 13895 1718 14144 1746
rect 14178 1718 14212 1752
rect 14248 1746 14495 1780
rect 14246 1718 14495 1746
rect 13895 1707 14495 1718
rect 13895 1673 14142 1707
rect 14176 1683 14214 1707
rect 13895 1649 14144 1673
rect 14178 1649 14212 1683
rect 14248 1673 14495 1707
rect 14246 1649 14495 1673
rect 13895 1634 14495 1649
rect 13895 1600 14142 1634
rect 14176 1614 14214 1634
rect 13895 1580 14144 1600
rect 14178 1580 14212 1614
rect 14248 1600 14495 1634
rect 14246 1580 14495 1600
rect 13895 1561 14495 1580
rect 13895 1527 14142 1561
rect 14176 1545 14214 1561
rect 13895 1511 14144 1527
rect 14178 1511 14212 1545
rect 14248 1527 14495 1561
rect 14246 1511 14495 1527
rect 13895 1488 14495 1511
rect 13895 1454 14142 1488
rect 14176 1476 14214 1488
rect 13895 1442 14144 1454
rect 14178 1442 14212 1476
rect 14248 1454 14495 1488
rect 14246 1442 14495 1454
rect 13895 1415 14495 1442
rect 13895 1381 14142 1415
rect 14176 1407 14214 1415
rect 13895 1373 14144 1381
rect 14178 1373 14212 1407
rect 14248 1381 14495 1415
rect 14246 1373 14495 1381
rect 13895 1342 14495 1373
rect 13895 1308 14142 1342
rect 14176 1338 14214 1342
rect 13895 1304 14144 1308
rect 14178 1304 14212 1338
rect 14248 1308 14495 1342
rect 14246 1304 14495 1308
rect 13895 1269 14495 1304
rect 13895 1235 14142 1269
rect 14178 1235 14212 1269
rect 14248 1235 14495 1269
rect 13895 1135 14495 1235
rect 14616 1777 14786 1812
rect 14650 1743 14684 1777
rect 14718 1743 14752 1777
rect 14616 1708 14786 1743
rect 14650 1674 14684 1708
rect 14718 1674 14752 1708
rect 14616 1639 14786 1674
rect 14650 1605 14684 1639
rect 14718 1605 14752 1639
rect 14616 1570 14786 1605
rect 14650 1536 14684 1570
rect 14718 1536 14752 1570
rect 14616 1501 14786 1536
rect 14650 1467 14684 1501
rect 14718 1467 14752 1501
rect 14616 1432 14786 1467
rect 14650 1398 14684 1432
rect 14718 1398 14752 1432
rect 14616 1363 14786 1398
rect 14650 1329 14684 1363
rect 14718 1329 14752 1363
rect 14616 1294 14786 1329
rect 14650 1260 14684 1294
rect 14718 1260 14752 1294
rect 14616 1225 14786 1260
rect 14650 1191 14684 1225
rect 14718 1191 14752 1225
rect 14616 1156 14786 1191
rect -4436 1087 -4266 1122
rect -4402 1053 -4368 1087
rect -4334 1053 -4300 1087
rect 14650 1122 14684 1156
rect 14718 1122 14752 1156
rect 14616 1087 14786 1122
rect -4436 1018 -4266 1053
rect -4402 984 -4368 1018
rect -4334 984 -4300 1018
rect -3658 1042 -3524 1058
rect -3658 1020 -3642 1042
rect -3658 992 -3644 1020
rect -3608 1008 -3574 1042
rect -3540 1020 -3524 1042
rect -3610 986 -3572 1008
rect -3538 992 -3524 1020
rect -2366 1042 -2232 1058
rect -2366 1008 -2352 1042
rect -2316 1008 -2282 1042
rect -2246 1008 -2232 1042
rect -2366 992 -2232 1008
rect -1854 1042 -1720 1058
rect -1854 1008 -1840 1042
rect -1804 1008 -1770 1042
rect -1734 1008 -1720 1042
rect -1854 992 -1720 1008
rect -562 1042 -428 1058
rect -562 1008 -548 1042
rect -512 1008 -478 1042
rect -442 1008 -428 1042
rect -562 992 -428 1008
rect -50 1042 84 1058
rect -50 1008 -36 1042
rect 0 1008 34 1042
rect 70 1008 84 1042
rect -50 992 84 1008
rect 1242 1042 1376 1058
rect 1242 1008 1256 1042
rect 1292 1008 1326 1042
rect 1362 1008 1376 1042
rect 1242 992 1376 1008
rect 1754 1042 1888 1058
rect 1754 1008 1768 1042
rect 1804 1008 1838 1042
rect 1874 1008 1888 1042
rect 1754 992 1888 1008
rect 3046 1042 3180 1058
rect 3046 1008 3060 1042
rect 3096 1008 3130 1042
rect 3166 1008 3180 1042
rect 3046 992 3180 1008
rect 3558 1042 3692 1058
rect 3558 1008 3572 1042
rect 3608 1008 3642 1042
rect 3678 1008 3692 1042
rect 3558 992 3692 1008
rect 4850 1042 4984 1058
rect 4850 1008 4864 1042
rect 4900 1008 4934 1042
rect 4970 1008 4984 1042
rect 4850 992 4984 1008
rect 5362 1042 5496 1058
rect 5362 1008 5376 1042
rect 5412 1008 5446 1042
rect 5482 1008 5496 1042
rect 5362 992 5496 1008
rect 6654 1042 6788 1058
rect 6654 1008 6668 1042
rect 6704 1008 6738 1042
rect 6774 1008 6788 1042
rect 6654 992 6788 1008
rect 7166 1042 7300 1058
rect 7166 1008 7180 1042
rect 7216 1008 7250 1042
rect 7286 1008 7300 1042
rect 7166 992 7300 1008
rect 8458 1042 8592 1058
rect 8458 1008 8472 1042
rect 8508 1008 8542 1042
rect 8578 1008 8592 1042
rect 8458 992 8592 1008
rect 8970 1042 9104 1058
rect 8970 1008 8984 1042
rect 9020 1008 9054 1042
rect 9090 1008 9104 1042
rect 8970 992 9104 1008
rect 10262 1042 10396 1058
rect 10262 1008 10276 1042
rect 10312 1008 10346 1042
rect 10382 1008 10396 1042
rect 10262 992 10396 1008
rect 10774 1042 10908 1058
rect 10774 1008 10788 1042
rect 10824 1008 10858 1042
rect 10894 1008 10908 1042
rect 10774 992 10908 1008
rect 12066 1042 12200 1058
rect 12066 1008 12080 1042
rect 12116 1008 12150 1042
rect 12186 1008 12200 1042
rect 12066 992 12200 1008
rect 12578 1042 12712 1058
rect 12578 1008 12592 1042
rect 12628 1008 12662 1042
rect 12698 1008 12712 1042
rect 12578 992 12712 1008
rect 13870 1042 14004 1058
rect 13870 1020 13886 1042
rect 13870 992 13884 1020
rect 13920 1008 13954 1042
rect 13988 1020 14004 1042
rect 13918 986 13956 1008
rect 13990 992 14004 1020
rect 14650 1053 14684 1087
rect 14718 1053 14752 1087
rect 14616 1018 14786 1053
rect -4436 949 -4266 984
rect -4402 915 -4368 949
rect -4334 915 -4300 949
rect -4436 880 -4266 915
rect -4402 846 -4368 880
rect -4334 846 -4300 880
rect -4436 811 -4266 846
rect -4402 777 -4368 811
rect -4334 777 -4300 811
rect -4436 742 -4266 777
rect -4402 708 -4368 742
rect -4334 708 -4300 742
rect -4436 640 -4266 708
rect 14650 984 14684 1018
rect 14718 984 14752 1018
rect 14616 949 14786 984
rect 14650 915 14684 949
rect 14718 915 14752 949
rect 14616 880 14786 915
rect 14650 846 14684 880
rect 14718 846 14752 880
rect 14616 811 14786 846
rect 14650 777 14684 811
rect 14718 777 14752 811
rect 14616 742 14786 777
rect 14650 708 14684 742
rect 14718 708 14752 742
rect 14616 640 14786 708
rect -4436 606 -4368 640
rect -4334 608 -4299 640
rect -4334 606 -4313 608
rect -4265 606 -4230 640
rect -4196 606 -4158 640
rect -4124 606 -4089 640
rect -4055 606 -4020 640
rect -3986 606 -3933 640
rect -3899 606 -3864 640
rect -3830 606 -3795 640
rect -3761 606 -3726 640
rect -3692 606 -3657 640
rect -3623 606 -3588 640
rect -3554 606 -3519 640
rect -3485 606 -3450 640
rect -3416 606 -3381 640
rect -3347 606 -3312 640
rect -3278 606 -3243 640
rect -3209 606 -3174 640
rect -3140 606 -3105 640
rect -3071 606 -3036 640
rect -3002 606 -2967 640
rect -2933 606 -2898 640
rect -2864 606 -2829 640
rect -2795 606 -2760 640
rect -2726 606 -2691 640
rect -2657 606 -2622 640
rect -2588 606 -2553 640
rect -2519 606 -2484 640
rect -2450 606 -2415 640
rect -2381 606 -2346 640
rect -2312 606 -2277 640
rect -2243 606 -2208 640
rect -2174 606 -2139 640
rect -2105 606 -2070 640
rect -2036 606 -2001 640
rect -1967 606 -1932 640
rect -1898 606 -1863 640
rect -1829 606 -1794 640
rect -4436 574 -4313 606
rect -4279 574 -1794 606
rect -4436 572 -1794 574
rect -4436 538 -4368 572
rect -4334 538 -4299 572
rect -4265 538 -4230 572
rect -4196 538 -4158 572
rect -4124 538 -4089 572
rect -4055 538 -4020 572
rect -3986 538 -3933 572
rect -3899 538 -3864 572
rect -3830 538 -3795 572
rect -3761 538 -3726 572
rect -3692 538 -3657 572
rect -3623 538 -3588 572
rect -3554 538 -3519 572
rect -3485 538 -3450 572
rect -3416 538 -3381 572
rect -3347 538 -3312 572
rect -3278 538 -3243 572
rect -3209 538 -3174 572
rect -3140 538 -3105 572
rect -3071 538 -3036 572
rect -3002 538 -2967 572
rect -2933 538 -2898 572
rect -2864 538 -2829 572
rect -2795 538 -2760 572
rect -2726 538 -2691 572
rect -2657 538 -2622 572
rect -2588 538 -2553 572
rect -2519 538 -2484 572
rect -2450 538 -2415 572
rect -2381 538 -2346 572
rect -2312 538 -2277 572
rect -2243 538 -2208 572
rect -2174 538 -2139 572
rect -2105 538 -2070 572
rect -2036 538 -2001 572
rect -1967 538 -1932 572
rect -1898 538 -1863 572
rect -1829 538 -1794 572
rect -4436 504 -1794 538
rect -4436 470 -4368 504
rect -4334 470 -4299 504
rect -4265 470 -4230 504
rect -4196 470 -4158 504
rect -4124 470 -4089 504
rect -4055 470 -4020 504
rect -3986 470 -3933 504
rect -3899 470 -3864 504
rect -3830 470 -3795 504
rect -3761 470 -3726 504
rect -3692 470 -3657 504
rect -3623 470 -3588 504
rect -3554 470 -3519 504
rect -3485 470 -3450 504
rect -3416 470 -3381 504
rect -3347 470 -3312 504
rect -3278 470 -3243 504
rect -3209 470 -3174 504
rect -3140 470 -3105 504
rect -3071 470 -3036 504
rect -3002 470 -2967 504
rect -2933 470 -2898 504
rect -2864 470 -2829 504
rect -2795 470 -2760 504
rect -2726 470 -2691 504
rect -2657 470 -2622 504
rect -2588 470 -2553 504
rect -2519 470 -2484 504
rect -2450 470 -2415 504
rect -2381 470 -2346 504
rect -2312 470 -2277 504
rect -2243 470 -2208 504
rect -2174 470 -2139 504
rect -2105 470 -2070 504
rect -2036 470 -2001 504
rect -1967 470 -1932 504
rect -1898 470 -1863 504
rect -1829 470 -1794 504
rect 824 606 859 640
rect 893 606 928 640
rect 962 606 997 640
rect 1031 606 1066 640
rect 1100 606 1135 640
rect 1169 606 1204 640
rect 1238 606 1273 640
rect 1307 606 1342 640
rect 1376 606 1411 640
rect 1445 606 1480 640
rect 1514 606 1549 640
rect 1583 606 1618 640
rect 1652 606 1687 640
rect 1721 606 1756 640
rect 1790 606 1825 640
rect 1859 606 1894 640
rect 1928 606 1963 640
rect 1997 606 2032 640
rect 2066 606 2101 640
rect 2135 606 2170 640
rect 2204 606 2239 640
rect 2273 606 2308 640
rect 824 572 2308 606
rect 824 538 859 572
rect 893 538 928 572
rect 962 538 997 572
rect 1031 538 1066 572
rect 1100 538 1135 572
rect 1169 538 1204 572
rect 1238 538 1273 572
rect 1307 538 1342 572
rect 1376 538 1411 572
rect 1445 538 1480 572
rect 1514 538 1549 572
rect 1583 538 1618 572
rect 1652 538 1687 572
rect 1721 538 1756 572
rect 1790 538 1825 572
rect 1859 538 1894 572
rect 1928 538 1963 572
rect 1997 538 2032 572
rect 2066 538 2101 572
rect 2135 538 2170 572
rect 2204 538 2239 572
rect 2273 538 2308 572
rect 824 504 2308 538
rect 824 470 859 504
rect 893 470 928 504
rect 962 470 997 504
rect 1031 470 1066 504
rect 1100 470 1135 504
rect 1169 470 1204 504
rect 1238 470 1273 504
rect 1307 470 1342 504
rect 1376 470 1411 504
rect 1445 470 1480 504
rect 1514 470 1549 504
rect 1583 470 1618 504
rect 1652 470 1687 504
rect 1721 470 1756 504
rect 1790 470 1825 504
rect 1859 470 1894 504
rect 1928 470 1963 504
rect 1997 470 2032 504
rect 2066 470 2101 504
rect 2135 470 2170 504
rect 2204 470 2239 504
rect 2273 470 2308 504
rect 14718 470 14786 640
rect 15100 11562 15270 11588
rect 15100 11543 15132 11562
rect 15166 11543 15204 11562
rect 15238 11543 15270 11562
rect 15166 11528 15168 11543
rect 15134 11509 15168 11528
rect 15202 11528 15204 11543
rect 15202 11509 15236 11528
rect 15100 11483 15270 11509
rect 15100 11464 15132 11483
rect 15238 11464 15270 11483
rect 15100 878 15132 890
rect 15166 878 15204 890
rect 15238 878 15270 890
rect 15100 855 15270 878
rect 15134 839 15168 855
rect 15166 821 15168 839
rect 15202 839 15236 855
rect 15202 821 15204 839
rect 15100 805 15132 821
rect 15166 805 15204 821
rect 15238 805 15270 821
rect 15100 786 15270 805
rect 15134 766 15168 786
rect 15166 752 15168 766
rect 15202 766 15236 786
rect 15202 752 15204 766
rect 15100 732 15132 752
rect 15166 732 15204 752
rect 15238 732 15270 752
rect 15100 717 15270 732
rect 15134 693 15168 717
rect 15166 683 15168 693
rect 15202 693 15236 717
rect 15202 683 15204 693
rect 15100 659 15132 683
rect 15166 659 15204 683
rect 15238 659 15270 683
rect 15100 648 15270 659
rect 15134 620 15168 648
rect 15166 614 15168 620
rect 15202 620 15236 648
rect 15202 614 15204 620
rect 15100 586 15132 614
rect 15166 586 15204 614
rect 15238 586 15270 614
rect 15100 579 15270 586
rect 15134 547 15168 579
rect 15166 545 15168 547
rect 15202 547 15236 579
rect 15202 545 15204 547
rect 15100 513 15132 545
rect 15166 513 15204 545
rect 15238 513 15270 545
rect 15100 510 15270 513
rect 15134 476 15168 510
rect 15202 476 15236 510
rect 15100 474 15270 476
rect -4854 440 -4852 441
rect -4886 407 -4852 440
rect -4818 440 -4816 441
rect -4818 407 -4784 440
rect -4920 401 -4750 407
rect -4920 372 -4888 401
rect -4854 372 -4816 401
rect -4782 372 -4750 401
rect -4854 367 -4852 372
rect -4886 338 -4852 367
rect -4818 367 -4816 372
rect -4818 338 -4784 367
rect -4920 270 -4750 338
rect 15100 441 15132 474
rect 15166 441 15204 474
rect 15238 441 15270 474
rect 15166 440 15168 441
rect 15134 407 15168 440
rect 15202 440 15204 441
rect 15202 407 15236 440
rect 15100 401 15270 407
rect 15100 372 15132 401
rect 15166 372 15204 401
rect 15238 372 15270 401
rect 15166 367 15168 372
rect 15134 338 15168 367
rect 15202 367 15204 372
rect 15202 338 15236 367
rect 15100 270 15270 338
rect -4920 236 -4852 270
rect -4818 236 -4783 270
rect -4749 236 -4703 270
rect -4669 236 -4634 270
rect -4600 236 -4565 270
rect -4531 236 -4496 270
rect -4462 236 -4427 270
rect -4393 236 -4358 270
rect -4324 236 -4289 270
rect -4255 236 -4220 270
rect -4186 236 -4151 270
rect -4117 236 -4082 270
rect -4048 236 -4013 270
rect -3979 236 -3913 270
rect -4920 202 -3913 236
rect -4920 168 -4852 202
rect -4818 168 -4783 202
rect -4749 168 -4703 202
rect -4669 168 -4634 202
rect -4600 168 -4565 202
rect -4531 168 -4496 202
rect -4462 168 -4427 202
rect -4393 168 -4358 202
rect -4324 168 -4289 202
rect -4255 168 -4220 202
rect -4186 168 -4151 202
rect -4117 168 -4082 202
rect -4048 168 -4013 202
rect -3979 168 -3913 202
rect -4920 134 -3913 168
rect -4920 100 -4852 134
rect -4818 100 -4783 134
rect -4749 100 -4703 134
rect -4669 100 -4634 134
rect -4600 100 -4565 134
rect -4531 100 -4496 134
rect -4462 100 -4427 134
rect -4393 100 -4358 134
rect -4324 100 -4289 134
rect -4255 100 -4220 134
rect -4186 100 -4151 134
rect -4117 100 -4082 134
rect -4048 100 -4013 134
rect -3979 100 -3913 134
rect -2995 236 -2960 270
rect -2926 236 -2891 270
rect -2857 236 -2822 270
rect -2995 202 -2822 236
rect -2995 168 -2960 202
rect -2926 168 -2891 202
rect -2857 168 -2822 202
rect -2995 134 -2822 168
rect -2995 100 -2960 134
rect -2926 100 -2891 134
rect -2857 100 -2822 134
rect 340 236 375 270
rect 409 236 444 270
rect 478 236 513 270
rect 547 236 582 270
rect 616 236 651 270
rect 685 236 720 270
rect 754 236 789 270
rect 823 236 858 270
rect 892 236 927 270
rect 961 236 996 270
rect 1030 236 1065 270
rect 1099 236 1134 270
rect 1168 236 1203 270
rect 1237 236 1272 270
rect 340 202 1272 236
rect 340 168 375 202
rect 409 168 444 202
rect 478 168 513 202
rect 547 168 582 202
rect 616 168 651 202
rect 685 168 720 202
rect 754 168 789 202
rect 823 168 858 202
rect 892 168 927 202
rect 961 168 996 202
rect 1030 168 1065 202
rect 1099 168 1134 202
rect 1168 168 1203 202
rect 1237 168 1272 202
rect 340 134 1272 168
rect 340 100 375 134
rect 409 100 444 134
rect 478 100 513 134
rect 547 100 582 134
rect 616 100 651 134
rect 685 100 720 134
rect 754 100 789 134
rect 823 100 858 134
rect 892 100 927 134
rect 961 100 996 134
rect 1030 100 1065 134
rect 1099 100 1134 134
rect 1168 100 1203 134
rect 1237 100 1272 134
rect 14974 100 15032 270
rect 15202 100 15270 270
<< viali >>
rect -4888 12726 -4782 12757
rect -4888 12692 -4886 12726
rect -4886 12692 -4852 12726
rect -4852 12692 -4818 12726
rect -4818 12692 -4784 12726
rect -4784 12692 -4782 12726
rect -4888 12650 -4782 12692
rect -4888 12616 -4886 12650
rect -4886 12616 -4852 12650
rect -4852 12616 -4818 12650
rect -4818 12616 -4784 12650
rect -4784 12616 -4782 12650
rect -4888 12574 -4782 12616
rect -4888 11931 -4782 12574
rect -4888 11611 -4782 11861
rect 15132 12726 15238 12757
rect 15132 12692 15134 12726
rect 15134 12692 15168 12726
rect 15168 12692 15202 12726
rect 15202 12692 15236 12726
rect 15236 12692 15238 12726
rect 15132 12650 15238 12692
rect 15132 12616 15134 12650
rect 15134 12616 15168 12650
rect 15168 12616 15202 12650
rect 15202 12616 15236 12650
rect 15236 12616 15238 12650
rect 15132 12574 15238 12616
rect 15132 11931 15238 12574
rect -4888 11543 -4854 11562
rect -4816 11543 -4782 11562
rect -4888 11528 -4886 11543
rect -4886 11528 -4854 11543
rect -4816 11528 -4784 11543
rect -4784 11528 -4782 11543
rect -4888 11464 -4782 11483
rect -4888 5185 -4782 11464
rect -4888 5112 -4854 5146
rect -4816 5112 -4782 5146
rect -4888 5039 -4854 5073
rect -4816 5039 -4782 5073
rect -4888 4966 -4854 5000
rect -4816 4966 -4782 5000
rect -4888 4893 -4854 4927
rect -4816 4893 -4782 4927
rect -4888 4820 -4854 4854
rect -4816 4820 -4782 4854
rect -4888 4747 -4854 4781
rect -4816 4747 -4782 4781
rect -4888 4674 -4854 4708
rect -4816 4674 -4782 4708
rect -4888 4601 -4854 4635
rect -4816 4601 -4782 4635
rect -4888 4528 -4854 4562
rect -4816 4528 -4782 4562
rect -4888 4455 -4854 4489
rect -4816 4455 -4782 4489
rect -4888 4382 -4854 4416
rect -4816 4382 -4782 4416
rect -4888 4309 -4854 4343
rect -4816 4309 -4782 4343
rect -4888 4236 -4854 4270
rect -4816 4236 -4782 4270
rect -4888 4163 -4854 4197
rect -4816 4163 -4782 4197
rect -4888 4090 -4854 4124
rect -4816 4090 -4782 4124
rect -4888 4017 -4854 4051
rect -4816 4017 -4782 4051
rect -4888 3944 -4854 3978
rect -4816 3944 -4782 3978
rect -4888 3871 -4854 3905
rect -4816 3871 -4782 3905
rect -4888 3798 -4854 3832
rect -4816 3798 -4782 3832
rect -4888 3725 -4854 3759
rect -4816 3725 -4782 3759
rect -4888 3652 -4854 3686
rect -4816 3652 -4782 3686
rect -4888 3579 -4854 3613
rect -4816 3579 -4782 3613
rect -4888 3506 -4854 3540
rect -4816 3506 -4782 3540
rect -4888 3433 -4854 3467
rect -4816 3433 -4782 3467
rect -4888 3360 -4854 3394
rect -4816 3360 -4782 3394
rect -4888 3287 -4854 3321
rect -4816 3287 -4782 3321
rect -4888 3214 -4854 3248
rect -4816 3214 -4782 3248
rect -4888 3141 -4854 3175
rect -4816 3141 -4782 3175
rect -4888 3068 -4854 3102
rect -4816 3068 -4782 3102
rect -4888 2995 -4854 3029
rect -4816 2995 -4782 3029
rect -4888 2922 -4854 2956
rect -4816 2922 -4782 2956
rect -4888 2849 -4854 2883
rect -4816 2849 -4782 2883
rect -4888 2776 -4854 2810
rect -4816 2776 -4782 2810
rect -4888 2703 -4854 2737
rect -4816 2703 -4782 2737
rect -4888 2630 -4854 2664
rect -4816 2630 -4782 2664
rect -4888 2557 -4854 2591
rect -4816 2557 -4782 2591
rect -4888 2484 -4854 2518
rect -4816 2484 -4782 2518
rect -4888 2411 -4854 2445
rect -4816 2411 -4782 2445
rect -4888 2338 -4854 2372
rect -4816 2338 -4782 2372
rect -4888 2265 -4854 2299
rect -4816 2265 -4782 2299
rect -4888 2192 -4854 2226
rect -4816 2192 -4782 2226
rect -4888 2119 -4854 2153
rect -4816 2119 -4782 2153
rect -4888 2046 -4854 2080
rect -4816 2046 -4782 2080
rect -4888 1973 -4854 2007
rect -4816 1973 -4782 2007
rect -4888 1900 -4854 1934
rect -4816 1900 -4782 1934
rect -4888 1827 -4854 1861
rect -4816 1827 -4782 1861
rect -4888 1754 -4854 1788
rect -4816 1754 -4782 1788
rect -4888 1681 -4854 1715
rect -4816 1681 -4782 1715
rect -4888 1608 -4854 1642
rect -4816 1608 -4782 1642
rect -4888 1535 -4854 1569
rect -4816 1535 -4782 1569
rect -4888 1462 -4854 1496
rect -4816 1462 -4782 1496
rect -4888 1389 -4854 1423
rect -4816 1389 -4782 1423
rect -4888 1316 -4854 1350
rect -4816 1316 -4782 1350
rect -4888 1243 -4854 1277
rect -4816 1243 -4782 1277
rect -4888 1170 -4854 1204
rect -4816 1170 -4782 1204
rect -4888 1097 -4854 1131
rect -4816 1097 -4782 1131
rect -4888 1024 -4854 1058
rect -4816 1024 -4782 1058
rect -4888 951 -4854 985
rect -4816 951 -4782 985
rect -4888 890 -4854 912
rect -4816 890 -4782 912
rect -4888 878 -4854 890
rect -4816 878 -4782 890
rect -4888 821 -4886 839
rect -4886 821 -4854 839
rect -4816 821 -4784 839
rect -4784 821 -4782 839
rect -4888 805 -4854 821
rect -4816 805 -4782 821
rect -4888 752 -4886 766
rect -4886 752 -4854 766
rect -4816 752 -4784 766
rect -4784 752 -4782 766
rect -4888 732 -4854 752
rect -4816 732 -4782 752
rect -4888 683 -4886 693
rect -4886 683 -4854 693
rect -4816 683 -4784 693
rect -4784 683 -4782 693
rect -4888 659 -4854 683
rect -4816 659 -4782 683
rect -4888 614 -4886 620
rect -4886 614 -4854 620
rect -4816 614 -4784 620
rect -4784 614 -4782 620
rect -4888 586 -4854 614
rect -4816 586 -4782 614
rect -4888 545 -4886 547
rect -4886 545 -4854 547
rect -4816 545 -4784 547
rect -4784 545 -4782 547
rect -4888 513 -4854 545
rect -4816 513 -4782 545
rect -4888 441 -4854 474
rect -4816 441 -4782 474
rect -3898 3719 -3896 11233
rect -3896 3719 -3794 11233
rect -3794 3719 -3792 11233
rect -3898 3684 -3792 3719
rect -3898 3650 -3896 3684
rect -3896 3650 -3862 3684
rect -3862 3650 -3828 3684
rect -3828 3650 -3794 3684
rect -3794 3650 -3792 3684
rect -3898 3615 -3792 3650
rect -3898 3581 -3896 3615
rect -3896 3581 -3862 3615
rect -3862 3581 -3828 3615
rect -3828 3581 -3794 3615
rect -3794 3581 -3792 3615
rect -3898 3546 -3792 3581
rect -3898 3512 -3896 3546
rect -3896 3512 -3862 3546
rect -3862 3512 -3828 3546
rect -3828 3512 -3794 3546
rect -3794 3512 -3792 3546
rect -3898 3477 -3792 3512
rect -3898 3443 -3896 3477
rect -3896 3443 -3862 3477
rect -3862 3443 -3828 3477
rect -3828 3443 -3794 3477
rect -3794 3443 -3792 3477
rect -3898 3408 -3792 3443
rect -3898 3374 -3896 3408
rect -3896 3374 -3862 3408
rect -3862 3374 -3828 3408
rect -3828 3374 -3794 3408
rect -3794 3374 -3792 3408
rect -3898 3339 -3792 3374
rect -3898 3305 -3896 3339
rect -3896 3305 -3862 3339
rect -3862 3305 -3828 3339
rect -3828 3305 -3794 3339
rect -3794 3305 -3792 3339
rect -3898 3279 -3792 3305
rect -3898 3236 -3896 3240
rect -3896 3236 -3864 3240
rect -3826 3236 -3794 3240
rect -3794 3236 -3792 3240
rect -3898 3206 -3864 3236
rect -3826 3206 -3792 3236
rect -3898 3133 -3864 3167
rect -3826 3133 -3792 3167
rect -3898 3063 -3864 3094
rect -3826 3063 -3792 3094
rect -3898 3060 -3896 3063
rect -3896 3060 -3864 3063
rect -3826 3060 -3794 3063
rect -3794 3060 -3792 3063
rect -3898 2994 -3864 3021
rect -3826 2994 -3792 3021
rect -3898 2987 -3896 2994
rect -3896 2987 -3864 2994
rect -3826 2987 -3794 2994
rect -3794 2987 -3792 2994
rect -3898 2925 -3864 2948
rect -3826 2925 -3792 2948
rect -3898 2914 -3896 2925
rect -3896 2914 -3864 2925
rect -3826 2914 -3794 2925
rect -3794 2914 -3792 2925
rect -3898 2856 -3864 2875
rect -3826 2856 -3792 2875
rect -3898 2841 -3896 2856
rect -3896 2841 -3864 2856
rect -3826 2841 -3794 2856
rect -3794 2841 -3792 2856
rect -3898 2787 -3864 2802
rect -3826 2787 -3792 2802
rect -3898 2768 -3896 2787
rect -3896 2768 -3864 2787
rect -3826 2768 -3794 2787
rect -3794 2768 -3792 2787
rect -3898 2718 -3864 2729
rect -3826 2718 -3792 2729
rect -3898 2695 -3896 2718
rect -3896 2695 -3864 2718
rect -3826 2695 -3794 2718
rect -3794 2695 -3792 2718
rect -3898 2649 -3864 2656
rect -3826 2649 -3792 2656
rect -3898 2622 -3896 2649
rect -3896 2622 -3864 2649
rect -3826 2622 -3794 2649
rect -3794 2622 -3792 2649
rect -3898 2580 -3864 2583
rect -3826 2580 -3792 2583
rect -3898 2549 -3896 2580
rect -3896 2549 -3864 2580
rect -3826 2549 -3794 2580
rect -3794 2549 -3792 2580
rect -3898 2477 -3896 2510
rect -3896 2477 -3864 2510
rect -3826 2477 -3794 2510
rect -3794 2477 -3792 2510
rect -3898 2476 -3864 2477
rect -3826 2476 -3792 2477
rect -3898 2408 -3896 2437
rect -3896 2408 -3864 2437
rect -3826 2408 -3794 2437
rect -3794 2408 -3792 2437
rect -3898 2403 -3864 2408
rect -3826 2403 -3792 2408
rect -3898 2339 -3896 2364
rect -3896 2339 -3864 2364
rect -3826 2339 -3794 2364
rect -3794 2339 -3792 2364
rect -3898 2330 -3864 2339
rect -3826 2330 -3792 2339
rect -3898 2270 -3896 2291
rect -3896 2270 -3864 2291
rect -3826 2270 -3794 2291
rect -3794 2270 -3792 2291
rect -3898 2257 -3864 2270
rect -3826 2257 -3792 2270
rect -3898 2201 -3896 2218
rect -3896 2201 -3864 2218
rect -3826 2201 -3794 2218
rect -3794 2201 -3792 2218
rect -3898 2184 -3864 2201
rect -3826 2184 -3792 2201
rect -3898 2132 -3896 2145
rect -3896 2132 -3864 2145
rect -3826 2132 -3794 2145
rect -3794 2132 -3792 2145
rect -3898 2111 -3864 2132
rect -3826 2111 -3792 2132
rect -3898 2063 -3896 2072
rect -3896 2063 -3864 2072
rect -3826 2063 -3794 2072
rect -3794 2063 -3792 2072
rect -3898 2038 -3864 2063
rect -3826 2038 -3792 2063
rect -3898 1994 -3896 1999
rect -3896 1994 -3864 1999
rect -3826 1994 -3794 1999
rect -3794 1994 -3792 1999
rect -3898 1965 -3864 1994
rect -3826 1965 -3792 1994
rect -3898 1925 -3896 1926
rect -3896 1925 -3864 1926
rect -3826 1925 -3794 1926
rect -3794 1925 -3792 1926
rect -3898 1892 -3864 1925
rect -3826 1892 -3792 1925
rect -3898 1821 -3864 1853
rect -3826 1821 -3792 1853
rect -3898 1819 -3896 1821
rect -3896 1819 -3864 1821
rect -3826 1819 -3794 1821
rect -3794 1819 -3792 1821
rect -3898 1752 -3864 1780
rect -3826 1752 -3792 1780
rect -3898 1746 -3896 1752
rect -3896 1746 -3864 1752
rect -3826 1746 -3794 1752
rect -3794 1746 -3792 1752
rect -3898 1683 -3864 1707
rect -3826 1683 -3792 1707
rect -3898 1673 -3896 1683
rect -3896 1673 -3864 1683
rect -3826 1673 -3794 1683
rect -3794 1673 -3792 1683
rect -3898 1614 -3864 1634
rect -3826 1614 -3792 1634
rect -3898 1600 -3896 1614
rect -3896 1600 -3864 1614
rect -3826 1600 -3794 1614
rect -3794 1600 -3792 1614
rect -3898 1545 -3864 1561
rect -3826 1545 -3792 1561
rect -3898 1527 -3896 1545
rect -3896 1527 -3864 1545
rect -3826 1527 -3794 1545
rect -3794 1527 -3792 1545
rect -3898 1476 -3864 1488
rect -3826 1476 -3792 1488
rect -3898 1454 -3896 1476
rect -3896 1454 -3864 1476
rect -3826 1454 -3794 1476
rect -3794 1454 -3792 1476
rect -3898 1407 -3864 1415
rect -3826 1407 -3792 1415
rect -3898 1381 -3896 1407
rect -3896 1381 -3864 1407
rect -3826 1381 -3794 1407
rect -3794 1381 -3792 1407
rect -3898 1338 -3864 1342
rect -3826 1338 -3792 1342
rect -3898 1308 -3896 1338
rect -3896 1308 -3864 1338
rect -3826 1308 -3794 1338
rect -3794 1308 -3792 1338
rect -3898 1235 -3896 1269
rect -3896 1235 -3864 1269
rect -3826 1235 -3794 1269
rect -3794 1235 -3792 1269
rect -2996 3719 -2994 11233
rect -2994 3719 -2892 11233
rect -2892 3719 -2890 11233
rect -2996 3684 -2890 3719
rect -2996 3650 -2994 3684
rect -2994 3650 -2960 3684
rect -2960 3650 -2926 3684
rect -2926 3650 -2892 3684
rect -2892 3650 -2890 3684
rect -2996 3615 -2890 3650
rect -2996 3581 -2994 3615
rect -2994 3581 -2960 3615
rect -2960 3581 -2926 3615
rect -2926 3581 -2892 3615
rect -2892 3581 -2890 3615
rect -2996 3546 -2890 3581
rect -2996 3512 -2994 3546
rect -2994 3512 -2960 3546
rect -2960 3512 -2926 3546
rect -2926 3512 -2892 3546
rect -2892 3512 -2890 3546
rect -2996 3477 -2890 3512
rect -2996 3443 -2994 3477
rect -2994 3443 -2960 3477
rect -2960 3443 -2926 3477
rect -2926 3443 -2892 3477
rect -2892 3443 -2890 3477
rect -2996 3408 -2890 3443
rect -2996 3374 -2994 3408
rect -2994 3374 -2960 3408
rect -2960 3374 -2926 3408
rect -2926 3374 -2892 3408
rect -2892 3374 -2890 3408
rect -2996 3339 -2890 3374
rect -2996 3305 -2994 3339
rect -2994 3305 -2960 3339
rect -2960 3305 -2926 3339
rect -2926 3305 -2892 3339
rect -2892 3305 -2890 3339
rect -2996 3279 -2890 3305
rect -2996 3236 -2994 3240
rect -2994 3236 -2962 3240
rect -2924 3236 -2892 3240
rect -2892 3236 -2890 3240
rect -2996 3206 -2962 3236
rect -2924 3206 -2890 3236
rect -2996 3133 -2962 3167
rect -2924 3133 -2890 3167
rect -2996 3063 -2962 3094
rect -2924 3063 -2890 3094
rect -2996 3060 -2994 3063
rect -2994 3060 -2962 3063
rect -2924 3060 -2892 3063
rect -2892 3060 -2890 3063
rect -2996 2994 -2962 3021
rect -2924 2994 -2890 3021
rect -2996 2987 -2994 2994
rect -2994 2987 -2962 2994
rect -2924 2987 -2892 2994
rect -2892 2987 -2890 2994
rect -2996 2925 -2962 2948
rect -2924 2925 -2890 2948
rect -2996 2914 -2994 2925
rect -2994 2914 -2962 2925
rect -2924 2914 -2892 2925
rect -2892 2914 -2890 2925
rect -2996 2856 -2962 2875
rect -2924 2856 -2890 2875
rect -2996 2841 -2994 2856
rect -2994 2841 -2962 2856
rect -2924 2841 -2892 2856
rect -2892 2841 -2890 2856
rect -2996 2787 -2962 2802
rect -2924 2787 -2890 2802
rect -2996 2768 -2994 2787
rect -2994 2768 -2962 2787
rect -2924 2768 -2892 2787
rect -2892 2768 -2890 2787
rect -2996 2718 -2962 2729
rect -2924 2718 -2890 2729
rect -2996 2695 -2994 2718
rect -2994 2695 -2962 2718
rect -2924 2695 -2892 2718
rect -2892 2695 -2890 2718
rect -2996 2649 -2962 2656
rect -2924 2649 -2890 2656
rect -2996 2622 -2994 2649
rect -2994 2622 -2962 2649
rect -2924 2622 -2892 2649
rect -2892 2622 -2890 2649
rect -2996 2580 -2962 2583
rect -2924 2580 -2890 2583
rect -2996 2549 -2994 2580
rect -2994 2549 -2962 2580
rect -2924 2549 -2892 2580
rect -2892 2549 -2890 2580
rect -2996 2477 -2994 2510
rect -2994 2477 -2962 2510
rect -2924 2477 -2892 2510
rect -2892 2477 -2890 2510
rect -2996 2476 -2962 2477
rect -2924 2476 -2890 2477
rect -2996 2408 -2994 2437
rect -2994 2408 -2962 2437
rect -2924 2408 -2892 2437
rect -2892 2408 -2890 2437
rect -2996 2403 -2962 2408
rect -2924 2403 -2890 2408
rect -2996 2339 -2994 2364
rect -2994 2339 -2962 2364
rect -2924 2339 -2892 2364
rect -2892 2339 -2890 2364
rect -2996 2330 -2962 2339
rect -2924 2330 -2890 2339
rect -2996 2270 -2994 2291
rect -2994 2270 -2962 2291
rect -2924 2270 -2892 2291
rect -2892 2270 -2890 2291
rect -2996 2257 -2962 2270
rect -2924 2257 -2890 2270
rect -2996 2201 -2994 2218
rect -2994 2201 -2962 2218
rect -2924 2201 -2892 2218
rect -2892 2201 -2890 2218
rect -2996 2184 -2962 2201
rect -2924 2184 -2890 2201
rect -2996 2132 -2994 2145
rect -2994 2132 -2962 2145
rect -2924 2132 -2892 2145
rect -2892 2132 -2890 2145
rect -2996 2111 -2962 2132
rect -2924 2111 -2890 2132
rect -2996 2063 -2994 2072
rect -2994 2063 -2962 2072
rect -2924 2063 -2892 2072
rect -2892 2063 -2890 2072
rect -2996 2038 -2962 2063
rect -2924 2038 -2890 2063
rect -2996 1994 -2994 1999
rect -2994 1994 -2962 1999
rect -2924 1994 -2892 1999
rect -2892 1994 -2890 1999
rect -2996 1965 -2962 1994
rect -2924 1965 -2890 1994
rect -2996 1925 -2994 1926
rect -2994 1925 -2962 1926
rect -2924 1925 -2892 1926
rect -2892 1925 -2890 1926
rect -2996 1892 -2962 1925
rect -2924 1892 -2890 1925
rect -2996 1821 -2962 1853
rect -2924 1821 -2890 1853
rect -2996 1819 -2994 1821
rect -2994 1819 -2962 1821
rect -2924 1819 -2892 1821
rect -2892 1819 -2890 1821
rect -2996 1752 -2962 1780
rect -2924 1752 -2890 1780
rect -2996 1746 -2994 1752
rect -2994 1746 -2962 1752
rect -2924 1746 -2892 1752
rect -2892 1746 -2890 1752
rect -2996 1683 -2962 1707
rect -2924 1683 -2890 1707
rect -2996 1673 -2994 1683
rect -2994 1673 -2962 1683
rect -2924 1673 -2892 1683
rect -2892 1673 -2890 1683
rect -2996 1614 -2962 1634
rect -2924 1614 -2890 1634
rect -2996 1600 -2994 1614
rect -2994 1600 -2962 1614
rect -2924 1600 -2892 1614
rect -2892 1600 -2890 1614
rect -2996 1545 -2962 1561
rect -2924 1545 -2890 1561
rect -2996 1527 -2994 1545
rect -2994 1527 -2962 1545
rect -2924 1527 -2892 1545
rect -2892 1527 -2890 1545
rect -2996 1476 -2962 1488
rect -2924 1476 -2890 1488
rect -2996 1454 -2994 1476
rect -2994 1454 -2962 1476
rect -2924 1454 -2892 1476
rect -2892 1454 -2890 1476
rect -2996 1407 -2962 1415
rect -2924 1407 -2890 1415
rect -2996 1381 -2994 1407
rect -2994 1381 -2962 1407
rect -2924 1381 -2892 1407
rect -2892 1381 -2890 1407
rect -2996 1338 -2962 1342
rect -2924 1338 -2890 1342
rect -2996 1308 -2994 1338
rect -2994 1308 -2962 1338
rect -2924 1308 -2892 1338
rect -2892 1308 -2890 1338
rect -2996 1235 -2994 1269
rect -2994 1235 -2962 1269
rect -2924 1235 -2892 1269
rect -2892 1235 -2890 1269
rect -2094 3719 -2092 11233
rect -2092 3719 -1990 11233
rect -1990 3719 -1988 11233
rect -2094 3684 -1988 3719
rect -2094 3650 -2092 3684
rect -2092 3650 -2058 3684
rect -2058 3650 -2024 3684
rect -2024 3650 -1990 3684
rect -1990 3650 -1988 3684
rect -2094 3615 -1988 3650
rect -2094 3581 -2092 3615
rect -2092 3581 -2058 3615
rect -2058 3581 -2024 3615
rect -2024 3581 -1990 3615
rect -1990 3581 -1988 3615
rect -2094 3546 -1988 3581
rect -2094 3512 -2092 3546
rect -2092 3512 -2058 3546
rect -2058 3512 -2024 3546
rect -2024 3512 -1990 3546
rect -1990 3512 -1988 3546
rect -2094 3477 -1988 3512
rect -2094 3443 -2092 3477
rect -2092 3443 -2058 3477
rect -2058 3443 -2024 3477
rect -2024 3443 -1990 3477
rect -1990 3443 -1988 3477
rect -2094 3408 -1988 3443
rect -2094 3374 -2092 3408
rect -2092 3374 -2058 3408
rect -2058 3374 -2024 3408
rect -2024 3374 -1990 3408
rect -1990 3374 -1988 3408
rect -2094 3339 -1988 3374
rect -2094 3305 -2092 3339
rect -2092 3305 -2058 3339
rect -2058 3305 -2024 3339
rect -2024 3305 -1990 3339
rect -1990 3305 -1988 3339
rect -2094 3279 -1988 3305
rect -2094 3236 -2092 3240
rect -2092 3236 -2060 3240
rect -2022 3236 -1990 3240
rect -1990 3236 -1988 3240
rect -2094 3206 -2060 3236
rect -2022 3206 -1988 3236
rect -2094 3133 -2060 3167
rect -2022 3133 -1988 3167
rect -2094 3063 -2060 3094
rect -2022 3063 -1988 3094
rect -2094 3060 -2092 3063
rect -2092 3060 -2060 3063
rect -2022 3060 -1990 3063
rect -1990 3060 -1988 3063
rect -2094 2994 -2060 3021
rect -2022 2994 -1988 3021
rect -2094 2987 -2092 2994
rect -2092 2987 -2060 2994
rect -2022 2987 -1990 2994
rect -1990 2987 -1988 2994
rect -2094 2925 -2060 2948
rect -2022 2925 -1988 2948
rect -2094 2914 -2092 2925
rect -2092 2914 -2060 2925
rect -2022 2914 -1990 2925
rect -1990 2914 -1988 2925
rect -2094 2856 -2060 2875
rect -2022 2856 -1988 2875
rect -2094 2841 -2092 2856
rect -2092 2841 -2060 2856
rect -2022 2841 -1990 2856
rect -1990 2841 -1988 2856
rect -2094 2787 -2060 2802
rect -2022 2787 -1988 2802
rect -2094 2768 -2092 2787
rect -2092 2768 -2060 2787
rect -2022 2768 -1990 2787
rect -1990 2768 -1988 2787
rect -2094 2718 -2060 2729
rect -2022 2718 -1988 2729
rect -2094 2695 -2092 2718
rect -2092 2695 -2060 2718
rect -2022 2695 -1990 2718
rect -1990 2695 -1988 2718
rect -2094 2649 -2060 2656
rect -2022 2649 -1988 2656
rect -2094 2622 -2092 2649
rect -2092 2622 -2060 2649
rect -2022 2622 -1990 2649
rect -1990 2622 -1988 2649
rect -2094 2580 -2060 2583
rect -2022 2580 -1988 2583
rect -2094 2549 -2092 2580
rect -2092 2549 -2060 2580
rect -2022 2549 -1990 2580
rect -1990 2549 -1988 2580
rect -2094 2477 -2092 2510
rect -2092 2477 -2060 2510
rect -2022 2477 -1990 2510
rect -1990 2477 -1988 2510
rect -2094 2476 -2060 2477
rect -2022 2476 -1988 2477
rect -2094 2408 -2092 2437
rect -2092 2408 -2060 2437
rect -2022 2408 -1990 2437
rect -1990 2408 -1988 2437
rect -2094 2403 -2060 2408
rect -2022 2403 -1988 2408
rect -2094 2339 -2092 2364
rect -2092 2339 -2060 2364
rect -2022 2339 -1990 2364
rect -1990 2339 -1988 2364
rect -2094 2330 -2060 2339
rect -2022 2330 -1988 2339
rect -2094 2270 -2092 2291
rect -2092 2270 -2060 2291
rect -2022 2270 -1990 2291
rect -1990 2270 -1988 2291
rect -2094 2257 -2060 2270
rect -2022 2257 -1988 2270
rect -2094 2201 -2092 2218
rect -2092 2201 -2060 2218
rect -2022 2201 -1990 2218
rect -1990 2201 -1988 2218
rect -2094 2184 -2060 2201
rect -2022 2184 -1988 2201
rect -2094 2132 -2092 2145
rect -2092 2132 -2060 2145
rect -2022 2132 -1990 2145
rect -1990 2132 -1988 2145
rect -2094 2111 -2060 2132
rect -2022 2111 -1988 2132
rect -2094 2063 -2092 2072
rect -2092 2063 -2060 2072
rect -2022 2063 -1990 2072
rect -1990 2063 -1988 2072
rect -2094 2038 -2060 2063
rect -2022 2038 -1988 2063
rect -2094 1994 -2092 1999
rect -2092 1994 -2060 1999
rect -2022 1994 -1990 1999
rect -1990 1994 -1988 1999
rect -2094 1965 -2060 1994
rect -2022 1965 -1988 1994
rect -2094 1925 -2092 1926
rect -2092 1925 -2060 1926
rect -2022 1925 -1990 1926
rect -1990 1925 -1988 1926
rect -2094 1892 -2060 1925
rect -2022 1892 -1988 1925
rect -2094 1821 -2060 1853
rect -2022 1821 -1988 1853
rect -2094 1819 -2092 1821
rect -2092 1819 -2060 1821
rect -2022 1819 -1990 1821
rect -1990 1819 -1988 1821
rect -2094 1752 -2060 1780
rect -2022 1752 -1988 1780
rect -2094 1746 -2092 1752
rect -2092 1746 -2060 1752
rect -2022 1746 -1990 1752
rect -1990 1746 -1988 1752
rect -2094 1683 -2060 1707
rect -2022 1683 -1988 1707
rect -2094 1673 -2092 1683
rect -2092 1673 -2060 1683
rect -2022 1673 -1990 1683
rect -1990 1673 -1988 1683
rect -2094 1614 -2060 1634
rect -2022 1614 -1988 1634
rect -2094 1600 -2092 1614
rect -2092 1600 -2060 1614
rect -2022 1600 -1990 1614
rect -1990 1600 -1988 1614
rect -2094 1545 -2060 1561
rect -2022 1545 -1988 1561
rect -2094 1527 -2092 1545
rect -2092 1527 -2060 1545
rect -2022 1527 -1990 1545
rect -1990 1527 -1988 1545
rect -2094 1476 -2060 1488
rect -2022 1476 -1988 1488
rect -2094 1454 -2092 1476
rect -2092 1454 -2060 1476
rect -2022 1454 -1990 1476
rect -1990 1454 -1988 1476
rect -2094 1407 -2060 1415
rect -2022 1407 -1988 1415
rect -2094 1381 -2092 1407
rect -2092 1381 -2060 1407
rect -2022 1381 -1990 1407
rect -1990 1381 -1988 1407
rect -2094 1338 -2060 1342
rect -2022 1338 -1988 1342
rect -2094 1308 -2092 1338
rect -2092 1308 -2060 1338
rect -2022 1308 -1990 1338
rect -1990 1308 -1988 1338
rect -2094 1235 -2092 1269
rect -2092 1235 -2060 1269
rect -2022 1235 -1990 1269
rect -1990 1235 -1988 1269
rect -1192 3719 -1190 11233
rect -1190 3719 -1088 11233
rect -1088 3719 -1086 11233
rect -1192 3684 -1086 3719
rect -1192 3650 -1190 3684
rect -1190 3650 -1156 3684
rect -1156 3650 -1122 3684
rect -1122 3650 -1088 3684
rect -1088 3650 -1086 3684
rect -1192 3615 -1086 3650
rect -1192 3581 -1190 3615
rect -1190 3581 -1156 3615
rect -1156 3581 -1122 3615
rect -1122 3581 -1088 3615
rect -1088 3581 -1086 3615
rect -1192 3546 -1086 3581
rect -1192 3512 -1190 3546
rect -1190 3512 -1156 3546
rect -1156 3512 -1122 3546
rect -1122 3512 -1088 3546
rect -1088 3512 -1086 3546
rect -1192 3477 -1086 3512
rect -1192 3443 -1190 3477
rect -1190 3443 -1156 3477
rect -1156 3443 -1122 3477
rect -1122 3443 -1088 3477
rect -1088 3443 -1086 3477
rect -1192 3408 -1086 3443
rect -1192 3374 -1190 3408
rect -1190 3374 -1156 3408
rect -1156 3374 -1122 3408
rect -1122 3374 -1088 3408
rect -1088 3374 -1086 3408
rect -1192 3339 -1086 3374
rect -1192 3305 -1190 3339
rect -1190 3305 -1156 3339
rect -1156 3305 -1122 3339
rect -1122 3305 -1088 3339
rect -1088 3305 -1086 3339
rect -1192 3279 -1086 3305
rect -1192 3236 -1190 3240
rect -1190 3236 -1158 3240
rect -1120 3236 -1088 3240
rect -1088 3236 -1086 3240
rect -1192 3206 -1158 3236
rect -1120 3206 -1086 3236
rect -1192 3133 -1158 3167
rect -1120 3133 -1086 3167
rect -1192 3063 -1158 3094
rect -1120 3063 -1086 3094
rect -1192 3060 -1190 3063
rect -1190 3060 -1158 3063
rect -1120 3060 -1088 3063
rect -1088 3060 -1086 3063
rect -1192 2994 -1158 3021
rect -1120 2994 -1086 3021
rect -1192 2987 -1190 2994
rect -1190 2987 -1158 2994
rect -1120 2987 -1088 2994
rect -1088 2987 -1086 2994
rect -1192 2925 -1158 2948
rect -1120 2925 -1086 2948
rect -1192 2914 -1190 2925
rect -1190 2914 -1158 2925
rect -1120 2914 -1088 2925
rect -1088 2914 -1086 2925
rect -1192 2856 -1158 2875
rect -1120 2856 -1086 2875
rect -1192 2841 -1190 2856
rect -1190 2841 -1158 2856
rect -1120 2841 -1088 2856
rect -1088 2841 -1086 2856
rect -1192 2787 -1158 2802
rect -1120 2787 -1086 2802
rect -1192 2768 -1190 2787
rect -1190 2768 -1158 2787
rect -1120 2768 -1088 2787
rect -1088 2768 -1086 2787
rect -1192 2718 -1158 2729
rect -1120 2718 -1086 2729
rect -1192 2695 -1190 2718
rect -1190 2695 -1158 2718
rect -1120 2695 -1088 2718
rect -1088 2695 -1086 2718
rect -1192 2649 -1158 2656
rect -1120 2649 -1086 2656
rect -1192 2622 -1190 2649
rect -1190 2622 -1158 2649
rect -1120 2622 -1088 2649
rect -1088 2622 -1086 2649
rect -1192 2580 -1158 2583
rect -1120 2580 -1086 2583
rect -1192 2549 -1190 2580
rect -1190 2549 -1158 2580
rect -1120 2549 -1088 2580
rect -1088 2549 -1086 2580
rect -1192 2477 -1190 2510
rect -1190 2477 -1158 2510
rect -1120 2477 -1088 2510
rect -1088 2477 -1086 2510
rect -1192 2476 -1158 2477
rect -1120 2476 -1086 2477
rect -1192 2408 -1190 2437
rect -1190 2408 -1158 2437
rect -1120 2408 -1088 2437
rect -1088 2408 -1086 2437
rect -1192 2403 -1158 2408
rect -1120 2403 -1086 2408
rect -1192 2339 -1190 2364
rect -1190 2339 -1158 2364
rect -1120 2339 -1088 2364
rect -1088 2339 -1086 2364
rect -1192 2330 -1158 2339
rect -1120 2330 -1086 2339
rect -1192 2270 -1190 2291
rect -1190 2270 -1158 2291
rect -1120 2270 -1088 2291
rect -1088 2270 -1086 2291
rect -1192 2257 -1158 2270
rect -1120 2257 -1086 2270
rect -1192 2201 -1190 2218
rect -1190 2201 -1158 2218
rect -1120 2201 -1088 2218
rect -1088 2201 -1086 2218
rect -1192 2184 -1158 2201
rect -1120 2184 -1086 2201
rect -1192 2132 -1190 2145
rect -1190 2132 -1158 2145
rect -1120 2132 -1088 2145
rect -1088 2132 -1086 2145
rect -1192 2111 -1158 2132
rect -1120 2111 -1086 2132
rect -1192 2063 -1190 2072
rect -1190 2063 -1158 2072
rect -1120 2063 -1088 2072
rect -1088 2063 -1086 2072
rect -1192 2038 -1158 2063
rect -1120 2038 -1086 2063
rect -1192 1994 -1190 1999
rect -1190 1994 -1158 1999
rect -1120 1994 -1088 1999
rect -1088 1994 -1086 1999
rect -1192 1965 -1158 1994
rect -1120 1965 -1086 1994
rect -1192 1925 -1190 1926
rect -1190 1925 -1158 1926
rect -1120 1925 -1088 1926
rect -1088 1925 -1086 1926
rect -1192 1892 -1158 1925
rect -1120 1892 -1086 1925
rect -1192 1821 -1158 1853
rect -1120 1821 -1086 1853
rect -1192 1819 -1190 1821
rect -1190 1819 -1158 1821
rect -1120 1819 -1088 1821
rect -1088 1819 -1086 1821
rect -1192 1752 -1158 1780
rect -1120 1752 -1086 1780
rect -1192 1746 -1190 1752
rect -1190 1746 -1158 1752
rect -1120 1746 -1088 1752
rect -1088 1746 -1086 1752
rect -1192 1683 -1158 1707
rect -1120 1683 -1086 1707
rect -1192 1673 -1190 1683
rect -1190 1673 -1158 1683
rect -1120 1673 -1088 1683
rect -1088 1673 -1086 1683
rect -1192 1614 -1158 1634
rect -1120 1614 -1086 1634
rect -1192 1600 -1190 1614
rect -1190 1600 -1158 1614
rect -1120 1600 -1088 1614
rect -1088 1600 -1086 1614
rect -1192 1545 -1158 1561
rect -1120 1545 -1086 1561
rect -1192 1527 -1190 1545
rect -1190 1527 -1158 1545
rect -1120 1527 -1088 1545
rect -1088 1527 -1086 1545
rect -1192 1476 -1158 1488
rect -1120 1476 -1086 1488
rect -1192 1454 -1190 1476
rect -1190 1454 -1158 1476
rect -1120 1454 -1088 1476
rect -1088 1454 -1086 1476
rect -1192 1407 -1158 1415
rect -1120 1407 -1086 1415
rect -1192 1381 -1190 1407
rect -1190 1381 -1158 1407
rect -1120 1381 -1088 1407
rect -1088 1381 -1086 1407
rect -1192 1338 -1158 1342
rect -1120 1338 -1086 1342
rect -1192 1308 -1190 1338
rect -1190 1308 -1158 1338
rect -1120 1308 -1088 1338
rect -1088 1308 -1086 1338
rect -1192 1235 -1190 1269
rect -1190 1235 -1158 1269
rect -1120 1235 -1088 1269
rect -1088 1235 -1086 1269
rect -290 3719 -288 11233
rect -288 3719 -186 11233
rect -186 3719 -184 11233
rect -290 3684 -184 3719
rect -290 3650 -288 3684
rect -288 3650 -254 3684
rect -254 3650 -220 3684
rect -220 3650 -186 3684
rect -186 3650 -184 3684
rect -290 3615 -184 3650
rect -290 3581 -288 3615
rect -288 3581 -254 3615
rect -254 3581 -220 3615
rect -220 3581 -186 3615
rect -186 3581 -184 3615
rect -290 3546 -184 3581
rect -290 3512 -288 3546
rect -288 3512 -254 3546
rect -254 3512 -220 3546
rect -220 3512 -186 3546
rect -186 3512 -184 3546
rect -290 3477 -184 3512
rect -290 3443 -288 3477
rect -288 3443 -254 3477
rect -254 3443 -220 3477
rect -220 3443 -186 3477
rect -186 3443 -184 3477
rect -290 3408 -184 3443
rect -290 3374 -288 3408
rect -288 3374 -254 3408
rect -254 3374 -220 3408
rect -220 3374 -186 3408
rect -186 3374 -184 3408
rect -290 3339 -184 3374
rect -290 3305 -288 3339
rect -288 3305 -254 3339
rect -254 3305 -220 3339
rect -220 3305 -186 3339
rect -186 3305 -184 3339
rect -290 3279 -184 3305
rect -290 3236 -288 3240
rect -288 3236 -256 3240
rect -218 3236 -186 3240
rect -186 3236 -184 3240
rect -290 3206 -256 3236
rect -218 3206 -184 3236
rect -290 3133 -256 3167
rect -218 3133 -184 3167
rect -290 3063 -256 3094
rect -218 3063 -184 3094
rect -290 3060 -288 3063
rect -288 3060 -256 3063
rect -218 3060 -186 3063
rect -186 3060 -184 3063
rect -290 2994 -256 3021
rect -218 2994 -184 3021
rect -290 2987 -288 2994
rect -288 2987 -256 2994
rect -218 2987 -186 2994
rect -186 2987 -184 2994
rect -290 2925 -256 2948
rect -218 2925 -184 2948
rect -290 2914 -288 2925
rect -288 2914 -256 2925
rect -218 2914 -186 2925
rect -186 2914 -184 2925
rect -290 2856 -256 2875
rect -218 2856 -184 2875
rect -290 2841 -288 2856
rect -288 2841 -256 2856
rect -218 2841 -186 2856
rect -186 2841 -184 2856
rect -290 2787 -256 2802
rect -218 2787 -184 2802
rect -290 2768 -288 2787
rect -288 2768 -256 2787
rect -218 2768 -186 2787
rect -186 2768 -184 2787
rect -290 2718 -256 2729
rect -218 2718 -184 2729
rect -290 2695 -288 2718
rect -288 2695 -256 2718
rect -218 2695 -186 2718
rect -186 2695 -184 2718
rect -290 2649 -256 2656
rect -218 2649 -184 2656
rect -290 2622 -288 2649
rect -288 2622 -256 2649
rect -218 2622 -186 2649
rect -186 2622 -184 2649
rect -290 2580 -256 2583
rect -218 2580 -184 2583
rect -290 2549 -288 2580
rect -288 2549 -256 2580
rect -218 2549 -186 2580
rect -186 2549 -184 2580
rect -290 2477 -288 2510
rect -288 2477 -256 2510
rect -218 2477 -186 2510
rect -186 2477 -184 2510
rect -290 2476 -256 2477
rect -218 2476 -184 2477
rect -290 2408 -288 2437
rect -288 2408 -256 2437
rect -218 2408 -186 2437
rect -186 2408 -184 2437
rect -290 2403 -256 2408
rect -218 2403 -184 2408
rect -290 2339 -288 2364
rect -288 2339 -256 2364
rect -218 2339 -186 2364
rect -186 2339 -184 2364
rect -290 2330 -256 2339
rect -218 2330 -184 2339
rect -290 2270 -288 2291
rect -288 2270 -256 2291
rect -218 2270 -186 2291
rect -186 2270 -184 2291
rect -290 2257 -256 2270
rect -218 2257 -184 2270
rect -290 2201 -288 2218
rect -288 2201 -256 2218
rect -218 2201 -186 2218
rect -186 2201 -184 2218
rect -290 2184 -256 2201
rect -218 2184 -184 2201
rect -290 2132 -288 2145
rect -288 2132 -256 2145
rect -218 2132 -186 2145
rect -186 2132 -184 2145
rect -290 2111 -256 2132
rect -218 2111 -184 2132
rect -290 2063 -288 2072
rect -288 2063 -256 2072
rect -218 2063 -186 2072
rect -186 2063 -184 2072
rect -290 2038 -256 2063
rect -218 2038 -184 2063
rect -290 1994 -288 1999
rect -288 1994 -256 1999
rect -218 1994 -186 1999
rect -186 1994 -184 1999
rect -290 1965 -256 1994
rect -218 1965 -184 1994
rect -290 1925 -288 1926
rect -288 1925 -256 1926
rect -218 1925 -186 1926
rect -186 1925 -184 1926
rect -290 1892 -256 1925
rect -218 1892 -184 1925
rect -290 1821 -256 1853
rect -218 1821 -184 1853
rect -290 1819 -288 1821
rect -288 1819 -256 1821
rect -218 1819 -186 1821
rect -186 1819 -184 1821
rect -290 1752 -256 1780
rect -218 1752 -184 1780
rect -290 1746 -288 1752
rect -288 1746 -256 1752
rect -218 1746 -186 1752
rect -186 1746 -184 1752
rect -290 1683 -256 1707
rect -218 1683 -184 1707
rect -290 1673 -288 1683
rect -288 1673 -256 1683
rect -218 1673 -186 1683
rect -186 1673 -184 1683
rect -290 1614 -256 1634
rect -218 1614 -184 1634
rect -290 1600 -288 1614
rect -288 1600 -256 1614
rect -218 1600 -186 1614
rect -186 1600 -184 1614
rect -290 1545 -256 1561
rect -218 1545 -184 1561
rect -290 1527 -288 1545
rect -288 1527 -256 1545
rect -218 1527 -186 1545
rect -186 1527 -184 1545
rect -290 1476 -256 1488
rect -218 1476 -184 1488
rect -290 1454 -288 1476
rect -288 1454 -256 1476
rect -218 1454 -186 1476
rect -186 1454 -184 1476
rect -290 1407 -256 1415
rect -218 1407 -184 1415
rect -290 1381 -288 1407
rect -288 1381 -256 1407
rect -218 1381 -186 1407
rect -186 1381 -184 1407
rect -290 1338 -256 1342
rect -218 1338 -184 1342
rect -290 1308 -288 1338
rect -288 1308 -256 1338
rect -218 1308 -186 1338
rect -186 1308 -184 1338
rect -290 1235 -288 1269
rect -288 1235 -256 1269
rect -218 1235 -186 1269
rect -186 1235 -184 1269
rect 612 3719 614 11233
rect 614 3719 716 11233
rect 716 3719 718 11233
rect 612 3684 718 3719
rect 612 3650 614 3684
rect 614 3650 648 3684
rect 648 3650 682 3684
rect 682 3650 716 3684
rect 716 3650 718 3684
rect 612 3615 718 3650
rect 612 3581 614 3615
rect 614 3581 648 3615
rect 648 3581 682 3615
rect 682 3581 716 3615
rect 716 3581 718 3615
rect 612 3546 718 3581
rect 612 3512 614 3546
rect 614 3512 648 3546
rect 648 3512 682 3546
rect 682 3512 716 3546
rect 716 3512 718 3546
rect 612 3477 718 3512
rect 612 3443 614 3477
rect 614 3443 648 3477
rect 648 3443 682 3477
rect 682 3443 716 3477
rect 716 3443 718 3477
rect 612 3408 718 3443
rect 612 3374 614 3408
rect 614 3374 648 3408
rect 648 3374 682 3408
rect 682 3374 716 3408
rect 716 3374 718 3408
rect 612 3339 718 3374
rect 612 3305 614 3339
rect 614 3305 648 3339
rect 648 3305 682 3339
rect 682 3305 716 3339
rect 716 3305 718 3339
rect 612 3279 718 3305
rect 612 3236 614 3240
rect 614 3236 646 3240
rect 684 3236 716 3240
rect 716 3236 718 3240
rect 612 3206 646 3236
rect 684 3206 718 3236
rect 612 3133 646 3167
rect 684 3133 718 3167
rect 612 3063 646 3094
rect 684 3063 718 3094
rect 612 3060 614 3063
rect 614 3060 646 3063
rect 684 3060 716 3063
rect 716 3060 718 3063
rect 612 2994 646 3021
rect 684 2994 718 3021
rect 612 2987 614 2994
rect 614 2987 646 2994
rect 684 2987 716 2994
rect 716 2987 718 2994
rect 612 2925 646 2948
rect 684 2925 718 2948
rect 612 2914 614 2925
rect 614 2914 646 2925
rect 684 2914 716 2925
rect 716 2914 718 2925
rect 612 2856 646 2875
rect 684 2856 718 2875
rect 612 2841 614 2856
rect 614 2841 646 2856
rect 684 2841 716 2856
rect 716 2841 718 2856
rect 612 2787 646 2802
rect 684 2787 718 2802
rect 612 2768 614 2787
rect 614 2768 646 2787
rect 684 2768 716 2787
rect 716 2768 718 2787
rect 612 2718 646 2729
rect 684 2718 718 2729
rect 612 2695 614 2718
rect 614 2695 646 2718
rect 684 2695 716 2718
rect 716 2695 718 2718
rect 612 2649 646 2656
rect 684 2649 718 2656
rect 612 2622 614 2649
rect 614 2622 646 2649
rect 684 2622 716 2649
rect 716 2622 718 2649
rect 612 2580 646 2583
rect 684 2580 718 2583
rect 612 2549 614 2580
rect 614 2549 646 2580
rect 684 2549 716 2580
rect 716 2549 718 2580
rect 612 2477 614 2510
rect 614 2477 646 2510
rect 684 2477 716 2510
rect 716 2477 718 2510
rect 612 2476 646 2477
rect 684 2476 718 2477
rect 612 2408 614 2437
rect 614 2408 646 2437
rect 684 2408 716 2437
rect 716 2408 718 2437
rect 612 2403 646 2408
rect 684 2403 718 2408
rect 612 2339 614 2364
rect 614 2339 646 2364
rect 684 2339 716 2364
rect 716 2339 718 2364
rect 612 2330 646 2339
rect 684 2330 718 2339
rect 612 2270 614 2291
rect 614 2270 646 2291
rect 684 2270 716 2291
rect 716 2270 718 2291
rect 612 2257 646 2270
rect 684 2257 718 2270
rect 612 2201 614 2218
rect 614 2201 646 2218
rect 684 2201 716 2218
rect 716 2201 718 2218
rect 612 2184 646 2201
rect 684 2184 718 2201
rect 612 2132 614 2145
rect 614 2132 646 2145
rect 684 2132 716 2145
rect 716 2132 718 2145
rect 612 2111 646 2132
rect 684 2111 718 2132
rect 612 2063 614 2072
rect 614 2063 646 2072
rect 684 2063 716 2072
rect 716 2063 718 2072
rect 612 2038 646 2063
rect 684 2038 718 2063
rect 612 1994 614 1999
rect 614 1994 646 1999
rect 684 1994 716 1999
rect 716 1994 718 1999
rect 612 1965 646 1994
rect 684 1965 718 1994
rect 612 1925 614 1926
rect 614 1925 646 1926
rect 684 1925 716 1926
rect 716 1925 718 1926
rect 612 1892 646 1925
rect 684 1892 718 1925
rect 612 1821 646 1853
rect 684 1821 718 1853
rect 612 1819 614 1821
rect 614 1819 646 1821
rect 684 1819 716 1821
rect 716 1819 718 1821
rect 612 1752 646 1780
rect 684 1752 718 1780
rect 612 1746 614 1752
rect 614 1746 646 1752
rect 684 1746 716 1752
rect 716 1746 718 1752
rect 612 1683 646 1707
rect 684 1683 718 1707
rect 612 1673 614 1683
rect 614 1673 646 1683
rect 684 1673 716 1683
rect 716 1673 718 1683
rect 612 1614 646 1634
rect 684 1614 718 1634
rect 612 1600 614 1614
rect 614 1600 646 1614
rect 684 1600 716 1614
rect 716 1600 718 1614
rect 612 1545 646 1561
rect 684 1545 718 1561
rect 612 1527 614 1545
rect 614 1527 646 1545
rect 684 1527 716 1545
rect 716 1527 718 1545
rect 612 1476 646 1488
rect 684 1476 718 1488
rect 612 1454 614 1476
rect 614 1454 646 1476
rect 684 1454 716 1476
rect 716 1454 718 1476
rect 612 1407 646 1415
rect 684 1407 718 1415
rect 612 1381 614 1407
rect 614 1381 646 1407
rect 684 1381 716 1407
rect 716 1381 718 1407
rect 612 1338 646 1342
rect 684 1338 718 1342
rect 612 1308 614 1338
rect 614 1308 646 1338
rect 684 1308 716 1338
rect 716 1308 718 1338
rect 612 1235 614 1269
rect 614 1235 646 1269
rect 684 1235 716 1269
rect 716 1235 718 1269
rect 1514 3719 1516 11233
rect 1516 3719 1618 11233
rect 1618 3719 1620 11233
rect 1514 3684 1620 3719
rect 1514 3650 1516 3684
rect 1516 3650 1550 3684
rect 1550 3650 1584 3684
rect 1584 3650 1618 3684
rect 1618 3650 1620 3684
rect 1514 3615 1620 3650
rect 1514 3581 1516 3615
rect 1516 3581 1550 3615
rect 1550 3581 1584 3615
rect 1584 3581 1618 3615
rect 1618 3581 1620 3615
rect 1514 3546 1620 3581
rect 1514 3512 1516 3546
rect 1516 3512 1550 3546
rect 1550 3512 1584 3546
rect 1584 3512 1618 3546
rect 1618 3512 1620 3546
rect 1514 3477 1620 3512
rect 1514 3443 1516 3477
rect 1516 3443 1550 3477
rect 1550 3443 1584 3477
rect 1584 3443 1618 3477
rect 1618 3443 1620 3477
rect 1514 3408 1620 3443
rect 1514 3374 1516 3408
rect 1516 3374 1550 3408
rect 1550 3374 1584 3408
rect 1584 3374 1618 3408
rect 1618 3374 1620 3408
rect 1514 3339 1620 3374
rect 1514 3305 1516 3339
rect 1516 3305 1550 3339
rect 1550 3305 1584 3339
rect 1584 3305 1618 3339
rect 1618 3305 1620 3339
rect 1514 3279 1620 3305
rect 1514 3236 1516 3240
rect 1516 3236 1548 3240
rect 1586 3236 1618 3240
rect 1618 3236 1620 3240
rect 1514 3206 1548 3236
rect 1586 3206 1620 3236
rect 1514 3133 1548 3167
rect 1586 3133 1620 3167
rect 1514 3063 1548 3094
rect 1586 3063 1620 3094
rect 1514 3060 1516 3063
rect 1516 3060 1548 3063
rect 1586 3060 1618 3063
rect 1618 3060 1620 3063
rect 1514 2994 1548 3021
rect 1586 2994 1620 3021
rect 1514 2987 1516 2994
rect 1516 2987 1548 2994
rect 1586 2987 1618 2994
rect 1618 2987 1620 2994
rect 1514 2925 1548 2948
rect 1586 2925 1620 2948
rect 1514 2914 1516 2925
rect 1516 2914 1548 2925
rect 1586 2914 1618 2925
rect 1618 2914 1620 2925
rect 1514 2856 1548 2875
rect 1586 2856 1620 2875
rect 1514 2841 1516 2856
rect 1516 2841 1548 2856
rect 1586 2841 1618 2856
rect 1618 2841 1620 2856
rect 1514 2787 1548 2802
rect 1586 2787 1620 2802
rect 1514 2768 1516 2787
rect 1516 2768 1548 2787
rect 1586 2768 1618 2787
rect 1618 2768 1620 2787
rect 1514 2718 1548 2729
rect 1586 2718 1620 2729
rect 1514 2695 1516 2718
rect 1516 2695 1548 2718
rect 1586 2695 1618 2718
rect 1618 2695 1620 2718
rect 1514 2649 1548 2656
rect 1586 2649 1620 2656
rect 1514 2622 1516 2649
rect 1516 2622 1548 2649
rect 1586 2622 1618 2649
rect 1618 2622 1620 2649
rect 1514 2580 1548 2583
rect 1586 2580 1620 2583
rect 1514 2549 1516 2580
rect 1516 2549 1548 2580
rect 1586 2549 1618 2580
rect 1618 2549 1620 2580
rect 1514 2477 1516 2510
rect 1516 2477 1548 2510
rect 1586 2477 1618 2510
rect 1618 2477 1620 2510
rect 1514 2476 1548 2477
rect 1586 2476 1620 2477
rect 1514 2408 1516 2437
rect 1516 2408 1548 2437
rect 1586 2408 1618 2437
rect 1618 2408 1620 2437
rect 1514 2403 1548 2408
rect 1586 2403 1620 2408
rect 1514 2339 1516 2364
rect 1516 2339 1548 2364
rect 1586 2339 1618 2364
rect 1618 2339 1620 2364
rect 1514 2330 1548 2339
rect 1586 2330 1620 2339
rect 1514 2270 1516 2291
rect 1516 2270 1548 2291
rect 1586 2270 1618 2291
rect 1618 2270 1620 2291
rect 1514 2257 1548 2270
rect 1586 2257 1620 2270
rect 1514 2201 1516 2218
rect 1516 2201 1548 2218
rect 1586 2201 1618 2218
rect 1618 2201 1620 2218
rect 1514 2184 1548 2201
rect 1586 2184 1620 2201
rect 1514 2132 1516 2145
rect 1516 2132 1548 2145
rect 1586 2132 1618 2145
rect 1618 2132 1620 2145
rect 1514 2111 1548 2132
rect 1586 2111 1620 2132
rect 1514 2063 1516 2072
rect 1516 2063 1548 2072
rect 1586 2063 1618 2072
rect 1618 2063 1620 2072
rect 1514 2038 1548 2063
rect 1586 2038 1620 2063
rect 1514 1994 1516 1999
rect 1516 1994 1548 1999
rect 1586 1994 1618 1999
rect 1618 1994 1620 1999
rect 1514 1965 1548 1994
rect 1586 1965 1620 1994
rect 1514 1925 1516 1926
rect 1516 1925 1548 1926
rect 1586 1925 1618 1926
rect 1618 1925 1620 1926
rect 1514 1892 1548 1925
rect 1586 1892 1620 1925
rect 1514 1821 1548 1853
rect 1586 1821 1620 1853
rect 1514 1819 1516 1821
rect 1516 1819 1548 1821
rect 1586 1819 1618 1821
rect 1618 1819 1620 1821
rect 1514 1752 1548 1780
rect 1586 1752 1620 1780
rect 1514 1746 1516 1752
rect 1516 1746 1548 1752
rect 1586 1746 1618 1752
rect 1618 1746 1620 1752
rect 1514 1683 1548 1707
rect 1586 1683 1620 1707
rect 1514 1673 1516 1683
rect 1516 1673 1548 1683
rect 1586 1673 1618 1683
rect 1618 1673 1620 1683
rect 1514 1614 1548 1634
rect 1586 1614 1620 1634
rect 1514 1600 1516 1614
rect 1516 1600 1548 1614
rect 1586 1600 1618 1614
rect 1618 1600 1620 1614
rect 1514 1545 1548 1561
rect 1586 1545 1620 1561
rect 1514 1527 1516 1545
rect 1516 1527 1548 1545
rect 1586 1527 1618 1545
rect 1618 1527 1620 1545
rect 1514 1476 1548 1488
rect 1586 1476 1620 1488
rect 1514 1454 1516 1476
rect 1516 1454 1548 1476
rect 1586 1454 1618 1476
rect 1618 1454 1620 1476
rect 1514 1407 1548 1415
rect 1586 1407 1620 1415
rect 1514 1381 1516 1407
rect 1516 1381 1548 1407
rect 1586 1381 1618 1407
rect 1618 1381 1620 1407
rect 1514 1338 1548 1342
rect 1586 1338 1620 1342
rect 1514 1308 1516 1338
rect 1516 1308 1548 1338
rect 1586 1308 1618 1338
rect 1618 1308 1620 1338
rect 1514 1235 1516 1269
rect 1516 1235 1548 1269
rect 1586 1235 1618 1269
rect 1618 1235 1620 1269
rect 2416 3719 2418 11233
rect 2418 3719 2520 11233
rect 2520 3719 2522 11233
rect 2416 3684 2522 3719
rect 2416 3650 2418 3684
rect 2418 3650 2452 3684
rect 2452 3650 2486 3684
rect 2486 3650 2520 3684
rect 2520 3650 2522 3684
rect 2416 3615 2522 3650
rect 2416 3581 2418 3615
rect 2418 3581 2452 3615
rect 2452 3581 2486 3615
rect 2486 3581 2520 3615
rect 2520 3581 2522 3615
rect 2416 3546 2522 3581
rect 2416 3512 2418 3546
rect 2418 3512 2452 3546
rect 2452 3512 2486 3546
rect 2486 3512 2520 3546
rect 2520 3512 2522 3546
rect 2416 3477 2522 3512
rect 2416 3443 2418 3477
rect 2418 3443 2452 3477
rect 2452 3443 2486 3477
rect 2486 3443 2520 3477
rect 2520 3443 2522 3477
rect 2416 3408 2522 3443
rect 2416 3374 2418 3408
rect 2418 3374 2452 3408
rect 2452 3374 2486 3408
rect 2486 3374 2520 3408
rect 2520 3374 2522 3408
rect 2416 3339 2522 3374
rect 2416 3305 2418 3339
rect 2418 3305 2452 3339
rect 2452 3305 2486 3339
rect 2486 3305 2520 3339
rect 2520 3305 2522 3339
rect 2416 3279 2522 3305
rect 2416 3236 2418 3240
rect 2418 3236 2450 3240
rect 2488 3236 2520 3240
rect 2520 3236 2522 3240
rect 2416 3206 2450 3236
rect 2488 3206 2522 3236
rect 2416 3133 2450 3167
rect 2488 3133 2522 3167
rect 2416 3063 2450 3094
rect 2488 3063 2522 3094
rect 2416 3060 2418 3063
rect 2418 3060 2450 3063
rect 2488 3060 2520 3063
rect 2520 3060 2522 3063
rect 2416 2994 2450 3021
rect 2488 2994 2522 3021
rect 2416 2987 2418 2994
rect 2418 2987 2450 2994
rect 2488 2987 2520 2994
rect 2520 2987 2522 2994
rect 2416 2925 2450 2948
rect 2488 2925 2522 2948
rect 2416 2914 2418 2925
rect 2418 2914 2450 2925
rect 2488 2914 2520 2925
rect 2520 2914 2522 2925
rect 2416 2856 2450 2875
rect 2488 2856 2522 2875
rect 2416 2841 2418 2856
rect 2418 2841 2450 2856
rect 2488 2841 2520 2856
rect 2520 2841 2522 2856
rect 2416 2787 2450 2802
rect 2488 2787 2522 2802
rect 2416 2768 2418 2787
rect 2418 2768 2450 2787
rect 2488 2768 2520 2787
rect 2520 2768 2522 2787
rect 2416 2718 2450 2729
rect 2488 2718 2522 2729
rect 2416 2695 2418 2718
rect 2418 2695 2450 2718
rect 2488 2695 2520 2718
rect 2520 2695 2522 2718
rect 2416 2649 2450 2656
rect 2488 2649 2522 2656
rect 2416 2622 2418 2649
rect 2418 2622 2450 2649
rect 2488 2622 2520 2649
rect 2520 2622 2522 2649
rect 2416 2580 2450 2583
rect 2488 2580 2522 2583
rect 2416 2549 2418 2580
rect 2418 2549 2450 2580
rect 2488 2549 2520 2580
rect 2520 2549 2522 2580
rect 2416 2477 2418 2510
rect 2418 2477 2450 2510
rect 2488 2477 2520 2510
rect 2520 2477 2522 2510
rect 2416 2476 2450 2477
rect 2488 2476 2522 2477
rect 2416 2408 2418 2437
rect 2418 2408 2450 2437
rect 2488 2408 2520 2437
rect 2520 2408 2522 2437
rect 2416 2403 2450 2408
rect 2488 2403 2522 2408
rect 2416 2339 2418 2364
rect 2418 2339 2450 2364
rect 2488 2339 2520 2364
rect 2520 2339 2522 2364
rect 2416 2330 2450 2339
rect 2488 2330 2522 2339
rect 2416 2270 2418 2291
rect 2418 2270 2450 2291
rect 2488 2270 2520 2291
rect 2520 2270 2522 2291
rect 2416 2257 2450 2270
rect 2488 2257 2522 2270
rect 2416 2201 2418 2218
rect 2418 2201 2450 2218
rect 2488 2201 2520 2218
rect 2520 2201 2522 2218
rect 2416 2184 2450 2201
rect 2488 2184 2522 2201
rect 2416 2132 2418 2145
rect 2418 2132 2450 2145
rect 2488 2132 2520 2145
rect 2520 2132 2522 2145
rect 2416 2111 2450 2132
rect 2488 2111 2522 2132
rect 2416 2063 2418 2072
rect 2418 2063 2450 2072
rect 2488 2063 2520 2072
rect 2520 2063 2522 2072
rect 2416 2038 2450 2063
rect 2488 2038 2522 2063
rect 2416 1994 2418 1999
rect 2418 1994 2450 1999
rect 2488 1994 2520 1999
rect 2520 1994 2522 1999
rect 2416 1965 2450 1994
rect 2488 1965 2522 1994
rect 2416 1925 2418 1926
rect 2418 1925 2450 1926
rect 2488 1925 2520 1926
rect 2520 1925 2522 1926
rect 2416 1892 2450 1925
rect 2488 1892 2522 1925
rect 2416 1821 2450 1853
rect 2488 1821 2522 1853
rect 2416 1819 2418 1821
rect 2418 1819 2450 1821
rect 2488 1819 2520 1821
rect 2520 1819 2522 1821
rect 2416 1752 2450 1780
rect 2488 1752 2522 1780
rect 2416 1746 2418 1752
rect 2418 1746 2450 1752
rect 2488 1746 2520 1752
rect 2520 1746 2522 1752
rect 2416 1683 2450 1707
rect 2488 1683 2522 1707
rect 2416 1673 2418 1683
rect 2418 1673 2450 1683
rect 2488 1673 2520 1683
rect 2520 1673 2522 1683
rect 2416 1614 2450 1634
rect 2488 1614 2522 1634
rect 2416 1600 2418 1614
rect 2418 1600 2450 1614
rect 2488 1600 2520 1614
rect 2520 1600 2522 1614
rect 2416 1545 2450 1561
rect 2488 1545 2522 1561
rect 2416 1527 2418 1545
rect 2418 1527 2450 1545
rect 2488 1527 2520 1545
rect 2520 1527 2522 1545
rect 2416 1476 2450 1488
rect 2488 1476 2522 1488
rect 2416 1454 2418 1476
rect 2418 1454 2450 1476
rect 2488 1454 2520 1476
rect 2520 1454 2522 1476
rect 2416 1407 2450 1415
rect 2488 1407 2522 1415
rect 2416 1381 2418 1407
rect 2418 1381 2450 1407
rect 2488 1381 2520 1407
rect 2520 1381 2522 1407
rect 2416 1338 2450 1342
rect 2488 1338 2522 1342
rect 2416 1308 2418 1338
rect 2418 1308 2450 1338
rect 2488 1308 2520 1338
rect 2520 1308 2522 1338
rect 2416 1235 2418 1269
rect 2418 1235 2450 1269
rect 2488 1235 2520 1269
rect 2520 1235 2522 1269
rect 3318 3719 3320 11233
rect 3320 3719 3422 11233
rect 3422 3719 3424 11233
rect 3318 3684 3424 3719
rect 3318 3650 3320 3684
rect 3320 3650 3354 3684
rect 3354 3650 3388 3684
rect 3388 3650 3422 3684
rect 3422 3650 3424 3684
rect 3318 3615 3424 3650
rect 3318 3581 3320 3615
rect 3320 3581 3354 3615
rect 3354 3581 3388 3615
rect 3388 3581 3422 3615
rect 3422 3581 3424 3615
rect 3318 3546 3424 3581
rect 3318 3512 3320 3546
rect 3320 3512 3354 3546
rect 3354 3512 3388 3546
rect 3388 3512 3422 3546
rect 3422 3512 3424 3546
rect 3318 3477 3424 3512
rect 3318 3443 3320 3477
rect 3320 3443 3354 3477
rect 3354 3443 3388 3477
rect 3388 3443 3422 3477
rect 3422 3443 3424 3477
rect 3318 3408 3424 3443
rect 3318 3374 3320 3408
rect 3320 3374 3354 3408
rect 3354 3374 3388 3408
rect 3388 3374 3422 3408
rect 3422 3374 3424 3408
rect 3318 3339 3424 3374
rect 3318 3305 3320 3339
rect 3320 3305 3354 3339
rect 3354 3305 3388 3339
rect 3388 3305 3422 3339
rect 3422 3305 3424 3339
rect 3318 3279 3424 3305
rect 3318 3236 3320 3240
rect 3320 3236 3352 3240
rect 3390 3236 3422 3240
rect 3422 3236 3424 3240
rect 3318 3206 3352 3236
rect 3390 3206 3424 3236
rect 3318 3133 3352 3167
rect 3390 3133 3424 3167
rect 3318 3063 3352 3094
rect 3390 3063 3424 3094
rect 3318 3060 3320 3063
rect 3320 3060 3352 3063
rect 3390 3060 3422 3063
rect 3422 3060 3424 3063
rect 3318 2994 3352 3021
rect 3390 2994 3424 3021
rect 3318 2987 3320 2994
rect 3320 2987 3352 2994
rect 3390 2987 3422 2994
rect 3422 2987 3424 2994
rect 3318 2925 3352 2948
rect 3390 2925 3424 2948
rect 3318 2914 3320 2925
rect 3320 2914 3352 2925
rect 3390 2914 3422 2925
rect 3422 2914 3424 2925
rect 3318 2856 3352 2875
rect 3390 2856 3424 2875
rect 3318 2841 3320 2856
rect 3320 2841 3352 2856
rect 3390 2841 3422 2856
rect 3422 2841 3424 2856
rect 3318 2787 3352 2802
rect 3390 2787 3424 2802
rect 3318 2768 3320 2787
rect 3320 2768 3352 2787
rect 3390 2768 3422 2787
rect 3422 2768 3424 2787
rect 3318 2718 3352 2729
rect 3390 2718 3424 2729
rect 3318 2695 3320 2718
rect 3320 2695 3352 2718
rect 3390 2695 3422 2718
rect 3422 2695 3424 2718
rect 3318 2649 3352 2656
rect 3390 2649 3424 2656
rect 3318 2622 3320 2649
rect 3320 2622 3352 2649
rect 3390 2622 3422 2649
rect 3422 2622 3424 2649
rect 3318 2580 3352 2583
rect 3390 2580 3424 2583
rect 3318 2549 3320 2580
rect 3320 2549 3352 2580
rect 3390 2549 3422 2580
rect 3422 2549 3424 2580
rect 3318 2477 3320 2510
rect 3320 2477 3352 2510
rect 3390 2477 3422 2510
rect 3422 2477 3424 2510
rect 3318 2476 3352 2477
rect 3390 2476 3424 2477
rect 3318 2408 3320 2437
rect 3320 2408 3352 2437
rect 3390 2408 3422 2437
rect 3422 2408 3424 2437
rect 3318 2403 3352 2408
rect 3390 2403 3424 2408
rect 3318 2339 3320 2364
rect 3320 2339 3352 2364
rect 3390 2339 3422 2364
rect 3422 2339 3424 2364
rect 3318 2330 3352 2339
rect 3390 2330 3424 2339
rect 3318 2270 3320 2291
rect 3320 2270 3352 2291
rect 3390 2270 3422 2291
rect 3422 2270 3424 2291
rect 3318 2257 3352 2270
rect 3390 2257 3424 2270
rect 3318 2201 3320 2218
rect 3320 2201 3352 2218
rect 3390 2201 3422 2218
rect 3422 2201 3424 2218
rect 3318 2184 3352 2201
rect 3390 2184 3424 2201
rect 3318 2132 3320 2145
rect 3320 2132 3352 2145
rect 3390 2132 3422 2145
rect 3422 2132 3424 2145
rect 3318 2111 3352 2132
rect 3390 2111 3424 2132
rect 3318 2063 3320 2072
rect 3320 2063 3352 2072
rect 3390 2063 3422 2072
rect 3422 2063 3424 2072
rect 3318 2038 3352 2063
rect 3390 2038 3424 2063
rect 3318 1994 3320 1999
rect 3320 1994 3352 1999
rect 3390 1994 3422 1999
rect 3422 1994 3424 1999
rect 3318 1965 3352 1994
rect 3390 1965 3424 1994
rect 3318 1925 3320 1926
rect 3320 1925 3352 1926
rect 3390 1925 3422 1926
rect 3422 1925 3424 1926
rect 3318 1892 3352 1925
rect 3390 1892 3424 1925
rect 3318 1821 3352 1853
rect 3390 1821 3424 1853
rect 3318 1819 3320 1821
rect 3320 1819 3352 1821
rect 3390 1819 3422 1821
rect 3422 1819 3424 1821
rect 3318 1752 3352 1780
rect 3390 1752 3424 1780
rect 3318 1746 3320 1752
rect 3320 1746 3352 1752
rect 3390 1746 3422 1752
rect 3422 1746 3424 1752
rect 3318 1683 3352 1707
rect 3390 1683 3424 1707
rect 3318 1673 3320 1683
rect 3320 1673 3352 1683
rect 3390 1673 3422 1683
rect 3422 1673 3424 1683
rect 3318 1614 3352 1634
rect 3390 1614 3424 1634
rect 3318 1600 3320 1614
rect 3320 1600 3352 1614
rect 3390 1600 3422 1614
rect 3422 1600 3424 1614
rect 3318 1545 3352 1561
rect 3390 1545 3424 1561
rect 3318 1527 3320 1545
rect 3320 1527 3352 1545
rect 3390 1527 3422 1545
rect 3422 1527 3424 1545
rect 3318 1476 3352 1488
rect 3390 1476 3424 1488
rect 3318 1454 3320 1476
rect 3320 1454 3352 1476
rect 3390 1454 3422 1476
rect 3422 1454 3424 1476
rect 3318 1407 3352 1415
rect 3390 1407 3424 1415
rect 3318 1381 3320 1407
rect 3320 1381 3352 1407
rect 3390 1381 3422 1407
rect 3422 1381 3424 1407
rect 3318 1338 3352 1342
rect 3390 1338 3424 1342
rect 3318 1308 3320 1338
rect 3320 1308 3352 1338
rect 3390 1308 3422 1338
rect 3422 1308 3424 1338
rect 3318 1235 3320 1269
rect 3320 1235 3352 1269
rect 3390 1235 3422 1269
rect 3422 1235 3424 1269
rect 4220 3719 4222 11233
rect 4222 3719 4324 11233
rect 4324 3719 4326 11233
rect 4220 3684 4326 3719
rect 4220 3650 4222 3684
rect 4222 3650 4256 3684
rect 4256 3650 4290 3684
rect 4290 3650 4324 3684
rect 4324 3650 4326 3684
rect 4220 3615 4326 3650
rect 4220 3581 4222 3615
rect 4222 3581 4256 3615
rect 4256 3581 4290 3615
rect 4290 3581 4324 3615
rect 4324 3581 4326 3615
rect 4220 3546 4326 3581
rect 4220 3512 4222 3546
rect 4222 3512 4256 3546
rect 4256 3512 4290 3546
rect 4290 3512 4324 3546
rect 4324 3512 4326 3546
rect 4220 3477 4326 3512
rect 4220 3443 4222 3477
rect 4222 3443 4256 3477
rect 4256 3443 4290 3477
rect 4290 3443 4324 3477
rect 4324 3443 4326 3477
rect 4220 3408 4326 3443
rect 4220 3374 4222 3408
rect 4222 3374 4256 3408
rect 4256 3374 4290 3408
rect 4290 3374 4324 3408
rect 4324 3374 4326 3408
rect 4220 3339 4326 3374
rect 4220 3305 4222 3339
rect 4222 3305 4256 3339
rect 4256 3305 4290 3339
rect 4290 3305 4324 3339
rect 4324 3305 4326 3339
rect 4220 3279 4326 3305
rect 4220 3236 4222 3240
rect 4222 3236 4254 3240
rect 4292 3236 4324 3240
rect 4324 3236 4326 3240
rect 4220 3206 4254 3236
rect 4292 3206 4326 3236
rect 4220 3133 4254 3167
rect 4292 3133 4326 3167
rect 4220 3063 4254 3094
rect 4292 3063 4326 3094
rect 4220 3060 4222 3063
rect 4222 3060 4254 3063
rect 4292 3060 4324 3063
rect 4324 3060 4326 3063
rect 4220 2994 4254 3021
rect 4292 2994 4326 3021
rect 4220 2987 4222 2994
rect 4222 2987 4254 2994
rect 4292 2987 4324 2994
rect 4324 2987 4326 2994
rect 4220 2925 4254 2948
rect 4292 2925 4326 2948
rect 4220 2914 4222 2925
rect 4222 2914 4254 2925
rect 4292 2914 4324 2925
rect 4324 2914 4326 2925
rect 4220 2856 4254 2875
rect 4292 2856 4326 2875
rect 4220 2841 4222 2856
rect 4222 2841 4254 2856
rect 4292 2841 4324 2856
rect 4324 2841 4326 2856
rect 4220 2787 4254 2802
rect 4292 2787 4326 2802
rect 4220 2768 4222 2787
rect 4222 2768 4254 2787
rect 4292 2768 4324 2787
rect 4324 2768 4326 2787
rect 4220 2718 4254 2729
rect 4292 2718 4326 2729
rect 4220 2695 4222 2718
rect 4222 2695 4254 2718
rect 4292 2695 4324 2718
rect 4324 2695 4326 2718
rect 4220 2649 4254 2656
rect 4292 2649 4326 2656
rect 4220 2622 4222 2649
rect 4222 2622 4254 2649
rect 4292 2622 4324 2649
rect 4324 2622 4326 2649
rect 4220 2580 4254 2583
rect 4292 2580 4326 2583
rect 4220 2549 4222 2580
rect 4222 2549 4254 2580
rect 4292 2549 4324 2580
rect 4324 2549 4326 2580
rect 4220 2477 4222 2510
rect 4222 2477 4254 2510
rect 4292 2477 4324 2510
rect 4324 2477 4326 2510
rect 4220 2476 4254 2477
rect 4292 2476 4326 2477
rect 4220 2408 4222 2437
rect 4222 2408 4254 2437
rect 4292 2408 4324 2437
rect 4324 2408 4326 2437
rect 4220 2403 4254 2408
rect 4292 2403 4326 2408
rect 4220 2339 4222 2364
rect 4222 2339 4254 2364
rect 4292 2339 4324 2364
rect 4324 2339 4326 2364
rect 4220 2330 4254 2339
rect 4292 2330 4326 2339
rect 4220 2270 4222 2291
rect 4222 2270 4254 2291
rect 4292 2270 4324 2291
rect 4324 2270 4326 2291
rect 4220 2257 4254 2270
rect 4292 2257 4326 2270
rect 4220 2201 4222 2218
rect 4222 2201 4254 2218
rect 4292 2201 4324 2218
rect 4324 2201 4326 2218
rect 4220 2184 4254 2201
rect 4292 2184 4326 2201
rect 4220 2132 4222 2145
rect 4222 2132 4254 2145
rect 4292 2132 4324 2145
rect 4324 2132 4326 2145
rect 4220 2111 4254 2132
rect 4292 2111 4326 2132
rect 4220 2063 4222 2072
rect 4222 2063 4254 2072
rect 4292 2063 4324 2072
rect 4324 2063 4326 2072
rect 4220 2038 4254 2063
rect 4292 2038 4326 2063
rect 4220 1994 4222 1999
rect 4222 1994 4254 1999
rect 4292 1994 4324 1999
rect 4324 1994 4326 1999
rect 4220 1965 4254 1994
rect 4292 1965 4326 1994
rect 4220 1925 4222 1926
rect 4222 1925 4254 1926
rect 4292 1925 4324 1926
rect 4324 1925 4326 1926
rect 4220 1892 4254 1925
rect 4292 1892 4326 1925
rect 4220 1821 4254 1853
rect 4292 1821 4326 1853
rect 4220 1819 4222 1821
rect 4222 1819 4254 1821
rect 4292 1819 4324 1821
rect 4324 1819 4326 1821
rect 4220 1752 4254 1780
rect 4292 1752 4326 1780
rect 4220 1746 4222 1752
rect 4222 1746 4254 1752
rect 4292 1746 4324 1752
rect 4324 1746 4326 1752
rect 4220 1683 4254 1707
rect 4292 1683 4326 1707
rect 4220 1673 4222 1683
rect 4222 1673 4254 1683
rect 4292 1673 4324 1683
rect 4324 1673 4326 1683
rect 4220 1614 4254 1634
rect 4292 1614 4326 1634
rect 4220 1600 4222 1614
rect 4222 1600 4254 1614
rect 4292 1600 4324 1614
rect 4324 1600 4326 1614
rect 4220 1545 4254 1561
rect 4292 1545 4326 1561
rect 4220 1527 4222 1545
rect 4222 1527 4254 1545
rect 4292 1527 4324 1545
rect 4324 1527 4326 1545
rect 4220 1476 4254 1488
rect 4292 1476 4326 1488
rect 4220 1454 4222 1476
rect 4222 1454 4254 1476
rect 4292 1454 4324 1476
rect 4324 1454 4326 1476
rect 4220 1407 4254 1415
rect 4292 1407 4326 1415
rect 4220 1381 4222 1407
rect 4222 1381 4254 1407
rect 4292 1381 4324 1407
rect 4324 1381 4326 1407
rect 4220 1338 4254 1342
rect 4292 1338 4326 1342
rect 4220 1308 4222 1338
rect 4222 1308 4254 1338
rect 4292 1308 4324 1338
rect 4324 1308 4326 1338
rect 4220 1235 4222 1269
rect 4222 1235 4254 1269
rect 4292 1235 4324 1269
rect 4324 1235 4326 1269
rect 5122 3719 5124 11233
rect 5124 3719 5226 11233
rect 5226 3719 5228 11233
rect 5122 3684 5228 3719
rect 5122 3650 5124 3684
rect 5124 3650 5158 3684
rect 5158 3650 5192 3684
rect 5192 3650 5226 3684
rect 5226 3650 5228 3684
rect 5122 3615 5228 3650
rect 5122 3581 5124 3615
rect 5124 3581 5158 3615
rect 5158 3581 5192 3615
rect 5192 3581 5226 3615
rect 5226 3581 5228 3615
rect 5122 3546 5228 3581
rect 5122 3512 5124 3546
rect 5124 3512 5158 3546
rect 5158 3512 5192 3546
rect 5192 3512 5226 3546
rect 5226 3512 5228 3546
rect 5122 3477 5228 3512
rect 5122 3443 5124 3477
rect 5124 3443 5158 3477
rect 5158 3443 5192 3477
rect 5192 3443 5226 3477
rect 5226 3443 5228 3477
rect 5122 3408 5228 3443
rect 5122 3374 5124 3408
rect 5124 3374 5158 3408
rect 5158 3374 5192 3408
rect 5192 3374 5226 3408
rect 5226 3374 5228 3408
rect 5122 3339 5228 3374
rect 5122 3305 5124 3339
rect 5124 3305 5158 3339
rect 5158 3305 5192 3339
rect 5192 3305 5226 3339
rect 5226 3305 5228 3339
rect 5122 3279 5228 3305
rect 5122 3236 5124 3240
rect 5124 3236 5156 3240
rect 5194 3236 5226 3240
rect 5226 3236 5228 3240
rect 5122 3206 5156 3236
rect 5194 3206 5228 3236
rect 5122 3133 5156 3167
rect 5194 3133 5228 3167
rect 5122 3063 5156 3094
rect 5194 3063 5228 3094
rect 5122 3060 5124 3063
rect 5124 3060 5156 3063
rect 5194 3060 5226 3063
rect 5226 3060 5228 3063
rect 5122 2994 5156 3021
rect 5194 2994 5228 3021
rect 5122 2987 5124 2994
rect 5124 2987 5156 2994
rect 5194 2987 5226 2994
rect 5226 2987 5228 2994
rect 5122 2925 5156 2948
rect 5194 2925 5228 2948
rect 5122 2914 5124 2925
rect 5124 2914 5156 2925
rect 5194 2914 5226 2925
rect 5226 2914 5228 2925
rect 5122 2856 5156 2875
rect 5194 2856 5228 2875
rect 5122 2841 5124 2856
rect 5124 2841 5156 2856
rect 5194 2841 5226 2856
rect 5226 2841 5228 2856
rect 5122 2787 5156 2802
rect 5194 2787 5228 2802
rect 5122 2768 5124 2787
rect 5124 2768 5156 2787
rect 5194 2768 5226 2787
rect 5226 2768 5228 2787
rect 5122 2718 5156 2729
rect 5194 2718 5228 2729
rect 5122 2695 5124 2718
rect 5124 2695 5156 2718
rect 5194 2695 5226 2718
rect 5226 2695 5228 2718
rect 5122 2649 5156 2656
rect 5194 2649 5228 2656
rect 5122 2622 5124 2649
rect 5124 2622 5156 2649
rect 5194 2622 5226 2649
rect 5226 2622 5228 2649
rect 5122 2580 5156 2583
rect 5194 2580 5228 2583
rect 5122 2549 5124 2580
rect 5124 2549 5156 2580
rect 5194 2549 5226 2580
rect 5226 2549 5228 2580
rect 5122 2477 5124 2510
rect 5124 2477 5156 2510
rect 5194 2477 5226 2510
rect 5226 2477 5228 2510
rect 5122 2476 5156 2477
rect 5194 2476 5228 2477
rect 5122 2408 5124 2437
rect 5124 2408 5156 2437
rect 5194 2408 5226 2437
rect 5226 2408 5228 2437
rect 5122 2403 5156 2408
rect 5194 2403 5228 2408
rect 5122 2339 5124 2364
rect 5124 2339 5156 2364
rect 5194 2339 5226 2364
rect 5226 2339 5228 2364
rect 5122 2330 5156 2339
rect 5194 2330 5228 2339
rect 5122 2270 5124 2291
rect 5124 2270 5156 2291
rect 5194 2270 5226 2291
rect 5226 2270 5228 2291
rect 5122 2257 5156 2270
rect 5194 2257 5228 2270
rect 5122 2201 5124 2218
rect 5124 2201 5156 2218
rect 5194 2201 5226 2218
rect 5226 2201 5228 2218
rect 5122 2184 5156 2201
rect 5194 2184 5228 2201
rect 5122 2132 5124 2145
rect 5124 2132 5156 2145
rect 5194 2132 5226 2145
rect 5226 2132 5228 2145
rect 5122 2111 5156 2132
rect 5194 2111 5228 2132
rect 5122 2063 5124 2072
rect 5124 2063 5156 2072
rect 5194 2063 5226 2072
rect 5226 2063 5228 2072
rect 5122 2038 5156 2063
rect 5194 2038 5228 2063
rect 5122 1994 5124 1999
rect 5124 1994 5156 1999
rect 5194 1994 5226 1999
rect 5226 1994 5228 1999
rect 5122 1965 5156 1994
rect 5194 1965 5228 1994
rect 5122 1925 5124 1926
rect 5124 1925 5156 1926
rect 5194 1925 5226 1926
rect 5226 1925 5228 1926
rect 5122 1892 5156 1925
rect 5194 1892 5228 1925
rect 5122 1821 5156 1853
rect 5194 1821 5228 1853
rect 5122 1819 5124 1821
rect 5124 1819 5156 1821
rect 5194 1819 5226 1821
rect 5226 1819 5228 1821
rect 5122 1752 5156 1780
rect 5194 1752 5228 1780
rect 5122 1746 5124 1752
rect 5124 1746 5156 1752
rect 5194 1746 5226 1752
rect 5226 1746 5228 1752
rect 5122 1683 5156 1707
rect 5194 1683 5228 1707
rect 5122 1673 5124 1683
rect 5124 1673 5156 1683
rect 5194 1673 5226 1683
rect 5226 1673 5228 1683
rect 5122 1614 5156 1634
rect 5194 1614 5228 1634
rect 5122 1600 5124 1614
rect 5124 1600 5156 1614
rect 5194 1600 5226 1614
rect 5226 1600 5228 1614
rect 5122 1545 5156 1561
rect 5194 1545 5228 1561
rect 5122 1527 5124 1545
rect 5124 1527 5156 1545
rect 5194 1527 5226 1545
rect 5226 1527 5228 1545
rect 5122 1476 5156 1488
rect 5194 1476 5228 1488
rect 5122 1454 5124 1476
rect 5124 1454 5156 1476
rect 5194 1454 5226 1476
rect 5226 1454 5228 1476
rect 5122 1407 5156 1415
rect 5194 1407 5228 1415
rect 5122 1381 5124 1407
rect 5124 1381 5156 1407
rect 5194 1381 5226 1407
rect 5226 1381 5228 1407
rect 5122 1338 5156 1342
rect 5194 1338 5228 1342
rect 5122 1308 5124 1338
rect 5124 1308 5156 1338
rect 5194 1308 5226 1338
rect 5226 1308 5228 1338
rect 5122 1235 5124 1269
rect 5124 1235 5156 1269
rect 5194 1235 5226 1269
rect 5226 1235 5228 1269
rect 6024 3719 6026 11233
rect 6026 3719 6128 11233
rect 6128 3719 6130 11233
rect 6024 3684 6130 3719
rect 6024 3650 6026 3684
rect 6026 3650 6060 3684
rect 6060 3650 6094 3684
rect 6094 3650 6128 3684
rect 6128 3650 6130 3684
rect 6024 3615 6130 3650
rect 6024 3581 6026 3615
rect 6026 3581 6060 3615
rect 6060 3581 6094 3615
rect 6094 3581 6128 3615
rect 6128 3581 6130 3615
rect 6024 3546 6130 3581
rect 6024 3512 6026 3546
rect 6026 3512 6060 3546
rect 6060 3512 6094 3546
rect 6094 3512 6128 3546
rect 6128 3512 6130 3546
rect 6024 3477 6130 3512
rect 6024 3443 6026 3477
rect 6026 3443 6060 3477
rect 6060 3443 6094 3477
rect 6094 3443 6128 3477
rect 6128 3443 6130 3477
rect 6024 3408 6130 3443
rect 6024 3374 6026 3408
rect 6026 3374 6060 3408
rect 6060 3374 6094 3408
rect 6094 3374 6128 3408
rect 6128 3374 6130 3408
rect 6024 3339 6130 3374
rect 6024 3305 6026 3339
rect 6026 3305 6060 3339
rect 6060 3305 6094 3339
rect 6094 3305 6128 3339
rect 6128 3305 6130 3339
rect 6024 3279 6130 3305
rect 6024 3236 6026 3240
rect 6026 3236 6058 3240
rect 6096 3236 6128 3240
rect 6128 3236 6130 3240
rect 6024 3206 6058 3236
rect 6096 3206 6130 3236
rect 6024 3133 6058 3167
rect 6096 3133 6130 3167
rect 6024 3063 6058 3094
rect 6096 3063 6130 3094
rect 6024 3060 6026 3063
rect 6026 3060 6058 3063
rect 6096 3060 6128 3063
rect 6128 3060 6130 3063
rect 6024 2994 6058 3021
rect 6096 2994 6130 3021
rect 6024 2987 6026 2994
rect 6026 2987 6058 2994
rect 6096 2987 6128 2994
rect 6128 2987 6130 2994
rect 6024 2925 6058 2948
rect 6096 2925 6130 2948
rect 6024 2914 6026 2925
rect 6026 2914 6058 2925
rect 6096 2914 6128 2925
rect 6128 2914 6130 2925
rect 6024 2856 6058 2875
rect 6096 2856 6130 2875
rect 6024 2841 6026 2856
rect 6026 2841 6058 2856
rect 6096 2841 6128 2856
rect 6128 2841 6130 2856
rect 6024 2787 6058 2802
rect 6096 2787 6130 2802
rect 6024 2768 6026 2787
rect 6026 2768 6058 2787
rect 6096 2768 6128 2787
rect 6128 2768 6130 2787
rect 6024 2718 6058 2729
rect 6096 2718 6130 2729
rect 6024 2695 6026 2718
rect 6026 2695 6058 2718
rect 6096 2695 6128 2718
rect 6128 2695 6130 2718
rect 6024 2649 6058 2656
rect 6096 2649 6130 2656
rect 6024 2622 6026 2649
rect 6026 2622 6058 2649
rect 6096 2622 6128 2649
rect 6128 2622 6130 2649
rect 6024 2580 6058 2583
rect 6096 2580 6130 2583
rect 6024 2549 6026 2580
rect 6026 2549 6058 2580
rect 6096 2549 6128 2580
rect 6128 2549 6130 2580
rect 6024 2477 6026 2510
rect 6026 2477 6058 2510
rect 6096 2477 6128 2510
rect 6128 2477 6130 2510
rect 6024 2476 6058 2477
rect 6096 2476 6130 2477
rect 6024 2408 6026 2437
rect 6026 2408 6058 2437
rect 6096 2408 6128 2437
rect 6128 2408 6130 2437
rect 6024 2403 6058 2408
rect 6096 2403 6130 2408
rect 6024 2339 6026 2364
rect 6026 2339 6058 2364
rect 6096 2339 6128 2364
rect 6128 2339 6130 2364
rect 6024 2330 6058 2339
rect 6096 2330 6130 2339
rect 6024 2270 6026 2291
rect 6026 2270 6058 2291
rect 6096 2270 6128 2291
rect 6128 2270 6130 2291
rect 6024 2257 6058 2270
rect 6096 2257 6130 2270
rect 6024 2201 6026 2218
rect 6026 2201 6058 2218
rect 6096 2201 6128 2218
rect 6128 2201 6130 2218
rect 6024 2184 6058 2201
rect 6096 2184 6130 2201
rect 6024 2132 6026 2145
rect 6026 2132 6058 2145
rect 6096 2132 6128 2145
rect 6128 2132 6130 2145
rect 6024 2111 6058 2132
rect 6096 2111 6130 2132
rect 6024 2063 6026 2072
rect 6026 2063 6058 2072
rect 6096 2063 6128 2072
rect 6128 2063 6130 2072
rect 6024 2038 6058 2063
rect 6096 2038 6130 2063
rect 6024 1994 6026 1999
rect 6026 1994 6058 1999
rect 6096 1994 6128 1999
rect 6128 1994 6130 1999
rect 6024 1965 6058 1994
rect 6096 1965 6130 1994
rect 6024 1925 6026 1926
rect 6026 1925 6058 1926
rect 6096 1925 6128 1926
rect 6128 1925 6130 1926
rect 6024 1892 6058 1925
rect 6096 1892 6130 1925
rect 6024 1821 6058 1853
rect 6096 1821 6130 1853
rect 6024 1819 6026 1821
rect 6026 1819 6058 1821
rect 6096 1819 6128 1821
rect 6128 1819 6130 1821
rect 6024 1752 6058 1780
rect 6096 1752 6130 1780
rect 6024 1746 6026 1752
rect 6026 1746 6058 1752
rect 6096 1746 6128 1752
rect 6128 1746 6130 1752
rect 6024 1683 6058 1707
rect 6096 1683 6130 1707
rect 6024 1673 6026 1683
rect 6026 1673 6058 1683
rect 6096 1673 6128 1683
rect 6128 1673 6130 1683
rect 6024 1614 6058 1634
rect 6096 1614 6130 1634
rect 6024 1600 6026 1614
rect 6026 1600 6058 1614
rect 6096 1600 6128 1614
rect 6128 1600 6130 1614
rect 6024 1545 6058 1561
rect 6096 1545 6130 1561
rect 6024 1527 6026 1545
rect 6026 1527 6058 1545
rect 6096 1527 6128 1545
rect 6128 1527 6130 1545
rect 6024 1476 6058 1488
rect 6096 1476 6130 1488
rect 6024 1454 6026 1476
rect 6026 1454 6058 1476
rect 6096 1454 6128 1476
rect 6128 1454 6130 1476
rect 6024 1407 6058 1415
rect 6096 1407 6130 1415
rect 6024 1381 6026 1407
rect 6026 1381 6058 1407
rect 6096 1381 6128 1407
rect 6128 1381 6130 1407
rect 6024 1338 6058 1342
rect 6096 1338 6130 1342
rect 6024 1308 6026 1338
rect 6026 1308 6058 1338
rect 6096 1308 6128 1338
rect 6128 1308 6130 1338
rect 6024 1235 6026 1269
rect 6026 1235 6058 1269
rect 6096 1235 6128 1269
rect 6128 1235 6130 1269
rect 6926 3719 6928 11233
rect 6928 3719 7030 11233
rect 7030 3719 7032 11233
rect 6926 3684 7032 3719
rect 6926 3650 6928 3684
rect 6928 3650 6962 3684
rect 6962 3650 6996 3684
rect 6996 3650 7030 3684
rect 7030 3650 7032 3684
rect 6926 3615 7032 3650
rect 6926 3581 6928 3615
rect 6928 3581 6962 3615
rect 6962 3581 6996 3615
rect 6996 3581 7030 3615
rect 7030 3581 7032 3615
rect 6926 3546 7032 3581
rect 6926 3512 6928 3546
rect 6928 3512 6962 3546
rect 6962 3512 6996 3546
rect 6996 3512 7030 3546
rect 7030 3512 7032 3546
rect 6926 3477 7032 3512
rect 6926 3443 6928 3477
rect 6928 3443 6962 3477
rect 6962 3443 6996 3477
rect 6996 3443 7030 3477
rect 7030 3443 7032 3477
rect 6926 3408 7032 3443
rect 6926 3374 6928 3408
rect 6928 3374 6962 3408
rect 6962 3374 6996 3408
rect 6996 3374 7030 3408
rect 7030 3374 7032 3408
rect 6926 3339 7032 3374
rect 6926 3305 6928 3339
rect 6928 3305 6962 3339
rect 6962 3305 6996 3339
rect 6996 3305 7030 3339
rect 7030 3305 7032 3339
rect 6926 3279 7032 3305
rect 6926 3236 6928 3240
rect 6928 3236 6960 3240
rect 6998 3236 7030 3240
rect 7030 3236 7032 3240
rect 6926 3206 6960 3236
rect 6998 3206 7032 3236
rect 6926 3133 6960 3167
rect 6998 3133 7032 3167
rect 6926 3063 6960 3094
rect 6998 3063 7032 3094
rect 6926 3060 6928 3063
rect 6928 3060 6960 3063
rect 6998 3060 7030 3063
rect 7030 3060 7032 3063
rect 6926 2994 6960 3021
rect 6998 2994 7032 3021
rect 6926 2987 6928 2994
rect 6928 2987 6960 2994
rect 6998 2987 7030 2994
rect 7030 2987 7032 2994
rect 6926 2925 6960 2948
rect 6998 2925 7032 2948
rect 6926 2914 6928 2925
rect 6928 2914 6960 2925
rect 6998 2914 7030 2925
rect 7030 2914 7032 2925
rect 6926 2856 6960 2875
rect 6998 2856 7032 2875
rect 6926 2841 6928 2856
rect 6928 2841 6960 2856
rect 6998 2841 7030 2856
rect 7030 2841 7032 2856
rect 6926 2787 6960 2802
rect 6998 2787 7032 2802
rect 6926 2768 6928 2787
rect 6928 2768 6960 2787
rect 6998 2768 7030 2787
rect 7030 2768 7032 2787
rect 6926 2718 6960 2729
rect 6998 2718 7032 2729
rect 6926 2695 6928 2718
rect 6928 2695 6960 2718
rect 6998 2695 7030 2718
rect 7030 2695 7032 2718
rect 6926 2649 6960 2656
rect 6998 2649 7032 2656
rect 6926 2622 6928 2649
rect 6928 2622 6960 2649
rect 6998 2622 7030 2649
rect 7030 2622 7032 2649
rect 6926 2580 6960 2583
rect 6998 2580 7032 2583
rect 6926 2549 6928 2580
rect 6928 2549 6960 2580
rect 6998 2549 7030 2580
rect 7030 2549 7032 2580
rect 6926 2477 6928 2510
rect 6928 2477 6960 2510
rect 6998 2477 7030 2510
rect 7030 2477 7032 2510
rect 6926 2476 6960 2477
rect 6998 2476 7032 2477
rect 6926 2408 6928 2437
rect 6928 2408 6960 2437
rect 6998 2408 7030 2437
rect 7030 2408 7032 2437
rect 6926 2403 6960 2408
rect 6998 2403 7032 2408
rect 6926 2339 6928 2364
rect 6928 2339 6960 2364
rect 6998 2339 7030 2364
rect 7030 2339 7032 2364
rect 6926 2330 6960 2339
rect 6998 2330 7032 2339
rect 6926 2270 6928 2291
rect 6928 2270 6960 2291
rect 6998 2270 7030 2291
rect 7030 2270 7032 2291
rect 6926 2257 6960 2270
rect 6998 2257 7032 2270
rect 6926 2201 6928 2218
rect 6928 2201 6960 2218
rect 6998 2201 7030 2218
rect 7030 2201 7032 2218
rect 6926 2184 6960 2201
rect 6998 2184 7032 2201
rect 6926 2132 6928 2145
rect 6928 2132 6960 2145
rect 6998 2132 7030 2145
rect 7030 2132 7032 2145
rect 6926 2111 6960 2132
rect 6998 2111 7032 2132
rect 6926 2063 6928 2072
rect 6928 2063 6960 2072
rect 6998 2063 7030 2072
rect 7030 2063 7032 2072
rect 6926 2038 6960 2063
rect 6998 2038 7032 2063
rect 6926 1994 6928 1999
rect 6928 1994 6960 1999
rect 6998 1994 7030 1999
rect 7030 1994 7032 1999
rect 6926 1965 6960 1994
rect 6998 1965 7032 1994
rect 6926 1925 6928 1926
rect 6928 1925 6960 1926
rect 6998 1925 7030 1926
rect 7030 1925 7032 1926
rect 6926 1892 6960 1925
rect 6998 1892 7032 1925
rect 6926 1821 6960 1853
rect 6998 1821 7032 1853
rect 6926 1819 6928 1821
rect 6928 1819 6960 1821
rect 6998 1819 7030 1821
rect 7030 1819 7032 1821
rect 6926 1752 6960 1780
rect 6998 1752 7032 1780
rect 6926 1746 6928 1752
rect 6928 1746 6960 1752
rect 6998 1746 7030 1752
rect 7030 1746 7032 1752
rect 6926 1683 6960 1707
rect 6998 1683 7032 1707
rect 6926 1673 6928 1683
rect 6928 1673 6960 1683
rect 6998 1673 7030 1683
rect 7030 1673 7032 1683
rect 6926 1614 6960 1634
rect 6998 1614 7032 1634
rect 6926 1600 6928 1614
rect 6928 1600 6960 1614
rect 6998 1600 7030 1614
rect 7030 1600 7032 1614
rect 6926 1545 6960 1561
rect 6998 1545 7032 1561
rect 6926 1527 6928 1545
rect 6928 1527 6960 1545
rect 6998 1527 7030 1545
rect 7030 1527 7032 1545
rect 6926 1476 6960 1488
rect 6998 1476 7032 1488
rect 6926 1454 6928 1476
rect 6928 1454 6960 1476
rect 6998 1454 7030 1476
rect 7030 1454 7032 1476
rect 6926 1407 6960 1415
rect 6998 1407 7032 1415
rect 6926 1381 6928 1407
rect 6928 1381 6960 1407
rect 6998 1381 7030 1407
rect 7030 1381 7032 1407
rect 6926 1338 6960 1342
rect 6998 1338 7032 1342
rect 6926 1308 6928 1338
rect 6928 1308 6960 1338
rect 6998 1308 7030 1338
rect 7030 1308 7032 1338
rect 6926 1235 6928 1269
rect 6928 1235 6960 1269
rect 6998 1235 7030 1269
rect 7030 1235 7032 1269
rect 7828 3719 7830 11233
rect 7830 3719 7932 11233
rect 7932 3719 7934 11233
rect 7828 3684 7934 3719
rect 7828 3650 7830 3684
rect 7830 3650 7864 3684
rect 7864 3650 7898 3684
rect 7898 3650 7932 3684
rect 7932 3650 7934 3684
rect 7828 3615 7934 3650
rect 7828 3581 7830 3615
rect 7830 3581 7864 3615
rect 7864 3581 7898 3615
rect 7898 3581 7932 3615
rect 7932 3581 7934 3615
rect 7828 3546 7934 3581
rect 7828 3512 7830 3546
rect 7830 3512 7864 3546
rect 7864 3512 7898 3546
rect 7898 3512 7932 3546
rect 7932 3512 7934 3546
rect 7828 3477 7934 3512
rect 7828 3443 7830 3477
rect 7830 3443 7864 3477
rect 7864 3443 7898 3477
rect 7898 3443 7932 3477
rect 7932 3443 7934 3477
rect 7828 3408 7934 3443
rect 7828 3374 7830 3408
rect 7830 3374 7864 3408
rect 7864 3374 7898 3408
rect 7898 3374 7932 3408
rect 7932 3374 7934 3408
rect 7828 3339 7934 3374
rect 7828 3305 7830 3339
rect 7830 3305 7864 3339
rect 7864 3305 7898 3339
rect 7898 3305 7932 3339
rect 7932 3305 7934 3339
rect 7828 3279 7934 3305
rect 7828 3236 7830 3240
rect 7830 3236 7862 3240
rect 7900 3236 7932 3240
rect 7932 3236 7934 3240
rect 7828 3206 7862 3236
rect 7900 3206 7934 3236
rect 7828 3133 7862 3167
rect 7900 3133 7934 3167
rect 7828 3063 7862 3094
rect 7900 3063 7934 3094
rect 7828 3060 7830 3063
rect 7830 3060 7862 3063
rect 7900 3060 7932 3063
rect 7932 3060 7934 3063
rect 7828 2994 7862 3021
rect 7900 2994 7934 3021
rect 7828 2987 7830 2994
rect 7830 2987 7862 2994
rect 7900 2987 7932 2994
rect 7932 2987 7934 2994
rect 7828 2925 7862 2948
rect 7900 2925 7934 2948
rect 7828 2914 7830 2925
rect 7830 2914 7862 2925
rect 7900 2914 7932 2925
rect 7932 2914 7934 2925
rect 7828 2856 7862 2875
rect 7900 2856 7934 2875
rect 7828 2841 7830 2856
rect 7830 2841 7862 2856
rect 7900 2841 7932 2856
rect 7932 2841 7934 2856
rect 7828 2787 7862 2802
rect 7900 2787 7934 2802
rect 7828 2768 7830 2787
rect 7830 2768 7862 2787
rect 7900 2768 7932 2787
rect 7932 2768 7934 2787
rect 7828 2718 7862 2729
rect 7900 2718 7934 2729
rect 7828 2695 7830 2718
rect 7830 2695 7862 2718
rect 7900 2695 7932 2718
rect 7932 2695 7934 2718
rect 7828 2649 7862 2656
rect 7900 2649 7934 2656
rect 7828 2622 7830 2649
rect 7830 2622 7862 2649
rect 7900 2622 7932 2649
rect 7932 2622 7934 2649
rect 7828 2580 7862 2583
rect 7900 2580 7934 2583
rect 7828 2549 7830 2580
rect 7830 2549 7862 2580
rect 7900 2549 7932 2580
rect 7932 2549 7934 2580
rect 7828 2477 7830 2510
rect 7830 2477 7862 2510
rect 7900 2477 7932 2510
rect 7932 2477 7934 2510
rect 7828 2476 7862 2477
rect 7900 2476 7934 2477
rect 7828 2408 7830 2437
rect 7830 2408 7862 2437
rect 7900 2408 7932 2437
rect 7932 2408 7934 2437
rect 7828 2403 7862 2408
rect 7900 2403 7934 2408
rect 7828 2339 7830 2364
rect 7830 2339 7862 2364
rect 7900 2339 7932 2364
rect 7932 2339 7934 2364
rect 7828 2330 7862 2339
rect 7900 2330 7934 2339
rect 7828 2270 7830 2291
rect 7830 2270 7862 2291
rect 7900 2270 7932 2291
rect 7932 2270 7934 2291
rect 7828 2257 7862 2270
rect 7900 2257 7934 2270
rect 7828 2201 7830 2218
rect 7830 2201 7862 2218
rect 7900 2201 7932 2218
rect 7932 2201 7934 2218
rect 7828 2184 7862 2201
rect 7900 2184 7934 2201
rect 7828 2132 7830 2145
rect 7830 2132 7862 2145
rect 7900 2132 7932 2145
rect 7932 2132 7934 2145
rect 7828 2111 7862 2132
rect 7900 2111 7934 2132
rect 7828 2063 7830 2072
rect 7830 2063 7862 2072
rect 7900 2063 7932 2072
rect 7932 2063 7934 2072
rect 7828 2038 7862 2063
rect 7900 2038 7934 2063
rect 7828 1994 7830 1999
rect 7830 1994 7862 1999
rect 7900 1994 7932 1999
rect 7932 1994 7934 1999
rect 7828 1965 7862 1994
rect 7900 1965 7934 1994
rect 7828 1925 7830 1926
rect 7830 1925 7862 1926
rect 7900 1925 7932 1926
rect 7932 1925 7934 1926
rect 7828 1892 7862 1925
rect 7900 1892 7934 1925
rect 7828 1821 7862 1853
rect 7900 1821 7934 1853
rect 7828 1819 7830 1821
rect 7830 1819 7862 1821
rect 7900 1819 7932 1821
rect 7932 1819 7934 1821
rect 7828 1752 7862 1780
rect 7900 1752 7934 1780
rect 7828 1746 7830 1752
rect 7830 1746 7862 1752
rect 7900 1746 7932 1752
rect 7932 1746 7934 1752
rect 7828 1683 7862 1707
rect 7900 1683 7934 1707
rect 7828 1673 7830 1683
rect 7830 1673 7862 1683
rect 7900 1673 7932 1683
rect 7932 1673 7934 1683
rect 7828 1614 7862 1634
rect 7900 1614 7934 1634
rect 7828 1600 7830 1614
rect 7830 1600 7862 1614
rect 7900 1600 7932 1614
rect 7932 1600 7934 1614
rect 7828 1545 7862 1561
rect 7900 1545 7934 1561
rect 7828 1527 7830 1545
rect 7830 1527 7862 1545
rect 7900 1527 7932 1545
rect 7932 1527 7934 1545
rect 7828 1476 7862 1488
rect 7900 1476 7934 1488
rect 7828 1454 7830 1476
rect 7830 1454 7862 1476
rect 7900 1454 7932 1476
rect 7932 1454 7934 1476
rect 7828 1407 7862 1415
rect 7900 1407 7934 1415
rect 7828 1381 7830 1407
rect 7830 1381 7862 1407
rect 7900 1381 7932 1407
rect 7932 1381 7934 1407
rect 7828 1338 7862 1342
rect 7900 1338 7934 1342
rect 7828 1308 7830 1338
rect 7830 1308 7862 1338
rect 7900 1308 7932 1338
rect 7932 1308 7934 1338
rect 7828 1235 7830 1269
rect 7830 1235 7862 1269
rect 7900 1235 7932 1269
rect 7932 1235 7934 1269
rect 8730 3719 8732 11233
rect 8732 3719 8834 11233
rect 8834 3719 8836 11233
rect 8730 3684 8836 3719
rect 8730 3650 8732 3684
rect 8732 3650 8766 3684
rect 8766 3650 8800 3684
rect 8800 3650 8834 3684
rect 8834 3650 8836 3684
rect 8730 3615 8836 3650
rect 8730 3581 8732 3615
rect 8732 3581 8766 3615
rect 8766 3581 8800 3615
rect 8800 3581 8834 3615
rect 8834 3581 8836 3615
rect 8730 3546 8836 3581
rect 8730 3512 8732 3546
rect 8732 3512 8766 3546
rect 8766 3512 8800 3546
rect 8800 3512 8834 3546
rect 8834 3512 8836 3546
rect 8730 3477 8836 3512
rect 8730 3443 8732 3477
rect 8732 3443 8766 3477
rect 8766 3443 8800 3477
rect 8800 3443 8834 3477
rect 8834 3443 8836 3477
rect 8730 3408 8836 3443
rect 8730 3374 8732 3408
rect 8732 3374 8766 3408
rect 8766 3374 8800 3408
rect 8800 3374 8834 3408
rect 8834 3374 8836 3408
rect 8730 3339 8836 3374
rect 8730 3305 8732 3339
rect 8732 3305 8766 3339
rect 8766 3305 8800 3339
rect 8800 3305 8834 3339
rect 8834 3305 8836 3339
rect 8730 3279 8836 3305
rect 8730 3236 8732 3240
rect 8732 3236 8764 3240
rect 8802 3236 8834 3240
rect 8834 3236 8836 3240
rect 8730 3206 8764 3236
rect 8802 3206 8836 3236
rect 8730 3133 8764 3167
rect 8802 3133 8836 3167
rect 8730 3063 8764 3094
rect 8802 3063 8836 3094
rect 8730 3060 8732 3063
rect 8732 3060 8764 3063
rect 8802 3060 8834 3063
rect 8834 3060 8836 3063
rect 8730 2994 8764 3021
rect 8802 2994 8836 3021
rect 8730 2987 8732 2994
rect 8732 2987 8764 2994
rect 8802 2987 8834 2994
rect 8834 2987 8836 2994
rect 8730 2925 8764 2948
rect 8802 2925 8836 2948
rect 8730 2914 8732 2925
rect 8732 2914 8764 2925
rect 8802 2914 8834 2925
rect 8834 2914 8836 2925
rect 8730 2856 8764 2875
rect 8802 2856 8836 2875
rect 8730 2841 8732 2856
rect 8732 2841 8764 2856
rect 8802 2841 8834 2856
rect 8834 2841 8836 2856
rect 8730 2787 8764 2802
rect 8802 2787 8836 2802
rect 8730 2768 8732 2787
rect 8732 2768 8764 2787
rect 8802 2768 8834 2787
rect 8834 2768 8836 2787
rect 8730 2718 8764 2729
rect 8802 2718 8836 2729
rect 8730 2695 8732 2718
rect 8732 2695 8764 2718
rect 8802 2695 8834 2718
rect 8834 2695 8836 2718
rect 8730 2649 8764 2656
rect 8802 2649 8836 2656
rect 8730 2622 8732 2649
rect 8732 2622 8764 2649
rect 8802 2622 8834 2649
rect 8834 2622 8836 2649
rect 8730 2580 8764 2583
rect 8802 2580 8836 2583
rect 8730 2549 8732 2580
rect 8732 2549 8764 2580
rect 8802 2549 8834 2580
rect 8834 2549 8836 2580
rect 8730 2477 8732 2510
rect 8732 2477 8764 2510
rect 8802 2477 8834 2510
rect 8834 2477 8836 2510
rect 8730 2476 8764 2477
rect 8802 2476 8836 2477
rect 8730 2408 8732 2437
rect 8732 2408 8764 2437
rect 8802 2408 8834 2437
rect 8834 2408 8836 2437
rect 8730 2403 8764 2408
rect 8802 2403 8836 2408
rect 8730 2339 8732 2364
rect 8732 2339 8764 2364
rect 8802 2339 8834 2364
rect 8834 2339 8836 2364
rect 8730 2330 8764 2339
rect 8802 2330 8836 2339
rect 8730 2270 8732 2291
rect 8732 2270 8764 2291
rect 8802 2270 8834 2291
rect 8834 2270 8836 2291
rect 8730 2257 8764 2270
rect 8802 2257 8836 2270
rect 8730 2201 8732 2218
rect 8732 2201 8764 2218
rect 8802 2201 8834 2218
rect 8834 2201 8836 2218
rect 8730 2184 8764 2201
rect 8802 2184 8836 2201
rect 8730 2132 8732 2145
rect 8732 2132 8764 2145
rect 8802 2132 8834 2145
rect 8834 2132 8836 2145
rect 8730 2111 8764 2132
rect 8802 2111 8836 2132
rect 8730 2063 8732 2072
rect 8732 2063 8764 2072
rect 8802 2063 8834 2072
rect 8834 2063 8836 2072
rect 8730 2038 8764 2063
rect 8802 2038 8836 2063
rect 8730 1994 8732 1999
rect 8732 1994 8764 1999
rect 8802 1994 8834 1999
rect 8834 1994 8836 1999
rect 8730 1965 8764 1994
rect 8802 1965 8836 1994
rect 8730 1925 8732 1926
rect 8732 1925 8764 1926
rect 8802 1925 8834 1926
rect 8834 1925 8836 1926
rect 8730 1892 8764 1925
rect 8802 1892 8836 1925
rect 8730 1821 8764 1853
rect 8802 1821 8836 1853
rect 8730 1819 8732 1821
rect 8732 1819 8764 1821
rect 8802 1819 8834 1821
rect 8834 1819 8836 1821
rect 8730 1752 8764 1780
rect 8802 1752 8836 1780
rect 8730 1746 8732 1752
rect 8732 1746 8764 1752
rect 8802 1746 8834 1752
rect 8834 1746 8836 1752
rect 8730 1683 8764 1707
rect 8802 1683 8836 1707
rect 8730 1673 8732 1683
rect 8732 1673 8764 1683
rect 8802 1673 8834 1683
rect 8834 1673 8836 1683
rect 8730 1614 8764 1634
rect 8802 1614 8836 1634
rect 8730 1600 8732 1614
rect 8732 1600 8764 1614
rect 8802 1600 8834 1614
rect 8834 1600 8836 1614
rect 8730 1545 8764 1561
rect 8802 1545 8836 1561
rect 8730 1527 8732 1545
rect 8732 1527 8764 1545
rect 8802 1527 8834 1545
rect 8834 1527 8836 1545
rect 8730 1476 8764 1488
rect 8802 1476 8836 1488
rect 8730 1454 8732 1476
rect 8732 1454 8764 1476
rect 8802 1454 8834 1476
rect 8834 1454 8836 1476
rect 8730 1407 8764 1415
rect 8802 1407 8836 1415
rect 8730 1381 8732 1407
rect 8732 1381 8764 1407
rect 8802 1381 8834 1407
rect 8834 1381 8836 1407
rect 8730 1338 8764 1342
rect 8802 1338 8836 1342
rect 8730 1308 8732 1338
rect 8732 1308 8764 1338
rect 8802 1308 8834 1338
rect 8834 1308 8836 1338
rect 8730 1235 8732 1269
rect 8732 1235 8764 1269
rect 8802 1235 8834 1269
rect 8834 1235 8836 1269
rect 9632 3719 9634 11233
rect 9634 3719 9736 11233
rect 9736 3719 9738 11233
rect 9632 3684 9738 3719
rect 9632 3650 9634 3684
rect 9634 3650 9668 3684
rect 9668 3650 9702 3684
rect 9702 3650 9736 3684
rect 9736 3650 9738 3684
rect 9632 3615 9738 3650
rect 9632 3581 9634 3615
rect 9634 3581 9668 3615
rect 9668 3581 9702 3615
rect 9702 3581 9736 3615
rect 9736 3581 9738 3615
rect 9632 3546 9738 3581
rect 9632 3512 9634 3546
rect 9634 3512 9668 3546
rect 9668 3512 9702 3546
rect 9702 3512 9736 3546
rect 9736 3512 9738 3546
rect 9632 3477 9738 3512
rect 9632 3443 9634 3477
rect 9634 3443 9668 3477
rect 9668 3443 9702 3477
rect 9702 3443 9736 3477
rect 9736 3443 9738 3477
rect 9632 3408 9738 3443
rect 9632 3374 9634 3408
rect 9634 3374 9668 3408
rect 9668 3374 9702 3408
rect 9702 3374 9736 3408
rect 9736 3374 9738 3408
rect 9632 3339 9738 3374
rect 9632 3305 9634 3339
rect 9634 3305 9668 3339
rect 9668 3305 9702 3339
rect 9702 3305 9736 3339
rect 9736 3305 9738 3339
rect 9632 3279 9738 3305
rect 9632 3236 9634 3240
rect 9634 3236 9666 3240
rect 9704 3236 9736 3240
rect 9736 3236 9738 3240
rect 9632 3206 9666 3236
rect 9704 3206 9738 3236
rect 9632 3133 9666 3167
rect 9704 3133 9738 3167
rect 9632 3063 9666 3094
rect 9704 3063 9738 3094
rect 9632 3060 9634 3063
rect 9634 3060 9666 3063
rect 9704 3060 9736 3063
rect 9736 3060 9738 3063
rect 9632 2994 9666 3021
rect 9704 2994 9738 3021
rect 9632 2987 9634 2994
rect 9634 2987 9666 2994
rect 9704 2987 9736 2994
rect 9736 2987 9738 2994
rect 9632 2925 9666 2948
rect 9704 2925 9738 2948
rect 9632 2914 9634 2925
rect 9634 2914 9666 2925
rect 9704 2914 9736 2925
rect 9736 2914 9738 2925
rect 9632 2856 9666 2875
rect 9704 2856 9738 2875
rect 9632 2841 9634 2856
rect 9634 2841 9666 2856
rect 9704 2841 9736 2856
rect 9736 2841 9738 2856
rect 9632 2787 9666 2802
rect 9704 2787 9738 2802
rect 9632 2768 9634 2787
rect 9634 2768 9666 2787
rect 9704 2768 9736 2787
rect 9736 2768 9738 2787
rect 9632 2718 9666 2729
rect 9704 2718 9738 2729
rect 9632 2695 9634 2718
rect 9634 2695 9666 2718
rect 9704 2695 9736 2718
rect 9736 2695 9738 2718
rect 9632 2649 9666 2656
rect 9704 2649 9738 2656
rect 9632 2622 9634 2649
rect 9634 2622 9666 2649
rect 9704 2622 9736 2649
rect 9736 2622 9738 2649
rect 9632 2580 9666 2583
rect 9704 2580 9738 2583
rect 9632 2549 9634 2580
rect 9634 2549 9666 2580
rect 9704 2549 9736 2580
rect 9736 2549 9738 2580
rect 9632 2477 9634 2510
rect 9634 2477 9666 2510
rect 9704 2477 9736 2510
rect 9736 2477 9738 2510
rect 9632 2476 9666 2477
rect 9704 2476 9738 2477
rect 9632 2408 9634 2437
rect 9634 2408 9666 2437
rect 9704 2408 9736 2437
rect 9736 2408 9738 2437
rect 9632 2403 9666 2408
rect 9704 2403 9738 2408
rect 9632 2339 9634 2364
rect 9634 2339 9666 2364
rect 9704 2339 9736 2364
rect 9736 2339 9738 2364
rect 9632 2330 9666 2339
rect 9704 2330 9738 2339
rect 9632 2270 9634 2291
rect 9634 2270 9666 2291
rect 9704 2270 9736 2291
rect 9736 2270 9738 2291
rect 9632 2257 9666 2270
rect 9704 2257 9738 2270
rect 9632 2201 9634 2218
rect 9634 2201 9666 2218
rect 9704 2201 9736 2218
rect 9736 2201 9738 2218
rect 9632 2184 9666 2201
rect 9704 2184 9738 2201
rect 9632 2132 9634 2145
rect 9634 2132 9666 2145
rect 9704 2132 9736 2145
rect 9736 2132 9738 2145
rect 9632 2111 9666 2132
rect 9704 2111 9738 2132
rect 9632 2063 9634 2072
rect 9634 2063 9666 2072
rect 9704 2063 9736 2072
rect 9736 2063 9738 2072
rect 9632 2038 9666 2063
rect 9704 2038 9738 2063
rect 9632 1994 9634 1999
rect 9634 1994 9666 1999
rect 9704 1994 9736 1999
rect 9736 1994 9738 1999
rect 9632 1965 9666 1994
rect 9704 1965 9738 1994
rect 9632 1925 9634 1926
rect 9634 1925 9666 1926
rect 9704 1925 9736 1926
rect 9736 1925 9738 1926
rect 9632 1892 9666 1925
rect 9704 1892 9738 1925
rect 9632 1821 9666 1853
rect 9704 1821 9738 1853
rect 9632 1819 9634 1821
rect 9634 1819 9666 1821
rect 9704 1819 9736 1821
rect 9736 1819 9738 1821
rect 9632 1752 9666 1780
rect 9704 1752 9738 1780
rect 9632 1746 9634 1752
rect 9634 1746 9666 1752
rect 9704 1746 9736 1752
rect 9736 1746 9738 1752
rect 9632 1683 9666 1707
rect 9704 1683 9738 1707
rect 9632 1673 9634 1683
rect 9634 1673 9666 1683
rect 9704 1673 9736 1683
rect 9736 1673 9738 1683
rect 9632 1614 9666 1634
rect 9704 1614 9738 1634
rect 9632 1600 9634 1614
rect 9634 1600 9666 1614
rect 9704 1600 9736 1614
rect 9736 1600 9738 1614
rect 9632 1545 9666 1561
rect 9704 1545 9738 1561
rect 9632 1527 9634 1545
rect 9634 1527 9666 1545
rect 9704 1527 9736 1545
rect 9736 1527 9738 1545
rect 9632 1476 9666 1488
rect 9704 1476 9738 1488
rect 9632 1454 9634 1476
rect 9634 1454 9666 1476
rect 9704 1454 9736 1476
rect 9736 1454 9738 1476
rect 9632 1407 9666 1415
rect 9704 1407 9738 1415
rect 9632 1381 9634 1407
rect 9634 1381 9666 1407
rect 9704 1381 9736 1407
rect 9736 1381 9738 1407
rect 9632 1338 9666 1342
rect 9704 1338 9738 1342
rect 9632 1308 9634 1338
rect 9634 1308 9666 1338
rect 9704 1308 9736 1338
rect 9736 1308 9738 1338
rect 9632 1235 9634 1269
rect 9634 1235 9666 1269
rect 9704 1235 9736 1269
rect 9736 1235 9738 1269
rect 10534 3719 10536 11233
rect 10536 3719 10638 11233
rect 10638 3719 10640 11233
rect 10534 3684 10640 3719
rect 10534 3650 10536 3684
rect 10536 3650 10570 3684
rect 10570 3650 10604 3684
rect 10604 3650 10638 3684
rect 10638 3650 10640 3684
rect 10534 3615 10640 3650
rect 10534 3581 10536 3615
rect 10536 3581 10570 3615
rect 10570 3581 10604 3615
rect 10604 3581 10638 3615
rect 10638 3581 10640 3615
rect 10534 3546 10640 3581
rect 10534 3512 10536 3546
rect 10536 3512 10570 3546
rect 10570 3512 10604 3546
rect 10604 3512 10638 3546
rect 10638 3512 10640 3546
rect 10534 3477 10640 3512
rect 10534 3443 10536 3477
rect 10536 3443 10570 3477
rect 10570 3443 10604 3477
rect 10604 3443 10638 3477
rect 10638 3443 10640 3477
rect 10534 3408 10640 3443
rect 10534 3374 10536 3408
rect 10536 3374 10570 3408
rect 10570 3374 10604 3408
rect 10604 3374 10638 3408
rect 10638 3374 10640 3408
rect 10534 3339 10640 3374
rect 10534 3305 10536 3339
rect 10536 3305 10570 3339
rect 10570 3305 10604 3339
rect 10604 3305 10638 3339
rect 10638 3305 10640 3339
rect 10534 3279 10640 3305
rect 10534 3236 10536 3240
rect 10536 3236 10568 3240
rect 10606 3236 10638 3240
rect 10638 3236 10640 3240
rect 10534 3206 10568 3236
rect 10606 3206 10640 3236
rect 10534 3133 10568 3167
rect 10606 3133 10640 3167
rect 10534 3063 10568 3094
rect 10606 3063 10640 3094
rect 10534 3060 10536 3063
rect 10536 3060 10568 3063
rect 10606 3060 10638 3063
rect 10638 3060 10640 3063
rect 10534 2994 10568 3021
rect 10606 2994 10640 3021
rect 10534 2987 10536 2994
rect 10536 2987 10568 2994
rect 10606 2987 10638 2994
rect 10638 2987 10640 2994
rect 10534 2925 10568 2948
rect 10606 2925 10640 2948
rect 10534 2914 10536 2925
rect 10536 2914 10568 2925
rect 10606 2914 10638 2925
rect 10638 2914 10640 2925
rect 10534 2856 10568 2875
rect 10606 2856 10640 2875
rect 10534 2841 10536 2856
rect 10536 2841 10568 2856
rect 10606 2841 10638 2856
rect 10638 2841 10640 2856
rect 10534 2787 10568 2802
rect 10606 2787 10640 2802
rect 10534 2768 10536 2787
rect 10536 2768 10568 2787
rect 10606 2768 10638 2787
rect 10638 2768 10640 2787
rect 10534 2718 10568 2729
rect 10606 2718 10640 2729
rect 10534 2695 10536 2718
rect 10536 2695 10568 2718
rect 10606 2695 10638 2718
rect 10638 2695 10640 2718
rect 10534 2649 10568 2656
rect 10606 2649 10640 2656
rect 10534 2622 10536 2649
rect 10536 2622 10568 2649
rect 10606 2622 10638 2649
rect 10638 2622 10640 2649
rect 10534 2580 10568 2583
rect 10606 2580 10640 2583
rect 10534 2549 10536 2580
rect 10536 2549 10568 2580
rect 10606 2549 10638 2580
rect 10638 2549 10640 2580
rect 10534 2477 10536 2510
rect 10536 2477 10568 2510
rect 10606 2477 10638 2510
rect 10638 2477 10640 2510
rect 10534 2476 10568 2477
rect 10606 2476 10640 2477
rect 10534 2408 10536 2437
rect 10536 2408 10568 2437
rect 10606 2408 10638 2437
rect 10638 2408 10640 2437
rect 10534 2403 10568 2408
rect 10606 2403 10640 2408
rect 10534 2339 10536 2364
rect 10536 2339 10568 2364
rect 10606 2339 10638 2364
rect 10638 2339 10640 2364
rect 10534 2330 10568 2339
rect 10606 2330 10640 2339
rect 10534 2270 10536 2291
rect 10536 2270 10568 2291
rect 10606 2270 10638 2291
rect 10638 2270 10640 2291
rect 10534 2257 10568 2270
rect 10606 2257 10640 2270
rect 10534 2201 10536 2218
rect 10536 2201 10568 2218
rect 10606 2201 10638 2218
rect 10638 2201 10640 2218
rect 10534 2184 10568 2201
rect 10606 2184 10640 2201
rect 10534 2132 10536 2145
rect 10536 2132 10568 2145
rect 10606 2132 10638 2145
rect 10638 2132 10640 2145
rect 10534 2111 10568 2132
rect 10606 2111 10640 2132
rect 10534 2063 10536 2072
rect 10536 2063 10568 2072
rect 10606 2063 10638 2072
rect 10638 2063 10640 2072
rect 10534 2038 10568 2063
rect 10606 2038 10640 2063
rect 10534 1994 10536 1999
rect 10536 1994 10568 1999
rect 10606 1994 10638 1999
rect 10638 1994 10640 1999
rect 10534 1965 10568 1994
rect 10606 1965 10640 1994
rect 10534 1925 10536 1926
rect 10536 1925 10568 1926
rect 10606 1925 10638 1926
rect 10638 1925 10640 1926
rect 10534 1892 10568 1925
rect 10606 1892 10640 1925
rect 10534 1821 10568 1853
rect 10606 1821 10640 1853
rect 10534 1819 10536 1821
rect 10536 1819 10568 1821
rect 10606 1819 10638 1821
rect 10638 1819 10640 1821
rect 10534 1752 10568 1780
rect 10606 1752 10640 1780
rect 10534 1746 10536 1752
rect 10536 1746 10568 1752
rect 10606 1746 10638 1752
rect 10638 1746 10640 1752
rect 10534 1683 10568 1707
rect 10606 1683 10640 1707
rect 10534 1673 10536 1683
rect 10536 1673 10568 1683
rect 10606 1673 10638 1683
rect 10638 1673 10640 1683
rect 10534 1614 10568 1634
rect 10606 1614 10640 1634
rect 10534 1600 10536 1614
rect 10536 1600 10568 1614
rect 10606 1600 10638 1614
rect 10638 1600 10640 1614
rect 10534 1545 10568 1561
rect 10606 1545 10640 1561
rect 10534 1527 10536 1545
rect 10536 1527 10568 1545
rect 10606 1527 10638 1545
rect 10638 1527 10640 1545
rect 10534 1476 10568 1488
rect 10606 1476 10640 1488
rect 10534 1454 10536 1476
rect 10536 1454 10568 1476
rect 10606 1454 10638 1476
rect 10638 1454 10640 1476
rect 10534 1407 10568 1415
rect 10606 1407 10640 1415
rect 10534 1381 10536 1407
rect 10536 1381 10568 1407
rect 10606 1381 10638 1407
rect 10638 1381 10640 1407
rect 10534 1338 10568 1342
rect 10606 1338 10640 1342
rect 10534 1308 10536 1338
rect 10536 1308 10568 1338
rect 10606 1308 10638 1338
rect 10638 1308 10640 1338
rect 10534 1235 10536 1269
rect 10536 1235 10568 1269
rect 10606 1235 10638 1269
rect 10638 1235 10640 1269
rect 11436 3719 11438 11233
rect 11438 3719 11540 11233
rect 11540 3719 11542 11233
rect 11436 3684 11542 3719
rect 11436 3650 11438 3684
rect 11438 3650 11472 3684
rect 11472 3650 11506 3684
rect 11506 3650 11540 3684
rect 11540 3650 11542 3684
rect 11436 3615 11542 3650
rect 11436 3581 11438 3615
rect 11438 3581 11472 3615
rect 11472 3581 11506 3615
rect 11506 3581 11540 3615
rect 11540 3581 11542 3615
rect 11436 3546 11542 3581
rect 11436 3512 11438 3546
rect 11438 3512 11472 3546
rect 11472 3512 11506 3546
rect 11506 3512 11540 3546
rect 11540 3512 11542 3546
rect 11436 3477 11542 3512
rect 11436 3443 11438 3477
rect 11438 3443 11472 3477
rect 11472 3443 11506 3477
rect 11506 3443 11540 3477
rect 11540 3443 11542 3477
rect 11436 3408 11542 3443
rect 11436 3374 11438 3408
rect 11438 3374 11472 3408
rect 11472 3374 11506 3408
rect 11506 3374 11540 3408
rect 11540 3374 11542 3408
rect 11436 3339 11542 3374
rect 11436 3305 11438 3339
rect 11438 3305 11472 3339
rect 11472 3305 11506 3339
rect 11506 3305 11540 3339
rect 11540 3305 11542 3339
rect 11436 3279 11542 3305
rect 11436 3236 11438 3240
rect 11438 3236 11470 3240
rect 11508 3236 11540 3240
rect 11540 3236 11542 3240
rect 11436 3206 11470 3236
rect 11508 3206 11542 3236
rect 11436 3133 11470 3167
rect 11508 3133 11542 3167
rect 11436 3063 11470 3094
rect 11508 3063 11542 3094
rect 11436 3060 11438 3063
rect 11438 3060 11470 3063
rect 11508 3060 11540 3063
rect 11540 3060 11542 3063
rect 11436 2994 11470 3021
rect 11508 2994 11542 3021
rect 11436 2987 11438 2994
rect 11438 2987 11470 2994
rect 11508 2987 11540 2994
rect 11540 2987 11542 2994
rect 11436 2925 11470 2948
rect 11508 2925 11542 2948
rect 11436 2914 11438 2925
rect 11438 2914 11470 2925
rect 11508 2914 11540 2925
rect 11540 2914 11542 2925
rect 11436 2856 11470 2875
rect 11508 2856 11542 2875
rect 11436 2841 11438 2856
rect 11438 2841 11470 2856
rect 11508 2841 11540 2856
rect 11540 2841 11542 2856
rect 11436 2787 11470 2802
rect 11508 2787 11542 2802
rect 11436 2768 11438 2787
rect 11438 2768 11470 2787
rect 11508 2768 11540 2787
rect 11540 2768 11542 2787
rect 11436 2718 11470 2729
rect 11508 2718 11542 2729
rect 11436 2695 11438 2718
rect 11438 2695 11470 2718
rect 11508 2695 11540 2718
rect 11540 2695 11542 2718
rect 11436 2649 11470 2656
rect 11508 2649 11542 2656
rect 11436 2622 11438 2649
rect 11438 2622 11470 2649
rect 11508 2622 11540 2649
rect 11540 2622 11542 2649
rect 11436 2580 11470 2583
rect 11508 2580 11542 2583
rect 11436 2549 11438 2580
rect 11438 2549 11470 2580
rect 11508 2549 11540 2580
rect 11540 2549 11542 2580
rect 11436 2477 11438 2510
rect 11438 2477 11470 2510
rect 11508 2477 11540 2510
rect 11540 2477 11542 2510
rect 11436 2476 11470 2477
rect 11508 2476 11542 2477
rect 11436 2408 11438 2437
rect 11438 2408 11470 2437
rect 11508 2408 11540 2437
rect 11540 2408 11542 2437
rect 11436 2403 11470 2408
rect 11508 2403 11542 2408
rect 11436 2339 11438 2364
rect 11438 2339 11470 2364
rect 11508 2339 11540 2364
rect 11540 2339 11542 2364
rect 11436 2330 11470 2339
rect 11508 2330 11542 2339
rect 11436 2270 11438 2291
rect 11438 2270 11470 2291
rect 11508 2270 11540 2291
rect 11540 2270 11542 2291
rect 11436 2257 11470 2270
rect 11508 2257 11542 2270
rect 11436 2201 11438 2218
rect 11438 2201 11470 2218
rect 11508 2201 11540 2218
rect 11540 2201 11542 2218
rect 11436 2184 11470 2201
rect 11508 2184 11542 2201
rect 11436 2132 11438 2145
rect 11438 2132 11470 2145
rect 11508 2132 11540 2145
rect 11540 2132 11542 2145
rect 11436 2111 11470 2132
rect 11508 2111 11542 2132
rect 11436 2063 11438 2072
rect 11438 2063 11470 2072
rect 11508 2063 11540 2072
rect 11540 2063 11542 2072
rect 11436 2038 11470 2063
rect 11508 2038 11542 2063
rect 11436 1994 11438 1999
rect 11438 1994 11470 1999
rect 11508 1994 11540 1999
rect 11540 1994 11542 1999
rect 11436 1965 11470 1994
rect 11508 1965 11542 1994
rect 11436 1925 11438 1926
rect 11438 1925 11470 1926
rect 11508 1925 11540 1926
rect 11540 1925 11542 1926
rect 11436 1892 11470 1925
rect 11508 1892 11542 1925
rect 11436 1821 11470 1853
rect 11508 1821 11542 1853
rect 11436 1819 11438 1821
rect 11438 1819 11470 1821
rect 11508 1819 11540 1821
rect 11540 1819 11542 1821
rect 11436 1752 11470 1780
rect 11508 1752 11542 1780
rect 11436 1746 11438 1752
rect 11438 1746 11470 1752
rect 11508 1746 11540 1752
rect 11540 1746 11542 1752
rect 11436 1683 11470 1707
rect 11508 1683 11542 1707
rect 11436 1673 11438 1683
rect 11438 1673 11470 1683
rect 11508 1673 11540 1683
rect 11540 1673 11542 1683
rect 11436 1614 11470 1634
rect 11508 1614 11542 1634
rect 11436 1600 11438 1614
rect 11438 1600 11470 1614
rect 11508 1600 11540 1614
rect 11540 1600 11542 1614
rect 11436 1545 11470 1561
rect 11508 1545 11542 1561
rect 11436 1527 11438 1545
rect 11438 1527 11470 1545
rect 11508 1527 11540 1545
rect 11540 1527 11542 1545
rect 11436 1476 11470 1488
rect 11508 1476 11542 1488
rect 11436 1454 11438 1476
rect 11438 1454 11470 1476
rect 11508 1454 11540 1476
rect 11540 1454 11542 1476
rect 11436 1407 11470 1415
rect 11508 1407 11542 1415
rect 11436 1381 11438 1407
rect 11438 1381 11470 1407
rect 11508 1381 11540 1407
rect 11540 1381 11542 1407
rect 11436 1338 11470 1342
rect 11508 1338 11542 1342
rect 11436 1308 11438 1338
rect 11438 1308 11470 1338
rect 11508 1308 11540 1338
rect 11540 1308 11542 1338
rect 11436 1235 11438 1269
rect 11438 1235 11470 1269
rect 11508 1235 11540 1269
rect 11540 1235 11542 1269
rect 12338 3719 12340 11233
rect 12340 3719 12442 11233
rect 12442 3719 12444 11233
rect 12338 3684 12444 3719
rect 12338 3650 12340 3684
rect 12340 3650 12374 3684
rect 12374 3650 12408 3684
rect 12408 3650 12442 3684
rect 12442 3650 12444 3684
rect 12338 3615 12444 3650
rect 12338 3581 12340 3615
rect 12340 3581 12374 3615
rect 12374 3581 12408 3615
rect 12408 3581 12442 3615
rect 12442 3581 12444 3615
rect 12338 3546 12444 3581
rect 12338 3512 12340 3546
rect 12340 3512 12374 3546
rect 12374 3512 12408 3546
rect 12408 3512 12442 3546
rect 12442 3512 12444 3546
rect 12338 3477 12444 3512
rect 12338 3443 12340 3477
rect 12340 3443 12374 3477
rect 12374 3443 12408 3477
rect 12408 3443 12442 3477
rect 12442 3443 12444 3477
rect 12338 3408 12444 3443
rect 12338 3374 12340 3408
rect 12340 3374 12374 3408
rect 12374 3374 12408 3408
rect 12408 3374 12442 3408
rect 12442 3374 12444 3408
rect 12338 3339 12444 3374
rect 12338 3305 12340 3339
rect 12340 3305 12374 3339
rect 12374 3305 12408 3339
rect 12408 3305 12442 3339
rect 12442 3305 12444 3339
rect 12338 3279 12444 3305
rect 12338 3236 12340 3240
rect 12340 3236 12372 3240
rect 12410 3236 12442 3240
rect 12442 3236 12444 3240
rect 12338 3206 12372 3236
rect 12410 3206 12444 3236
rect 12338 3133 12372 3167
rect 12410 3133 12444 3167
rect 12338 3063 12372 3094
rect 12410 3063 12444 3094
rect 12338 3060 12340 3063
rect 12340 3060 12372 3063
rect 12410 3060 12442 3063
rect 12442 3060 12444 3063
rect 12338 2994 12372 3021
rect 12410 2994 12444 3021
rect 12338 2987 12340 2994
rect 12340 2987 12372 2994
rect 12410 2987 12442 2994
rect 12442 2987 12444 2994
rect 12338 2925 12372 2948
rect 12410 2925 12444 2948
rect 12338 2914 12340 2925
rect 12340 2914 12372 2925
rect 12410 2914 12442 2925
rect 12442 2914 12444 2925
rect 12338 2856 12372 2875
rect 12410 2856 12444 2875
rect 12338 2841 12340 2856
rect 12340 2841 12372 2856
rect 12410 2841 12442 2856
rect 12442 2841 12444 2856
rect 12338 2787 12372 2802
rect 12410 2787 12444 2802
rect 12338 2768 12340 2787
rect 12340 2768 12372 2787
rect 12410 2768 12442 2787
rect 12442 2768 12444 2787
rect 12338 2718 12372 2729
rect 12410 2718 12444 2729
rect 12338 2695 12340 2718
rect 12340 2695 12372 2718
rect 12410 2695 12442 2718
rect 12442 2695 12444 2718
rect 12338 2649 12372 2656
rect 12410 2649 12444 2656
rect 12338 2622 12340 2649
rect 12340 2622 12372 2649
rect 12410 2622 12442 2649
rect 12442 2622 12444 2649
rect 12338 2580 12372 2583
rect 12410 2580 12444 2583
rect 12338 2549 12340 2580
rect 12340 2549 12372 2580
rect 12410 2549 12442 2580
rect 12442 2549 12444 2580
rect 12338 2477 12340 2510
rect 12340 2477 12372 2510
rect 12410 2477 12442 2510
rect 12442 2477 12444 2510
rect 12338 2476 12372 2477
rect 12410 2476 12444 2477
rect 12338 2408 12340 2437
rect 12340 2408 12372 2437
rect 12410 2408 12442 2437
rect 12442 2408 12444 2437
rect 12338 2403 12372 2408
rect 12410 2403 12444 2408
rect 12338 2339 12340 2364
rect 12340 2339 12372 2364
rect 12410 2339 12442 2364
rect 12442 2339 12444 2364
rect 12338 2330 12372 2339
rect 12410 2330 12444 2339
rect 12338 2270 12340 2291
rect 12340 2270 12372 2291
rect 12410 2270 12442 2291
rect 12442 2270 12444 2291
rect 12338 2257 12372 2270
rect 12410 2257 12444 2270
rect 12338 2201 12340 2218
rect 12340 2201 12372 2218
rect 12410 2201 12442 2218
rect 12442 2201 12444 2218
rect 12338 2184 12372 2201
rect 12410 2184 12444 2201
rect 12338 2132 12340 2145
rect 12340 2132 12372 2145
rect 12410 2132 12442 2145
rect 12442 2132 12444 2145
rect 12338 2111 12372 2132
rect 12410 2111 12444 2132
rect 12338 2063 12340 2072
rect 12340 2063 12372 2072
rect 12410 2063 12442 2072
rect 12442 2063 12444 2072
rect 12338 2038 12372 2063
rect 12410 2038 12444 2063
rect 12338 1994 12340 1999
rect 12340 1994 12372 1999
rect 12410 1994 12442 1999
rect 12442 1994 12444 1999
rect 12338 1965 12372 1994
rect 12410 1965 12444 1994
rect 12338 1925 12340 1926
rect 12340 1925 12372 1926
rect 12410 1925 12442 1926
rect 12442 1925 12444 1926
rect 12338 1892 12372 1925
rect 12410 1892 12444 1925
rect 12338 1821 12372 1853
rect 12410 1821 12444 1853
rect 12338 1819 12340 1821
rect 12340 1819 12372 1821
rect 12410 1819 12442 1821
rect 12442 1819 12444 1821
rect 12338 1752 12372 1780
rect 12410 1752 12444 1780
rect 12338 1746 12340 1752
rect 12340 1746 12372 1752
rect 12410 1746 12442 1752
rect 12442 1746 12444 1752
rect 12338 1683 12372 1707
rect 12410 1683 12444 1707
rect 12338 1673 12340 1683
rect 12340 1673 12372 1683
rect 12410 1673 12442 1683
rect 12442 1673 12444 1683
rect 12338 1614 12372 1634
rect 12410 1614 12444 1634
rect 12338 1600 12340 1614
rect 12340 1600 12372 1614
rect 12410 1600 12442 1614
rect 12442 1600 12444 1614
rect 12338 1545 12372 1561
rect 12410 1545 12444 1561
rect 12338 1527 12340 1545
rect 12340 1527 12372 1545
rect 12410 1527 12442 1545
rect 12442 1527 12444 1545
rect 12338 1476 12372 1488
rect 12410 1476 12444 1488
rect 12338 1454 12340 1476
rect 12340 1454 12372 1476
rect 12410 1454 12442 1476
rect 12442 1454 12444 1476
rect 12338 1407 12372 1415
rect 12410 1407 12444 1415
rect 12338 1381 12340 1407
rect 12340 1381 12372 1407
rect 12410 1381 12442 1407
rect 12442 1381 12444 1407
rect 12338 1338 12372 1342
rect 12410 1338 12444 1342
rect 12338 1308 12340 1338
rect 12340 1308 12372 1338
rect 12410 1308 12442 1338
rect 12442 1308 12444 1338
rect 12338 1235 12340 1269
rect 12340 1235 12372 1269
rect 12410 1235 12442 1269
rect 12442 1235 12444 1269
rect 13240 3719 13242 11233
rect 13242 3719 13344 11233
rect 13344 3719 13346 11233
rect 13240 3684 13346 3719
rect 13240 3650 13242 3684
rect 13242 3650 13276 3684
rect 13276 3650 13310 3684
rect 13310 3650 13344 3684
rect 13344 3650 13346 3684
rect 13240 3615 13346 3650
rect 13240 3581 13242 3615
rect 13242 3581 13276 3615
rect 13276 3581 13310 3615
rect 13310 3581 13344 3615
rect 13344 3581 13346 3615
rect 13240 3546 13346 3581
rect 13240 3512 13242 3546
rect 13242 3512 13276 3546
rect 13276 3512 13310 3546
rect 13310 3512 13344 3546
rect 13344 3512 13346 3546
rect 13240 3477 13346 3512
rect 13240 3443 13242 3477
rect 13242 3443 13276 3477
rect 13276 3443 13310 3477
rect 13310 3443 13344 3477
rect 13344 3443 13346 3477
rect 13240 3408 13346 3443
rect 13240 3374 13242 3408
rect 13242 3374 13276 3408
rect 13276 3374 13310 3408
rect 13310 3374 13344 3408
rect 13344 3374 13346 3408
rect 13240 3339 13346 3374
rect 13240 3305 13242 3339
rect 13242 3305 13276 3339
rect 13276 3305 13310 3339
rect 13310 3305 13344 3339
rect 13344 3305 13346 3339
rect 13240 3279 13346 3305
rect 13240 3236 13242 3240
rect 13242 3236 13274 3240
rect 13312 3236 13344 3240
rect 13344 3236 13346 3240
rect 13240 3206 13274 3236
rect 13312 3206 13346 3236
rect 13240 3133 13274 3167
rect 13312 3133 13346 3167
rect 13240 3063 13274 3094
rect 13312 3063 13346 3094
rect 13240 3060 13242 3063
rect 13242 3060 13274 3063
rect 13312 3060 13344 3063
rect 13344 3060 13346 3063
rect 13240 2994 13274 3021
rect 13312 2994 13346 3021
rect 13240 2987 13242 2994
rect 13242 2987 13274 2994
rect 13312 2987 13344 2994
rect 13344 2987 13346 2994
rect 13240 2925 13274 2948
rect 13312 2925 13346 2948
rect 13240 2914 13242 2925
rect 13242 2914 13274 2925
rect 13312 2914 13344 2925
rect 13344 2914 13346 2925
rect 13240 2856 13274 2875
rect 13312 2856 13346 2875
rect 13240 2841 13242 2856
rect 13242 2841 13274 2856
rect 13312 2841 13344 2856
rect 13344 2841 13346 2856
rect 13240 2787 13274 2802
rect 13312 2787 13346 2802
rect 13240 2768 13242 2787
rect 13242 2768 13274 2787
rect 13312 2768 13344 2787
rect 13344 2768 13346 2787
rect 13240 2718 13274 2729
rect 13312 2718 13346 2729
rect 13240 2695 13242 2718
rect 13242 2695 13274 2718
rect 13312 2695 13344 2718
rect 13344 2695 13346 2718
rect 13240 2649 13274 2656
rect 13312 2649 13346 2656
rect 13240 2622 13242 2649
rect 13242 2622 13274 2649
rect 13312 2622 13344 2649
rect 13344 2622 13346 2649
rect 13240 2580 13274 2583
rect 13312 2580 13346 2583
rect 13240 2549 13242 2580
rect 13242 2549 13274 2580
rect 13312 2549 13344 2580
rect 13344 2549 13346 2580
rect 13240 2477 13242 2510
rect 13242 2477 13274 2510
rect 13312 2477 13344 2510
rect 13344 2477 13346 2510
rect 13240 2476 13274 2477
rect 13312 2476 13346 2477
rect 13240 2408 13242 2437
rect 13242 2408 13274 2437
rect 13312 2408 13344 2437
rect 13344 2408 13346 2437
rect 13240 2403 13274 2408
rect 13312 2403 13346 2408
rect 13240 2339 13242 2364
rect 13242 2339 13274 2364
rect 13312 2339 13344 2364
rect 13344 2339 13346 2364
rect 13240 2330 13274 2339
rect 13312 2330 13346 2339
rect 13240 2270 13242 2291
rect 13242 2270 13274 2291
rect 13312 2270 13344 2291
rect 13344 2270 13346 2291
rect 13240 2257 13274 2270
rect 13312 2257 13346 2270
rect 13240 2201 13242 2218
rect 13242 2201 13274 2218
rect 13312 2201 13344 2218
rect 13344 2201 13346 2218
rect 13240 2184 13274 2201
rect 13312 2184 13346 2201
rect 13240 2132 13242 2145
rect 13242 2132 13274 2145
rect 13312 2132 13344 2145
rect 13344 2132 13346 2145
rect 13240 2111 13274 2132
rect 13312 2111 13346 2132
rect 13240 2063 13242 2072
rect 13242 2063 13274 2072
rect 13312 2063 13344 2072
rect 13344 2063 13346 2072
rect 13240 2038 13274 2063
rect 13312 2038 13346 2063
rect 13240 1994 13242 1999
rect 13242 1994 13274 1999
rect 13312 1994 13344 1999
rect 13344 1994 13346 1999
rect 13240 1965 13274 1994
rect 13312 1965 13346 1994
rect 13240 1925 13242 1926
rect 13242 1925 13274 1926
rect 13312 1925 13344 1926
rect 13344 1925 13346 1926
rect 13240 1892 13274 1925
rect 13312 1892 13346 1925
rect 13240 1821 13274 1853
rect 13312 1821 13346 1853
rect 13240 1819 13242 1821
rect 13242 1819 13274 1821
rect 13312 1819 13344 1821
rect 13344 1819 13346 1821
rect 13240 1752 13274 1780
rect 13312 1752 13346 1780
rect 13240 1746 13242 1752
rect 13242 1746 13274 1752
rect 13312 1746 13344 1752
rect 13344 1746 13346 1752
rect 13240 1683 13274 1707
rect 13312 1683 13346 1707
rect 13240 1673 13242 1683
rect 13242 1673 13274 1683
rect 13312 1673 13344 1683
rect 13344 1673 13346 1683
rect 13240 1614 13274 1634
rect 13312 1614 13346 1634
rect 13240 1600 13242 1614
rect 13242 1600 13274 1614
rect 13312 1600 13344 1614
rect 13344 1600 13346 1614
rect 13240 1545 13274 1561
rect 13312 1545 13346 1561
rect 13240 1527 13242 1545
rect 13242 1527 13274 1545
rect 13312 1527 13344 1545
rect 13344 1527 13346 1545
rect 13240 1476 13274 1488
rect 13312 1476 13346 1488
rect 13240 1454 13242 1476
rect 13242 1454 13274 1476
rect 13312 1454 13344 1476
rect 13344 1454 13346 1476
rect 13240 1407 13274 1415
rect 13312 1407 13346 1415
rect 13240 1381 13242 1407
rect 13242 1381 13274 1407
rect 13312 1381 13344 1407
rect 13344 1381 13346 1407
rect 13240 1338 13274 1342
rect 13312 1338 13346 1342
rect 13240 1308 13242 1338
rect 13242 1308 13274 1338
rect 13312 1308 13344 1338
rect 13344 1308 13346 1338
rect 13240 1235 13242 1269
rect 13242 1235 13274 1269
rect 13312 1235 13344 1269
rect 13344 1235 13346 1269
rect 14142 3719 14144 11233
rect 14144 3719 14246 11233
rect 14246 3719 14248 11233
rect 14142 3684 14248 3719
rect 14142 3650 14144 3684
rect 14144 3650 14178 3684
rect 14178 3650 14212 3684
rect 14212 3650 14246 3684
rect 14246 3650 14248 3684
rect 14142 3615 14248 3650
rect 14142 3581 14144 3615
rect 14144 3581 14178 3615
rect 14178 3581 14212 3615
rect 14212 3581 14246 3615
rect 14246 3581 14248 3615
rect 14142 3546 14248 3581
rect 14142 3512 14144 3546
rect 14144 3512 14178 3546
rect 14178 3512 14212 3546
rect 14212 3512 14246 3546
rect 14246 3512 14248 3546
rect 14142 3477 14248 3512
rect 14142 3443 14144 3477
rect 14144 3443 14178 3477
rect 14178 3443 14212 3477
rect 14212 3443 14246 3477
rect 14246 3443 14248 3477
rect 14142 3408 14248 3443
rect 14142 3374 14144 3408
rect 14144 3374 14178 3408
rect 14178 3374 14212 3408
rect 14212 3374 14246 3408
rect 14246 3374 14248 3408
rect 14142 3339 14248 3374
rect 14142 3305 14144 3339
rect 14144 3305 14178 3339
rect 14178 3305 14212 3339
rect 14212 3305 14246 3339
rect 14246 3305 14248 3339
rect 14142 3279 14248 3305
rect 14142 3236 14144 3240
rect 14144 3236 14176 3240
rect 14214 3236 14246 3240
rect 14246 3236 14248 3240
rect 14142 3206 14176 3236
rect 14214 3206 14248 3236
rect 14142 3133 14176 3167
rect 14214 3133 14248 3167
rect 14142 3063 14176 3094
rect 14214 3063 14248 3094
rect 14142 3060 14144 3063
rect 14144 3060 14176 3063
rect 14214 3060 14246 3063
rect 14246 3060 14248 3063
rect 14142 2994 14176 3021
rect 14214 2994 14248 3021
rect 14142 2987 14144 2994
rect 14144 2987 14176 2994
rect 14214 2987 14246 2994
rect 14246 2987 14248 2994
rect 14142 2925 14176 2948
rect 14214 2925 14248 2948
rect 14142 2914 14144 2925
rect 14144 2914 14176 2925
rect 14214 2914 14246 2925
rect 14246 2914 14248 2925
rect 14142 2856 14176 2875
rect 14214 2856 14248 2875
rect 14142 2841 14144 2856
rect 14144 2841 14176 2856
rect 14214 2841 14246 2856
rect 14246 2841 14248 2856
rect 14142 2787 14176 2802
rect 14214 2787 14248 2802
rect 14142 2768 14144 2787
rect 14144 2768 14176 2787
rect 14214 2768 14246 2787
rect 14246 2768 14248 2787
rect 14142 2718 14176 2729
rect 14214 2718 14248 2729
rect 14142 2695 14144 2718
rect 14144 2695 14176 2718
rect 14214 2695 14246 2718
rect 14246 2695 14248 2718
rect 14142 2649 14176 2656
rect 14214 2649 14248 2656
rect 14142 2622 14144 2649
rect 14144 2622 14176 2649
rect 14214 2622 14246 2649
rect 14246 2622 14248 2649
rect 14142 2580 14176 2583
rect 14214 2580 14248 2583
rect 14142 2549 14144 2580
rect 14144 2549 14176 2580
rect 14214 2549 14246 2580
rect 14246 2549 14248 2580
rect 14142 2477 14144 2510
rect 14144 2477 14176 2510
rect 14214 2477 14246 2510
rect 14246 2477 14248 2510
rect 14142 2476 14176 2477
rect 14214 2476 14248 2477
rect 14142 2408 14144 2437
rect 14144 2408 14176 2437
rect 14214 2408 14246 2437
rect 14246 2408 14248 2437
rect 14142 2403 14176 2408
rect 14214 2403 14248 2408
rect 14142 2339 14144 2364
rect 14144 2339 14176 2364
rect 14214 2339 14246 2364
rect 14246 2339 14248 2364
rect 14142 2330 14176 2339
rect 14214 2330 14248 2339
rect 14142 2270 14144 2291
rect 14144 2270 14176 2291
rect 14214 2270 14246 2291
rect 14246 2270 14248 2291
rect 14142 2257 14176 2270
rect 14214 2257 14248 2270
rect 14142 2201 14144 2218
rect 14144 2201 14176 2218
rect 14214 2201 14246 2218
rect 14246 2201 14248 2218
rect 14142 2184 14176 2201
rect 14214 2184 14248 2201
rect 14142 2132 14144 2145
rect 14144 2132 14176 2145
rect 14214 2132 14246 2145
rect 14246 2132 14248 2145
rect 14142 2111 14176 2132
rect 14214 2111 14248 2132
rect 14142 2063 14144 2072
rect 14144 2063 14176 2072
rect 14214 2063 14246 2072
rect 14246 2063 14248 2072
rect 14142 2038 14176 2063
rect 14214 2038 14248 2063
rect 14142 1994 14144 1999
rect 14144 1994 14176 1999
rect 14214 1994 14246 1999
rect 14246 1994 14248 1999
rect 14142 1965 14176 1994
rect 14214 1965 14248 1994
rect 14142 1925 14144 1926
rect 14144 1925 14176 1926
rect 14214 1925 14246 1926
rect 14246 1925 14248 1926
rect 14142 1892 14176 1925
rect 14214 1892 14248 1925
rect 14142 1821 14176 1853
rect 14214 1821 14248 1853
rect 14142 1819 14144 1821
rect 14144 1819 14176 1821
rect 14214 1819 14246 1821
rect 14246 1819 14248 1821
rect 14142 1752 14176 1780
rect 14214 1752 14248 1780
rect 14142 1746 14144 1752
rect 14144 1746 14176 1752
rect 14214 1746 14246 1752
rect 14246 1746 14248 1752
rect 14142 1683 14176 1707
rect 14214 1683 14248 1707
rect 14142 1673 14144 1683
rect 14144 1673 14176 1683
rect 14214 1673 14246 1683
rect 14246 1673 14248 1683
rect 14142 1614 14176 1634
rect 14214 1614 14248 1634
rect 14142 1600 14144 1614
rect 14144 1600 14176 1614
rect 14214 1600 14246 1614
rect 14246 1600 14248 1614
rect 14142 1545 14176 1561
rect 14214 1545 14248 1561
rect 14142 1527 14144 1545
rect 14144 1527 14176 1545
rect 14214 1527 14246 1545
rect 14246 1527 14248 1545
rect 14142 1476 14176 1488
rect 14214 1476 14248 1488
rect 14142 1454 14144 1476
rect 14144 1454 14176 1476
rect 14214 1454 14246 1476
rect 14246 1454 14248 1476
rect 14142 1407 14176 1415
rect 14214 1407 14248 1415
rect 14142 1381 14144 1407
rect 14144 1381 14176 1407
rect 14214 1381 14246 1407
rect 14246 1381 14248 1407
rect 14142 1338 14176 1342
rect 14214 1338 14248 1342
rect 14142 1308 14144 1338
rect 14144 1308 14176 1338
rect 14214 1308 14246 1338
rect 14246 1308 14248 1338
rect 14142 1235 14144 1269
rect 14144 1235 14176 1269
rect 14214 1235 14246 1269
rect 14246 1235 14248 1269
rect -3644 1008 -3642 1020
rect -3642 1008 -3610 1020
rect -3572 1008 -3540 1020
rect -3540 1008 -3538 1020
rect -3644 986 -3610 1008
rect -3572 986 -3538 1008
rect -2352 1008 -2350 1042
rect -2350 1008 -2318 1042
rect -2280 1008 -2248 1042
rect -2248 1008 -2246 1042
rect -1840 1008 -1838 1042
rect -1838 1008 -1806 1042
rect -1768 1008 -1736 1042
rect -1736 1008 -1734 1042
rect -548 1008 -546 1042
rect -546 1008 -514 1042
rect -476 1008 -444 1042
rect -444 1008 -442 1042
rect -36 1008 -34 1042
rect -34 1008 -2 1042
rect 36 1008 68 1042
rect 68 1008 70 1042
rect 1256 1008 1258 1042
rect 1258 1008 1290 1042
rect 1328 1008 1360 1042
rect 1360 1008 1362 1042
rect 1768 1008 1770 1042
rect 1770 1008 1802 1042
rect 1840 1008 1872 1042
rect 1872 1008 1874 1042
rect 3060 1008 3062 1042
rect 3062 1008 3094 1042
rect 3132 1008 3164 1042
rect 3164 1008 3166 1042
rect 3572 1008 3574 1042
rect 3574 1008 3606 1042
rect 3644 1008 3676 1042
rect 3676 1008 3678 1042
rect 4864 1008 4866 1042
rect 4866 1008 4898 1042
rect 4936 1008 4968 1042
rect 4968 1008 4970 1042
rect 5376 1008 5378 1042
rect 5378 1008 5410 1042
rect 5448 1008 5480 1042
rect 5480 1008 5482 1042
rect 6668 1008 6670 1042
rect 6670 1008 6702 1042
rect 6740 1008 6772 1042
rect 6772 1008 6774 1042
rect 7180 1008 7182 1042
rect 7182 1008 7214 1042
rect 7252 1008 7284 1042
rect 7284 1008 7286 1042
rect 8472 1008 8474 1042
rect 8474 1008 8506 1042
rect 8544 1008 8576 1042
rect 8576 1008 8578 1042
rect 8984 1008 8986 1042
rect 8986 1008 9018 1042
rect 9056 1008 9088 1042
rect 9088 1008 9090 1042
rect 10276 1008 10278 1042
rect 10278 1008 10310 1042
rect 10348 1008 10380 1042
rect 10380 1008 10382 1042
rect 10788 1008 10790 1042
rect 10790 1008 10822 1042
rect 10860 1008 10892 1042
rect 10892 1008 10894 1042
rect 12080 1008 12082 1042
rect 12082 1008 12114 1042
rect 12152 1008 12184 1042
rect 12184 1008 12186 1042
rect 12592 1008 12594 1042
rect 12594 1008 12626 1042
rect 12664 1008 12696 1042
rect 12696 1008 12698 1042
rect 13884 1008 13886 1020
rect 13886 1008 13918 1020
rect 13956 1008 13988 1020
rect 13988 1008 13990 1020
rect 13884 986 13918 1008
rect 13956 986 13990 1008
rect -4313 606 -4299 608
rect -4299 606 -4279 608
rect -4313 574 -4279 606
rect 14603 574 14637 608
rect 15132 11611 15238 11861
rect 15132 11543 15166 11562
rect 15204 11543 15238 11562
rect 15132 11528 15134 11543
rect 15134 11528 15166 11543
rect 15204 11528 15236 11543
rect 15236 11528 15238 11543
rect 15132 11464 15238 11483
rect 15132 5185 15238 11464
rect 15132 5112 15166 5146
rect 15204 5112 15238 5146
rect 15132 5039 15166 5073
rect 15204 5039 15238 5073
rect 15132 4966 15166 5000
rect 15204 4966 15238 5000
rect 15132 4893 15166 4927
rect 15204 4893 15238 4927
rect 15132 4820 15166 4854
rect 15204 4820 15238 4854
rect 15132 4747 15166 4781
rect 15204 4747 15238 4781
rect 15132 4674 15166 4708
rect 15204 4674 15238 4708
rect 15132 4601 15166 4635
rect 15204 4601 15238 4635
rect 15132 4528 15166 4562
rect 15204 4528 15238 4562
rect 15132 4455 15166 4489
rect 15204 4455 15238 4489
rect 15132 4382 15166 4416
rect 15204 4382 15238 4416
rect 15132 4309 15166 4343
rect 15204 4309 15238 4343
rect 15132 4236 15166 4270
rect 15204 4236 15238 4270
rect 15132 4163 15166 4197
rect 15204 4163 15238 4197
rect 15132 4090 15166 4124
rect 15204 4090 15238 4124
rect 15132 4017 15166 4051
rect 15204 4017 15238 4051
rect 15132 3944 15166 3978
rect 15204 3944 15238 3978
rect 15132 3871 15166 3905
rect 15204 3871 15238 3905
rect 15132 3798 15166 3832
rect 15204 3798 15238 3832
rect 15132 3725 15166 3759
rect 15204 3725 15238 3759
rect 15132 3652 15166 3686
rect 15204 3652 15238 3686
rect 15132 3579 15166 3613
rect 15204 3579 15238 3613
rect 15132 3506 15166 3540
rect 15204 3506 15238 3540
rect 15132 3433 15166 3467
rect 15204 3433 15238 3467
rect 15132 3360 15166 3394
rect 15204 3360 15238 3394
rect 15132 3287 15166 3321
rect 15204 3287 15238 3321
rect 15132 3214 15166 3248
rect 15204 3214 15238 3248
rect 15132 3141 15166 3175
rect 15204 3141 15238 3175
rect 15132 3068 15166 3102
rect 15204 3068 15238 3102
rect 15132 2995 15166 3029
rect 15204 2995 15238 3029
rect 15132 2922 15166 2956
rect 15204 2922 15238 2956
rect 15132 2849 15166 2883
rect 15204 2849 15238 2883
rect 15132 2776 15166 2810
rect 15204 2776 15238 2810
rect 15132 2703 15166 2737
rect 15204 2703 15238 2737
rect 15132 2630 15166 2664
rect 15204 2630 15238 2664
rect 15132 2557 15166 2591
rect 15204 2557 15238 2591
rect 15132 2484 15166 2518
rect 15204 2484 15238 2518
rect 15132 2411 15166 2445
rect 15204 2411 15238 2445
rect 15132 2338 15166 2372
rect 15204 2338 15238 2372
rect 15132 2265 15166 2299
rect 15204 2265 15238 2299
rect 15132 2192 15166 2226
rect 15204 2192 15238 2226
rect 15132 2119 15166 2153
rect 15204 2119 15238 2153
rect 15132 2046 15166 2080
rect 15204 2046 15238 2080
rect 15132 1973 15166 2007
rect 15204 1973 15238 2007
rect 15132 1900 15166 1934
rect 15204 1900 15238 1934
rect 15132 1827 15166 1861
rect 15204 1827 15238 1861
rect 15132 1754 15166 1788
rect 15204 1754 15238 1788
rect 15132 1681 15166 1715
rect 15204 1681 15238 1715
rect 15132 1608 15166 1642
rect 15204 1608 15238 1642
rect 15132 1535 15166 1569
rect 15204 1535 15238 1569
rect 15132 1462 15166 1496
rect 15204 1462 15238 1496
rect 15132 1389 15166 1423
rect 15204 1389 15238 1423
rect 15132 1316 15166 1350
rect 15204 1316 15238 1350
rect 15132 1243 15166 1277
rect 15204 1243 15238 1277
rect 15132 1170 15166 1204
rect 15204 1170 15238 1204
rect 15132 1097 15166 1131
rect 15204 1097 15238 1131
rect 15132 1024 15166 1058
rect 15204 1024 15238 1058
rect 15132 951 15166 985
rect 15204 951 15238 985
rect 15132 890 15166 912
rect 15204 890 15238 912
rect 15132 878 15166 890
rect 15204 878 15238 890
rect 15132 821 15134 839
rect 15134 821 15166 839
rect 15204 821 15236 839
rect 15236 821 15238 839
rect 15132 805 15166 821
rect 15204 805 15238 821
rect 15132 752 15134 766
rect 15134 752 15166 766
rect 15204 752 15236 766
rect 15236 752 15238 766
rect 15132 732 15166 752
rect 15204 732 15238 752
rect 15132 683 15134 693
rect 15134 683 15166 693
rect 15204 683 15236 693
rect 15236 683 15238 693
rect 15132 659 15166 683
rect 15204 659 15238 683
rect 15132 614 15134 620
rect 15134 614 15166 620
rect 15204 614 15236 620
rect 15236 614 15238 620
rect 15132 586 15166 614
rect 15204 586 15238 614
rect 15132 545 15134 547
rect 15134 545 15166 547
rect 15204 545 15236 547
rect 15236 545 15238 547
rect 15132 513 15166 545
rect 15204 513 15238 545
rect -4888 440 -4886 441
rect -4886 440 -4854 441
rect -4816 440 -4784 441
rect -4784 440 -4782 441
rect -4888 372 -4854 401
rect -4816 372 -4782 401
rect -4888 367 -4886 372
rect -4886 367 -4854 372
rect -4816 367 -4784 372
rect -4784 367 -4782 372
rect 15132 441 15166 474
rect 15204 441 15238 474
rect 15132 440 15134 441
rect 15134 440 15166 441
rect 15204 440 15236 441
rect 15236 440 15238 441
rect 15132 372 15166 401
rect 15204 372 15238 401
rect 15132 367 15134 372
rect 15134 367 15166 372
rect 15204 367 15236 372
rect 15236 367 15238 372
<< metal1 >>
tri -4965 12850 -4835 12980 se
rect -4835 12850 15185 12980
tri 15185 12850 15315 12980 sw
rect -4965 12757 15315 12850
rect -4965 11931 -4888 12757
rect -4782 12480 15132 12757
rect -4782 11931 -4770 12480
tri -4770 12270 -4560 12480 nw
tri 14910 12270 15120 12480 ne
tri -4165 11931 -3916 12180 se
rect -3916 11931 14266 12180
tri 14266 11931 14515 12180 sw
rect 15120 11931 15132 12480
rect 15238 11931 15315 12757
rect -4965 11861 -4770 11931
tri -4235 11861 -4165 11931 se
rect -4165 11861 14515 11931
tri 14515 11861 14585 11931 sw
rect 15120 11861 15315 11931
rect -4965 11611 -4888 11861
rect -4782 11611 -4770 11861
rect -4965 11562 -4770 11611
rect -4965 11528 -4888 11562
rect -4854 11528 -4816 11562
rect -4782 11528 -4770 11562
rect -4965 11483 -4770 11528
rect -4965 5185 -4888 11483
rect -4782 5185 -4770 11483
rect -4965 5146 -4770 5185
rect -4965 5112 -4888 5146
rect -4854 5112 -4816 5146
rect -4782 5112 -4770 5146
rect -4965 5073 -4770 5112
rect -4965 5039 -4888 5073
rect -4854 5039 -4816 5073
rect -4782 5039 -4770 5073
rect -4965 5000 -4770 5039
rect -4965 4966 -4888 5000
rect -4854 4966 -4816 5000
rect -4782 4966 -4770 5000
rect -4965 4927 -4770 4966
rect -4965 4893 -4888 4927
rect -4854 4893 -4816 4927
rect -4782 4893 -4770 4927
rect -4965 4854 -4770 4893
rect -4965 4820 -4888 4854
rect -4854 4820 -4816 4854
rect -4782 4820 -4770 4854
rect -4965 4781 -4770 4820
rect -4965 4747 -4888 4781
rect -4854 4747 -4816 4781
rect -4782 4747 -4770 4781
rect -4965 4708 -4770 4747
rect -4965 4674 -4888 4708
rect -4854 4674 -4816 4708
rect -4782 4674 -4770 4708
rect -4965 4635 -4770 4674
rect -4965 4601 -4888 4635
rect -4854 4601 -4816 4635
rect -4782 4601 -4770 4635
rect -4965 4562 -4770 4601
rect -4965 4528 -4888 4562
rect -4854 4528 -4816 4562
rect -4782 4528 -4770 4562
rect -4965 4489 -4770 4528
rect -4965 4455 -4888 4489
rect -4854 4455 -4816 4489
rect -4782 4455 -4770 4489
rect -4965 4416 -4770 4455
rect -4965 4382 -4888 4416
rect -4854 4382 -4816 4416
rect -4782 4382 -4770 4416
rect -4965 4343 -4770 4382
rect -4965 4309 -4888 4343
rect -4854 4309 -4816 4343
rect -4782 4309 -4770 4343
rect -4965 4270 -4770 4309
rect -4965 4236 -4888 4270
rect -4854 4236 -4816 4270
rect -4782 4236 -4770 4270
rect -4965 4197 -4770 4236
rect -4965 4163 -4888 4197
rect -4854 4163 -4816 4197
rect -4782 4163 -4770 4197
rect -4965 4124 -4770 4163
rect -4965 4090 -4888 4124
rect -4854 4090 -4816 4124
rect -4782 4090 -4770 4124
rect -4965 4051 -4770 4090
rect -4965 4017 -4888 4051
rect -4854 4017 -4816 4051
rect -4782 4017 -4770 4051
rect -4965 3978 -4770 4017
rect -4965 3944 -4888 3978
rect -4854 3944 -4816 3978
rect -4782 3944 -4770 3978
rect -4965 3905 -4770 3944
rect -4965 3871 -4888 3905
rect -4854 3871 -4816 3905
rect -4782 3871 -4770 3905
rect -4965 3832 -4770 3871
rect -4965 3798 -4888 3832
rect -4854 3798 -4816 3832
rect -4782 3798 -4770 3832
rect -4965 3759 -4770 3798
rect -4965 3725 -4888 3759
rect -4854 3725 -4816 3759
rect -4782 3725 -4770 3759
rect -4965 3686 -4770 3725
rect -4965 3652 -4888 3686
rect -4854 3652 -4816 3686
rect -4782 3652 -4770 3686
rect -4965 3613 -4770 3652
rect -4965 3579 -4888 3613
rect -4854 3579 -4816 3613
rect -4782 3579 -4770 3613
rect -4965 3540 -4770 3579
rect -4965 3506 -4888 3540
rect -4854 3506 -4816 3540
rect -4782 3506 -4770 3540
rect -4965 3467 -4770 3506
rect -4965 3433 -4888 3467
rect -4854 3433 -4816 3467
rect -4782 3433 -4770 3467
rect -4965 3394 -4770 3433
rect -4965 3360 -4888 3394
rect -4854 3360 -4816 3394
rect -4782 3360 -4770 3394
rect -4965 3321 -4770 3360
rect -4965 3287 -4888 3321
rect -4854 3287 -4816 3321
rect -4782 3287 -4770 3321
rect -4965 3248 -4770 3287
rect -4965 3214 -4888 3248
rect -4854 3214 -4816 3248
rect -4782 3214 -4770 3248
rect -4965 3175 -4770 3214
rect -4965 3141 -4888 3175
rect -4854 3141 -4816 3175
rect -4782 3141 -4770 3175
rect -4965 3102 -4770 3141
rect -4965 3068 -4888 3102
rect -4854 3068 -4816 3102
rect -4782 3068 -4770 3102
rect -4965 3029 -4770 3068
rect -4965 2995 -4888 3029
rect -4854 2995 -4816 3029
rect -4782 2995 -4770 3029
rect -4965 2956 -4770 2995
rect -4965 2922 -4888 2956
rect -4854 2922 -4816 2956
rect -4782 2922 -4770 2956
rect -4965 2883 -4770 2922
rect -4965 2849 -4888 2883
rect -4854 2849 -4816 2883
rect -4782 2849 -4770 2883
rect -4965 2810 -4770 2849
rect -4965 2776 -4888 2810
rect -4854 2776 -4816 2810
rect -4782 2776 -4770 2810
rect -4965 2737 -4770 2776
rect -4965 2703 -4888 2737
rect -4854 2703 -4816 2737
rect -4782 2703 -4770 2737
rect -4965 2664 -4770 2703
rect -4965 2630 -4888 2664
rect -4854 2630 -4816 2664
rect -4782 2630 -4770 2664
rect -4965 2591 -4770 2630
rect -4965 2557 -4888 2591
rect -4854 2557 -4816 2591
rect -4782 2557 -4770 2591
rect -4965 2518 -4770 2557
rect -4965 2484 -4888 2518
rect -4854 2484 -4816 2518
rect -4782 2484 -4770 2518
rect -4965 2445 -4770 2484
rect -4965 2411 -4888 2445
rect -4854 2411 -4816 2445
rect -4782 2411 -4770 2445
rect -4965 2372 -4770 2411
rect -4965 2338 -4888 2372
rect -4854 2338 -4816 2372
rect -4782 2338 -4770 2372
rect -4965 2299 -4770 2338
rect -4965 2265 -4888 2299
rect -4854 2265 -4816 2299
rect -4782 2265 -4770 2299
rect -4965 2226 -4770 2265
rect -4965 2192 -4888 2226
rect -4854 2192 -4816 2226
rect -4782 2192 -4770 2226
rect -4965 2153 -4770 2192
rect -4965 2119 -4888 2153
rect -4854 2119 -4816 2153
rect -4782 2119 -4770 2153
rect -4965 2080 -4770 2119
rect -4965 2046 -4888 2080
rect -4854 2046 -4816 2080
rect -4782 2046 -4770 2080
rect -4965 2007 -4770 2046
rect -4965 1973 -4888 2007
rect -4854 1973 -4816 2007
rect -4782 1973 -4770 2007
rect -4965 1934 -4770 1973
rect -4965 1900 -4888 1934
rect -4854 1900 -4816 1934
rect -4782 1900 -4770 1934
rect -4965 1861 -4770 1900
rect -4965 1827 -4888 1861
rect -4854 1827 -4816 1861
rect -4782 1827 -4770 1861
rect -4965 1788 -4770 1827
rect -4965 1754 -4888 1788
rect -4854 1754 -4816 1788
rect -4782 1754 -4770 1788
rect -4965 1715 -4770 1754
rect -4965 1681 -4888 1715
rect -4854 1681 -4816 1715
rect -4782 1681 -4770 1715
rect -4965 1642 -4770 1681
rect -4965 1608 -4888 1642
rect -4854 1608 -4816 1642
rect -4782 1608 -4770 1642
rect -4965 1569 -4770 1608
rect -4965 1535 -4888 1569
rect -4854 1535 -4816 1569
rect -4782 1535 -4770 1569
rect -4965 1496 -4770 1535
rect -4965 1462 -4888 1496
rect -4854 1462 -4816 1496
rect -4782 1462 -4770 1496
rect -4965 1423 -4770 1462
rect -4965 1389 -4888 1423
rect -4854 1389 -4816 1423
rect -4782 1389 -4770 1423
rect -4965 1350 -4770 1389
rect -4965 1316 -4888 1350
rect -4854 1316 -4816 1350
rect -4782 1316 -4770 1350
rect -4965 1277 -4770 1316
rect -4965 1243 -4888 1277
rect -4854 1243 -4816 1277
rect -4782 1243 -4770 1277
rect -4965 1204 -4770 1243
rect -4965 1170 -4888 1204
rect -4854 1170 -4816 1204
rect -4782 1170 -4770 1204
rect -4965 1131 -4770 1170
rect -4965 1097 -4888 1131
rect -4854 1097 -4816 1131
rect -4782 1097 -4770 1131
rect -4965 1058 -4770 1097
rect -4965 1024 -4888 1058
rect -4854 1024 -4816 1058
rect -4782 1024 -4770 1058
rect -4965 985 -4770 1024
rect -4965 951 -4888 985
rect -4854 951 -4816 985
rect -4782 951 -4770 985
rect -4965 912 -4770 951
rect -4965 878 -4888 912
rect -4854 878 -4816 912
rect -4782 878 -4770 912
rect -4965 839 -4770 878
rect -4965 805 -4888 839
rect -4854 805 -4816 839
rect -4782 805 -4770 839
rect -4965 766 -4770 805
rect -4965 732 -4888 766
rect -4854 732 -4816 766
rect -4782 732 -4770 766
rect -4965 693 -4770 732
rect -4965 659 -4888 693
rect -4854 659 -4816 693
rect -4782 659 -4770 693
rect -4965 620 -4770 659
rect -4965 586 -4888 620
rect -4854 586 -4816 620
rect -4782 586 -4770 620
tri -4416 11680 -4235 11861 se
rect -4235 11680 14585 11861
tri 14585 11680 14766 11861 sw
rect -4416 11611 -4065 11680
tri -4065 11611 -3996 11680 nw
tri 13606 11611 13675 11680 ne
rect 13675 11611 14766 11680
rect -4416 11562 -4114 11611
tri -4114 11562 -4065 11611 nw
tri 13675 11562 13724 11611 ne
rect 13724 11562 14766 11611
rect -4416 11528 -4148 11562
tri -4148 11528 -4114 11562 nw
tri 13724 11528 13758 11562 ne
rect 13758 11528 14766 11562
rect -4416 11483 -4193 11528
tri -4193 11483 -4148 11528 nw
tri 13758 11483 13803 11528 ne
rect 13803 11483 14766 11528
rect -4416 693 -4286 11483
tri -4286 11390 -4193 11483 nw
tri 13803 11390 13896 11483 ne
tri -4145 11333 -4098 11380 se
rect -4098 11333 -3592 11380
tri -3592 11333 -3545 11380 sw
rect -4145 11233 -3545 11333
rect -4145 3279 -3898 11233
rect -3792 3279 -3545 11233
rect -4145 3240 -3545 3279
rect -4145 3206 -3898 3240
rect -3864 3206 -3826 3240
rect -3792 3206 -3545 3240
rect -4145 3167 -3545 3206
rect -4145 3133 -3898 3167
rect -3864 3133 -3826 3167
rect -3792 3133 -3545 3167
rect -4145 3094 -3545 3133
rect -4145 3060 -3898 3094
rect -3864 3060 -3826 3094
rect -3792 3060 -3545 3094
rect -4145 3021 -3545 3060
rect -4145 2987 -3898 3021
rect -3864 2987 -3826 3021
rect -3792 2987 -3545 3021
rect -4145 2948 -3545 2987
rect -4145 2914 -3898 2948
rect -3864 2914 -3826 2948
rect -3792 2914 -3545 2948
rect -4145 2875 -3545 2914
rect -4145 2841 -3898 2875
rect -3864 2841 -3826 2875
rect -3792 2841 -3545 2875
rect -4145 2802 -3545 2841
rect -4145 2768 -3898 2802
rect -3864 2768 -3826 2802
rect -3792 2768 -3545 2802
rect -4145 2729 -3545 2768
rect -4145 2695 -3898 2729
rect -3864 2695 -3826 2729
rect -3792 2695 -3545 2729
rect -4145 2656 -3545 2695
rect -4145 2622 -3898 2656
rect -3864 2622 -3826 2656
rect -3792 2622 -3545 2656
rect -4145 2583 -3545 2622
rect -4145 2549 -3898 2583
rect -3864 2549 -3826 2583
rect -3792 2549 -3545 2583
rect -4145 2510 -3545 2549
rect -4145 2476 -3898 2510
rect -3864 2476 -3826 2510
rect -3792 2476 -3545 2510
rect -4145 2437 -3545 2476
rect -4145 2403 -3898 2437
rect -3864 2403 -3826 2437
rect -3792 2403 -3545 2437
rect -4145 2364 -3545 2403
rect -4145 2330 -3898 2364
rect -3864 2330 -3826 2364
rect -3792 2330 -3545 2364
rect -4145 2291 -3545 2330
rect -4145 2257 -3898 2291
rect -3864 2257 -3826 2291
rect -3792 2257 -3545 2291
rect -4145 2218 -3545 2257
rect -4145 2184 -3898 2218
rect -3864 2184 -3826 2218
rect -3792 2184 -3545 2218
rect -4145 2145 -3545 2184
rect -4145 2111 -3898 2145
rect -3864 2111 -3826 2145
rect -3792 2111 -3545 2145
rect -4145 2072 -3545 2111
rect -4145 2038 -3898 2072
rect -3864 2038 -3826 2072
rect -3792 2038 -3545 2072
rect -4145 1999 -3545 2038
rect -4145 1965 -3898 1999
rect -3864 1965 -3826 1999
rect -3792 1965 -3545 1999
rect -4145 1926 -3545 1965
rect -4145 1892 -3898 1926
rect -3864 1892 -3826 1926
rect -3792 1892 -3545 1926
rect -4145 1853 -3545 1892
rect -4145 1819 -3898 1853
rect -3864 1819 -3826 1853
rect -3792 1819 -3545 1853
rect -4145 1780 -3545 1819
rect -4145 1746 -3898 1780
rect -3864 1746 -3826 1780
rect -3792 1746 -3545 1780
rect -4145 1707 -3545 1746
rect -4145 1673 -3898 1707
rect -3864 1673 -3826 1707
rect -3792 1673 -3545 1707
rect -4145 1634 -3545 1673
rect -4145 1600 -3898 1634
rect -3864 1600 -3826 1634
rect -3792 1600 -3545 1634
rect -4145 1561 -3545 1600
rect -4145 1527 -3898 1561
rect -3864 1527 -3826 1561
rect -3792 1527 -3545 1561
rect -4145 1488 -3545 1527
rect -4145 1454 -3898 1488
rect -3864 1454 -3826 1488
rect -3792 1454 -3545 1488
rect -4145 1415 -3545 1454
rect -4145 1381 -3898 1415
rect -3864 1381 -3826 1415
rect -3792 1381 -3545 1415
rect -4145 1342 -3545 1381
rect -4145 1308 -3898 1342
rect -3864 1308 -3826 1342
rect -3792 1308 -3545 1342
rect -4145 1269 -3545 1308
rect -4145 1235 -3898 1269
rect -3864 1235 -3826 1269
rect -3792 1235 -3545 1269
rect -4145 1135 -3545 1235
tri -4145 1131 -4141 1135 ne
rect -4141 1131 -3549 1135
tri -3549 1131 -3545 1135 nw
tri -3243 11333 -3196 11380 se
rect -3196 11333 -2690 11380
tri -2690 11333 -2643 11380 sw
rect -3243 11233 -2643 11333
rect -3243 3279 -2996 11233
rect -2890 3279 -2643 11233
rect -3243 3240 -2643 3279
rect -3243 3206 -2996 3240
rect -2962 3206 -2924 3240
rect -2890 3206 -2643 3240
rect -3243 3167 -2643 3206
rect -3243 3133 -2996 3167
rect -2962 3133 -2924 3167
rect -2890 3133 -2643 3167
rect -3243 3094 -2643 3133
rect -3243 3060 -2996 3094
rect -2962 3060 -2924 3094
rect -2890 3060 -2643 3094
rect -3243 3021 -2643 3060
rect -3243 2987 -2996 3021
rect -2962 2987 -2924 3021
rect -2890 2987 -2643 3021
rect -3243 2948 -2643 2987
rect -3243 2914 -2996 2948
rect -2962 2914 -2924 2948
rect -2890 2914 -2643 2948
rect -3243 2875 -2643 2914
rect -3243 2841 -2996 2875
rect -2962 2841 -2924 2875
rect -2890 2841 -2643 2875
rect -3243 2802 -2643 2841
rect -3243 2768 -2996 2802
rect -2962 2768 -2924 2802
rect -2890 2768 -2643 2802
rect -3243 2729 -2643 2768
rect -3243 2695 -2996 2729
rect -2962 2695 -2924 2729
rect -2890 2695 -2643 2729
rect -3243 2656 -2643 2695
rect -3243 2622 -2996 2656
rect -2962 2622 -2924 2656
rect -2890 2622 -2643 2656
rect -3243 2583 -2643 2622
rect -3243 2549 -2996 2583
rect -2962 2549 -2924 2583
rect -2890 2549 -2643 2583
rect -3243 2510 -2643 2549
rect -3243 2476 -2996 2510
rect -2962 2476 -2924 2510
rect -2890 2476 -2643 2510
rect -3243 2437 -2643 2476
rect -3243 2403 -2996 2437
rect -2962 2403 -2924 2437
rect -2890 2403 -2643 2437
rect -3243 2364 -2643 2403
rect -3243 2330 -2996 2364
rect -2962 2330 -2924 2364
rect -2890 2330 -2643 2364
rect -3243 2291 -2643 2330
rect -3243 2257 -2996 2291
rect -2962 2257 -2924 2291
rect -2890 2257 -2643 2291
rect -3243 2218 -2643 2257
rect -3243 2184 -2996 2218
rect -2962 2184 -2924 2218
rect -2890 2184 -2643 2218
rect -3243 2145 -2643 2184
rect -3243 2111 -2996 2145
rect -2962 2111 -2924 2145
rect -2890 2111 -2643 2145
rect -3243 2072 -2643 2111
rect -3243 2038 -2996 2072
rect -2962 2038 -2924 2072
rect -2890 2038 -2643 2072
rect -3243 1999 -2643 2038
rect -3243 1965 -2996 1999
rect -2962 1965 -2924 1999
rect -2890 1965 -2643 1999
rect -3243 1926 -2643 1965
rect -3243 1892 -2996 1926
rect -2962 1892 -2924 1926
rect -2890 1892 -2643 1926
rect -3243 1853 -2643 1892
rect -3243 1819 -2996 1853
rect -2962 1819 -2924 1853
rect -2890 1819 -2643 1853
rect -3243 1780 -2643 1819
rect -3243 1746 -2996 1780
rect -2962 1746 -2924 1780
rect -2890 1746 -2643 1780
rect -3243 1707 -2643 1746
rect -3243 1673 -2996 1707
rect -2962 1673 -2924 1707
rect -2890 1673 -2643 1707
rect -3243 1634 -2643 1673
rect -3243 1600 -2996 1634
rect -2962 1600 -2924 1634
rect -2890 1600 -2643 1634
rect -3243 1561 -2643 1600
rect -3243 1527 -2996 1561
rect -2962 1527 -2924 1561
rect -2890 1527 -2643 1561
rect -3243 1488 -2643 1527
rect -3243 1454 -2996 1488
rect -2962 1454 -2924 1488
rect -2890 1454 -2643 1488
rect -3243 1415 -2643 1454
rect -3243 1381 -2996 1415
rect -2962 1381 -2924 1415
rect -2890 1381 -2643 1415
rect -3243 1342 -2643 1381
rect -3243 1308 -2996 1342
rect -2962 1308 -2924 1342
rect -2890 1308 -2643 1342
rect -3243 1269 -2643 1308
rect -3243 1235 -2996 1269
rect -2962 1235 -2924 1269
rect -2890 1235 -2643 1269
rect -3243 1135 -2643 1235
tri -3243 1131 -3239 1135 ne
rect -3239 1131 -2647 1135
tri -2647 1131 -2643 1135 nw
tri -2341 11333 -2294 11380 se
rect -2294 11333 -1788 11380
tri -1788 11333 -1741 11380 sw
rect -2341 11233 -1741 11333
rect -2341 3279 -2094 11233
rect -1988 3279 -1741 11233
rect -2341 3240 -1741 3279
rect -2341 3206 -2094 3240
rect -2060 3206 -2022 3240
rect -1988 3206 -1741 3240
rect -2341 3167 -1741 3206
rect -2341 3133 -2094 3167
rect -2060 3133 -2022 3167
rect -1988 3133 -1741 3167
rect -2341 3094 -1741 3133
rect -2341 3060 -2094 3094
rect -2060 3060 -2022 3094
rect -1988 3060 -1741 3094
rect -2341 3021 -1741 3060
rect -2341 2987 -2094 3021
rect -2060 2987 -2022 3021
rect -1988 2987 -1741 3021
rect -2341 2948 -1741 2987
rect -2341 2914 -2094 2948
rect -2060 2914 -2022 2948
rect -1988 2914 -1741 2948
rect -2341 2875 -1741 2914
rect -2341 2841 -2094 2875
rect -2060 2841 -2022 2875
rect -1988 2841 -1741 2875
rect -2341 2802 -1741 2841
rect -2341 2768 -2094 2802
rect -2060 2768 -2022 2802
rect -1988 2768 -1741 2802
rect -2341 2729 -1741 2768
rect -2341 2695 -2094 2729
rect -2060 2695 -2022 2729
rect -1988 2695 -1741 2729
rect -2341 2656 -1741 2695
rect -2341 2622 -2094 2656
rect -2060 2622 -2022 2656
rect -1988 2622 -1741 2656
rect -2341 2583 -1741 2622
rect -2341 2549 -2094 2583
rect -2060 2549 -2022 2583
rect -1988 2549 -1741 2583
rect -2341 2510 -1741 2549
rect -2341 2476 -2094 2510
rect -2060 2476 -2022 2510
rect -1988 2476 -1741 2510
rect -2341 2437 -1741 2476
rect -2341 2403 -2094 2437
rect -2060 2403 -2022 2437
rect -1988 2403 -1741 2437
rect -2341 2364 -1741 2403
rect -2341 2330 -2094 2364
rect -2060 2330 -2022 2364
rect -1988 2330 -1741 2364
rect -2341 2291 -1741 2330
rect -2341 2257 -2094 2291
rect -2060 2257 -2022 2291
rect -1988 2257 -1741 2291
rect -2341 2218 -1741 2257
rect -2341 2184 -2094 2218
rect -2060 2184 -2022 2218
rect -1988 2184 -1741 2218
rect -2341 2145 -1741 2184
rect -2341 2111 -2094 2145
rect -2060 2111 -2022 2145
rect -1988 2111 -1741 2145
rect -2341 2072 -1741 2111
rect -2341 2038 -2094 2072
rect -2060 2038 -2022 2072
rect -1988 2038 -1741 2072
rect -2341 1999 -1741 2038
rect -2341 1965 -2094 1999
rect -2060 1965 -2022 1999
rect -1988 1965 -1741 1999
rect -2341 1926 -1741 1965
rect -2341 1892 -2094 1926
rect -2060 1892 -2022 1926
rect -1988 1892 -1741 1926
rect -2341 1853 -1741 1892
rect -2341 1819 -2094 1853
rect -2060 1819 -2022 1853
rect -1988 1819 -1741 1853
rect -2341 1780 -1741 1819
rect -2341 1746 -2094 1780
rect -2060 1746 -2022 1780
rect -1988 1746 -1741 1780
rect -2341 1707 -1741 1746
rect -2341 1673 -2094 1707
rect -2060 1673 -2022 1707
rect -1988 1673 -1741 1707
rect -2341 1634 -1741 1673
rect -2341 1600 -2094 1634
rect -2060 1600 -2022 1634
rect -1988 1600 -1741 1634
rect -2341 1561 -1741 1600
rect -2341 1527 -2094 1561
rect -2060 1527 -2022 1561
rect -1988 1527 -1741 1561
rect -2341 1488 -1741 1527
rect -2341 1454 -2094 1488
rect -2060 1454 -2022 1488
rect -1988 1454 -1741 1488
rect -2341 1415 -1741 1454
rect -2341 1381 -2094 1415
rect -2060 1381 -2022 1415
rect -1988 1381 -1741 1415
rect -2341 1342 -1741 1381
rect -2341 1308 -2094 1342
rect -2060 1308 -2022 1342
rect -1988 1308 -1741 1342
rect -2341 1269 -1741 1308
rect -2341 1235 -2094 1269
rect -2060 1235 -2022 1269
rect -1988 1235 -1741 1269
rect -2341 1135 -1741 1235
tri -2341 1131 -2337 1135 ne
rect -2337 1131 -1745 1135
tri -1745 1131 -1741 1135 nw
tri -1439 11333 -1392 11380 se
rect -1392 11333 -886 11380
tri -886 11333 -839 11380 sw
rect -1439 11233 -839 11333
rect -1439 3279 -1192 11233
rect -1086 3279 -839 11233
rect -1439 3240 -839 3279
rect -1439 3206 -1192 3240
rect -1158 3206 -1120 3240
rect -1086 3206 -839 3240
rect -1439 3167 -839 3206
rect -1439 3133 -1192 3167
rect -1158 3133 -1120 3167
rect -1086 3133 -839 3167
rect -1439 3094 -839 3133
rect -1439 3060 -1192 3094
rect -1158 3060 -1120 3094
rect -1086 3060 -839 3094
rect -1439 3021 -839 3060
rect -1439 2987 -1192 3021
rect -1158 2987 -1120 3021
rect -1086 2987 -839 3021
rect -1439 2948 -839 2987
rect -1439 2914 -1192 2948
rect -1158 2914 -1120 2948
rect -1086 2914 -839 2948
rect -1439 2875 -839 2914
rect -1439 2841 -1192 2875
rect -1158 2841 -1120 2875
rect -1086 2841 -839 2875
rect -1439 2802 -839 2841
rect -1439 2768 -1192 2802
rect -1158 2768 -1120 2802
rect -1086 2768 -839 2802
rect -1439 2729 -839 2768
rect -1439 2695 -1192 2729
rect -1158 2695 -1120 2729
rect -1086 2695 -839 2729
rect -1439 2656 -839 2695
rect -1439 2622 -1192 2656
rect -1158 2622 -1120 2656
rect -1086 2622 -839 2656
rect -1439 2583 -839 2622
rect -1439 2549 -1192 2583
rect -1158 2549 -1120 2583
rect -1086 2549 -839 2583
rect -1439 2510 -839 2549
rect -1439 2476 -1192 2510
rect -1158 2476 -1120 2510
rect -1086 2476 -839 2510
rect -1439 2437 -839 2476
rect -1439 2403 -1192 2437
rect -1158 2403 -1120 2437
rect -1086 2403 -839 2437
rect -1439 2364 -839 2403
rect -1439 2330 -1192 2364
rect -1158 2330 -1120 2364
rect -1086 2330 -839 2364
rect -1439 2291 -839 2330
rect -1439 2257 -1192 2291
rect -1158 2257 -1120 2291
rect -1086 2257 -839 2291
rect -1439 2218 -839 2257
rect -1439 2184 -1192 2218
rect -1158 2184 -1120 2218
rect -1086 2184 -839 2218
rect -1439 2145 -839 2184
rect -1439 2111 -1192 2145
rect -1158 2111 -1120 2145
rect -1086 2111 -839 2145
rect -1439 2072 -839 2111
rect -1439 2038 -1192 2072
rect -1158 2038 -1120 2072
rect -1086 2038 -839 2072
rect -1439 1999 -839 2038
rect -1439 1965 -1192 1999
rect -1158 1965 -1120 1999
rect -1086 1965 -839 1999
rect -1439 1926 -839 1965
rect -1439 1892 -1192 1926
rect -1158 1892 -1120 1926
rect -1086 1892 -839 1926
rect -1439 1853 -839 1892
rect -1439 1819 -1192 1853
rect -1158 1819 -1120 1853
rect -1086 1819 -839 1853
rect -1439 1780 -839 1819
rect -1439 1746 -1192 1780
rect -1158 1746 -1120 1780
rect -1086 1746 -839 1780
rect -1439 1707 -839 1746
rect -1439 1673 -1192 1707
rect -1158 1673 -1120 1707
rect -1086 1673 -839 1707
rect -1439 1634 -839 1673
rect -1439 1600 -1192 1634
rect -1158 1600 -1120 1634
rect -1086 1600 -839 1634
rect -1439 1561 -839 1600
rect -1439 1527 -1192 1561
rect -1158 1527 -1120 1561
rect -1086 1527 -839 1561
rect -1439 1488 -839 1527
rect -1439 1454 -1192 1488
rect -1158 1454 -1120 1488
rect -1086 1454 -839 1488
rect -1439 1415 -839 1454
rect -1439 1381 -1192 1415
rect -1158 1381 -1120 1415
rect -1086 1381 -839 1415
rect -1439 1342 -839 1381
rect -1439 1308 -1192 1342
rect -1158 1308 -1120 1342
rect -1086 1308 -839 1342
rect -1439 1269 -839 1308
rect -1439 1235 -1192 1269
rect -1158 1235 -1120 1269
rect -1086 1235 -839 1269
rect -1439 1135 -839 1235
tri -1439 1131 -1435 1135 ne
rect -1435 1131 -843 1135
tri -843 1131 -839 1135 nw
tri -537 11333 -490 11380 se
rect -490 11333 16 11380
tri 16 11333 63 11380 sw
rect -537 11233 63 11333
rect -537 3279 -290 11233
rect -184 3279 63 11233
rect -537 3240 63 3279
rect -537 3206 -290 3240
rect -256 3206 -218 3240
rect -184 3206 63 3240
rect -537 3167 63 3206
rect -537 3133 -290 3167
rect -256 3133 -218 3167
rect -184 3133 63 3167
rect -537 3094 63 3133
rect -537 3060 -290 3094
rect -256 3060 -218 3094
rect -184 3060 63 3094
rect -537 3021 63 3060
rect -537 2987 -290 3021
rect -256 2987 -218 3021
rect -184 2987 63 3021
rect -537 2948 63 2987
rect -537 2914 -290 2948
rect -256 2914 -218 2948
rect -184 2914 63 2948
rect -537 2875 63 2914
rect -537 2841 -290 2875
rect -256 2841 -218 2875
rect -184 2841 63 2875
rect -537 2802 63 2841
rect -537 2768 -290 2802
rect -256 2768 -218 2802
rect -184 2768 63 2802
rect -537 2729 63 2768
rect -537 2695 -290 2729
rect -256 2695 -218 2729
rect -184 2695 63 2729
rect -537 2656 63 2695
rect -537 2622 -290 2656
rect -256 2622 -218 2656
rect -184 2622 63 2656
rect -537 2583 63 2622
rect -537 2549 -290 2583
rect -256 2549 -218 2583
rect -184 2549 63 2583
rect -537 2510 63 2549
rect -537 2476 -290 2510
rect -256 2476 -218 2510
rect -184 2476 63 2510
rect -537 2437 63 2476
rect -537 2403 -290 2437
rect -256 2403 -218 2437
rect -184 2403 63 2437
rect -537 2364 63 2403
rect -537 2330 -290 2364
rect -256 2330 -218 2364
rect -184 2330 63 2364
rect -537 2291 63 2330
rect -537 2257 -290 2291
rect -256 2257 -218 2291
rect -184 2257 63 2291
rect -537 2218 63 2257
rect -537 2184 -290 2218
rect -256 2184 -218 2218
rect -184 2184 63 2218
rect -537 2145 63 2184
rect -537 2111 -290 2145
rect -256 2111 -218 2145
rect -184 2111 63 2145
rect -537 2072 63 2111
rect -537 2038 -290 2072
rect -256 2038 -218 2072
rect -184 2038 63 2072
rect -537 1999 63 2038
rect -537 1965 -290 1999
rect -256 1965 -218 1999
rect -184 1965 63 1999
rect -537 1926 63 1965
rect -537 1892 -290 1926
rect -256 1892 -218 1926
rect -184 1892 63 1926
rect -537 1853 63 1892
rect -537 1819 -290 1853
rect -256 1819 -218 1853
rect -184 1819 63 1853
rect -537 1780 63 1819
rect -537 1746 -290 1780
rect -256 1746 -218 1780
rect -184 1746 63 1780
rect -537 1707 63 1746
rect -537 1673 -290 1707
rect -256 1673 -218 1707
rect -184 1673 63 1707
rect -537 1634 63 1673
rect -537 1600 -290 1634
rect -256 1600 -218 1634
rect -184 1600 63 1634
rect -537 1561 63 1600
rect -537 1527 -290 1561
rect -256 1527 -218 1561
rect -184 1527 63 1561
rect -537 1488 63 1527
rect -537 1454 -290 1488
rect -256 1454 -218 1488
rect -184 1454 63 1488
rect -537 1415 63 1454
rect -537 1381 -290 1415
rect -256 1381 -218 1415
rect -184 1381 63 1415
rect -537 1342 63 1381
rect -537 1308 -290 1342
rect -256 1308 -218 1342
rect -184 1308 63 1342
rect -537 1269 63 1308
rect -537 1235 -290 1269
rect -256 1235 -218 1269
rect -184 1235 63 1269
rect -537 1135 63 1235
tri -537 1131 -533 1135 ne
rect -533 1131 59 1135
tri 59 1131 63 1135 nw
tri 365 11333 412 11380 se
rect 412 11333 918 11380
tri 918 11333 965 11380 sw
rect 365 11233 965 11333
rect 365 3279 612 11233
rect 718 3279 965 11233
rect 365 3240 965 3279
rect 365 3206 612 3240
rect 646 3206 684 3240
rect 718 3206 965 3240
rect 365 3167 965 3206
rect 365 3133 612 3167
rect 646 3133 684 3167
rect 718 3133 965 3167
rect 365 3094 965 3133
rect 365 3060 612 3094
rect 646 3060 684 3094
rect 718 3060 965 3094
rect 365 3021 965 3060
rect 365 2987 612 3021
rect 646 2987 684 3021
rect 718 2987 965 3021
rect 365 2948 965 2987
rect 365 2914 612 2948
rect 646 2914 684 2948
rect 718 2914 965 2948
rect 365 2875 965 2914
rect 365 2841 612 2875
rect 646 2841 684 2875
rect 718 2841 965 2875
rect 365 2802 965 2841
rect 365 2768 612 2802
rect 646 2768 684 2802
rect 718 2768 965 2802
rect 365 2729 965 2768
rect 365 2695 612 2729
rect 646 2695 684 2729
rect 718 2695 965 2729
rect 365 2656 965 2695
rect 365 2622 612 2656
rect 646 2622 684 2656
rect 718 2622 965 2656
rect 365 2583 965 2622
rect 365 2549 612 2583
rect 646 2549 684 2583
rect 718 2549 965 2583
rect 365 2510 965 2549
rect 365 2476 612 2510
rect 646 2476 684 2510
rect 718 2476 965 2510
rect 365 2437 965 2476
rect 365 2403 612 2437
rect 646 2403 684 2437
rect 718 2403 965 2437
rect 365 2364 965 2403
rect 365 2330 612 2364
rect 646 2330 684 2364
rect 718 2330 965 2364
rect 365 2291 965 2330
rect 365 2257 612 2291
rect 646 2257 684 2291
rect 718 2257 965 2291
rect 365 2218 965 2257
rect 365 2184 612 2218
rect 646 2184 684 2218
rect 718 2184 965 2218
rect 365 2145 965 2184
rect 365 2111 612 2145
rect 646 2111 684 2145
rect 718 2111 965 2145
rect 365 2072 965 2111
rect 365 2038 612 2072
rect 646 2038 684 2072
rect 718 2038 965 2072
rect 365 1999 965 2038
rect 365 1965 612 1999
rect 646 1965 684 1999
rect 718 1965 965 1999
rect 365 1926 965 1965
rect 365 1892 612 1926
rect 646 1892 684 1926
rect 718 1892 965 1926
rect 365 1853 965 1892
rect 365 1819 612 1853
rect 646 1819 684 1853
rect 718 1819 965 1853
rect 365 1780 965 1819
rect 365 1746 612 1780
rect 646 1746 684 1780
rect 718 1746 965 1780
rect 365 1707 965 1746
rect 365 1673 612 1707
rect 646 1673 684 1707
rect 718 1673 965 1707
rect 365 1634 965 1673
rect 365 1600 612 1634
rect 646 1600 684 1634
rect 718 1600 965 1634
rect 365 1561 965 1600
rect 365 1527 612 1561
rect 646 1527 684 1561
rect 718 1527 965 1561
rect 365 1488 965 1527
rect 365 1454 612 1488
rect 646 1454 684 1488
rect 718 1454 965 1488
rect 365 1415 965 1454
rect 365 1381 612 1415
rect 646 1381 684 1415
rect 718 1381 965 1415
rect 365 1342 965 1381
rect 365 1308 612 1342
rect 646 1308 684 1342
rect 718 1308 965 1342
rect 365 1269 965 1308
rect 365 1235 612 1269
rect 646 1235 684 1269
rect 718 1235 965 1269
rect 365 1135 965 1235
tri 365 1131 369 1135 ne
rect 369 1131 961 1135
tri 961 1131 965 1135 nw
tri 1267 11333 1314 11380 se
rect 1314 11333 1820 11380
tri 1820 11333 1867 11380 sw
rect 1267 11233 1867 11333
rect 1267 3279 1514 11233
rect 1620 3279 1867 11233
rect 1267 3240 1867 3279
rect 1267 3206 1514 3240
rect 1548 3206 1586 3240
rect 1620 3206 1867 3240
rect 1267 3167 1867 3206
rect 1267 3133 1514 3167
rect 1548 3133 1586 3167
rect 1620 3133 1867 3167
rect 1267 3094 1867 3133
rect 1267 3060 1514 3094
rect 1548 3060 1586 3094
rect 1620 3060 1867 3094
rect 1267 3021 1867 3060
rect 1267 2987 1514 3021
rect 1548 2987 1586 3021
rect 1620 2987 1867 3021
rect 1267 2948 1867 2987
rect 1267 2914 1514 2948
rect 1548 2914 1586 2948
rect 1620 2914 1867 2948
rect 1267 2875 1867 2914
rect 1267 2841 1514 2875
rect 1548 2841 1586 2875
rect 1620 2841 1867 2875
rect 1267 2802 1867 2841
rect 1267 2768 1514 2802
rect 1548 2768 1586 2802
rect 1620 2768 1867 2802
rect 1267 2729 1867 2768
rect 1267 2695 1514 2729
rect 1548 2695 1586 2729
rect 1620 2695 1867 2729
rect 1267 2656 1867 2695
rect 1267 2622 1514 2656
rect 1548 2622 1586 2656
rect 1620 2622 1867 2656
rect 1267 2583 1867 2622
rect 1267 2549 1514 2583
rect 1548 2549 1586 2583
rect 1620 2549 1867 2583
rect 1267 2510 1867 2549
rect 1267 2476 1514 2510
rect 1548 2476 1586 2510
rect 1620 2476 1867 2510
rect 1267 2437 1867 2476
rect 1267 2403 1514 2437
rect 1548 2403 1586 2437
rect 1620 2403 1867 2437
rect 1267 2364 1867 2403
rect 1267 2330 1514 2364
rect 1548 2330 1586 2364
rect 1620 2330 1867 2364
rect 1267 2291 1867 2330
rect 1267 2257 1514 2291
rect 1548 2257 1586 2291
rect 1620 2257 1867 2291
rect 1267 2218 1867 2257
rect 1267 2184 1514 2218
rect 1548 2184 1586 2218
rect 1620 2184 1867 2218
rect 1267 2145 1867 2184
rect 1267 2111 1514 2145
rect 1548 2111 1586 2145
rect 1620 2111 1867 2145
rect 1267 2072 1867 2111
rect 1267 2038 1514 2072
rect 1548 2038 1586 2072
rect 1620 2038 1867 2072
rect 1267 1999 1867 2038
rect 1267 1965 1514 1999
rect 1548 1965 1586 1999
rect 1620 1965 1867 1999
rect 1267 1926 1867 1965
rect 1267 1892 1514 1926
rect 1548 1892 1586 1926
rect 1620 1892 1867 1926
rect 1267 1853 1867 1892
rect 1267 1819 1514 1853
rect 1548 1819 1586 1853
rect 1620 1819 1867 1853
rect 1267 1780 1867 1819
rect 1267 1746 1514 1780
rect 1548 1746 1586 1780
rect 1620 1746 1867 1780
rect 1267 1707 1867 1746
rect 1267 1673 1514 1707
rect 1548 1673 1586 1707
rect 1620 1673 1867 1707
rect 1267 1634 1867 1673
rect 1267 1600 1514 1634
rect 1548 1600 1586 1634
rect 1620 1600 1867 1634
rect 1267 1561 1867 1600
rect 1267 1527 1514 1561
rect 1548 1527 1586 1561
rect 1620 1527 1867 1561
rect 1267 1488 1867 1527
rect 1267 1454 1514 1488
rect 1548 1454 1586 1488
rect 1620 1454 1867 1488
rect 1267 1415 1867 1454
rect 1267 1381 1514 1415
rect 1548 1381 1586 1415
rect 1620 1381 1867 1415
rect 1267 1342 1867 1381
rect 1267 1308 1514 1342
rect 1548 1308 1586 1342
rect 1620 1308 1867 1342
rect 1267 1269 1867 1308
rect 1267 1235 1514 1269
rect 1548 1235 1586 1269
rect 1620 1235 1867 1269
rect 1267 1135 1867 1235
tri 1267 1131 1271 1135 ne
rect 1271 1131 1863 1135
tri 1863 1131 1867 1135 nw
tri 2169 11333 2216 11380 se
rect 2216 11333 2722 11380
tri 2722 11333 2769 11380 sw
rect 2169 11233 2769 11333
rect 2169 3279 2416 11233
rect 2522 3279 2769 11233
rect 2169 3240 2769 3279
rect 2169 3206 2416 3240
rect 2450 3206 2488 3240
rect 2522 3206 2769 3240
rect 2169 3167 2769 3206
rect 2169 3133 2416 3167
rect 2450 3133 2488 3167
rect 2522 3133 2769 3167
rect 2169 3094 2769 3133
rect 2169 3060 2416 3094
rect 2450 3060 2488 3094
rect 2522 3060 2769 3094
rect 2169 3021 2769 3060
rect 2169 2987 2416 3021
rect 2450 2987 2488 3021
rect 2522 2987 2769 3021
rect 2169 2948 2769 2987
rect 2169 2914 2416 2948
rect 2450 2914 2488 2948
rect 2522 2914 2769 2948
rect 2169 2875 2769 2914
rect 2169 2841 2416 2875
rect 2450 2841 2488 2875
rect 2522 2841 2769 2875
rect 2169 2802 2769 2841
rect 2169 2768 2416 2802
rect 2450 2768 2488 2802
rect 2522 2768 2769 2802
rect 2169 2729 2769 2768
rect 2169 2695 2416 2729
rect 2450 2695 2488 2729
rect 2522 2695 2769 2729
rect 2169 2656 2769 2695
rect 2169 2622 2416 2656
rect 2450 2622 2488 2656
rect 2522 2622 2769 2656
rect 2169 2583 2769 2622
rect 2169 2549 2416 2583
rect 2450 2549 2488 2583
rect 2522 2549 2769 2583
rect 2169 2510 2769 2549
rect 2169 2476 2416 2510
rect 2450 2476 2488 2510
rect 2522 2476 2769 2510
rect 2169 2437 2769 2476
rect 2169 2403 2416 2437
rect 2450 2403 2488 2437
rect 2522 2403 2769 2437
rect 2169 2364 2769 2403
rect 2169 2330 2416 2364
rect 2450 2330 2488 2364
rect 2522 2330 2769 2364
rect 2169 2291 2769 2330
rect 2169 2257 2416 2291
rect 2450 2257 2488 2291
rect 2522 2257 2769 2291
rect 2169 2218 2769 2257
rect 2169 2184 2416 2218
rect 2450 2184 2488 2218
rect 2522 2184 2769 2218
rect 2169 2145 2769 2184
rect 2169 2111 2416 2145
rect 2450 2111 2488 2145
rect 2522 2111 2769 2145
rect 2169 2072 2769 2111
rect 2169 2038 2416 2072
rect 2450 2038 2488 2072
rect 2522 2038 2769 2072
rect 2169 1999 2769 2038
rect 2169 1965 2416 1999
rect 2450 1965 2488 1999
rect 2522 1965 2769 1999
rect 2169 1926 2769 1965
rect 2169 1892 2416 1926
rect 2450 1892 2488 1926
rect 2522 1892 2769 1926
rect 2169 1853 2769 1892
rect 2169 1819 2416 1853
rect 2450 1819 2488 1853
rect 2522 1819 2769 1853
rect 2169 1780 2769 1819
rect 2169 1746 2416 1780
rect 2450 1746 2488 1780
rect 2522 1746 2769 1780
rect 2169 1707 2769 1746
rect 2169 1673 2416 1707
rect 2450 1673 2488 1707
rect 2522 1673 2769 1707
rect 2169 1634 2769 1673
rect 2169 1600 2416 1634
rect 2450 1600 2488 1634
rect 2522 1600 2769 1634
rect 2169 1561 2769 1600
rect 2169 1527 2416 1561
rect 2450 1527 2488 1561
rect 2522 1527 2769 1561
rect 2169 1488 2769 1527
rect 2169 1454 2416 1488
rect 2450 1454 2488 1488
rect 2522 1454 2769 1488
rect 2169 1415 2769 1454
rect 2169 1381 2416 1415
rect 2450 1381 2488 1415
rect 2522 1381 2769 1415
rect 2169 1342 2769 1381
rect 2169 1308 2416 1342
rect 2450 1308 2488 1342
rect 2522 1308 2769 1342
rect 2169 1269 2769 1308
rect 2169 1235 2416 1269
rect 2450 1235 2488 1269
rect 2522 1235 2769 1269
rect 2169 1135 2769 1235
tri 2169 1131 2173 1135 ne
rect 2173 1131 2765 1135
tri 2765 1131 2769 1135 nw
tri 3071 11333 3118 11380 se
rect 3118 11333 3624 11380
tri 3624 11333 3671 11380 sw
rect 3071 11233 3671 11333
rect 3071 3279 3318 11233
rect 3424 3279 3671 11233
rect 3071 3240 3671 3279
rect 3071 3206 3318 3240
rect 3352 3206 3390 3240
rect 3424 3206 3671 3240
rect 3071 3167 3671 3206
rect 3071 3133 3318 3167
rect 3352 3133 3390 3167
rect 3424 3133 3671 3167
rect 3071 3094 3671 3133
rect 3071 3060 3318 3094
rect 3352 3060 3390 3094
rect 3424 3060 3671 3094
rect 3071 3021 3671 3060
rect 3071 2987 3318 3021
rect 3352 2987 3390 3021
rect 3424 2987 3671 3021
rect 3071 2948 3671 2987
rect 3071 2914 3318 2948
rect 3352 2914 3390 2948
rect 3424 2914 3671 2948
rect 3071 2875 3671 2914
rect 3071 2841 3318 2875
rect 3352 2841 3390 2875
rect 3424 2841 3671 2875
rect 3071 2802 3671 2841
rect 3071 2768 3318 2802
rect 3352 2768 3390 2802
rect 3424 2768 3671 2802
rect 3071 2729 3671 2768
rect 3071 2695 3318 2729
rect 3352 2695 3390 2729
rect 3424 2695 3671 2729
rect 3071 2656 3671 2695
rect 3071 2622 3318 2656
rect 3352 2622 3390 2656
rect 3424 2622 3671 2656
rect 3071 2583 3671 2622
rect 3071 2549 3318 2583
rect 3352 2549 3390 2583
rect 3424 2549 3671 2583
rect 3071 2510 3671 2549
rect 3071 2476 3318 2510
rect 3352 2476 3390 2510
rect 3424 2476 3671 2510
rect 3071 2437 3671 2476
rect 3071 2403 3318 2437
rect 3352 2403 3390 2437
rect 3424 2403 3671 2437
rect 3071 2364 3671 2403
rect 3071 2330 3318 2364
rect 3352 2330 3390 2364
rect 3424 2330 3671 2364
rect 3071 2291 3671 2330
rect 3071 2257 3318 2291
rect 3352 2257 3390 2291
rect 3424 2257 3671 2291
rect 3071 2218 3671 2257
rect 3071 2184 3318 2218
rect 3352 2184 3390 2218
rect 3424 2184 3671 2218
rect 3071 2145 3671 2184
rect 3071 2111 3318 2145
rect 3352 2111 3390 2145
rect 3424 2111 3671 2145
rect 3071 2072 3671 2111
rect 3071 2038 3318 2072
rect 3352 2038 3390 2072
rect 3424 2038 3671 2072
rect 3071 1999 3671 2038
rect 3071 1965 3318 1999
rect 3352 1965 3390 1999
rect 3424 1965 3671 1999
rect 3071 1926 3671 1965
rect 3071 1892 3318 1926
rect 3352 1892 3390 1926
rect 3424 1892 3671 1926
rect 3071 1853 3671 1892
rect 3071 1819 3318 1853
rect 3352 1819 3390 1853
rect 3424 1819 3671 1853
rect 3071 1780 3671 1819
rect 3071 1746 3318 1780
rect 3352 1746 3390 1780
rect 3424 1746 3671 1780
rect 3071 1707 3671 1746
rect 3071 1673 3318 1707
rect 3352 1673 3390 1707
rect 3424 1673 3671 1707
rect 3071 1634 3671 1673
rect 3071 1600 3318 1634
rect 3352 1600 3390 1634
rect 3424 1600 3671 1634
rect 3071 1561 3671 1600
rect 3071 1527 3318 1561
rect 3352 1527 3390 1561
rect 3424 1527 3671 1561
rect 3071 1488 3671 1527
rect 3071 1454 3318 1488
rect 3352 1454 3390 1488
rect 3424 1454 3671 1488
rect 3071 1415 3671 1454
rect 3071 1381 3318 1415
rect 3352 1381 3390 1415
rect 3424 1381 3671 1415
rect 3071 1342 3671 1381
rect 3071 1308 3318 1342
rect 3352 1308 3390 1342
rect 3424 1308 3671 1342
rect 3071 1269 3671 1308
rect 3071 1235 3318 1269
rect 3352 1235 3390 1269
rect 3424 1235 3671 1269
rect 3071 1135 3671 1235
tri 3071 1131 3075 1135 ne
rect 3075 1131 3667 1135
tri 3667 1131 3671 1135 nw
tri 3973 11333 4020 11380 se
rect 4020 11333 4526 11380
tri 4526 11333 4573 11380 sw
rect 3973 11233 4573 11333
rect 3973 3279 4220 11233
rect 4326 3279 4573 11233
rect 3973 3240 4573 3279
rect 3973 3206 4220 3240
rect 4254 3206 4292 3240
rect 4326 3206 4573 3240
rect 3973 3167 4573 3206
rect 3973 3133 4220 3167
rect 4254 3133 4292 3167
rect 4326 3133 4573 3167
rect 3973 3094 4573 3133
rect 3973 3060 4220 3094
rect 4254 3060 4292 3094
rect 4326 3060 4573 3094
rect 3973 3021 4573 3060
rect 3973 2987 4220 3021
rect 4254 2987 4292 3021
rect 4326 2987 4573 3021
rect 3973 2948 4573 2987
rect 3973 2914 4220 2948
rect 4254 2914 4292 2948
rect 4326 2914 4573 2948
rect 3973 2875 4573 2914
rect 3973 2841 4220 2875
rect 4254 2841 4292 2875
rect 4326 2841 4573 2875
rect 3973 2802 4573 2841
rect 3973 2768 4220 2802
rect 4254 2768 4292 2802
rect 4326 2768 4573 2802
rect 3973 2729 4573 2768
rect 3973 2695 4220 2729
rect 4254 2695 4292 2729
rect 4326 2695 4573 2729
rect 3973 2656 4573 2695
rect 3973 2622 4220 2656
rect 4254 2622 4292 2656
rect 4326 2622 4573 2656
rect 3973 2583 4573 2622
rect 3973 2549 4220 2583
rect 4254 2549 4292 2583
rect 4326 2549 4573 2583
rect 3973 2510 4573 2549
rect 3973 2476 4220 2510
rect 4254 2476 4292 2510
rect 4326 2476 4573 2510
rect 3973 2437 4573 2476
rect 3973 2403 4220 2437
rect 4254 2403 4292 2437
rect 4326 2403 4573 2437
rect 3973 2364 4573 2403
rect 3973 2330 4220 2364
rect 4254 2330 4292 2364
rect 4326 2330 4573 2364
rect 3973 2291 4573 2330
rect 3973 2257 4220 2291
rect 4254 2257 4292 2291
rect 4326 2257 4573 2291
rect 3973 2218 4573 2257
rect 3973 2184 4220 2218
rect 4254 2184 4292 2218
rect 4326 2184 4573 2218
rect 3973 2145 4573 2184
rect 3973 2111 4220 2145
rect 4254 2111 4292 2145
rect 4326 2111 4573 2145
rect 3973 2072 4573 2111
rect 3973 2038 4220 2072
rect 4254 2038 4292 2072
rect 4326 2038 4573 2072
rect 3973 1999 4573 2038
rect 3973 1965 4220 1999
rect 4254 1965 4292 1999
rect 4326 1965 4573 1999
rect 3973 1926 4573 1965
rect 3973 1892 4220 1926
rect 4254 1892 4292 1926
rect 4326 1892 4573 1926
rect 3973 1853 4573 1892
rect 3973 1819 4220 1853
rect 4254 1819 4292 1853
rect 4326 1819 4573 1853
rect 3973 1780 4573 1819
rect 3973 1746 4220 1780
rect 4254 1746 4292 1780
rect 4326 1746 4573 1780
rect 3973 1707 4573 1746
rect 3973 1673 4220 1707
rect 4254 1673 4292 1707
rect 4326 1673 4573 1707
rect 3973 1634 4573 1673
rect 3973 1600 4220 1634
rect 4254 1600 4292 1634
rect 4326 1600 4573 1634
rect 3973 1561 4573 1600
rect 3973 1527 4220 1561
rect 4254 1527 4292 1561
rect 4326 1527 4573 1561
rect 3973 1488 4573 1527
rect 3973 1454 4220 1488
rect 4254 1454 4292 1488
rect 4326 1454 4573 1488
rect 3973 1415 4573 1454
rect 3973 1381 4220 1415
rect 4254 1381 4292 1415
rect 4326 1381 4573 1415
rect 3973 1342 4573 1381
rect 3973 1308 4220 1342
rect 4254 1308 4292 1342
rect 4326 1308 4573 1342
rect 3973 1269 4573 1308
rect 3973 1235 4220 1269
rect 4254 1235 4292 1269
rect 4326 1235 4573 1269
rect 3973 1135 4573 1235
tri 3973 1131 3977 1135 ne
rect 3977 1131 4569 1135
tri 4569 1131 4573 1135 nw
tri 4875 11333 4922 11380 se
rect 4922 11333 5428 11380
tri 5428 11333 5475 11380 sw
rect 4875 11233 5475 11333
rect 4875 3279 5122 11233
rect 5228 3279 5475 11233
rect 4875 3240 5475 3279
rect 4875 3206 5122 3240
rect 5156 3206 5194 3240
rect 5228 3206 5475 3240
rect 4875 3167 5475 3206
rect 4875 3133 5122 3167
rect 5156 3133 5194 3167
rect 5228 3133 5475 3167
rect 4875 3094 5475 3133
rect 4875 3060 5122 3094
rect 5156 3060 5194 3094
rect 5228 3060 5475 3094
rect 4875 3021 5475 3060
rect 4875 2987 5122 3021
rect 5156 2987 5194 3021
rect 5228 2987 5475 3021
rect 4875 2948 5475 2987
rect 4875 2914 5122 2948
rect 5156 2914 5194 2948
rect 5228 2914 5475 2948
rect 4875 2875 5475 2914
rect 4875 2841 5122 2875
rect 5156 2841 5194 2875
rect 5228 2841 5475 2875
rect 4875 2802 5475 2841
rect 4875 2768 5122 2802
rect 5156 2768 5194 2802
rect 5228 2768 5475 2802
rect 4875 2729 5475 2768
rect 4875 2695 5122 2729
rect 5156 2695 5194 2729
rect 5228 2695 5475 2729
rect 4875 2656 5475 2695
rect 4875 2622 5122 2656
rect 5156 2622 5194 2656
rect 5228 2622 5475 2656
rect 4875 2583 5475 2622
rect 4875 2549 5122 2583
rect 5156 2549 5194 2583
rect 5228 2549 5475 2583
rect 4875 2510 5475 2549
rect 4875 2476 5122 2510
rect 5156 2476 5194 2510
rect 5228 2476 5475 2510
rect 4875 2437 5475 2476
rect 4875 2403 5122 2437
rect 5156 2403 5194 2437
rect 5228 2403 5475 2437
rect 4875 2364 5475 2403
rect 4875 2330 5122 2364
rect 5156 2330 5194 2364
rect 5228 2330 5475 2364
rect 4875 2291 5475 2330
rect 4875 2257 5122 2291
rect 5156 2257 5194 2291
rect 5228 2257 5475 2291
rect 4875 2218 5475 2257
rect 4875 2184 5122 2218
rect 5156 2184 5194 2218
rect 5228 2184 5475 2218
rect 4875 2145 5475 2184
rect 4875 2111 5122 2145
rect 5156 2111 5194 2145
rect 5228 2111 5475 2145
rect 4875 2072 5475 2111
rect 4875 2038 5122 2072
rect 5156 2038 5194 2072
rect 5228 2038 5475 2072
rect 4875 1999 5475 2038
rect 4875 1965 5122 1999
rect 5156 1965 5194 1999
rect 5228 1965 5475 1999
rect 4875 1926 5475 1965
rect 4875 1892 5122 1926
rect 5156 1892 5194 1926
rect 5228 1892 5475 1926
rect 4875 1853 5475 1892
rect 4875 1819 5122 1853
rect 5156 1819 5194 1853
rect 5228 1819 5475 1853
rect 4875 1780 5475 1819
rect 4875 1746 5122 1780
rect 5156 1746 5194 1780
rect 5228 1746 5475 1780
rect 4875 1707 5475 1746
rect 4875 1673 5122 1707
rect 5156 1673 5194 1707
rect 5228 1673 5475 1707
rect 4875 1634 5475 1673
rect 4875 1600 5122 1634
rect 5156 1600 5194 1634
rect 5228 1600 5475 1634
rect 4875 1561 5475 1600
rect 4875 1527 5122 1561
rect 5156 1527 5194 1561
rect 5228 1527 5475 1561
rect 4875 1488 5475 1527
rect 4875 1454 5122 1488
rect 5156 1454 5194 1488
rect 5228 1454 5475 1488
rect 4875 1415 5475 1454
rect 4875 1381 5122 1415
rect 5156 1381 5194 1415
rect 5228 1381 5475 1415
rect 4875 1342 5475 1381
rect 4875 1308 5122 1342
rect 5156 1308 5194 1342
rect 5228 1308 5475 1342
rect 4875 1269 5475 1308
rect 4875 1235 5122 1269
rect 5156 1235 5194 1269
rect 5228 1235 5475 1269
rect 4875 1135 5475 1235
tri 4875 1131 4879 1135 ne
rect 4879 1131 5471 1135
tri 5471 1131 5475 1135 nw
tri 5777 11333 5824 11380 se
rect 5824 11333 6330 11380
tri 6330 11333 6377 11380 sw
rect 5777 11233 6377 11333
rect 5777 3279 6024 11233
rect 6130 3279 6377 11233
rect 5777 3240 6377 3279
rect 5777 3206 6024 3240
rect 6058 3206 6096 3240
rect 6130 3206 6377 3240
rect 5777 3167 6377 3206
rect 5777 3133 6024 3167
rect 6058 3133 6096 3167
rect 6130 3133 6377 3167
rect 5777 3094 6377 3133
rect 5777 3060 6024 3094
rect 6058 3060 6096 3094
rect 6130 3060 6377 3094
rect 5777 3021 6377 3060
rect 5777 2987 6024 3021
rect 6058 2987 6096 3021
rect 6130 2987 6377 3021
rect 5777 2948 6377 2987
rect 5777 2914 6024 2948
rect 6058 2914 6096 2948
rect 6130 2914 6377 2948
rect 5777 2875 6377 2914
rect 5777 2841 6024 2875
rect 6058 2841 6096 2875
rect 6130 2841 6377 2875
rect 5777 2802 6377 2841
rect 5777 2768 6024 2802
rect 6058 2768 6096 2802
rect 6130 2768 6377 2802
rect 5777 2729 6377 2768
rect 5777 2695 6024 2729
rect 6058 2695 6096 2729
rect 6130 2695 6377 2729
rect 5777 2656 6377 2695
rect 5777 2622 6024 2656
rect 6058 2622 6096 2656
rect 6130 2622 6377 2656
rect 5777 2583 6377 2622
rect 5777 2549 6024 2583
rect 6058 2549 6096 2583
rect 6130 2549 6377 2583
rect 5777 2510 6377 2549
rect 5777 2476 6024 2510
rect 6058 2476 6096 2510
rect 6130 2476 6377 2510
rect 5777 2437 6377 2476
rect 5777 2403 6024 2437
rect 6058 2403 6096 2437
rect 6130 2403 6377 2437
rect 5777 2364 6377 2403
rect 5777 2330 6024 2364
rect 6058 2330 6096 2364
rect 6130 2330 6377 2364
rect 5777 2291 6377 2330
rect 5777 2257 6024 2291
rect 6058 2257 6096 2291
rect 6130 2257 6377 2291
rect 5777 2218 6377 2257
rect 5777 2184 6024 2218
rect 6058 2184 6096 2218
rect 6130 2184 6377 2218
rect 5777 2145 6377 2184
rect 5777 2111 6024 2145
rect 6058 2111 6096 2145
rect 6130 2111 6377 2145
rect 5777 2072 6377 2111
rect 5777 2038 6024 2072
rect 6058 2038 6096 2072
rect 6130 2038 6377 2072
rect 5777 1999 6377 2038
rect 5777 1965 6024 1999
rect 6058 1965 6096 1999
rect 6130 1965 6377 1999
rect 5777 1926 6377 1965
rect 5777 1892 6024 1926
rect 6058 1892 6096 1926
rect 6130 1892 6377 1926
rect 5777 1853 6377 1892
rect 5777 1819 6024 1853
rect 6058 1819 6096 1853
rect 6130 1819 6377 1853
rect 5777 1780 6377 1819
rect 5777 1746 6024 1780
rect 6058 1746 6096 1780
rect 6130 1746 6377 1780
rect 5777 1707 6377 1746
rect 5777 1673 6024 1707
rect 6058 1673 6096 1707
rect 6130 1673 6377 1707
rect 5777 1634 6377 1673
rect 5777 1600 6024 1634
rect 6058 1600 6096 1634
rect 6130 1600 6377 1634
rect 5777 1561 6377 1600
rect 5777 1527 6024 1561
rect 6058 1527 6096 1561
rect 6130 1527 6377 1561
rect 5777 1488 6377 1527
rect 5777 1454 6024 1488
rect 6058 1454 6096 1488
rect 6130 1454 6377 1488
rect 5777 1415 6377 1454
rect 5777 1381 6024 1415
rect 6058 1381 6096 1415
rect 6130 1381 6377 1415
rect 5777 1342 6377 1381
rect 5777 1308 6024 1342
rect 6058 1308 6096 1342
rect 6130 1308 6377 1342
rect 5777 1269 6377 1308
rect 5777 1235 6024 1269
rect 6058 1235 6096 1269
rect 6130 1235 6377 1269
rect 5777 1135 6377 1235
tri 5777 1131 5781 1135 ne
rect 5781 1131 6373 1135
tri 6373 1131 6377 1135 nw
tri 6679 11333 6726 11380 se
rect 6726 11333 7232 11380
tri 7232 11333 7279 11380 sw
rect 6679 11233 7279 11333
rect 6679 3279 6926 11233
rect 7032 3279 7279 11233
rect 6679 3240 7279 3279
rect 6679 3206 6926 3240
rect 6960 3206 6998 3240
rect 7032 3206 7279 3240
rect 6679 3167 7279 3206
rect 6679 3133 6926 3167
rect 6960 3133 6998 3167
rect 7032 3133 7279 3167
rect 6679 3094 7279 3133
rect 6679 3060 6926 3094
rect 6960 3060 6998 3094
rect 7032 3060 7279 3094
rect 6679 3021 7279 3060
rect 6679 2987 6926 3021
rect 6960 2987 6998 3021
rect 7032 2987 7279 3021
rect 6679 2948 7279 2987
rect 6679 2914 6926 2948
rect 6960 2914 6998 2948
rect 7032 2914 7279 2948
rect 6679 2875 7279 2914
rect 6679 2841 6926 2875
rect 6960 2841 6998 2875
rect 7032 2841 7279 2875
rect 6679 2802 7279 2841
rect 6679 2768 6926 2802
rect 6960 2768 6998 2802
rect 7032 2768 7279 2802
rect 6679 2729 7279 2768
rect 6679 2695 6926 2729
rect 6960 2695 6998 2729
rect 7032 2695 7279 2729
rect 6679 2656 7279 2695
rect 6679 2622 6926 2656
rect 6960 2622 6998 2656
rect 7032 2622 7279 2656
rect 6679 2583 7279 2622
rect 6679 2549 6926 2583
rect 6960 2549 6998 2583
rect 7032 2549 7279 2583
rect 6679 2510 7279 2549
rect 6679 2476 6926 2510
rect 6960 2476 6998 2510
rect 7032 2476 7279 2510
rect 6679 2437 7279 2476
rect 6679 2403 6926 2437
rect 6960 2403 6998 2437
rect 7032 2403 7279 2437
rect 6679 2364 7279 2403
rect 6679 2330 6926 2364
rect 6960 2330 6998 2364
rect 7032 2330 7279 2364
rect 6679 2291 7279 2330
rect 6679 2257 6926 2291
rect 6960 2257 6998 2291
rect 7032 2257 7279 2291
rect 6679 2218 7279 2257
rect 6679 2184 6926 2218
rect 6960 2184 6998 2218
rect 7032 2184 7279 2218
rect 6679 2145 7279 2184
rect 6679 2111 6926 2145
rect 6960 2111 6998 2145
rect 7032 2111 7279 2145
rect 6679 2072 7279 2111
rect 6679 2038 6926 2072
rect 6960 2038 6998 2072
rect 7032 2038 7279 2072
rect 6679 1999 7279 2038
rect 6679 1965 6926 1999
rect 6960 1965 6998 1999
rect 7032 1965 7279 1999
rect 6679 1926 7279 1965
rect 6679 1892 6926 1926
rect 6960 1892 6998 1926
rect 7032 1892 7279 1926
rect 6679 1853 7279 1892
rect 6679 1819 6926 1853
rect 6960 1819 6998 1853
rect 7032 1819 7279 1853
rect 6679 1780 7279 1819
rect 6679 1746 6926 1780
rect 6960 1746 6998 1780
rect 7032 1746 7279 1780
rect 6679 1707 7279 1746
rect 6679 1673 6926 1707
rect 6960 1673 6998 1707
rect 7032 1673 7279 1707
rect 6679 1634 7279 1673
rect 6679 1600 6926 1634
rect 6960 1600 6998 1634
rect 7032 1600 7279 1634
rect 6679 1561 7279 1600
rect 6679 1527 6926 1561
rect 6960 1527 6998 1561
rect 7032 1527 7279 1561
rect 6679 1488 7279 1527
rect 6679 1454 6926 1488
rect 6960 1454 6998 1488
rect 7032 1454 7279 1488
rect 6679 1415 7279 1454
rect 6679 1381 6926 1415
rect 6960 1381 6998 1415
rect 7032 1381 7279 1415
rect 6679 1342 7279 1381
rect 6679 1308 6926 1342
rect 6960 1308 6998 1342
rect 7032 1308 7279 1342
rect 6679 1269 7279 1308
rect 6679 1235 6926 1269
rect 6960 1235 6998 1269
rect 7032 1235 7279 1269
rect 6679 1135 7279 1235
tri 6679 1131 6683 1135 ne
rect 6683 1131 7275 1135
tri 7275 1131 7279 1135 nw
tri 7581 11333 7628 11380 se
rect 7628 11333 8134 11380
tri 8134 11333 8181 11380 sw
rect 7581 11233 8181 11333
rect 7581 3279 7828 11233
rect 7934 3279 8181 11233
rect 7581 3240 8181 3279
rect 7581 3206 7828 3240
rect 7862 3206 7900 3240
rect 7934 3206 8181 3240
rect 7581 3167 8181 3206
rect 7581 3133 7828 3167
rect 7862 3133 7900 3167
rect 7934 3133 8181 3167
rect 7581 3094 8181 3133
rect 7581 3060 7828 3094
rect 7862 3060 7900 3094
rect 7934 3060 8181 3094
rect 7581 3021 8181 3060
rect 7581 2987 7828 3021
rect 7862 2987 7900 3021
rect 7934 2987 8181 3021
rect 7581 2948 8181 2987
rect 7581 2914 7828 2948
rect 7862 2914 7900 2948
rect 7934 2914 8181 2948
rect 7581 2875 8181 2914
rect 7581 2841 7828 2875
rect 7862 2841 7900 2875
rect 7934 2841 8181 2875
rect 7581 2802 8181 2841
rect 7581 2768 7828 2802
rect 7862 2768 7900 2802
rect 7934 2768 8181 2802
rect 7581 2729 8181 2768
rect 7581 2695 7828 2729
rect 7862 2695 7900 2729
rect 7934 2695 8181 2729
rect 7581 2656 8181 2695
rect 7581 2622 7828 2656
rect 7862 2622 7900 2656
rect 7934 2622 8181 2656
rect 7581 2583 8181 2622
rect 7581 2549 7828 2583
rect 7862 2549 7900 2583
rect 7934 2549 8181 2583
rect 7581 2510 8181 2549
rect 7581 2476 7828 2510
rect 7862 2476 7900 2510
rect 7934 2476 8181 2510
rect 7581 2437 8181 2476
rect 7581 2403 7828 2437
rect 7862 2403 7900 2437
rect 7934 2403 8181 2437
rect 7581 2364 8181 2403
rect 7581 2330 7828 2364
rect 7862 2330 7900 2364
rect 7934 2330 8181 2364
rect 7581 2291 8181 2330
rect 7581 2257 7828 2291
rect 7862 2257 7900 2291
rect 7934 2257 8181 2291
rect 7581 2218 8181 2257
rect 7581 2184 7828 2218
rect 7862 2184 7900 2218
rect 7934 2184 8181 2218
rect 7581 2145 8181 2184
rect 7581 2111 7828 2145
rect 7862 2111 7900 2145
rect 7934 2111 8181 2145
rect 7581 2072 8181 2111
rect 7581 2038 7828 2072
rect 7862 2038 7900 2072
rect 7934 2038 8181 2072
rect 7581 1999 8181 2038
rect 7581 1965 7828 1999
rect 7862 1965 7900 1999
rect 7934 1965 8181 1999
rect 7581 1926 8181 1965
rect 7581 1892 7828 1926
rect 7862 1892 7900 1926
rect 7934 1892 8181 1926
rect 7581 1853 8181 1892
rect 7581 1819 7828 1853
rect 7862 1819 7900 1853
rect 7934 1819 8181 1853
rect 7581 1780 8181 1819
rect 7581 1746 7828 1780
rect 7862 1746 7900 1780
rect 7934 1746 8181 1780
rect 7581 1707 8181 1746
rect 7581 1673 7828 1707
rect 7862 1673 7900 1707
rect 7934 1673 8181 1707
rect 7581 1634 8181 1673
rect 7581 1600 7828 1634
rect 7862 1600 7900 1634
rect 7934 1600 8181 1634
rect 7581 1561 8181 1600
rect 7581 1527 7828 1561
rect 7862 1527 7900 1561
rect 7934 1527 8181 1561
rect 7581 1488 8181 1527
rect 7581 1454 7828 1488
rect 7862 1454 7900 1488
rect 7934 1454 8181 1488
rect 7581 1415 8181 1454
rect 7581 1381 7828 1415
rect 7862 1381 7900 1415
rect 7934 1381 8181 1415
rect 7581 1342 8181 1381
rect 7581 1308 7828 1342
rect 7862 1308 7900 1342
rect 7934 1308 8181 1342
rect 7581 1269 8181 1308
rect 7581 1235 7828 1269
rect 7862 1235 7900 1269
rect 7934 1235 8181 1269
rect 7581 1135 8181 1235
tri 7581 1131 7585 1135 ne
rect 7585 1131 8177 1135
tri 8177 1131 8181 1135 nw
tri 8483 11333 8530 11380 se
rect 8530 11333 9036 11380
tri 9036 11333 9083 11380 sw
rect 8483 11233 9083 11333
rect 8483 3279 8730 11233
rect 8836 3279 9083 11233
rect 8483 3240 9083 3279
rect 8483 3206 8730 3240
rect 8764 3206 8802 3240
rect 8836 3206 9083 3240
rect 8483 3167 9083 3206
rect 8483 3133 8730 3167
rect 8764 3133 8802 3167
rect 8836 3133 9083 3167
rect 8483 3094 9083 3133
rect 8483 3060 8730 3094
rect 8764 3060 8802 3094
rect 8836 3060 9083 3094
rect 8483 3021 9083 3060
rect 8483 2987 8730 3021
rect 8764 2987 8802 3021
rect 8836 2987 9083 3021
rect 8483 2948 9083 2987
rect 8483 2914 8730 2948
rect 8764 2914 8802 2948
rect 8836 2914 9083 2948
rect 8483 2875 9083 2914
rect 8483 2841 8730 2875
rect 8764 2841 8802 2875
rect 8836 2841 9083 2875
rect 8483 2802 9083 2841
rect 8483 2768 8730 2802
rect 8764 2768 8802 2802
rect 8836 2768 9083 2802
rect 8483 2729 9083 2768
rect 8483 2695 8730 2729
rect 8764 2695 8802 2729
rect 8836 2695 9083 2729
rect 8483 2656 9083 2695
rect 8483 2622 8730 2656
rect 8764 2622 8802 2656
rect 8836 2622 9083 2656
rect 8483 2583 9083 2622
rect 8483 2549 8730 2583
rect 8764 2549 8802 2583
rect 8836 2549 9083 2583
rect 8483 2510 9083 2549
rect 8483 2476 8730 2510
rect 8764 2476 8802 2510
rect 8836 2476 9083 2510
rect 8483 2437 9083 2476
rect 8483 2403 8730 2437
rect 8764 2403 8802 2437
rect 8836 2403 9083 2437
rect 8483 2364 9083 2403
rect 8483 2330 8730 2364
rect 8764 2330 8802 2364
rect 8836 2330 9083 2364
rect 8483 2291 9083 2330
rect 8483 2257 8730 2291
rect 8764 2257 8802 2291
rect 8836 2257 9083 2291
rect 8483 2218 9083 2257
rect 8483 2184 8730 2218
rect 8764 2184 8802 2218
rect 8836 2184 9083 2218
rect 8483 2145 9083 2184
rect 8483 2111 8730 2145
rect 8764 2111 8802 2145
rect 8836 2111 9083 2145
rect 8483 2072 9083 2111
rect 8483 2038 8730 2072
rect 8764 2038 8802 2072
rect 8836 2038 9083 2072
rect 8483 1999 9083 2038
rect 8483 1965 8730 1999
rect 8764 1965 8802 1999
rect 8836 1965 9083 1999
rect 8483 1926 9083 1965
rect 8483 1892 8730 1926
rect 8764 1892 8802 1926
rect 8836 1892 9083 1926
rect 8483 1853 9083 1892
rect 8483 1819 8730 1853
rect 8764 1819 8802 1853
rect 8836 1819 9083 1853
rect 8483 1780 9083 1819
rect 8483 1746 8730 1780
rect 8764 1746 8802 1780
rect 8836 1746 9083 1780
rect 8483 1707 9083 1746
rect 8483 1673 8730 1707
rect 8764 1673 8802 1707
rect 8836 1673 9083 1707
rect 8483 1634 9083 1673
rect 8483 1600 8730 1634
rect 8764 1600 8802 1634
rect 8836 1600 9083 1634
rect 8483 1561 9083 1600
rect 8483 1527 8730 1561
rect 8764 1527 8802 1561
rect 8836 1527 9083 1561
rect 8483 1488 9083 1527
rect 8483 1454 8730 1488
rect 8764 1454 8802 1488
rect 8836 1454 9083 1488
rect 8483 1415 9083 1454
rect 8483 1381 8730 1415
rect 8764 1381 8802 1415
rect 8836 1381 9083 1415
rect 8483 1342 9083 1381
rect 8483 1308 8730 1342
rect 8764 1308 8802 1342
rect 8836 1308 9083 1342
rect 8483 1269 9083 1308
rect 8483 1235 8730 1269
rect 8764 1235 8802 1269
rect 8836 1235 9083 1269
rect 8483 1135 9083 1235
tri 8483 1131 8487 1135 ne
rect 8487 1131 9079 1135
tri 9079 1131 9083 1135 nw
tri 9385 11333 9432 11380 se
rect 9432 11333 9938 11380
tri 9938 11333 9985 11380 sw
rect 9385 11233 9985 11333
rect 9385 3279 9632 11233
rect 9738 3279 9985 11233
rect 9385 3240 9985 3279
rect 9385 3206 9632 3240
rect 9666 3206 9704 3240
rect 9738 3206 9985 3240
rect 9385 3167 9985 3206
rect 9385 3133 9632 3167
rect 9666 3133 9704 3167
rect 9738 3133 9985 3167
rect 9385 3094 9985 3133
rect 9385 3060 9632 3094
rect 9666 3060 9704 3094
rect 9738 3060 9985 3094
rect 9385 3021 9985 3060
rect 9385 2987 9632 3021
rect 9666 2987 9704 3021
rect 9738 2987 9985 3021
rect 9385 2948 9985 2987
rect 9385 2914 9632 2948
rect 9666 2914 9704 2948
rect 9738 2914 9985 2948
rect 9385 2875 9985 2914
rect 9385 2841 9632 2875
rect 9666 2841 9704 2875
rect 9738 2841 9985 2875
rect 9385 2802 9985 2841
rect 9385 2768 9632 2802
rect 9666 2768 9704 2802
rect 9738 2768 9985 2802
rect 9385 2729 9985 2768
rect 9385 2695 9632 2729
rect 9666 2695 9704 2729
rect 9738 2695 9985 2729
rect 9385 2656 9985 2695
rect 9385 2622 9632 2656
rect 9666 2622 9704 2656
rect 9738 2622 9985 2656
rect 9385 2583 9985 2622
rect 9385 2549 9632 2583
rect 9666 2549 9704 2583
rect 9738 2549 9985 2583
rect 9385 2510 9985 2549
rect 9385 2476 9632 2510
rect 9666 2476 9704 2510
rect 9738 2476 9985 2510
rect 9385 2437 9985 2476
rect 9385 2403 9632 2437
rect 9666 2403 9704 2437
rect 9738 2403 9985 2437
rect 9385 2364 9985 2403
rect 9385 2330 9632 2364
rect 9666 2330 9704 2364
rect 9738 2330 9985 2364
rect 9385 2291 9985 2330
rect 9385 2257 9632 2291
rect 9666 2257 9704 2291
rect 9738 2257 9985 2291
rect 9385 2218 9985 2257
rect 9385 2184 9632 2218
rect 9666 2184 9704 2218
rect 9738 2184 9985 2218
rect 9385 2145 9985 2184
rect 9385 2111 9632 2145
rect 9666 2111 9704 2145
rect 9738 2111 9985 2145
rect 9385 2072 9985 2111
rect 9385 2038 9632 2072
rect 9666 2038 9704 2072
rect 9738 2038 9985 2072
rect 9385 1999 9985 2038
rect 9385 1965 9632 1999
rect 9666 1965 9704 1999
rect 9738 1965 9985 1999
rect 9385 1926 9985 1965
rect 9385 1892 9632 1926
rect 9666 1892 9704 1926
rect 9738 1892 9985 1926
rect 9385 1853 9985 1892
rect 9385 1819 9632 1853
rect 9666 1819 9704 1853
rect 9738 1819 9985 1853
rect 9385 1780 9985 1819
rect 9385 1746 9632 1780
rect 9666 1746 9704 1780
rect 9738 1746 9985 1780
rect 9385 1707 9985 1746
rect 9385 1673 9632 1707
rect 9666 1673 9704 1707
rect 9738 1673 9985 1707
rect 9385 1634 9985 1673
rect 9385 1600 9632 1634
rect 9666 1600 9704 1634
rect 9738 1600 9985 1634
rect 9385 1561 9985 1600
rect 9385 1527 9632 1561
rect 9666 1527 9704 1561
rect 9738 1527 9985 1561
rect 9385 1488 9985 1527
rect 9385 1454 9632 1488
rect 9666 1454 9704 1488
rect 9738 1454 9985 1488
rect 9385 1415 9985 1454
rect 9385 1381 9632 1415
rect 9666 1381 9704 1415
rect 9738 1381 9985 1415
rect 9385 1342 9985 1381
rect 9385 1308 9632 1342
rect 9666 1308 9704 1342
rect 9738 1308 9985 1342
rect 9385 1269 9985 1308
rect 9385 1235 9632 1269
rect 9666 1235 9704 1269
rect 9738 1235 9985 1269
rect 9385 1135 9985 1235
tri 9385 1131 9389 1135 ne
rect 9389 1131 9981 1135
tri 9981 1131 9985 1135 nw
tri 10287 11333 10334 11380 se
rect 10334 11333 10840 11380
tri 10840 11333 10887 11380 sw
rect 10287 11233 10887 11333
rect 10287 3279 10534 11233
rect 10640 3279 10887 11233
rect 10287 3240 10887 3279
rect 10287 3206 10534 3240
rect 10568 3206 10606 3240
rect 10640 3206 10887 3240
rect 10287 3167 10887 3206
rect 10287 3133 10534 3167
rect 10568 3133 10606 3167
rect 10640 3133 10887 3167
rect 10287 3094 10887 3133
rect 10287 3060 10534 3094
rect 10568 3060 10606 3094
rect 10640 3060 10887 3094
rect 10287 3021 10887 3060
rect 10287 2987 10534 3021
rect 10568 2987 10606 3021
rect 10640 2987 10887 3021
rect 10287 2948 10887 2987
rect 10287 2914 10534 2948
rect 10568 2914 10606 2948
rect 10640 2914 10887 2948
rect 10287 2875 10887 2914
rect 10287 2841 10534 2875
rect 10568 2841 10606 2875
rect 10640 2841 10887 2875
rect 10287 2802 10887 2841
rect 10287 2768 10534 2802
rect 10568 2768 10606 2802
rect 10640 2768 10887 2802
rect 10287 2729 10887 2768
rect 10287 2695 10534 2729
rect 10568 2695 10606 2729
rect 10640 2695 10887 2729
rect 10287 2656 10887 2695
rect 10287 2622 10534 2656
rect 10568 2622 10606 2656
rect 10640 2622 10887 2656
rect 10287 2583 10887 2622
rect 10287 2549 10534 2583
rect 10568 2549 10606 2583
rect 10640 2549 10887 2583
rect 10287 2510 10887 2549
rect 10287 2476 10534 2510
rect 10568 2476 10606 2510
rect 10640 2476 10887 2510
rect 10287 2437 10887 2476
rect 10287 2403 10534 2437
rect 10568 2403 10606 2437
rect 10640 2403 10887 2437
rect 10287 2364 10887 2403
rect 10287 2330 10534 2364
rect 10568 2330 10606 2364
rect 10640 2330 10887 2364
rect 10287 2291 10887 2330
rect 10287 2257 10534 2291
rect 10568 2257 10606 2291
rect 10640 2257 10887 2291
rect 10287 2218 10887 2257
rect 10287 2184 10534 2218
rect 10568 2184 10606 2218
rect 10640 2184 10887 2218
rect 10287 2145 10887 2184
rect 10287 2111 10534 2145
rect 10568 2111 10606 2145
rect 10640 2111 10887 2145
rect 10287 2072 10887 2111
rect 10287 2038 10534 2072
rect 10568 2038 10606 2072
rect 10640 2038 10887 2072
rect 10287 1999 10887 2038
rect 10287 1965 10534 1999
rect 10568 1965 10606 1999
rect 10640 1965 10887 1999
rect 10287 1926 10887 1965
rect 10287 1892 10534 1926
rect 10568 1892 10606 1926
rect 10640 1892 10887 1926
rect 10287 1853 10887 1892
rect 10287 1819 10534 1853
rect 10568 1819 10606 1853
rect 10640 1819 10887 1853
rect 10287 1780 10887 1819
rect 10287 1746 10534 1780
rect 10568 1746 10606 1780
rect 10640 1746 10887 1780
rect 10287 1707 10887 1746
rect 10287 1673 10534 1707
rect 10568 1673 10606 1707
rect 10640 1673 10887 1707
rect 10287 1634 10887 1673
rect 10287 1600 10534 1634
rect 10568 1600 10606 1634
rect 10640 1600 10887 1634
rect 10287 1561 10887 1600
rect 10287 1527 10534 1561
rect 10568 1527 10606 1561
rect 10640 1527 10887 1561
rect 10287 1488 10887 1527
rect 10287 1454 10534 1488
rect 10568 1454 10606 1488
rect 10640 1454 10887 1488
rect 10287 1415 10887 1454
rect 10287 1381 10534 1415
rect 10568 1381 10606 1415
rect 10640 1381 10887 1415
rect 10287 1342 10887 1381
rect 10287 1308 10534 1342
rect 10568 1308 10606 1342
rect 10640 1308 10887 1342
rect 10287 1269 10887 1308
rect 10287 1235 10534 1269
rect 10568 1235 10606 1269
rect 10640 1235 10887 1269
rect 10287 1135 10887 1235
tri 10287 1131 10291 1135 ne
rect 10291 1131 10883 1135
tri 10883 1131 10887 1135 nw
tri 11189 11333 11236 11380 se
rect 11236 11333 11742 11380
tri 11742 11333 11789 11380 sw
rect 11189 11233 11789 11333
rect 11189 3279 11436 11233
rect 11542 3279 11789 11233
rect 11189 3240 11789 3279
rect 11189 3206 11436 3240
rect 11470 3206 11508 3240
rect 11542 3206 11789 3240
rect 11189 3167 11789 3206
rect 11189 3133 11436 3167
rect 11470 3133 11508 3167
rect 11542 3133 11789 3167
rect 11189 3094 11789 3133
rect 11189 3060 11436 3094
rect 11470 3060 11508 3094
rect 11542 3060 11789 3094
rect 11189 3021 11789 3060
rect 11189 2987 11436 3021
rect 11470 2987 11508 3021
rect 11542 2987 11789 3021
rect 11189 2948 11789 2987
rect 11189 2914 11436 2948
rect 11470 2914 11508 2948
rect 11542 2914 11789 2948
rect 11189 2875 11789 2914
rect 11189 2841 11436 2875
rect 11470 2841 11508 2875
rect 11542 2841 11789 2875
rect 11189 2802 11789 2841
rect 11189 2768 11436 2802
rect 11470 2768 11508 2802
rect 11542 2768 11789 2802
rect 11189 2729 11789 2768
rect 11189 2695 11436 2729
rect 11470 2695 11508 2729
rect 11542 2695 11789 2729
rect 11189 2656 11789 2695
rect 11189 2622 11436 2656
rect 11470 2622 11508 2656
rect 11542 2622 11789 2656
rect 11189 2583 11789 2622
rect 11189 2549 11436 2583
rect 11470 2549 11508 2583
rect 11542 2549 11789 2583
rect 11189 2510 11789 2549
rect 11189 2476 11436 2510
rect 11470 2476 11508 2510
rect 11542 2476 11789 2510
rect 11189 2437 11789 2476
rect 11189 2403 11436 2437
rect 11470 2403 11508 2437
rect 11542 2403 11789 2437
rect 11189 2364 11789 2403
rect 11189 2330 11436 2364
rect 11470 2330 11508 2364
rect 11542 2330 11789 2364
rect 11189 2291 11789 2330
rect 11189 2257 11436 2291
rect 11470 2257 11508 2291
rect 11542 2257 11789 2291
rect 11189 2218 11789 2257
rect 11189 2184 11436 2218
rect 11470 2184 11508 2218
rect 11542 2184 11789 2218
rect 11189 2145 11789 2184
rect 11189 2111 11436 2145
rect 11470 2111 11508 2145
rect 11542 2111 11789 2145
rect 11189 2072 11789 2111
rect 11189 2038 11436 2072
rect 11470 2038 11508 2072
rect 11542 2038 11789 2072
rect 11189 1999 11789 2038
rect 11189 1965 11436 1999
rect 11470 1965 11508 1999
rect 11542 1965 11789 1999
rect 11189 1926 11789 1965
rect 11189 1892 11436 1926
rect 11470 1892 11508 1926
rect 11542 1892 11789 1926
rect 11189 1853 11789 1892
rect 11189 1819 11436 1853
rect 11470 1819 11508 1853
rect 11542 1819 11789 1853
rect 11189 1780 11789 1819
rect 11189 1746 11436 1780
rect 11470 1746 11508 1780
rect 11542 1746 11789 1780
rect 11189 1707 11789 1746
rect 11189 1673 11436 1707
rect 11470 1673 11508 1707
rect 11542 1673 11789 1707
rect 11189 1634 11789 1673
rect 11189 1600 11436 1634
rect 11470 1600 11508 1634
rect 11542 1600 11789 1634
rect 11189 1561 11789 1600
rect 11189 1527 11436 1561
rect 11470 1527 11508 1561
rect 11542 1527 11789 1561
rect 11189 1488 11789 1527
rect 11189 1454 11436 1488
rect 11470 1454 11508 1488
rect 11542 1454 11789 1488
rect 11189 1415 11789 1454
rect 11189 1381 11436 1415
rect 11470 1381 11508 1415
rect 11542 1381 11789 1415
rect 11189 1342 11789 1381
rect 11189 1308 11436 1342
rect 11470 1308 11508 1342
rect 11542 1308 11789 1342
rect 11189 1269 11789 1308
rect 11189 1235 11436 1269
rect 11470 1235 11508 1269
rect 11542 1235 11789 1269
rect 11189 1135 11789 1235
tri 11189 1131 11193 1135 ne
rect 11193 1131 11785 1135
tri 11785 1131 11789 1135 nw
tri 12091 11333 12138 11380 se
rect 12138 11333 12644 11380
tri 12644 11333 12691 11380 sw
rect 12091 11233 12691 11333
rect 12091 3279 12338 11233
rect 12444 3279 12691 11233
rect 12091 3240 12691 3279
rect 12091 3206 12338 3240
rect 12372 3206 12410 3240
rect 12444 3206 12691 3240
rect 12091 3167 12691 3206
rect 12091 3133 12338 3167
rect 12372 3133 12410 3167
rect 12444 3133 12691 3167
rect 12091 3094 12691 3133
rect 12091 3060 12338 3094
rect 12372 3060 12410 3094
rect 12444 3060 12691 3094
rect 12091 3021 12691 3060
rect 12091 2987 12338 3021
rect 12372 2987 12410 3021
rect 12444 2987 12691 3021
rect 12091 2948 12691 2987
rect 12091 2914 12338 2948
rect 12372 2914 12410 2948
rect 12444 2914 12691 2948
rect 12091 2875 12691 2914
rect 12091 2841 12338 2875
rect 12372 2841 12410 2875
rect 12444 2841 12691 2875
rect 12091 2802 12691 2841
rect 12091 2768 12338 2802
rect 12372 2768 12410 2802
rect 12444 2768 12691 2802
rect 12091 2729 12691 2768
rect 12091 2695 12338 2729
rect 12372 2695 12410 2729
rect 12444 2695 12691 2729
rect 12091 2656 12691 2695
rect 12091 2622 12338 2656
rect 12372 2622 12410 2656
rect 12444 2622 12691 2656
rect 12091 2583 12691 2622
rect 12091 2549 12338 2583
rect 12372 2549 12410 2583
rect 12444 2549 12691 2583
rect 12091 2510 12691 2549
rect 12091 2476 12338 2510
rect 12372 2476 12410 2510
rect 12444 2476 12691 2510
rect 12091 2437 12691 2476
rect 12091 2403 12338 2437
rect 12372 2403 12410 2437
rect 12444 2403 12691 2437
rect 12091 2364 12691 2403
rect 12091 2330 12338 2364
rect 12372 2330 12410 2364
rect 12444 2330 12691 2364
rect 12091 2291 12691 2330
rect 12091 2257 12338 2291
rect 12372 2257 12410 2291
rect 12444 2257 12691 2291
rect 12091 2218 12691 2257
rect 12091 2184 12338 2218
rect 12372 2184 12410 2218
rect 12444 2184 12691 2218
rect 12091 2145 12691 2184
rect 12091 2111 12338 2145
rect 12372 2111 12410 2145
rect 12444 2111 12691 2145
rect 12091 2072 12691 2111
rect 12091 2038 12338 2072
rect 12372 2038 12410 2072
rect 12444 2038 12691 2072
rect 12091 1999 12691 2038
rect 12091 1965 12338 1999
rect 12372 1965 12410 1999
rect 12444 1965 12691 1999
rect 12091 1926 12691 1965
rect 12091 1892 12338 1926
rect 12372 1892 12410 1926
rect 12444 1892 12691 1926
rect 12091 1853 12691 1892
rect 12091 1819 12338 1853
rect 12372 1819 12410 1853
rect 12444 1819 12691 1853
rect 12091 1780 12691 1819
rect 12091 1746 12338 1780
rect 12372 1746 12410 1780
rect 12444 1746 12691 1780
rect 12091 1707 12691 1746
rect 12091 1673 12338 1707
rect 12372 1673 12410 1707
rect 12444 1673 12691 1707
rect 12091 1634 12691 1673
rect 12091 1600 12338 1634
rect 12372 1600 12410 1634
rect 12444 1600 12691 1634
rect 12091 1561 12691 1600
rect 12091 1527 12338 1561
rect 12372 1527 12410 1561
rect 12444 1527 12691 1561
rect 12091 1488 12691 1527
rect 12091 1454 12338 1488
rect 12372 1454 12410 1488
rect 12444 1454 12691 1488
rect 12091 1415 12691 1454
rect 12091 1381 12338 1415
rect 12372 1381 12410 1415
rect 12444 1381 12691 1415
rect 12091 1342 12691 1381
rect 12091 1308 12338 1342
rect 12372 1308 12410 1342
rect 12444 1308 12691 1342
rect 12091 1269 12691 1308
rect 12091 1235 12338 1269
rect 12372 1235 12410 1269
rect 12444 1235 12691 1269
rect 12091 1135 12691 1235
tri 12091 1131 12095 1135 ne
rect 12095 1131 12687 1135
tri 12687 1131 12691 1135 nw
tri 12993 11333 13040 11380 se
rect 13040 11333 13546 11380
tri 13546 11333 13593 11380 sw
rect 12993 11233 13593 11333
rect 12993 3279 13240 11233
rect 13346 3279 13593 11233
rect 12993 3240 13593 3279
rect 12993 3206 13240 3240
rect 13274 3206 13312 3240
rect 13346 3206 13593 3240
rect 12993 3167 13593 3206
rect 12993 3133 13240 3167
rect 13274 3133 13312 3167
rect 13346 3133 13593 3167
rect 12993 3094 13593 3133
rect 12993 3060 13240 3094
rect 13274 3060 13312 3094
rect 13346 3060 13593 3094
rect 12993 3021 13593 3060
rect 12993 2987 13240 3021
rect 13274 2987 13312 3021
rect 13346 2987 13593 3021
rect 12993 2948 13593 2987
rect 12993 2914 13240 2948
rect 13274 2914 13312 2948
rect 13346 2914 13593 2948
rect 12993 2875 13593 2914
rect 12993 2841 13240 2875
rect 13274 2841 13312 2875
rect 13346 2841 13593 2875
rect 12993 2802 13593 2841
rect 12993 2768 13240 2802
rect 13274 2768 13312 2802
rect 13346 2768 13593 2802
rect 12993 2729 13593 2768
rect 12993 2695 13240 2729
rect 13274 2695 13312 2729
rect 13346 2695 13593 2729
rect 12993 2656 13593 2695
rect 12993 2622 13240 2656
rect 13274 2622 13312 2656
rect 13346 2622 13593 2656
rect 12993 2583 13593 2622
rect 12993 2549 13240 2583
rect 13274 2549 13312 2583
rect 13346 2549 13593 2583
rect 12993 2510 13593 2549
rect 12993 2476 13240 2510
rect 13274 2476 13312 2510
rect 13346 2476 13593 2510
rect 12993 2437 13593 2476
rect 12993 2403 13240 2437
rect 13274 2403 13312 2437
rect 13346 2403 13593 2437
rect 12993 2364 13593 2403
rect 12993 2330 13240 2364
rect 13274 2330 13312 2364
rect 13346 2330 13593 2364
rect 12993 2291 13593 2330
rect 12993 2257 13240 2291
rect 13274 2257 13312 2291
rect 13346 2257 13593 2291
rect 12993 2218 13593 2257
rect 12993 2184 13240 2218
rect 13274 2184 13312 2218
rect 13346 2184 13593 2218
rect 12993 2145 13593 2184
rect 12993 2111 13240 2145
rect 13274 2111 13312 2145
rect 13346 2111 13593 2145
rect 12993 2072 13593 2111
rect 12993 2038 13240 2072
rect 13274 2038 13312 2072
rect 13346 2038 13593 2072
rect 12993 1999 13593 2038
rect 12993 1965 13240 1999
rect 13274 1965 13312 1999
rect 13346 1965 13593 1999
rect 12993 1926 13593 1965
rect 12993 1892 13240 1926
rect 13274 1892 13312 1926
rect 13346 1892 13593 1926
rect 12993 1853 13593 1892
rect 12993 1819 13240 1853
rect 13274 1819 13312 1853
rect 13346 1819 13593 1853
rect 12993 1780 13593 1819
rect 12993 1746 13240 1780
rect 13274 1746 13312 1780
rect 13346 1746 13593 1780
rect 12993 1707 13593 1746
rect 12993 1673 13240 1707
rect 13274 1673 13312 1707
rect 13346 1673 13593 1707
rect 12993 1634 13593 1673
rect 12993 1600 13240 1634
rect 13274 1600 13312 1634
rect 13346 1600 13593 1634
rect 12993 1561 13593 1600
rect 12993 1527 13240 1561
rect 13274 1527 13312 1561
rect 13346 1527 13593 1561
rect 12993 1488 13593 1527
rect 12993 1454 13240 1488
rect 13274 1454 13312 1488
rect 13346 1454 13593 1488
rect 12993 1415 13593 1454
rect 12993 1381 13240 1415
rect 13274 1381 13312 1415
rect 13346 1381 13593 1415
rect 12993 1342 13593 1381
rect 12993 1308 13240 1342
rect 13274 1308 13312 1342
rect 13346 1308 13593 1342
rect 12993 1269 13593 1308
rect 12993 1235 13240 1269
rect 13274 1235 13312 1269
rect 13346 1235 13593 1269
rect 12993 1135 13593 1235
tri 12993 1131 12997 1135 ne
rect 12997 1131 13589 1135
tri 13589 1131 13593 1135 nw
tri 13895 11333 13896 11334 se
rect 13896 11333 14766 11483
rect 13895 11233 14766 11333
rect 13895 3279 14142 11233
rect 14248 3279 14766 11233
rect 13895 3240 14766 3279
rect 13895 3206 14142 3240
rect 14176 3206 14214 3240
rect 14248 3206 14766 3240
rect 13895 3167 14766 3206
rect 13895 3133 14142 3167
rect 14176 3133 14214 3167
rect 14248 3133 14766 3167
rect 13895 3094 14766 3133
rect 13895 3060 14142 3094
rect 14176 3060 14214 3094
rect 14248 3060 14766 3094
rect 13895 3021 14766 3060
rect 13895 2987 14142 3021
rect 14176 2987 14214 3021
rect 14248 2987 14766 3021
rect 13895 2948 14766 2987
rect 13895 2914 14142 2948
rect 14176 2914 14214 2948
rect 14248 2914 14766 2948
rect 13895 2875 14766 2914
rect 13895 2841 14142 2875
rect 14176 2841 14214 2875
rect 14248 2841 14766 2875
rect 13895 2802 14766 2841
rect 13895 2768 14142 2802
rect 14176 2768 14214 2802
rect 14248 2768 14766 2802
rect 13895 2729 14766 2768
rect 13895 2695 14142 2729
rect 14176 2695 14214 2729
rect 14248 2695 14766 2729
rect 13895 2656 14766 2695
rect 13895 2622 14142 2656
rect 14176 2622 14214 2656
rect 14248 2622 14766 2656
rect 13895 2583 14766 2622
rect 13895 2549 14142 2583
rect 14176 2549 14214 2583
rect 14248 2549 14766 2583
rect 13895 2510 14766 2549
rect 13895 2476 14142 2510
rect 14176 2476 14214 2510
rect 14248 2476 14766 2510
rect 13895 2437 14766 2476
rect 13895 2403 14142 2437
rect 14176 2403 14214 2437
rect 14248 2403 14766 2437
rect 13895 2364 14766 2403
rect 13895 2330 14142 2364
rect 14176 2330 14214 2364
rect 14248 2330 14766 2364
rect 13895 2291 14766 2330
rect 13895 2257 14142 2291
rect 14176 2257 14214 2291
rect 14248 2257 14766 2291
rect 13895 2218 14766 2257
rect 13895 2184 14142 2218
rect 14176 2184 14214 2218
rect 14248 2184 14766 2218
rect 13895 2145 14766 2184
rect 13895 2111 14142 2145
rect 14176 2111 14214 2145
rect 14248 2111 14766 2145
rect 13895 2072 14766 2111
rect 13895 2038 14142 2072
rect 14176 2038 14214 2072
rect 14248 2038 14766 2072
rect 13895 1999 14766 2038
rect 13895 1965 14142 1999
rect 14176 1965 14214 1999
rect 14248 1965 14766 1999
rect 13895 1926 14766 1965
rect 13895 1892 14142 1926
rect 14176 1892 14214 1926
rect 14248 1892 14766 1926
rect 13895 1853 14766 1892
rect 13895 1819 14142 1853
rect 14176 1819 14214 1853
rect 14248 1819 14766 1853
rect 13895 1780 14766 1819
rect 13895 1746 14142 1780
rect 14176 1746 14214 1780
rect 14248 1746 14766 1780
rect 13895 1707 14766 1746
rect 13895 1673 14142 1707
rect 14176 1673 14214 1707
rect 14248 1673 14766 1707
rect 13895 1634 14766 1673
rect 13895 1600 14142 1634
rect 14176 1600 14214 1634
rect 14248 1600 14766 1634
rect 13895 1561 14766 1600
rect 13895 1527 14142 1561
rect 14176 1527 14214 1561
rect 14248 1527 14766 1561
rect 13895 1488 14766 1527
rect 13895 1454 14142 1488
rect 14176 1454 14214 1488
rect 14248 1454 14766 1488
rect 13895 1415 14766 1454
rect 13895 1381 14142 1415
rect 14176 1381 14214 1415
rect 14248 1381 14766 1415
rect 13895 1342 14766 1381
rect 13895 1308 14142 1342
rect 14176 1308 14214 1342
rect 14248 1308 14766 1342
rect 13895 1269 14766 1308
rect 13895 1235 14142 1269
rect 14176 1235 14214 1269
rect 14248 1235 14766 1269
rect 13895 1135 14766 1235
tri 13895 1134 13896 1135 ne
rect 13896 1134 14766 1135
tri 13896 1131 13899 1134 ne
rect 13899 1131 14766 1134
tri -4141 1097 -4107 1131 ne
rect -4107 1097 -3583 1131
tri -3583 1097 -3549 1131 nw
tri -3239 1097 -3205 1131 ne
rect -3205 1097 -2681 1131
tri -2681 1097 -2647 1131 nw
tri -2337 1097 -2303 1131 ne
rect -2303 1097 -1779 1131
tri -1779 1097 -1745 1131 nw
tri -1435 1097 -1401 1131 ne
rect -1401 1097 -877 1131
tri -877 1097 -843 1131 nw
tri -533 1097 -499 1131 ne
rect -499 1097 25 1131
tri 25 1097 59 1131 nw
tri 369 1097 403 1131 ne
rect 403 1097 927 1131
tri 927 1097 961 1131 nw
tri 1271 1097 1305 1131 ne
rect 1305 1097 1829 1131
tri 1829 1097 1863 1131 nw
tri 2173 1097 2207 1131 ne
rect 2207 1097 2731 1131
tri 2731 1097 2765 1131 nw
tri 3075 1097 3109 1131 ne
rect 3109 1097 3633 1131
tri 3633 1097 3667 1131 nw
tri 3977 1097 4011 1131 ne
rect 4011 1097 4535 1131
tri 4535 1097 4569 1131 nw
tri 4879 1097 4913 1131 ne
rect 4913 1097 5437 1131
tri 5437 1097 5471 1131 nw
tri 5781 1097 5815 1131 ne
rect 5815 1097 6339 1131
tri 6339 1097 6373 1131 nw
tri 6683 1097 6717 1131 ne
rect 6717 1097 7241 1131
tri 7241 1097 7275 1131 nw
tri 7585 1097 7619 1131 ne
rect 7619 1097 8143 1131
tri 8143 1097 8177 1131 nw
tri 8487 1097 8521 1131 ne
rect 8521 1097 9045 1131
tri 9045 1097 9079 1131 nw
tri 9389 1097 9423 1131 ne
rect 9423 1097 9947 1131
tri 9947 1097 9981 1131 nw
tri 10291 1097 10325 1131 ne
rect 10325 1097 10849 1131
tri 10849 1097 10883 1131 nw
tri 11193 1097 11227 1131 ne
rect 11227 1097 11751 1131
tri 11751 1097 11785 1131 nw
tri 12095 1097 12129 1131 ne
rect 12129 1097 12653 1131
tri 12653 1097 12687 1131 nw
tri 12997 1097 13031 1131 ne
rect 13031 1097 13555 1131
tri 13555 1097 13589 1131 nw
tri 13899 1127 13903 1131 ne
rect 13903 1127 14766 1131
tri 13903 1120 13910 1127 ne
rect 13910 1120 14766 1127
tri 13910 1113 13917 1120 ne
rect 13917 1113 14766 1120
tri 13917 1109 13921 1113 ne
rect 13921 1109 14766 1113
tri 13921 1102 13928 1109 ne
rect 13928 1102 14766 1109
tri 13928 1097 13933 1102 ne
rect 13933 1097 14766 1102
tri -4107 1088 -4098 1097 ne
rect -4098 1088 -3592 1097
tri -3592 1088 -3583 1097 nw
tri -3205 1088 -3196 1097 ne
rect -3196 1088 -2690 1097
tri -2690 1088 -2681 1097 nw
tri -2303 1088 -2294 1097 ne
rect -2294 1088 -1788 1097
tri -1788 1088 -1779 1097 nw
tri -1401 1088 -1392 1097 ne
rect -1392 1088 -886 1097
tri -886 1088 -877 1097 nw
tri -499 1088 -490 1097 ne
rect -490 1088 16 1097
tri 16 1088 25 1097 nw
tri 403 1088 412 1097 ne
rect 412 1088 918 1097
tri 918 1088 927 1097 nw
tri 1305 1088 1314 1097 ne
rect 1314 1088 1820 1097
tri 1820 1088 1829 1097 nw
tri 2207 1088 2216 1097 ne
rect 2216 1088 2722 1097
tri 2722 1088 2731 1097 nw
tri 3109 1088 3118 1097 ne
rect 3118 1088 3624 1097
tri 3624 1088 3633 1097 nw
tri 4011 1088 4020 1097 ne
rect 4020 1088 4526 1097
tri 4526 1088 4535 1097 nw
tri 4913 1088 4922 1097 ne
rect 4922 1088 5428 1097
tri 5428 1088 5437 1097 nw
tri 5815 1088 5824 1097 ne
rect 5824 1088 6330 1097
tri 6330 1088 6339 1097 nw
tri 6717 1088 6726 1097 ne
rect 6726 1088 7232 1097
tri 7232 1088 7241 1097 nw
tri 7619 1088 7628 1097 ne
rect 7628 1088 8134 1097
tri 8134 1088 8143 1097 nw
tri 8521 1088 8530 1097 ne
rect 8530 1088 9036 1097
tri 9036 1088 9045 1097 nw
tri 9423 1088 9432 1097 ne
rect 9432 1088 9938 1097
tri 9938 1088 9947 1097 nw
tri 10325 1088 10334 1097 ne
rect 10334 1088 10840 1097
tri 10840 1088 10849 1097 nw
tri 11227 1088 11236 1097 ne
rect 11236 1088 11742 1097
tri 11742 1088 11751 1097 nw
tri 12129 1088 12138 1097 ne
rect 12138 1088 12644 1097
tri 12644 1088 12653 1097 nw
tri 13031 1088 13040 1097 ne
rect 13040 1088 13546 1097
tri 13546 1088 13555 1097 nw
tri 13933 1095 13935 1097 ne
rect 13935 1095 14766 1097
tri 13935 1088 13942 1095 ne
rect 13942 1088 14766 1095
tri 14587 1058 14617 1088 ne
rect 14617 1058 14766 1088
tri 14617 1054 14621 1058 ne
rect 14621 1054 14766 1058
rect -2364 1050 -2234 1054
rect -2364 1042 -2232 1050
rect -3656 1020 -3443 1032
rect -3656 986 -3644 1020
rect -3610 986 -3572 1020
rect -3538 986 -3443 1020
rect -2364 1008 -2352 1042
rect -2318 1008 -2280 1042
rect -2246 1008 -2232 1042
rect -2364 996 -2232 1008
rect -1852 1042 -1722 1054
rect -1852 1008 -1840 1042
rect -1806 1008 -1768 1042
rect -1734 1008 -1722 1042
rect -1852 996 -1722 1008
rect -560 1050 -430 1054
rect -560 1042 -428 1050
rect -560 1008 -548 1042
rect -514 1008 -476 1042
rect -442 1008 -428 1042
rect -560 996 -428 1008
rect -48 1042 82 1054
rect -48 1008 -36 1042
rect -2 1008 36 1042
rect 70 1008 82 1042
rect -48 996 82 1008
rect 1244 1050 1374 1054
rect 1244 1042 1378 1050
rect 1244 1008 1256 1042
rect 1290 1008 1328 1042
rect 1362 1008 1378 1042
rect 1244 996 1378 1008
rect 1756 1042 1886 1054
rect 1756 1008 1768 1042
rect 1802 1008 1840 1042
rect 1874 1008 1886 1042
rect 1756 996 1886 1008
rect 3048 1042 3178 1054
rect 3048 1008 3060 1042
rect 3094 1008 3132 1042
rect 3166 1008 3178 1042
rect 3048 996 3178 1008
rect 3560 1042 3690 1054
rect 3560 1008 3572 1042
rect 3606 1008 3644 1042
rect 3678 1008 3690 1042
rect 3560 996 3690 1008
rect 4852 1050 4982 1054
rect 4852 1042 4984 1050
rect 4852 1008 4864 1042
rect 4898 1008 4936 1042
rect 4970 1008 4984 1042
rect 4852 996 4984 1008
rect 5364 1042 5494 1054
rect 5364 1008 5376 1042
rect 5410 1008 5448 1042
rect 5482 1008 5494 1042
rect 5364 996 5494 1008
rect 6656 1042 6786 1054
rect 6656 1008 6668 1042
rect 6702 1008 6740 1042
rect 6774 1008 6786 1042
rect 6656 996 6786 1008
rect 7168 1042 7298 1054
rect 7168 1008 7180 1042
rect 7214 1008 7252 1042
rect 7286 1008 7298 1042
rect 7168 996 7298 1008
rect 8460 1042 8590 1054
rect 8460 1008 8472 1042
rect 8506 1008 8544 1042
rect 8578 1008 8590 1042
rect 8460 996 8590 1008
rect 8972 1042 9102 1054
rect 8972 1008 8984 1042
rect 9018 1008 9056 1042
rect 9090 1008 9102 1042
rect 8972 996 9102 1008
rect 10264 1042 10394 1054
rect 10264 1008 10276 1042
rect 10310 1008 10348 1042
rect 10382 1008 10394 1042
rect 10264 996 10394 1008
rect 10776 1042 10906 1054
rect 10776 1008 10788 1042
rect 10822 1008 10860 1042
rect 10894 1008 10906 1042
rect 10776 996 10906 1008
rect 12068 1042 12198 1054
rect 12068 1008 12080 1042
rect 12114 1008 12152 1042
rect 12186 1008 12198 1042
rect 12068 996 12198 1008
rect 12580 1042 12710 1054
rect 12580 1008 12592 1042
rect 12626 1008 12664 1042
rect 12698 1008 12710 1042
tri 14621 1039 14636 1054 ne
rect 12580 996 12710 1008
rect 13872 1020 14002 1032
rect -2290 992 -2232 996
rect -1831 992 -1779 996
rect -486 992 -428 996
rect -28 992 28 996
rect 1319 992 1378 996
rect 1778 992 1833 996
rect 3124 992 3177 996
rect 3579 992 3636 996
rect 4929 992 4984 996
rect -3656 974 -3443 986
rect 13872 986 13884 1020
rect 13918 986 13956 1020
rect 13990 986 14002 1020
rect 13872 974 14002 986
tri -4286 693 -4262 717 sw
tri 14624 693 14636 705 se
rect 14636 693 14766 1054
rect -4416 659 -4262 693
tri -4262 659 -4228 693 sw
tri 14590 659 14624 693 se
rect 14624 659 14766 693
rect -4416 620 -4228 659
tri -4228 620 -4189 659 sw
tri 14551 620 14590 659 se
rect 14590 620 14766 659
tri -4416 608 -4404 620 ne
rect -4404 608 -1663 620
rect -4965 547 -4770 586
tri -4404 574 -4370 608 ne
rect -4370 574 -4313 608
rect -4279 574 -1663 608
tri -4370 562 -4358 574 ne
rect -4358 562 -1663 574
tri -4358 547 -4343 562 ne
rect -4343 547 -1663 562
rect -4965 513 -4888 547
rect -4854 513 -4816 547
rect -4782 513 -4770 547
tri -4343 513 -4309 547 ne
rect -4309 513 -1663 547
rect -4965 474 -4770 513
tri -4309 490 -4286 513 ne
rect -4286 490 -1663 513
rect 13896 608 14732 620
rect 13896 574 14603 608
rect 14637 586 14732 608
tri 14732 586 14766 620 nw
rect 15120 11611 15132 11861
rect 15238 11611 15315 11861
rect 15120 11562 15315 11611
rect 15120 11528 15132 11562
rect 15166 11528 15204 11562
rect 15238 11528 15315 11562
rect 15120 11483 15315 11528
rect 15120 5185 15132 11483
rect 15238 5185 15315 11483
rect 15120 5146 15315 5185
rect 15120 5112 15132 5146
rect 15166 5112 15204 5146
rect 15238 5112 15315 5146
rect 15120 5073 15315 5112
rect 15120 5039 15132 5073
rect 15166 5039 15204 5073
rect 15238 5039 15315 5073
rect 15120 5000 15315 5039
rect 15120 4966 15132 5000
rect 15166 4966 15204 5000
rect 15238 4966 15315 5000
rect 15120 4927 15315 4966
rect 15120 4893 15132 4927
rect 15166 4893 15204 4927
rect 15238 4893 15315 4927
rect 15120 4854 15315 4893
rect 15120 4820 15132 4854
rect 15166 4820 15204 4854
rect 15238 4820 15315 4854
rect 15120 4781 15315 4820
rect 15120 4747 15132 4781
rect 15166 4747 15204 4781
rect 15238 4747 15315 4781
rect 15120 4708 15315 4747
rect 15120 4674 15132 4708
rect 15166 4674 15204 4708
rect 15238 4674 15315 4708
rect 15120 4635 15315 4674
rect 15120 4601 15132 4635
rect 15166 4601 15204 4635
rect 15238 4601 15315 4635
rect 15120 4562 15315 4601
rect 15120 4528 15132 4562
rect 15166 4528 15204 4562
rect 15238 4528 15315 4562
rect 15120 4489 15315 4528
rect 15120 4455 15132 4489
rect 15166 4455 15204 4489
rect 15238 4455 15315 4489
rect 15120 4416 15315 4455
rect 15120 4382 15132 4416
rect 15166 4382 15204 4416
rect 15238 4382 15315 4416
rect 15120 4343 15315 4382
rect 15120 4309 15132 4343
rect 15166 4309 15204 4343
rect 15238 4309 15315 4343
rect 15120 4270 15315 4309
rect 15120 4236 15132 4270
rect 15166 4236 15204 4270
rect 15238 4236 15315 4270
rect 15120 4197 15315 4236
rect 15120 4163 15132 4197
rect 15166 4163 15204 4197
rect 15238 4163 15315 4197
rect 15120 4124 15315 4163
rect 15120 4090 15132 4124
rect 15166 4090 15204 4124
rect 15238 4090 15315 4124
rect 15120 4051 15315 4090
rect 15120 4017 15132 4051
rect 15166 4017 15204 4051
rect 15238 4017 15315 4051
rect 15120 3978 15315 4017
rect 15120 3944 15132 3978
rect 15166 3944 15204 3978
rect 15238 3944 15315 3978
rect 15120 3905 15315 3944
rect 15120 3871 15132 3905
rect 15166 3871 15204 3905
rect 15238 3871 15315 3905
rect 15120 3832 15315 3871
rect 15120 3798 15132 3832
rect 15166 3798 15204 3832
rect 15238 3798 15315 3832
rect 15120 3759 15315 3798
rect 15120 3725 15132 3759
rect 15166 3725 15204 3759
rect 15238 3725 15315 3759
rect 15120 3686 15315 3725
rect 15120 3652 15132 3686
rect 15166 3652 15204 3686
rect 15238 3652 15315 3686
rect 15120 3613 15315 3652
rect 15120 3579 15132 3613
rect 15166 3579 15204 3613
rect 15238 3579 15315 3613
rect 15120 3540 15315 3579
rect 15120 3506 15132 3540
rect 15166 3506 15204 3540
rect 15238 3506 15315 3540
rect 15120 3467 15315 3506
rect 15120 3433 15132 3467
rect 15166 3433 15204 3467
rect 15238 3433 15315 3467
rect 15120 3394 15315 3433
rect 15120 3360 15132 3394
rect 15166 3360 15204 3394
rect 15238 3360 15315 3394
rect 15120 3321 15315 3360
rect 15120 3287 15132 3321
rect 15166 3287 15204 3321
rect 15238 3287 15315 3321
rect 15120 3248 15315 3287
rect 15120 3214 15132 3248
rect 15166 3214 15204 3248
rect 15238 3214 15315 3248
rect 15120 3175 15315 3214
rect 15120 3141 15132 3175
rect 15166 3141 15204 3175
rect 15238 3141 15315 3175
rect 15120 3102 15315 3141
rect 15120 3068 15132 3102
rect 15166 3068 15204 3102
rect 15238 3068 15315 3102
rect 15120 3029 15315 3068
rect 15120 2995 15132 3029
rect 15166 2995 15204 3029
rect 15238 2995 15315 3029
rect 15120 2956 15315 2995
rect 15120 2922 15132 2956
rect 15166 2922 15204 2956
rect 15238 2922 15315 2956
rect 15120 2883 15315 2922
rect 15120 2849 15132 2883
rect 15166 2849 15204 2883
rect 15238 2849 15315 2883
rect 15120 2810 15315 2849
rect 15120 2776 15132 2810
rect 15166 2776 15204 2810
rect 15238 2776 15315 2810
rect 15120 2737 15315 2776
rect 15120 2703 15132 2737
rect 15166 2703 15204 2737
rect 15238 2703 15315 2737
rect 15120 2664 15315 2703
rect 15120 2630 15132 2664
rect 15166 2630 15204 2664
rect 15238 2630 15315 2664
rect 15120 2591 15315 2630
rect 15120 2557 15132 2591
rect 15166 2557 15204 2591
rect 15238 2557 15315 2591
rect 15120 2518 15315 2557
rect 15120 2484 15132 2518
rect 15166 2484 15204 2518
rect 15238 2484 15315 2518
rect 15120 2445 15315 2484
rect 15120 2411 15132 2445
rect 15166 2411 15204 2445
rect 15238 2411 15315 2445
rect 15120 2372 15315 2411
rect 15120 2338 15132 2372
rect 15166 2338 15204 2372
rect 15238 2338 15315 2372
rect 15120 2299 15315 2338
rect 15120 2265 15132 2299
rect 15166 2265 15204 2299
rect 15238 2265 15315 2299
rect 15120 2226 15315 2265
rect 15120 2192 15132 2226
rect 15166 2192 15204 2226
rect 15238 2192 15315 2226
rect 15120 2153 15315 2192
rect 15120 2119 15132 2153
rect 15166 2119 15204 2153
rect 15238 2119 15315 2153
rect 15120 2080 15315 2119
rect 15120 2046 15132 2080
rect 15166 2046 15204 2080
rect 15238 2046 15315 2080
rect 15120 2007 15315 2046
rect 15120 1973 15132 2007
rect 15166 1973 15204 2007
rect 15238 1973 15315 2007
rect 15120 1934 15315 1973
rect 15120 1900 15132 1934
rect 15166 1900 15204 1934
rect 15238 1900 15315 1934
rect 15120 1861 15315 1900
rect 15120 1827 15132 1861
rect 15166 1827 15204 1861
rect 15238 1827 15315 1861
rect 15120 1788 15315 1827
rect 15120 1754 15132 1788
rect 15166 1754 15204 1788
rect 15238 1754 15315 1788
rect 15120 1715 15315 1754
rect 15120 1681 15132 1715
rect 15166 1681 15204 1715
rect 15238 1681 15315 1715
rect 15120 1642 15315 1681
rect 15120 1608 15132 1642
rect 15166 1608 15204 1642
rect 15238 1608 15315 1642
rect 15120 1569 15315 1608
rect 15120 1535 15132 1569
rect 15166 1535 15204 1569
rect 15238 1535 15315 1569
rect 15120 1496 15315 1535
rect 15120 1462 15132 1496
rect 15166 1462 15204 1496
rect 15238 1462 15315 1496
rect 15120 1423 15315 1462
rect 15120 1389 15132 1423
rect 15166 1389 15204 1423
rect 15238 1389 15315 1423
rect 15120 1350 15315 1389
rect 15120 1316 15132 1350
rect 15166 1316 15204 1350
rect 15238 1316 15315 1350
rect 15120 1277 15315 1316
rect 15120 1243 15132 1277
rect 15166 1243 15204 1277
rect 15238 1243 15315 1277
rect 15120 1204 15315 1243
rect 15120 1170 15132 1204
rect 15166 1170 15204 1204
rect 15238 1170 15315 1204
rect 15120 1131 15315 1170
rect 15120 1097 15132 1131
rect 15166 1097 15204 1131
rect 15238 1097 15315 1131
rect 15120 1058 15315 1097
rect 15120 1024 15132 1058
rect 15166 1024 15204 1058
rect 15238 1024 15315 1058
rect 15120 985 15315 1024
rect 15120 951 15132 985
rect 15166 951 15204 985
rect 15238 951 15315 985
rect 15120 912 15315 951
rect 15120 878 15132 912
rect 15166 878 15204 912
rect 15238 878 15315 912
rect 15120 839 15315 878
rect 15120 805 15132 839
rect 15166 805 15204 839
rect 15238 805 15315 839
rect 15120 766 15315 805
rect 15120 732 15132 766
rect 15166 732 15204 766
rect 15238 732 15315 766
rect 15120 693 15315 732
rect 15120 659 15132 693
rect 15166 659 15204 693
rect 15238 659 15315 693
rect 15120 620 15315 659
rect 15120 586 15132 620
rect 15166 586 15204 620
rect 15238 586 15315 620
rect 14637 574 14708 586
rect 13896 562 14708 574
tri 14708 562 14732 586 nw
rect 13896 547 14693 562
tri 14693 547 14708 562 nw
rect 15120 547 15315 586
rect 13896 513 14659 547
tri 14659 513 14693 547 nw
rect 15120 513 15132 547
rect 15166 513 15204 547
rect 15238 513 15315 547
rect 13896 490 14636 513
tri 14636 490 14659 513 nw
rect -4965 440 -4888 474
rect -4854 440 -4816 474
rect -4782 440 -4770 474
rect 15120 474 15315 513
tri -4770 440 -4744 466 sw
tri 15094 440 15120 466 se
rect 15120 440 15132 474
rect 15166 440 15204 474
rect 15238 440 15315 474
rect -4965 401 -4744 440
tri -4744 401 -4705 440 sw
tri 15055 401 15094 440 se
rect 15094 401 15315 440
rect -4965 367 -4888 401
rect -4854 367 -4816 401
rect -4782 367 -4705 401
tri -4705 367 -4671 401 sw
tri 15021 367 15055 401 se
rect 15055 367 15132 401
rect 15166 367 15204 401
rect 15238 367 15315 401
rect -4965 250 -4671 367
tri -4671 250 -4554 367 sw
tri 14904 250 15021 367 se
rect 15021 250 15315 367
tri -4965 120 -4835 250 ne
rect -4835 164 -3923 250
rect -4835 120 -4622 164
tri -4622 120 -4578 164 nw
tri -4488 120 -4444 164 ne
rect -4444 120 -3923 164
rect 14904 247 15229 250
rect 14903 164 15229 247
tri 15229 164 15315 250 nw
rect 14903 120 15185 164
tri 15185 120 15229 164 nw
<< rmetal1 >>
rect 14903 247 14904 250
use L1M1_C_CDNS_5246887918513  L1M1_C_CDNS_5246887918513_0
timestamp 1707688321
transform 1 0 13937 0 -1 1003
box 0 0 1 1
use L1M1_C_CDNS_5246887918513  L1M1_C_CDNS_5246887918513_1
timestamp 1707688321
transform 1 0 4917 0 -1 1025
box 0 0 1 1
use L1M1_C_CDNS_5246887918513  L1M1_C_CDNS_5246887918513_2
timestamp 1707688321
transform 1 0 3113 0 -1 1025
box 0 0 1 1
use L1M1_C_CDNS_5246887918513  L1M1_C_CDNS_5246887918513_3
timestamp 1707688321
transform 1 0 3625 0 -1 1025
box 0 0 1 1
use L1M1_C_CDNS_5246887918513  L1M1_C_CDNS_5246887918513_4
timestamp 1707688321
transform 1 0 1309 0 -1 1025
box 0 0 1 1
use L1M1_C_CDNS_5246887918513  L1M1_C_CDNS_5246887918513_5
timestamp 1707688321
transform 1 0 1821 0 -1 1025
box 0 0 1 1
use L1M1_C_CDNS_5246887918513  L1M1_C_CDNS_5246887918513_6
timestamp 1707688321
transform 1 0 17 0 -1 1025
box 0 0 1 1
use L1M1_C_CDNS_5246887918513  L1M1_C_CDNS_5246887918513_7
timestamp 1707688321
transform 1 0 -495 0 -1 1025
box 0 0 1 1
use L1M1_C_CDNS_5246887918513  L1M1_C_CDNS_5246887918513_8
timestamp 1707688321
transform 1 0 -2299 0 -1 1025
box 0 0 1 1
use L1M1_C_CDNS_5246887918513  L1M1_C_CDNS_5246887918513_9
timestamp 1707688321
transform 1 0 -1787 0 -1 1025
box 0 0 1 1
use L1M1_C_CDNS_5246887918513  L1M1_C_CDNS_5246887918513_10
timestamp 1707688321
transform 1 0 -3591 0 -1 1003
box 0 0 1 1
use L1M1_C_CDNS_5246887918513  L1M1_C_CDNS_5246887918513_11
timestamp 1707688321
transform 1 0 12133 0 -1 1025
box 0 0 1 1
use L1M1_C_CDNS_5246887918513  L1M1_C_CDNS_5246887918513_12
timestamp 1707688321
transform 1 0 12645 0 -1 1025
box 0 0 1 1
use L1M1_C_CDNS_5246887918513  L1M1_C_CDNS_5246887918513_13
timestamp 1707688321
transform 1 0 10329 0 -1 1025
box 0 0 1 1
use L1M1_C_CDNS_5246887918513  L1M1_C_CDNS_5246887918513_14
timestamp 1707688321
transform 1 0 10841 0 -1 1025
box 0 0 1 1
use L1M1_C_CDNS_5246887918513  L1M1_C_CDNS_5246887918513_15
timestamp 1707688321
transform 1 0 9037 0 -1 1025
box 0 0 1 1
use L1M1_C_CDNS_5246887918513  L1M1_C_CDNS_5246887918513_16
timestamp 1707688321
transform 1 0 8525 0 -1 1025
box 0 0 1 1
use L1M1_C_CDNS_5246887918513  L1M1_C_CDNS_5246887918513_17
timestamp 1707688321
transform 1 0 6721 0 -1 1025
box 0 0 1 1
use L1M1_C_CDNS_5246887918513  L1M1_C_CDNS_5246887918513_18
timestamp 1707688321
transform 1 0 7233 0 -1 1025
box 0 0 1 1
use L1M1_C_CDNS_5246887918513  L1M1_C_CDNS_5246887918513_19
timestamp 1707688321
transform 1 0 5429 0 -1 1025
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_0
timestamp 1707688321
transform 0 -1 14637 1 0 574
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_1
timestamp 1707688321
transform 0 -1 -4279 1 0 574
box 0 0 1 1
use L1M1_CDNS_524688791851534  L1M1_CDNS_524688791851534_0
timestamp 1707688321
transform 0 1 -4249 1 0 11692
box -12 -6 118 18688
use L1M1_CDNS_524688791851535  L1M1_CDNS_524688791851535_0
timestamp 1707688321
transform 0 1 -4217 -1 0 608
box -12 -6 118 18760
use L1M1_CDNS_524688791851536  L1M1_CDNS_524688791851536_0
timestamp 1707688321
transform 0 1 -3917 -1 0 238
box -12 -6 118 19048
use L1M1_CDNS_524688791851537  L1M1_CDNS_524688791851537_0
timestamp 1707688321
transform 1 0 14648 0 1 711
box -12 -6 118 10840
use L1M1_CDNS_524688791851537  L1M1_CDNS_524688791851537_1
timestamp 1707688321
transform 1 0 -4404 0 1 711
box -12 -6 118 10840
use L1M1_CDNS_524688791851538  L1M1_CDNS_524688791851538_0
timestamp 1707688321
transform 0 1 218 -1 0 12968
box -12 -6 118 14944
use PYL1_C_CDNS_5246887918514  PYL1_C_CDNS_5246887918514_0
timestamp 1707688321
transform 1 0 4917 0 -1 1025
box 0 0 1 1
use PYL1_C_CDNS_5246887918514  PYL1_C_CDNS_5246887918514_1
timestamp 1707688321
transform 1 0 3113 0 -1 1025
box 0 0 1 1
use PYL1_C_CDNS_5246887918514  PYL1_C_CDNS_5246887918514_2
timestamp 1707688321
transform 1 0 3625 0 -1 1025
box 0 0 1 1
use PYL1_C_CDNS_5246887918514  PYL1_C_CDNS_5246887918514_3
timestamp 1707688321
transform 1 0 1309 0 -1 1025
box 0 0 1 1
use PYL1_C_CDNS_5246887918514  PYL1_C_CDNS_5246887918514_4
timestamp 1707688321
transform 1 0 1821 0 -1 1025
box 0 0 1 1
use PYL1_C_CDNS_5246887918514  PYL1_C_CDNS_5246887918514_5
timestamp 1707688321
transform 1 0 17 0 -1 1025
box 0 0 1 1
use PYL1_C_CDNS_5246887918514  PYL1_C_CDNS_5246887918514_6
timestamp 1707688321
transform 1 0 -495 0 -1 1025
box 0 0 1 1
use PYL1_C_CDNS_5246887918514  PYL1_C_CDNS_5246887918514_7
timestamp 1707688321
transform 1 0 -2299 0 -1 1025
box 0 0 1 1
use PYL1_C_CDNS_5246887918514  PYL1_C_CDNS_5246887918514_8
timestamp 1707688321
transform 1 0 -1787 0 -1 1025
box 0 0 1 1
use PYL1_C_CDNS_5246887918514  PYL1_C_CDNS_5246887918514_9
timestamp 1707688321
transform 1 0 -3591 0 -1 1025
box 0 0 1 1
use PYL1_C_CDNS_5246887918514  PYL1_C_CDNS_5246887918514_10
timestamp 1707688321
transform 1 0 12133 0 -1 1025
box 0 0 1 1
use PYL1_C_CDNS_5246887918514  PYL1_C_CDNS_5246887918514_11
timestamp 1707688321
transform 1 0 12645 0 -1 1025
box 0 0 1 1
use PYL1_C_CDNS_5246887918514  PYL1_C_CDNS_5246887918514_12
timestamp 1707688321
transform 1 0 13937 0 -1 1025
box 0 0 1 1
use PYL1_C_CDNS_5246887918514  PYL1_C_CDNS_5246887918514_13
timestamp 1707688321
transform 1 0 10329 0 -1 1025
box 0 0 1 1
use PYL1_C_CDNS_5246887918514  PYL1_C_CDNS_5246887918514_14
timestamp 1707688321
transform 1 0 10841 0 -1 1025
box 0 0 1 1
use PYL1_C_CDNS_5246887918514  PYL1_C_CDNS_5246887918514_15
timestamp 1707688321
transform 1 0 9037 0 -1 1025
box 0 0 1 1
use PYL1_C_CDNS_5246887918514  PYL1_C_CDNS_5246887918514_16
timestamp 1707688321
transform 1 0 8525 0 -1 1025
box 0 0 1 1
use PYL1_C_CDNS_5246887918514  PYL1_C_CDNS_5246887918514_17
timestamp 1707688321
transform 1 0 6721 0 -1 1025
box 0 0 1 1
use PYL1_C_CDNS_5246887918514  PYL1_C_CDNS_5246887918514_18
timestamp 1707688321
transform 1 0 7233 0 -1 1025
box 0 0 1 1
use PYL1_C_CDNS_5246887918514  PYL1_C_CDNS_5246887918514_19
timestamp 1707688321
transform 1 0 5429 0 -1 1025
box 0 0 1 1
<< labels >>
flabel comment s 2595 11881 2595 11881 0 FreeSans 1000 0 0 0 condiode
flabel metal1 s 5055 11257 5315 11380 0 FreeSans 1000 180 0 0 gnd
port 1 nsew
flabel metal1 s 5956 11257 6216 11380 0 FreeSans 1000 180 0 0 pad
port 2 nsew
flabel metal1 s 6874 11257 7134 11380 0 FreeSans 1000 180 0 0 gnd
port 1 nsew
flabel metal1 s 7762 11257 8022 11380 0 FreeSans 1000 180 0 0 pad
port 2 nsew
flabel metal1 s 8667 11257 8927 11380 0 FreeSans 1000 180 0 0 gnd
port 1 nsew
flabel metal1 s 9577 11257 9837 11380 0 FreeSans 1000 180 0 0 pad
port 2 nsew
flabel metal1 s 10467 11257 10727 11380 0 FreeSans 1000 180 0 0 gnd
port 1 nsew
flabel metal1 s 11373 11257 11633 11380 0 FreeSans 1000 180 0 0 pad
port 2 nsew
flabel metal1 s 12264 11257 12524 11380 0 FreeSans 1000 180 0 0 gnd
port 1 nsew
flabel metal1 s 13140 11257 13400 11380 0 FreeSans 1000 180 0 0 pad
port 2 nsew
flabel metal1 s 14018 11257 14278 11380 0 FreeSans 1000 180 0 0 gnd
port 1 nsew
flabel metal1 s -4897 11038 -4797 11238 0 FreeSans 300 90 0 0 nwellRing
port 3 nsew
flabel metal1 s -4398 11039 -4298 11239 0 FreeSans 300 90 0 0 gnd
port 1 nsew
flabel metal1 s 6717 996 6775 1054 0 FreeSans 400 0 0 0 gate<11>
port 5 nsew
flabel metal1 s 7176 996 7228 1054 0 FreeSans 400 0 0 0 gate<12>
port 6 nsew
flabel metal1 s 8521 996 8579 1054 0 FreeSans 400 0 0 0 gate<13>
port 7 nsew
flabel metal1 s 8979 996 9035 1054 0 FreeSans 400 0 0 0 gate<14>
port 8 nsew
flabel metal1 s 10326 996 10385 1054 0 FreeSans 400 0 0 0 gate<15>
port 9 nsew
flabel metal1 s 10785 996 10840 1054 0 FreeSans 400 0 0 0 gate<16>
port 10 nsew
flabel metal1 s 12131 996 12184 1054 0 FreeSans 400 0 0 0 gate<17>
port 11 nsew
flabel metal1 s 12586 996 12643 1054 0 FreeSans 400 0 0 0 gate<18>
port 12 nsew
flabel metal1 s 13936 974 13991 1032 0 FreeSans 400 0 0 0 gate<19>
port 14 nsew
flabel metal1 s 5372 996 5425 1054 0 FreeSans 400 0 0 0 gate<10>
port 4 nsew
flabel metal1 s -3635 974 -3582 1032 0 FreeSans 400 0 0 0 gate<0>
port 15 nsew
flabel metal1 s -2290 992 -2232 1050 0 FreeSans 400 0 0 0 gate<1>
port 19 nsew
flabel metal1 s 1778 992 1833 1050 0 FreeSans 400 0 0 0 gate<6>
port 20 nsew
flabel metal1 s 1319 992 1378 1050 0 FreeSans 400 0 0 0 gate<5>
port 13 nsew
flabel metal1 s -28 992 28 1050 0 FreeSans 400 0 0 0 gate<4>
port 18 nsew
flabel metal1 s -486 992 -428 1050 0 FreeSans 400 0 0 0 gate<3>
port 17 nsew
flabel metal1 s -1831 992 -1779 1050 0 FreeSans 400 0 0 0 gate<2>
port 16 nsew
flabel metal1 s 4929 992 4984 1050 0 FreeSans 400 0 0 0 gate<9>
port 23 nsew
flabel metal1 s 3579 992 3636 1050 0 FreeSans 400 0 0 0 gate<8>
port 22 nsew
flabel metal1 s 3124 992 3177 1050 0 FreeSans 400 0 0 0 gate<7>
port 21 nsew
flabel metal1 s 4132 11257 4392 11380 0 FreeSans 1000 0 0 0 pad
port 2 nsew
flabel metal1 s 3180 11257 3440 11380 0 FreeSans 1000 0 0 0 gnd
port 1 nsew
flabel metal1 s 2292 11257 2552 11380 0 FreeSans 1000 0 0 0 pad
port 2 nsew
flabel metal1 s 1387 11257 1647 11380 0 FreeSans 1000 0 0 0 gnd
port 1 nsew
flabel metal1 s 477 11257 737 11380 0 FreeSans 1000 0 0 0 pad
port 2 nsew
flabel metal1 s -413 11257 -153 11380 0 FreeSans 1000 0 0 0 gnd
port 1 nsew
flabel metal1 s -1319 11257 -1059 11380 0 FreeSans 1000 0 0 0 pad
port 2 nsew
flabel metal1 s -2210 11257 -1950 11380 0 FreeSans 1000 0 0 0 gnd
port 1 nsew
flabel metal1 s -3086 11257 -2826 11380 0 FreeSans 1000 0 0 0 pad
port 2 nsew
flabel metal1 s -3964 11257 -3704 11380 0 FreeSans 1000 0 0 0 gnd
port 1 nsew
<< properties >>
string GDS_END 93352904
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 92165670
<< end >>
