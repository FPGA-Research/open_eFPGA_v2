magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -107 515 487 1337
<< pwell >>
rect -67 367 67 455
rect 313 367 447 455
<< mvpsubdiff >>
rect -41 427 41 429
rect -41 393 -17 427
rect 17 393 41 427
rect 339 427 421 429
rect 339 393 363 427
rect 397 393 421 427
<< mvnsubdiff >>
rect -41 583 -17 617
rect 17 583 41 617
rect -41 581 41 583
rect 339 583 363 617
rect 397 583 421 617
rect 339 581 421 583
<< mvpsubdiffcont >>
rect -17 393 17 427
rect 363 393 397 427
<< mvnsubdiffcont >>
rect -17 583 17 617
rect 363 583 397 617
<< poly >>
rect 35 1353 169 1369
rect 35 1319 51 1353
rect 85 1319 119 1353
rect 153 1319 169 1353
rect 35 1297 169 1319
rect 211 1353 345 1369
rect 211 1319 227 1353
rect 261 1319 295 1353
rect 329 1319 345 1353
rect 211 1297 345 1319
rect 52 557 162 645
rect 52 523 89 557
rect 123 523 162 557
rect 52 489 162 523
rect 52 455 89 489
rect 123 455 162 489
rect 52 345 162 455
rect 218 557 328 645
rect 218 523 257 557
rect 291 523 328 557
rect 218 489 328 523
rect 218 455 257 489
rect 291 455 328 489
rect 218 345 328 455
rect 35 71 169 93
rect 35 37 51 71
rect 85 37 119 71
rect 153 37 169 71
rect 35 21 169 37
rect 211 71 345 93
rect 211 37 227 71
rect 261 37 295 71
rect 329 37 345 71
rect 211 21 345 37
<< polycont >>
rect 51 1319 85 1353
rect 119 1319 153 1353
rect 227 1319 261 1353
rect 295 1319 329 1353
rect 89 523 123 557
rect 89 455 123 489
rect 257 523 291 557
rect 257 455 291 489
rect 51 37 85 71
rect 119 37 153 71
rect 227 37 261 71
rect 295 37 329 71
<< locali >>
rect 51 1353 153 1369
rect 85 1319 119 1353
rect 51 1303 153 1319
rect 227 1353 329 1369
rect 261 1319 295 1353
rect 227 1303 329 1319
rect -17 785 17 823
rect -17 713 17 751
rect -17 667 17 679
rect -17 567 17 583
rect 65 557 139 1303
rect 65 523 89 557
rect 123 523 139 557
rect 65 489 139 523
rect 65 455 89 489
rect 123 455 139 489
rect -17 427 17 443
rect -17 259 17 297
rect -17 187 17 225
rect 65 87 139 455
rect 173 943 207 1013
rect 173 121 207 909
rect 241 557 315 1303
rect 363 943 397 1270
rect 363 673 397 909
rect 363 567 397 583
rect 241 523 257 557
rect 291 523 315 557
rect 241 489 315 523
rect 241 455 257 489
rect 291 455 315 489
rect 241 87 315 455
rect 363 427 397 443
rect 363 259 397 297
rect 363 187 397 225
rect 51 71 153 87
rect 85 37 119 71
rect 51 21 153 37
rect 227 71 329 87
rect 261 37 295 71
rect 227 21 329 37
<< viali >>
rect -17 823 17 857
rect -17 751 17 785
rect -17 679 17 713
rect -17 617 17 633
rect -17 599 17 617
rect -17 393 17 411
rect -17 377 17 393
rect -17 297 17 331
rect -17 225 17 259
rect -17 153 17 187
rect 173 909 207 943
rect 363 909 397 943
rect 363 617 397 633
rect 363 599 397 617
rect 363 393 397 411
rect 363 377 397 393
rect 363 297 397 331
rect 363 225 397 259
rect 363 153 397 187
<< metal1 >>
rect 167 943 403 955
rect 167 909 173 943
rect 207 909 363 943
rect 397 909 403 943
rect 167 897 403 909
rect -29 857 409 869
rect -29 823 -17 857
rect 17 823 409 857
rect -29 785 409 823
rect -29 751 -17 785
rect 17 751 409 785
rect -29 713 409 751
rect -29 679 -17 713
rect 17 679 409 713
rect -29 667 409 679
rect -29 633 409 639
rect -29 599 -17 633
rect 17 599 363 633
rect 397 599 409 633
rect -29 593 409 599
rect -29 411 409 417
rect -29 377 -17 411
rect 17 377 363 411
rect 397 377 409 411
rect -29 371 409 377
rect -29 331 409 343
rect -29 297 -17 331
rect 17 297 363 331
rect 397 297 409 331
rect -29 259 409 297
rect -29 225 -17 259
rect 17 225 363 259
rect 397 225 409 259
rect -29 187 409 225
rect -29 153 -17 187
rect 17 153 363 187
rect 397 153 409 187
rect -29 141 409 153
use hvnTran_CDNS_52468879185364  hvnTran_CDNS_52468879185364_0
timestamp 1707688321
transform 1 0 42 0 -1 319
box -93 -26 389 226
use hvpTran_CDNS_52468879185361  hvpTran_CDNS_52468879185361_0
timestamp 1707688321
transform -1 0 338 0 1 671
box -133 -66 236 666
use hvpTran_CDNS_52468879185361  hvpTran_CDNS_52468879185361_1
timestamp 1707688321
transform 1 0 42 0 1 671
box -133 -66 236 666
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1707688321
transform 0 -1 397 -1 0 331
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1707688321
transform 0 -1 17 -1 0 331
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_2
timestamp 1707688321
transform 0 -1 17 1 0 679
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_0
timestamp 1707688321
transform -1 0 17 0 -1 633
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_1
timestamp 1707688321
transform 0 -1 207 1 0 909
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_2
timestamp 1707688321
transform 0 -1 397 1 0 909
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_3
timestamp 1707688321
transform 1 0 363 0 -1 411
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_4
timestamp 1707688321
transform 1 0 -17 0 -1 411
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_5
timestamp 1707688321
transform 1 0 363 0 -1 633
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_0
timestamp 1707688321
transform 0 -1 139 1 0 439
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_1
timestamp 1707688321
transform 0 -1 307 1 0 439
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_2
timestamp 1707688321
transform 1 0 211 0 1 21
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_3
timestamp 1707688321
transform 1 0 35 0 1 21
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_4
timestamp 1707688321
transform 1 0 35 0 1 1303
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_5
timestamp 1707688321
transform 1 0 211 0 1 1303
box 0 0 1 1
<< labels >>
flabel metal1 s 0 667 23 869 3 FreeSans 200 0 0 0 vpwr
port 1 nsew
flabel metal1 s 0 593 23 639 3 FreeSans 200 0 0 0 vpb
port 2 nsew
flabel metal1 s 0 371 23 417 3 FreeSans 200 0 0 0 vnb
port 3 nsew
flabel metal1 s 0 141 23 343 3 FreeSans 200 0 0 0 vgnd
port 4 nsew
flabel metal1 s 357 141 380 343 7 FreeSans 200 0 0 0 vgnd
port 4 nsew
flabel metal1 s 357 371 380 417 7 FreeSans 200 0 0 0 vnb
port 3 nsew
flabel metal1 s 357 593 380 639 7 FreeSans 200 0 0 0 vpb
port 2 nsew
flabel metal1 s 357 667 380 869 7 FreeSans 200 0 0 0 vpwr
port 1 nsew
flabel locali s 363 1209 397 1270 0 FreeSans 200 0 0 0 out
port 6 nsew
flabel locali s 85 1303 119 1369 0 FreeSans 200 0 0 0 in0
port 7 nsew
flabel locali s 261 1303 295 1369 0 FreeSans 200 0 0 0 in1
port 8 nsew
flabel locali s 86 21 119 87 0 FreeSans 200 0 0 0 in0
port 7 nsew
flabel locali s 261 21 295 87 0 FreeSans 200 0 0 0 in1
port 8 nsew
<< properties >>
string GDS_END 87674976
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87669814
<< end >>
