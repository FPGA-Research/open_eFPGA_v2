magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -88 17172 1318 17258
rect -88 -2 -2 17172
rect 616 12879 768 17172
rect 1078 8586 1318 17172
rect 1232 -2 1318 8586
rect -88 -88 1318 -2
<< ndiff >>
rect 642 17136 742 17144
rect 642 17102 675 17136
rect 709 17102 742 17136
rect 642 16834 742 17102
rect 642 16800 675 16834
rect 709 16800 742 16834
rect 642 16532 742 16800
rect 642 16498 675 16532
rect 709 16498 742 16532
rect 642 16230 742 16498
rect 642 16196 675 16230
rect 709 16196 742 16230
rect 642 15928 742 16196
rect 642 15894 675 15928
rect 709 15894 742 15928
rect 642 15626 742 15894
rect 642 15592 675 15626
rect 709 15592 742 15626
rect 642 15324 742 15592
rect 642 15290 675 15324
rect 709 15290 742 15324
rect 642 15022 742 15290
rect 642 14988 675 15022
rect 709 14988 742 15022
rect 642 14720 742 14988
rect 642 14686 675 14720
rect 709 14686 742 14720
rect 642 14418 742 14686
rect 642 14384 675 14418
rect 709 14384 742 14418
rect 642 14116 742 14384
rect 642 14082 675 14116
rect 709 14082 742 14116
rect 642 13814 742 14082
rect 642 13780 675 13814
rect 709 13780 742 13814
rect 642 13512 742 13780
rect 642 13478 675 13512
rect 709 13478 742 13512
rect 642 13210 742 13478
rect 642 13176 675 13210
rect 709 13176 742 13210
rect 642 12905 742 13176
rect 1104 17136 1204 17144
rect 1104 17102 1137 17136
rect 1171 17102 1204 17136
rect 1104 16834 1204 17102
rect 1104 16800 1137 16834
rect 1171 16800 1204 16834
rect 1104 16532 1204 16800
rect 1104 16498 1137 16532
rect 1171 16498 1204 16532
rect 1104 16230 1204 16498
rect 1104 16196 1137 16230
rect 1171 16196 1204 16230
rect 1104 15928 1204 16196
rect 1104 15894 1137 15928
rect 1171 15894 1204 15928
rect 1104 15626 1204 15894
rect 1104 15592 1137 15626
rect 1171 15592 1204 15626
rect 1104 15324 1204 15592
rect 1104 15290 1137 15324
rect 1171 15290 1204 15324
rect 1104 15022 1204 15290
rect 1104 14988 1137 15022
rect 1171 14988 1204 15022
rect 1104 14720 1204 14988
rect 1104 14686 1137 14720
rect 1171 14686 1204 14720
rect 1104 14418 1204 14686
rect 1104 14384 1137 14418
rect 1171 14384 1204 14418
rect 1104 14116 1204 14384
rect 1104 14082 1137 14116
rect 1171 14082 1204 14116
rect 1104 13814 1204 14082
rect 1104 13780 1137 13814
rect 1171 13780 1204 13814
rect 1104 13512 1204 13780
rect 1104 13478 1137 13512
rect 1171 13478 1204 13512
rect 1104 13210 1204 13478
rect 1104 13176 1137 13210
rect 1171 13176 1204 13210
rect 1104 12908 1204 13176
rect 1104 12874 1137 12908
rect 1171 12874 1204 12908
rect 1104 12606 1204 12874
rect 1104 12572 1137 12606
rect 1171 12572 1204 12606
rect 1104 12304 1204 12572
rect 1104 12270 1137 12304
rect 1171 12270 1204 12304
rect 1104 12002 1204 12270
rect 1104 11968 1137 12002
rect 1171 11968 1204 12002
rect 1104 11700 1204 11968
rect 1104 11666 1137 11700
rect 1171 11666 1204 11700
rect 1104 11398 1204 11666
rect 1104 11364 1137 11398
rect 1171 11364 1204 11398
rect 1104 11096 1204 11364
rect 1104 11062 1137 11096
rect 1171 11062 1204 11096
rect 1104 10794 1204 11062
rect 1104 10760 1137 10794
rect 1171 10760 1204 10794
rect 1104 10492 1204 10760
rect 1104 10458 1137 10492
rect 1171 10458 1204 10492
rect 1104 10190 1204 10458
rect 1104 10156 1137 10190
rect 1171 10156 1204 10190
rect 1104 9888 1204 10156
rect 1104 9854 1137 9888
rect 1171 9854 1204 9888
rect 1104 9586 1204 9854
rect 1104 9552 1137 9586
rect 1171 9552 1204 9586
rect 1104 9284 1204 9552
rect 1104 9250 1137 9284
rect 1171 9250 1204 9284
rect 1104 8982 1204 9250
rect 1104 8948 1137 8982
rect 1171 8948 1204 8982
rect 1104 8612 1204 8948
<< ndiffc >>
rect 675 17102 709 17136
rect 675 16800 709 16834
rect 675 16498 709 16532
rect 675 16196 709 16230
rect 675 15894 709 15928
rect 675 15592 709 15626
rect 675 15290 709 15324
rect 675 14988 709 15022
rect 675 14686 709 14720
rect 675 14384 709 14418
rect 675 14082 709 14116
rect 675 13780 709 13814
rect 675 13478 709 13512
rect 675 13176 709 13210
rect 1137 17102 1171 17136
rect 1137 16800 1171 16834
rect 1137 16498 1171 16532
rect 1137 16196 1171 16230
rect 1137 15894 1171 15928
rect 1137 15592 1171 15626
rect 1137 15290 1171 15324
rect 1137 14988 1171 15022
rect 1137 14686 1171 14720
rect 1137 14384 1171 14418
rect 1137 14082 1171 14116
rect 1137 13780 1171 13814
rect 1137 13478 1171 13512
rect 1137 13176 1171 13210
rect 1137 12874 1171 12908
rect 1137 12572 1171 12606
rect 1137 12270 1171 12304
rect 1137 11968 1171 12002
rect 1137 11666 1171 11700
rect 1137 11364 1171 11398
rect 1137 11062 1171 11096
rect 1137 10760 1171 10794
rect 1137 10458 1171 10492
rect 1137 10156 1171 10190
rect 1137 9854 1171 9888
rect 1137 9552 1171 9586
rect 1137 9250 1171 9284
rect 1137 8948 1171 8982
<< psubdiff >>
rect -62 17198 34 17232
rect 68 17198 102 17232
rect 136 17198 170 17232
rect 204 17198 238 17232
rect 272 17198 306 17232
rect 340 17198 374 17232
rect 408 17198 442 17232
rect 476 17198 510 17232
rect 544 17198 578 17232
rect 612 17198 646 17232
rect 680 17198 714 17232
rect 748 17198 782 17232
rect 816 17198 850 17232
rect 884 17198 918 17232
rect 952 17198 986 17232
rect 1020 17198 1054 17232
rect 1088 17198 1122 17232
rect 1156 17198 1190 17232
rect 1224 17198 1292 17232
rect -62 17164 -28 17198
rect -62 17096 -28 17130
rect -62 17028 -28 17062
rect -62 16960 -28 16994
rect -62 16892 -28 16926
rect -62 16824 -28 16858
rect -62 16756 -28 16790
rect -62 16688 -28 16722
rect -62 16620 -28 16654
rect -62 16552 -28 16586
rect -62 16484 -28 16518
rect -62 16416 -28 16450
rect -62 16348 -28 16382
rect -62 16280 -28 16314
rect -62 16212 -28 16246
rect -62 16144 -28 16178
rect -62 16076 -28 16110
rect -62 16008 -28 16042
rect -62 15940 -28 15974
rect -62 15872 -28 15906
rect -62 15804 -28 15838
rect -62 15736 -28 15770
rect -62 15668 -28 15702
rect -62 15600 -28 15634
rect -62 15532 -28 15566
rect -62 15464 -28 15498
rect -62 15396 -28 15430
rect -62 15328 -28 15362
rect -62 15260 -28 15294
rect -62 15192 -28 15226
rect -62 15124 -28 15158
rect -62 15056 -28 15090
rect -62 14988 -28 15022
rect -62 14920 -28 14954
rect -62 14852 -28 14886
rect -62 14784 -28 14818
rect -62 14716 -28 14750
rect -62 14648 -28 14682
rect -62 14580 -28 14614
rect -62 14512 -28 14546
rect -62 14444 -28 14478
rect -62 14376 -28 14410
rect -62 14308 -28 14342
rect -62 14240 -28 14274
rect -62 14172 -28 14206
rect -62 14104 -28 14138
rect -62 14036 -28 14070
rect -62 13968 -28 14002
rect -62 13900 -28 13934
rect -62 13832 -28 13866
rect -62 13764 -28 13798
rect -62 13696 -28 13730
rect -62 13628 -28 13662
rect -62 13560 -28 13594
rect -62 13492 -28 13526
rect -62 13424 -28 13458
rect -62 13356 -28 13390
rect -62 13288 -28 13322
rect -62 13220 -28 13254
rect -62 13152 -28 13186
rect -62 13084 -28 13118
rect -62 13016 -28 13050
rect -62 12948 -28 12982
rect -62 12880 -28 12914
rect -62 12812 -28 12846
rect -62 12744 -28 12778
rect -62 12676 -28 12710
rect -62 12608 -28 12642
rect -62 12540 -28 12574
rect -62 12472 -28 12506
rect -62 12404 -28 12438
rect -62 12336 -28 12370
rect -62 12268 -28 12302
rect -62 12200 -28 12234
rect -62 12132 -28 12166
rect -62 12064 -28 12098
rect -62 11996 -28 12030
rect -62 11928 -28 11962
rect -62 11860 -28 11894
rect -62 11792 -28 11826
rect -62 11724 -28 11758
rect -62 11656 -28 11690
rect -62 11588 -28 11622
rect -62 11520 -28 11554
rect -62 11452 -28 11486
rect -62 11384 -28 11418
rect -62 11316 -28 11350
rect -62 11248 -28 11282
rect -62 11180 -28 11214
rect -62 11112 -28 11146
rect -62 11044 -28 11078
rect -62 10976 -28 11010
rect -62 10908 -28 10942
rect -62 10840 -28 10874
rect -62 10772 -28 10806
rect -62 10704 -28 10738
rect -62 10636 -28 10670
rect -62 10568 -28 10602
rect -62 10500 -28 10534
rect -62 10432 -28 10466
rect -62 10364 -28 10398
rect -62 10296 -28 10330
rect -62 10228 -28 10262
rect -62 10160 -28 10194
rect -62 10092 -28 10126
rect -62 10024 -28 10058
rect -62 9956 -28 9990
rect -62 9888 -28 9922
rect -62 9820 -28 9854
rect -62 9752 -28 9786
rect -62 9684 -28 9718
rect -62 9616 -28 9650
rect -62 9548 -28 9582
rect -62 9480 -28 9514
rect -62 9412 -28 9446
rect -62 9344 -28 9378
rect -62 9276 -28 9310
rect -62 9208 -28 9242
rect -62 9140 -28 9174
rect -62 9072 -28 9106
rect -62 9004 -28 9038
rect -62 8936 -28 8970
rect -62 8868 -28 8902
rect -62 8800 -28 8834
rect -62 8732 -28 8766
rect -62 8664 -28 8698
rect -62 8596 -28 8630
rect 1258 17108 1292 17198
rect 1258 17040 1292 17074
rect 1258 16972 1292 17006
rect 1258 16904 1292 16938
rect 1258 16836 1292 16870
rect 1258 16768 1292 16802
rect 1258 16700 1292 16734
rect 1258 16632 1292 16666
rect 1258 16564 1292 16598
rect 1258 16496 1292 16530
rect 1258 16428 1292 16462
rect 1258 16360 1292 16394
rect 1258 16292 1292 16326
rect 1258 16224 1292 16258
rect 1258 16156 1292 16190
rect 1258 16088 1292 16122
rect 1258 16020 1292 16054
rect 1258 15952 1292 15986
rect 1258 15884 1292 15918
rect 1258 15816 1292 15850
rect 1258 15748 1292 15782
rect 1258 15680 1292 15714
rect 1258 15612 1292 15646
rect 1258 15544 1292 15578
rect 1258 15476 1292 15510
rect 1258 15408 1292 15442
rect 1258 15340 1292 15374
rect 1258 15272 1292 15306
rect 1258 15204 1292 15238
rect 1258 15136 1292 15170
rect 1258 15068 1292 15102
rect 1258 15000 1292 15034
rect 1258 14932 1292 14966
rect 1258 14864 1292 14898
rect 1258 14796 1292 14830
rect 1258 14728 1292 14762
rect 1258 14660 1292 14694
rect 1258 14592 1292 14626
rect 1258 14524 1292 14558
rect 1258 14456 1292 14490
rect 1258 14388 1292 14422
rect 1258 14320 1292 14354
rect 1258 14252 1292 14286
rect 1258 14184 1292 14218
rect 1258 14116 1292 14150
rect 1258 14048 1292 14082
rect 1258 13980 1292 14014
rect 1258 13912 1292 13946
rect 1258 13844 1292 13878
rect 1258 13776 1292 13810
rect 1258 13708 1292 13742
rect 1258 13640 1292 13674
rect 1258 13572 1292 13606
rect 1258 13504 1292 13538
rect 1258 13436 1292 13470
rect 1258 13368 1292 13402
rect 1258 13300 1292 13334
rect 1258 13232 1292 13266
rect 1258 13164 1292 13198
rect 1258 13096 1292 13130
rect 1258 13028 1292 13062
rect 1258 12960 1292 12994
rect 1258 12892 1292 12926
rect 1258 12824 1292 12858
rect 1258 12756 1292 12790
rect 1258 12688 1292 12722
rect 1258 12620 1292 12654
rect 1258 12552 1292 12586
rect 1258 12484 1292 12518
rect 1258 12416 1292 12450
rect 1258 12348 1292 12382
rect 1258 12280 1292 12314
rect 1258 12212 1292 12246
rect 1258 12144 1292 12178
rect 1258 12076 1292 12110
rect 1258 12008 1292 12042
rect 1258 11940 1292 11974
rect 1258 11872 1292 11906
rect 1258 11804 1292 11838
rect 1258 11736 1292 11770
rect 1258 11668 1292 11702
rect 1258 11600 1292 11634
rect 1258 11532 1292 11566
rect 1258 11464 1292 11498
rect 1258 11396 1292 11430
rect 1258 11328 1292 11362
rect 1258 11260 1292 11294
rect 1258 11192 1292 11226
rect 1258 11124 1292 11158
rect 1258 11056 1292 11090
rect 1258 10988 1292 11022
rect 1258 10920 1292 10954
rect 1258 10852 1292 10886
rect 1258 10784 1292 10818
rect 1258 10716 1292 10750
rect 1258 10648 1292 10682
rect 1258 10580 1292 10614
rect 1258 10512 1292 10546
rect 1258 10444 1292 10478
rect 1258 10376 1292 10410
rect 1258 10308 1292 10342
rect 1258 10240 1292 10274
rect 1258 10172 1292 10206
rect 1258 10104 1292 10138
rect 1258 10036 1292 10070
rect 1258 9968 1292 10002
rect 1258 9900 1292 9934
rect 1258 9832 1292 9866
rect 1258 9764 1292 9798
rect 1258 9696 1292 9730
rect 1258 9628 1292 9662
rect 1258 9560 1292 9594
rect 1258 9492 1292 9526
rect 1258 9424 1292 9458
rect 1258 9356 1292 9390
rect 1258 9288 1292 9322
rect 1258 9220 1292 9254
rect 1258 9152 1292 9186
rect 1258 9084 1292 9118
rect 1258 9016 1292 9050
rect 1258 8948 1292 8982
rect 1258 8880 1292 8914
rect 1258 8812 1292 8846
rect 1258 8744 1292 8778
rect 1258 8676 1292 8710
rect -62 8528 -28 8562
rect -62 8460 -28 8494
rect -62 8392 -28 8426
rect -62 8324 -28 8358
rect -62 8256 -28 8290
rect -62 8188 -28 8222
rect -62 8120 -28 8154
rect -62 8052 -28 8086
rect -62 7984 -28 8018
rect -62 7916 -28 7950
rect -62 7848 -28 7882
rect -62 7780 -28 7814
rect -62 7712 -28 7746
rect -62 7644 -28 7678
rect -62 7576 -28 7610
rect -62 7508 -28 7542
rect -62 7440 -28 7474
rect -62 7372 -28 7406
rect -62 7304 -28 7338
rect -62 7236 -28 7270
rect -62 7168 -28 7202
rect -62 7100 -28 7134
rect -62 7032 -28 7066
rect -62 6964 -28 6998
rect -62 6896 -28 6930
rect -62 6828 -28 6862
rect -62 6760 -28 6794
rect -62 6692 -28 6726
rect -62 6624 -28 6658
rect -62 6556 -28 6590
rect -62 6488 -28 6522
rect -62 6420 -28 6454
rect -62 6352 -28 6386
rect -62 6284 -28 6318
rect -62 6216 -28 6250
rect -62 6148 -28 6182
rect -62 6080 -28 6114
rect -62 6012 -28 6046
rect -62 5944 -28 5978
rect -62 5876 -28 5910
rect -62 5808 -28 5842
rect -62 5740 -28 5774
rect -62 5672 -28 5706
rect -62 5604 -28 5638
rect -62 5536 -28 5570
rect -62 5468 -28 5502
rect -62 5400 -28 5434
rect -62 5332 -28 5366
rect -62 5264 -28 5298
rect -62 5196 -28 5230
rect -62 5128 -28 5162
rect -62 5060 -28 5094
rect -62 4992 -28 5026
rect -62 4924 -28 4958
rect -62 4856 -28 4890
rect -62 4788 -28 4822
rect -62 4720 -28 4754
rect -62 4652 -28 4686
rect -62 4584 -28 4618
rect -62 4516 -28 4550
rect -62 4448 -28 4482
rect -62 4380 -28 4414
rect -62 4312 -28 4346
rect -62 4244 -28 4278
rect -62 4176 -28 4210
rect -62 4108 -28 4142
rect -62 4040 -28 4074
rect -62 3972 -28 4006
rect -62 3904 -28 3938
rect -62 3836 -28 3870
rect -62 3768 -28 3802
rect -62 3700 -28 3734
rect -62 3632 -28 3666
rect -62 3564 -28 3598
rect -62 3496 -28 3530
rect -62 3428 -28 3462
rect -62 3360 -28 3394
rect -62 3292 -28 3326
rect -62 3224 -28 3258
rect -62 3156 -28 3190
rect -62 3088 -28 3122
rect -62 3020 -28 3054
rect -62 2952 -28 2986
rect -62 2884 -28 2918
rect -62 2816 -28 2850
rect -62 2748 -28 2782
rect -62 2680 -28 2714
rect -62 2612 -28 2646
rect -62 2544 -28 2578
rect -62 2476 -28 2510
rect -62 2408 -28 2442
rect -62 2340 -28 2374
rect -62 2272 -28 2306
rect -62 2204 -28 2238
rect -62 2136 -28 2170
rect -62 2068 -28 2102
rect -62 2000 -28 2034
rect -62 1932 -28 1966
rect -62 1864 -28 1898
rect -62 1796 -28 1830
rect -62 1728 -28 1762
rect -62 1660 -28 1694
rect -62 1592 -28 1626
rect -62 1524 -28 1558
rect -62 1456 -28 1490
rect -62 1388 -28 1422
rect -62 1320 -28 1354
rect -62 1252 -28 1286
rect -62 1184 -28 1218
rect -62 1116 -28 1150
rect -62 1048 -28 1082
rect -62 980 -28 1014
rect -62 912 -28 946
rect -62 844 -28 878
rect -62 776 -28 810
rect -62 708 -28 742
rect -62 640 -28 674
rect -62 572 -28 606
rect -62 504 -28 538
rect -62 436 -28 470
rect -62 368 -28 402
rect -62 300 -28 334
rect -62 232 -28 266
rect -62 164 -28 198
rect -62 96 -28 130
rect -62 -28 -28 62
rect 1258 8608 1292 8642
rect 1258 8540 1292 8574
rect 1258 8472 1292 8506
rect 1258 8404 1292 8438
rect 1258 8336 1292 8370
rect 1258 8268 1292 8302
rect 1258 8200 1292 8234
rect 1258 8132 1292 8166
rect 1258 8064 1292 8098
rect 1258 7996 1292 8030
rect 1258 7928 1292 7962
rect 1258 7860 1292 7894
rect 1258 7792 1292 7826
rect 1258 7724 1292 7758
rect 1258 7656 1292 7690
rect 1258 7588 1292 7622
rect 1258 7520 1292 7554
rect 1258 7452 1292 7486
rect 1258 7384 1292 7418
rect 1258 7316 1292 7350
rect 1258 7248 1292 7282
rect 1258 7180 1292 7214
rect 1258 7112 1292 7146
rect 1258 7044 1292 7078
rect 1258 6976 1292 7010
rect 1258 6908 1292 6942
rect 1258 6840 1292 6874
rect 1258 6772 1292 6806
rect 1258 6704 1292 6738
rect 1258 6636 1292 6670
rect 1258 6568 1292 6602
rect 1258 6500 1292 6534
rect 1258 6432 1292 6466
rect 1258 6364 1292 6398
rect 1258 6296 1292 6330
rect 1258 6228 1292 6262
rect 1258 6160 1292 6194
rect 1258 6092 1292 6126
rect 1258 6024 1292 6058
rect 1258 5956 1292 5990
rect 1258 5888 1292 5922
rect 1258 5820 1292 5854
rect 1258 5752 1292 5786
rect 1258 5684 1292 5718
rect 1258 5616 1292 5650
rect 1258 5548 1292 5582
rect 1258 5480 1292 5514
rect 1258 5412 1292 5446
rect 1258 5344 1292 5378
rect 1258 5276 1292 5310
rect 1258 5208 1292 5242
rect 1258 5140 1292 5174
rect 1258 5072 1292 5106
rect 1258 5004 1292 5038
rect 1258 4936 1292 4970
rect 1258 4868 1292 4902
rect 1258 4800 1292 4834
rect 1258 4732 1292 4766
rect 1258 4664 1292 4698
rect 1258 4596 1292 4630
rect 1258 4528 1292 4562
rect 1258 4460 1292 4494
rect 1258 4392 1292 4426
rect 1258 4324 1292 4358
rect 1258 4256 1292 4290
rect 1258 4188 1292 4222
rect 1258 4120 1292 4154
rect 1258 4052 1292 4086
rect 1258 3984 1292 4018
rect 1258 3916 1292 3950
rect 1258 3848 1292 3882
rect 1258 3780 1292 3814
rect 1258 3712 1292 3746
rect 1258 3644 1292 3678
rect 1258 3576 1292 3610
rect 1258 3508 1292 3542
rect 1258 3440 1292 3474
rect 1258 3372 1292 3406
rect 1258 3304 1292 3338
rect 1258 3236 1292 3270
rect 1258 3168 1292 3202
rect 1258 3100 1292 3134
rect 1258 3032 1292 3066
rect 1258 2964 1292 2998
rect 1258 2896 1292 2930
rect 1258 2828 1292 2862
rect 1258 2760 1292 2794
rect 1258 2692 1292 2726
rect 1258 2624 1292 2658
rect 1258 2556 1292 2590
rect 1258 2488 1292 2522
rect 1258 2420 1292 2454
rect 1258 2352 1292 2386
rect 1258 2284 1292 2318
rect 1258 2216 1292 2250
rect 1258 2148 1292 2182
rect 1258 2080 1292 2114
rect 1258 2012 1292 2046
rect 1258 1944 1292 1978
rect 1258 1876 1292 1910
rect 1258 1808 1292 1842
rect 1258 1740 1292 1774
rect 1258 1672 1292 1706
rect 1258 1604 1292 1638
rect 1258 1536 1292 1570
rect 1258 1468 1292 1502
rect 1258 1400 1292 1434
rect 1258 1332 1292 1366
rect 1258 1264 1292 1298
rect 1258 1196 1292 1230
rect 1258 1128 1292 1162
rect 1258 1060 1292 1094
rect 1258 992 1292 1026
rect 1258 924 1292 958
rect 1258 856 1292 890
rect 1258 788 1292 822
rect 1258 720 1292 754
rect 1258 652 1292 686
rect 1258 584 1292 618
rect 1258 516 1292 550
rect 1258 448 1292 482
rect 1258 380 1292 414
rect 1258 312 1292 346
rect 1258 244 1292 278
rect 1258 176 1292 210
rect 1258 108 1292 142
rect 1258 40 1292 74
rect 1258 -28 1292 6
rect -62 -62 6 -28
rect 40 -62 74 -28
rect 108 -62 142 -28
rect 176 -62 210 -28
rect 244 -62 278 -28
rect 312 -62 346 -28
rect 380 -62 414 -28
rect 448 -62 482 -28
rect 516 -62 550 -28
rect 584 -62 618 -28
rect 652 -62 686 -28
rect 720 -62 754 -28
rect 788 -62 822 -28
rect 856 -62 890 -28
rect 924 -62 958 -28
rect 992 -62 1026 -28
rect 1060 -62 1094 -28
rect 1128 -62 1162 -28
rect 1196 -62 1292 -28
<< psubdiffcont >>
rect 34 17198 68 17232
rect 102 17198 136 17232
rect 170 17198 204 17232
rect 238 17198 272 17232
rect 306 17198 340 17232
rect 374 17198 408 17232
rect 442 17198 476 17232
rect 510 17198 544 17232
rect 578 17198 612 17232
rect 646 17198 680 17232
rect 714 17198 748 17232
rect 782 17198 816 17232
rect 850 17198 884 17232
rect 918 17198 952 17232
rect 986 17198 1020 17232
rect 1054 17198 1088 17232
rect 1122 17198 1156 17232
rect 1190 17198 1224 17232
rect -62 17130 -28 17164
rect -62 17062 -28 17096
rect -62 16994 -28 17028
rect -62 16926 -28 16960
rect -62 16858 -28 16892
rect -62 16790 -28 16824
rect -62 16722 -28 16756
rect -62 16654 -28 16688
rect -62 16586 -28 16620
rect -62 16518 -28 16552
rect -62 16450 -28 16484
rect -62 16382 -28 16416
rect -62 16314 -28 16348
rect -62 16246 -28 16280
rect -62 16178 -28 16212
rect -62 16110 -28 16144
rect -62 16042 -28 16076
rect -62 15974 -28 16008
rect -62 15906 -28 15940
rect -62 15838 -28 15872
rect -62 15770 -28 15804
rect -62 15702 -28 15736
rect -62 15634 -28 15668
rect -62 15566 -28 15600
rect -62 15498 -28 15532
rect -62 15430 -28 15464
rect -62 15362 -28 15396
rect -62 15294 -28 15328
rect -62 15226 -28 15260
rect -62 15158 -28 15192
rect -62 15090 -28 15124
rect -62 15022 -28 15056
rect -62 14954 -28 14988
rect -62 14886 -28 14920
rect -62 14818 -28 14852
rect -62 14750 -28 14784
rect -62 14682 -28 14716
rect -62 14614 -28 14648
rect -62 14546 -28 14580
rect -62 14478 -28 14512
rect -62 14410 -28 14444
rect -62 14342 -28 14376
rect -62 14274 -28 14308
rect -62 14206 -28 14240
rect -62 14138 -28 14172
rect -62 14070 -28 14104
rect -62 14002 -28 14036
rect -62 13934 -28 13968
rect -62 13866 -28 13900
rect -62 13798 -28 13832
rect -62 13730 -28 13764
rect -62 13662 -28 13696
rect -62 13594 -28 13628
rect -62 13526 -28 13560
rect -62 13458 -28 13492
rect -62 13390 -28 13424
rect -62 13322 -28 13356
rect -62 13254 -28 13288
rect -62 13186 -28 13220
rect -62 13118 -28 13152
rect -62 13050 -28 13084
rect -62 12982 -28 13016
rect -62 12914 -28 12948
rect -62 12846 -28 12880
rect -62 12778 -28 12812
rect -62 12710 -28 12744
rect -62 12642 -28 12676
rect -62 12574 -28 12608
rect -62 12506 -28 12540
rect -62 12438 -28 12472
rect -62 12370 -28 12404
rect -62 12302 -28 12336
rect -62 12234 -28 12268
rect -62 12166 -28 12200
rect -62 12098 -28 12132
rect -62 12030 -28 12064
rect -62 11962 -28 11996
rect -62 11894 -28 11928
rect -62 11826 -28 11860
rect -62 11758 -28 11792
rect -62 11690 -28 11724
rect -62 11622 -28 11656
rect -62 11554 -28 11588
rect -62 11486 -28 11520
rect -62 11418 -28 11452
rect -62 11350 -28 11384
rect -62 11282 -28 11316
rect -62 11214 -28 11248
rect -62 11146 -28 11180
rect -62 11078 -28 11112
rect -62 11010 -28 11044
rect -62 10942 -28 10976
rect -62 10874 -28 10908
rect -62 10806 -28 10840
rect -62 10738 -28 10772
rect -62 10670 -28 10704
rect -62 10602 -28 10636
rect -62 10534 -28 10568
rect -62 10466 -28 10500
rect -62 10398 -28 10432
rect -62 10330 -28 10364
rect -62 10262 -28 10296
rect -62 10194 -28 10228
rect -62 10126 -28 10160
rect -62 10058 -28 10092
rect -62 9990 -28 10024
rect -62 9922 -28 9956
rect -62 9854 -28 9888
rect -62 9786 -28 9820
rect -62 9718 -28 9752
rect -62 9650 -28 9684
rect -62 9582 -28 9616
rect -62 9514 -28 9548
rect -62 9446 -28 9480
rect -62 9378 -28 9412
rect -62 9310 -28 9344
rect -62 9242 -28 9276
rect -62 9174 -28 9208
rect -62 9106 -28 9140
rect -62 9038 -28 9072
rect -62 8970 -28 9004
rect -62 8902 -28 8936
rect -62 8834 -28 8868
rect -62 8766 -28 8800
rect -62 8698 -28 8732
rect -62 8630 -28 8664
rect 1258 17074 1292 17108
rect 1258 17006 1292 17040
rect 1258 16938 1292 16972
rect 1258 16870 1292 16904
rect 1258 16802 1292 16836
rect 1258 16734 1292 16768
rect 1258 16666 1292 16700
rect 1258 16598 1292 16632
rect 1258 16530 1292 16564
rect 1258 16462 1292 16496
rect 1258 16394 1292 16428
rect 1258 16326 1292 16360
rect 1258 16258 1292 16292
rect 1258 16190 1292 16224
rect 1258 16122 1292 16156
rect 1258 16054 1292 16088
rect 1258 15986 1292 16020
rect 1258 15918 1292 15952
rect 1258 15850 1292 15884
rect 1258 15782 1292 15816
rect 1258 15714 1292 15748
rect 1258 15646 1292 15680
rect 1258 15578 1292 15612
rect 1258 15510 1292 15544
rect 1258 15442 1292 15476
rect 1258 15374 1292 15408
rect 1258 15306 1292 15340
rect 1258 15238 1292 15272
rect 1258 15170 1292 15204
rect 1258 15102 1292 15136
rect 1258 15034 1292 15068
rect 1258 14966 1292 15000
rect 1258 14898 1292 14932
rect 1258 14830 1292 14864
rect 1258 14762 1292 14796
rect 1258 14694 1292 14728
rect 1258 14626 1292 14660
rect 1258 14558 1292 14592
rect 1258 14490 1292 14524
rect 1258 14422 1292 14456
rect 1258 14354 1292 14388
rect 1258 14286 1292 14320
rect 1258 14218 1292 14252
rect 1258 14150 1292 14184
rect 1258 14082 1292 14116
rect 1258 14014 1292 14048
rect 1258 13946 1292 13980
rect 1258 13878 1292 13912
rect 1258 13810 1292 13844
rect 1258 13742 1292 13776
rect 1258 13674 1292 13708
rect 1258 13606 1292 13640
rect 1258 13538 1292 13572
rect 1258 13470 1292 13504
rect 1258 13402 1292 13436
rect 1258 13334 1292 13368
rect 1258 13266 1292 13300
rect 1258 13198 1292 13232
rect 1258 13130 1292 13164
rect 1258 13062 1292 13096
rect 1258 12994 1292 13028
rect 1258 12926 1292 12960
rect 1258 12858 1292 12892
rect 1258 12790 1292 12824
rect 1258 12722 1292 12756
rect 1258 12654 1292 12688
rect 1258 12586 1292 12620
rect 1258 12518 1292 12552
rect 1258 12450 1292 12484
rect 1258 12382 1292 12416
rect 1258 12314 1292 12348
rect 1258 12246 1292 12280
rect 1258 12178 1292 12212
rect 1258 12110 1292 12144
rect 1258 12042 1292 12076
rect 1258 11974 1292 12008
rect 1258 11906 1292 11940
rect 1258 11838 1292 11872
rect 1258 11770 1292 11804
rect 1258 11702 1292 11736
rect 1258 11634 1292 11668
rect 1258 11566 1292 11600
rect 1258 11498 1292 11532
rect 1258 11430 1292 11464
rect 1258 11362 1292 11396
rect 1258 11294 1292 11328
rect 1258 11226 1292 11260
rect 1258 11158 1292 11192
rect 1258 11090 1292 11124
rect 1258 11022 1292 11056
rect 1258 10954 1292 10988
rect 1258 10886 1292 10920
rect 1258 10818 1292 10852
rect 1258 10750 1292 10784
rect 1258 10682 1292 10716
rect 1258 10614 1292 10648
rect 1258 10546 1292 10580
rect 1258 10478 1292 10512
rect 1258 10410 1292 10444
rect 1258 10342 1292 10376
rect 1258 10274 1292 10308
rect 1258 10206 1292 10240
rect 1258 10138 1292 10172
rect 1258 10070 1292 10104
rect 1258 10002 1292 10036
rect 1258 9934 1292 9968
rect 1258 9866 1292 9900
rect 1258 9798 1292 9832
rect 1258 9730 1292 9764
rect 1258 9662 1292 9696
rect 1258 9594 1292 9628
rect 1258 9526 1292 9560
rect 1258 9458 1292 9492
rect 1258 9390 1292 9424
rect 1258 9322 1292 9356
rect 1258 9254 1292 9288
rect 1258 9186 1292 9220
rect 1258 9118 1292 9152
rect 1258 9050 1292 9084
rect 1258 8982 1292 9016
rect 1258 8914 1292 8948
rect 1258 8846 1292 8880
rect 1258 8778 1292 8812
rect 1258 8710 1292 8744
rect 1258 8642 1292 8676
rect -62 8562 -28 8596
rect -62 8494 -28 8528
rect -62 8426 -28 8460
rect -62 8358 -28 8392
rect -62 8290 -28 8324
rect -62 8222 -28 8256
rect -62 8154 -28 8188
rect -62 8086 -28 8120
rect -62 8018 -28 8052
rect -62 7950 -28 7984
rect -62 7882 -28 7916
rect -62 7814 -28 7848
rect -62 7746 -28 7780
rect -62 7678 -28 7712
rect -62 7610 -28 7644
rect -62 7542 -28 7576
rect -62 7474 -28 7508
rect -62 7406 -28 7440
rect -62 7338 -28 7372
rect -62 7270 -28 7304
rect -62 7202 -28 7236
rect -62 7134 -28 7168
rect -62 7066 -28 7100
rect -62 6998 -28 7032
rect -62 6930 -28 6964
rect -62 6862 -28 6896
rect -62 6794 -28 6828
rect -62 6726 -28 6760
rect -62 6658 -28 6692
rect -62 6590 -28 6624
rect -62 6522 -28 6556
rect -62 6454 -28 6488
rect -62 6386 -28 6420
rect -62 6318 -28 6352
rect -62 6250 -28 6284
rect -62 6182 -28 6216
rect -62 6114 -28 6148
rect -62 6046 -28 6080
rect -62 5978 -28 6012
rect -62 5910 -28 5944
rect -62 5842 -28 5876
rect -62 5774 -28 5808
rect -62 5706 -28 5740
rect -62 5638 -28 5672
rect -62 5570 -28 5604
rect -62 5502 -28 5536
rect -62 5434 -28 5468
rect -62 5366 -28 5400
rect -62 5298 -28 5332
rect -62 5230 -28 5264
rect -62 5162 -28 5196
rect -62 5094 -28 5128
rect -62 5026 -28 5060
rect -62 4958 -28 4992
rect -62 4890 -28 4924
rect -62 4822 -28 4856
rect -62 4754 -28 4788
rect -62 4686 -28 4720
rect -62 4618 -28 4652
rect -62 4550 -28 4584
rect -62 4482 -28 4516
rect -62 4414 -28 4448
rect -62 4346 -28 4380
rect -62 4278 -28 4312
rect -62 4210 -28 4244
rect -62 4142 -28 4176
rect -62 4074 -28 4108
rect -62 4006 -28 4040
rect -62 3938 -28 3972
rect -62 3870 -28 3904
rect -62 3802 -28 3836
rect -62 3734 -28 3768
rect -62 3666 -28 3700
rect -62 3598 -28 3632
rect -62 3530 -28 3564
rect -62 3462 -28 3496
rect -62 3394 -28 3428
rect -62 3326 -28 3360
rect -62 3258 -28 3292
rect -62 3190 -28 3224
rect -62 3122 -28 3156
rect -62 3054 -28 3088
rect -62 2986 -28 3020
rect -62 2918 -28 2952
rect -62 2850 -28 2884
rect -62 2782 -28 2816
rect -62 2714 -28 2748
rect -62 2646 -28 2680
rect -62 2578 -28 2612
rect -62 2510 -28 2544
rect -62 2442 -28 2476
rect -62 2374 -28 2408
rect -62 2306 -28 2340
rect -62 2238 -28 2272
rect -62 2170 -28 2204
rect -62 2102 -28 2136
rect -62 2034 -28 2068
rect -62 1966 -28 2000
rect -62 1898 -28 1932
rect -62 1830 -28 1864
rect -62 1762 -28 1796
rect -62 1694 -28 1728
rect -62 1626 -28 1660
rect -62 1558 -28 1592
rect -62 1490 -28 1524
rect -62 1422 -28 1456
rect -62 1354 -28 1388
rect -62 1286 -28 1320
rect -62 1218 -28 1252
rect -62 1150 -28 1184
rect -62 1082 -28 1116
rect -62 1014 -28 1048
rect -62 946 -28 980
rect -62 878 -28 912
rect -62 810 -28 844
rect -62 742 -28 776
rect -62 674 -28 708
rect -62 606 -28 640
rect -62 538 -28 572
rect -62 470 -28 504
rect -62 402 -28 436
rect -62 334 -28 368
rect -62 266 -28 300
rect -62 198 -28 232
rect -62 130 -28 164
rect -62 62 -28 96
rect 1258 8574 1292 8608
rect 1258 8506 1292 8540
rect 1258 8438 1292 8472
rect 1258 8370 1292 8404
rect 1258 8302 1292 8336
rect 1258 8234 1292 8268
rect 1258 8166 1292 8200
rect 1258 8098 1292 8132
rect 1258 8030 1292 8064
rect 1258 7962 1292 7996
rect 1258 7894 1292 7928
rect 1258 7826 1292 7860
rect 1258 7758 1292 7792
rect 1258 7690 1292 7724
rect 1258 7622 1292 7656
rect 1258 7554 1292 7588
rect 1258 7486 1292 7520
rect 1258 7418 1292 7452
rect 1258 7350 1292 7384
rect 1258 7282 1292 7316
rect 1258 7214 1292 7248
rect 1258 7146 1292 7180
rect 1258 7078 1292 7112
rect 1258 7010 1292 7044
rect 1258 6942 1292 6976
rect 1258 6874 1292 6908
rect 1258 6806 1292 6840
rect 1258 6738 1292 6772
rect 1258 6670 1292 6704
rect 1258 6602 1292 6636
rect 1258 6534 1292 6568
rect 1258 6466 1292 6500
rect 1258 6398 1292 6432
rect 1258 6330 1292 6364
rect 1258 6262 1292 6296
rect 1258 6194 1292 6228
rect 1258 6126 1292 6160
rect 1258 6058 1292 6092
rect 1258 5990 1292 6024
rect 1258 5922 1292 5956
rect 1258 5854 1292 5888
rect 1258 5786 1292 5820
rect 1258 5718 1292 5752
rect 1258 5650 1292 5684
rect 1258 5582 1292 5616
rect 1258 5514 1292 5548
rect 1258 5446 1292 5480
rect 1258 5378 1292 5412
rect 1258 5310 1292 5344
rect 1258 5242 1292 5276
rect 1258 5174 1292 5208
rect 1258 5106 1292 5140
rect 1258 5038 1292 5072
rect 1258 4970 1292 5004
rect 1258 4902 1292 4936
rect 1258 4834 1292 4868
rect 1258 4766 1292 4800
rect 1258 4698 1292 4732
rect 1258 4630 1292 4664
rect 1258 4562 1292 4596
rect 1258 4494 1292 4528
rect 1258 4426 1292 4460
rect 1258 4358 1292 4392
rect 1258 4290 1292 4324
rect 1258 4222 1292 4256
rect 1258 4154 1292 4188
rect 1258 4086 1292 4120
rect 1258 4018 1292 4052
rect 1258 3950 1292 3984
rect 1258 3882 1292 3916
rect 1258 3814 1292 3848
rect 1258 3746 1292 3780
rect 1258 3678 1292 3712
rect 1258 3610 1292 3644
rect 1258 3542 1292 3576
rect 1258 3474 1292 3508
rect 1258 3406 1292 3440
rect 1258 3338 1292 3372
rect 1258 3270 1292 3304
rect 1258 3202 1292 3236
rect 1258 3134 1292 3168
rect 1258 3066 1292 3100
rect 1258 2998 1292 3032
rect 1258 2930 1292 2964
rect 1258 2862 1292 2896
rect 1258 2794 1292 2828
rect 1258 2726 1292 2760
rect 1258 2658 1292 2692
rect 1258 2590 1292 2624
rect 1258 2522 1292 2556
rect 1258 2454 1292 2488
rect 1258 2386 1292 2420
rect 1258 2318 1292 2352
rect 1258 2250 1292 2284
rect 1258 2182 1292 2216
rect 1258 2114 1292 2148
rect 1258 2046 1292 2080
rect 1258 1978 1292 2012
rect 1258 1910 1292 1944
rect 1258 1842 1292 1876
rect 1258 1774 1292 1808
rect 1258 1706 1292 1740
rect 1258 1638 1292 1672
rect 1258 1570 1292 1604
rect 1258 1502 1292 1536
rect 1258 1434 1292 1468
rect 1258 1366 1292 1400
rect 1258 1298 1292 1332
rect 1258 1230 1292 1264
rect 1258 1162 1292 1196
rect 1258 1094 1292 1128
rect 1258 1026 1292 1060
rect 1258 958 1292 992
rect 1258 890 1292 924
rect 1258 822 1292 856
rect 1258 754 1292 788
rect 1258 686 1292 720
rect 1258 618 1292 652
rect 1258 550 1292 584
rect 1258 482 1292 516
rect 1258 414 1292 448
rect 1258 346 1292 380
rect 1258 278 1292 312
rect 1258 210 1292 244
rect 1258 142 1292 176
rect 1258 74 1292 108
rect 1258 6 1292 40
rect 6 -62 40 -28
rect 74 -62 108 -28
rect 142 -62 176 -28
rect 210 -62 244 -28
rect 278 -62 312 -28
rect 346 -62 380 -28
rect 414 -62 448 -28
rect 482 -62 516 -28
rect 550 -62 584 -28
rect 618 -62 652 -28
rect 686 -62 720 -28
rect 754 -62 788 -28
rect 822 -62 856 -28
rect 890 -62 924 -28
rect 958 -62 992 -28
rect 1026 -62 1060 -28
rect 1094 -62 1128 -28
rect 1162 -62 1196 -28
<< locali >>
rect -62 17198 34 17232
rect 68 17198 102 17232
rect 136 17198 170 17232
rect 204 17198 238 17232
rect 272 17198 306 17232
rect 340 17198 374 17232
rect 408 17198 442 17232
rect 476 17198 510 17232
rect 544 17198 578 17232
rect 612 17198 646 17232
rect 680 17198 714 17232
rect 748 17198 782 17232
rect 816 17198 850 17232
rect 884 17198 918 17232
rect 952 17198 986 17232
rect 1020 17198 1054 17232
rect 1088 17198 1122 17232
rect 1156 17198 1190 17232
rect 1224 17198 1292 17232
rect -62 17164 -28 17198
rect 642 17136 742 17198
rect -62 17096 -28 17130
rect 77 17102 136 17136
rect 170 17102 229 17136
rect 385 17102 444 17136
rect 478 17102 537 17136
rect 642 17102 675 17136
rect 709 17102 742 17136
rect -62 17028 -28 17062
rect -62 16960 -28 16994
rect -62 16892 -28 16926
rect -62 16824 -28 16858
rect -62 16756 -28 16790
rect -62 16688 -28 16722
rect -62 16620 -28 16654
rect -62 16552 -28 16586
rect -62 16484 -28 16518
rect -62 16416 -28 16450
rect -62 16348 -28 16382
rect -62 16280 -28 16314
rect -62 16212 -28 16246
rect -62 16144 -28 16178
rect -62 16076 -28 16110
rect -62 16008 -28 16042
rect -62 15940 -28 15974
rect -62 15872 -28 15906
rect -62 15804 -28 15838
rect 642 16834 742 17102
rect 813 17053 1033 17144
rect 1104 17136 1204 17198
rect 1104 17102 1137 17136
rect 1171 17102 1204 17136
rect 642 16800 675 16834
rect 709 16800 742 16834
rect 642 16532 742 16800
rect 642 16498 675 16532
rect 709 16498 742 16532
rect 642 16230 742 16498
rect 642 16196 675 16230
rect 709 16196 742 16230
rect 642 15928 742 16196
rect 642 15894 675 15928
rect 709 15894 742 15928
rect -62 15736 -28 15770
rect 43 15705 109 15775
rect 197 15705 263 15775
rect 351 15705 417 15775
rect 505 15705 571 15775
rect -62 15668 -28 15702
rect -62 15600 -28 15634
rect -62 15532 -28 15566
rect -62 15464 -28 15498
rect -62 15396 -28 15430
rect -62 15328 -28 15362
rect -62 15260 -28 15294
rect -62 15192 -28 15226
rect -62 15124 -28 15158
rect -62 15056 -28 15090
rect -62 14988 -28 15022
rect -62 14920 -28 14954
rect -62 14852 -28 14886
rect -62 14784 -28 14818
rect -62 14716 -28 14750
rect -62 14648 -28 14682
rect -62 14580 -28 14614
rect -62 14512 -28 14546
rect -62 14444 -28 14478
rect -62 14376 -28 14410
rect 642 15626 742 15894
rect 1104 16834 1204 17102
rect 1104 16800 1137 16834
rect 1171 16800 1204 16834
rect 1104 16532 1204 16800
rect 1104 16498 1137 16532
rect 1171 16498 1204 16532
rect 1104 16230 1204 16498
rect 1104 16196 1137 16230
rect 1171 16196 1204 16230
rect 1104 15928 1204 16196
rect 1104 15894 1137 15928
rect 1171 15894 1204 15928
rect 813 15705 879 15775
rect 967 15705 1033 15775
rect 642 15592 675 15626
rect 709 15592 742 15626
rect 642 15324 742 15592
rect 642 15290 675 15324
rect 709 15290 742 15324
rect 642 15022 742 15290
rect 642 14988 675 15022
rect 709 14988 742 15022
rect 642 14720 742 14988
rect 642 14686 675 14720
rect 709 14686 742 14720
rect 642 14418 742 14686
rect 642 14384 675 14418
rect 709 14384 742 14418
rect -62 14308 -28 14342
rect 43 14274 109 14344
rect 197 14274 263 14344
rect 351 14274 417 14344
rect 505 14343 521 14344
rect 555 14343 571 14344
rect 505 14275 571 14343
rect 505 14274 521 14275
rect -62 14240 -28 14274
rect 555 14274 571 14275
rect -62 14172 -28 14206
rect -62 14104 -28 14138
rect -62 14036 -28 14070
rect -62 13968 -28 14002
rect -62 13900 -28 13934
rect -62 13832 -28 13866
rect -62 13764 -28 13798
rect -62 13696 -28 13730
rect -62 13628 -28 13662
rect -62 13560 -28 13594
rect -62 13492 -28 13526
rect -62 13424 -28 13458
rect -62 13356 -28 13390
rect -62 13288 -28 13322
rect -62 13220 -28 13254
rect -62 13152 -28 13186
rect -62 13084 -28 13118
rect 642 14116 742 14384
rect 1104 15626 1204 15894
rect 1104 15592 1137 15626
rect 1171 15592 1204 15626
rect 1104 15324 1204 15592
rect 1104 15290 1137 15324
rect 1171 15290 1204 15324
rect 1104 15022 1204 15290
rect 1104 14988 1137 15022
rect 1171 14988 1204 15022
rect 1104 14720 1204 14988
rect 1104 14686 1137 14720
rect 1171 14686 1204 14720
rect 1104 14418 1204 14686
rect 1104 14384 1137 14418
rect 1171 14384 1204 14418
rect 813 14274 879 14344
rect 967 14274 1033 14344
rect 980 14240 1018 14274
rect 642 14082 675 14116
rect 709 14082 742 14116
rect 642 13814 742 14082
rect 642 13780 675 13814
rect 709 13780 742 13814
rect 642 13512 742 13780
rect 642 13478 675 13512
rect 709 13478 742 13512
rect 642 13210 742 13478
rect 642 13176 675 13210
rect 709 13176 742 13210
rect 642 13058 742 13176
rect 1104 14116 1204 14384
rect 1104 14082 1137 14116
rect 1171 14082 1204 14116
rect 1104 13814 1204 14082
rect 1104 13780 1137 13814
rect 1171 13780 1204 13814
rect 1104 13512 1204 13780
rect 1104 13478 1137 13512
rect 1171 13478 1204 13512
rect 1104 13210 1204 13478
rect 1104 13176 1137 13210
rect 1171 13176 1204 13210
rect -62 13016 -28 13050
rect -62 12948 -28 12982
rect -62 12880 -28 12914
rect -62 12812 -28 12846
rect 43 12843 109 12913
rect 197 12843 263 12913
rect 351 12843 417 12913
rect 488 12877 588 12947
rect 813 12896 827 12913
rect 861 12896 879 12913
rect 488 12786 742 12877
rect 813 12858 879 12896
rect 813 12843 827 12858
rect 861 12843 879 12858
rect 967 12843 1033 12913
rect 1104 12908 1204 13176
rect 1104 12874 1137 12908
rect 1171 12874 1204 12908
rect -62 12744 -28 12778
rect -62 12676 -28 12710
rect -62 12608 -28 12642
rect -62 12540 -28 12574
rect -62 12472 -28 12506
rect -62 12404 -28 12438
rect -62 12336 -28 12370
rect -62 12268 -28 12302
rect -62 12200 -28 12234
rect -62 12132 -28 12166
rect -62 12064 -28 12098
rect -62 11996 -28 12030
rect -62 11928 -28 11962
rect -62 11860 -28 11894
rect -62 11792 -28 11826
rect -62 11724 -28 11758
rect -62 11656 -28 11690
rect -62 11588 -28 11622
rect -62 11520 -28 11554
rect 1104 12606 1204 12874
rect 1104 12572 1137 12606
rect 1171 12572 1204 12606
rect 1104 12304 1204 12572
rect 1104 12270 1137 12304
rect 1171 12270 1204 12304
rect 1104 12002 1204 12270
rect 1104 11968 1137 12002
rect 1171 11968 1204 12002
rect 1104 11700 1204 11968
rect 1104 11666 1137 11700
rect 1171 11666 1204 11700
rect -62 11452 -28 11486
rect -62 11384 -28 11418
rect 43 11412 109 11482
rect 197 11412 263 11482
rect 368 11431 402 11469
rect 488 11464 742 11516
rect 488 11430 559 11464
rect 593 11430 631 11464
rect 665 11430 742 11464
rect 488 11378 742 11430
rect 813 11412 879 11482
rect 967 11412 1033 11482
rect 1104 11398 1204 11666
rect -62 11316 -28 11350
rect -62 11248 -28 11282
rect -62 11180 -28 11214
rect -62 11112 -28 11146
rect -62 11044 -28 11078
rect -62 10976 -28 11010
rect -62 10908 -28 10942
rect -62 10840 -28 10874
rect -62 10772 -28 10806
rect -62 10704 -28 10738
rect -62 10636 -28 10670
rect -62 10568 -28 10602
rect -62 10500 -28 10534
rect -62 10432 -28 10466
rect -62 10364 -28 10398
rect -62 10296 -28 10330
rect -62 10228 -28 10262
rect -62 10160 -28 10194
rect -62 10092 -28 10126
rect 1104 11364 1137 11398
rect 1171 11364 1204 11398
rect 1104 11096 1204 11364
rect 1104 11062 1137 11096
rect 1171 11062 1204 11096
rect 1104 10794 1204 11062
rect 1104 10760 1137 10794
rect 1171 10760 1204 10794
rect 1104 10492 1204 10760
rect 1104 10458 1137 10492
rect 1171 10458 1204 10492
rect 1104 10190 1204 10458
rect 1104 10156 1137 10190
rect 1171 10156 1204 10190
rect -62 10024 -28 10058
rect -62 9956 -28 9990
rect 43 9981 109 10051
rect 197 9981 263 10051
rect 351 9981 417 10051
rect 488 10043 742 10093
rect 488 9947 588 10043
rect -62 9888 -28 9922
rect -62 9820 -28 9854
rect -62 9752 -28 9786
rect -62 9684 -28 9718
rect -62 9616 -28 9650
rect 642 9586 742 9989
rect 813 9981 879 10051
rect 967 9981 1033 10051
rect -62 9548 -28 9582
rect -62 9480 -28 9514
rect -62 9412 -28 9446
rect -62 9344 -28 9378
rect -62 9276 -28 9310
rect -62 9208 -28 9242
rect -62 9140 -28 9174
rect -62 9072 -28 9106
rect -62 9004 -28 9038
rect -62 8936 -28 8970
rect -62 8868 -28 8902
rect -62 8800 -28 8834
rect -62 8732 -28 8766
rect -62 8664 -28 8698
rect 488 9497 742 9586
rect 1104 9888 1204 10156
rect 1104 9854 1137 9888
rect 1171 9854 1204 9888
rect 1104 9586 1204 9854
rect 1104 9552 1137 9586
rect 1171 9552 1204 9586
rect -62 8596 -28 8630
rect 212 8620 250 8654
rect -62 8528 -28 8562
rect 43 8550 109 8620
rect 197 8550 263 8620
rect 330 8558 434 8680
rect 488 8612 588 9497
rect 1104 9284 1204 9552
rect 1104 9250 1137 9284
rect 1171 9250 1204 9284
rect 1104 8982 1204 9250
rect 1104 8948 1137 8982
rect 1171 8948 1204 8982
rect 1104 8771 1204 8948
rect 1258 17108 1292 17198
rect 1258 17040 1292 17074
rect 1258 16972 1292 17006
rect 1258 16904 1292 16938
rect 1258 16836 1292 16870
rect 1258 16768 1292 16802
rect 1258 16700 1292 16734
rect 1258 16632 1292 16666
rect 1258 16564 1292 16598
rect 1258 16496 1292 16530
rect 1258 16428 1292 16462
rect 1258 16360 1292 16394
rect 1258 16292 1292 16326
rect 1258 16224 1292 16258
rect 1258 16156 1292 16190
rect 1258 16088 1292 16122
rect 1258 16020 1292 16054
rect 1258 15952 1292 15986
rect 1258 15884 1292 15918
rect 1258 15816 1292 15850
rect 1258 15748 1292 15782
rect 1258 15680 1292 15714
rect 1258 15612 1292 15646
rect 1258 15544 1292 15578
rect 1258 15476 1292 15510
rect 1258 15408 1292 15442
rect 1258 15340 1292 15374
rect 1258 15272 1292 15306
rect 1258 15204 1292 15238
rect 1258 15136 1292 15170
rect 1258 15068 1292 15102
rect 1258 15000 1292 15034
rect 1258 14932 1292 14966
rect 1258 14864 1292 14898
rect 1258 14796 1292 14830
rect 1258 14728 1292 14762
rect 1258 14660 1292 14694
rect 1258 14592 1292 14626
rect 1258 14524 1292 14558
rect 1258 14456 1292 14490
rect 1258 14388 1292 14422
rect 1258 14320 1292 14354
rect 1258 14252 1292 14286
rect 1258 14184 1292 14218
rect 1258 14116 1292 14150
rect 1258 14048 1292 14082
rect 1258 13980 1292 14014
rect 1258 13912 1292 13946
rect 1258 13844 1292 13878
rect 1258 13776 1292 13810
rect 1258 13708 1292 13742
rect 1258 13640 1292 13674
rect 1258 13572 1292 13606
rect 1258 13504 1292 13538
rect 1258 13436 1292 13470
rect 1258 13368 1292 13402
rect 1258 13300 1292 13334
rect 1258 13232 1292 13266
rect 1258 13164 1292 13198
rect 1258 13096 1292 13130
rect 1258 13028 1292 13062
rect 1258 12960 1292 12994
rect 1258 12892 1292 12926
rect 1258 12824 1292 12858
rect 1258 12756 1292 12790
rect 1258 12688 1292 12722
rect 1258 12620 1292 12654
rect 1258 12552 1292 12586
rect 1258 12484 1292 12518
rect 1258 12416 1292 12450
rect 1258 12348 1292 12382
rect 1258 12280 1292 12314
rect 1258 12212 1292 12246
rect 1258 12144 1292 12178
rect 1258 12076 1292 12110
rect 1258 12008 1292 12042
rect 1258 11940 1292 11974
rect 1258 11872 1292 11906
rect 1258 11804 1292 11838
rect 1258 11736 1292 11770
rect 1258 11668 1292 11702
rect 1258 11600 1292 11634
rect 1258 11532 1292 11566
rect 1258 11464 1292 11498
rect 1258 11396 1292 11430
rect 1258 11328 1292 11362
rect 1258 11260 1292 11294
rect 1258 11192 1292 11226
rect 1258 11124 1292 11158
rect 1258 11056 1292 11090
rect 1258 10988 1292 11022
rect 1258 10920 1292 10954
rect 1258 10852 1292 10886
rect 1258 10784 1292 10818
rect 1258 10716 1292 10750
rect 1258 10648 1292 10682
rect 1258 10580 1292 10614
rect 1258 10512 1292 10546
rect 1258 10444 1292 10478
rect 1258 10376 1292 10410
rect 1258 10308 1292 10342
rect 1258 10240 1292 10274
rect 1258 10172 1292 10206
rect 1258 10104 1292 10138
rect 1258 10036 1292 10070
rect 1258 9968 1292 10002
rect 1258 9900 1292 9934
rect 1258 9832 1292 9866
rect 1258 9764 1292 9798
rect 1258 9696 1292 9730
rect 1258 9628 1292 9662
rect 1258 9560 1292 9594
rect 1258 9492 1292 9526
rect 1258 9424 1292 9458
rect 1258 9356 1292 9390
rect 1258 9288 1292 9322
rect 1258 9220 1292 9254
rect 1258 9152 1292 9186
rect 1258 9084 1292 9118
rect 1258 9016 1292 9050
rect 1258 8948 1292 8982
rect 1258 8880 1292 8914
rect 1258 8812 1292 8846
rect 1258 8744 1292 8778
rect 1258 8676 1292 8710
rect -62 8460 -28 8494
rect 330 8481 588 8558
rect 659 8550 725 8620
rect 813 8550 879 8620
rect 967 8550 1033 8620
rect 1258 8608 1292 8642
rect 1132 8516 1170 8550
rect 1258 8540 1292 8574
rect -62 8392 -28 8426
rect -62 8324 -28 8358
rect -62 8256 -28 8290
rect -62 8188 -28 8222
rect -62 8120 -28 8154
rect -62 8052 -28 8086
rect -62 7984 -28 8018
rect -62 7916 -28 7950
rect -62 7848 -28 7882
rect -62 7780 -28 7814
rect -62 7712 -28 7746
rect -62 7644 -28 7678
rect -62 7576 -28 7610
rect -62 7508 -28 7542
rect -62 7440 -28 7474
rect -62 7372 -28 7406
rect -62 7304 -28 7338
rect -62 7236 -28 7270
rect 1258 8472 1292 8506
rect 1258 8404 1292 8438
rect 1258 8336 1292 8370
rect 1258 8268 1292 8302
rect 1258 8200 1292 8234
rect 1258 8132 1292 8166
rect 1258 8064 1292 8098
rect 1258 7996 1292 8030
rect 1258 7928 1292 7962
rect 1258 7860 1292 7894
rect 1258 7792 1292 7826
rect 1258 7724 1292 7758
rect 1258 7656 1292 7690
rect 1258 7588 1292 7622
rect 1258 7520 1292 7554
rect 1258 7452 1292 7486
rect 1258 7384 1292 7418
rect 1258 7316 1292 7350
rect -62 7168 -28 7202
rect -62 7100 -28 7134
rect 43 7119 109 7189
rect 197 7119 263 7189
rect 351 7143 571 7223
rect 659 7181 879 7249
rect 1258 7248 1292 7282
rect -62 7032 -28 7066
rect 351 7024 879 7143
rect 967 7119 1033 7189
rect 1121 7119 1187 7189
rect 1258 7180 1292 7214
rect 1258 7112 1292 7146
rect 1258 7044 1292 7078
rect -62 6964 -28 6998
rect -62 6896 -28 6930
rect -62 6828 -28 6862
rect -62 6760 -28 6794
rect -62 6692 -28 6726
rect -62 6624 -28 6658
rect -62 6556 -28 6590
rect -62 6488 -28 6522
rect -62 6420 -28 6454
rect -62 6352 -28 6386
rect -62 6284 -28 6318
rect -62 6216 -28 6250
rect -62 6148 -28 6182
rect -62 6080 -28 6114
rect -62 6012 -28 6046
rect -62 5944 -28 5978
rect -62 5876 -28 5910
rect -62 5808 -28 5842
rect 1258 6976 1292 7010
rect 1258 6908 1292 6942
rect 1258 6840 1292 6874
rect 1258 6772 1292 6806
rect 1258 6704 1292 6738
rect 1258 6636 1292 6670
rect 1258 6568 1292 6602
rect 1258 6500 1292 6534
rect 1258 6432 1292 6466
rect 1258 6364 1292 6398
rect 1258 6296 1292 6330
rect 1258 6228 1292 6262
rect 1258 6160 1292 6194
rect 1258 6092 1292 6126
rect 1258 6024 1292 6058
rect 1258 5956 1292 5990
rect 1258 5888 1292 5922
rect 1258 5820 1292 5854
rect -62 5740 -28 5774
rect -62 5672 -28 5706
rect 43 5688 109 5758
rect 197 5688 263 5758
rect 351 5739 879 5792
rect 351 5705 379 5739
rect 413 5705 451 5739
rect 485 5705 879 5739
rect 351 5654 879 5705
rect 967 5688 1033 5758
rect 1121 5688 1187 5758
rect 1258 5752 1292 5786
rect 1258 5684 1292 5718
rect -62 5604 -28 5638
rect -62 5536 -28 5570
rect -62 5468 -28 5502
rect -62 5400 -28 5434
rect -62 5332 -28 5366
rect -62 5264 -28 5298
rect -62 5196 -28 5230
rect -62 5128 -28 5162
rect -62 5060 -28 5094
rect -62 4992 -28 5026
rect -62 4924 -28 4958
rect -62 4856 -28 4890
rect -62 4788 -28 4822
rect -62 4720 -28 4754
rect -62 4652 -28 4686
rect -62 4584 -28 4618
rect -62 4516 -28 4550
rect -62 4448 -28 4482
rect 1258 5616 1292 5650
rect 1258 5548 1292 5582
rect 1258 5480 1292 5514
rect 1258 5412 1292 5446
rect 1258 5344 1292 5378
rect 1258 5276 1292 5310
rect 1258 5208 1292 5242
rect 1258 5140 1292 5174
rect 1258 5072 1292 5106
rect 1258 5004 1292 5038
rect 1258 4936 1292 4970
rect 1258 4868 1292 4902
rect 1258 4800 1292 4834
rect 1258 4732 1292 4766
rect 1258 4664 1292 4698
rect 1258 4596 1292 4630
rect 1258 4528 1292 4562
rect 1258 4460 1292 4494
rect -62 4380 -28 4414
rect -62 4312 -28 4346
rect -62 4244 -28 4278
rect 43 4257 109 4327
rect 197 4257 263 4327
rect 334 4301 879 4426
rect 1258 4392 1292 4426
rect 977 4327 1015 4361
rect 1121 4313 1138 4327
rect 1172 4313 1187 4327
rect 334 4213 434 4301
rect 1121 4275 1187 4313
rect -62 4176 -28 4210
rect 505 4163 725 4265
rect 813 4163 1033 4265
rect 1121 4257 1138 4275
rect 1172 4257 1187 4275
rect 1258 4324 1292 4358
rect 1258 4256 1292 4290
rect 1258 4188 1292 4222
rect -62 4108 -28 4142
rect -62 4040 -28 4074
rect -62 3972 -28 4006
rect -62 3904 -28 3938
rect -62 3836 -28 3870
rect -62 3768 -28 3802
rect -62 3700 -28 3734
rect -62 3632 -28 3666
rect -62 3564 -28 3598
rect -62 3496 -28 3530
rect -62 3428 -28 3462
rect -62 3360 -28 3394
rect -62 3292 -28 3326
rect -62 3224 -28 3258
rect -62 3156 -28 3190
rect -62 3088 -28 3122
rect -62 3020 -28 3054
rect -62 2952 -28 2986
rect -62 2884 -28 2918
rect 1258 4120 1292 4154
rect 1258 4052 1292 4086
rect 1258 3984 1292 4018
rect 1258 3916 1292 3950
rect 1258 3848 1292 3882
rect 1258 3780 1292 3814
rect 1258 3712 1292 3746
rect 1258 3644 1292 3678
rect 1258 3576 1292 3610
rect 1258 3508 1292 3542
rect 1258 3440 1292 3474
rect 1258 3372 1292 3406
rect 1258 3304 1292 3338
rect 1258 3236 1292 3270
rect 1258 3168 1292 3202
rect 1258 3100 1292 3134
rect 1258 3032 1292 3066
rect 1258 2964 1292 2998
rect 1258 2896 1292 2930
rect -62 2816 -28 2850
rect 43 2826 109 2896
rect 197 2826 263 2896
rect 351 2826 417 2896
rect 505 2826 571 2896
rect 659 2826 725 2896
rect 813 2826 879 2896
rect 967 2826 1033 2896
rect 1121 2826 1187 2896
rect 1258 2828 1292 2862
rect -62 2748 -28 2782
rect -62 2680 -28 2714
rect -62 2612 -28 2646
rect -62 2544 -28 2578
rect -62 2476 -28 2510
rect -62 2408 -28 2442
rect -62 2340 -28 2374
rect -62 2272 -28 2306
rect -62 2204 -28 2238
rect -62 2136 -28 2170
rect -62 2068 -28 2102
rect -62 2000 -28 2034
rect -62 1932 -28 1966
rect -62 1864 -28 1898
rect -62 1796 -28 1830
rect -62 1728 -28 1762
rect -62 1660 -28 1694
rect -62 1592 -28 1626
rect -62 1524 -28 1558
rect -62 1456 -28 1490
rect 1258 2760 1292 2794
rect 1258 2692 1292 2726
rect 1258 2624 1292 2658
rect 1258 2556 1292 2590
rect 1258 2488 1292 2522
rect 1258 2420 1292 2454
rect 1258 2352 1292 2386
rect 1258 2284 1292 2318
rect 1258 2216 1292 2250
rect 1258 2148 1292 2182
rect 1258 2080 1292 2114
rect 1258 2012 1292 2046
rect 1258 1944 1292 1978
rect 1258 1876 1292 1910
rect 1258 1808 1292 1842
rect 1258 1740 1292 1774
rect 1258 1672 1292 1706
rect 1258 1604 1292 1638
rect 1258 1536 1292 1570
rect 1258 1468 1292 1502
rect -62 1388 -28 1422
rect 43 1395 109 1465
rect 197 1395 263 1465
rect 351 1395 417 1465
rect 505 1395 571 1465
rect 659 1395 725 1465
rect 813 1395 879 1465
rect 967 1395 1033 1465
rect 1121 1395 1187 1465
rect 1258 1400 1292 1434
rect -62 1320 -28 1354
rect -62 1252 -28 1286
rect -62 1184 -28 1218
rect -62 1116 -28 1150
rect -62 1048 -28 1082
rect -62 980 -28 1014
rect -62 912 -28 946
rect -62 844 -28 878
rect -62 776 -28 810
rect -62 708 -28 742
rect -62 640 -28 674
rect -62 572 -28 606
rect -62 504 -28 538
rect -62 436 -28 470
rect -62 368 -28 402
rect -62 300 -28 334
rect -62 232 -28 266
rect -62 164 -28 198
rect -62 96 -28 130
rect 1258 1332 1292 1366
rect 1258 1264 1292 1298
rect 1258 1196 1292 1230
rect 1258 1128 1292 1162
rect 1258 1060 1292 1094
rect 1258 992 1292 1026
rect 1258 924 1292 958
rect 1258 856 1292 890
rect 1258 788 1292 822
rect 1258 720 1292 754
rect 1258 652 1292 686
rect 1258 584 1292 618
rect 1258 516 1292 550
rect 1258 448 1292 482
rect 1258 380 1292 414
rect 1258 312 1292 346
rect 1258 244 1292 278
rect 1258 176 1292 210
rect -62 -28 -28 62
rect 54 34 92 68
rect 231 34 290 68
rect 324 34 383 68
rect 518 34 556 68
rect 659 22 879 124
rect 967 21 1187 123
rect 1258 108 1292 142
rect 1258 40 1292 74
rect 1258 -28 1292 6
rect -62 -62 6 -28
rect 40 -62 74 -28
rect 108 -62 142 -28
rect 176 -62 210 -28
rect 244 -62 278 -28
rect 312 -62 346 -28
rect 380 -62 414 -28
rect 448 -62 482 -28
rect 516 -62 550 -28
rect 584 -62 618 -28
rect 652 -62 686 -28
rect 720 -62 754 -28
rect 788 -62 822 -28
rect 856 -62 890 -28
rect 924 -62 958 -28
rect 992 -62 1026 -28
rect 1060 -62 1094 -28
rect 1128 -62 1162 -28
rect 1196 -62 1292 -28
<< viali >>
rect 43 17102 77 17136
rect 136 17102 170 17136
rect 229 17102 263 17136
rect 351 17102 385 17136
rect 444 17102 478 17136
rect 537 17102 571 17136
rect 521 14343 555 14377
rect 521 14241 555 14275
rect 946 14240 980 14274
rect 1018 14240 1052 14274
rect 827 12896 861 12930
rect 827 12824 861 12858
rect 368 11469 402 11503
rect 368 11397 402 11431
rect 559 11430 593 11464
rect 631 11430 665 11464
rect 178 8620 212 8654
rect 250 8620 284 8654
rect 1098 8516 1132 8550
rect 1170 8516 1204 8550
rect 379 5705 413 5739
rect 451 5705 485 5739
rect 943 4327 977 4361
rect 1015 4327 1049 4361
rect 1138 4313 1172 4347
rect 1138 4241 1172 4275
rect 20 34 54 68
rect 92 34 126 68
rect 197 34 231 68
rect 290 34 324 68
rect 383 34 417 68
rect 484 34 518 68
rect 556 34 590 68
<< metal1 >>
rect 31 17136 275 17142
rect 31 17102 43 17136
rect 77 17102 136 17136
rect 170 17102 229 17136
rect 263 17102 275 17136
rect 31 17096 275 17102
rect 339 17136 583 17142
rect 339 17102 351 17136
rect 385 17102 444 17136
rect 478 17102 537 17136
rect 571 17102 583 17136
rect 339 17096 583 17102
rect 515 14377 561 14389
rect 515 14343 521 14377
rect 555 14343 561 14377
rect 515 14275 561 14343
rect 515 14241 521 14275
rect 555 14241 561 14275
rect 515 14229 561 14241
rect 934 14274 1064 14280
rect 934 14240 946 14274
rect 980 14240 1018 14274
rect 1052 14240 1064 14274
rect 934 14234 1064 14240
rect 821 12930 867 12942
rect 821 12896 827 12930
rect 861 12896 867 12930
rect 821 12858 867 12896
rect 821 12824 827 12858
rect 861 12824 867 12858
rect 821 12812 867 12824
rect 362 11503 408 11515
rect 362 11469 368 11503
rect 402 11469 408 11503
rect 362 11431 408 11469
rect 362 11397 368 11431
rect 402 11397 408 11431
rect 547 11464 677 11470
rect 547 11430 559 11464
rect 593 11430 631 11464
rect 665 11430 677 11464
rect 547 11424 677 11430
rect 362 11385 408 11397
rect 166 8654 296 8660
rect 166 8620 178 8654
rect 212 8620 250 8654
rect 284 8620 296 8654
rect 166 8614 296 8620
rect 977 8550 1216 8556
rect 977 8516 1098 8550
rect 1132 8516 1170 8550
rect 1204 8516 1216 8550
rect 977 8510 1216 8516
rect 367 5739 497 5745
rect 367 5705 379 5739
rect 413 5705 451 5739
rect 485 5705 497 5739
rect 367 5699 497 5705
rect 977 4367 1023 8510
rect 931 4361 1061 4367
rect 931 4327 943 4361
rect 977 4327 1015 4361
rect 1049 4327 1061 4361
rect 931 4321 1061 4327
rect 1132 4347 1178 4359
rect 1132 4313 1138 4347
rect 1172 4313 1178 4347
rect 1132 4275 1178 4313
rect 1132 4241 1138 4275
rect 1172 4241 1178 4275
rect 1132 4229 1178 4241
rect 472 117 602 158
rect 8 68 138 74
rect 8 34 20 68
rect 54 34 92 68
rect 126 34 138 68
rect 8 28 138 34
rect 185 68 429 74
rect 185 34 197 68
rect 231 34 290 68
rect 324 34 383 68
rect 417 34 429 68
rect 185 28 429 34
rect 472 68 602 115
rect 472 34 484 68
rect 518 34 556 68
rect 590 34 602 68
rect 472 28 602 34
<< rmetal1 >>
rect 472 115 602 117
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_0
timestamp 1707688321
transform 0 1 1125 -1 0 8990
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_1
timestamp 1707688321
transform 0 1 1125 -1 0 9896
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_2
timestamp 1707688321
transform 0 1 1125 -1 0 9594
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_3
timestamp 1707688321
transform 0 1 1125 -1 0 9292
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_4
timestamp 1707688321
transform 0 1 1125 -1 0 10198
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_5
timestamp 1707688321
transform 0 1 1125 -1 0 10500
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_6
timestamp 1707688321
transform 0 1 1125 -1 0 10802
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_7
timestamp 1707688321
transform 0 1 1125 -1 0 11104
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_8
timestamp 1707688321
transform 0 1 1125 -1 0 11406
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_9
timestamp 1707688321
transform 0 1 1125 -1 0 11708
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_10
timestamp 1707688321
transform 0 1 1125 -1 0 12010
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_11
timestamp 1707688321
transform 0 1 1125 -1 0 12312
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_12
timestamp 1707688321
transform 0 1 1125 -1 0 12614
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_13
timestamp 1707688321
transform 0 1 1125 -1 0 12916
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_14
timestamp 1707688321
transform 0 1 1125 -1 0 17144
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_15
timestamp 1707688321
transform 0 1 1125 -1 0 16842
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_16
timestamp 1707688321
transform 0 1 1125 -1 0 16540
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_17
timestamp 1707688321
transform 0 1 1125 -1 0 16238
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_18
timestamp 1707688321
transform 0 1 1125 -1 0 15936
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_19
timestamp 1707688321
transform 0 1 1125 -1 0 15634
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_20
timestamp 1707688321
transform 0 1 1125 -1 0 15332
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_21
timestamp 1707688321
transform 0 1 1125 -1 0 15030
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_22
timestamp 1707688321
transform 0 1 1125 -1 0 14728
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_23
timestamp 1707688321
transform 0 1 1125 -1 0 14426
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_24
timestamp 1707688321
transform 0 1 1125 -1 0 14124
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_25
timestamp 1707688321
transform 0 1 1125 -1 0 13218
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_26
timestamp 1707688321
transform 0 1 1125 -1 0 13520
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_27
timestamp 1707688321
transform 0 1 1125 -1 0 13822
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_28
timestamp 1707688321
transform 0 1 663 -1 0 13822
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_29
timestamp 1707688321
transform 0 1 663 -1 0 13520
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_30
timestamp 1707688321
transform 0 1 663 -1 0 13218
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_31
timestamp 1707688321
transform 0 1 663 -1 0 14124
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_32
timestamp 1707688321
transform 0 1 663 -1 0 14426
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_33
timestamp 1707688321
transform 0 1 663 -1 0 17144
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_34
timestamp 1707688321
transform 0 1 663 -1 0 16842
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_35
timestamp 1707688321
transform 0 1 663 -1 0 16540
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_36
timestamp 1707688321
transform 0 1 663 -1 0 15936
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_37
timestamp 1707688321
transform 0 1 663 -1 0 14728
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_38
timestamp 1707688321
transform 0 1 663 -1 0 15030
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_39
timestamp 1707688321
transform 0 1 663 -1 0 16238
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_40
timestamp 1707688321
transform 0 1 663 -1 0 15332
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_41
timestamp 1707688321
transform 0 1 663 -1 0 15634
box 0 0 1 1
use M1short_CDNS_524688791851141  M1short_CDNS_524688791851141_0
timestamp 1707688321
transform 0 -1 602 -1 0 130
box 0 0 1 1
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_0
timestamp 1707688321
transform 0 -1 126 1 0 68
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_1
timestamp 1707688321
transform 0 -1 126 1 0 1499
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_2
timestamp 1707688321
transform 0 -1 126 1 0 2930
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_3
timestamp 1707688321
transform 0 -1 126 1 0 4361
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_4
timestamp 1707688321
transform 0 -1 126 1 0 5792
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_5
timestamp 1707688321
transform 0 -1 126 1 0 7223
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_6
timestamp 1707688321
transform 0 -1 126 1 0 8654
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_7
timestamp 1707688321
transform 0 -1 126 1 0 10085
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_8
timestamp 1707688321
transform 0 -1 126 1 0 11516
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_9
timestamp 1707688321
transform 0 -1 126 1 0 12947
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_10
timestamp 1707688321
transform 0 -1 126 1 0 14378
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_11
timestamp 1707688321
transform 0 -1 126 1 0 15809
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_12
timestamp 1707688321
transform 0 -1 280 1 0 15809
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_13
timestamp 1707688321
transform 0 -1 280 1 0 14378
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_14
timestamp 1707688321
transform 0 -1 280 1 0 12947
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_15
timestamp 1707688321
transform 0 -1 280 1 0 11516
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_16
timestamp 1707688321
transform 0 -1 280 1 0 10085
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_17
timestamp 1707688321
transform 0 -1 280 1 0 68
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_18
timestamp 1707688321
transform 0 -1 280 1 0 1499
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_19
timestamp 1707688321
transform 0 -1 280 1 0 2930
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_20
timestamp 1707688321
transform 0 -1 280 1 0 4361
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_21
timestamp 1707688321
transform 0 -1 280 1 0 5792
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_22
timestamp 1707688321
transform 0 -1 280 1 0 7223
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_23
timestamp 1707688321
transform 0 -1 280 1 0 8654
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_24
timestamp 1707688321
transform 0 -1 588 1 0 8654
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_25
timestamp 1707688321
transform 0 -1 588 1 0 7223
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_26
timestamp 1707688321
transform 0 -1 588 1 0 5792
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_27
timestamp 1707688321
transform 0 -1 588 1 0 4361
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_28
timestamp 1707688321
transform 0 -1 588 1 0 2930
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_29
timestamp 1707688321
transform 0 -1 588 1 0 1499
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_30
timestamp 1707688321
transform 0 -1 588 1 0 68
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_31
timestamp 1707688321
transform 0 -1 588 1 0 10085
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_32
timestamp 1707688321
transform 0 -1 588 1 0 11516
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_33
timestamp 1707688321
transform 0 -1 588 1 0 12947
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_34
timestamp 1707688321
transform 0 -1 588 1 0 14378
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_35
timestamp 1707688321
transform 0 -1 588 1 0 15809
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_36
timestamp 1707688321
transform 0 -1 434 1 0 15809
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_37
timestamp 1707688321
transform 0 -1 434 1 0 14378
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_38
timestamp 1707688321
transform 0 -1 434 1 0 12947
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_39
timestamp 1707688321
transform 0 -1 434 1 0 11516
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_40
timestamp 1707688321
transform 0 -1 434 1 0 10085
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_41
timestamp 1707688321
transform 0 -1 434 1 0 68
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_42
timestamp 1707688321
transform 0 -1 434 1 0 1499
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_43
timestamp 1707688321
transform 0 -1 434 1 0 2930
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_44
timestamp 1707688321
transform 0 -1 434 1 0 4361
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_45
timestamp 1707688321
transform 0 -1 434 1 0 5792
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_46
timestamp 1707688321
transform 0 -1 434 1 0 7223
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_47
timestamp 1707688321
transform 0 -1 434 1 0 8654
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_48
timestamp 1707688321
transform 0 -1 1050 1 0 8654
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_49
timestamp 1707688321
transform 0 -1 1050 1 0 7223
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_50
timestamp 1707688321
transform 0 -1 1050 1 0 5792
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_51
timestamp 1707688321
transform 0 -1 1050 1 0 4361
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_52
timestamp 1707688321
transform 0 -1 1050 1 0 2930
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_53
timestamp 1707688321
transform 0 -1 1050 1 0 1499
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_54
timestamp 1707688321
transform 0 -1 1050 1 0 68
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_55
timestamp 1707688321
transform 0 -1 1050 1 0 10085
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_56
timestamp 1707688321
transform 0 -1 1050 1 0 11516
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_57
timestamp 1707688321
transform 0 -1 1050 1 0 12947
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_58
timestamp 1707688321
transform 0 -1 1050 1 0 14378
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_59
timestamp 1707688321
transform 0 -1 1050 1 0 15809
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_60
timestamp 1707688321
transform 0 -1 1204 1 0 68
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_61
timestamp 1707688321
transform 0 -1 1204 1 0 1499
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_62
timestamp 1707688321
transform 0 -1 1204 1 0 2930
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_63
timestamp 1707688321
transform 0 -1 1204 1 0 4361
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_64
timestamp 1707688321
transform 0 -1 1204 1 0 5792
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_65
timestamp 1707688321
transform 0 -1 1204 1 0 7223
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_66
timestamp 1707688321
transform 0 -1 896 1 0 8654
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_67
timestamp 1707688321
transform 0 -1 896 1 0 7223
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_68
timestamp 1707688321
transform 0 -1 896 1 0 5792
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_69
timestamp 1707688321
transform 0 -1 896 1 0 4361
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_70
timestamp 1707688321
transform 0 -1 896 1 0 2930
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_71
timestamp 1707688321
transform 0 -1 896 1 0 1499
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_72
timestamp 1707688321
transform 0 -1 896 1 0 68
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_73
timestamp 1707688321
transform 0 -1 896 1 0 10085
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_74
timestamp 1707688321
transform 0 -1 896 1 0 11516
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_75
timestamp 1707688321
transform 0 -1 896 1 0 12947
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_76
timestamp 1707688321
transform 0 -1 896 1 0 14378
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_77
timestamp 1707688321
transform 0 -1 896 1 0 15809
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_78
timestamp 1707688321
transform 0 -1 742 1 0 11516
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_79
timestamp 1707688321
transform 0 -1 742 1 0 10085
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_80
timestamp 1707688321
transform 0 -1 742 1 0 68
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_81
timestamp 1707688321
transform 0 -1 742 1 0 1499
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_82
timestamp 1707688321
transform 0 -1 742 1 0 2930
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_83
timestamp 1707688321
transform 0 -1 742 1 0 4361
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_84
timestamp 1707688321
transform 0 -1 742 1 0 5792
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_85
timestamp 1707688321
transform 0 -1 742 1 0 7223
box -68 -26 1361 126
use nDFres_CDNS_524688791851142  nDFres_CDNS_524688791851142_86
timestamp 1707688321
transform 0 -1 742 1 0 8654
box -68 -26 1361 126
<< labels >>
flabel metal1 s 498 140 579 152 0 FreeSans 200 0 0 0 fb_out
port 1 nsew
<< properties >>
string GDS_END 79506792
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 79453912
string path -1.125 -0.050 -1.125 -1.125 31.875 -1.125 31.875 430.375 -1.125 430.375 -1.125 -0.050 
<< end >>
