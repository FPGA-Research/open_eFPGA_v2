magic
tech sky130B
timestamp 1707688321
<< poly >>
rect 0 5907 33 5915
rect 0 5890 8 5907
rect 25 5890 33 5907
rect 0 5873 33 5890
rect 0 5856 8 5873
rect 25 5856 33 5873
rect 0 5839 33 5856
rect 0 5822 8 5839
rect 25 5822 33 5839
rect 0 5805 33 5822
rect 0 5788 8 5805
rect 25 5788 33 5805
rect 0 5771 33 5788
rect 0 5754 8 5771
rect 25 5754 33 5771
rect 0 5737 33 5754
rect 0 5720 8 5737
rect 25 5720 33 5737
rect 0 5703 33 5720
rect 0 5686 8 5703
rect 25 5686 33 5703
rect 0 5669 33 5686
rect 0 5652 8 5669
rect 25 5652 33 5669
rect 0 5635 33 5652
rect 0 5618 8 5635
rect 25 5618 33 5635
rect 0 5601 33 5618
rect 0 5584 8 5601
rect 25 5584 33 5601
rect 0 5567 33 5584
rect 0 5550 8 5567
rect 25 5550 33 5567
rect 0 5533 33 5550
rect 0 5516 8 5533
rect 25 5516 33 5533
rect 0 5499 33 5516
rect 0 5482 8 5499
rect 25 5482 33 5499
rect 0 5465 33 5482
rect 0 5448 8 5465
rect 25 5448 33 5465
rect 0 5431 33 5448
rect 0 5414 8 5431
rect 25 5414 33 5431
rect 0 5397 33 5414
rect 0 5380 8 5397
rect 25 5380 33 5397
rect 0 5363 33 5380
rect 0 5346 8 5363
rect 25 5346 33 5363
rect 0 5329 33 5346
rect 0 5312 8 5329
rect 25 5312 33 5329
rect 0 5295 33 5312
rect 0 5278 8 5295
rect 25 5278 33 5295
rect 0 5261 33 5278
rect 0 5244 8 5261
rect 25 5244 33 5261
rect 0 5227 33 5244
rect 0 5210 8 5227
rect 25 5210 33 5227
rect 0 5193 33 5210
rect 0 5176 8 5193
rect 25 5176 33 5193
rect 0 5159 33 5176
rect 0 5142 8 5159
rect 25 5142 33 5159
rect 0 5125 33 5142
rect 0 5108 8 5125
rect 25 5108 33 5125
rect 0 5091 33 5108
rect 0 5074 8 5091
rect 25 5074 33 5091
rect 0 5057 33 5074
rect 0 5040 8 5057
rect 25 5040 33 5057
rect 0 5023 33 5040
rect 0 5006 8 5023
rect 25 5006 33 5023
rect 0 4989 33 5006
rect 0 4972 8 4989
rect 25 4972 33 4989
rect 0 4955 33 4972
rect 0 4938 8 4955
rect 25 4938 33 4955
rect 0 4921 33 4938
rect 0 4904 8 4921
rect 25 4904 33 4921
rect 0 4887 33 4904
rect 0 4870 8 4887
rect 25 4870 33 4887
rect 0 4853 33 4870
rect 0 4836 8 4853
rect 25 4836 33 4853
rect 0 4819 33 4836
rect 0 4802 8 4819
rect 25 4802 33 4819
rect 0 4785 33 4802
rect 0 4768 8 4785
rect 25 4768 33 4785
rect 0 4751 33 4768
rect 0 4734 8 4751
rect 25 4734 33 4751
rect 0 4717 33 4734
rect 0 4700 8 4717
rect 25 4700 33 4717
rect 0 4683 33 4700
rect 0 4666 8 4683
rect 25 4666 33 4683
rect 0 4649 33 4666
rect 0 4632 8 4649
rect 25 4632 33 4649
rect 0 4615 33 4632
rect 0 4598 8 4615
rect 25 4598 33 4615
rect 0 4581 33 4598
rect 0 4564 8 4581
rect 25 4564 33 4581
rect 0 4547 33 4564
rect 0 4530 8 4547
rect 25 4530 33 4547
rect 0 4513 33 4530
rect 0 4496 8 4513
rect 25 4496 33 4513
rect 0 4479 33 4496
rect 0 4462 8 4479
rect 25 4462 33 4479
rect 0 4445 33 4462
rect 0 4428 8 4445
rect 25 4428 33 4445
rect 0 4411 33 4428
rect 0 4394 8 4411
rect 25 4394 33 4411
rect 0 4377 33 4394
rect 0 4360 8 4377
rect 25 4360 33 4377
rect 0 4343 33 4360
rect 0 4326 8 4343
rect 25 4326 33 4343
rect 0 4309 33 4326
rect 0 4292 8 4309
rect 25 4292 33 4309
rect 0 4275 33 4292
rect 0 4258 8 4275
rect 25 4258 33 4275
rect 0 4241 33 4258
rect 0 4224 8 4241
rect 25 4224 33 4241
rect 0 4207 33 4224
rect 0 4190 8 4207
rect 25 4190 33 4207
rect 0 4173 33 4190
rect 0 4156 8 4173
rect 25 4156 33 4173
rect 0 4139 33 4156
rect 0 4122 8 4139
rect 25 4122 33 4139
rect 0 4105 33 4122
rect 0 4088 8 4105
rect 25 4088 33 4105
rect 0 4071 33 4088
rect 0 4054 8 4071
rect 25 4054 33 4071
rect 0 4037 33 4054
rect 0 4020 8 4037
rect 25 4020 33 4037
rect 0 4003 33 4020
rect 0 3986 8 4003
rect 25 3986 33 4003
rect 0 3969 33 3986
rect 0 3952 8 3969
rect 25 3952 33 3969
rect 0 3935 33 3952
rect 0 3918 8 3935
rect 25 3918 33 3935
rect 0 3901 33 3918
rect 0 3884 8 3901
rect 25 3884 33 3901
rect 0 3867 33 3884
rect 0 3850 8 3867
rect 25 3850 33 3867
rect 0 3833 33 3850
rect 0 3816 8 3833
rect 25 3816 33 3833
rect 0 3799 33 3816
rect 0 3782 8 3799
rect 25 3782 33 3799
rect 0 3765 33 3782
rect 0 3748 8 3765
rect 25 3748 33 3765
rect 0 3731 33 3748
rect 0 3714 8 3731
rect 25 3714 33 3731
rect 0 3697 33 3714
rect 0 3680 8 3697
rect 25 3680 33 3697
rect 0 3663 33 3680
rect 0 3646 8 3663
rect 25 3646 33 3663
rect 0 3629 33 3646
rect 0 3612 8 3629
rect 25 3612 33 3629
rect 0 3595 33 3612
rect 0 3578 8 3595
rect 25 3578 33 3595
rect 0 3561 33 3578
rect 0 3544 8 3561
rect 25 3544 33 3561
rect 0 3527 33 3544
rect 0 3510 8 3527
rect 25 3510 33 3527
rect 0 3493 33 3510
rect 0 3476 8 3493
rect 25 3476 33 3493
rect 0 3459 33 3476
rect 0 3442 8 3459
rect 25 3442 33 3459
rect 0 3425 33 3442
rect 0 3408 8 3425
rect 25 3408 33 3425
rect 0 3391 33 3408
rect 0 3374 8 3391
rect 25 3374 33 3391
rect 0 3357 33 3374
rect 0 3340 8 3357
rect 25 3340 33 3357
rect 0 3323 33 3340
rect 0 3306 8 3323
rect 25 3306 33 3323
rect 0 3289 33 3306
rect 0 3272 8 3289
rect 25 3272 33 3289
rect 0 3255 33 3272
rect 0 3238 8 3255
rect 25 3238 33 3255
rect 0 3221 33 3238
rect 0 3204 8 3221
rect 25 3204 33 3221
rect 0 3187 33 3204
rect 0 3170 8 3187
rect 25 3170 33 3187
rect 0 3153 33 3170
rect 0 3136 8 3153
rect 25 3136 33 3153
rect 0 3119 33 3136
rect 0 3102 8 3119
rect 25 3102 33 3119
rect 0 3085 33 3102
rect 0 3068 8 3085
rect 25 3068 33 3085
rect 0 3051 33 3068
rect 0 3034 8 3051
rect 25 3034 33 3051
rect 0 3017 33 3034
rect 0 3000 8 3017
rect 25 3000 33 3017
rect 0 2983 33 3000
rect 0 2966 8 2983
rect 25 2966 33 2983
rect 0 2949 33 2966
rect 0 2932 8 2949
rect 25 2932 33 2949
rect 0 2915 33 2932
rect 0 2898 8 2915
rect 25 2898 33 2915
rect 0 2881 33 2898
rect 0 2864 8 2881
rect 25 2864 33 2881
rect 0 2847 33 2864
rect 0 2830 8 2847
rect 25 2830 33 2847
rect 0 2813 33 2830
rect 0 2796 8 2813
rect 25 2796 33 2813
rect 0 2779 33 2796
rect 0 2762 8 2779
rect 25 2762 33 2779
rect 0 2745 33 2762
rect 0 2728 8 2745
rect 25 2728 33 2745
rect 0 2711 33 2728
rect 0 2694 8 2711
rect 25 2694 33 2711
rect 0 2677 33 2694
rect 0 2660 8 2677
rect 25 2660 33 2677
rect 0 2643 33 2660
rect 0 2626 8 2643
rect 25 2626 33 2643
rect 0 2609 33 2626
rect 0 2592 8 2609
rect 25 2592 33 2609
rect 0 2575 33 2592
rect 0 2558 8 2575
rect 25 2558 33 2575
rect 0 2541 33 2558
rect 0 2524 8 2541
rect 25 2524 33 2541
rect 0 2507 33 2524
rect 0 2490 8 2507
rect 25 2490 33 2507
rect 0 2473 33 2490
rect 0 2456 8 2473
rect 25 2456 33 2473
rect 0 2439 33 2456
rect 0 2422 8 2439
rect 25 2422 33 2439
rect 0 2405 33 2422
rect 0 2388 8 2405
rect 25 2388 33 2405
rect 0 2371 33 2388
rect 0 2354 8 2371
rect 25 2354 33 2371
rect 0 2337 33 2354
rect 0 2320 8 2337
rect 25 2320 33 2337
rect 0 2303 33 2320
rect 0 2286 8 2303
rect 25 2286 33 2303
rect 0 2269 33 2286
rect 0 2252 8 2269
rect 25 2252 33 2269
rect 0 2235 33 2252
rect 0 2218 8 2235
rect 25 2218 33 2235
rect 0 2201 33 2218
rect 0 2184 8 2201
rect 25 2184 33 2201
rect 0 2167 33 2184
rect 0 2150 8 2167
rect 25 2150 33 2167
rect 0 2133 33 2150
rect 0 2116 8 2133
rect 25 2116 33 2133
rect 0 2099 33 2116
rect 0 2082 8 2099
rect 25 2082 33 2099
rect 0 2065 33 2082
rect 0 2048 8 2065
rect 25 2048 33 2065
rect 0 2031 33 2048
rect 0 2014 8 2031
rect 25 2014 33 2031
rect 0 1997 33 2014
rect 0 1980 8 1997
rect 25 1980 33 1997
rect 0 1963 33 1980
rect 0 1946 8 1963
rect 25 1946 33 1963
rect 0 1929 33 1946
rect 0 1912 8 1929
rect 25 1912 33 1929
rect 0 1895 33 1912
rect 0 1878 8 1895
rect 25 1878 33 1895
rect 0 1861 33 1878
rect 0 1844 8 1861
rect 25 1844 33 1861
rect 0 1827 33 1844
rect 0 1810 8 1827
rect 25 1810 33 1827
rect 0 1793 33 1810
rect 0 1776 8 1793
rect 25 1776 33 1793
rect 0 1759 33 1776
rect 0 1742 8 1759
rect 25 1742 33 1759
rect 0 1725 33 1742
rect 0 1708 8 1725
rect 25 1708 33 1725
rect 0 1691 33 1708
rect 0 1674 8 1691
rect 25 1674 33 1691
rect 0 1657 33 1674
rect 0 1640 8 1657
rect 25 1640 33 1657
rect 0 1623 33 1640
rect 0 1606 8 1623
rect 25 1606 33 1623
rect 0 1589 33 1606
rect 0 1572 8 1589
rect 25 1572 33 1589
rect 0 1555 33 1572
rect 0 1538 8 1555
rect 25 1538 33 1555
rect 0 1521 33 1538
rect 0 1504 8 1521
rect 25 1504 33 1521
rect 0 1487 33 1504
rect 0 1470 8 1487
rect 25 1470 33 1487
rect 0 1453 33 1470
rect 0 1436 8 1453
rect 25 1436 33 1453
rect 0 1419 33 1436
rect 0 1402 8 1419
rect 25 1402 33 1419
rect 0 1385 33 1402
rect 0 1368 8 1385
rect 25 1368 33 1385
rect 0 1351 33 1368
rect 0 1334 8 1351
rect 25 1334 33 1351
rect 0 1317 33 1334
rect 0 1300 8 1317
rect 25 1300 33 1317
rect 0 1283 33 1300
rect 0 1266 8 1283
rect 25 1266 33 1283
rect 0 1249 33 1266
rect 0 1232 8 1249
rect 25 1232 33 1249
rect 0 1215 33 1232
rect 0 1198 8 1215
rect 25 1198 33 1215
rect 0 1181 33 1198
rect 0 1164 8 1181
rect 25 1164 33 1181
rect 0 1147 33 1164
rect 0 1130 8 1147
rect 25 1130 33 1147
rect 0 1113 33 1130
rect 0 1096 8 1113
rect 25 1096 33 1113
rect 0 1079 33 1096
rect 0 1062 8 1079
rect 25 1062 33 1079
rect 0 1045 33 1062
rect 0 1028 8 1045
rect 25 1028 33 1045
rect 0 1011 33 1028
rect 0 994 8 1011
rect 25 994 33 1011
rect 0 977 33 994
rect 0 960 8 977
rect 25 960 33 977
rect 0 943 33 960
rect 0 926 8 943
rect 25 926 33 943
rect 0 909 33 926
rect 0 892 8 909
rect 25 892 33 909
rect 0 875 33 892
rect 0 858 8 875
rect 25 858 33 875
rect 0 841 33 858
rect 0 824 8 841
rect 25 824 33 841
rect 0 807 33 824
rect 0 790 8 807
rect 25 790 33 807
rect 0 773 33 790
rect 0 756 8 773
rect 25 756 33 773
rect 0 739 33 756
rect 0 722 8 739
rect 25 722 33 739
rect 0 705 33 722
rect 0 688 8 705
rect 25 688 33 705
rect 0 671 33 688
rect 0 654 8 671
rect 25 654 33 671
rect 0 637 33 654
rect 0 620 8 637
rect 25 620 33 637
rect 0 603 33 620
rect 0 586 8 603
rect 25 586 33 603
rect 0 569 33 586
rect 0 552 8 569
rect 25 552 33 569
rect 0 535 33 552
rect 0 518 8 535
rect 25 518 33 535
rect 0 501 33 518
rect 0 484 8 501
rect 25 484 33 501
rect 0 467 33 484
rect 0 450 8 467
rect 25 450 33 467
rect 0 433 33 450
rect 0 416 8 433
rect 25 416 33 433
rect 0 399 33 416
rect 0 382 8 399
rect 25 382 33 399
rect 0 365 33 382
rect 0 348 8 365
rect 25 348 33 365
rect 0 331 33 348
rect 0 314 8 331
rect 25 314 33 331
rect 0 297 33 314
rect 0 280 8 297
rect 25 280 33 297
rect 0 263 33 280
rect 0 246 8 263
rect 25 246 33 263
rect 0 229 33 246
rect 0 212 8 229
rect 25 212 33 229
rect 0 195 33 212
rect 0 178 8 195
rect 25 178 33 195
rect 0 161 33 178
rect 0 144 8 161
rect 25 144 33 161
rect 0 127 33 144
rect 0 110 8 127
rect 25 110 33 127
rect 0 93 33 110
rect 0 76 8 93
rect 25 76 33 93
rect 0 59 33 76
rect 0 42 8 59
rect 25 42 33 59
rect 0 25 33 42
rect 0 8 8 25
rect 25 8 33 25
rect 0 0 33 8
<< polycont >>
rect 8 5890 25 5907
rect 8 5856 25 5873
rect 8 5822 25 5839
rect 8 5788 25 5805
rect 8 5754 25 5771
rect 8 5720 25 5737
rect 8 5686 25 5703
rect 8 5652 25 5669
rect 8 5618 25 5635
rect 8 5584 25 5601
rect 8 5550 25 5567
rect 8 5516 25 5533
rect 8 5482 25 5499
rect 8 5448 25 5465
rect 8 5414 25 5431
rect 8 5380 25 5397
rect 8 5346 25 5363
rect 8 5312 25 5329
rect 8 5278 25 5295
rect 8 5244 25 5261
rect 8 5210 25 5227
rect 8 5176 25 5193
rect 8 5142 25 5159
rect 8 5108 25 5125
rect 8 5074 25 5091
rect 8 5040 25 5057
rect 8 5006 25 5023
rect 8 4972 25 4989
rect 8 4938 25 4955
rect 8 4904 25 4921
rect 8 4870 25 4887
rect 8 4836 25 4853
rect 8 4802 25 4819
rect 8 4768 25 4785
rect 8 4734 25 4751
rect 8 4700 25 4717
rect 8 4666 25 4683
rect 8 4632 25 4649
rect 8 4598 25 4615
rect 8 4564 25 4581
rect 8 4530 25 4547
rect 8 4496 25 4513
rect 8 4462 25 4479
rect 8 4428 25 4445
rect 8 4394 25 4411
rect 8 4360 25 4377
rect 8 4326 25 4343
rect 8 4292 25 4309
rect 8 4258 25 4275
rect 8 4224 25 4241
rect 8 4190 25 4207
rect 8 4156 25 4173
rect 8 4122 25 4139
rect 8 4088 25 4105
rect 8 4054 25 4071
rect 8 4020 25 4037
rect 8 3986 25 4003
rect 8 3952 25 3969
rect 8 3918 25 3935
rect 8 3884 25 3901
rect 8 3850 25 3867
rect 8 3816 25 3833
rect 8 3782 25 3799
rect 8 3748 25 3765
rect 8 3714 25 3731
rect 8 3680 25 3697
rect 8 3646 25 3663
rect 8 3612 25 3629
rect 8 3578 25 3595
rect 8 3544 25 3561
rect 8 3510 25 3527
rect 8 3476 25 3493
rect 8 3442 25 3459
rect 8 3408 25 3425
rect 8 3374 25 3391
rect 8 3340 25 3357
rect 8 3306 25 3323
rect 8 3272 25 3289
rect 8 3238 25 3255
rect 8 3204 25 3221
rect 8 3170 25 3187
rect 8 3136 25 3153
rect 8 3102 25 3119
rect 8 3068 25 3085
rect 8 3034 25 3051
rect 8 3000 25 3017
rect 8 2966 25 2983
rect 8 2932 25 2949
rect 8 2898 25 2915
rect 8 2864 25 2881
rect 8 2830 25 2847
rect 8 2796 25 2813
rect 8 2762 25 2779
rect 8 2728 25 2745
rect 8 2694 25 2711
rect 8 2660 25 2677
rect 8 2626 25 2643
rect 8 2592 25 2609
rect 8 2558 25 2575
rect 8 2524 25 2541
rect 8 2490 25 2507
rect 8 2456 25 2473
rect 8 2422 25 2439
rect 8 2388 25 2405
rect 8 2354 25 2371
rect 8 2320 25 2337
rect 8 2286 25 2303
rect 8 2252 25 2269
rect 8 2218 25 2235
rect 8 2184 25 2201
rect 8 2150 25 2167
rect 8 2116 25 2133
rect 8 2082 25 2099
rect 8 2048 25 2065
rect 8 2014 25 2031
rect 8 1980 25 1997
rect 8 1946 25 1963
rect 8 1912 25 1929
rect 8 1878 25 1895
rect 8 1844 25 1861
rect 8 1810 25 1827
rect 8 1776 25 1793
rect 8 1742 25 1759
rect 8 1708 25 1725
rect 8 1674 25 1691
rect 8 1640 25 1657
rect 8 1606 25 1623
rect 8 1572 25 1589
rect 8 1538 25 1555
rect 8 1504 25 1521
rect 8 1470 25 1487
rect 8 1436 25 1453
rect 8 1402 25 1419
rect 8 1368 25 1385
rect 8 1334 25 1351
rect 8 1300 25 1317
rect 8 1266 25 1283
rect 8 1232 25 1249
rect 8 1198 25 1215
rect 8 1164 25 1181
rect 8 1130 25 1147
rect 8 1096 25 1113
rect 8 1062 25 1079
rect 8 1028 25 1045
rect 8 994 25 1011
rect 8 960 25 977
rect 8 926 25 943
rect 8 892 25 909
rect 8 858 25 875
rect 8 824 25 841
rect 8 790 25 807
rect 8 756 25 773
rect 8 722 25 739
rect 8 688 25 705
rect 8 654 25 671
rect 8 620 25 637
rect 8 586 25 603
rect 8 552 25 569
rect 8 518 25 535
rect 8 484 25 501
rect 8 450 25 467
rect 8 416 25 433
rect 8 382 25 399
rect 8 348 25 365
rect 8 314 25 331
rect 8 280 25 297
rect 8 246 25 263
rect 8 212 25 229
rect 8 178 25 195
rect 8 144 25 161
rect 8 110 25 127
rect 8 76 25 93
rect 8 42 25 59
rect 8 8 25 25
<< locali >>
rect 8 5907 25 5915
rect 8 5873 25 5890
rect 8 5839 25 5856
rect 8 5805 25 5822
rect 8 5771 25 5788
rect 8 5737 25 5754
rect 8 5703 25 5720
rect 8 5669 25 5686
rect 8 5635 25 5652
rect 8 5601 25 5618
rect 8 5567 25 5584
rect 8 5533 25 5550
rect 8 5499 25 5516
rect 8 5465 25 5482
rect 8 5431 25 5448
rect 8 5397 25 5414
rect 8 5363 25 5380
rect 8 5329 25 5346
rect 8 5295 25 5312
rect 8 5261 25 5278
rect 8 5227 25 5244
rect 8 5193 25 5210
rect 8 5159 25 5176
rect 8 5125 25 5142
rect 8 5091 25 5108
rect 8 5057 25 5074
rect 8 5023 25 5040
rect 8 4989 25 5006
rect 8 4955 25 4972
rect 8 4921 25 4938
rect 8 4887 25 4904
rect 8 4853 25 4870
rect 8 4819 25 4836
rect 8 4785 25 4802
rect 8 4751 25 4768
rect 8 4717 25 4734
rect 8 4683 25 4700
rect 8 4649 25 4666
rect 8 4615 25 4632
rect 8 4581 25 4598
rect 8 4547 25 4564
rect 8 4513 25 4530
rect 8 4479 25 4496
rect 8 4445 25 4462
rect 8 4411 25 4428
rect 8 4377 25 4394
rect 8 4343 25 4360
rect 8 4309 25 4326
rect 8 4275 25 4292
rect 8 4241 25 4258
rect 8 4207 25 4224
rect 8 4173 25 4190
rect 8 4139 25 4156
rect 8 4105 25 4122
rect 8 4071 25 4088
rect 8 4037 25 4054
rect 8 4003 25 4020
rect 8 3969 25 3986
rect 8 3935 25 3952
rect 8 3901 25 3918
rect 8 3867 25 3884
rect 8 3833 25 3850
rect 8 3799 25 3816
rect 8 3765 25 3782
rect 8 3731 25 3748
rect 8 3697 25 3714
rect 8 3663 25 3680
rect 8 3629 25 3646
rect 8 3595 25 3612
rect 8 3561 25 3578
rect 8 3527 25 3544
rect 8 3493 25 3510
rect 8 3459 25 3476
rect 8 3425 25 3442
rect 8 3391 25 3408
rect 8 3357 25 3374
rect 8 3323 25 3340
rect 8 3289 25 3306
rect 8 3255 25 3272
rect 8 3221 25 3238
rect 8 3187 25 3204
rect 8 3153 25 3170
rect 8 3119 25 3136
rect 8 3085 25 3102
rect 8 3051 25 3068
rect 8 3017 25 3034
rect 8 2983 25 3000
rect 8 2949 25 2966
rect 8 2915 25 2932
rect 8 2881 25 2898
rect 8 2847 25 2864
rect 8 2813 25 2830
rect 8 2779 25 2796
rect 8 2745 25 2762
rect 8 2711 25 2728
rect 8 2677 25 2694
rect 8 2643 25 2660
rect 8 2609 25 2626
rect 8 2575 25 2592
rect 8 2541 25 2558
rect 8 2507 25 2524
rect 8 2473 25 2490
rect 8 2439 25 2456
rect 8 2405 25 2422
rect 8 2371 25 2388
rect 8 2337 25 2354
rect 8 2303 25 2320
rect 8 2269 25 2286
rect 8 2235 25 2252
rect 8 2201 25 2218
rect 8 2167 25 2184
rect 8 2133 25 2150
rect 8 2099 25 2116
rect 8 2065 25 2082
rect 8 2031 25 2048
rect 8 1997 25 2014
rect 8 1963 25 1980
rect 8 1929 25 1946
rect 8 1895 25 1912
rect 8 1861 25 1878
rect 8 1827 25 1844
rect 8 1793 25 1810
rect 8 1759 25 1776
rect 8 1725 25 1742
rect 8 1691 25 1708
rect 8 1657 25 1674
rect 8 1623 25 1640
rect 8 1589 25 1606
rect 8 1555 25 1572
rect 8 1521 25 1538
rect 8 1487 25 1504
rect 8 1453 25 1470
rect 8 1419 25 1436
rect 8 1385 25 1402
rect 8 1351 25 1368
rect 8 1317 25 1334
rect 8 1283 25 1300
rect 8 1249 25 1266
rect 8 1215 25 1232
rect 8 1181 25 1198
rect 8 1147 25 1164
rect 8 1113 25 1130
rect 8 1079 25 1096
rect 8 1045 25 1062
rect 8 1011 25 1028
rect 8 977 25 994
rect 8 943 25 960
rect 8 909 25 926
rect 8 875 25 892
rect 8 841 25 858
rect 8 807 25 824
rect 8 773 25 790
rect 8 739 25 756
rect 8 705 25 722
rect 8 671 25 688
rect 8 637 25 654
rect 8 603 25 620
rect 8 569 25 586
rect 8 535 25 552
rect 8 501 25 518
rect 8 467 25 484
rect 8 433 25 450
rect 8 399 25 416
rect 8 365 25 382
rect 8 331 25 348
rect 8 297 25 314
rect 8 263 25 280
rect 8 229 25 246
rect 8 195 25 212
rect 8 161 25 178
rect 8 127 25 144
rect 8 93 25 110
rect 8 59 25 76
rect 8 25 25 42
rect 8 0 25 8
<< properties >>
string GDS_END 80380088
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 80368756
<< end >>
