magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -89 -36 217 636
<< pmos >>
rect 0 0 36 600
rect 92 0 128 600
<< pdiff >>
rect -50 0 0 600
rect 128 0 178 600
<< poly >>
rect 0 600 36 626
rect 0 -26 36 0
rect 92 600 128 626
rect 92 -26 128 0
<< locali >>
rect -45 -4 -11 538
rect 47 -4 81 538
rect 139 -4 173 538
use hvDFL1sd2_CDNS_52468879185138  hvDFL1sd2_CDNS_52468879185138_0
timestamp 1707688321
transform 1 0 36 0 1 0
box -36 -36 92 636
use hvDFL1sd_CDNS_52468879185135  hvDFL1sd_CDNS_52468879185135_0
timestamp 1707688321
transform -1 0 0 0 1 0
box -36 -36 89 636
use hvDFL1sd_CDNS_52468879185135  hvDFL1sd_CDNS_52468879185135_1
timestamp 1707688321
transform 1 0 128 0 1 0
box -36 -36 89 636
<< labels >>
flabel comment s -28 267 -28 267 0 FreeSans 300 0 0 0 S
flabel comment s 64 267 64 267 0 FreeSans 300 0 0 0 D
flabel comment s 156 267 156 267 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 79586246
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 79584856
<< end >>
