magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< poly >>
rect -50 50 0 66
rect -50 16 -34 50
rect -50 0 0 16
rect 1137 50 1187 66
rect 1171 16 1187 50
rect 1137 0 1187 16
<< polycont >>
rect -34 16 0 50
rect 1137 16 1171 50
<< npolyres >>
rect 0 0 1137 66
<< locali >>
rect -34 50 0 66
rect -34 0 0 16
rect 1137 50 1171 66
rect 1137 0 1171 16
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_0
timestamp 1707688321
transform -1 0 16 0 1 0
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_1
timestamp 1707688321
transform 1 0 1121 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 86903924
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86903490
<< end >>
