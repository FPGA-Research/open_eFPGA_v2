magic
tech sky130B
timestamp 1707688321
<< properties >>
string GDS_END 86902300
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86901976
<< end >>
