magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< pwell >>
rect 10 66 1950 1536
<< mvnmos >>
rect 228 92 328 1510
rect 384 92 484 1510
rect 540 92 640 1510
rect 696 92 796 1510
rect 852 92 952 1510
rect 1008 92 1108 1510
rect 1164 92 1264 1510
rect 1320 92 1420 1510
rect 1476 92 1576 1510
rect 1632 92 1732 1510
<< mvndiff >>
rect 172 1498 228 1510
rect 172 1464 183 1498
rect 217 1464 228 1498
rect 172 1430 228 1464
rect 172 1396 183 1430
rect 217 1396 228 1430
rect 172 1362 228 1396
rect 172 1328 183 1362
rect 217 1328 228 1362
rect 172 1294 228 1328
rect 172 1260 183 1294
rect 217 1260 228 1294
rect 172 1226 228 1260
rect 172 1192 183 1226
rect 217 1192 228 1226
rect 172 1158 228 1192
rect 172 1124 183 1158
rect 217 1124 228 1158
rect 172 1090 228 1124
rect 172 1056 183 1090
rect 217 1056 228 1090
rect 172 1022 228 1056
rect 172 988 183 1022
rect 217 988 228 1022
rect 172 954 228 988
rect 172 920 183 954
rect 217 920 228 954
rect 172 886 228 920
rect 172 852 183 886
rect 217 852 228 886
rect 172 818 228 852
rect 172 784 183 818
rect 217 784 228 818
rect 172 750 228 784
rect 172 716 183 750
rect 217 716 228 750
rect 172 682 228 716
rect 172 648 183 682
rect 217 648 228 682
rect 172 614 228 648
rect 172 580 183 614
rect 217 580 228 614
rect 172 546 228 580
rect 172 512 183 546
rect 217 512 228 546
rect 172 478 228 512
rect 172 444 183 478
rect 217 444 228 478
rect 172 410 228 444
rect 172 376 183 410
rect 217 376 228 410
rect 172 342 228 376
rect 172 308 183 342
rect 217 308 228 342
rect 172 274 228 308
rect 172 240 183 274
rect 217 240 228 274
rect 172 206 228 240
rect 172 172 183 206
rect 217 172 228 206
rect 172 138 228 172
rect 172 104 183 138
rect 217 104 228 138
rect 172 92 228 104
rect 328 1498 384 1510
rect 328 1464 339 1498
rect 373 1464 384 1498
rect 328 1430 384 1464
rect 328 1396 339 1430
rect 373 1396 384 1430
rect 328 1362 384 1396
rect 328 1328 339 1362
rect 373 1328 384 1362
rect 328 1294 384 1328
rect 328 1260 339 1294
rect 373 1260 384 1294
rect 328 1226 384 1260
rect 328 1192 339 1226
rect 373 1192 384 1226
rect 328 1158 384 1192
rect 328 1124 339 1158
rect 373 1124 384 1158
rect 328 1090 384 1124
rect 328 1056 339 1090
rect 373 1056 384 1090
rect 328 1022 384 1056
rect 328 988 339 1022
rect 373 988 384 1022
rect 328 954 384 988
rect 328 920 339 954
rect 373 920 384 954
rect 328 886 384 920
rect 328 852 339 886
rect 373 852 384 886
rect 328 818 384 852
rect 328 784 339 818
rect 373 784 384 818
rect 328 750 384 784
rect 328 716 339 750
rect 373 716 384 750
rect 328 682 384 716
rect 328 648 339 682
rect 373 648 384 682
rect 328 614 384 648
rect 328 580 339 614
rect 373 580 384 614
rect 328 546 384 580
rect 328 512 339 546
rect 373 512 384 546
rect 328 478 384 512
rect 328 444 339 478
rect 373 444 384 478
rect 328 410 384 444
rect 328 376 339 410
rect 373 376 384 410
rect 328 342 384 376
rect 328 308 339 342
rect 373 308 384 342
rect 328 274 384 308
rect 328 240 339 274
rect 373 240 384 274
rect 328 206 384 240
rect 328 172 339 206
rect 373 172 384 206
rect 328 138 384 172
rect 328 104 339 138
rect 373 104 384 138
rect 328 92 384 104
rect 484 1498 540 1510
rect 484 1464 495 1498
rect 529 1464 540 1498
rect 484 1430 540 1464
rect 484 1396 495 1430
rect 529 1396 540 1430
rect 484 1362 540 1396
rect 484 1328 495 1362
rect 529 1328 540 1362
rect 484 1294 540 1328
rect 484 1260 495 1294
rect 529 1260 540 1294
rect 484 1226 540 1260
rect 484 1192 495 1226
rect 529 1192 540 1226
rect 484 1158 540 1192
rect 484 1124 495 1158
rect 529 1124 540 1158
rect 484 1090 540 1124
rect 484 1056 495 1090
rect 529 1056 540 1090
rect 484 1022 540 1056
rect 484 988 495 1022
rect 529 988 540 1022
rect 484 954 540 988
rect 484 920 495 954
rect 529 920 540 954
rect 484 886 540 920
rect 484 852 495 886
rect 529 852 540 886
rect 484 818 540 852
rect 484 784 495 818
rect 529 784 540 818
rect 484 750 540 784
rect 484 716 495 750
rect 529 716 540 750
rect 484 682 540 716
rect 484 648 495 682
rect 529 648 540 682
rect 484 614 540 648
rect 484 580 495 614
rect 529 580 540 614
rect 484 546 540 580
rect 484 512 495 546
rect 529 512 540 546
rect 484 478 540 512
rect 484 444 495 478
rect 529 444 540 478
rect 484 410 540 444
rect 484 376 495 410
rect 529 376 540 410
rect 484 342 540 376
rect 484 308 495 342
rect 529 308 540 342
rect 484 274 540 308
rect 484 240 495 274
rect 529 240 540 274
rect 484 206 540 240
rect 484 172 495 206
rect 529 172 540 206
rect 484 138 540 172
rect 484 104 495 138
rect 529 104 540 138
rect 484 92 540 104
rect 640 1498 696 1510
rect 640 1464 651 1498
rect 685 1464 696 1498
rect 640 1430 696 1464
rect 640 1396 651 1430
rect 685 1396 696 1430
rect 640 1362 696 1396
rect 640 1328 651 1362
rect 685 1328 696 1362
rect 640 1294 696 1328
rect 640 1260 651 1294
rect 685 1260 696 1294
rect 640 1226 696 1260
rect 640 1192 651 1226
rect 685 1192 696 1226
rect 640 1158 696 1192
rect 640 1124 651 1158
rect 685 1124 696 1158
rect 640 1090 696 1124
rect 640 1056 651 1090
rect 685 1056 696 1090
rect 640 1022 696 1056
rect 640 988 651 1022
rect 685 988 696 1022
rect 640 954 696 988
rect 640 920 651 954
rect 685 920 696 954
rect 640 886 696 920
rect 640 852 651 886
rect 685 852 696 886
rect 640 818 696 852
rect 640 784 651 818
rect 685 784 696 818
rect 640 750 696 784
rect 640 716 651 750
rect 685 716 696 750
rect 640 682 696 716
rect 640 648 651 682
rect 685 648 696 682
rect 640 614 696 648
rect 640 580 651 614
rect 685 580 696 614
rect 640 546 696 580
rect 640 512 651 546
rect 685 512 696 546
rect 640 478 696 512
rect 640 444 651 478
rect 685 444 696 478
rect 640 410 696 444
rect 640 376 651 410
rect 685 376 696 410
rect 640 342 696 376
rect 640 308 651 342
rect 685 308 696 342
rect 640 274 696 308
rect 640 240 651 274
rect 685 240 696 274
rect 640 206 696 240
rect 640 172 651 206
rect 685 172 696 206
rect 640 138 696 172
rect 640 104 651 138
rect 685 104 696 138
rect 640 92 696 104
rect 796 1498 852 1510
rect 796 1464 807 1498
rect 841 1464 852 1498
rect 796 1430 852 1464
rect 796 1396 807 1430
rect 841 1396 852 1430
rect 796 1362 852 1396
rect 796 1328 807 1362
rect 841 1328 852 1362
rect 796 1294 852 1328
rect 796 1260 807 1294
rect 841 1260 852 1294
rect 796 1226 852 1260
rect 796 1192 807 1226
rect 841 1192 852 1226
rect 796 1158 852 1192
rect 796 1124 807 1158
rect 841 1124 852 1158
rect 796 1090 852 1124
rect 796 1056 807 1090
rect 841 1056 852 1090
rect 796 1022 852 1056
rect 796 988 807 1022
rect 841 988 852 1022
rect 796 954 852 988
rect 796 920 807 954
rect 841 920 852 954
rect 796 886 852 920
rect 796 852 807 886
rect 841 852 852 886
rect 796 818 852 852
rect 796 784 807 818
rect 841 784 852 818
rect 796 750 852 784
rect 796 716 807 750
rect 841 716 852 750
rect 796 682 852 716
rect 796 648 807 682
rect 841 648 852 682
rect 796 614 852 648
rect 796 580 807 614
rect 841 580 852 614
rect 796 546 852 580
rect 796 512 807 546
rect 841 512 852 546
rect 796 478 852 512
rect 796 444 807 478
rect 841 444 852 478
rect 796 410 852 444
rect 796 376 807 410
rect 841 376 852 410
rect 796 342 852 376
rect 796 308 807 342
rect 841 308 852 342
rect 796 274 852 308
rect 796 240 807 274
rect 841 240 852 274
rect 796 206 852 240
rect 796 172 807 206
rect 841 172 852 206
rect 796 138 852 172
rect 796 104 807 138
rect 841 104 852 138
rect 796 92 852 104
rect 952 1498 1008 1510
rect 952 1464 963 1498
rect 997 1464 1008 1498
rect 952 1430 1008 1464
rect 952 1396 963 1430
rect 997 1396 1008 1430
rect 952 1362 1008 1396
rect 952 1328 963 1362
rect 997 1328 1008 1362
rect 952 1294 1008 1328
rect 952 1260 963 1294
rect 997 1260 1008 1294
rect 952 1226 1008 1260
rect 952 1192 963 1226
rect 997 1192 1008 1226
rect 952 1158 1008 1192
rect 952 1124 963 1158
rect 997 1124 1008 1158
rect 952 1090 1008 1124
rect 952 1056 963 1090
rect 997 1056 1008 1090
rect 952 1022 1008 1056
rect 952 988 963 1022
rect 997 988 1008 1022
rect 952 954 1008 988
rect 952 920 963 954
rect 997 920 1008 954
rect 952 886 1008 920
rect 952 852 963 886
rect 997 852 1008 886
rect 952 818 1008 852
rect 952 784 963 818
rect 997 784 1008 818
rect 952 750 1008 784
rect 952 716 963 750
rect 997 716 1008 750
rect 952 682 1008 716
rect 952 648 963 682
rect 997 648 1008 682
rect 952 614 1008 648
rect 952 580 963 614
rect 997 580 1008 614
rect 952 546 1008 580
rect 952 512 963 546
rect 997 512 1008 546
rect 952 478 1008 512
rect 952 444 963 478
rect 997 444 1008 478
rect 952 410 1008 444
rect 952 376 963 410
rect 997 376 1008 410
rect 952 342 1008 376
rect 952 308 963 342
rect 997 308 1008 342
rect 952 274 1008 308
rect 952 240 963 274
rect 997 240 1008 274
rect 952 206 1008 240
rect 952 172 963 206
rect 997 172 1008 206
rect 952 138 1008 172
rect 952 104 963 138
rect 997 104 1008 138
rect 952 92 1008 104
rect 1108 1498 1164 1510
rect 1108 1464 1119 1498
rect 1153 1464 1164 1498
rect 1108 1430 1164 1464
rect 1108 1396 1119 1430
rect 1153 1396 1164 1430
rect 1108 1362 1164 1396
rect 1108 1328 1119 1362
rect 1153 1328 1164 1362
rect 1108 1294 1164 1328
rect 1108 1260 1119 1294
rect 1153 1260 1164 1294
rect 1108 1226 1164 1260
rect 1108 1192 1119 1226
rect 1153 1192 1164 1226
rect 1108 1158 1164 1192
rect 1108 1124 1119 1158
rect 1153 1124 1164 1158
rect 1108 1090 1164 1124
rect 1108 1056 1119 1090
rect 1153 1056 1164 1090
rect 1108 1022 1164 1056
rect 1108 988 1119 1022
rect 1153 988 1164 1022
rect 1108 954 1164 988
rect 1108 920 1119 954
rect 1153 920 1164 954
rect 1108 886 1164 920
rect 1108 852 1119 886
rect 1153 852 1164 886
rect 1108 818 1164 852
rect 1108 784 1119 818
rect 1153 784 1164 818
rect 1108 750 1164 784
rect 1108 716 1119 750
rect 1153 716 1164 750
rect 1108 682 1164 716
rect 1108 648 1119 682
rect 1153 648 1164 682
rect 1108 614 1164 648
rect 1108 580 1119 614
rect 1153 580 1164 614
rect 1108 546 1164 580
rect 1108 512 1119 546
rect 1153 512 1164 546
rect 1108 478 1164 512
rect 1108 444 1119 478
rect 1153 444 1164 478
rect 1108 410 1164 444
rect 1108 376 1119 410
rect 1153 376 1164 410
rect 1108 342 1164 376
rect 1108 308 1119 342
rect 1153 308 1164 342
rect 1108 274 1164 308
rect 1108 240 1119 274
rect 1153 240 1164 274
rect 1108 206 1164 240
rect 1108 172 1119 206
rect 1153 172 1164 206
rect 1108 138 1164 172
rect 1108 104 1119 138
rect 1153 104 1164 138
rect 1108 92 1164 104
rect 1264 1498 1320 1510
rect 1264 1464 1275 1498
rect 1309 1464 1320 1498
rect 1264 1430 1320 1464
rect 1264 1396 1275 1430
rect 1309 1396 1320 1430
rect 1264 1362 1320 1396
rect 1264 1328 1275 1362
rect 1309 1328 1320 1362
rect 1264 1294 1320 1328
rect 1264 1260 1275 1294
rect 1309 1260 1320 1294
rect 1264 1226 1320 1260
rect 1264 1192 1275 1226
rect 1309 1192 1320 1226
rect 1264 1158 1320 1192
rect 1264 1124 1275 1158
rect 1309 1124 1320 1158
rect 1264 1090 1320 1124
rect 1264 1056 1275 1090
rect 1309 1056 1320 1090
rect 1264 1022 1320 1056
rect 1264 988 1275 1022
rect 1309 988 1320 1022
rect 1264 954 1320 988
rect 1264 920 1275 954
rect 1309 920 1320 954
rect 1264 886 1320 920
rect 1264 852 1275 886
rect 1309 852 1320 886
rect 1264 818 1320 852
rect 1264 784 1275 818
rect 1309 784 1320 818
rect 1264 750 1320 784
rect 1264 716 1275 750
rect 1309 716 1320 750
rect 1264 682 1320 716
rect 1264 648 1275 682
rect 1309 648 1320 682
rect 1264 614 1320 648
rect 1264 580 1275 614
rect 1309 580 1320 614
rect 1264 546 1320 580
rect 1264 512 1275 546
rect 1309 512 1320 546
rect 1264 478 1320 512
rect 1264 444 1275 478
rect 1309 444 1320 478
rect 1264 410 1320 444
rect 1264 376 1275 410
rect 1309 376 1320 410
rect 1264 342 1320 376
rect 1264 308 1275 342
rect 1309 308 1320 342
rect 1264 274 1320 308
rect 1264 240 1275 274
rect 1309 240 1320 274
rect 1264 206 1320 240
rect 1264 172 1275 206
rect 1309 172 1320 206
rect 1264 138 1320 172
rect 1264 104 1275 138
rect 1309 104 1320 138
rect 1264 92 1320 104
rect 1420 1498 1476 1510
rect 1420 1464 1431 1498
rect 1465 1464 1476 1498
rect 1420 1430 1476 1464
rect 1420 1396 1431 1430
rect 1465 1396 1476 1430
rect 1420 1362 1476 1396
rect 1420 1328 1431 1362
rect 1465 1328 1476 1362
rect 1420 1294 1476 1328
rect 1420 1260 1431 1294
rect 1465 1260 1476 1294
rect 1420 1226 1476 1260
rect 1420 1192 1431 1226
rect 1465 1192 1476 1226
rect 1420 1158 1476 1192
rect 1420 1124 1431 1158
rect 1465 1124 1476 1158
rect 1420 1090 1476 1124
rect 1420 1056 1431 1090
rect 1465 1056 1476 1090
rect 1420 1022 1476 1056
rect 1420 988 1431 1022
rect 1465 988 1476 1022
rect 1420 954 1476 988
rect 1420 920 1431 954
rect 1465 920 1476 954
rect 1420 886 1476 920
rect 1420 852 1431 886
rect 1465 852 1476 886
rect 1420 818 1476 852
rect 1420 784 1431 818
rect 1465 784 1476 818
rect 1420 750 1476 784
rect 1420 716 1431 750
rect 1465 716 1476 750
rect 1420 682 1476 716
rect 1420 648 1431 682
rect 1465 648 1476 682
rect 1420 614 1476 648
rect 1420 580 1431 614
rect 1465 580 1476 614
rect 1420 546 1476 580
rect 1420 512 1431 546
rect 1465 512 1476 546
rect 1420 478 1476 512
rect 1420 444 1431 478
rect 1465 444 1476 478
rect 1420 410 1476 444
rect 1420 376 1431 410
rect 1465 376 1476 410
rect 1420 342 1476 376
rect 1420 308 1431 342
rect 1465 308 1476 342
rect 1420 274 1476 308
rect 1420 240 1431 274
rect 1465 240 1476 274
rect 1420 206 1476 240
rect 1420 172 1431 206
rect 1465 172 1476 206
rect 1420 138 1476 172
rect 1420 104 1431 138
rect 1465 104 1476 138
rect 1420 92 1476 104
rect 1576 1498 1632 1510
rect 1576 1464 1587 1498
rect 1621 1464 1632 1498
rect 1576 1430 1632 1464
rect 1576 1396 1587 1430
rect 1621 1396 1632 1430
rect 1576 1362 1632 1396
rect 1576 1328 1587 1362
rect 1621 1328 1632 1362
rect 1576 1294 1632 1328
rect 1576 1260 1587 1294
rect 1621 1260 1632 1294
rect 1576 1226 1632 1260
rect 1576 1192 1587 1226
rect 1621 1192 1632 1226
rect 1576 1158 1632 1192
rect 1576 1124 1587 1158
rect 1621 1124 1632 1158
rect 1576 1090 1632 1124
rect 1576 1056 1587 1090
rect 1621 1056 1632 1090
rect 1576 1022 1632 1056
rect 1576 988 1587 1022
rect 1621 988 1632 1022
rect 1576 954 1632 988
rect 1576 920 1587 954
rect 1621 920 1632 954
rect 1576 886 1632 920
rect 1576 852 1587 886
rect 1621 852 1632 886
rect 1576 818 1632 852
rect 1576 784 1587 818
rect 1621 784 1632 818
rect 1576 750 1632 784
rect 1576 716 1587 750
rect 1621 716 1632 750
rect 1576 682 1632 716
rect 1576 648 1587 682
rect 1621 648 1632 682
rect 1576 614 1632 648
rect 1576 580 1587 614
rect 1621 580 1632 614
rect 1576 546 1632 580
rect 1576 512 1587 546
rect 1621 512 1632 546
rect 1576 478 1632 512
rect 1576 444 1587 478
rect 1621 444 1632 478
rect 1576 410 1632 444
rect 1576 376 1587 410
rect 1621 376 1632 410
rect 1576 342 1632 376
rect 1576 308 1587 342
rect 1621 308 1632 342
rect 1576 274 1632 308
rect 1576 240 1587 274
rect 1621 240 1632 274
rect 1576 206 1632 240
rect 1576 172 1587 206
rect 1621 172 1632 206
rect 1576 138 1632 172
rect 1576 104 1587 138
rect 1621 104 1632 138
rect 1576 92 1632 104
rect 1732 1498 1788 1510
rect 1732 1464 1743 1498
rect 1777 1464 1788 1498
rect 1732 1430 1788 1464
rect 1732 1396 1743 1430
rect 1777 1396 1788 1430
rect 1732 1362 1788 1396
rect 1732 1328 1743 1362
rect 1777 1328 1788 1362
rect 1732 1294 1788 1328
rect 1732 1260 1743 1294
rect 1777 1260 1788 1294
rect 1732 1226 1788 1260
rect 1732 1192 1743 1226
rect 1777 1192 1788 1226
rect 1732 1158 1788 1192
rect 1732 1124 1743 1158
rect 1777 1124 1788 1158
rect 1732 1090 1788 1124
rect 1732 1056 1743 1090
rect 1777 1056 1788 1090
rect 1732 1022 1788 1056
rect 1732 988 1743 1022
rect 1777 988 1788 1022
rect 1732 954 1788 988
rect 1732 920 1743 954
rect 1777 920 1788 954
rect 1732 886 1788 920
rect 1732 852 1743 886
rect 1777 852 1788 886
rect 1732 818 1788 852
rect 1732 784 1743 818
rect 1777 784 1788 818
rect 1732 750 1788 784
rect 1732 716 1743 750
rect 1777 716 1788 750
rect 1732 682 1788 716
rect 1732 648 1743 682
rect 1777 648 1788 682
rect 1732 614 1788 648
rect 1732 580 1743 614
rect 1777 580 1788 614
rect 1732 546 1788 580
rect 1732 512 1743 546
rect 1777 512 1788 546
rect 1732 478 1788 512
rect 1732 444 1743 478
rect 1777 444 1788 478
rect 1732 410 1788 444
rect 1732 376 1743 410
rect 1777 376 1788 410
rect 1732 342 1788 376
rect 1732 308 1743 342
rect 1777 308 1788 342
rect 1732 274 1788 308
rect 1732 240 1743 274
rect 1777 240 1788 274
rect 1732 206 1788 240
rect 1732 172 1743 206
rect 1777 172 1788 206
rect 1732 138 1788 172
rect 1732 104 1743 138
rect 1777 104 1788 138
rect 1732 92 1788 104
<< mvndiffc >>
rect 183 1464 217 1498
rect 183 1396 217 1430
rect 183 1328 217 1362
rect 183 1260 217 1294
rect 183 1192 217 1226
rect 183 1124 217 1158
rect 183 1056 217 1090
rect 183 988 217 1022
rect 183 920 217 954
rect 183 852 217 886
rect 183 784 217 818
rect 183 716 217 750
rect 183 648 217 682
rect 183 580 217 614
rect 183 512 217 546
rect 183 444 217 478
rect 183 376 217 410
rect 183 308 217 342
rect 183 240 217 274
rect 183 172 217 206
rect 183 104 217 138
rect 339 1464 373 1498
rect 339 1396 373 1430
rect 339 1328 373 1362
rect 339 1260 373 1294
rect 339 1192 373 1226
rect 339 1124 373 1158
rect 339 1056 373 1090
rect 339 988 373 1022
rect 339 920 373 954
rect 339 852 373 886
rect 339 784 373 818
rect 339 716 373 750
rect 339 648 373 682
rect 339 580 373 614
rect 339 512 373 546
rect 339 444 373 478
rect 339 376 373 410
rect 339 308 373 342
rect 339 240 373 274
rect 339 172 373 206
rect 339 104 373 138
rect 495 1464 529 1498
rect 495 1396 529 1430
rect 495 1328 529 1362
rect 495 1260 529 1294
rect 495 1192 529 1226
rect 495 1124 529 1158
rect 495 1056 529 1090
rect 495 988 529 1022
rect 495 920 529 954
rect 495 852 529 886
rect 495 784 529 818
rect 495 716 529 750
rect 495 648 529 682
rect 495 580 529 614
rect 495 512 529 546
rect 495 444 529 478
rect 495 376 529 410
rect 495 308 529 342
rect 495 240 529 274
rect 495 172 529 206
rect 495 104 529 138
rect 651 1464 685 1498
rect 651 1396 685 1430
rect 651 1328 685 1362
rect 651 1260 685 1294
rect 651 1192 685 1226
rect 651 1124 685 1158
rect 651 1056 685 1090
rect 651 988 685 1022
rect 651 920 685 954
rect 651 852 685 886
rect 651 784 685 818
rect 651 716 685 750
rect 651 648 685 682
rect 651 580 685 614
rect 651 512 685 546
rect 651 444 685 478
rect 651 376 685 410
rect 651 308 685 342
rect 651 240 685 274
rect 651 172 685 206
rect 651 104 685 138
rect 807 1464 841 1498
rect 807 1396 841 1430
rect 807 1328 841 1362
rect 807 1260 841 1294
rect 807 1192 841 1226
rect 807 1124 841 1158
rect 807 1056 841 1090
rect 807 988 841 1022
rect 807 920 841 954
rect 807 852 841 886
rect 807 784 841 818
rect 807 716 841 750
rect 807 648 841 682
rect 807 580 841 614
rect 807 512 841 546
rect 807 444 841 478
rect 807 376 841 410
rect 807 308 841 342
rect 807 240 841 274
rect 807 172 841 206
rect 807 104 841 138
rect 963 1464 997 1498
rect 963 1396 997 1430
rect 963 1328 997 1362
rect 963 1260 997 1294
rect 963 1192 997 1226
rect 963 1124 997 1158
rect 963 1056 997 1090
rect 963 988 997 1022
rect 963 920 997 954
rect 963 852 997 886
rect 963 784 997 818
rect 963 716 997 750
rect 963 648 997 682
rect 963 580 997 614
rect 963 512 997 546
rect 963 444 997 478
rect 963 376 997 410
rect 963 308 997 342
rect 963 240 997 274
rect 963 172 997 206
rect 963 104 997 138
rect 1119 1464 1153 1498
rect 1119 1396 1153 1430
rect 1119 1328 1153 1362
rect 1119 1260 1153 1294
rect 1119 1192 1153 1226
rect 1119 1124 1153 1158
rect 1119 1056 1153 1090
rect 1119 988 1153 1022
rect 1119 920 1153 954
rect 1119 852 1153 886
rect 1119 784 1153 818
rect 1119 716 1153 750
rect 1119 648 1153 682
rect 1119 580 1153 614
rect 1119 512 1153 546
rect 1119 444 1153 478
rect 1119 376 1153 410
rect 1119 308 1153 342
rect 1119 240 1153 274
rect 1119 172 1153 206
rect 1119 104 1153 138
rect 1275 1464 1309 1498
rect 1275 1396 1309 1430
rect 1275 1328 1309 1362
rect 1275 1260 1309 1294
rect 1275 1192 1309 1226
rect 1275 1124 1309 1158
rect 1275 1056 1309 1090
rect 1275 988 1309 1022
rect 1275 920 1309 954
rect 1275 852 1309 886
rect 1275 784 1309 818
rect 1275 716 1309 750
rect 1275 648 1309 682
rect 1275 580 1309 614
rect 1275 512 1309 546
rect 1275 444 1309 478
rect 1275 376 1309 410
rect 1275 308 1309 342
rect 1275 240 1309 274
rect 1275 172 1309 206
rect 1275 104 1309 138
rect 1431 1464 1465 1498
rect 1431 1396 1465 1430
rect 1431 1328 1465 1362
rect 1431 1260 1465 1294
rect 1431 1192 1465 1226
rect 1431 1124 1465 1158
rect 1431 1056 1465 1090
rect 1431 988 1465 1022
rect 1431 920 1465 954
rect 1431 852 1465 886
rect 1431 784 1465 818
rect 1431 716 1465 750
rect 1431 648 1465 682
rect 1431 580 1465 614
rect 1431 512 1465 546
rect 1431 444 1465 478
rect 1431 376 1465 410
rect 1431 308 1465 342
rect 1431 240 1465 274
rect 1431 172 1465 206
rect 1431 104 1465 138
rect 1587 1464 1621 1498
rect 1587 1396 1621 1430
rect 1587 1328 1621 1362
rect 1587 1260 1621 1294
rect 1587 1192 1621 1226
rect 1587 1124 1621 1158
rect 1587 1056 1621 1090
rect 1587 988 1621 1022
rect 1587 920 1621 954
rect 1587 852 1621 886
rect 1587 784 1621 818
rect 1587 716 1621 750
rect 1587 648 1621 682
rect 1587 580 1621 614
rect 1587 512 1621 546
rect 1587 444 1621 478
rect 1587 376 1621 410
rect 1587 308 1621 342
rect 1587 240 1621 274
rect 1587 172 1621 206
rect 1587 104 1621 138
rect 1743 1464 1777 1498
rect 1743 1396 1777 1430
rect 1743 1328 1777 1362
rect 1743 1260 1777 1294
rect 1743 1192 1777 1226
rect 1743 1124 1777 1158
rect 1743 1056 1777 1090
rect 1743 988 1777 1022
rect 1743 920 1777 954
rect 1743 852 1777 886
rect 1743 784 1777 818
rect 1743 716 1777 750
rect 1743 648 1777 682
rect 1743 580 1777 614
rect 1743 512 1777 546
rect 1743 444 1777 478
rect 1743 376 1777 410
rect 1743 308 1777 342
rect 1743 240 1777 274
rect 1743 172 1777 206
rect 1743 104 1777 138
<< mvpsubdiff >>
rect 36 1464 94 1510
rect 36 1430 48 1464
rect 82 1430 94 1464
rect 36 1396 94 1430
rect 36 1362 48 1396
rect 82 1362 94 1396
rect 36 1328 94 1362
rect 36 1294 48 1328
rect 82 1294 94 1328
rect 36 1260 94 1294
rect 36 1226 48 1260
rect 82 1226 94 1260
rect 36 1192 94 1226
rect 36 1158 48 1192
rect 82 1158 94 1192
rect 36 1124 94 1158
rect 36 1090 48 1124
rect 82 1090 94 1124
rect 36 1056 94 1090
rect 36 1022 48 1056
rect 82 1022 94 1056
rect 36 988 94 1022
rect 36 954 48 988
rect 82 954 94 988
rect 36 920 94 954
rect 36 886 48 920
rect 82 886 94 920
rect 36 852 94 886
rect 36 818 48 852
rect 82 818 94 852
rect 36 784 94 818
rect 36 750 48 784
rect 82 750 94 784
rect 36 716 94 750
rect 36 682 48 716
rect 82 682 94 716
rect 36 648 94 682
rect 36 614 48 648
rect 82 614 94 648
rect 36 580 94 614
rect 36 546 48 580
rect 82 546 94 580
rect 36 512 94 546
rect 36 478 48 512
rect 82 478 94 512
rect 36 444 94 478
rect 36 410 48 444
rect 82 410 94 444
rect 36 376 94 410
rect 36 342 48 376
rect 82 342 94 376
rect 36 308 94 342
rect 36 274 48 308
rect 82 274 94 308
rect 36 240 94 274
rect 36 206 48 240
rect 82 206 94 240
rect 36 172 94 206
rect 36 138 48 172
rect 82 138 94 172
rect 36 92 94 138
rect 1866 1464 1924 1510
rect 1866 1430 1878 1464
rect 1912 1430 1924 1464
rect 1866 1396 1924 1430
rect 1866 1362 1878 1396
rect 1912 1362 1924 1396
rect 1866 1328 1924 1362
rect 1866 1294 1878 1328
rect 1912 1294 1924 1328
rect 1866 1260 1924 1294
rect 1866 1226 1878 1260
rect 1912 1226 1924 1260
rect 1866 1192 1924 1226
rect 1866 1158 1878 1192
rect 1912 1158 1924 1192
rect 1866 1124 1924 1158
rect 1866 1090 1878 1124
rect 1912 1090 1924 1124
rect 1866 1056 1924 1090
rect 1866 1022 1878 1056
rect 1912 1022 1924 1056
rect 1866 988 1924 1022
rect 1866 954 1878 988
rect 1912 954 1924 988
rect 1866 920 1924 954
rect 1866 886 1878 920
rect 1912 886 1924 920
rect 1866 852 1924 886
rect 1866 818 1878 852
rect 1912 818 1924 852
rect 1866 784 1924 818
rect 1866 750 1878 784
rect 1912 750 1924 784
rect 1866 716 1924 750
rect 1866 682 1878 716
rect 1912 682 1924 716
rect 1866 648 1924 682
rect 1866 614 1878 648
rect 1912 614 1924 648
rect 1866 580 1924 614
rect 1866 546 1878 580
rect 1912 546 1924 580
rect 1866 512 1924 546
rect 1866 478 1878 512
rect 1912 478 1924 512
rect 1866 444 1924 478
rect 1866 410 1878 444
rect 1912 410 1924 444
rect 1866 376 1924 410
rect 1866 342 1878 376
rect 1912 342 1924 376
rect 1866 308 1924 342
rect 1866 274 1878 308
rect 1912 274 1924 308
rect 1866 240 1924 274
rect 1866 206 1878 240
rect 1912 206 1924 240
rect 1866 172 1924 206
rect 1866 138 1878 172
rect 1912 138 1924 172
rect 1866 92 1924 138
<< mvpsubdiffcont >>
rect 48 1430 82 1464
rect 48 1362 82 1396
rect 48 1294 82 1328
rect 48 1226 82 1260
rect 48 1158 82 1192
rect 48 1090 82 1124
rect 48 1022 82 1056
rect 48 954 82 988
rect 48 886 82 920
rect 48 818 82 852
rect 48 750 82 784
rect 48 682 82 716
rect 48 614 82 648
rect 48 546 82 580
rect 48 478 82 512
rect 48 410 82 444
rect 48 342 82 376
rect 48 274 82 308
rect 48 206 82 240
rect 48 138 82 172
rect 1878 1430 1912 1464
rect 1878 1362 1912 1396
rect 1878 1294 1912 1328
rect 1878 1226 1912 1260
rect 1878 1158 1912 1192
rect 1878 1090 1912 1124
rect 1878 1022 1912 1056
rect 1878 954 1912 988
rect 1878 886 1912 920
rect 1878 818 1912 852
rect 1878 750 1912 784
rect 1878 682 1912 716
rect 1878 614 1912 648
rect 1878 546 1912 580
rect 1878 478 1912 512
rect 1878 410 1912 444
rect 1878 342 1912 376
rect 1878 274 1912 308
rect 1878 206 1912 240
rect 1878 138 1912 172
<< poly >>
rect 199 1582 1761 1602
rect 199 1548 215 1582
rect 249 1548 283 1582
rect 317 1548 351 1582
rect 385 1548 419 1582
rect 453 1548 487 1582
rect 521 1548 555 1582
rect 589 1548 623 1582
rect 657 1548 691 1582
rect 725 1548 759 1582
rect 793 1548 827 1582
rect 861 1548 895 1582
rect 929 1548 963 1582
rect 997 1548 1031 1582
rect 1065 1548 1099 1582
rect 1133 1548 1167 1582
rect 1201 1548 1235 1582
rect 1269 1548 1303 1582
rect 1337 1548 1371 1582
rect 1405 1548 1439 1582
rect 1473 1548 1507 1582
rect 1541 1548 1575 1582
rect 1609 1548 1643 1582
rect 1677 1548 1711 1582
rect 1745 1548 1761 1582
rect 199 1532 1761 1548
rect 228 1510 328 1532
rect 384 1510 484 1532
rect 540 1510 640 1532
rect 696 1510 796 1532
rect 852 1510 952 1532
rect 1008 1510 1108 1532
rect 1164 1510 1264 1532
rect 1320 1510 1420 1532
rect 1476 1510 1576 1532
rect 1632 1510 1732 1532
rect 228 70 328 92
rect 384 70 484 92
rect 540 70 640 92
rect 696 70 796 92
rect 852 70 952 92
rect 1008 70 1108 92
rect 1164 70 1264 92
rect 1320 70 1420 92
rect 1476 70 1576 92
rect 1632 70 1732 92
rect 199 54 1761 70
rect 199 20 215 54
rect 249 20 283 54
rect 317 20 351 54
rect 385 20 419 54
rect 453 20 487 54
rect 521 20 555 54
rect 589 20 623 54
rect 657 20 691 54
rect 725 20 759 54
rect 793 20 827 54
rect 861 20 895 54
rect 929 20 963 54
rect 997 20 1031 54
rect 1065 20 1099 54
rect 1133 20 1167 54
rect 1201 20 1235 54
rect 1269 20 1303 54
rect 1337 20 1371 54
rect 1405 20 1439 54
rect 1473 20 1507 54
rect 1541 20 1575 54
rect 1609 20 1643 54
rect 1677 20 1711 54
rect 1745 20 1761 54
rect 199 0 1761 20
<< polycont >>
rect 215 1548 249 1582
rect 283 1548 317 1582
rect 351 1548 385 1582
rect 419 1548 453 1582
rect 487 1548 521 1582
rect 555 1548 589 1582
rect 623 1548 657 1582
rect 691 1548 725 1582
rect 759 1548 793 1582
rect 827 1548 861 1582
rect 895 1548 929 1582
rect 963 1548 997 1582
rect 1031 1548 1065 1582
rect 1099 1548 1133 1582
rect 1167 1548 1201 1582
rect 1235 1548 1269 1582
rect 1303 1548 1337 1582
rect 1371 1548 1405 1582
rect 1439 1548 1473 1582
rect 1507 1548 1541 1582
rect 1575 1548 1609 1582
rect 1643 1548 1677 1582
rect 1711 1548 1745 1582
rect 215 20 249 54
rect 283 20 317 54
rect 351 20 385 54
rect 419 20 453 54
rect 487 20 521 54
rect 555 20 589 54
rect 623 20 657 54
rect 691 20 725 54
rect 759 20 793 54
rect 827 20 861 54
rect 895 20 929 54
rect 963 20 997 54
rect 1031 20 1065 54
rect 1099 20 1133 54
rect 1167 20 1201 54
rect 1235 20 1269 54
rect 1303 20 1337 54
rect 1371 20 1405 54
rect 1439 20 1473 54
rect 1507 20 1541 54
rect 1575 20 1609 54
rect 1643 20 1677 54
rect 1711 20 1745 54
<< locali >>
rect 199 1548 207 1582
rect 249 1548 279 1582
rect 317 1548 351 1582
rect 385 1548 419 1582
rect 457 1548 487 1582
rect 529 1548 555 1582
rect 601 1548 623 1582
rect 673 1548 691 1582
rect 745 1548 759 1582
rect 817 1548 827 1582
rect 889 1548 895 1582
rect 961 1548 963 1582
rect 997 1548 999 1582
rect 1065 1548 1071 1582
rect 1133 1548 1143 1582
rect 1201 1548 1215 1582
rect 1269 1548 1287 1582
rect 1337 1548 1359 1582
rect 1405 1548 1431 1582
rect 1473 1548 1503 1582
rect 1541 1548 1575 1582
rect 1609 1548 1643 1582
rect 1681 1548 1711 1582
rect 1753 1548 1761 1582
rect 48 1466 82 1514
rect 48 1396 82 1430
rect 48 1328 82 1360
rect 48 1260 82 1288
rect 48 1192 82 1216
rect 48 1124 82 1144
rect 48 1056 82 1072
rect 48 988 82 1000
rect 48 920 82 928
rect 48 852 82 856
rect 48 746 82 750
rect 48 674 82 682
rect 48 602 82 614
rect 48 530 82 546
rect 48 458 82 478
rect 48 386 82 410
rect 48 314 82 342
rect 48 242 82 274
rect 48 172 82 206
rect 48 88 82 136
rect 183 1498 217 1514
rect 183 1430 217 1432
rect 183 1394 217 1396
rect 183 1322 217 1328
rect 183 1250 217 1260
rect 183 1178 217 1192
rect 183 1106 217 1124
rect 183 1034 217 1056
rect 183 962 217 988
rect 183 890 217 920
rect 183 818 217 852
rect 183 750 217 784
rect 183 682 217 712
rect 183 614 217 640
rect 183 546 217 568
rect 183 478 217 496
rect 183 410 217 424
rect 183 342 217 352
rect 183 274 217 280
rect 183 206 217 208
rect 183 170 217 172
rect 183 88 217 104
rect 339 1498 373 1514
rect 339 1430 373 1432
rect 339 1394 373 1396
rect 339 1322 373 1328
rect 339 1250 373 1260
rect 339 1178 373 1192
rect 339 1106 373 1124
rect 339 1034 373 1056
rect 339 962 373 988
rect 339 890 373 920
rect 339 818 373 852
rect 339 750 373 784
rect 339 682 373 712
rect 339 614 373 640
rect 339 546 373 568
rect 339 478 373 496
rect 339 410 373 424
rect 339 342 373 352
rect 339 274 373 280
rect 339 206 373 208
rect 339 170 373 172
rect 339 88 373 104
rect 495 1498 529 1514
rect 495 1430 529 1432
rect 495 1394 529 1396
rect 495 1322 529 1328
rect 495 1250 529 1260
rect 495 1178 529 1192
rect 495 1106 529 1124
rect 495 1034 529 1056
rect 495 962 529 988
rect 495 890 529 920
rect 495 818 529 852
rect 495 750 529 784
rect 495 682 529 712
rect 495 614 529 640
rect 495 546 529 568
rect 495 478 529 496
rect 495 410 529 424
rect 495 342 529 352
rect 495 274 529 280
rect 495 206 529 208
rect 495 170 529 172
rect 495 88 529 104
rect 651 1498 685 1514
rect 651 1430 685 1432
rect 651 1394 685 1396
rect 651 1322 685 1328
rect 651 1250 685 1260
rect 651 1178 685 1192
rect 651 1106 685 1124
rect 651 1034 685 1056
rect 651 962 685 988
rect 651 890 685 920
rect 651 818 685 852
rect 651 750 685 784
rect 651 682 685 712
rect 651 614 685 640
rect 651 546 685 568
rect 651 478 685 496
rect 651 410 685 424
rect 651 342 685 352
rect 651 274 685 280
rect 651 206 685 208
rect 651 170 685 172
rect 651 88 685 104
rect 807 1498 841 1514
rect 807 1430 841 1432
rect 807 1394 841 1396
rect 807 1322 841 1328
rect 807 1250 841 1260
rect 807 1178 841 1192
rect 807 1106 841 1124
rect 807 1034 841 1056
rect 807 962 841 988
rect 807 890 841 920
rect 807 818 841 852
rect 807 750 841 784
rect 807 682 841 712
rect 807 614 841 640
rect 807 546 841 568
rect 807 478 841 496
rect 807 410 841 424
rect 807 342 841 352
rect 807 274 841 280
rect 807 206 841 208
rect 807 170 841 172
rect 807 88 841 104
rect 963 1498 997 1514
rect 963 1430 997 1432
rect 963 1394 997 1396
rect 963 1322 997 1328
rect 963 1250 997 1260
rect 963 1178 997 1192
rect 963 1106 997 1124
rect 963 1034 997 1056
rect 963 962 997 988
rect 963 890 997 920
rect 963 818 997 852
rect 963 750 997 784
rect 963 682 997 712
rect 963 614 997 640
rect 963 546 997 568
rect 963 478 997 496
rect 963 410 997 424
rect 963 342 997 352
rect 963 274 997 280
rect 963 206 997 208
rect 963 170 997 172
rect 963 88 997 104
rect 1119 1498 1153 1514
rect 1119 1430 1153 1432
rect 1119 1394 1153 1396
rect 1119 1322 1153 1328
rect 1119 1250 1153 1260
rect 1119 1178 1153 1192
rect 1119 1106 1153 1124
rect 1119 1034 1153 1056
rect 1119 962 1153 988
rect 1119 890 1153 920
rect 1119 818 1153 852
rect 1119 750 1153 784
rect 1119 682 1153 712
rect 1119 614 1153 640
rect 1119 546 1153 568
rect 1119 478 1153 496
rect 1119 410 1153 424
rect 1119 342 1153 352
rect 1119 274 1153 280
rect 1119 206 1153 208
rect 1119 170 1153 172
rect 1119 88 1153 104
rect 1275 1498 1309 1514
rect 1275 1430 1309 1432
rect 1275 1394 1309 1396
rect 1275 1322 1309 1328
rect 1275 1250 1309 1260
rect 1275 1178 1309 1192
rect 1275 1106 1309 1124
rect 1275 1034 1309 1056
rect 1275 962 1309 988
rect 1275 890 1309 920
rect 1275 818 1309 852
rect 1275 750 1309 784
rect 1275 682 1309 712
rect 1275 614 1309 640
rect 1275 546 1309 568
rect 1275 478 1309 496
rect 1275 410 1309 424
rect 1275 342 1309 352
rect 1275 274 1309 280
rect 1275 206 1309 208
rect 1275 170 1309 172
rect 1275 88 1309 104
rect 1431 1498 1465 1514
rect 1431 1430 1465 1432
rect 1431 1394 1465 1396
rect 1431 1322 1465 1328
rect 1431 1250 1465 1260
rect 1431 1178 1465 1192
rect 1431 1106 1465 1124
rect 1431 1034 1465 1056
rect 1431 962 1465 988
rect 1431 890 1465 920
rect 1431 818 1465 852
rect 1431 750 1465 784
rect 1431 682 1465 712
rect 1431 614 1465 640
rect 1431 546 1465 568
rect 1431 478 1465 496
rect 1431 410 1465 424
rect 1431 342 1465 352
rect 1431 274 1465 280
rect 1431 206 1465 208
rect 1431 170 1465 172
rect 1431 88 1465 104
rect 1587 1498 1621 1514
rect 1587 1430 1621 1432
rect 1587 1394 1621 1396
rect 1587 1322 1621 1328
rect 1587 1250 1621 1260
rect 1587 1178 1621 1192
rect 1587 1106 1621 1124
rect 1587 1034 1621 1056
rect 1587 962 1621 988
rect 1587 890 1621 920
rect 1587 818 1621 852
rect 1587 750 1621 784
rect 1587 682 1621 712
rect 1587 614 1621 640
rect 1587 546 1621 568
rect 1587 478 1621 496
rect 1587 410 1621 424
rect 1587 342 1621 352
rect 1587 274 1621 280
rect 1587 206 1621 208
rect 1587 170 1621 172
rect 1587 88 1621 104
rect 1743 1498 1777 1514
rect 1743 1430 1777 1432
rect 1743 1394 1777 1396
rect 1743 1322 1777 1328
rect 1743 1250 1777 1260
rect 1743 1178 1777 1192
rect 1743 1106 1777 1124
rect 1743 1034 1777 1056
rect 1743 962 1777 988
rect 1743 890 1777 920
rect 1743 818 1777 852
rect 1743 750 1777 784
rect 1743 682 1777 712
rect 1743 614 1777 640
rect 1743 546 1777 568
rect 1743 478 1777 496
rect 1743 410 1777 424
rect 1743 342 1777 352
rect 1743 274 1777 280
rect 1743 206 1777 208
rect 1743 170 1777 172
rect 1743 88 1777 104
rect 1878 1466 1912 1514
rect 1878 1396 1912 1430
rect 1878 1328 1912 1360
rect 1878 1260 1912 1288
rect 1878 1192 1912 1216
rect 1878 1124 1912 1144
rect 1878 1056 1912 1072
rect 1878 988 1912 1000
rect 1878 920 1912 928
rect 1878 852 1912 856
rect 1878 746 1912 750
rect 1878 674 1912 682
rect 1878 602 1912 614
rect 1878 530 1912 546
rect 1878 458 1912 478
rect 1878 386 1912 410
rect 1878 314 1912 342
rect 1878 242 1912 274
rect 1878 172 1912 206
rect 1878 88 1912 136
rect 199 20 207 54
rect 249 20 279 54
rect 317 20 351 54
rect 385 20 419 54
rect 457 20 487 54
rect 529 20 555 54
rect 601 20 623 54
rect 673 20 691 54
rect 745 20 759 54
rect 817 20 827 54
rect 889 20 895 54
rect 961 20 963 54
rect 997 20 999 54
rect 1065 20 1071 54
rect 1133 20 1143 54
rect 1201 20 1215 54
rect 1269 20 1287 54
rect 1337 20 1359 54
rect 1405 20 1431 54
rect 1473 20 1503 54
rect 1541 20 1575 54
rect 1609 20 1643 54
rect 1681 20 1711 54
rect 1753 20 1761 54
<< viali >>
rect 207 1548 215 1582
rect 215 1548 241 1582
rect 279 1548 283 1582
rect 283 1548 313 1582
rect 351 1548 385 1582
rect 423 1548 453 1582
rect 453 1548 457 1582
rect 495 1548 521 1582
rect 521 1548 529 1582
rect 567 1548 589 1582
rect 589 1548 601 1582
rect 639 1548 657 1582
rect 657 1548 673 1582
rect 711 1548 725 1582
rect 725 1548 745 1582
rect 783 1548 793 1582
rect 793 1548 817 1582
rect 855 1548 861 1582
rect 861 1548 889 1582
rect 927 1548 929 1582
rect 929 1548 961 1582
rect 999 1548 1031 1582
rect 1031 1548 1033 1582
rect 1071 1548 1099 1582
rect 1099 1548 1105 1582
rect 1143 1548 1167 1582
rect 1167 1548 1177 1582
rect 1215 1548 1235 1582
rect 1235 1548 1249 1582
rect 1287 1548 1303 1582
rect 1303 1548 1321 1582
rect 1359 1548 1371 1582
rect 1371 1548 1393 1582
rect 1431 1548 1439 1582
rect 1439 1548 1465 1582
rect 1503 1548 1507 1582
rect 1507 1548 1537 1582
rect 1575 1548 1609 1582
rect 1647 1548 1677 1582
rect 1677 1548 1681 1582
rect 1719 1548 1745 1582
rect 1745 1548 1753 1582
rect 48 1464 82 1466
rect 48 1432 82 1464
rect 48 1362 82 1394
rect 48 1360 82 1362
rect 48 1294 82 1322
rect 48 1288 82 1294
rect 48 1226 82 1250
rect 48 1216 82 1226
rect 48 1158 82 1178
rect 48 1144 82 1158
rect 48 1090 82 1106
rect 48 1072 82 1090
rect 48 1022 82 1034
rect 48 1000 82 1022
rect 48 954 82 962
rect 48 928 82 954
rect 48 886 82 890
rect 48 856 82 886
rect 48 784 82 818
rect 48 716 82 746
rect 48 712 82 716
rect 48 648 82 674
rect 48 640 82 648
rect 48 580 82 602
rect 48 568 82 580
rect 48 512 82 530
rect 48 496 82 512
rect 48 444 82 458
rect 48 424 82 444
rect 48 376 82 386
rect 48 352 82 376
rect 48 308 82 314
rect 48 280 82 308
rect 48 240 82 242
rect 48 208 82 240
rect 48 138 82 170
rect 48 136 82 138
rect 183 1464 217 1466
rect 183 1432 217 1464
rect 183 1362 217 1394
rect 183 1360 217 1362
rect 183 1294 217 1322
rect 183 1288 217 1294
rect 183 1226 217 1250
rect 183 1216 217 1226
rect 183 1158 217 1178
rect 183 1144 217 1158
rect 183 1090 217 1106
rect 183 1072 217 1090
rect 183 1022 217 1034
rect 183 1000 217 1022
rect 183 954 217 962
rect 183 928 217 954
rect 183 886 217 890
rect 183 856 217 886
rect 183 784 217 818
rect 183 716 217 746
rect 183 712 217 716
rect 183 648 217 674
rect 183 640 217 648
rect 183 580 217 602
rect 183 568 217 580
rect 183 512 217 530
rect 183 496 217 512
rect 183 444 217 458
rect 183 424 217 444
rect 183 376 217 386
rect 183 352 217 376
rect 183 308 217 314
rect 183 280 217 308
rect 183 240 217 242
rect 183 208 217 240
rect 183 138 217 170
rect 183 136 217 138
rect 339 1464 373 1466
rect 339 1432 373 1464
rect 339 1362 373 1394
rect 339 1360 373 1362
rect 339 1294 373 1322
rect 339 1288 373 1294
rect 339 1226 373 1250
rect 339 1216 373 1226
rect 339 1158 373 1178
rect 339 1144 373 1158
rect 339 1090 373 1106
rect 339 1072 373 1090
rect 339 1022 373 1034
rect 339 1000 373 1022
rect 339 954 373 962
rect 339 928 373 954
rect 339 886 373 890
rect 339 856 373 886
rect 339 784 373 818
rect 339 716 373 746
rect 339 712 373 716
rect 339 648 373 674
rect 339 640 373 648
rect 339 580 373 602
rect 339 568 373 580
rect 339 512 373 530
rect 339 496 373 512
rect 339 444 373 458
rect 339 424 373 444
rect 339 376 373 386
rect 339 352 373 376
rect 339 308 373 314
rect 339 280 373 308
rect 339 240 373 242
rect 339 208 373 240
rect 339 138 373 170
rect 339 136 373 138
rect 495 1464 529 1466
rect 495 1432 529 1464
rect 495 1362 529 1394
rect 495 1360 529 1362
rect 495 1294 529 1322
rect 495 1288 529 1294
rect 495 1226 529 1250
rect 495 1216 529 1226
rect 495 1158 529 1178
rect 495 1144 529 1158
rect 495 1090 529 1106
rect 495 1072 529 1090
rect 495 1022 529 1034
rect 495 1000 529 1022
rect 495 954 529 962
rect 495 928 529 954
rect 495 886 529 890
rect 495 856 529 886
rect 495 784 529 818
rect 495 716 529 746
rect 495 712 529 716
rect 495 648 529 674
rect 495 640 529 648
rect 495 580 529 602
rect 495 568 529 580
rect 495 512 529 530
rect 495 496 529 512
rect 495 444 529 458
rect 495 424 529 444
rect 495 376 529 386
rect 495 352 529 376
rect 495 308 529 314
rect 495 280 529 308
rect 495 240 529 242
rect 495 208 529 240
rect 495 138 529 170
rect 495 136 529 138
rect 651 1464 685 1466
rect 651 1432 685 1464
rect 651 1362 685 1394
rect 651 1360 685 1362
rect 651 1294 685 1322
rect 651 1288 685 1294
rect 651 1226 685 1250
rect 651 1216 685 1226
rect 651 1158 685 1178
rect 651 1144 685 1158
rect 651 1090 685 1106
rect 651 1072 685 1090
rect 651 1022 685 1034
rect 651 1000 685 1022
rect 651 954 685 962
rect 651 928 685 954
rect 651 886 685 890
rect 651 856 685 886
rect 651 784 685 818
rect 651 716 685 746
rect 651 712 685 716
rect 651 648 685 674
rect 651 640 685 648
rect 651 580 685 602
rect 651 568 685 580
rect 651 512 685 530
rect 651 496 685 512
rect 651 444 685 458
rect 651 424 685 444
rect 651 376 685 386
rect 651 352 685 376
rect 651 308 685 314
rect 651 280 685 308
rect 651 240 685 242
rect 651 208 685 240
rect 651 138 685 170
rect 651 136 685 138
rect 807 1464 841 1466
rect 807 1432 841 1464
rect 807 1362 841 1394
rect 807 1360 841 1362
rect 807 1294 841 1322
rect 807 1288 841 1294
rect 807 1226 841 1250
rect 807 1216 841 1226
rect 807 1158 841 1178
rect 807 1144 841 1158
rect 807 1090 841 1106
rect 807 1072 841 1090
rect 807 1022 841 1034
rect 807 1000 841 1022
rect 807 954 841 962
rect 807 928 841 954
rect 807 886 841 890
rect 807 856 841 886
rect 807 784 841 818
rect 807 716 841 746
rect 807 712 841 716
rect 807 648 841 674
rect 807 640 841 648
rect 807 580 841 602
rect 807 568 841 580
rect 807 512 841 530
rect 807 496 841 512
rect 807 444 841 458
rect 807 424 841 444
rect 807 376 841 386
rect 807 352 841 376
rect 807 308 841 314
rect 807 280 841 308
rect 807 240 841 242
rect 807 208 841 240
rect 807 138 841 170
rect 807 136 841 138
rect 963 1464 997 1466
rect 963 1432 997 1464
rect 963 1362 997 1394
rect 963 1360 997 1362
rect 963 1294 997 1322
rect 963 1288 997 1294
rect 963 1226 997 1250
rect 963 1216 997 1226
rect 963 1158 997 1178
rect 963 1144 997 1158
rect 963 1090 997 1106
rect 963 1072 997 1090
rect 963 1022 997 1034
rect 963 1000 997 1022
rect 963 954 997 962
rect 963 928 997 954
rect 963 886 997 890
rect 963 856 997 886
rect 963 784 997 818
rect 963 716 997 746
rect 963 712 997 716
rect 963 648 997 674
rect 963 640 997 648
rect 963 580 997 602
rect 963 568 997 580
rect 963 512 997 530
rect 963 496 997 512
rect 963 444 997 458
rect 963 424 997 444
rect 963 376 997 386
rect 963 352 997 376
rect 963 308 997 314
rect 963 280 997 308
rect 963 240 997 242
rect 963 208 997 240
rect 963 138 997 170
rect 963 136 997 138
rect 1119 1464 1153 1466
rect 1119 1432 1153 1464
rect 1119 1362 1153 1394
rect 1119 1360 1153 1362
rect 1119 1294 1153 1322
rect 1119 1288 1153 1294
rect 1119 1226 1153 1250
rect 1119 1216 1153 1226
rect 1119 1158 1153 1178
rect 1119 1144 1153 1158
rect 1119 1090 1153 1106
rect 1119 1072 1153 1090
rect 1119 1022 1153 1034
rect 1119 1000 1153 1022
rect 1119 954 1153 962
rect 1119 928 1153 954
rect 1119 886 1153 890
rect 1119 856 1153 886
rect 1119 784 1153 818
rect 1119 716 1153 746
rect 1119 712 1153 716
rect 1119 648 1153 674
rect 1119 640 1153 648
rect 1119 580 1153 602
rect 1119 568 1153 580
rect 1119 512 1153 530
rect 1119 496 1153 512
rect 1119 444 1153 458
rect 1119 424 1153 444
rect 1119 376 1153 386
rect 1119 352 1153 376
rect 1119 308 1153 314
rect 1119 280 1153 308
rect 1119 240 1153 242
rect 1119 208 1153 240
rect 1119 138 1153 170
rect 1119 136 1153 138
rect 1275 1464 1309 1466
rect 1275 1432 1309 1464
rect 1275 1362 1309 1394
rect 1275 1360 1309 1362
rect 1275 1294 1309 1322
rect 1275 1288 1309 1294
rect 1275 1226 1309 1250
rect 1275 1216 1309 1226
rect 1275 1158 1309 1178
rect 1275 1144 1309 1158
rect 1275 1090 1309 1106
rect 1275 1072 1309 1090
rect 1275 1022 1309 1034
rect 1275 1000 1309 1022
rect 1275 954 1309 962
rect 1275 928 1309 954
rect 1275 886 1309 890
rect 1275 856 1309 886
rect 1275 784 1309 818
rect 1275 716 1309 746
rect 1275 712 1309 716
rect 1275 648 1309 674
rect 1275 640 1309 648
rect 1275 580 1309 602
rect 1275 568 1309 580
rect 1275 512 1309 530
rect 1275 496 1309 512
rect 1275 444 1309 458
rect 1275 424 1309 444
rect 1275 376 1309 386
rect 1275 352 1309 376
rect 1275 308 1309 314
rect 1275 280 1309 308
rect 1275 240 1309 242
rect 1275 208 1309 240
rect 1275 138 1309 170
rect 1275 136 1309 138
rect 1431 1464 1465 1466
rect 1431 1432 1465 1464
rect 1431 1362 1465 1394
rect 1431 1360 1465 1362
rect 1431 1294 1465 1322
rect 1431 1288 1465 1294
rect 1431 1226 1465 1250
rect 1431 1216 1465 1226
rect 1431 1158 1465 1178
rect 1431 1144 1465 1158
rect 1431 1090 1465 1106
rect 1431 1072 1465 1090
rect 1431 1022 1465 1034
rect 1431 1000 1465 1022
rect 1431 954 1465 962
rect 1431 928 1465 954
rect 1431 886 1465 890
rect 1431 856 1465 886
rect 1431 784 1465 818
rect 1431 716 1465 746
rect 1431 712 1465 716
rect 1431 648 1465 674
rect 1431 640 1465 648
rect 1431 580 1465 602
rect 1431 568 1465 580
rect 1431 512 1465 530
rect 1431 496 1465 512
rect 1431 444 1465 458
rect 1431 424 1465 444
rect 1431 376 1465 386
rect 1431 352 1465 376
rect 1431 308 1465 314
rect 1431 280 1465 308
rect 1431 240 1465 242
rect 1431 208 1465 240
rect 1431 138 1465 170
rect 1431 136 1465 138
rect 1587 1464 1621 1466
rect 1587 1432 1621 1464
rect 1587 1362 1621 1394
rect 1587 1360 1621 1362
rect 1587 1294 1621 1322
rect 1587 1288 1621 1294
rect 1587 1226 1621 1250
rect 1587 1216 1621 1226
rect 1587 1158 1621 1178
rect 1587 1144 1621 1158
rect 1587 1090 1621 1106
rect 1587 1072 1621 1090
rect 1587 1022 1621 1034
rect 1587 1000 1621 1022
rect 1587 954 1621 962
rect 1587 928 1621 954
rect 1587 886 1621 890
rect 1587 856 1621 886
rect 1587 784 1621 818
rect 1587 716 1621 746
rect 1587 712 1621 716
rect 1587 648 1621 674
rect 1587 640 1621 648
rect 1587 580 1621 602
rect 1587 568 1621 580
rect 1587 512 1621 530
rect 1587 496 1621 512
rect 1587 444 1621 458
rect 1587 424 1621 444
rect 1587 376 1621 386
rect 1587 352 1621 376
rect 1587 308 1621 314
rect 1587 280 1621 308
rect 1587 240 1621 242
rect 1587 208 1621 240
rect 1587 138 1621 170
rect 1587 136 1621 138
rect 1743 1464 1777 1466
rect 1743 1432 1777 1464
rect 1743 1362 1777 1394
rect 1743 1360 1777 1362
rect 1743 1294 1777 1322
rect 1743 1288 1777 1294
rect 1743 1226 1777 1250
rect 1743 1216 1777 1226
rect 1743 1158 1777 1178
rect 1743 1144 1777 1158
rect 1743 1090 1777 1106
rect 1743 1072 1777 1090
rect 1743 1022 1777 1034
rect 1743 1000 1777 1022
rect 1743 954 1777 962
rect 1743 928 1777 954
rect 1743 886 1777 890
rect 1743 856 1777 886
rect 1743 784 1777 818
rect 1743 716 1777 746
rect 1743 712 1777 716
rect 1743 648 1777 674
rect 1743 640 1777 648
rect 1743 580 1777 602
rect 1743 568 1777 580
rect 1743 512 1777 530
rect 1743 496 1777 512
rect 1743 444 1777 458
rect 1743 424 1777 444
rect 1743 376 1777 386
rect 1743 352 1777 376
rect 1743 308 1777 314
rect 1743 280 1777 308
rect 1743 240 1777 242
rect 1743 208 1777 240
rect 1743 138 1777 170
rect 1743 136 1777 138
rect 1878 1464 1912 1466
rect 1878 1432 1912 1464
rect 1878 1362 1912 1394
rect 1878 1360 1912 1362
rect 1878 1294 1912 1322
rect 1878 1288 1912 1294
rect 1878 1226 1912 1250
rect 1878 1216 1912 1226
rect 1878 1158 1912 1178
rect 1878 1144 1912 1158
rect 1878 1090 1912 1106
rect 1878 1072 1912 1090
rect 1878 1022 1912 1034
rect 1878 1000 1912 1022
rect 1878 954 1912 962
rect 1878 928 1912 954
rect 1878 886 1912 890
rect 1878 856 1912 886
rect 1878 784 1912 818
rect 1878 716 1912 746
rect 1878 712 1912 716
rect 1878 648 1912 674
rect 1878 640 1912 648
rect 1878 580 1912 602
rect 1878 568 1912 580
rect 1878 512 1912 530
rect 1878 496 1912 512
rect 1878 444 1912 458
rect 1878 424 1912 444
rect 1878 376 1912 386
rect 1878 352 1912 376
rect 1878 308 1912 314
rect 1878 280 1912 308
rect 1878 240 1912 242
rect 1878 208 1912 240
rect 1878 138 1912 170
rect 1878 136 1912 138
rect 207 20 215 54
rect 215 20 241 54
rect 279 20 283 54
rect 283 20 313 54
rect 351 20 385 54
rect 423 20 453 54
rect 453 20 457 54
rect 495 20 521 54
rect 521 20 529 54
rect 567 20 589 54
rect 589 20 601 54
rect 639 20 657 54
rect 657 20 673 54
rect 711 20 725 54
rect 725 20 745 54
rect 783 20 793 54
rect 793 20 817 54
rect 855 20 861 54
rect 861 20 889 54
rect 927 20 929 54
rect 929 20 961 54
rect 999 20 1031 54
rect 1031 20 1033 54
rect 1071 20 1099 54
rect 1099 20 1105 54
rect 1143 20 1167 54
rect 1167 20 1177 54
rect 1215 20 1235 54
rect 1235 20 1249 54
rect 1287 20 1303 54
rect 1303 20 1321 54
rect 1359 20 1371 54
rect 1371 20 1393 54
rect 1431 20 1439 54
rect 1439 20 1465 54
rect 1503 20 1507 54
rect 1507 20 1537 54
rect 1575 20 1609 54
rect 1647 20 1677 54
rect 1677 20 1681 54
rect 1719 20 1745 54
rect 1745 20 1753 54
<< metal1 >>
rect 195 1582 1765 1602
rect 195 1548 207 1582
rect 241 1548 279 1582
rect 313 1548 351 1582
rect 385 1548 423 1582
rect 457 1548 495 1582
rect 529 1548 567 1582
rect 601 1548 639 1582
rect 673 1548 711 1582
rect 745 1548 783 1582
rect 817 1548 855 1582
rect 889 1548 927 1582
rect 961 1548 999 1582
rect 1033 1548 1071 1582
rect 1105 1548 1143 1582
rect 1177 1548 1215 1582
rect 1249 1548 1287 1582
rect 1321 1548 1359 1582
rect 1393 1548 1431 1582
rect 1465 1548 1503 1582
rect 1537 1548 1575 1582
rect 1609 1548 1647 1582
rect 1681 1548 1719 1582
rect 1753 1548 1765 1582
rect 195 1536 1765 1548
rect 36 1466 94 1497
rect 36 1432 48 1466
rect 82 1432 94 1466
rect 36 1394 94 1432
rect 36 1360 48 1394
rect 82 1360 94 1394
rect 36 1322 94 1360
rect 36 1288 48 1322
rect 82 1288 94 1322
rect 36 1250 94 1288
rect 36 1216 48 1250
rect 82 1216 94 1250
rect 36 1178 94 1216
rect 36 1144 48 1178
rect 82 1144 94 1178
rect 36 1106 94 1144
rect 36 1072 48 1106
rect 82 1072 94 1106
rect 36 1034 94 1072
rect 36 1000 48 1034
rect 82 1000 94 1034
rect 36 962 94 1000
rect 36 928 48 962
rect 82 928 94 962
rect 36 890 94 928
rect 36 856 48 890
rect 82 856 94 890
rect 36 818 94 856
rect 36 784 48 818
rect 82 784 94 818
rect 36 746 94 784
rect 36 712 48 746
rect 82 712 94 746
rect 36 674 94 712
rect 36 640 48 674
rect 82 640 94 674
rect 36 602 94 640
rect 36 568 48 602
rect 82 568 94 602
rect 36 530 94 568
rect 36 496 48 530
rect 82 496 94 530
rect 36 458 94 496
rect 36 424 48 458
rect 82 424 94 458
rect 36 386 94 424
rect 36 352 48 386
rect 82 352 94 386
rect 36 314 94 352
rect 36 280 48 314
rect 82 280 94 314
rect 36 242 94 280
rect 36 208 48 242
rect 82 208 94 242
rect 36 170 94 208
rect 36 136 48 170
rect 82 136 94 170
rect 36 105 94 136
rect 174 1491 226 1497
rect 174 1432 183 1439
rect 217 1432 226 1439
rect 174 1427 226 1432
rect 174 1363 183 1375
rect 217 1363 226 1375
rect 174 1299 183 1311
rect 217 1299 226 1311
rect 174 1235 183 1247
rect 217 1235 226 1247
rect 174 1178 226 1183
rect 174 1144 183 1178
rect 217 1144 226 1178
rect 174 1106 226 1144
rect 174 1072 183 1106
rect 217 1072 226 1106
rect 174 1034 226 1072
rect 174 1000 183 1034
rect 217 1000 226 1034
rect 174 962 226 1000
rect 174 928 183 962
rect 217 928 226 962
rect 174 890 226 928
rect 174 856 183 890
rect 217 856 226 890
rect 174 818 226 856
rect 174 784 183 818
rect 217 784 226 818
rect 174 746 226 784
rect 174 712 183 746
rect 217 712 226 746
rect 174 674 226 712
rect 174 640 183 674
rect 217 640 226 674
rect 174 602 226 640
rect 174 568 183 602
rect 217 568 226 602
rect 174 530 226 568
rect 174 496 183 530
rect 217 496 226 530
rect 174 458 226 496
rect 174 424 183 458
rect 217 424 226 458
rect 174 419 226 424
rect 174 355 183 367
rect 217 355 226 367
rect 174 291 183 303
rect 217 291 226 303
rect 174 227 183 239
rect 217 227 226 239
rect 174 170 226 175
rect 174 163 183 170
rect 217 163 226 170
rect 174 105 226 111
rect 330 1466 382 1497
rect 330 1432 339 1466
rect 373 1432 382 1466
rect 330 1394 382 1432
rect 330 1360 339 1394
rect 373 1360 382 1394
rect 330 1322 382 1360
rect 330 1288 339 1322
rect 373 1288 382 1322
rect 330 1250 382 1288
rect 330 1216 339 1250
rect 373 1216 382 1250
rect 330 1178 382 1216
rect 330 1144 339 1178
rect 373 1144 382 1178
rect 330 1115 382 1144
rect 330 1051 382 1063
rect 330 987 382 999
rect 330 928 339 935
rect 373 928 382 935
rect 330 923 382 928
rect 330 859 339 871
rect 373 859 382 871
rect 330 795 339 807
rect 373 795 382 807
rect 330 731 339 743
rect 373 731 382 743
rect 330 674 382 679
rect 330 667 339 674
rect 373 667 382 674
rect 330 603 382 615
rect 330 539 382 551
rect 330 458 382 487
rect 330 424 339 458
rect 373 424 382 458
rect 330 386 382 424
rect 330 352 339 386
rect 373 352 382 386
rect 330 314 382 352
rect 330 280 339 314
rect 373 280 382 314
rect 330 242 382 280
rect 330 208 339 242
rect 373 208 382 242
rect 330 170 382 208
rect 330 136 339 170
rect 373 136 382 170
rect 330 105 382 136
rect 486 1491 538 1497
rect 486 1432 495 1439
rect 529 1432 538 1439
rect 486 1427 538 1432
rect 486 1363 495 1375
rect 529 1363 538 1375
rect 486 1299 495 1311
rect 529 1299 538 1311
rect 486 1235 495 1247
rect 529 1235 538 1247
rect 486 1178 538 1183
rect 486 1144 495 1178
rect 529 1144 538 1178
rect 486 1106 538 1144
rect 486 1072 495 1106
rect 529 1072 538 1106
rect 486 1034 538 1072
rect 486 1000 495 1034
rect 529 1000 538 1034
rect 486 962 538 1000
rect 486 928 495 962
rect 529 928 538 962
rect 486 890 538 928
rect 486 856 495 890
rect 529 856 538 890
rect 486 818 538 856
rect 486 784 495 818
rect 529 784 538 818
rect 486 746 538 784
rect 486 712 495 746
rect 529 712 538 746
rect 486 674 538 712
rect 486 640 495 674
rect 529 640 538 674
rect 486 602 538 640
rect 486 568 495 602
rect 529 568 538 602
rect 486 530 538 568
rect 486 496 495 530
rect 529 496 538 530
rect 486 458 538 496
rect 486 424 495 458
rect 529 424 538 458
rect 486 419 538 424
rect 486 355 495 367
rect 529 355 538 367
rect 486 291 495 303
rect 529 291 538 303
rect 486 227 495 239
rect 529 227 538 239
rect 486 170 538 175
rect 486 163 495 170
rect 529 163 538 170
rect 486 105 538 111
rect 642 1466 694 1497
rect 642 1432 651 1466
rect 685 1432 694 1466
rect 642 1394 694 1432
rect 642 1360 651 1394
rect 685 1360 694 1394
rect 642 1322 694 1360
rect 642 1288 651 1322
rect 685 1288 694 1322
rect 642 1250 694 1288
rect 642 1216 651 1250
rect 685 1216 694 1250
rect 642 1178 694 1216
rect 642 1144 651 1178
rect 685 1144 694 1178
rect 642 1115 694 1144
rect 642 1051 694 1063
rect 642 987 694 999
rect 642 928 651 935
rect 685 928 694 935
rect 642 923 694 928
rect 642 859 651 871
rect 685 859 694 871
rect 642 795 651 807
rect 685 795 694 807
rect 642 731 651 743
rect 685 731 694 743
rect 642 674 694 679
rect 642 667 651 674
rect 685 667 694 674
rect 642 603 694 615
rect 642 539 694 551
rect 642 458 694 487
rect 642 424 651 458
rect 685 424 694 458
rect 642 386 694 424
rect 642 352 651 386
rect 685 352 694 386
rect 642 314 694 352
rect 642 280 651 314
rect 685 280 694 314
rect 642 242 694 280
rect 642 208 651 242
rect 685 208 694 242
rect 642 170 694 208
rect 642 136 651 170
rect 685 136 694 170
rect 642 105 694 136
rect 798 1491 850 1497
rect 798 1432 807 1439
rect 841 1432 850 1439
rect 798 1427 850 1432
rect 798 1363 807 1375
rect 841 1363 850 1375
rect 798 1299 807 1311
rect 841 1299 850 1311
rect 798 1235 807 1247
rect 841 1235 850 1247
rect 798 1178 850 1183
rect 798 1144 807 1178
rect 841 1144 850 1178
rect 798 1106 850 1144
rect 798 1072 807 1106
rect 841 1072 850 1106
rect 798 1034 850 1072
rect 798 1000 807 1034
rect 841 1000 850 1034
rect 798 962 850 1000
rect 798 928 807 962
rect 841 928 850 962
rect 798 890 850 928
rect 798 856 807 890
rect 841 856 850 890
rect 798 818 850 856
rect 798 784 807 818
rect 841 784 850 818
rect 798 746 850 784
rect 798 712 807 746
rect 841 712 850 746
rect 798 674 850 712
rect 798 640 807 674
rect 841 640 850 674
rect 798 602 850 640
rect 798 568 807 602
rect 841 568 850 602
rect 798 530 850 568
rect 798 496 807 530
rect 841 496 850 530
rect 798 458 850 496
rect 798 424 807 458
rect 841 424 850 458
rect 798 419 850 424
rect 798 355 807 367
rect 841 355 850 367
rect 798 291 807 303
rect 841 291 850 303
rect 798 227 807 239
rect 841 227 850 239
rect 798 170 850 175
rect 798 163 807 170
rect 841 163 850 170
rect 798 105 850 111
rect 954 1466 1006 1497
rect 954 1432 963 1466
rect 997 1432 1006 1466
rect 954 1394 1006 1432
rect 954 1360 963 1394
rect 997 1360 1006 1394
rect 954 1322 1006 1360
rect 954 1288 963 1322
rect 997 1288 1006 1322
rect 954 1250 1006 1288
rect 954 1216 963 1250
rect 997 1216 1006 1250
rect 954 1178 1006 1216
rect 954 1144 963 1178
rect 997 1144 1006 1178
rect 954 1115 1006 1144
rect 954 1051 1006 1063
rect 954 987 1006 999
rect 954 928 963 935
rect 997 928 1006 935
rect 954 923 1006 928
rect 954 859 963 871
rect 997 859 1006 871
rect 954 795 963 807
rect 997 795 1006 807
rect 954 731 963 743
rect 997 731 1006 743
rect 954 674 1006 679
rect 954 667 963 674
rect 997 667 1006 674
rect 954 603 1006 615
rect 954 539 1006 551
rect 954 458 1006 487
rect 954 424 963 458
rect 997 424 1006 458
rect 954 386 1006 424
rect 954 352 963 386
rect 997 352 1006 386
rect 954 314 1006 352
rect 954 280 963 314
rect 997 280 1006 314
rect 954 242 1006 280
rect 954 208 963 242
rect 997 208 1006 242
rect 954 170 1006 208
rect 954 136 963 170
rect 997 136 1006 170
rect 954 105 1006 136
rect 1110 1491 1162 1497
rect 1110 1432 1119 1439
rect 1153 1432 1162 1439
rect 1110 1427 1162 1432
rect 1110 1363 1119 1375
rect 1153 1363 1162 1375
rect 1110 1299 1119 1311
rect 1153 1299 1162 1311
rect 1110 1235 1119 1247
rect 1153 1235 1162 1247
rect 1110 1178 1162 1183
rect 1110 1144 1119 1178
rect 1153 1144 1162 1178
rect 1110 1106 1162 1144
rect 1110 1072 1119 1106
rect 1153 1072 1162 1106
rect 1110 1034 1162 1072
rect 1110 1000 1119 1034
rect 1153 1000 1162 1034
rect 1110 962 1162 1000
rect 1110 928 1119 962
rect 1153 928 1162 962
rect 1110 890 1162 928
rect 1110 856 1119 890
rect 1153 856 1162 890
rect 1110 818 1162 856
rect 1110 784 1119 818
rect 1153 784 1162 818
rect 1110 746 1162 784
rect 1110 712 1119 746
rect 1153 712 1162 746
rect 1110 674 1162 712
rect 1110 640 1119 674
rect 1153 640 1162 674
rect 1110 602 1162 640
rect 1110 568 1119 602
rect 1153 568 1162 602
rect 1110 530 1162 568
rect 1110 496 1119 530
rect 1153 496 1162 530
rect 1110 458 1162 496
rect 1110 424 1119 458
rect 1153 424 1162 458
rect 1110 419 1162 424
rect 1110 355 1119 367
rect 1153 355 1162 367
rect 1110 291 1119 303
rect 1153 291 1162 303
rect 1110 227 1119 239
rect 1153 227 1162 239
rect 1110 170 1162 175
rect 1110 163 1119 170
rect 1153 163 1162 170
rect 1110 105 1162 111
rect 1266 1466 1318 1497
rect 1266 1432 1275 1466
rect 1309 1432 1318 1466
rect 1266 1394 1318 1432
rect 1266 1360 1275 1394
rect 1309 1360 1318 1394
rect 1266 1322 1318 1360
rect 1266 1288 1275 1322
rect 1309 1288 1318 1322
rect 1266 1250 1318 1288
rect 1266 1216 1275 1250
rect 1309 1216 1318 1250
rect 1266 1178 1318 1216
rect 1266 1144 1275 1178
rect 1309 1144 1318 1178
rect 1266 1115 1318 1144
rect 1266 1051 1318 1063
rect 1266 987 1318 999
rect 1266 928 1275 935
rect 1309 928 1318 935
rect 1266 923 1318 928
rect 1266 859 1275 871
rect 1309 859 1318 871
rect 1266 795 1275 807
rect 1309 795 1318 807
rect 1266 731 1275 743
rect 1309 731 1318 743
rect 1266 674 1318 679
rect 1266 667 1275 674
rect 1309 667 1318 674
rect 1266 603 1318 615
rect 1266 539 1318 551
rect 1266 458 1318 487
rect 1266 424 1275 458
rect 1309 424 1318 458
rect 1266 386 1318 424
rect 1266 352 1275 386
rect 1309 352 1318 386
rect 1266 314 1318 352
rect 1266 280 1275 314
rect 1309 280 1318 314
rect 1266 242 1318 280
rect 1266 208 1275 242
rect 1309 208 1318 242
rect 1266 170 1318 208
rect 1266 136 1275 170
rect 1309 136 1318 170
rect 1266 105 1318 136
rect 1422 1491 1474 1497
rect 1422 1432 1431 1439
rect 1465 1432 1474 1439
rect 1422 1427 1474 1432
rect 1422 1363 1431 1375
rect 1465 1363 1474 1375
rect 1422 1299 1431 1311
rect 1465 1299 1474 1311
rect 1422 1235 1431 1247
rect 1465 1235 1474 1247
rect 1422 1178 1474 1183
rect 1422 1144 1431 1178
rect 1465 1144 1474 1178
rect 1422 1106 1474 1144
rect 1422 1072 1431 1106
rect 1465 1072 1474 1106
rect 1422 1034 1474 1072
rect 1422 1000 1431 1034
rect 1465 1000 1474 1034
rect 1422 962 1474 1000
rect 1422 928 1431 962
rect 1465 928 1474 962
rect 1422 890 1474 928
rect 1422 856 1431 890
rect 1465 856 1474 890
rect 1422 818 1474 856
rect 1422 784 1431 818
rect 1465 784 1474 818
rect 1422 746 1474 784
rect 1422 712 1431 746
rect 1465 712 1474 746
rect 1422 674 1474 712
rect 1422 640 1431 674
rect 1465 640 1474 674
rect 1422 602 1474 640
rect 1422 568 1431 602
rect 1465 568 1474 602
rect 1422 530 1474 568
rect 1422 496 1431 530
rect 1465 496 1474 530
rect 1422 458 1474 496
rect 1422 424 1431 458
rect 1465 424 1474 458
rect 1422 419 1474 424
rect 1422 355 1431 367
rect 1465 355 1474 367
rect 1422 291 1431 303
rect 1465 291 1474 303
rect 1422 227 1431 239
rect 1465 227 1474 239
rect 1422 170 1474 175
rect 1422 163 1431 170
rect 1465 163 1474 170
rect 1422 105 1474 111
rect 1578 1466 1630 1497
rect 1578 1432 1587 1466
rect 1621 1432 1630 1466
rect 1578 1394 1630 1432
rect 1578 1360 1587 1394
rect 1621 1360 1630 1394
rect 1578 1322 1630 1360
rect 1578 1288 1587 1322
rect 1621 1288 1630 1322
rect 1578 1250 1630 1288
rect 1578 1216 1587 1250
rect 1621 1216 1630 1250
rect 1578 1178 1630 1216
rect 1578 1144 1587 1178
rect 1621 1144 1630 1178
rect 1578 1115 1630 1144
rect 1578 1051 1630 1063
rect 1578 987 1630 999
rect 1578 928 1587 935
rect 1621 928 1630 935
rect 1578 923 1630 928
rect 1578 859 1587 871
rect 1621 859 1630 871
rect 1578 795 1587 807
rect 1621 795 1630 807
rect 1578 731 1587 743
rect 1621 731 1630 743
rect 1578 674 1630 679
rect 1578 667 1587 674
rect 1621 667 1630 674
rect 1578 603 1630 615
rect 1578 539 1630 551
rect 1578 458 1630 487
rect 1578 424 1587 458
rect 1621 424 1630 458
rect 1578 386 1630 424
rect 1578 352 1587 386
rect 1621 352 1630 386
rect 1578 314 1630 352
rect 1578 280 1587 314
rect 1621 280 1630 314
rect 1578 242 1630 280
rect 1578 208 1587 242
rect 1621 208 1630 242
rect 1578 170 1630 208
rect 1578 136 1587 170
rect 1621 136 1630 170
rect 1578 105 1630 136
rect 1734 1491 1786 1497
rect 1734 1432 1743 1439
rect 1777 1432 1786 1439
rect 1734 1427 1786 1432
rect 1734 1363 1743 1375
rect 1777 1363 1786 1375
rect 1734 1299 1743 1311
rect 1777 1299 1786 1311
rect 1734 1235 1743 1247
rect 1777 1235 1786 1247
rect 1734 1178 1786 1183
rect 1734 1144 1743 1178
rect 1777 1144 1786 1178
rect 1734 1106 1786 1144
rect 1734 1072 1743 1106
rect 1777 1072 1786 1106
rect 1734 1034 1786 1072
rect 1734 1000 1743 1034
rect 1777 1000 1786 1034
rect 1734 962 1786 1000
rect 1734 928 1743 962
rect 1777 928 1786 962
rect 1734 890 1786 928
rect 1734 856 1743 890
rect 1777 856 1786 890
rect 1734 818 1786 856
rect 1734 784 1743 818
rect 1777 784 1786 818
rect 1734 746 1786 784
rect 1734 712 1743 746
rect 1777 712 1786 746
rect 1734 674 1786 712
rect 1734 640 1743 674
rect 1777 640 1786 674
rect 1734 602 1786 640
rect 1734 568 1743 602
rect 1777 568 1786 602
rect 1734 530 1786 568
rect 1734 496 1743 530
rect 1777 496 1786 530
rect 1734 458 1786 496
rect 1734 424 1743 458
rect 1777 424 1786 458
rect 1734 419 1786 424
rect 1734 355 1743 367
rect 1777 355 1786 367
rect 1734 291 1743 303
rect 1777 291 1786 303
rect 1734 227 1743 239
rect 1777 227 1786 239
rect 1734 170 1786 175
rect 1734 163 1743 170
rect 1777 163 1786 170
rect 1734 105 1786 111
rect 1866 1466 1924 1497
rect 1866 1432 1878 1466
rect 1912 1432 1924 1466
rect 1866 1394 1924 1432
rect 1866 1360 1878 1394
rect 1912 1360 1924 1394
rect 1866 1322 1924 1360
rect 1866 1288 1878 1322
rect 1912 1288 1924 1322
rect 1866 1250 1924 1288
rect 1866 1216 1878 1250
rect 1912 1216 1924 1250
rect 1866 1178 1924 1216
rect 1866 1144 1878 1178
rect 1912 1144 1924 1178
rect 1866 1106 1924 1144
rect 1866 1072 1878 1106
rect 1912 1072 1924 1106
rect 1866 1034 1924 1072
rect 1866 1000 1878 1034
rect 1912 1000 1924 1034
rect 1866 962 1924 1000
rect 1866 928 1878 962
rect 1912 928 1924 962
rect 1866 890 1924 928
rect 1866 856 1878 890
rect 1912 856 1924 890
rect 1866 818 1924 856
rect 1866 784 1878 818
rect 1912 784 1924 818
rect 1866 746 1924 784
rect 1866 712 1878 746
rect 1912 712 1924 746
rect 1866 674 1924 712
rect 1866 640 1878 674
rect 1912 640 1924 674
rect 1866 602 1924 640
rect 1866 568 1878 602
rect 1912 568 1924 602
rect 1866 530 1924 568
rect 1866 496 1878 530
rect 1912 496 1924 530
rect 1866 458 1924 496
rect 1866 424 1878 458
rect 1912 424 1924 458
rect 1866 386 1924 424
rect 1866 352 1878 386
rect 1912 352 1924 386
rect 1866 314 1924 352
rect 1866 280 1878 314
rect 1912 280 1924 314
rect 1866 242 1924 280
rect 1866 208 1878 242
rect 1912 208 1924 242
rect 1866 170 1924 208
rect 1866 136 1878 170
rect 1912 136 1924 170
rect 1866 105 1924 136
rect 195 54 1765 66
rect 195 20 207 54
rect 241 20 279 54
rect 313 20 351 54
rect 385 20 423 54
rect 457 20 495 54
rect 529 20 567 54
rect 601 20 639 54
rect 673 20 711 54
rect 745 20 783 54
rect 817 20 855 54
rect 889 20 927 54
rect 961 20 999 54
rect 1033 20 1071 54
rect 1105 20 1143 54
rect 1177 20 1215 54
rect 1249 20 1287 54
rect 1321 20 1359 54
rect 1393 20 1431 54
rect 1465 20 1503 54
rect 1537 20 1575 54
rect 1609 20 1647 54
rect 1681 20 1719 54
rect 1753 20 1765 54
rect 195 0 1765 20
<< via1 >>
rect 174 1466 226 1491
rect 174 1439 183 1466
rect 183 1439 217 1466
rect 217 1439 226 1466
rect 174 1394 226 1427
rect 174 1375 183 1394
rect 183 1375 217 1394
rect 217 1375 226 1394
rect 174 1360 183 1363
rect 183 1360 217 1363
rect 217 1360 226 1363
rect 174 1322 226 1360
rect 174 1311 183 1322
rect 183 1311 217 1322
rect 217 1311 226 1322
rect 174 1288 183 1299
rect 183 1288 217 1299
rect 217 1288 226 1299
rect 174 1250 226 1288
rect 174 1247 183 1250
rect 183 1247 217 1250
rect 217 1247 226 1250
rect 174 1216 183 1235
rect 183 1216 217 1235
rect 217 1216 226 1235
rect 174 1183 226 1216
rect 174 386 226 419
rect 174 367 183 386
rect 183 367 217 386
rect 217 367 226 386
rect 174 352 183 355
rect 183 352 217 355
rect 217 352 226 355
rect 174 314 226 352
rect 174 303 183 314
rect 183 303 217 314
rect 217 303 226 314
rect 174 280 183 291
rect 183 280 217 291
rect 217 280 226 291
rect 174 242 226 280
rect 174 239 183 242
rect 183 239 217 242
rect 217 239 226 242
rect 174 208 183 227
rect 183 208 217 227
rect 217 208 226 227
rect 174 175 226 208
rect 174 136 183 163
rect 183 136 217 163
rect 217 136 226 163
rect 174 111 226 136
rect 330 1106 382 1115
rect 330 1072 339 1106
rect 339 1072 373 1106
rect 373 1072 382 1106
rect 330 1063 382 1072
rect 330 1034 382 1051
rect 330 1000 339 1034
rect 339 1000 373 1034
rect 373 1000 382 1034
rect 330 999 382 1000
rect 330 962 382 987
rect 330 935 339 962
rect 339 935 373 962
rect 373 935 382 962
rect 330 890 382 923
rect 330 871 339 890
rect 339 871 373 890
rect 373 871 382 890
rect 330 856 339 859
rect 339 856 373 859
rect 373 856 382 859
rect 330 818 382 856
rect 330 807 339 818
rect 339 807 373 818
rect 373 807 382 818
rect 330 784 339 795
rect 339 784 373 795
rect 373 784 382 795
rect 330 746 382 784
rect 330 743 339 746
rect 339 743 373 746
rect 373 743 382 746
rect 330 712 339 731
rect 339 712 373 731
rect 373 712 382 731
rect 330 679 382 712
rect 330 640 339 667
rect 339 640 373 667
rect 373 640 382 667
rect 330 615 382 640
rect 330 602 382 603
rect 330 568 339 602
rect 339 568 373 602
rect 373 568 382 602
rect 330 551 382 568
rect 330 530 382 539
rect 330 496 339 530
rect 339 496 373 530
rect 373 496 382 530
rect 330 487 382 496
rect 486 1466 538 1491
rect 486 1439 495 1466
rect 495 1439 529 1466
rect 529 1439 538 1466
rect 486 1394 538 1427
rect 486 1375 495 1394
rect 495 1375 529 1394
rect 529 1375 538 1394
rect 486 1360 495 1363
rect 495 1360 529 1363
rect 529 1360 538 1363
rect 486 1322 538 1360
rect 486 1311 495 1322
rect 495 1311 529 1322
rect 529 1311 538 1322
rect 486 1288 495 1299
rect 495 1288 529 1299
rect 529 1288 538 1299
rect 486 1250 538 1288
rect 486 1247 495 1250
rect 495 1247 529 1250
rect 529 1247 538 1250
rect 486 1216 495 1235
rect 495 1216 529 1235
rect 529 1216 538 1235
rect 486 1183 538 1216
rect 486 386 538 419
rect 486 367 495 386
rect 495 367 529 386
rect 529 367 538 386
rect 486 352 495 355
rect 495 352 529 355
rect 529 352 538 355
rect 486 314 538 352
rect 486 303 495 314
rect 495 303 529 314
rect 529 303 538 314
rect 486 280 495 291
rect 495 280 529 291
rect 529 280 538 291
rect 486 242 538 280
rect 486 239 495 242
rect 495 239 529 242
rect 529 239 538 242
rect 486 208 495 227
rect 495 208 529 227
rect 529 208 538 227
rect 486 175 538 208
rect 486 136 495 163
rect 495 136 529 163
rect 529 136 538 163
rect 486 111 538 136
rect 642 1106 694 1115
rect 642 1072 651 1106
rect 651 1072 685 1106
rect 685 1072 694 1106
rect 642 1063 694 1072
rect 642 1034 694 1051
rect 642 1000 651 1034
rect 651 1000 685 1034
rect 685 1000 694 1034
rect 642 999 694 1000
rect 642 962 694 987
rect 642 935 651 962
rect 651 935 685 962
rect 685 935 694 962
rect 642 890 694 923
rect 642 871 651 890
rect 651 871 685 890
rect 685 871 694 890
rect 642 856 651 859
rect 651 856 685 859
rect 685 856 694 859
rect 642 818 694 856
rect 642 807 651 818
rect 651 807 685 818
rect 685 807 694 818
rect 642 784 651 795
rect 651 784 685 795
rect 685 784 694 795
rect 642 746 694 784
rect 642 743 651 746
rect 651 743 685 746
rect 685 743 694 746
rect 642 712 651 731
rect 651 712 685 731
rect 685 712 694 731
rect 642 679 694 712
rect 642 640 651 667
rect 651 640 685 667
rect 685 640 694 667
rect 642 615 694 640
rect 642 602 694 603
rect 642 568 651 602
rect 651 568 685 602
rect 685 568 694 602
rect 642 551 694 568
rect 642 530 694 539
rect 642 496 651 530
rect 651 496 685 530
rect 685 496 694 530
rect 642 487 694 496
rect 798 1466 850 1491
rect 798 1439 807 1466
rect 807 1439 841 1466
rect 841 1439 850 1466
rect 798 1394 850 1427
rect 798 1375 807 1394
rect 807 1375 841 1394
rect 841 1375 850 1394
rect 798 1360 807 1363
rect 807 1360 841 1363
rect 841 1360 850 1363
rect 798 1322 850 1360
rect 798 1311 807 1322
rect 807 1311 841 1322
rect 841 1311 850 1322
rect 798 1288 807 1299
rect 807 1288 841 1299
rect 841 1288 850 1299
rect 798 1250 850 1288
rect 798 1247 807 1250
rect 807 1247 841 1250
rect 841 1247 850 1250
rect 798 1216 807 1235
rect 807 1216 841 1235
rect 841 1216 850 1235
rect 798 1183 850 1216
rect 798 386 850 419
rect 798 367 807 386
rect 807 367 841 386
rect 841 367 850 386
rect 798 352 807 355
rect 807 352 841 355
rect 841 352 850 355
rect 798 314 850 352
rect 798 303 807 314
rect 807 303 841 314
rect 841 303 850 314
rect 798 280 807 291
rect 807 280 841 291
rect 841 280 850 291
rect 798 242 850 280
rect 798 239 807 242
rect 807 239 841 242
rect 841 239 850 242
rect 798 208 807 227
rect 807 208 841 227
rect 841 208 850 227
rect 798 175 850 208
rect 798 136 807 163
rect 807 136 841 163
rect 841 136 850 163
rect 798 111 850 136
rect 954 1106 1006 1115
rect 954 1072 963 1106
rect 963 1072 997 1106
rect 997 1072 1006 1106
rect 954 1063 1006 1072
rect 954 1034 1006 1051
rect 954 1000 963 1034
rect 963 1000 997 1034
rect 997 1000 1006 1034
rect 954 999 1006 1000
rect 954 962 1006 987
rect 954 935 963 962
rect 963 935 997 962
rect 997 935 1006 962
rect 954 890 1006 923
rect 954 871 963 890
rect 963 871 997 890
rect 997 871 1006 890
rect 954 856 963 859
rect 963 856 997 859
rect 997 856 1006 859
rect 954 818 1006 856
rect 954 807 963 818
rect 963 807 997 818
rect 997 807 1006 818
rect 954 784 963 795
rect 963 784 997 795
rect 997 784 1006 795
rect 954 746 1006 784
rect 954 743 963 746
rect 963 743 997 746
rect 997 743 1006 746
rect 954 712 963 731
rect 963 712 997 731
rect 997 712 1006 731
rect 954 679 1006 712
rect 954 640 963 667
rect 963 640 997 667
rect 997 640 1006 667
rect 954 615 1006 640
rect 954 602 1006 603
rect 954 568 963 602
rect 963 568 997 602
rect 997 568 1006 602
rect 954 551 1006 568
rect 954 530 1006 539
rect 954 496 963 530
rect 963 496 997 530
rect 997 496 1006 530
rect 954 487 1006 496
rect 1110 1466 1162 1491
rect 1110 1439 1119 1466
rect 1119 1439 1153 1466
rect 1153 1439 1162 1466
rect 1110 1394 1162 1427
rect 1110 1375 1119 1394
rect 1119 1375 1153 1394
rect 1153 1375 1162 1394
rect 1110 1360 1119 1363
rect 1119 1360 1153 1363
rect 1153 1360 1162 1363
rect 1110 1322 1162 1360
rect 1110 1311 1119 1322
rect 1119 1311 1153 1322
rect 1153 1311 1162 1322
rect 1110 1288 1119 1299
rect 1119 1288 1153 1299
rect 1153 1288 1162 1299
rect 1110 1250 1162 1288
rect 1110 1247 1119 1250
rect 1119 1247 1153 1250
rect 1153 1247 1162 1250
rect 1110 1216 1119 1235
rect 1119 1216 1153 1235
rect 1153 1216 1162 1235
rect 1110 1183 1162 1216
rect 1110 386 1162 419
rect 1110 367 1119 386
rect 1119 367 1153 386
rect 1153 367 1162 386
rect 1110 352 1119 355
rect 1119 352 1153 355
rect 1153 352 1162 355
rect 1110 314 1162 352
rect 1110 303 1119 314
rect 1119 303 1153 314
rect 1153 303 1162 314
rect 1110 280 1119 291
rect 1119 280 1153 291
rect 1153 280 1162 291
rect 1110 242 1162 280
rect 1110 239 1119 242
rect 1119 239 1153 242
rect 1153 239 1162 242
rect 1110 208 1119 227
rect 1119 208 1153 227
rect 1153 208 1162 227
rect 1110 175 1162 208
rect 1110 136 1119 163
rect 1119 136 1153 163
rect 1153 136 1162 163
rect 1110 111 1162 136
rect 1266 1106 1318 1115
rect 1266 1072 1275 1106
rect 1275 1072 1309 1106
rect 1309 1072 1318 1106
rect 1266 1063 1318 1072
rect 1266 1034 1318 1051
rect 1266 1000 1275 1034
rect 1275 1000 1309 1034
rect 1309 1000 1318 1034
rect 1266 999 1318 1000
rect 1266 962 1318 987
rect 1266 935 1275 962
rect 1275 935 1309 962
rect 1309 935 1318 962
rect 1266 890 1318 923
rect 1266 871 1275 890
rect 1275 871 1309 890
rect 1309 871 1318 890
rect 1266 856 1275 859
rect 1275 856 1309 859
rect 1309 856 1318 859
rect 1266 818 1318 856
rect 1266 807 1275 818
rect 1275 807 1309 818
rect 1309 807 1318 818
rect 1266 784 1275 795
rect 1275 784 1309 795
rect 1309 784 1318 795
rect 1266 746 1318 784
rect 1266 743 1275 746
rect 1275 743 1309 746
rect 1309 743 1318 746
rect 1266 712 1275 731
rect 1275 712 1309 731
rect 1309 712 1318 731
rect 1266 679 1318 712
rect 1266 640 1275 667
rect 1275 640 1309 667
rect 1309 640 1318 667
rect 1266 615 1318 640
rect 1266 602 1318 603
rect 1266 568 1275 602
rect 1275 568 1309 602
rect 1309 568 1318 602
rect 1266 551 1318 568
rect 1266 530 1318 539
rect 1266 496 1275 530
rect 1275 496 1309 530
rect 1309 496 1318 530
rect 1266 487 1318 496
rect 1422 1466 1474 1491
rect 1422 1439 1431 1466
rect 1431 1439 1465 1466
rect 1465 1439 1474 1466
rect 1422 1394 1474 1427
rect 1422 1375 1431 1394
rect 1431 1375 1465 1394
rect 1465 1375 1474 1394
rect 1422 1360 1431 1363
rect 1431 1360 1465 1363
rect 1465 1360 1474 1363
rect 1422 1322 1474 1360
rect 1422 1311 1431 1322
rect 1431 1311 1465 1322
rect 1465 1311 1474 1322
rect 1422 1288 1431 1299
rect 1431 1288 1465 1299
rect 1465 1288 1474 1299
rect 1422 1250 1474 1288
rect 1422 1247 1431 1250
rect 1431 1247 1465 1250
rect 1465 1247 1474 1250
rect 1422 1216 1431 1235
rect 1431 1216 1465 1235
rect 1465 1216 1474 1235
rect 1422 1183 1474 1216
rect 1422 386 1474 419
rect 1422 367 1431 386
rect 1431 367 1465 386
rect 1465 367 1474 386
rect 1422 352 1431 355
rect 1431 352 1465 355
rect 1465 352 1474 355
rect 1422 314 1474 352
rect 1422 303 1431 314
rect 1431 303 1465 314
rect 1465 303 1474 314
rect 1422 280 1431 291
rect 1431 280 1465 291
rect 1465 280 1474 291
rect 1422 242 1474 280
rect 1422 239 1431 242
rect 1431 239 1465 242
rect 1465 239 1474 242
rect 1422 208 1431 227
rect 1431 208 1465 227
rect 1465 208 1474 227
rect 1422 175 1474 208
rect 1422 136 1431 163
rect 1431 136 1465 163
rect 1465 136 1474 163
rect 1422 111 1474 136
rect 1578 1106 1630 1115
rect 1578 1072 1587 1106
rect 1587 1072 1621 1106
rect 1621 1072 1630 1106
rect 1578 1063 1630 1072
rect 1578 1034 1630 1051
rect 1578 1000 1587 1034
rect 1587 1000 1621 1034
rect 1621 1000 1630 1034
rect 1578 999 1630 1000
rect 1578 962 1630 987
rect 1578 935 1587 962
rect 1587 935 1621 962
rect 1621 935 1630 962
rect 1578 890 1630 923
rect 1578 871 1587 890
rect 1587 871 1621 890
rect 1621 871 1630 890
rect 1578 856 1587 859
rect 1587 856 1621 859
rect 1621 856 1630 859
rect 1578 818 1630 856
rect 1578 807 1587 818
rect 1587 807 1621 818
rect 1621 807 1630 818
rect 1578 784 1587 795
rect 1587 784 1621 795
rect 1621 784 1630 795
rect 1578 746 1630 784
rect 1578 743 1587 746
rect 1587 743 1621 746
rect 1621 743 1630 746
rect 1578 712 1587 731
rect 1587 712 1621 731
rect 1621 712 1630 731
rect 1578 679 1630 712
rect 1578 640 1587 667
rect 1587 640 1621 667
rect 1621 640 1630 667
rect 1578 615 1630 640
rect 1578 602 1630 603
rect 1578 568 1587 602
rect 1587 568 1621 602
rect 1621 568 1630 602
rect 1578 551 1630 568
rect 1578 530 1630 539
rect 1578 496 1587 530
rect 1587 496 1621 530
rect 1621 496 1630 530
rect 1578 487 1630 496
rect 1734 1466 1786 1491
rect 1734 1439 1743 1466
rect 1743 1439 1777 1466
rect 1777 1439 1786 1466
rect 1734 1394 1786 1427
rect 1734 1375 1743 1394
rect 1743 1375 1777 1394
rect 1777 1375 1786 1394
rect 1734 1360 1743 1363
rect 1743 1360 1777 1363
rect 1777 1360 1786 1363
rect 1734 1322 1786 1360
rect 1734 1311 1743 1322
rect 1743 1311 1777 1322
rect 1777 1311 1786 1322
rect 1734 1288 1743 1299
rect 1743 1288 1777 1299
rect 1777 1288 1786 1299
rect 1734 1250 1786 1288
rect 1734 1247 1743 1250
rect 1743 1247 1777 1250
rect 1777 1247 1786 1250
rect 1734 1216 1743 1235
rect 1743 1216 1777 1235
rect 1777 1216 1786 1235
rect 1734 1183 1786 1216
rect 1734 386 1786 419
rect 1734 367 1743 386
rect 1743 367 1777 386
rect 1777 367 1786 386
rect 1734 352 1743 355
rect 1743 352 1777 355
rect 1777 352 1786 355
rect 1734 314 1786 352
rect 1734 303 1743 314
rect 1743 303 1777 314
rect 1777 303 1786 314
rect 1734 280 1743 291
rect 1743 280 1777 291
rect 1777 280 1786 291
rect 1734 242 1786 280
rect 1734 239 1743 242
rect 1743 239 1777 242
rect 1777 239 1786 242
rect 1734 208 1743 227
rect 1743 208 1777 227
rect 1777 208 1786 227
rect 1734 175 1786 208
rect 1734 136 1743 163
rect 1743 136 1777 163
rect 1777 136 1786 163
rect 1734 111 1786 136
<< metal2 >>
rect 10 1491 1950 1497
rect 10 1439 174 1491
rect 226 1439 486 1491
rect 538 1439 798 1491
rect 850 1439 1110 1491
rect 1162 1439 1422 1491
rect 1474 1439 1734 1491
rect 1786 1439 1950 1491
rect 10 1427 1950 1439
rect 10 1375 174 1427
rect 226 1375 486 1427
rect 538 1375 798 1427
rect 850 1375 1110 1427
rect 1162 1375 1422 1427
rect 1474 1375 1734 1427
rect 1786 1375 1950 1427
rect 10 1363 1950 1375
rect 10 1311 174 1363
rect 226 1311 486 1363
rect 538 1311 798 1363
rect 850 1311 1110 1363
rect 1162 1311 1422 1363
rect 1474 1311 1734 1363
rect 1786 1311 1950 1363
rect 10 1299 1950 1311
rect 10 1247 174 1299
rect 226 1247 486 1299
rect 538 1247 798 1299
rect 850 1247 1110 1299
rect 1162 1247 1422 1299
rect 1474 1247 1734 1299
rect 1786 1247 1950 1299
rect 10 1235 1950 1247
rect 10 1183 174 1235
rect 226 1183 486 1235
rect 538 1183 798 1235
rect 850 1183 1110 1235
rect 1162 1183 1422 1235
rect 1474 1183 1734 1235
rect 1786 1183 1950 1235
rect 10 1177 1950 1183
rect 10 1115 1950 1121
rect 10 1063 330 1115
rect 382 1063 642 1115
rect 694 1063 954 1115
rect 1006 1063 1266 1115
rect 1318 1063 1578 1115
rect 1630 1063 1950 1115
rect 10 1051 1950 1063
rect 10 999 330 1051
rect 382 999 642 1051
rect 694 999 954 1051
rect 1006 999 1266 1051
rect 1318 999 1578 1051
rect 1630 999 1950 1051
rect 10 987 1950 999
rect 10 935 330 987
rect 382 935 642 987
rect 694 935 954 987
rect 1006 935 1266 987
rect 1318 935 1578 987
rect 1630 935 1950 987
rect 10 923 1950 935
rect 10 871 330 923
rect 382 871 642 923
rect 694 871 954 923
rect 1006 871 1266 923
rect 1318 871 1578 923
rect 1630 871 1950 923
rect 10 859 1950 871
rect 10 807 330 859
rect 382 807 642 859
rect 694 807 954 859
rect 1006 807 1266 859
rect 1318 807 1578 859
rect 1630 807 1950 859
rect 10 795 1950 807
rect 10 743 330 795
rect 382 743 642 795
rect 694 743 954 795
rect 1006 743 1266 795
rect 1318 743 1578 795
rect 1630 743 1950 795
rect 10 731 1950 743
rect 10 679 330 731
rect 382 679 642 731
rect 694 679 954 731
rect 1006 679 1266 731
rect 1318 679 1578 731
rect 1630 679 1950 731
rect 10 667 1950 679
rect 10 615 330 667
rect 382 615 642 667
rect 694 615 954 667
rect 1006 615 1266 667
rect 1318 615 1578 667
rect 1630 615 1950 667
rect 10 603 1950 615
rect 10 551 330 603
rect 382 551 642 603
rect 694 551 954 603
rect 1006 551 1266 603
rect 1318 551 1578 603
rect 1630 551 1950 603
rect 10 539 1950 551
rect 10 487 330 539
rect 382 487 642 539
rect 694 487 954 539
rect 1006 487 1266 539
rect 1318 487 1578 539
rect 1630 487 1950 539
rect 10 481 1950 487
rect 10 419 1950 425
rect 10 367 174 419
rect 226 367 486 419
rect 538 367 798 419
rect 850 367 1110 419
rect 1162 367 1422 419
rect 1474 367 1734 419
rect 1786 367 1950 419
rect 10 355 1950 367
rect 10 303 174 355
rect 226 303 486 355
rect 538 303 798 355
rect 850 303 1110 355
rect 1162 303 1422 355
rect 1474 303 1734 355
rect 1786 303 1950 355
rect 10 291 1950 303
rect 10 239 174 291
rect 226 239 486 291
rect 538 239 798 291
rect 850 239 1110 291
rect 1162 239 1422 291
rect 1474 239 1734 291
rect 1786 239 1950 291
rect 10 227 1950 239
rect 10 175 174 227
rect 226 175 486 227
rect 538 175 798 227
rect 850 175 1110 227
rect 1162 175 1422 227
rect 1474 175 1734 227
rect 1786 175 1950 227
rect 10 163 1950 175
rect 10 111 174 163
rect 226 111 486 163
rect 538 111 798 163
rect 850 111 1110 163
rect 1162 111 1422 163
rect 1474 111 1734 163
rect 1786 111 1950 163
rect 10 105 1950 111
<< labels >>
flabel comment s 200 801 200 801 0 FreeSans 300 0 0 0 S
flabel comment s 200 801 200 801 0 FreeSans 300 0 0 0 S
flabel comment s 356 801 356 801 0 FreeSans 300 0 0 0 S
flabel comment s 356 801 356 801 0 FreeSans 300 0 0 0 D
flabel comment s 512 801 512 801 0 FreeSans 300 0 0 0 S
flabel comment s 512 801 512 801 0 FreeSans 300 0 0 0 S
flabel comment s 668 801 668 801 0 FreeSans 300 0 0 0 S
flabel comment s 668 801 668 801 0 FreeSans 300 0 0 0 D
flabel comment s 824 801 824 801 0 FreeSans 300 0 0 0 S
flabel comment s 824 801 824 801 0 FreeSans 300 0 0 0 D
flabel comment s 980 801 980 801 0 FreeSans 300 0 0 0 S
flabel comment s 980 801 980 801 0 FreeSans 300 0 0 0 S
flabel comment s 1136 801 1136 801 0 FreeSans 300 0 0 0 S
flabel comment s 1136 801 1136 801 0 FreeSans 300 0 0 0 D
flabel comment s 1292 801 1292 801 0 FreeSans 300 0 0 0 D
flabel comment s 1292 801 1292 801 0 FreeSans 300 0 0 0 S
flabel comment s 1448 801 1448 801 0 FreeSans 300 0 0 0 S
flabel comment s 1448 801 1448 801 0 FreeSans 300 0 0 0 S
flabel comment s 1604 801 1604 801 0 FreeSans 300 0 0 0 D
flabel comment s 1604 801 1604 801 0 FreeSans 300 0 0 0 S
flabel comment s 1760 801 1760 801 0 FreeSans 300 0 0 0 S
flabel metal2 s 41 701 86 925 0 FreeSans 200 90 0 0 DRAIN
port 2 nsew
flabel metal2 s 41 1265 83 1417 0 FreeSans 200 90 0 0 SOURCE
port 3 nsew
flabel metal2 s 41 176 80 367 0 FreeSans 200 90 0 0 SOURCE
port 3 nsew
flabel metal1 s 1878 1086 1907 1205 0 FreeSans 200 90 0 0 SUBSTRATE
port 4 nsew
flabel metal1 s 909 1548 1064 1587 0 FreeSans 200 0 0 0 GATE
port 5 nsew
flabel metal1 s 906 15 1064 54 0 FreeSans 200 0 0 0 GATE
port 5 nsew
flabel metal1 s 47 1077 80 1205 0 FreeSans 200 90 0 0 SUBSTRATE
port 4 nsew
<< properties >>
string GDS_END 7971292
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 7914840
<< end >>
