magic
tech sky130A
timestamp 1707688321
<< poly >>
rect 0 331 67 339
rect 0 8 8 331
rect 59 8 67 331
rect 0 0 67 8
<< polycont >>
rect 8 8 59 331
<< locali >>
rect 8 331 59 339
rect 8 0 59 8
<< properties >>
string GDS_END 87772416
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87770940
<< end >>
