magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -38 261 1418 582
<< pwell >>
rect 1 21 1339 203
rect 29 -17 63 21
<< locali >>
rect 29 215 130 323
rect 96 199 130 215
rect 312 341 545 407
rect 312 317 572 341
rect 514 179 572 317
rect 606 296 1290 341
rect 606 213 675 296
rect 709 213 994 262
rect 1041 215 1290 296
rect 514 173 977 179
rect 255 139 977 173
rect 255 123 465 139
rect 651 135 977 139
rect 255 74 293 123
rect 427 51 465 123
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 25 401 91 493
rect 125 435 177 527
rect 232 443 619 493
rect 653 455 719 527
rect 825 455 891 527
rect 25 357 198 401
rect 232 359 271 443
rect 387 441 619 443
rect 579 421 619 441
rect 925 421 963 493
rect 997 455 1063 527
rect 1097 421 1133 493
rect 1169 455 1235 527
rect 1269 421 1321 493
rect 164 269 198 357
rect 579 375 1321 421
rect 164 207 480 269
rect 164 159 221 207
rect 18 123 221 159
rect 1011 147 1235 181
rect 18 51 89 123
rect 144 17 221 89
rect 327 17 393 89
rect 499 17 617 105
rect 1011 101 1063 147
rect 653 51 1063 101
rect 1097 17 1135 113
rect 1169 51 1235 147
rect 1269 17 1321 177
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
<< metal1 >>
rect 0 561 1380 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 0 496 1380 527
rect 0 17 1380 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
rect 0 -48 1380 -17
<< labels >>
rlabel locali s 709 213 994 262 6 A1
port 1 nsew signal input
rlabel locali s 1041 215 1290 296 6 A2
port 2 nsew signal input
rlabel locali s 606 213 675 296 6 A2
port 2 nsew signal input
rlabel locali s 606 296 1290 341 6 A2
port 2 nsew signal input
rlabel locali s 96 199 130 215 6 B1_N
port 3 nsew signal input
rlabel locali s 29 215 130 323 6 B1_N
port 3 nsew signal input
rlabel metal1 s 0 -48 1380 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 1339 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 1418 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 1380 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 427 51 465 123 6 Y
port 8 nsew signal output
rlabel locali s 255 74 293 123 6 Y
port 8 nsew signal output
rlabel locali s 651 135 977 139 6 Y
port 8 nsew signal output
rlabel locali s 255 123 465 139 6 Y
port 8 nsew signal output
rlabel locali s 255 139 977 173 6 Y
port 8 nsew signal output
rlabel locali s 514 173 977 179 6 Y
port 8 nsew signal output
rlabel locali s 514 179 572 317 6 Y
port 8 nsew signal output
rlabel locali s 312 317 572 341 6 Y
port 8 nsew signal output
rlabel locali s 312 341 545 407 6 Y
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1380 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 4010510
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 4001078
<< end >>
