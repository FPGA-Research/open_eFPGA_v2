magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -89 -36 125 236
<< pmoshvt >>
rect 0 0 36 200
<< pdiff >>
rect -50 0 0 200
rect 36 0 86 200
<< poly >>
rect 0 200 36 226
rect 0 -26 36 0
<< metal1 >>
rect -51 -16 -5 186
rect 41 -16 87 186
use hvDFM1sd_CDNS_52468879185130  hvDFM1sd_CDNS_52468879185130_0
timestamp 1707688321
transform -1 0 0 0 1 0
box -36 -36 89 236
use hvDFM1sd_CDNS_52468879185130  hvDFM1sd_CDNS_52468879185130_1
timestamp 1707688321
transform 1 0 36 0 1 0
box -36 -36 89 236
<< labels >>
flabel comment s -28 85 -28 85 0 FreeSans 300 0 0 0 S
flabel comment s 64 85 64 85 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 86829724
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86828770
<< end >>
