magic
tech sky130A
timestamp 1707688321
<< metal1 >>
rect 0 0 3 186
rect 61 0 64 186
<< via1 >>
rect 3 0 61 186
<< metal2 >>
rect 0 0 3 186
rect 61 0 64 186
<< properties >>
string GDS_END 79997126
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 79996226
<< end >>
