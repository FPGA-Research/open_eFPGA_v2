magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< locali >>
rect 248 961 382 980
rect 248 855 262 961
rect 368 855 382 961
rect 248 841 382 855
rect 248 125 382 139
rect 248 19 262 125
rect 368 19 382 125
rect 248 0 382 19
<< viali >>
rect 262 855 368 961
rect 262 19 368 125
<< obsli1 >>
rect 120 817 186 883
rect 444 817 510 883
rect 120 795 160 817
rect 470 795 510 817
rect 41 759 160 795
rect 41 725 60 759
rect 94 725 160 759
rect 41 687 160 725
rect 41 653 60 687
rect 94 653 160 687
rect 41 615 160 653
rect 41 581 60 615
rect 94 581 160 615
rect 41 543 160 581
rect 41 509 60 543
rect 94 509 160 543
rect 41 471 160 509
rect 41 437 60 471
rect 94 437 160 471
rect 41 399 160 437
rect 41 365 60 399
rect 94 365 160 399
rect 41 327 160 365
rect 41 293 60 327
rect 94 293 160 327
rect 41 255 160 293
rect 41 221 60 255
rect 94 221 160 255
rect 41 185 160 221
rect 212 185 246 795
rect 298 185 332 795
rect 384 185 418 795
rect 470 759 589 795
rect 470 725 536 759
rect 570 725 589 759
rect 470 687 589 725
rect 470 653 536 687
rect 570 653 589 687
rect 470 615 589 653
rect 470 581 536 615
rect 570 581 589 615
rect 470 543 589 581
rect 470 509 536 543
rect 570 509 589 543
rect 470 471 589 509
rect 470 437 536 471
rect 570 437 589 471
rect 470 399 589 437
rect 470 365 536 399
rect 570 365 589 399
rect 470 327 589 365
rect 470 293 536 327
rect 570 293 589 327
rect 470 255 589 293
rect 470 221 536 255
rect 570 221 589 255
rect 470 185 589 221
rect 120 163 160 185
rect 470 163 510 185
rect 120 97 186 163
rect 444 97 510 163
<< obsli1c >>
rect 60 725 94 759
rect 60 653 94 687
rect 60 581 94 615
rect 60 509 94 543
rect 60 437 94 471
rect 60 365 94 399
rect 60 293 94 327
rect 60 221 94 255
rect 536 725 570 759
rect 536 653 570 687
rect 536 581 570 615
rect 536 509 570 543
rect 536 437 570 471
rect 536 365 570 399
rect 536 293 570 327
rect 536 221 570 255
<< metal1 >>
rect 250 961 380 980
rect 250 855 262 961
rect 368 855 380 961
rect 250 843 380 855
rect 41 759 100 771
rect 41 725 60 759
rect 94 725 100 759
rect 41 687 100 725
rect 41 653 60 687
rect 94 653 100 687
rect 41 615 100 653
rect 41 581 60 615
rect 94 581 100 615
rect 41 543 100 581
rect 41 509 60 543
rect 94 509 100 543
rect 41 471 100 509
rect 41 437 60 471
rect 94 437 100 471
rect 41 399 100 437
rect 41 365 60 399
rect 94 365 100 399
rect 41 327 100 365
rect 41 293 60 327
rect 94 293 100 327
rect 41 255 100 293
rect 41 221 60 255
rect 94 221 100 255
rect 41 209 100 221
rect 530 759 589 771
rect 530 725 536 759
rect 570 725 589 759
rect 530 687 589 725
rect 530 653 536 687
rect 570 653 589 687
rect 530 615 589 653
rect 530 581 536 615
rect 570 581 589 615
rect 530 543 589 581
rect 530 509 536 543
rect 570 509 589 543
rect 530 471 589 509
rect 530 437 536 471
rect 570 437 589 471
rect 530 399 589 437
rect 530 365 536 399
rect 570 365 589 399
rect 530 327 589 365
rect 530 293 536 327
rect 570 293 589 327
rect 530 255 589 293
rect 530 221 536 255
rect 570 221 589 255
rect 530 209 589 221
rect 250 125 380 137
rect 250 19 262 125
rect 368 19 380 125
rect 250 0 380 19
<< obsm1 >>
rect 203 209 255 771
rect 289 209 341 771
rect 375 209 427 771
<< metal2 >>
rect 14 515 616 771
rect 14 209 616 465
<< labels >>
rlabel metal2 s 14 515 616 771 6 DRAIN
port 1 nsew
rlabel viali s 262 855 368 961 6 GATE
port 2 nsew
rlabel viali s 262 19 368 125 6 GATE
port 2 nsew
rlabel locali s 248 841 382 980 6 GATE
port 2 nsew
rlabel locali s 248 0 382 139 6 GATE
port 2 nsew
rlabel metal1 s 250 843 380 980 6 GATE
port 2 nsew
rlabel metal1 s 250 0 380 137 6 GATE
port 2 nsew
rlabel metal2 s 14 209 616 465 6 SOURCE
port 3 nsew
rlabel metal1 s 41 209 100 771 6 SUBSTRATE
port 4 nsew
rlabel metal1 s 530 209 589 771 6 SUBSTRATE
port 4 nsew
<< properties >>
string FIXED_BBOX 14 0 616 980
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6545994
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 6533130
<< end >>
