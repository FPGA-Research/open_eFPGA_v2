magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< pwell >>
rect 78 373 88 389
<< obsli1 >>
rect 83 447 217 463
rect 83 413 97 447
rect 131 413 169 447
rect 203 413 217 447
rect 83 397 217 413
rect 47 329 81 357
rect 47 257 81 295
rect 47 185 81 223
rect 47 113 81 151
rect 47 51 81 79
rect 133 51 167 357
rect 219 329 253 357
rect 219 257 253 295
rect 219 185 253 223
rect 219 113 253 151
rect 219 51 253 79
<< obsli1c >>
rect 97 413 131 447
rect 169 413 203 447
rect 47 295 81 329
rect 47 223 81 257
rect 47 151 81 185
rect 47 79 81 113
rect 219 295 253 329
rect 219 223 253 257
rect 219 151 253 185
rect 219 79 253 113
<< metal1 >>
rect 85 447 215 459
rect 85 413 97 447
rect 131 413 169 447
rect 203 413 215 447
rect 85 401 215 413
rect 41 329 87 357
rect 41 295 47 329
rect 81 295 87 329
rect 41 257 87 295
rect 41 223 47 257
rect 81 223 87 257
rect 41 185 87 223
rect 41 151 47 185
rect 81 151 87 185
rect 41 113 87 151
rect 41 79 47 113
rect 81 79 87 113
rect 41 -29 87 79
rect 213 329 259 357
rect 213 295 219 329
rect 253 295 259 329
rect 213 257 259 295
rect 213 223 219 257
rect 253 223 259 257
rect 213 185 259 223
rect 213 151 219 185
rect 253 151 259 185
rect 213 113 259 151
rect 213 79 219 113
rect 253 79 259 113
rect 213 -29 259 79
rect 41 -89 259 -29
<< obsm1 >>
rect 124 51 176 357
<< metal2 >>
rect 124 224 176 352
<< labels >>
rlabel metal2 s 124 224 176 352 6 DRAIN
port 1 nsew
rlabel metal1 s 85 401 215 459 6 GATE
port 2 nsew
rlabel metal1 s 213 -29 259 357 6 SOURCE
port 3 nsew
rlabel metal1 s 41 -29 87 357 6 SOURCE
port 3 nsew
rlabel metal1 s 41 -89 259 -29 8 SOURCE
port 3 nsew
rlabel pwell s 78 373 88 389 6 SUBSTRATE
port 4 nsew
<< properties >>
string FIXED_BBOX 36 -89 264 463
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 5769084
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 5764462
<< end >>
