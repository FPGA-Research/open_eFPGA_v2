magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 156 163 815 203
rect 1 27 815 163
rect 29 21 815 27
rect 29 -17 63 21
<< scnmos >>
rect 79 53 109 137
rect 259 47 289 177
rect 343 47 373 177
rect 441 47 471 177
rect 525 47 555 177
rect 609 47 639 177
rect 693 47 723 177
<< scpmoshvt >>
rect 79 413 109 497
rect 271 297 301 497
rect 343 297 373 497
rect 441 297 471 497
rect 525 297 555 497
rect 609 297 639 497
rect 693 297 723 497
<< ndiff >>
rect 182 137 259 177
rect 27 106 79 137
rect 27 72 35 106
rect 69 72 79 106
rect 27 53 79 72
rect 109 97 259 137
rect 109 63 119 97
rect 153 63 215 97
rect 249 63 259 97
rect 109 53 259 63
rect 182 47 259 53
rect 289 165 343 177
rect 289 131 299 165
rect 333 131 343 165
rect 289 97 343 131
rect 289 63 299 97
rect 333 63 343 97
rect 289 47 343 63
rect 373 165 441 177
rect 373 131 397 165
rect 431 131 441 165
rect 373 97 441 131
rect 373 63 397 97
rect 431 63 441 97
rect 373 47 441 63
rect 471 165 525 177
rect 471 131 481 165
rect 515 131 525 165
rect 471 97 525 131
rect 471 63 481 97
rect 515 63 525 97
rect 471 47 525 63
rect 555 94 609 177
rect 555 60 565 94
rect 599 60 609 94
rect 555 47 609 60
rect 639 165 693 177
rect 639 131 649 165
rect 683 131 693 165
rect 639 97 693 131
rect 639 63 649 97
rect 683 63 693 97
rect 639 47 693 63
rect 723 94 789 177
rect 723 60 733 94
rect 767 60 789 94
rect 723 47 789 60
<< pdiff >>
rect 27 475 79 497
rect 27 441 35 475
rect 69 441 79 475
rect 27 413 79 441
rect 109 457 165 497
rect 109 423 119 457
rect 153 423 165 457
rect 109 413 165 423
rect 219 479 271 497
rect 219 445 227 479
rect 261 445 271 479
rect 219 411 271 445
rect 219 377 227 411
rect 261 377 271 411
rect 219 343 271 377
rect 219 309 227 343
rect 261 309 271 343
rect 219 297 271 309
rect 301 297 343 497
rect 373 485 441 497
rect 373 451 396 485
rect 430 451 441 485
rect 373 417 441 451
rect 373 383 396 417
rect 430 383 441 417
rect 373 297 441 383
rect 471 477 525 497
rect 471 443 481 477
rect 515 443 525 477
rect 471 409 525 443
rect 471 375 481 409
rect 515 375 525 409
rect 471 297 525 375
rect 555 477 609 497
rect 555 443 565 477
rect 599 443 609 477
rect 555 297 609 443
rect 639 477 693 497
rect 639 443 649 477
rect 683 443 693 477
rect 639 409 693 443
rect 639 375 649 409
rect 683 375 693 409
rect 639 341 693 375
rect 639 307 649 341
rect 683 307 693 341
rect 639 297 693 307
rect 723 477 782 497
rect 723 443 733 477
rect 767 443 782 477
rect 723 409 782 443
rect 723 375 733 409
rect 767 375 782 409
rect 723 297 782 375
<< ndiffc >>
rect 35 72 69 106
rect 119 63 153 97
rect 215 63 249 97
rect 299 131 333 165
rect 299 63 333 97
rect 397 131 431 165
rect 397 63 431 97
rect 481 131 515 165
rect 481 63 515 97
rect 565 60 599 94
rect 649 131 683 165
rect 649 63 683 97
rect 733 60 767 94
<< pdiffc >>
rect 35 441 69 475
rect 119 423 153 457
rect 227 445 261 479
rect 227 377 261 411
rect 227 309 261 343
rect 396 451 430 485
rect 396 383 430 417
rect 481 443 515 477
rect 481 375 515 409
rect 565 443 599 477
rect 649 443 683 477
rect 649 375 683 409
rect 649 307 683 341
rect 733 443 767 477
rect 733 375 767 409
<< poly >>
rect 79 497 109 523
rect 271 497 301 523
rect 343 497 373 523
rect 441 497 471 523
rect 525 497 555 523
rect 609 497 639 523
rect 693 497 723 523
rect 79 265 109 413
rect 271 265 301 297
rect 22 249 109 265
rect 22 215 35 249
rect 69 215 109 249
rect 22 199 109 215
rect 174 249 301 265
rect 174 215 184 249
rect 218 215 301 249
rect 174 199 301 215
rect 343 265 373 297
rect 441 265 471 297
rect 525 265 555 297
rect 609 265 639 297
rect 693 265 723 297
rect 343 249 397 265
rect 343 215 353 249
rect 387 215 397 249
rect 343 199 397 215
rect 441 249 723 265
rect 441 215 514 249
rect 548 215 582 249
rect 616 215 650 249
rect 684 215 723 249
rect 441 199 723 215
rect 79 137 109 199
rect 259 177 289 199
rect 343 177 373 199
rect 441 177 471 199
rect 525 177 555 199
rect 609 177 639 199
rect 693 177 723 199
rect 79 27 109 53
rect 259 21 289 47
rect 343 21 373 47
rect 441 21 471 47
rect 525 21 555 47
rect 609 21 639 47
rect 693 21 723 47
<< polycont >>
rect 35 215 69 249
rect 184 215 218 249
rect 353 215 387 249
rect 514 215 548 249
rect 582 215 616 249
rect 650 215 684 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 18 475 69 527
rect 18 441 35 475
rect 18 425 69 441
rect 119 457 153 493
rect 18 249 85 391
rect 18 215 35 249
rect 69 215 85 249
rect 119 265 153 423
rect 198 479 292 493
rect 198 445 227 479
rect 261 445 292 479
rect 198 411 292 445
rect 198 377 227 411
rect 261 377 292 411
rect 198 343 292 377
rect 383 485 439 527
rect 383 451 396 485
rect 430 451 439 485
rect 383 417 439 451
rect 383 383 396 417
rect 430 383 439 417
rect 383 367 439 383
rect 473 477 523 493
rect 473 443 481 477
rect 515 443 523 477
rect 473 409 523 443
rect 557 477 607 527
rect 557 443 565 477
rect 599 443 607 477
rect 557 427 607 443
rect 641 477 691 493
rect 641 443 649 477
rect 683 443 691 477
rect 473 375 481 409
rect 515 391 523 409
rect 641 409 691 443
rect 641 391 649 409
rect 515 375 649 391
rect 683 375 691 409
rect 473 357 691 375
rect 725 477 775 527
rect 725 443 733 477
rect 767 443 775 477
rect 725 409 775 443
rect 725 375 733 409
rect 767 375 775 409
rect 725 359 775 375
rect 198 309 227 343
rect 261 323 292 343
rect 566 341 691 357
rect 261 309 532 323
rect 198 299 532 309
rect 258 289 532 299
rect 566 307 649 341
rect 683 323 691 341
rect 683 307 811 323
rect 566 289 811 307
rect 119 249 224 265
rect 119 215 184 249
rect 218 215 224 249
rect 119 199 224 215
rect 119 181 169 199
rect 22 147 169 181
rect 258 181 292 289
rect 326 249 464 255
rect 326 215 353 249
rect 387 215 464 249
rect 498 249 532 289
rect 498 215 514 249
rect 548 215 582 249
rect 616 215 650 249
rect 684 215 700 249
rect 734 181 811 289
rect 258 165 349 181
rect 258 147 299 165
rect 22 106 84 147
rect 283 131 299 147
rect 333 131 349 165
rect 22 72 35 106
rect 69 72 84 106
rect 22 53 84 72
rect 118 97 249 113
rect 118 63 119 97
rect 153 63 215 97
rect 118 17 249 63
rect 283 97 349 131
rect 283 63 299 97
rect 333 63 349 97
rect 283 61 349 63
rect 396 165 431 181
rect 396 131 397 165
rect 396 97 431 131
rect 396 63 397 97
rect 396 17 431 63
rect 465 165 811 181
rect 465 131 481 165
rect 515 147 649 165
rect 515 131 531 147
rect 465 97 531 131
rect 633 131 649 147
rect 683 147 811 165
rect 683 131 699 147
rect 465 63 481 97
rect 515 63 531 97
rect 465 58 531 63
rect 565 94 599 110
rect 565 17 599 60
rect 633 97 699 131
rect 633 63 649 97
rect 683 63 699 97
rect 633 58 699 63
rect 733 94 767 110
rect 733 17 767 60
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel locali s 397 221 431 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 29 221 63 255 0 FreeSans 400 0 0 0 B_N
port 2 nsew signal input
flabel locali s 765 289 799 323 0 FreeSans 400 0 0 0 X
port 7 nsew signal output
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 or2b_4
rlabel metal1 s 0 -48 828 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 828 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_END 1011720
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1004944
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 4.140 0.000 
<< end >>
