magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -76 -26 1676 626
<< mvnmos >>
rect 0 0 1600 600
<< mvndiff >>
rect -50 0 0 600
rect 1600 0 1650 600
<< poly >>
rect 0 600 1600 632
rect 0 -32 1600 0
<< metal1 >>
rect -51 -16 -5 546
rect 1605 -16 1651 546
use hvDFM1sd2_CDNS_52468879185154  hvDFM1sd2_CDNS_52468879185154_0
timestamp 1707688321
transform -1 0 0 0 1 0
box -26 -26 82 626
use hvDFM1sd2_CDNS_52468879185154  hvDFM1sd2_CDNS_52468879185154_1
timestamp 1707688321
transform 1 0 1600 0 1 0
box -26 -26 82 626
<< labels >>
flabel comment s -28 265 -28 265 0 FreeSans 300 0 0 0 S
flabel comment s 1628 265 1628 265 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 6115406
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 6114512
<< end >>
