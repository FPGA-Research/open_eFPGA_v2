magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 1 21 557 203
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 177
rect 155 47 185 177
rect 279 47 309 177
rect 353 47 383 177
rect 449 47 479 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 279 297 309 497
rect 363 297 393 497
rect 449 297 479 497
<< ndiff >>
rect 27 93 79 177
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 47 155 177
rect 185 123 279 177
rect 185 89 199 123
rect 233 89 279 123
rect 185 47 279 89
rect 309 47 353 177
rect 383 47 449 177
rect 479 161 531 177
rect 479 127 489 161
rect 523 127 531 161
rect 479 93 531 127
rect 479 59 489 93
rect 523 59 531 93
rect 479 47 531 59
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 297 79 383
rect 109 417 163 497
rect 109 383 119 417
rect 153 383 163 417
rect 109 297 163 383
rect 193 477 279 497
rect 193 443 235 477
rect 269 443 279 477
rect 193 391 279 443
rect 193 357 235 391
rect 269 357 279 391
rect 193 297 279 357
rect 309 477 363 497
rect 309 443 319 477
rect 353 443 363 477
rect 309 297 363 443
rect 393 477 449 497
rect 393 443 403 477
rect 437 443 449 477
rect 393 399 449 443
rect 393 365 403 399
rect 437 365 449 399
rect 393 297 449 365
rect 479 485 531 497
rect 479 451 489 485
rect 523 451 531 485
rect 479 417 531 451
rect 479 383 489 417
rect 523 383 531 417
rect 479 349 531 383
rect 479 315 489 349
rect 523 315 531 349
rect 479 297 531 315
<< ndiffc >>
rect 35 59 69 93
rect 199 89 233 123
rect 489 127 523 161
rect 489 59 523 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 119 383 153 417
rect 235 443 269 477
rect 235 357 269 391
rect 319 443 353 477
rect 403 443 437 477
rect 403 365 437 399
rect 489 451 523 485
rect 489 383 523 417
rect 489 315 523 349
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 279 497 309 523
rect 363 497 393 523
rect 449 497 479 523
rect 79 265 109 297
rect 163 265 193 297
rect 279 265 309 297
rect 363 282 393 297
rect 449 282 479 297
rect 21 249 109 265
rect 21 215 31 249
rect 65 215 109 249
rect 21 199 109 215
rect 151 249 215 265
rect 151 215 171 249
rect 205 215 215 249
rect 151 199 215 215
rect 257 249 311 265
rect 257 215 267 249
rect 301 215 311 249
rect 257 199 311 215
rect 353 249 407 282
rect 353 215 363 249
rect 397 215 407 249
rect 79 177 109 199
rect 155 177 185 199
rect 279 177 309 199
rect 353 192 407 215
rect 449 249 537 282
rect 449 215 485 249
rect 519 215 537 249
rect 449 192 537 215
rect 353 177 383 192
rect 449 177 479 192
rect 79 21 109 47
rect 155 21 185 47
rect 279 21 309 47
rect 353 21 383 47
rect 449 21 479 47
<< polycont >>
rect 31 215 65 249
rect 171 215 205 249
rect 267 215 301 249
rect 363 215 397 249
rect 485 215 519 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 17 485 269 493
rect 17 451 35 485
rect 69 477 269 485
rect 69 451 235 477
rect 17 417 69 451
rect 219 443 235 451
rect 17 383 35 417
rect 17 367 69 383
rect 103 383 119 417
rect 153 383 173 417
rect 103 357 173 383
rect 219 391 269 443
rect 311 477 361 527
rect 311 443 319 477
rect 353 443 361 477
rect 311 427 361 443
rect 403 477 437 493
rect 403 399 437 443
rect 219 357 235 391
rect 269 365 403 391
rect 269 357 437 365
rect 17 249 69 265
rect 17 215 31 249
rect 65 215 69 249
rect 17 199 69 215
rect 103 161 137 357
rect 403 349 437 357
rect 471 485 539 527
rect 471 451 489 485
rect 523 451 539 485
rect 471 417 539 451
rect 471 383 489 417
rect 523 383 539 417
rect 471 349 539 383
rect 171 285 251 323
rect 471 315 489 349
rect 523 315 539 349
rect 471 299 539 315
rect 171 249 205 285
rect 246 249 319 251
rect 246 215 267 249
rect 301 215 319 249
rect 171 199 205 215
rect 103 127 233 161
rect 183 123 233 127
rect 19 59 35 93
rect 69 59 85 93
rect 183 89 199 123
rect 183 59 233 89
rect 281 153 319 215
rect 361 249 433 265
rect 361 215 363 249
rect 397 215 433 249
rect 361 199 433 215
rect 467 249 550 265
rect 467 215 485 249
rect 519 215 550 249
rect 467 203 550 215
rect 281 69 341 153
rect 393 83 433 199
rect 471 127 489 161
rect 523 127 539 161
rect 471 93 539 127
rect 471 59 489 93
rect 523 59 539 93
rect 19 17 85 59
rect 471 17 539 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel locali s 399 85 433 119 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 119 357 153 391 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 307 85 341 119 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 B2
port 5 nsew signal input
flabel locali s 215 289 249 323 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 399 153 433 187 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 399 221 433 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 493 221 527 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 a32oi_1
rlabel metal1 s 0 -48 644 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_END 3473666
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3467700
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 16.100 0.000 
<< end >>
