magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< obsli1 >>
rect 366 40 10828 39895
<< metal1 >>
rect 1296 11892 1324 11920
rect 1296 11858 1358 11892
rect 1296 1252 1324 11858
rect 1579 13795 1707 13847
rect 1579 13761 1641 13795
rect 1579 11892 1607 13761
rect 1576 11440 1604 11468
rect 1576 11406 1638 11440
rect 1576 2137 1604 11406
rect 1859 12835 1987 12887
rect 1859 12801 1921 12835
rect 1859 11440 1887 12801
rect 1576 2085 1704 2137
rect 1618 2051 1704 2085
rect 1296 1200 1467 1252
rect 1381 1166 1467 1200
rect 282 0 334 128
rect 1415 0 1467 1166
rect 1652 0 1704 2051
rect 1733 1814 1785 11043
rect 1813 1996 1865 10236
rect 2087 2165 2215 2217
rect 2129 2131 2215 2165
rect 1909 1814 1961 1866
rect 1875 1780 1961 1814
rect 1909 0 1961 1780
rect 2163 0 2215 2131
rect 2483 0 2561 128
rect 6843 0 6895 128
rect 8176 792 8228 844
rect 8176 758 8262 792
rect 8176 0 8228 758
rect 8388 792 8440 948
rect 8469 0 8521 128
rect 8701 0 8753 128
rect 8918 0 8970 128
rect 9232 300 9284 352
rect 9232 266 9318 300
rect 9232 0 9284 266
rect 9492 300 9544 952
rect 9652 291 9704 12268
rect 9784 291 9836 343
rect 9750 257 9836 291
rect 9572 0 9624 128
rect 9784 0 9836 257
rect 10031 0 10083 128
rect 10263 0 10315 128
<< obsm1 >>
rect 282 13903 10828 39895
rect 282 11976 1523 13903
rect 282 1144 1240 11976
rect 1380 11948 1523 11976
rect 1414 11836 1523 11948
rect 1763 13739 10828 13903
rect 1697 13705 10828 13739
rect 1663 12943 10828 13705
rect 1663 11836 1803 12943
rect 1414 11802 1803 11836
rect 1380 11524 1803 11802
rect 1380 2029 1520 11524
rect 1660 11496 1803 11524
rect 1694 11384 1803 11496
rect 2043 12779 10828 12943
rect 1977 12745 10828 12779
rect 1943 12324 10828 12745
rect 1943 11384 9596 12324
rect 1694 11350 9596 11384
rect 1660 11099 9596 11350
rect 1660 2193 1677 11099
rect 1380 1995 1562 2029
rect 1380 1308 1596 1995
rect 282 1110 1325 1144
rect 282 184 1359 1110
rect 282 128 334 184
rect 390 0 1359 184
rect 1523 0 1596 1308
rect 1841 10292 9596 11099
rect 1921 2273 9596 10292
rect 1921 2109 2031 2273
rect 1921 2075 2073 2109
rect 1921 1940 2107 2075
rect 1841 1922 2107 1940
rect 1841 1870 1853 1922
rect 1760 1724 1819 1758
rect 1760 0 1853 1724
rect 2017 0 2107 1922
rect 2271 1008 9596 2273
rect 2271 1004 9436 1008
rect 2271 900 8332 1004
rect 2271 184 8120 900
rect 8284 848 8332 900
rect 2271 0 2427 184
rect 2617 0 6787 184
rect 6951 0 8120 184
rect 8318 736 8332 848
rect 8496 736 9436 1004
rect 8318 702 9436 736
rect 8284 408 9436 702
rect 8284 184 9176 408
rect 9340 356 9436 408
rect 8284 0 8413 184
rect 8577 0 8645 184
rect 8809 0 8862 184
rect 9026 0 9176 184
rect 9374 244 9436 356
rect 9760 399 10828 12324
rect 9374 235 9596 244
rect 9374 210 9694 235
rect 9340 201 9694 210
rect 9340 184 9728 201
rect 9340 0 9516 184
rect 9680 0 9728 184
rect 9892 184 10828 399
rect 9892 0 9975 184
rect 10139 0 10207 184
rect 10371 0 10828 184
<< metal2 >>
rect 282 0 334 128
rect 1415 0 1467 128
rect 1652 0 1704 128
rect 1909 0 1961 128
rect 2163 0 2215 128
rect 2483 0 2561 128
rect 6843 0 6895 128
rect 8176 0 8228 128
rect 8469 0 8521 128
rect 8701 0 8753 128
rect 8918 0 8970 128
rect 9232 0 9284 128
rect 9572 0 9624 128
rect 9784 0 9836 128
rect 10031 0 10083 128
rect 10263 0 10315 128
<< obsm2 >>
rect 282 184 10828 39725
rect 390 0 1359 184
rect 1523 0 1596 184
rect 1760 0 1853 184
rect 2017 0 2107 184
rect 2271 0 2427 184
rect 2617 0 6787 184
rect 6951 0 8120 184
rect 8284 0 8413 184
rect 8577 0 8645 184
rect 8809 0 8862 184
rect 9026 0 9176 184
rect 9340 0 9516 184
rect 9680 0 9728 184
rect 9892 0 9975 184
rect 10139 0 10207 184
rect 10371 0 10828 184
<< metal3 >>
rect 1583 27485 2501 40000
rect 2661 38979 3543 40000
rect 3703 28185 4503 40000
rect 4663 39267 5663 40000
rect 282 0 1423 631
rect 1583 0 2383 25153
rect 5823 22133 6623 40000
rect 6733 27282 7908 40000
rect 2661 0 3543 6774
rect 3703 0 4503 1208
rect 4663 0 5663 7287
rect 5823 0 6725 994
rect 7000 0 7918 1655
<< obsm3 >>
rect 282 27405 1503 40000
rect 2581 28105 3623 38899
rect 4583 28105 5743 39187
rect 2581 27405 5743 28105
rect 282 25233 5743 27405
rect 282 711 1503 25233
rect 2463 22053 5743 25233
rect 7988 27202 10856 40000
rect 6703 22053 10856 27202
rect 2463 7367 10856 22053
rect 2463 6854 4583 7367
rect 2463 0 2581 6854
rect 3623 1288 4583 6854
rect 5743 1735 10856 7367
rect 5743 1074 6920 1735
rect 6805 0 6920 1074
rect 7998 0 10856 1735
<< labels >>
rlabel metal1 s 9232 0 9284 128 6 in1_vddd_hv
port 1 nsew signal input
rlabel metal2 s 9232 0 9284 128 6 in1_vddd_hv
port 1 nsew signal input
rlabel metal1 s 9492 386 9544 952 6 in1_vddd_hv
port 1 nsew signal input
rlabel metal1 s 9492 300 9544 386 6 in1_vddd_hv
port 1 nsew signal input
rlabel metal1 s 9284 266 9318 300 6 in1_vddd_hv
port 1 nsew signal input
rlabel metal1 s 9232 128 9284 352 6 in1_vddd_hv
port 1 nsew signal input
rlabel metal1 s 9572 0 9624 128 6 in2_vddd_hv
port 2 nsew signal input
rlabel metal2 s 9572 0 9624 128 6 in2_vddd_hv
port 2 nsew signal input
rlabel metal1 s 6843 0 6895 128 6 out3_vddio_hv
port 3 nsew signal output
rlabel metal2 s 6843 0 6895 128 6 out3_vddio_hv
port 3 nsew signal output
rlabel metal1 s 8918 0 8970 128 6 out1_vddio_hv
port 4 nsew signal output
rlabel metal2 s 8918 0 8970 128 6 out1_vddio_hv
port 4 nsew signal output
rlabel metal1 s 10263 0 10315 128 6 out2_vddio_hv
port 5 nsew signal output
rlabel metal2 s 10263 0 10315 128 6 out2_vddio_hv
port 5 nsew signal output
rlabel metal1 s 8701 0 8753 128 6 out2_vddd_hv
port 6 nsew signal output
rlabel metal2 s 8701 0 8753 128 6 out2_vddd_hv
port 6 nsew signal output
rlabel metal1 s 10031 0 10083 128 6 out1_vddd_hv
port 7 nsew signal output
rlabel metal2 s 10031 0 10083 128 6 out1_vddd_hv
port 7 nsew signal output
rlabel metal1 s 9784 0 9836 128 6 in1_vddio_hv
port 8 nsew signal input
rlabel metal2 s 9784 0 9836 128 6 in1_vddio_hv
port 8 nsew signal input
rlabel metal1 s 9652 377 9704 12268 6 in1_vddio_hv
port 8 nsew signal input
rlabel metal1 s 9652 291 9704 377 6 in1_vddio_hv
port 8 nsew signal input
rlabel metal1 s 9750 257 9784 291 6 in1_vddio_hv
port 8 nsew signal input
rlabel metal1 s 9784 128 9836 343 6 in1_vddio_hv
port 8 nsew signal input
rlabel metal1 s 8176 0 8228 128 6 vddio_present_vddd_hv
port 9 nsew signal output
rlabel metal2 s 8176 0 8228 128 6 vddio_present_vddd_hv
port 9 nsew signal output
rlabel metal1 s 8388 792 8440 948 6 vddio_present_vddd_hv
port 9 nsew signal output
rlabel metal1 s 8228 758 8262 792 6 vddio_present_vddd_hv
port 9 nsew signal output
rlabel metal1 s 8176 128 8228 844 6 vddio_present_vddd_hv
port 9 nsew signal output
rlabel metal1 s 1909 0 1961 128 6 vddd_present_vddio_hv
port 10 nsew signal output
rlabel metal2 s 1909 0 1961 128 6 vddd_present_vddio_hv
port 10 nsew signal output
rlabel metal1 s 1733 1900 1785 11043 6 vddd_present_vddio_hv
port 10 nsew signal output
rlabel metal1 s 1733 1814 1785 1900 6 vddd_present_vddio_hv
port 10 nsew signal output
rlabel metal1 s 1875 1780 1909 1814 6 vddd_present_vddio_hv
port 10 nsew signal output
rlabel metal1 s 1909 128 1961 1866 6 vddd_present_vddio_hv
port 10 nsew signal output
rlabel metal1 s 2483 0 2561 128 6 tie_lo_esd
port 11 nsew signal output
rlabel metal2 s 2483 0 2561 128 6 tie_lo_esd
port 11 nsew signal output
rlabel metal1 s 282 0 334 128 6 rst_por_hv_n
port 12 nsew signal input
rlabel metal2 s 282 0 334 128 6 rst_por_hv_n
port 12 nsew signal input
rlabel metal1 s 8469 0 8521 128 6 out3_vddd_hv
port 13 nsew signal output
rlabel metal2 s 8469 0 8521 128 6 out3_vddd_hv
port 13 nsew signal output
rlabel metal1 s 1415 0 1467 128 6 in3_vddio_hv
port 14 nsew signal input
rlabel metal2 s 1415 0 1467 128 6 in3_vddio_hv
port 14 nsew signal input
rlabel metal1 s 1607 13761 1641 13795 6 in3_vddio_hv
port 14 nsew signal input
rlabel metal1 s 1579 11892 1607 13795 6 in3_vddio_hv
port 14 nsew signal input
rlabel metal1 s 1324 11858 1358 11892 6 in3_vddio_hv
port 14 nsew signal input
rlabel metal1 s 1296 1252 1324 11920 6 in3_vddio_hv
port 14 nsew signal input
rlabel metal1 s 1381 1166 1415 1200 6 in3_vddio_hv
port 14 nsew signal input
rlabel metal1 s 1415 128 1467 1200 6 in3_vddio_hv
port 14 nsew signal input
rlabel metal1 s 1296 1200 1467 1252 6 in3_vddio_hv
port 14 nsew signal input
rlabel metal1 s 1579 13795 1707 13847 6 in3_vddio_hv
port 14 nsew signal input
rlabel metal1 s 1652 0 1704 128 6 in2_vddio_hv
port 15 nsew signal input
rlabel metal2 s 1652 0 1704 128 6 in2_vddio_hv
port 15 nsew signal input
rlabel metal1 s 1887 12801 1921 12835 6 in2_vddio_hv
port 15 nsew signal input
rlabel metal1 s 1859 11440 1887 12835 6 in2_vddio_hv
port 15 nsew signal input
rlabel metal1 s 1604 11406 1638 11440 6 in2_vddio_hv
port 15 nsew signal input
rlabel metal1 s 1576 2137 1604 11468 6 in2_vddio_hv
port 15 nsew signal input
rlabel metal1 s 1618 2051 1652 2085 6 in2_vddio_hv
port 15 nsew signal input
rlabel metal1 s 1652 128 1704 2085 6 in2_vddio_hv
port 15 nsew signal input
rlabel metal1 s 1859 12835 1987 12887 6 in2_vddio_hv
port 15 nsew signal input
rlabel metal1 s 1576 2085 1704 2137 6 in2_vddio_hv
port 15 nsew signal input
rlabel metal1 s 2163 0 2215 128 6 in3_vddd_hv
port 16 nsew signal input
rlabel metal2 s 2163 0 2215 128 6 in3_vddd_hv
port 16 nsew signal input
rlabel metal1 s 1813 1996 1865 10236 6 in3_vddd_hv
port 16 nsew signal input
rlabel metal1 s 2129 2131 2163 2165 6 in3_vddd_hv
port 16 nsew signal input
rlabel metal1 s 2163 128 2215 2165 6 in3_vddd_hv
port 16 nsew signal input
rlabel metal1 s 2087 2165 2215 2217 6 in3_vddd_hv
port 16 nsew signal input
rlabel metal3 s 282 0 1423 631 6 vssio_q
port 17 nsew ground bidirectional
rlabel metal3 s 1583 0 2383 25153 6 vccd
port 18 nsew power bidirectional
rlabel metal3 s 1583 27485 2501 40000 6 vccd
port 18 nsew power bidirectional
rlabel metal3 s 3703 0 4503 1208 6 vddd1
port 19 nsew power bidirectional
rlabel metal3 s 3703 28185 4503 40000 6 vddd1
port 19 nsew power bidirectional
rlabel metal3 s 4663 0 5663 7287 6 vssa
port 20 nsew ground bidirectional
rlabel metal3 s 4663 39267 5663 40000 6 vssa
port 20 nsew ground bidirectional
rlabel metal3 s 5823 0 6725 994 6 vddio_q
port 21 nsew power bidirectional
rlabel metal3 s 5823 22133 6623 40000 6 vddio_q
port 21 nsew power bidirectional
rlabel metal3 s 7000 0 7918 1655 6 vddd2
port 22 nsew power bidirectional
rlabel metal3 s 6733 27282 7908 40000 6 vddd2
port 22 nsew power bidirectional
rlabel metal3 s 2661 0 3543 6774 6 vssd
port 23 nsew ground bidirectional
rlabel metal3 s 2661 38979 3543 40000 6 vssd
port 23 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 11200 40000
string LEFclass BLOCK
string LEFsymmetry R90
string LEFview TRUE
string GDS_END 8293100
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7616778
<< end >>
