magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< pwell >>
rect -79 -26 195 226
<< nmoslvt >>
rect 0 0 30 200
rect 86 0 116 200
<< ndiff >>
rect -53 182 0 200
rect -53 148 -45 182
rect -11 148 0 182
rect -53 114 0 148
rect -53 80 -45 114
rect -11 80 0 114
rect -53 46 0 80
rect -53 12 -45 46
rect -11 12 0 46
rect -53 0 0 12
rect 30 182 86 200
rect 30 148 41 182
rect 75 148 86 182
rect 30 114 86 148
rect 30 80 41 114
rect 75 80 86 114
rect 30 46 86 80
rect 30 12 41 46
rect 75 12 86 46
rect 30 0 86 12
rect 116 182 169 200
rect 116 148 127 182
rect 161 148 169 182
rect 116 114 169 148
rect 116 80 127 114
rect 161 80 169 114
rect 116 46 169 80
rect 116 12 127 46
rect 161 12 169 46
rect 116 0 169 12
<< ndiffc >>
rect -45 148 -11 182
rect -45 80 -11 114
rect -45 12 -11 46
rect 41 148 75 182
rect 41 80 75 114
rect 41 12 75 46
rect 127 148 161 182
rect 127 80 161 114
rect 127 12 161 46
<< poly >>
rect 0 200 30 226
rect 86 200 116 226
rect 0 -26 30 0
rect 86 -26 116 0
<< locali >>
rect -45 182 -11 198
rect -45 114 -11 148
rect -45 46 -11 80
rect -45 -4 -11 12
rect 41 182 75 198
rect 41 114 75 148
rect 41 46 75 80
rect 41 -4 75 12
rect 127 182 161 198
rect 127 114 161 148
rect 127 46 161 80
rect 127 -4 161 12
use hvDFL1sd2_CDNS_52468879185133  hvDFL1sd2_CDNS_52468879185133_0
timestamp 1707688321
transform 1 0 30 0 1 0
box 0 0 1 1
use hvDFL1sd_CDNS_52468879185132  hvDFL1sd_CDNS_52468879185132_0
timestamp 1707688321
transform -1 0 0 0 1 0
box 0 0 1 1
use hvDFL1sd_CDNS_52468879185132  hvDFL1sd_CDNS_52468879185132_1
timestamp 1707688321
transform 1 0 116 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 97 -28 97 0 FreeSans 300 0 0 0 D
flabel comment s 58 97 58 97 0 FreeSans 300 0 0 0 S
flabel comment s 144 97 144 97 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 87524230
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87522840
<< end >>
