magic
tech sky130B
timestamp 1707688321
<< viali >>
rect 0 0 845 53
<< metal1 >>
rect -6 53 851 56
rect -6 0 0 53
rect 845 0 851 53
rect -6 -3 851 0
<< properties >>
string GDS_END 79754770
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 79751566
<< end >>
