##
## LEF for PtnCells ;
## created by Innovus v15.20-p005_1 on Mon Jun 14 18:10:40 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO RAM_IO
  CLASS BLOCK ;
  SIZE 100.2800 BY 219.6400 ;
  FOREIGN RAM_IO 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.43225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.685 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 12.538 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 62.643 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.3915 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.7865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.4058 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 87.968 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 7.9650 219.3100 8.1350 219.6400 ;
    END
  END N1BEG[3]
  PIN N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3952 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.455 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 46.0356 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 246.464 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 7.0450 219.3100 7.2150 219.6400 ;
    END
  END N1BEG[2]
  PIN N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.0664 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.2545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3191 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.436 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.792 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.1958 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 230.848 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 6.1250 219.3100 6.2950 219.6400 ;
    END
  END N1BEG[1]
  PIN N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.5036 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.4405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6232 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.88 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 5.2050 219.3100 5.3750 219.6400 ;
    END
  END N1BEG[0]
  PIN N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9748 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7965 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.5236 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.264 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 16.7050 219.3100 16.8750 219.6400 ;
    END
  END N2BEG[7]
  PIN N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.8904 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.3745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2511 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.0845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.562 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.7108 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 94.928 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 15.3250 219.3100 15.4950 219.6400 ;
    END
  END N2BEG[6]
  PIN N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.14325 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.345 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7816 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.2597 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.1275 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.471 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.4248 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 194.736 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 14.4050 219.3100 14.5750 219.6400 ;
    END
  END N2BEG[5]
  PIN N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.20105 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.413 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.0712 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.12 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 13.4850 219.3100 13.6550 219.6400 ;
    END
  END N2BEG[4]
  PIN N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.0695 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.1765 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.3168 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.16 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 12.1050 219.3100 12.2750 219.6400 ;
    END
  END N2BEG[3]
  PIN N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.49 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.3725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1335 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.369 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.768 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.3308 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 231.568 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 11.1850 219.3100 11.3550 219.6400 ;
    END
  END N2BEG[2]
  PIN N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.35745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.2683 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.0525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.7718 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 89.92 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 10.2650 219.3100 10.4350 219.6400 ;
    END
  END N2BEG[1]
  PIN N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.91205 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.073 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.1357 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.5075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.368 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.9518 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 90.88 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 9.3450 219.3100 9.5150 219.6400 ;
    END
  END N2BEG[0]
  PIN N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.77905 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.093 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.6528 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.8376 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 49.07 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 24.9850 219.3100 25.1550 219.6400 ;
    END
  END N2BEGb[7]
  PIN N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.81985 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.141 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.0332 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.092 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 24.0650 219.3100 24.2350 219.6400 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.3254 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.553 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 22.6850 219.3100 22.8550 219.6400 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.3748 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.7965 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.3444 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.604 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 21.7650 219.3100 21.9350 219.6400 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.7648 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 63.588 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 20.8450 219.3100 21.0150 219.6400 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5095 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3765 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 46.8156 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 250.624 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 19.4650 219.3100 19.6350 219.6400 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1517 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 56.3718 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 301.12 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 18.5450 219.3100 18.7150 219.6400 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1852 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.8485 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.7029 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.3435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.023 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.5524 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.024 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 17.6250 219.3100 17.7950 219.6400 ;
    END
  END N2BEGb[0]
  PIN N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.77905 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.093 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0732 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3149 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.781 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.4418 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 264.16 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 41.5450 219.3100 41.7150 219.6400 ;
    END
  END N4BEG[15]
  PIN N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.4496 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 27.1705 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4353 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.7338 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 244.384 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 40.6250 219.3100 40.7950 219.6400 ;
    END
  END N4BEG[14]
  PIN N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.8256 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.0505 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3047 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3525 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.0608 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 214.128 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 39.7050 219.3100 39.8750 219.6400 ;
    END
  END N4BEG[13]
  PIN N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.6832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.3385 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8679 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.1685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.99 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.08 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.6278 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 137.152 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 38.7850 219.3100 38.9550 219.6400 ;
    END
  END N4BEG[12]
  PIN N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.246 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.1525 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9557 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.6075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.687 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.1896 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 17.952 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 37.4050 219.3100 37.5750 219.6400 ;
    END
  END N4BEG[11]
  PIN N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.6256 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 33.0505 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.964 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.702 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 36.4850 219.3100 36.6550 219.6400 ;
    END
  END N4BEG[10]
  PIN N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.83725 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.985 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 7.0274 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 35.063 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 35.5650 219.3100 35.7350 219.6400 ;
    END
  END N4BEG[9]
  PIN N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.3276 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.5605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.2016 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.89 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 34.1850 219.3100 34.3550 219.6400 ;
    END
  END N4BEG[8]
  PIN N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.16 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.4356 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 27.1005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.5492 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.628 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 33.2650 219.3100 33.4350 219.6400 ;
    END
  END N4BEG[7]
  PIN N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2239 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 61.4718 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 328.32 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 32.3450 219.3100 32.5150 219.6400 ;
    END
  END N4BEG[6]
  PIN N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1959 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.8085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.6178 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 318.432 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 31.4250 219.3100 31.5950 219.6400 ;
    END
  END N4BEG[5]
  PIN N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.77905 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.093 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.88 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1212 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.488 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 30.0450 219.3100 30.2150 219.6400 ;
    END
  END N4BEG[4]
  PIN N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.93545 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.277 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7404 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.584 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 29.1250 219.3100 29.2950 219.6400 ;
    END
  END N4BEG[3]
  PIN N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.8768 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.3065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.09 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.332 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 28.2050 219.3100 28.3750 219.6400 ;
    END
  END N4BEG[2]
  PIN N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.461 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3308 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1572 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.668 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 26.8250 219.3100 26.9950 219.6400 ;
    END
  END N4BEG[1]
  PIN N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2496 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.13 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 25.9050 219.3100 26.0750 219.6400 ;
    END
  END N4BEG[0]
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.72125 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.025 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.562 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.936 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.4615 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 270.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 441.406 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2322.26 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 7.9650 0.0000 8.1350 0.3300 ;
    END
  END N1END[3]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.1124 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.897 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0578 LAYER mcon  ;
    ANTENNADIFFAREA 0.1872 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 6.7037 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 33.2185 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0675 LAYER via  ;
    ANTENNADIFFAREA 0.936 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.066 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 129.514 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 169.819 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 827.827 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 7.0450 0.0000 7.2150 0.3300 ;
    END
  END N1END[2]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9752 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.7985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.936 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 14.4784 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 71.596 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 101.22 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 484.277 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.46478 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 6.1250 0.0000 6.2950 0.3300 ;
    END
  END N1END[1]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.0288 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 29.925 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met1  ;
    ANTENNAMAXAREACAR 41.584 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 190.893 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via  ;
    ANTENNADIFFAREA 0.936 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.96 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 53.984 LAYER met2  ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 110.515 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 530.415 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 5.2050 0.0000 5.3750 0.3300 ;
    END
  END N1END[0]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 0.1872 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.79 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.8355 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4072 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.918 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 0.956768 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 3.48013 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 16.7050 0.0000 16.8750 0.3300 ;
    END
  END N2MID[7]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.5752 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.65 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 8.90343 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 42.9771 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 15.3250 0.0000 15.4950 0.3300 ;
    END
  END N2MID[6]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.70425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.7176 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.352 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.71589 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 35.8869 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0995286 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 14.4050 0.0000 14.5750 0.3300 ;
    END
  END N2MID[5]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6868 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2183 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.1872 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 58.4568 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 312.24 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 97.2275 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 516.533 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.207273 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 13.4850 0.0000 13.6550 0.3300 ;
    END
  END N2MID[4]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1872 LAYER li1  ;
    ANTENNAPARTIALMETALAREA 24.0676 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 28.282 LAYER li1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER li1  ;
    ANTENNAMAXAREACAR 32.4143 LAYER li1  ;
    ANTENNAMAXSIDEAREACAR 38.0902 LAYER li1  ;
    PORT
      LAYER li1 ;
        RECT 12.1050 0.0000 12.2750 0.3300 ;
    END
  END N2MID[3]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.3244 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.5445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.004 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.784 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.87838 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.6929 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0995286 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 11.1850 0.0000 11.3550 0.3300 ;
    END
  END N2MID[2]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.81145 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.837 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.5437 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.5735 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met1  ;
    ANTENNAMAXAREACAR 5.40667 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 24.4155 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.8832 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.298 LAYER met2  ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.59616 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 30.204 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 10.2650 0.0000 10.4350 0.3300 ;
    END
  END N2MID[1]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3952 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4769 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2135 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.506 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.1872 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.8318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 282.24 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 94.2916 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 500.129 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 9.3450 0.0000 9.5150 0.3300 ;
    END
  END N2MID[0]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08545 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.277 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2729 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.1908 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.1458 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 209.248 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 24.9850 0.0000 25.1550 0.3300 ;
    END
  END N2END[7]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.7512 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.2984 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.374 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 24.0650 0.0000 24.2350 0.3300 ;
    END
  END N2END[6]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.7816 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.7104 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.434 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 22.6850 0.0000 22.8550 0.3300 ;
    END
  END N2END[5]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.29965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.5208 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.5265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3107 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3825 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.161 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.1908 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.6214 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 127.392 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 21.7650 0.0000 21.9350 0.3300 ;
    END
  END N2END[4]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6001 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8295 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.1908 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.4688 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 152.304 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 20.8450 0.0000 21.0150 0.3300 ;
    END
  END N2END[3]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.20105 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.413 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.6978 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.4115 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.978 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.772 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 19.4650 0.0000 19.6350 0.3300 ;
    END
  END N2END[2]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.6296 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.03 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 18.5450 0.0000 18.7150 0.3300 ;
    END
  END N2END[1]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.6408 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.0895 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1829 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1908 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.3268 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.88 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 17.6250 0.0000 17.7950 0.3300 ;
    END
  END N2END[0]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.461 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.9812 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 34.8285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 27.2928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 136.346 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 39.2124 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 194.667 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 41.5450 0.0000 41.7150 0.3300 ;
    END
  END N4END[15]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.3508 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 36.6765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 15.2974 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 76.251 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 23.172 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 114.306 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 40.6250 0.0000 40.7950 0.3300 ;
    END
  END N4END[14]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.461 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.0224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.5492 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.628 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.25623 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 33.8929 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 39.7050 0.0000 39.8750 0.3300 ;
    END
  END N4END[13]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.524 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.8227 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 43.9425 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 40.2438 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 215.104 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 56.0768 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 298.541 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 38.7850 0.0000 38.9550 0.3300 ;
    END
  END N4END[12]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1569 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5985 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 52.5594 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 281.728 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 78.6652 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 418.187 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 37.4050 0.0000 37.5750 0.3300 ;
    END
  END N4END[11]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2164 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.964 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 2.0466 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 8.92929 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 36.4850 0.0000 36.6550 0.3300 ;
    END
  END N4END[10]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.748 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6625 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.678 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.272 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.38027 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.2013 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 35.5650 0.0000 35.7350 0.3300 ;
    END
  END N4END[9]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.8513 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.9675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 34.5066 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 184.976 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 55.3836 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 294.1 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 34.1850 0.0000 34.3550 0.3300 ;
    END
  END N4END[8]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.47305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5884 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1073 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.7024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.824 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 20.196 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 101.674 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 33.2650 0.0000 33.4350 0.3300 ;
    END
  END N4END[7]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.0528 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.1865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 9.2731 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.9585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 30.9816 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 166.176 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 49.7956 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 263.467 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 32.3450 0.0000 32.5150 0.3300 ;
    END
  END N4END[6]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.992 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.539 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 50.5638 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 270.144 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 78.8928 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 417.321 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 31.4250 0.0000 31.5950 0.3300 ;
    END
  END N4END[5]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3191 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.6676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 100.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.7658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.888 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 15.9471 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 84.6451 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 30.0450 0.0000 30.2150 0.3300 ;
    END
  END N4END[4]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6607 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.5286 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 147.76 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 262.437 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1379 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 29.1250 0.0000 29.2950 0.3300 ;
    END
  END N4END[3]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96985 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.141 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.7645 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 28.637 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.045 LAYER via  ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.255 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 35.707 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 0.1908 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.6688 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.504 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 76.4211 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 391.057 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.7087 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 254.912 LAYER met4  ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 376.476 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1994.28 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 28.2050 0.0000 28.3750 0.3300 ;
    END
  END N4END[2]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.3816 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.1876 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 55.454 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 80.9412 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 384.846 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via2  ;
    ANTENNADIFFAREA 0.7632 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.6708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.048 LAYER met3  ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 85.1601 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 410.305 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 26.8250 0.0000 26.9950 0.3300 ;
    END
  END N4END[1]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.08545 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.277 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2977 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.7766 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 218.416 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.492 LAYER met4  ;
    ANTENNAMAXAREACAR 107.425 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 561.645 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.312805 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 25.9050 0.0000 26.0750 0.3300 ;
    END
  END N4END[0]
  PIN E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5553 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.6685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5161 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.4095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.783 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.976 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3104 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.1539 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 195.168 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 84.7600 0.5950 84.9000 ;
    END
  END E1END[3]
  PIN E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0384 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.084 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.3744 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.025 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.728 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3744 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.381 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.832 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3104 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5186 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.04 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 83.4000 0.5950 83.5400 ;
    END
  END E1END[2]
  PIN E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2641 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3905 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7815 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.3104 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.5567 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.768 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 81.3600 0.5950 81.5000 ;
    END
  END E1END[1]
  PIN E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3317 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5505 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.3104 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 19.8636 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 98.168 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 80.3400 0.5950 80.4800 ;
    END
  END E1END[0]
  PIN E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7765 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.7745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5616 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.5808 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.432 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 96.6600 0.5950 96.8000 ;
    END
  END E2MID[7]
  PIN E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0537 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.1605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3803 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7305 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3744 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.8818 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 85.64 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5616 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.0346 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 59.792 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 94.9600 0.5950 95.1000 ;
    END
  END E2MID[6]
  PIN E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4741 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2625 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5616 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.097 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 93.6000 0.5950 93.7400 ;
    END
  END E2MID[5]
  PIN E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3417 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.6005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.3744 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.881 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.782 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5616 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.0278 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.952 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 92.2400 0.5950 92.3800 ;
    END
  END E2MID[4]
  PIN E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3621 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.7025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.4119 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.8885 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5652 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.4648 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.616 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 90.2000 0.5950 90.3400 ;
    END
  END E2MID[3]
  PIN E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6537 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5652 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.8984 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 48.902 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 88.8400 0.5950 88.9800 ;
    END
  END E2MID[2]
  PIN E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2129 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.9565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.4353 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.7665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5652 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.5198 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.576 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 87.8200 0.5950 87.9600 ;
    END
  END E2MID[1]
  PIN E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6337 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.0605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.6411 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.0345 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.298 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.056 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5652 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.5958 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.648 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 86.1200 0.5950 86.2600 ;
    END
  END E2MID[0]
  PIN E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2343 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.0635 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.5075 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.3665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.895 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.24 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5724 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.6166 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.896 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 108.2200 0.5950 108.3600 ;
    END
  END E2END[7]
  PIN E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1689 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7365 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.2381 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.0195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.048 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.056 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5724 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.1318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.84 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 106.5200 0.5950 106.6600 ;
    END
  END E2END[6]
  PIN E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.6101 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.9425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2007 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.8325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5724 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.3628 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 29.072 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 105.5000 0.5950 105.6400 ;
    END
  END E2END[5]
  PIN E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.7837 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 28.7735 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5724 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.0662 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 19.761 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 103.8000 0.5950 103.9400 ;
    END
  END E2END[4]
  PIN E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8877 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.3305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5688 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.3868 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.472 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 102.4400 0.5950 102.5800 ;
    END
  END E2END[3]
  PIN E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3085 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.4345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.6681 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 33.1695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.5958 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 19.648 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 101.0800 0.5950 101.2200 ;
    END
  END E2END[2]
  PIN E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7625 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.7045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2459 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5688 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 23.6535 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 127.088 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 99.3800 0.5950 99.5200 ;
    END
  END E2END[1]
  PIN E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6537 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.7999 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.8285 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.8516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 58.816 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 98.0200 0.5950 98.1600 ;
    END
  END E2END[0]
  PIN EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6537 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 8.5369 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 42.3955 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1908 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.9678 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.3986 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 40.4 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 132.0200 0.5950 132.1600 ;
    END
  END EE4END[15]
  PIN EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1872 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.1547 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.561 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.378 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.2365 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.9035 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.378 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.129 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 86.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5688 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.0676 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.968 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 130.3200 0.5950 130.4600 ;
    END
  END EE4END[14]
  PIN EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1385 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.378 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.1113 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 55.1495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5688 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.3168 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.16 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 128.9600 0.5950 129.1000 ;
    END
  END EE4END[13]
  PIN EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7407 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.5585 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5688 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.9322 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.199 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 127.6000 0.5950 127.7400 ;
    END
  END EE4END[12]
  PIN EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7973 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.7705 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.045 LAYER via  ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3815 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.6185 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3816 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 17.2278 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 92.352 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 125.9000 0.5950 126.0400 ;
    END
  END EE4END[11]
  PIN EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3929 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8931 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3816 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.5592 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 148.864 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 124.5400 0.5950 124.6800 ;
    END
  END EE4END[10]
  PIN EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4265 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.3816 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.9984 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.638 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 123.1800 0.5950 123.3200 ;
    END
  END EE4END[9]
  PIN EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2981 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.3816 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.3544 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 46.536 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 121.4800 0.5950 121.6200 ;
    END
  END EE4END[8]
  PIN EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2435 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7485 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.5715 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.8508 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.378 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.6895 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 47.28 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 120.1200 0.5950 120.2600 ;
    END
  END EE4END[7]
  PIN EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2505 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.378 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.1744 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 45.528 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 118.7600 0.5950 118.9000 ;
    END
  END EE4END[6]
  PIN EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9057 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.3835 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.1747 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.5945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1908 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.815 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.48 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.378 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.2168 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 6.96 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 117.0600 0.5950 117.2000 ;
    END
  END EE4END[5]
  PIN EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1872 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.4546 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.0605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.378 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5284 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.406 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 115.7000 0.5950 115.8400 ;
    END
  END EE4END[4]
  PIN EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8173 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.8705 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.045 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.0475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5652 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 19.6188 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 105.104 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 114.3400 0.5950 114.4800 ;
    END
  END EE4END[3]
  PIN EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3929 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.1445 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.5515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.505 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.16 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.5652 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.4934 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 41.376 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 112.6400 0.5950 112.7800 ;
    END
  END EE4END[2]
  PIN EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.1085 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.4345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5652 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.7944 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.52 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 111.2800 0.5950 111.4200 ;
    END
  END EE4END[1]
  PIN EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9633 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.6715 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5652 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.0764 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.812 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 109.9200 0.5950 110.0600 ;
    END
  END EE4END[0]
  PIN E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3317 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5505 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4699 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.1785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7524 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.5268 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 83.28 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 149.7000 0.5950 149.8400 ;
    END
  END E6END[11]
  PIN E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8437 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6361 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.14 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7524 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 10.0008 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 53.808 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 148.0000 0.5950 148.1400 ;
    END
  END E6END[10]
  PIN E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5293 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.5015 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5652 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.4415 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.4665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.5652 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.3578 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.512 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7524 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.7788 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 20.624 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 146.6400 0.5950 146.7800 ;
    END
  END E6END[9]
  PIN E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1825 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.8045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6649 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1535 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7524 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.9148 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.016 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 145.2800 0.5950 145.4200 ;
    END
  END E6END[8]
  PIN E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.1872 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.2972 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.2365 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.7405 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.5315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3744 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 22.0679 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 118.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNADIFFAREA 0.7524 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 39.0576 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 209.248 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 143.5800 0.5950 143.7200 ;
    END
  END E6END[7]
  PIN E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3317 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5505 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.378 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.8415 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.6925 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.378 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7524 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.2668 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 28.56 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 142.2200 0.5950 142.3600 ;
    END
  END E6END[6]
  PIN E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2473 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.1285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.9681 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 29.6695 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.665 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7524 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.7296 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 68.832 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 140.8600 0.5950 141.0000 ;
    END
  END E6END[5]
  PIN E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4573 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.1785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.5616 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 11.5163 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.4865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.7524 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 139.1600 0.5950 139.3000 ;
    END
  END E6END[4]
  PIN E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4701 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.0975 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.045 LAYER via  ;
    ANTENNADIFFAREA 0.3744 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.8012 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.438 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNADIFFAREA 0.5652 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.3967 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.056 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.756 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.8938 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 95.904 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 137.8000 0.5950 137.9400 ;
    END
  END E6END[3]
  PIN E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0197 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.9905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.3013 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.2175 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1872 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.9821 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.756 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 136.4400 0.5950 136.5800 ;
    END
  END E6END[2]
  PIN E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.4329 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 26.9115 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.045 LAYER via  ;
    ANTENNADIFFAREA 0.378 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8005 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.4875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.756 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.6387 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.872 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 134.7400 0.5950 134.8800 ;
    END
  END E6END[1]
  PIN E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.5141 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 27.3175 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.045 LAYER via  ;
    ANTENNADIFFAREA 0.5688 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.2572 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.632 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.756 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.3268 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.88 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 133.3800 0.5950 133.5200 ;
    END
  END E6END[0]
  PIN S1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.16 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.1036 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.4405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.3005 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.285 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.4538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 88.224 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 45.6850 0.0000 45.8550 0.3300 ;
    END
  END S1BEG[3]
  PIN S1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.43225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.685 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 0.368 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 7.5916 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 37.884 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 44.7650 0.0000 44.9350 0.3300 ;
    END
  END S1BEG[2]
  PIN S1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.12625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.6528 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1865 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 12.422 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 61.992 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 43.8450 0.0000 44.0150 0.3300 ;
    END
  END S1BEG[1]
  PIN S1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3135 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.4 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.8668 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 239.76 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 42.9250 0.0000 43.0950 0.3300 ;
    END
  END S1BEG[0]
  PIN S2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2183 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9205 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.78 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 41.5008 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 221.808 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 62.7050 0.0000 62.8750 0.3300 ;
    END
  END S2BEG[7]
  PIN S2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96985 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.141 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 0.368 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.87 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 24.276 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 61.7850 0.0000 61.9550 0.3300 ;
    END
  END S2BEG[6]
  PIN S2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.1004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.8816 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.29 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 60.4050 0.0000 60.5750 0.3300 ;
    END
  END S2BEG[5]
  PIN S2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1208 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2659 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.677 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.3768 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 194.48 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 59.4850 0.0000 59.6550 0.3300 ;
    END
  END S2BEG[4]
  PIN S2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.41525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3863 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7605 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.0328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 155.312 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 58.5650 0.0000 58.7350 0.3300 ;
    END
  END S2BEG[3]
  PIN S2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.31665 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.549 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.524 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.368 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.36 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.682 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 57.6450 0.0000 57.8150 0.3300 ;
    END
  END S2BEG[2]
  PIN S2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.20105 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.413 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9454 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.6495 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8987 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.263 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.2468 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 87.12 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 56.2650 0.0000 56.4350 0.3300 ;
    END
  END S2BEG[1]
  PIN S2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.31665 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.549 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8511 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0845 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.987 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.368 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.4768 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 237.68 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 55.3450 0.0000 55.5150 0.3300 ;
    END
  END S2BEG[0]
  PIN S2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8315 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.9865 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.333 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.5668 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 126.16 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 54.4250 0.0000 54.5950 0.3300 ;
    END
  END S2BEGb[7]
  PIN S2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.3104 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.4745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.406 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.912 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 53.0450 0.0000 53.2150 0.3300 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.16065 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.189 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.5014 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 27.4295 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.8676 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.22 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 52.1250 0.0000 52.2950 0.3300 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.91205 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.073 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2664 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4195 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.9265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.125 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.5158 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 253.888 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 51.2050 0.0000 51.3750 0.3300 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.91205 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.073 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.3444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4157 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.9075 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.481 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.032 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.1028 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 134.352 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 50.2850 0.0000 50.4550 0.3300 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.6928 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.346 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 48.9050 0.0000 49.0750 0.3300 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.44965 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.529 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.0496 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.1705 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.7396 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.58 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 47.9850 0.0000 48.1550 0.3300 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5884 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2109 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.8835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.817 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.824 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 51.9798 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 277.696 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 47.0650 0.0000 47.2350 0.3300 ;
    END
  END S2BEGb[0]
  PIN S4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.64645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0079 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.8685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 32.5578 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 174.112 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 79.2650 0.0000 79.4350 0.3300 ;
    END
  END S4BEG[15]
  PIN S4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.0932 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 40.348 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 78.3450 0.0000 78.5150 0.3300 ;
    END
  END S4BEG[14]
  PIN S4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.4224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.0863 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2605 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.987 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.4676 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 152.768 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 77.4250 0.0000 77.5950 0.3300 ;
    END
  END S4BEG[13]
  PIN S4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.37445 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.617 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.6224 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9743 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.7005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.953 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.4818 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 131.04 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 76.5050 0.0000 76.6750 0.3300 ;
    END
  END S4BEG[12]
  PIN S4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.31665 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.549 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.142 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.5955 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1855 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6755 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.5928 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.632 LAYER met3  ;
    PORT
      LAYER li1 ;
        RECT 75.1250 0.0000 75.2950 0.3300 ;
    END
  END S4BEG[11]
  PIN S4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.1376 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9472 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.618 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 74.2050 0.0000 74.3750 0.3300 ;
    END
  END S4BEG[10]
  PIN S4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7083 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.3705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 54.5178 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 291.232 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 73.2850 0.0000 73.4550 0.3300 ;
    END
  END S4BEG[9]
  PIN S4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.02765 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.209 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.3385 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.394 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 72.3650 0.0000 72.5350 0.3300 ;
    END
  END S4BEG[8]
  PIN S4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.31665 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.549 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1507 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5825 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 49.5768 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 264.88 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 70.9850 0.0000 71.1550 0.3300 ;
    END
  END S4BEG[7]
  PIN S4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.5508 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.6765 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2284 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.906 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 70.0650 0.0000 70.2350 0.3300 ;
    END
  END S4BEG[6]
  PIN S4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.54785 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.821 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.9748 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7965 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.4072 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.918 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 69.1450 0.0000 69.3150 0.3300 ;
    END
  END S4BEG[5]
  PIN S4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.14325 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.345 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.582 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.8325 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4815 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 53.0538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 283.424 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 67.7650 0.0000 67.9350 0.3300 ;
    END
  END S4BEG[4]
  PIN S4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.14325 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.345 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.0664 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.2545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0904 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.334 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 66.8450 0.0000 67.0150 0.3300 ;
    END
  END S4BEG[3]
  PIN S4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.62305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 7.5734 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 37.793 LAYER met1  ;
    PORT
      LAYER li1 ;
        RECT 65.9250 0.0000 66.0950 0.3300 ;
    END
  END S4BEG[2]
  PIN S4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.79645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.5172 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.5085 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.2024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.894 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 65.0050 0.0000 65.1750 0.3300 ;
    END
  END S4BEG[1]
  PIN S4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.49005 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.753 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.3596 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.68 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 63.6250 0.0000 63.7950 0.3300 ;
    END
  END S4BEG[0]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.1952 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.8985 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1929 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.6665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1872 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.936 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.3295 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 141.36 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 171.621 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 916.164 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 45.6850 219.3100 45.8550 219.6400 ;
    END
  END S1END[3]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.27625 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.325 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0732 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.2315 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.7605 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1872 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.126 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.936 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.7153 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 271.888 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 383.009 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 2046.36 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 44.7650 219.3100 44.9350 219.6400 ;
    END
  END S1END[2]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.33405 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.393 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.504 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.4425 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.6679 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.1685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.021 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.936 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.7388 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 137.744 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 219.736 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1149.01 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.10943 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 43.8450 219.3100 44.0150 219.6400 ;
    END
  END S1END[1]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.25885 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.481 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4607 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1872 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.936 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.4498 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 29.536 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 71.4365 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 380.079 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 42.9250 219.3100 43.0950 219.6400 ;
    END
  END S1END[0]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.77905 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.093 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.5867 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.6445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.932 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.104 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.1872 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.4258 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 29.408 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 11.3865 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 59.4774 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 62.7050 219.3100 62.8750 219.6400 ;
    END
  END S2MID[7]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.14325 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.345 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 4.4504 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.1375 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 26.8724 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 134.008 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 37.9976 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 188.275 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 61.7850 219.3100 61.9550 219.6400 ;
    END
  END S2MID[6]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.47305 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.733 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 7.0456 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 35.1505 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.6313 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.8675 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.78 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.1872 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.9988 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 32.464 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 12.2512 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 64.0889 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 60.4050 219.3100 60.5750 219.6400 ;
    END
  END S2MID[5]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.8156 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.0005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1872 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.0448 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.752 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 9.84599 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 46.2195 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0995286 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 59.4850 219.3100 59.6550 219.6400 ;
    END
  END S2MID[4]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.77905 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.093 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.6283 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.9705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.092 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.624 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.1872 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 26.2999 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 134.896 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 58.5650 219.3100 58.7350 219.6400 ;
    END
  END S2MID[3]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.461 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1673 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6265 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.1872 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 60.3498 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 322.336 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 84.5665 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 449.464 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 57.6450 219.3100 57.8150 219.6400 ;
    END
  END S2MID[2]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.64645 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.937 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4936 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.3905 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7237 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4475 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.1872 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 44.5236 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 238.4 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 72.8047 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 384.859 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 56.2650 219.3100 56.4350 219.6400 ;
    END
  END S2MID[1]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.77905 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.093 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8917 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.1872 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.5036 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.96 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 11.789 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 62.1145 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 55.3450 219.3100 55.5150 219.6400 ;
    END
  END S2MID[0]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.10585 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.301 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.9452 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 34.6115 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.026 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.012 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 54.4250 219.3100 54.5950 219.6400 ;
    END
  END S2END[7]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3191 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.1908 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.5866 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 270.736 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 53.0450 219.3100 53.2150 219.6400 ;
    END
  END S2END[6]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.45265 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.709 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.9712 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.7785 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0996 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.262 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 52.1250 219.3100 52.2950 219.6400 ;
    END
  END S2END[5]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.41225 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.485 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.5884 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.8645 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.292 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.224 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 51.2050 219.3100 51.3750 219.6400 ;
    END
  END S2END[4]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.56825 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.845 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.8764 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.3045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4332 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.93 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 50.2850 219.3100 50.4550 219.6400 ;
    END
  END S2END[3]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.77905 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.093 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.4292 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0685 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7667 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6625 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.1908 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 53.2368 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 284.4 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 48.9050 219.3100 49.0750 219.6400 ;
    END
  END S2END[2]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.85425 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.005 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.236 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1025 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8031 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8445 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.224 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.1908 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.2906 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 231.824 LAYER met4  ;
    PORT
      LAYER li1 ;
        RECT 47.9850 219.3100 48.1550 219.6400 ;
    END
  END S2END[1]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.2768 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.3065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.6232 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.88 LAYER met2  ;
    PORT
      LAYER li1 ;
        RECT 47.0650 219.3100 47.2350 219.6400 ;
    END
  END S2END[0]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 6.2896 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 31.3705 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2636 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.2 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.57603 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 16.4855 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 79.2650 219.3100 79.4350 219.6400 ;
    END
  END S4END[15]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.10285 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.121 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.0088 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.9665 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1335 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5355 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.538 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.336 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 51.2718 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 273.92 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 77.716 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 412.345 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 78.3450 219.3100 78.5150 219.6400 ;
    END
  END S4END[14]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.31665 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.549 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.2496 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.1705 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.9304 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.534 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.64256 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 26.8182 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 77.4250 219.3100 77.5950 219.6400 ;
    END
  END S4END[13]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.136 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.16 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.4848 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 12.3095 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4557 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.9895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 37.8408 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 202.288 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 58.3912 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 311.434 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 76.5050 219.3100 76.6750 219.6400 ;
    END
  END S4END[12]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.03105 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.213 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 2.1988 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.9165 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.7876 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.82 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 3.36828 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 14.4532 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 75.1250 219.3100 75.2950 219.6400 ;
    END
  END S4END[11]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.73865 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.869 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 3.3748 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.7965 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 16.0453 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 80.0555 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.781 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 31.5318 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 168.64 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 50.7766 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 267.946 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 74.2050 219.3100 74.3750 219.6400 ;
    END
  END S4END[10]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.77905 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.093 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.1716 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.1727 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.6925 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 51.1998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 273.536 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 77.9341 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 412.226 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 73.2850 219.3100 73.4550 219.6400 ;
    END
  END S4END[9]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.68085 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.801 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.9444 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.6445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.6472 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.118 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.17939 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 19.5024 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 72.3650 219.3100 72.5350 219.6400 ;
    END
  END S4END[8]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56525 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.665 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3004 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.7925 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.7915 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.171 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.712 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 53.5788 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 286.224 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 79.8193 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 422.362 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 70.9850 219.3100 71.1550 219.6400 ;
    END
  END S4END[7]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.21845 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.257 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.3784 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8145 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.5512 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.638 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.7437 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 32.3239 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 70.0650 219.3100 70.2350 219.6400 ;
    END
  END S4END[6]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50745 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.597 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 5.2012 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 25.8545 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.5697 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.2872 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 126.08 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 33.3119 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 178.173 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER li1 ;
        RECT 69.1450 219.3100 69.3150 219.6400 ;
    END
  END S4END[5]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.96985 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.141 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 9.6976 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 48.3735 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 19.1252 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 95.508 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 26.8057 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 132.634 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 67.7650 219.3100 67.9350 219.6400 ;
    END
  END S4END[4]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.66345 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.957 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.0832 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.406 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.6419 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.0385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3816 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.2549 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.488 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.3996 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 66.592 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 87.3094 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 462.557 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 66.8450 219.3100 67.0150 219.6400 ;
    END
  END S4END[3]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.56825 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.845 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0578 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 10.4152 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 51.884 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.045 LAYER via  ;
    ANTENNADIFFAREA 0.1908 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 18.5313 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 92.2495 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 123.757 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 610.28 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via2  ;
    ANTENNADIFFAREA 0.1908 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.992 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.424 LAYER met3  ;
    ANTENNAGATEAREA 0.159 LAYER met3  ;
    ANTENNAMAXAREACAR 199.178 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 1015.46 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.5663 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 73.76 LAYER met4  ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 284.501 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1479.36 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.967925 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 65.9250 219.3100 66.0950 219.6400 ;
    END
  END S4END[2]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.31665 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.549 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 1.958 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2459 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.297 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7632 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.0918 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 144.96 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 265.692 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1393.63 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.10943 LAYER via4  ;
    PORT
      LAYER li1 ;
        RECT 65.0050 219.3100 65.1750 219.6400 ;
    END
  END S4END[1]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.39185 LAYER li1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.461 LAYER li1  ;
    ANTENNAPARTIALCUTAREA 0.0289 LAYER mcon  ;
    ANTENNAPARTIALMETALAREA 0.3648 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 0.7632 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 10.2222 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.197 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.492 LAYER met2  ;
    ANTENNAMAXAREACAR 22.5464 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 109.874 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.104472 LAYER via2  ;
    PORT
      LAYER li1 ;
        RECT 63.6250 219.3100 63.7950 219.6400 ;
    END
  END S4END[0]
  PIN W1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7181 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4535 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0965 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.536 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 125.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.1528 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 139.952 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 14.0400 0.5950 14.1800 ;
    END
  END W1BEG[3]
  PIN W1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2029 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.8073 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.909 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 90.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.8638 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 15.744 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 12.6800 0.5950 12.8200 ;
    END
  END W1BEG[2]
  PIN W1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9665 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 19.6875 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.6452 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 38.108 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 11.3200 0.5950 11.4600 ;
    END
  END W1BEG[1]
  PIN W1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6133 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 52.9585 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.932 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.542 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 9.9600 0.5950 10.1000 ;
    END
  END W1BEG[0]
  PIN W2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.1321 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.556 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 25.9400 0.5950 26.0800 ;
    END
  END W2BEG[7]
  PIN W2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3217 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 21.5005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9308 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.536 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 24.5800 0.5950 24.7200 ;
    END
  END W2BEG[6]
  PIN W2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7181 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9657 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.5395 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.6166 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.896 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 22.8800 0.5950 23.0200 ;
    END
  END W2BEG[5]
  PIN W2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0384 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.084 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 14.8677 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 74.0495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.953 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.8776 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 80.288 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 21.5200 0.5950 21.6600 ;
    END
  END W2BEG[4]
  PIN W2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3317 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5505 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3331 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.4945 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.635 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.5208 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 163.248 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 20.1600 0.5950 20.3000 ;
    END
  END W2BEG[3]
  PIN W2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.0941 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 30.3625 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.7468 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.38 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 18.4600 0.5950 18.6000 ;
    END
  END W2BEG[2]
  PIN W2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2129 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.9565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2841 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2495 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.127 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.8186 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 106.64 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 17.1000 0.5950 17.2400 ;
    END
  END W2BEG[1]
  PIN W2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3961 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6145 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.9015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.125 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 45.3198 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 242.176 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 15.7400 0.5950 15.8800 ;
    END
  END W2BEG[0]
  PIN W2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3929 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1439 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.253 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.816 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 36.8148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 196.816 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 37.8400 0.5950 37.9800 ;
    END
  END W2BEGb[7]
  PIN W2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.9137 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.464 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 36.1400 0.5950 36.2800 ;
    END
  END W2BEGb[6]
  PIN W2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5625 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.7045 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.2644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.204 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 34.7800 0.5950 34.9200 ;
    END
  END W2BEGb[5]
  PIN W2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1045 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4145 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1829 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.1862 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 216.208 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 33.4200 0.5950 33.5600 ;
    END
  END W2BEGb[4]
  PIN W2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1385 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6789 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.2235 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.992 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.972 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 167.536 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 31.7200 0.5950 31.8600 ;
    END
  END W2BEGb[3]
  PIN W2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.2917 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 11.354 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 30.3600 0.5950 30.5000 ;
    END
  END W2BEGb[2]
  PIN W2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4677 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.2305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2239 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.543 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.5116 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 78.336 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 29.0000 0.5950 29.1400 ;
    END
  END W2BEGb[1]
  PIN W2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6537 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.8707 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.1825 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.376 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.9492 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 166.944 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 27.3000 0.5950 27.4400 ;
    END
  END W2BEGb[0]
  PIN WW4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7489 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6365 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2953 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.818 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 47.496 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.3086 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 135.92 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 61.3000 0.5950 61.4400 ;
    END
  END WW4BEG[15]
  PIN WW4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.8577 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.184 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 59.9400 0.5950 60.0800 ;
    END
  END WW4BEG[14]
  PIN WW4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 9.1797 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 45.794 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 58.2400 0.5950 58.3800 ;
    END
  END WW4BEG[13]
  PIN WW4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2505 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.4541 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.0995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.06 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 54.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.0372 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.08 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 56.8800 0.5950 57.0200 ;
    END
  END WW4BEG[12]
  PIN WW4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2029 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3359 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.7958 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 90.048 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 55.5200 0.5950 55.6600 ;
    END
  END WW4BEG[11]
  PIN WW4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0677 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 10.2305 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2361 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.607 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.3518 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 23.68 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 53.8200 0.5950 53.9600 ;
    END
  END WW4BEG[10]
  PIN WW4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7135 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.4225 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6523 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.0905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.425 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 77.4 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.9878 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.072 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 52.4600 0.5950 52.6000 ;
    END
  END WW4BEG[9]
  PIN WW4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1045 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4145 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.4065 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.8615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 29.8434 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 160.576 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 51.1000 0.5950 51.2400 ;
    END
  END WW4BEG[8]
  PIN WW4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.5979 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.885 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 49.4000 0.5950 49.5400 ;
    END
  END WW4BEG[7]
  PIN WW4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.6105 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.948 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 48.0400 0.5950 48.1800 ;
    END
  END WW4BEG[6]
  PIN WW4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7593 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.6885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.0243 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.9505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.139 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 49.208 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.8204 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 11.12 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 46.6800 0.5950 46.8200 ;
    END
  END WW4BEG[5]
  PIN WW4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3317 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5505 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4451 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 88.328 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 11.2818 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 60.64 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 44.9800 0.5950 45.1200 ;
    END
  END WW4BEG[4]
  PIN WW4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6537 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1059 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.3585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.401 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.272 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.8678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 74.432 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 43.6200 0.5950 43.7600 ;
    END
  END WW4BEG[3]
  PIN WW4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6469 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 18.1265 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.1212 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.488 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 42.2600 0.5950 42.4000 ;
    END
  END WW4BEG[2]
  PIN WW4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6977 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.3805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4087 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.8725 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1905 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 6.2766 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 34.416 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 40.5600 0.5950 40.7000 ;
    END
  END WW4BEG[1]
  PIN WW4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3929 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6565 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1115 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.852 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.344 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.4794 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 179.968 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 39.2000 0.5950 39.3400 ;
    END
  END WW4BEG[0]
  PIN W6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9669 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 14.6895 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2351 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0045 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 10.012 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.8464 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 32.592 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 78.9800 0.5950 79.1200 ;
    END
  END W6BEG[11]
  PIN W6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3285 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.2605 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.1315 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.6968 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 57.52 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 77.6200 0.5950 77.7600 ;
    END
  END W6BEG[10]
  PIN W6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4097 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.9405 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.1745 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 21.9876 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 118.208 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 75.9200 0.5950 76.0600 ;
    END
  END W6BEG[9]
  PIN W6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2437 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.1105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.3791 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.7245 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.37 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 50.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.4188 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 98.704 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 74.5600 0.5950 74.7000 ;
    END
  END W6BEG[8]
  PIN W6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0401 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.0925 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9785 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.7215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.345 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.64 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.0378 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 64.672 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 73.2000 0.5950 73.3400 ;
    END
  END W6BEG[7]
  PIN W6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1385 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.3567 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.6125 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.874 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.128 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 71.5000 0.5950 71.6400 ;
    END
  END W6BEG[6]
  PIN W6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3093 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.4015 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1075 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4655 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.8108 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 90.128 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 70.1400 0.5950 70.2800 ;
    END
  END W6BEG[5]
  PIN W6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1045 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.4145 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 7.3415 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 36.5365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.473 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.656 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.4266 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 83.216 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 68.7800 0.5950 68.9200 ;
    END
  END W6BEG[4]
  PIN W6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0709 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.2465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.6719 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1885 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.195 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.84 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.3538 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 45.024 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 67.0800 0.5950 67.2200 ;
    END
  END W6BEG[3]
  PIN W6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3929 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.9421 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.5395 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 21.442 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 114.824 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.5828 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.912 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 65.7200 0.5950 65.8600 ;
    END
  END W6BEG[2]
  PIN W6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3317 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5505 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.6445 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.0515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.597 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.984 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.3998 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 7.936 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 64.3600 0.5950 64.5000 ;
    END
  END W6BEG[1]
  PIN W6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9705 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.7075 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2743 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2005 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.096 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 27.2508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 145.808 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 0.0000 62.3200 0.5950 62.4600 ;
    END
  END W6BEG[0]
  PIN RAM2FAB_D0_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3285 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.5265 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.4615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.0316 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.776 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 57.0591 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 279.558 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 45.3200 100.2800 45.4600 ;
    END
  END RAM2FAB_D0_I0
  PIN RAM2FAB_D0_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.0734 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 20.195 LAYER met1  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met1  ;
    ANTENNAMAXAREACAR 18.7028 LAYER met1  ;
    ANTENNAMAXSIDEAREACAR 82.4246 LAYER met1  ;
    ANTENNAMAXCUTCAR 0.229365 LAYER via  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 48.3800 100.2800 48.5200 ;
    END
  END RAM2FAB_D0_I1
  PIN RAM2FAB_D0_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4673 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.2285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2651 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.0515 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.0498 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.736 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 42.2198 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 208.538 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 51.4400 100.2800 51.5800 ;
    END
  END RAM2FAB_D0_I2
  PIN RAM2FAB_D0_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2673 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.2285 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 3.6175 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.9165 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 23.2618 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 125 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.7328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 57.712 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 60.7671 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 308.903 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 54.5000 100.2800 54.6400 ;
    END
  END RAM2FAB_D0_I3
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.2556 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 102.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.6938 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.504 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.608 LAYER met4  ;
    ANTENNAMAXAREACAR 1.54431 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 7.46452 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.0473307 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 80.5800 0.0000 80.8800 0.8000 ;
    END
  END UserCLK
  PIN RAM2FAB_D1_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3317 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5505 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 11.2741 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 56.1995 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.816 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.5868 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 67.6 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 66.2766 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 342.169 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 33.4200 100.2800 33.5600 ;
    END
  END RAM2FAB_D1_I0
  PIN RAM2FAB_D1_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4237 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.6309 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.186 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 70.792 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 14.0321 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 63.4802 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 36.4800 100.2800 36.6200 ;
    END
  END RAM2FAB_D1_I1
  PIN RAM2FAB_D1_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5249 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.5165 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3513 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5855 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 15.898 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 85.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 9.6252 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 53.216 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 54.1913 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 281.772 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 39.5400 100.2800 39.6800 ;
    END
  END RAM2FAB_D1_I2
  PIN RAM2FAB_D1_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2505 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1445 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.2679 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.1685 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 14.0554 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.84 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.2844 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.928 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 75.6417 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 390.28 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 42.6000 100.2800 42.7400 ;
    END
  END RAM2FAB_D1_I3
  PIN RAM2FAB_D2_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2029 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9065 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.3505 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 26.4635 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.32 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.392 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 72.8718 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 367.423 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.745238 LAYER via3  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 21.5200 100.2800 21.6600 ;
    END
  END RAM2FAB_D2_I0
  PIN RAM2FAB_D2_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1385 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 10.292 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.988 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 51.1802 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 243.952 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 24.5800 100.2800 24.7200 ;
    END
  END RAM2FAB_D2_I1
  PIN RAM2FAB_D2_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9757 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.7705 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2225 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.9415 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.8328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 138.712 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 13.5968 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 59.756 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 27.6400 100.2800 27.7800 ;
    END
  END RAM2FAB_D2_I2
  PIN RAM2FAB_D2_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8753 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.2315 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.3059 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 21.1225 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.5218 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.72 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 1.8846 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 10.992 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 88.5984 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 441.405 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.38016 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 30.7000 100.2800 30.8400 ;
    END
  END RAM2FAB_D2_I3
  PIN RAM2FAB_D3_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5533 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 2.6215 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.8448 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.87 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 47.7563 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 227.008 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 9.9600 100.2800 10.1000 ;
    END
  END RAM2FAB_D3_I0
  PIN RAM2FAB_D3_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2129 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.9565 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4402 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.965 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met2  ;
    ANTENNAMAXAREACAR 36.7591 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 170.98 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.586508 LAYER via2  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 12.6800 100.2800 12.8200 ;
    END
  END RAM2FAB_D3_I1
  PIN RAM2FAB_D3_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.1209 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 45.4965 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 4.6197 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 22.8095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 16.4058 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 87.968 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 93.0913 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 484.689 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 15.7400 100.2800 15.8800 ;
    END
  END RAM2FAB_D3_I2
  PIN RAM2FAB_D3_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7181 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 6.5195 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.3085 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.019 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.568 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.9736 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 64.8 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 121.765 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 636.966 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.903968 LAYER via4  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 18.8000 100.2800 18.9400 ;
    END
  END RAM2FAB_D3_I3
  PIN FAB2RAM_D0_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9865 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.8245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.2781 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 15.0396 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 81.152 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 140.5200 100.2800 140.6600 ;
    END
  END FAB2RAM_D0_O0
  PIN FAB2RAM_D0_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2641 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.7321 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4895 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.7808 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 73.968 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 143.5800 100.2800 143.7200 ;
    END
  END FAB2RAM_D0_O1
  PIN FAB2RAM_D0_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3285 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.5345 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4381 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.0195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.61 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 35.72 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.4846 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 206.192 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 146.3000 100.2800 146.4400 ;
    END
  END FAB2RAM_D0_O2
  PIN FAB2RAM_D0_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1961 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.8725 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.5812 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.788 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 149.7000 100.2800 149.8400 ;
    END
  END FAB2RAM_D0_O3
  PIN FAB2RAM_D1_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6537 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.1605 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 9.6246 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 47.887 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 128.6200 100.2800 128.7600 ;
    END
  END FAB2RAM_D1_O0
  PIN FAB2RAM_D1_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.7909 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.813 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 131.6800 100.2800 131.8200 ;
    END
  END FAB2RAM_D1_O1
  PIN FAB2RAM_D1_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9061 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.3855 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.7048 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.288 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 134.7400 100.2800 134.8800 ;
    END
  END FAB2RAM_D1_O2
  PIN FAB2RAM_D1_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2165 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.9745 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1179 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.4935 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.99 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.08 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 8.1708 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 44.048 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 137.8000 100.2800 137.9400 ;
    END
  END FAB2RAM_D1_O3
  PIN FAB2RAM_D2_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2977 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.3805 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.5889 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.7735 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.883 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.3286 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 77.36 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 116.7200 100.2800 116.8600 ;
    END
  END FAB2RAM_D2_O0
  PIN FAB2RAM_D2_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1373 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.572 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2407 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.0325 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.4328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.112 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 119.7800 100.2800 119.9200 ;
    END
  END FAB2RAM_D2_O1
  PIN FAB2RAM_D2_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0349 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 5.0295 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3863 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.7605 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.646 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 51.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.8028 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 20.752 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 122.5000 100.2800 122.6400 ;
    END
  END FAB2RAM_D2_O2
  PIN FAB2RAM_D2_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8437 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1105 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2636 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.2 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 125.9000 100.2800 126.0400 ;
    END
  END FAB2RAM_D2_O3
  PIN FAB2RAM_D3_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9705 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 4.7075 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.2659 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.1585 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.8608 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 111.728 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 104.8200 100.2800 104.9600 ;
    END
  END FAB2RAM_D3_O0
  PIN FAB2RAM_D3_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1385 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 0.5845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.5336 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 32.55 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 107.8800 100.2800 108.0200 ;
    END
  END FAB2RAM_D3_O1
  PIN FAB2RAM_D3_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5385 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5845 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.6724 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 28.126 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 110.9400 100.2800 111.0800 ;
    END
  END FAB2RAM_D3_O2
  PIN FAB2RAM_D3_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2641 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 6.2125 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3471 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.2598 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.856 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 114.0000 100.2800 114.1400 ;
    END
  END FAB2RAM_D3_O3
  PIN FAB2RAM_A0_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 3.3571 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 16.681 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 92.9200 100.2800 93.0600 ;
    END
  END FAB2RAM_A0_O0
  PIN FAB2RAM_A0_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5793 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.7885 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.788 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.822 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 95.9800 100.2800 96.1200 ;
    END
  END FAB2RAM_A0_O1
  PIN FAB2RAM_A0_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8605 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 9.1945 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 5.1323 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.4905 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.2436 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 82.24 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 98.7000 100.2800 98.8400 ;
    END
  END FAB2RAM_A0_O2
  PIN FAB2RAM_A0_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3317 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5505 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 1.4153 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.9055 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.16 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.3148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.816 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 102.1000 100.2800 102.2400 ;
    END
  END FAB2RAM_A0_O3
  PIN FAB2RAM_A1_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7181 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4825 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 2.4891 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.2745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 11.0208 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.248 LAYER met3  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 81.0200 100.2800 81.1600 ;
    END
  END FAB2RAM_A1_O0
  PIN FAB2RAM_A1_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5601 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 22.6555 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.0048 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.788 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 84.0800 100.2800 84.2200 ;
    END
  END FAB2RAM_A1_O1
  PIN FAB2RAM_A1_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5217 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.5005 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.3636 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.464 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 87.1400 100.2800 87.2800 ;
    END
  END FAB2RAM_A1_O2
  PIN FAB2RAM_A1_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4265 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.0245 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.1932 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.73 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 90.2000 100.2800 90.3400 ;
    END
  END FAB2RAM_A1_O3
  PIN FAB2RAM_C_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 1.6981 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 8.386 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 69.1200 100.2800 69.2600 ;
    END
  END FAB2RAM_C_O0
  PIN FAB2RAM_C_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 4.7739 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 23.765 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 72.1800 100.2800 72.3200 ;
    END
  END FAB2RAM_C_O1
  PIN FAB2RAM_C_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3317 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 1.5505 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.4815 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 2.2365 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 11.161 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 59.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.4336 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.92 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 75.2400 100.2800 75.3800 ;
    END
  END FAB2RAM_C_O2
  PIN FAB2RAM_C_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7055 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 3.4195 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.8672 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 44.1 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 78.3000 100.2800 78.4400 ;
    END
  END FAB2RAM_C_O3
  PIN Config_accessC_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5465 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 17.5875 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.3709 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6835 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 13.003 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 69.816 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 5.2428 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 28.432 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 57.2200 100.2800 57.3600 ;
    END
  END Config_accessC_bit0
  PIN Config_accessC_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2077 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 15.8935 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNAPARTIALMETALAREA 0.1917 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7875 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 9.094 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 1.7658 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 9.888 LAYER met4  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 60.2800 100.2800 60.4200 ;
    END
  END Config_accessC_bit1
  PIN Config_accessC_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met1  ;
    ANTENNAPARTIALMETALAREA 2.7712 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 13.7515 LAYER met1  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 63.3400 100.2800 63.4800 ;
    END
  END Config_accessC_bit2
  PIN Config_accessC_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4909 LAYER met1  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3465 LAYER met1  ;
    ANTENNAPARTIALCUTAREA 0.0225 LAYER via  ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 7.9622 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.221 LAYER met2  ;
    PORT
      LAYER met1 ;
        RECT 99.6850 66.0600 100.2800 66.2000 ;
    END
  END Config_accessC_bit3
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.7746 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 89.456 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.1008 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 97.008 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1735 LAYER met4  ;
    ANTENNAMAXAREACAR 43.4302 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 216.31 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.667808 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 209.3500 0.8000 209.6500 ;
    END
  END FrameData[31]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.4686 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.824 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.1794 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 98.368 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1735 LAYER met4  ;
    ANTENNAMAXAREACAR 27.679 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 138.253 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.593246 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 207.5200 0.8000 207.8200 ;
    END
  END FrameData[30]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.575 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 105.336 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1735 LAYER met3  ;
    ANTENNAMAXAREACAR 46.9277 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 232.832 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.706918 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 205.6900 0.8000 205.9900 ;
    END
  END FrameData[29]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2386 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.0342 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 146.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1735 LAYER met4  ;
    ANTENNAMAXAREACAR 45.8895 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 230.574 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.80021 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 203.8600 0.8000 204.1600 ;
    END
  END FrameData[28]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9406 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 23.5026 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 126.288 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1735 LAYER met4  ;
    ANTENNAMAXAREACAR 31.7689 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 159.892 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.590566 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 202.0300 0.8000 202.3300 ;
    END
  END FrameData[27]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.2577 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 87.64 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met3  ;
    ANTENNAMAXAREACAR 57.4138 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 302.552 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.700629 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.8017 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 31.408 LAYER met4  ;
    ANTENNAGATEAREA 2.1735 LAYER met4  ;
    ANTENNAMAXAREACAR 60.0831 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 317.002 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.849993 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 200.2000 0.8000 200.5000 ;
    END
  END FrameData[26]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.284 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.816 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.8555 LAYER met3  ;
    ANTENNAMAXAREACAR 26.3247 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 127.398 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.649404 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.8508 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 5.008 LAYER met4  ;
    ANTENNAGATEAREA 2.1735 LAYER met4  ;
    ANTENNAMAXAREACAR 26.7161 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 129.702 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 198.3700 0.8000 198.6700 ;
    END
  END FrameData[25]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.8802 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.96 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.954 LAYER met3  ;
    ANTENNAMAXAREACAR 35.7866 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 177.129 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.868344 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.6478 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 62.592 LAYER met4  ;
    ANTENNAGATEAREA 2.1735 LAYER met4  ;
    ANTENNAMAXAREACAR 41.1456 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 205.927 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.868344 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 196.5400 0.8000 196.8400 ;
    END
  END FrameData[24]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3642 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.408 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1735 LAYER met3  ;
    ANTENNAMAXAREACAR 28.8453 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 140.015 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.511936 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 195.3200 0.8000 195.6200 ;
    END
  END FrameData[23]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3596 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.5576 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 41.248 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1735 LAYER met4  ;
    ANTENNAMAXAREACAR 38.0116 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 192.57 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.574843 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 193.4900 0.8000 193.7900 ;
    END
  END FrameData[22]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4456 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.7952 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.456 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1735 LAYER met4  ;
    ANTENNAMAXAREACAR 30.1711 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 150.89 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 191.6600 0.8000 191.9600 ;
    END
  END FrameData[21]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.9662 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 80.752 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.636 LAYER met3  ;
    ANTENNAMAXAREACAR 44.0204 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 223.009 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.779245 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.0468 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.72 LAYER met4  ;
    ANTENNAGATEAREA 2.1735 LAYER met4  ;
    ANTENNAMAXAREACAR 45.4222 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 230.702 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.779245 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 189.8300 0.8000 190.1300 ;
    END
  END FrameData[20]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1716 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.24 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 24.9426 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 133.968 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1735 LAYER met4  ;
    ANTENNAMAXAREACAR 35.9566 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 179.886 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.25921 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 188.0000 0.8000 188.3000 ;
    END
  END FrameData[19]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.9224 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.048 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.2511 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 147.216 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1735 LAYER met4  ;
    ANTENNAMAXAREACAR 61.609 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 325.597 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.2195 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 186.1700 0.8000 186.4700 ;
    END
  END FrameData[18]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4456 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.3884 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 104.816 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1735 LAYER met4  ;
    ANTENNAMAXAREACAR 30.0334 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 150.068 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.632495 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 184.3400 0.8000 184.6400 ;
    END
  END FrameData[17]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8626 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.8464 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 32.592 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1735 LAYER met4  ;
    ANTENNAMAXAREACAR 33.7226 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 177.388 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 182.5100 0.8000 182.8100 ;
    END
  END FrameData[16]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.4664 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 61.616 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5375 LAYER met3  ;
    ANTENNAMAXAREACAR 27.4294 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 135.096 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.472074 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAGATEAREA 2.1735 LAYER met4  ;
    ANTENNAMAXAREACAR 27.7367 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 136.951 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.590566 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 181.2900 0.8000 181.5900 ;
    END
  END FrameData[15]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.735 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.656 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9015 LAYER met3  ;
    ANTENNAMAXAREACAR 10.0291 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 47.6628 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.870786 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.4778 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 72.352 LAYER met4  ;
    ANTENNAGATEAREA 2.1735 LAYER met4  ;
    ANTENNAMAXAREACAR 34.122 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 169.801 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.870786 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 179.4600 0.8000 179.7600 ;
    END
  END FrameData[14]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4456 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 43.4742 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 235.616 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1735 LAYER met4  ;
    ANTENNAMAXAREACAR 75.7529 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 395.762 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.47107 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 177.6300 0.8000 177.9300 ;
    END
  END FrameData[13]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.2859 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.968 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.477 LAYER met3  ;
    ANTENNAMAXAREACAR 45.9524 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 229.057 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.857862 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.6524 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 58.224 LAYER met4  ;
    ANTENNAGATEAREA 2.1735 LAYER met4  ;
    ANTENNAMAXAREACAR 103.257 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 521.996 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 175.8000 0.8000 176.1000 ;
    END
  END FrameData[12]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1261 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.6 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3785 LAYER met3  ;
    ANTENNAMAXAREACAR 40.8842 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 202.602 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.619583 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.5238 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 35.264 LAYER met4  ;
    ANTENNAGATEAREA 2.1735 LAYER met4  ;
    ANTENNAMAXAREACAR 43.8857 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 218.827 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.619583 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 173.9700 0.8000 174.2700 ;
    END
  END FrameData[11]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.608 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1735 LAYER met3  ;
    ANTENNAMAXAREACAR 34.9967 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 170.081 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.483183 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 172.1400 0.8000 172.4400 ;
    END
  END FrameData[10]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.0456 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 37.568 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.8126 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 26.608 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1735 LAYER met4  ;
    ANTENNAMAXAREACAR 37.3914 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 184.961 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.568845 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 170.3100 0.8000 170.6100 ;
    END
  END FrameData[9]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.8976 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.112 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 21.9582 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 118.992 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.1735 LAYER met4  ;
    ANTENNAMAXAREACAR 31.4915 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 158.289 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04597 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 168.4800 0.8000 168.7800 ;
    END
  END FrameData[8]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4916 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 21.48 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 116.912 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.0145 LAYER met4  ;
    ANTENNAMAXAREACAR 53.1113 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 277.584 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.993373 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 167.2600 0.8000 167.5600 ;
    END
  END FrameData[7]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2386 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 11.2818 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 60.64 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.0145 LAYER met4  ;
    ANTENNAMAXAREACAR 35.3495 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 177.096 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.504492 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 165.4300 0.8000 165.7300 ;
    END
  END FrameData[6]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.5933 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 88.488 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.0145 LAYER met3  ;
    ANTENNAMAXAREACAR 33.0275 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 162.005 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.629867 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 163.6000 0.8000 163.9000 ;
    END
  END FrameData[5]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.3713 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.104 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.477 LAYER met3  ;
    ANTENNAMAXAREACAR 53.9455 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 270.284 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.941719 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 33.1134 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 178.016 LAYER met4  ;
    ANTENNAGATEAREA 2.0145 LAYER met4  ;
    ANTENNAMAXAREACAR 70.383 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 358.651 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.941719 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 161.7700 0.8000 162.0700 ;
    END
  END FrameData[4]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8206 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 14.8776 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 80.288 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.0145 LAYER met4  ;
    ANTENNAMAXAREACAR 24.5048 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 124.148 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 159.9400 0.8000 160.2400 ;
    END
  END FrameData[3]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7034 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 20.7372 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 112 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.0145 LAYER met4  ;
    ANTENNAMAXAREACAR 39.8581 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 208.001 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 158.1100 0.8000 158.4100 ;
    END
  END FrameData[2]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7988 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.0145 LAYER met3  ;
    ANTENNAMAXAREACAR 42.1806 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 208.071 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.716352 LAYER via3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 156.2800 0.8000 156.5800 ;
    END
  END FrameData[1]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.886 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.712 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.636 LAYER met3  ;
    ANTENNAMAXAREACAR 35.369 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 175.991 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.449057 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 13.1118 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 70.4 LAYER met4  ;
    ANTENNAGATEAREA 2.0145 LAYER met4  ;
    ANTENNAMAXAREACAR 41.8777 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 210.938 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.449057 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 155.0600 0.8000 155.3600 ;
    END
  END FrameData[0]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 1.4064 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.496 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 99.4800 209.3500 100.2800 209.6500 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7916 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.88 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.7758 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 164.608 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.4800 207.5200 100.2800 207.8200 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6976 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.712 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.9348 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 165.456 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.4800 205.6900 100.2800 205.9900 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0076 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.032 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 30.8628 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 165.072 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.4800 203.8600 100.2800 204.1600 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4126 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.192 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 22.4994 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 121.408 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.4800 202.0300 100.2800 202.3300 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.0099 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.048 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 99.4800 200.2000 100.2800 200.5000 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3076 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.0906 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 177.424 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.4800 198.3700 100.2800 198.6700 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.0696 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 69.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.6856 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 127.264 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.4800 196.5400 100.2800 196.8400 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1816 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 26.8992 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 145.344 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.4800 195.3200 100.2800 195.6200 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.6876 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.992 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 23.9088 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 127.984 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.4800 193.4900 100.2800 193.7900 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.5156 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 45.408 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 50.3394 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 269.888 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.4800 191.6600 100.2800 191.9600 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.2576 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 92.032 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.9504 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 118.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.4800 189.8300 100.2800 190.1300 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.2896 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.8244 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 69.808 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.4800 188.0000 100.2800 188.3000 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3426 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.152 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.3528 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 84.704 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.4800 186.1700 100.2800 186.4700 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.1194 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 64.632 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 99.4800 184.3400 100.2800 184.6400 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.344 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 99.4800 182.5100 100.2800 182.8100 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 24.8926 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 132.752 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.2358 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 97.728 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.4800 181.2900 100.2800 181.5900 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.2546 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 60.016 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 7.9236 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 43.2 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.4800 179.4600 100.2800 179.7600 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3776 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 12.672 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.5158 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 253.888 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.4800 177.6300 100.2800 177.9300 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.2636 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 76.064 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 14.2098 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 76.256 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.4800 175.8000 100.2800 176.1000 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.2866 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.52 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 19.2294 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 103.968 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.4800 173.9700 100.2800 174.2700 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3076 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 31.1178 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 166.432 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.4800 172.1400 100.2800 172.4400 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.608 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 99.4800 170.3100 100.2800 170.6100 ;
    END
  END FrameData_O[9]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.344 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 99.4800 168.4800 100.2800 168.7800 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.344 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 99.4800 167.2600 100.2800 167.5600 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.0099 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.048 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 99.4800 165.4300 100.2800 165.7300 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.608 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 99.4800 163.6000 100.2800 163.9000 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4404 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.344 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 99.4800 161.7700 100.2800 162.0700 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6826 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 16.0398 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 86.016 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.4800 159.9400 100.2800 160.2400 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.7356 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.248 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 43.5138 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 232.544 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.4800 157.5000 100.2800 157.8000 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.8006 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.928 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 4.1352 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 23.936 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.4800 156.2800 100.2800 156.5800 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.7816 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 52.16 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 15.4506 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 83.344 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 99.4800 155.0600 100.2800 155.3600 ;
    END
  END FrameData_O[0]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.0246 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.962 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.195 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.84 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 42.2952 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 227.456 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 70.4791 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 376.718 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 97.2200 0.0000 97.3600 0.4850 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0663 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.2235 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 5.45603 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 25.899 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 96.7600 0.0000 96.9000 0.4850 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0724 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.201 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 30.2988 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 162.064 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 54.2321 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 284.657 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 95.8400 0.0000 95.9800 0.4850 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9206 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 24.206 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 27.1866 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 145.936 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 41.0859 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 218.39 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 94.9200 0.0000 95.0600 0.4850 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4423 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.9855 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 7.56943 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 36.3071 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 94.4600 0.0000 94.6000 0.4850 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3038 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.358 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.6268 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 46.48 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 19.6314 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 101.197 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 92.6200 0.0000 92.7600 0.4850 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.0121 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 54.3095 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.8898 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.216 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 7.96835 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 40.7556 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 92.1600 0.0000 92.3000 0.4850 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1067 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.3075 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 4.05859 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 18.7529 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 91.2400 0.0000 91.3800 0.4850 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1539 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.5435 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 6.05347 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 28.7273 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 90.3200 0.0000 90.4600 0.4850 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.4723 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.1355 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met2  ;
    ANTENNAMAXAREACAR 9.39084 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 45.4141 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0692256 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 89.4000 0.0000 89.5400 0.4850 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 27.1052 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 135.247 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.08 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.56 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.5108 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 24.528 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met4  ;
    ANTENNAMAXAREACAR 9.1468 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 47.7037 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.17697 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 88.9400 0.0000 89.0800 0.4850 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.2148 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.333 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.477 LAYER met2  ;
    ANTENNAMAXAREACAR 19.2822 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 85.6499 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.730398 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAGATEAREA 0.477 LAYER met3  ;
    ANTENNAMAXAREACAR 19.8314 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 89.5577 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.814256 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 23.1162 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 124.688 LAYER met4  ;
    ANTENNAGATEAREA 4.0125 LAYER met4  ;
    ANTENNAMAXAREACAR 36.5846 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 185.117 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 88.0200 0.0000 88.1600 0.4850 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.0862 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 215.915 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.293 LAYER met2  ;
    ANTENNAMAXAREACAR 35.4159 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 170.364 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.655858 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.228 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.016 LAYER met3  ;
    ANTENNAGATEAREA 4.293 LAYER met3  ;
    ANTENNAMAXAREACAR 35.7019 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 171.998 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.665176 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.6938 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 25.504 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 36.5901 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 176.824 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.665176 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 87.1000 0.0000 87.2400 0.4850 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2222 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.95 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.714 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 41.608 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 10.8288 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 58.224 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 26.5082 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 123.637 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.772009 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 86.6400 0.0000 86.7800 0.4850 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.5288 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.247 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.4508 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.208 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met3  ;
    ANTENNAMAXAREACAR 20.377 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 96.2918 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.472349 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 85.7200 0.0000 85.8600 0.4850 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.9722 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 162.204 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.021 LAYER met2  ;
    ANTENNAMAXAREACAR 27.003 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 129.395 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.61953 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 5.9325 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.576 LAYER met3  ;
    ANTENNAGATEAREA 5.2845 LAYER met3  ;
    ANTENNAMAXAREACAR 28.1256 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 135.559 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 84.8000 0.0000 84.9400 0.4850 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.7334 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 52.71 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.636 LAYER met2  ;
    ANTENNAMAXAREACAR 21.8676 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 103.274 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.527673 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 8.9164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 48.016 LAYER met3  ;
    ANTENNAGATEAREA 0.954 LAYER met3  ;
    ANTENNAMAXAREACAR 31.2139 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 153.605 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.569602 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.4336 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.92 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 32.0456 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 156.239 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.86457 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 84.3400 0.0000 84.4800 0.4850 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 43.611 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 213.703 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.6485 LAYER met2  ;
    ANTENNAMAXAREACAR 30.5534 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 146.847 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.80526 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.2495 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.6 LAYER met3  ;
    ANTENNAGATEAREA 5.2845 LAYER met3  ;
    ANTENNAMAXAREACAR 31.3576 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 151.313 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.80526 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 83.4200 0.0000 83.5600 0.4850 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.1882 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 39.984 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.272 LAYER met2  ;
    ANTENNAMAXAREACAR 14.3542 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 61.6195 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.496226 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAGATEAREA 1.272 LAYER met3  ;
    ANTENNAMAXAREACAR 14.4524 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 62.5126 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.527673 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.8472 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 86.4 LAYER met4  ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 42.0016 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 217.796 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.07799 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 82.5000 0.0000 82.6400 0.4850 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5862 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.77 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.331 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 12.5565 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 67.904 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.2845 LAYER met4  ;
    ANTENNAMAXAREACAR 36.6195 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 180.622 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.705547 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 82.0400 0.0000 82.1800 0.4850 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.0619 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.0835 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 97.6800 219.1550 97.8200 219.6400 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8773 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.2785 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 96.7600 219.1550 96.9000 219.6400 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.3991 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.8875 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 95.8400 219.1550 95.9800 219.6400 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2327 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.9375 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 94.9200 219.1550 95.0600 219.6400 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.063 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.154 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.056 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.432 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.8728 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 319.792 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 94.0000 219.1550 94.1400 219.6400 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.6502 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 27.972 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.469 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.968 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 17.1378 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 91.872 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 93.5400 219.1550 93.6800 219.6400 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.2871 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.3275 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 92.6200 219.1550 92.7600 219.6400 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3268 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.473 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.952 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 5.544 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 55.4088 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 295.984 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 91.7000 219.1550 91.8400 219.6400 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8043 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.7955 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 90.7800 219.1550 90.9200 219.6400 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.7967 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.8755 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 89.8600 219.1550 90.0000 219.6400 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5187 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.3675 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 89.4000 219.1550 89.5400 219.6400 ;
    END
  END FrameStrobe_O[9]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.3971 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8775 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 88.4800 219.1550 88.6200 219.6400 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.633 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.768 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.745 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 3.4128 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.672 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 87.5600 219.1550 87.7000 219.6400 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.198 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.829 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.507 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.504 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 24.0276 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 129.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 86.6400 219.1550 86.7800 219.6400 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3192 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.435 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.498 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 88.456 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 20.1378 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 107.872 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 85.7200 219.1550 85.8600 219.6400 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.203 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.854 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 16.753 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 89.816 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 85.2600 219.1550 85.4000 219.6400 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 5.1543 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 25.4275 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 83.8800 219.1550 84.0200 219.6400 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 6.2435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 30.8735 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 83.4200 219.1550 83.5600 219.6400 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.7751 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 23.6495 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 82.9600 219.1550 83.1000 219.6400 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7054 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.248 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.918 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 10.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 57.5886 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 308.08 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 82.0400 219.1550 82.1800 219.6400 ;
    END
  END FrameStrobe_O[0]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 5.5600 5.4300 94.7200 6.9300 ;
        RECT 5.5600 212.0300 94.7200 213.5300 ;
        RECT 5.5600 12.3400 7.0600 12.8200 ;
        RECT 5.5600 17.7800 7.0600 18.2600 ;
        RECT 5.5600 23.2200 7.0600 23.7000 ;
        RECT 5.5600 28.6600 7.0600 29.1400 ;
        RECT 5.5600 34.1000 7.0600 34.5800 ;
        RECT 5.5600 39.5400 7.0600 40.0200 ;
        RECT 5.5600 44.9800 7.0600 45.4600 ;
        RECT 5.5600 50.4200 7.0600 50.9000 ;
        RECT 5.5600 55.8600 7.0600 56.3400 ;
        RECT 5.5600 61.3000 7.0600 61.7800 ;
        RECT 5.5600 66.7400 7.0600 67.2200 ;
        RECT 5.5600 72.1800 7.0600 72.6600 ;
        RECT 5.5600 77.6200 7.0600 78.1000 ;
        RECT 5.5600 83.0600 7.0600 83.5400 ;
        RECT 5.5600 88.5000 7.0600 88.9800 ;
        RECT 5.5600 93.9400 7.0600 94.4200 ;
        RECT 5.5600 99.3800 7.0600 99.8600 ;
        RECT 5.5600 104.8200 7.0600 105.3000 ;
        RECT 93.2200 12.3400 94.7200 12.8200 ;
        RECT 93.2200 17.7800 94.7200 18.2600 ;
        RECT 93.2200 23.2200 94.7200 23.7000 ;
        RECT 93.2200 28.6600 94.7200 29.1400 ;
        RECT 93.2200 34.1000 94.7200 34.5800 ;
        RECT 93.2200 39.5400 94.7200 40.0200 ;
        RECT 93.2200 44.9800 94.7200 45.4600 ;
        RECT 93.2200 50.4200 94.7200 50.9000 ;
        RECT 93.2200 55.8600 94.7200 56.3400 ;
        RECT 93.2200 61.3000 94.7200 61.7800 ;
        RECT 93.2200 66.7400 94.7200 67.2200 ;
        RECT 93.2200 72.1800 94.7200 72.6600 ;
        RECT 93.2200 77.6200 94.7200 78.1000 ;
        RECT 93.2200 83.0600 94.7200 83.5400 ;
        RECT 93.2200 88.5000 94.7200 88.9800 ;
        RECT 93.2200 93.9400 94.7200 94.4200 ;
        RECT 93.2200 99.3800 94.7200 99.8600 ;
        RECT 93.2200 104.8200 94.7200 105.3000 ;
        RECT 5.5600 164.6600 7.0600 165.1400 ;
        RECT 5.5600 110.2600 7.0600 110.7400 ;
        RECT 5.5600 115.7000 7.0600 116.1800 ;
        RECT 5.5600 121.1400 7.0600 121.6200 ;
        RECT 5.5600 126.5800 7.0600 127.0600 ;
        RECT 5.5600 132.0200 7.0600 132.5000 ;
        RECT 5.5600 137.4600 7.0600 137.9400 ;
        RECT 5.5600 142.9000 7.0600 143.3800 ;
        RECT 5.5600 148.3400 7.0600 148.8200 ;
        RECT 5.5600 153.7800 7.0600 154.2600 ;
        RECT 5.5600 159.2200 7.0600 159.7000 ;
        RECT 5.5600 191.8600 7.0600 192.3400 ;
        RECT 5.5600 170.1000 7.0600 170.5800 ;
        RECT 5.5600 175.5400 7.0600 176.0200 ;
        RECT 5.5600 180.9800 7.0600 181.4600 ;
        RECT 5.5600 186.4200 7.0600 186.9000 ;
        RECT 5.5600 197.3000 7.0600 197.7800 ;
        RECT 5.5600 202.7400 7.0600 203.2200 ;
        RECT 5.5600 208.1800 7.0600 208.6600 ;
        RECT 93.2200 164.6600 94.7200 165.1400 ;
        RECT 93.2200 110.2600 94.7200 110.7400 ;
        RECT 93.2200 115.7000 94.7200 116.1800 ;
        RECT 93.2200 121.1400 94.7200 121.6200 ;
        RECT 93.2200 126.5800 94.7200 127.0600 ;
        RECT 93.2200 132.0200 94.7200 132.5000 ;
        RECT 93.2200 137.4600 94.7200 137.9400 ;
        RECT 93.2200 142.9000 94.7200 143.3800 ;
        RECT 93.2200 148.3400 94.7200 148.8200 ;
        RECT 93.2200 153.7800 94.7200 154.2600 ;
        RECT 93.2200 159.2200 94.7200 159.7000 ;
        RECT 93.2200 191.8600 94.7200 192.3400 ;
        RECT 93.2200 170.1000 94.7200 170.5800 ;
        RECT 93.2200 175.5400 94.7200 176.0200 ;
        RECT 93.2200 180.9800 94.7200 181.4600 ;
        RECT 93.2200 186.4200 94.7200 186.9000 ;
        RECT 93.2200 197.3000 94.7200 197.7800 ;
        RECT 93.2200 202.7400 94.7200 203.2200 ;
        RECT 93.2200 208.1800 94.7200 208.6600 ;
      LAYER met4 ;
        RECT 93.2200 5.4300 94.7200 213.5300 ;
        RECT 5.5600 5.4300 7.0600 213.5300 ;
    END
# end of P/G power stripe data as pin

  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 3.0600 2.9300 97.2200 4.4300 ;
        RECT 3.0600 214.5300 97.2200 216.0300 ;
        RECT 3.0600 9.6200 4.5600 10.1000 ;
        RECT 3.0600 15.0600 4.5600 15.5400 ;
        RECT 3.0600 20.5000 4.5600 20.9800 ;
        RECT 3.0600 25.9400 4.5600 26.4200 ;
        RECT 3.0600 31.3800 4.5600 31.8600 ;
        RECT 3.0600 36.8200 4.5600 37.3000 ;
        RECT 3.0600 42.2600 4.5600 42.7400 ;
        RECT 3.0600 47.7000 4.5600 48.1800 ;
        RECT 3.0600 53.1400 4.5600 53.6200 ;
        RECT 3.0600 58.5800 4.5600 59.0600 ;
        RECT 3.0600 64.0200 4.5600 64.5000 ;
        RECT 3.0600 69.4600 4.5600 69.9400 ;
        RECT 3.0600 74.9000 4.5600 75.3800 ;
        RECT 3.0600 80.3400 4.5600 80.8200 ;
        RECT 3.0600 85.7800 4.5600 86.2600 ;
        RECT 3.0600 91.2200 4.5600 91.7000 ;
        RECT 3.0600 96.6600 4.5600 97.1400 ;
        RECT 3.0600 102.1000 4.5600 102.5800 ;
        RECT 3.0600 107.5400 4.5600 108.0200 ;
        RECT 95.7200 9.6200 97.2200 10.1000 ;
        RECT 95.7200 15.0600 97.2200 15.5400 ;
        RECT 95.7200 20.5000 97.2200 20.9800 ;
        RECT 95.7200 25.9400 97.2200 26.4200 ;
        RECT 95.7200 31.3800 97.2200 31.8600 ;
        RECT 95.7200 36.8200 97.2200 37.3000 ;
        RECT 95.7200 42.2600 97.2200 42.7400 ;
        RECT 95.7200 47.7000 97.2200 48.1800 ;
        RECT 95.7200 53.1400 97.2200 53.6200 ;
        RECT 95.7200 58.5800 97.2200 59.0600 ;
        RECT 95.7200 64.0200 97.2200 64.5000 ;
        RECT 95.7200 69.4600 97.2200 69.9400 ;
        RECT 95.7200 74.9000 97.2200 75.3800 ;
        RECT 95.7200 80.3400 97.2200 80.8200 ;
        RECT 95.7200 85.7800 97.2200 86.2600 ;
        RECT 95.7200 91.2200 97.2200 91.7000 ;
        RECT 95.7200 96.6600 97.2200 97.1400 ;
        RECT 95.7200 102.1000 97.2200 102.5800 ;
        RECT 95.7200 107.5400 97.2200 108.0200 ;
        RECT 3.0600 112.9800 4.5600 113.4600 ;
        RECT 3.0600 118.4200 4.5600 118.9000 ;
        RECT 3.0600 123.8600 4.5600 124.3400 ;
        RECT 3.0600 129.3000 4.5600 129.7800 ;
        RECT 3.0600 134.7400 4.5600 135.2200 ;
        RECT 3.0600 140.1800 4.5600 140.6600 ;
        RECT 3.0600 145.6200 4.5600 146.1000 ;
        RECT 3.0600 151.0600 4.5600 151.5400 ;
        RECT 3.0600 156.5000 4.5600 156.9800 ;
        RECT 3.0600 161.9400 4.5600 162.4200 ;
        RECT 3.0600 178.2600 4.5600 178.7400 ;
        RECT 3.0600 167.3800 4.5600 167.8600 ;
        RECT 3.0600 172.8200 4.5600 173.3000 ;
        RECT 3.0600 183.7000 4.5600 184.1800 ;
        RECT 3.0600 189.1400 4.5600 189.6200 ;
        RECT 3.0600 205.4600 4.5600 205.9400 ;
        RECT 3.0600 194.5800 4.5600 195.0600 ;
        RECT 3.0600 200.0200 4.5600 200.5000 ;
        RECT 95.7200 112.9800 97.2200 113.4600 ;
        RECT 95.7200 118.4200 97.2200 118.9000 ;
        RECT 95.7200 123.8600 97.2200 124.3400 ;
        RECT 95.7200 129.3000 97.2200 129.7800 ;
        RECT 95.7200 134.7400 97.2200 135.2200 ;
        RECT 95.7200 140.1800 97.2200 140.6600 ;
        RECT 95.7200 145.6200 97.2200 146.1000 ;
        RECT 95.7200 151.0600 97.2200 151.5400 ;
        RECT 95.7200 156.5000 97.2200 156.9800 ;
        RECT 95.7200 161.9400 97.2200 162.4200 ;
        RECT 95.7200 178.2600 97.2200 178.7400 ;
        RECT 95.7200 167.3800 97.2200 167.8600 ;
        RECT 95.7200 172.8200 97.2200 173.3000 ;
        RECT 95.7200 183.7000 97.2200 184.1800 ;
        RECT 95.7200 189.1400 97.2200 189.6200 ;
        RECT 95.7200 205.4600 97.2200 205.9400 ;
        RECT 95.7200 194.5800 97.2200 195.0600 ;
        RECT 95.7200 200.0200 97.2200 200.5000 ;
      LAYER met4 ;
        RECT 95.7200 2.9300 97.2200 216.0300 ;
        RECT 3.0600 2.9300 4.5600 216.0300 ;
    END
# end of P/G power stripe data as pin

  END VPWR
  OBS
    LAYER li1 ;
      RECT 79.6050 219.1400 100.2800 219.6400 ;
      RECT 78.6850 219.1400 79.0950 219.6400 ;
      RECT 77.7650 219.1400 78.1750 219.6400 ;
      RECT 76.8450 219.1400 77.2550 219.6400 ;
      RECT 75.4650 219.1400 76.3350 219.6400 ;
      RECT 74.5450 219.1400 74.9550 219.6400 ;
      RECT 73.6250 219.1400 74.0350 219.6400 ;
      RECT 72.7050 219.1400 73.1150 219.6400 ;
      RECT 71.3250 219.1400 72.1950 219.6400 ;
      RECT 70.4050 219.1400 70.8150 219.6400 ;
      RECT 69.4850 219.1400 69.8950 219.6400 ;
      RECT 68.1050 219.1400 68.9750 219.6400 ;
      RECT 67.1850 219.1400 67.5950 219.6400 ;
      RECT 66.2650 219.1400 66.6750 219.6400 ;
      RECT 65.3450 219.1400 65.7550 219.6400 ;
      RECT 63.9650 219.1400 64.8350 219.6400 ;
      RECT 63.0450 219.1400 63.4550 219.6400 ;
      RECT 62.1250 219.1400 62.5350 219.6400 ;
      RECT 60.7450 219.1400 61.6150 219.6400 ;
      RECT 59.8250 219.1400 60.2350 219.6400 ;
      RECT 58.9050 219.1400 59.3150 219.6400 ;
      RECT 57.9850 219.1400 58.3950 219.6400 ;
      RECT 56.6050 219.1400 57.4750 219.6400 ;
      RECT 55.6850 219.1400 56.0950 219.6400 ;
      RECT 54.7650 219.1400 55.1750 219.6400 ;
      RECT 53.3850 219.1400 54.2550 219.6400 ;
      RECT 52.4650 219.1400 52.8750 219.6400 ;
      RECT 51.5450 219.1400 51.9550 219.6400 ;
      RECT 50.6250 219.1400 51.0350 219.6400 ;
      RECT 49.2450 219.1400 50.1150 219.6400 ;
      RECT 48.3250 219.1400 48.7350 219.6400 ;
      RECT 47.4050 219.1400 47.8150 219.6400 ;
      RECT 46.0250 219.1400 46.8950 219.6400 ;
      RECT 45.1050 219.1400 45.5150 219.6400 ;
      RECT 44.1850 219.1400 44.5950 219.6400 ;
      RECT 43.2650 219.1400 43.6750 219.6400 ;
      RECT 41.8850 219.1400 42.7550 219.6400 ;
      RECT 40.9650 219.1400 41.3750 219.6400 ;
      RECT 40.0450 219.1400 40.4550 219.6400 ;
      RECT 39.1250 219.1400 39.5350 219.6400 ;
      RECT 37.7450 219.1400 38.6150 219.6400 ;
      RECT 36.8250 219.1400 37.2350 219.6400 ;
      RECT 35.9050 219.1400 36.3150 219.6400 ;
      RECT 34.5250 219.1400 35.3950 219.6400 ;
      RECT 33.6050 219.1400 34.0150 219.6400 ;
      RECT 32.6850 219.1400 33.0950 219.6400 ;
      RECT 31.7650 219.1400 32.1750 219.6400 ;
      RECT 30.3850 219.1400 31.2550 219.6400 ;
      RECT 29.4650 219.1400 29.8750 219.6400 ;
      RECT 28.5450 219.1400 28.9550 219.6400 ;
      RECT 27.1650 219.1400 28.0350 219.6400 ;
      RECT 26.2450 219.1400 26.6550 219.6400 ;
      RECT 25.3250 219.1400 25.7350 219.6400 ;
      RECT 24.4050 219.1400 24.8150 219.6400 ;
      RECT 23.0250 219.1400 23.8950 219.6400 ;
      RECT 22.1050 219.1400 22.5150 219.6400 ;
      RECT 21.1850 219.1400 21.5950 219.6400 ;
      RECT 19.8050 219.1400 20.6750 219.6400 ;
      RECT 18.8850 219.1400 19.2950 219.6400 ;
      RECT 17.9650 219.1400 18.3750 219.6400 ;
      RECT 17.0450 219.1400 17.4550 219.6400 ;
      RECT 15.6650 219.1400 16.5350 219.6400 ;
      RECT 14.7450 219.1400 15.1550 219.6400 ;
      RECT 13.8250 219.1400 14.2350 219.6400 ;
      RECT 12.4450 219.1400 13.3150 219.6400 ;
      RECT 11.5250 219.1400 11.9350 219.6400 ;
      RECT 10.6050 219.1400 11.0150 219.6400 ;
      RECT 9.6850 219.1400 10.0950 219.6400 ;
      RECT 8.3050 219.1400 9.1750 219.6400 ;
      RECT 7.3850 219.1400 7.7950 219.6400 ;
      RECT 6.4650 219.1400 6.8750 219.6400 ;
      RECT 5.5450 219.1400 5.9550 219.6400 ;
      RECT 0.0000 219.1400 5.0350 219.6400 ;
      RECT 0.0000 0.5000 100.2800 219.1400 ;
      RECT 79.6050 0.0000 100.2800 0.5000 ;
      RECT 78.6850 0.0000 79.0950 0.5000 ;
      RECT 77.7650 0.0000 78.1750 0.5000 ;
      RECT 76.8450 0.0000 77.2550 0.5000 ;
      RECT 75.4650 0.0000 76.3350 0.5000 ;
      RECT 74.5450 0.0000 74.9550 0.5000 ;
      RECT 73.6250 0.0000 74.0350 0.5000 ;
      RECT 72.7050 0.0000 73.1150 0.5000 ;
      RECT 71.3250 0.0000 72.1950 0.5000 ;
      RECT 70.4050 0.0000 70.8150 0.5000 ;
      RECT 69.4850 0.0000 69.8950 0.5000 ;
      RECT 68.1050 0.0000 68.9750 0.5000 ;
      RECT 67.1850 0.0000 67.5950 0.5000 ;
      RECT 66.2650 0.0000 66.6750 0.5000 ;
      RECT 65.3450 0.0000 65.7550 0.5000 ;
      RECT 63.9650 0.0000 64.8350 0.5000 ;
      RECT 63.0450 0.0000 63.4550 0.5000 ;
      RECT 62.1250 0.0000 62.5350 0.5000 ;
      RECT 60.7450 0.0000 61.6150 0.5000 ;
      RECT 59.8250 0.0000 60.2350 0.5000 ;
      RECT 58.9050 0.0000 59.3150 0.5000 ;
      RECT 57.9850 0.0000 58.3950 0.5000 ;
      RECT 56.6050 0.0000 57.4750 0.5000 ;
      RECT 55.6850 0.0000 56.0950 0.5000 ;
      RECT 54.7650 0.0000 55.1750 0.5000 ;
      RECT 53.3850 0.0000 54.2550 0.5000 ;
      RECT 52.4650 0.0000 52.8750 0.5000 ;
      RECT 51.5450 0.0000 51.9550 0.5000 ;
      RECT 50.6250 0.0000 51.0350 0.5000 ;
      RECT 49.2450 0.0000 50.1150 0.5000 ;
      RECT 48.3250 0.0000 48.7350 0.5000 ;
      RECT 47.4050 0.0000 47.8150 0.5000 ;
      RECT 46.0250 0.0000 46.8950 0.5000 ;
      RECT 45.1050 0.0000 45.5150 0.5000 ;
      RECT 44.1850 0.0000 44.5950 0.5000 ;
      RECT 43.2650 0.0000 43.6750 0.5000 ;
      RECT 41.8850 0.0000 42.7550 0.5000 ;
      RECT 40.9650 0.0000 41.3750 0.5000 ;
      RECT 40.0450 0.0000 40.4550 0.5000 ;
      RECT 39.1250 0.0000 39.5350 0.5000 ;
      RECT 37.7450 0.0000 38.6150 0.5000 ;
      RECT 36.8250 0.0000 37.2350 0.5000 ;
      RECT 35.9050 0.0000 36.3150 0.5000 ;
      RECT 34.5250 0.0000 35.3950 0.5000 ;
      RECT 33.6050 0.0000 34.0150 0.5000 ;
      RECT 32.6850 0.0000 33.0950 0.5000 ;
      RECT 31.7650 0.0000 32.1750 0.5000 ;
      RECT 30.3850 0.0000 31.2550 0.5000 ;
      RECT 29.4650 0.0000 29.8750 0.5000 ;
      RECT 28.5450 0.0000 28.9550 0.5000 ;
      RECT 27.1650 0.0000 28.0350 0.5000 ;
      RECT 26.2450 0.0000 26.6550 0.5000 ;
      RECT 25.3250 0.0000 25.7350 0.5000 ;
      RECT 24.4050 0.0000 24.8150 0.5000 ;
      RECT 23.0250 0.0000 23.8950 0.5000 ;
      RECT 22.1050 0.0000 22.5150 0.5000 ;
      RECT 21.1850 0.0000 21.5950 0.5000 ;
      RECT 19.8050 0.0000 20.6750 0.5000 ;
      RECT 18.8850 0.0000 19.2950 0.5000 ;
      RECT 17.9650 0.0000 18.3750 0.5000 ;
      RECT 17.0450 0.0000 17.4550 0.5000 ;
      RECT 15.6650 0.0000 16.5350 0.5000 ;
      RECT 14.7450 0.0000 15.1550 0.5000 ;
      RECT 13.8250 0.0000 14.2350 0.5000 ;
      RECT 12.4450 0.0000 13.3150 0.5000 ;
      RECT 11.5250 0.0000 11.9350 0.5000 ;
      RECT 10.6050 0.0000 11.0150 0.5000 ;
      RECT 9.6850 0.0000 10.0950 0.5000 ;
      RECT 8.3050 0.0000 9.1750 0.5000 ;
      RECT 7.3850 0.0000 7.7950 0.5000 ;
      RECT 6.4650 0.0000 6.8750 0.5000 ;
      RECT 5.5450 0.0000 5.9550 0.5000 ;
      RECT 0.0000 0.0000 5.0350 0.5000 ;
    LAYER met1 ;
      RECT 0.0000 149.9800 100.2800 219.6400 ;
      RECT 0.7350 149.5600 99.5450 149.9800 ;
      RECT 0.0000 148.2800 100.2800 149.5600 ;
      RECT 0.7350 147.8600 100.2800 148.2800 ;
      RECT 0.0000 146.9200 100.2800 147.8600 ;
      RECT 0.7350 146.5800 100.2800 146.9200 ;
      RECT 0.7350 146.5000 99.5450 146.5800 ;
      RECT 0.0000 146.1600 99.5450 146.5000 ;
      RECT 0.0000 145.5600 100.2800 146.1600 ;
      RECT 0.7350 145.1400 100.2800 145.5600 ;
      RECT 0.0000 143.8600 100.2800 145.1400 ;
      RECT 0.7350 143.4400 99.5450 143.8600 ;
      RECT 0.0000 142.5000 100.2800 143.4400 ;
      RECT 0.7350 142.0800 100.2800 142.5000 ;
      RECT 0.0000 141.1400 100.2800 142.0800 ;
      RECT 0.7350 140.8000 100.2800 141.1400 ;
      RECT 0.7350 140.7200 99.5450 140.8000 ;
      RECT 0.0000 140.3800 99.5450 140.7200 ;
      RECT 0.0000 139.4400 100.2800 140.3800 ;
      RECT 0.7350 139.0200 100.2800 139.4400 ;
      RECT 0.0000 138.0800 100.2800 139.0200 ;
      RECT 0.7350 137.6600 99.5450 138.0800 ;
      RECT 0.0000 136.7200 100.2800 137.6600 ;
      RECT 0.7350 136.3000 100.2800 136.7200 ;
      RECT 0.0000 135.0200 100.2800 136.3000 ;
      RECT 0.7350 134.6000 99.5450 135.0200 ;
      RECT 0.0000 133.6600 100.2800 134.6000 ;
      RECT 0.7350 133.2400 100.2800 133.6600 ;
      RECT 0.0000 132.3000 100.2800 133.2400 ;
      RECT 0.7350 131.9600 100.2800 132.3000 ;
      RECT 0.7350 131.8800 99.5450 131.9600 ;
      RECT 0.0000 131.5400 99.5450 131.8800 ;
      RECT 0.0000 130.6000 100.2800 131.5400 ;
      RECT 0.7350 130.1800 100.2800 130.6000 ;
      RECT 0.0000 129.2400 100.2800 130.1800 ;
      RECT 0.7350 128.9000 100.2800 129.2400 ;
      RECT 0.7350 128.8200 99.5450 128.9000 ;
      RECT 0.0000 128.4800 99.5450 128.8200 ;
      RECT 0.0000 127.8800 100.2800 128.4800 ;
      RECT 0.7350 127.4600 100.2800 127.8800 ;
      RECT 0.0000 126.1800 100.2800 127.4600 ;
      RECT 0.7350 125.7600 99.5450 126.1800 ;
      RECT 0.0000 124.8200 100.2800 125.7600 ;
      RECT 0.7350 124.4000 100.2800 124.8200 ;
      RECT 0.0000 123.4600 100.2800 124.4000 ;
      RECT 0.7350 123.0400 100.2800 123.4600 ;
      RECT 0.0000 122.7800 100.2800 123.0400 ;
      RECT 0.0000 122.3600 99.5450 122.7800 ;
      RECT 0.0000 121.7600 100.2800 122.3600 ;
      RECT 0.7350 121.3400 100.2800 121.7600 ;
      RECT 0.0000 120.4000 100.2800 121.3400 ;
      RECT 0.7350 120.0600 100.2800 120.4000 ;
      RECT 0.7350 119.9800 99.5450 120.0600 ;
      RECT 0.0000 119.6400 99.5450 119.9800 ;
      RECT 0.0000 119.0400 100.2800 119.6400 ;
      RECT 0.7350 118.6200 100.2800 119.0400 ;
      RECT 0.0000 117.3400 100.2800 118.6200 ;
      RECT 0.7350 117.0000 100.2800 117.3400 ;
      RECT 0.7350 116.9200 99.5450 117.0000 ;
      RECT 0.0000 116.5800 99.5450 116.9200 ;
      RECT 0.0000 115.9800 100.2800 116.5800 ;
      RECT 0.7350 115.5600 100.2800 115.9800 ;
      RECT 0.0000 114.6200 100.2800 115.5600 ;
      RECT 0.7350 114.2800 100.2800 114.6200 ;
      RECT 0.7350 114.2000 99.5450 114.2800 ;
      RECT 0.0000 113.8600 99.5450 114.2000 ;
      RECT 0.0000 112.9200 100.2800 113.8600 ;
      RECT 0.7350 112.5000 100.2800 112.9200 ;
      RECT 0.0000 111.5600 100.2800 112.5000 ;
      RECT 0.7350 111.2200 100.2800 111.5600 ;
      RECT 0.7350 111.1400 99.5450 111.2200 ;
      RECT 0.0000 110.8000 99.5450 111.1400 ;
      RECT 0.0000 110.2000 100.2800 110.8000 ;
      RECT 0.7350 109.7800 100.2800 110.2000 ;
      RECT 0.0000 108.5000 100.2800 109.7800 ;
      RECT 0.7350 108.1600 100.2800 108.5000 ;
      RECT 0.7350 108.0800 99.5450 108.1600 ;
      RECT 0.0000 107.7400 99.5450 108.0800 ;
      RECT 0.0000 106.8000 100.2800 107.7400 ;
      RECT 0.7350 106.3800 100.2800 106.8000 ;
      RECT 0.0000 105.7800 100.2800 106.3800 ;
      RECT 0.7350 105.3600 100.2800 105.7800 ;
      RECT 0.0000 105.1000 100.2800 105.3600 ;
      RECT 0.0000 104.6800 99.5450 105.1000 ;
      RECT 0.0000 104.0800 100.2800 104.6800 ;
      RECT 0.7350 103.6600 100.2800 104.0800 ;
      RECT 0.0000 102.7200 100.2800 103.6600 ;
      RECT 0.7350 102.3800 100.2800 102.7200 ;
      RECT 0.7350 102.3000 99.5450 102.3800 ;
      RECT 0.0000 101.9600 99.5450 102.3000 ;
      RECT 0.0000 101.3600 100.2800 101.9600 ;
      RECT 0.7350 100.9400 100.2800 101.3600 ;
      RECT 0.0000 99.6600 100.2800 100.9400 ;
      RECT 0.7350 99.2400 100.2800 99.6600 ;
      RECT 0.0000 98.9800 100.2800 99.2400 ;
      RECT 0.0000 98.5600 99.5450 98.9800 ;
      RECT 0.0000 98.3000 100.2800 98.5600 ;
      RECT 0.7350 97.8800 100.2800 98.3000 ;
      RECT 0.0000 96.9400 100.2800 97.8800 ;
      RECT 0.7350 96.5200 100.2800 96.9400 ;
      RECT 0.0000 96.2600 100.2800 96.5200 ;
      RECT 0.0000 95.8400 99.5450 96.2600 ;
      RECT 0.0000 95.2400 100.2800 95.8400 ;
      RECT 0.7350 94.8200 100.2800 95.2400 ;
      RECT 0.0000 93.8800 100.2800 94.8200 ;
      RECT 0.7350 93.4600 100.2800 93.8800 ;
      RECT 0.0000 93.2000 100.2800 93.4600 ;
      RECT 0.0000 92.7800 99.5450 93.2000 ;
      RECT 0.0000 92.5200 100.2800 92.7800 ;
      RECT 0.7350 92.1000 100.2800 92.5200 ;
      RECT 0.0000 90.4800 100.2800 92.1000 ;
      RECT 0.7350 90.0600 99.5450 90.4800 ;
      RECT 0.0000 89.1200 100.2800 90.0600 ;
      RECT 0.7350 88.7000 100.2800 89.1200 ;
      RECT 0.0000 88.1000 100.2800 88.7000 ;
      RECT 0.7350 87.6800 100.2800 88.1000 ;
      RECT 0.0000 87.4200 100.2800 87.6800 ;
      RECT 0.0000 87.0000 99.5450 87.4200 ;
      RECT 0.0000 86.4000 100.2800 87.0000 ;
      RECT 0.7350 85.9800 100.2800 86.4000 ;
      RECT 0.0000 85.0400 100.2800 85.9800 ;
      RECT 0.7350 84.6200 100.2800 85.0400 ;
      RECT 0.0000 84.3600 100.2800 84.6200 ;
      RECT 0.0000 83.9400 99.5450 84.3600 ;
      RECT 0.0000 83.6800 100.2800 83.9400 ;
      RECT 0.7350 83.2600 100.2800 83.6800 ;
      RECT 0.0000 81.6400 100.2800 83.2600 ;
      RECT 0.7350 81.3000 100.2800 81.6400 ;
      RECT 0.7350 81.2200 99.5450 81.3000 ;
      RECT 0.0000 80.8800 99.5450 81.2200 ;
      RECT 0.0000 80.6200 100.2800 80.8800 ;
      RECT 0.7350 80.2000 100.2800 80.6200 ;
      RECT 0.0000 79.2600 100.2800 80.2000 ;
      RECT 0.7350 78.8400 100.2800 79.2600 ;
      RECT 0.0000 78.5800 100.2800 78.8400 ;
      RECT 0.0000 78.1600 99.5450 78.5800 ;
      RECT 0.0000 77.9000 100.2800 78.1600 ;
      RECT 0.7350 77.4800 100.2800 77.9000 ;
      RECT 0.0000 76.2000 100.2800 77.4800 ;
      RECT 0.7350 75.7800 100.2800 76.2000 ;
      RECT 0.0000 75.5200 100.2800 75.7800 ;
      RECT 0.0000 75.1000 99.5450 75.5200 ;
      RECT 0.0000 74.8400 100.2800 75.1000 ;
      RECT 0.7350 74.4200 100.2800 74.8400 ;
      RECT 0.0000 73.4800 100.2800 74.4200 ;
      RECT 0.7350 73.0600 100.2800 73.4800 ;
      RECT 0.0000 72.4600 100.2800 73.0600 ;
      RECT 0.0000 72.0400 99.5450 72.4600 ;
      RECT 0.0000 71.7800 100.2800 72.0400 ;
      RECT 0.7350 71.3600 100.2800 71.7800 ;
      RECT 0.0000 70.4200 100.2800 71.3600 ;
      RECT 0.7350 70.0000 100.2800 70.4200 ;
      RECT 0.0000 69.4000 100.2800 70.0000 ;
      RECT 0.0000 69.0600 99.5450 69.4000 ;
      RECT 0.7350 68.9800 99.5450 69.0600 ;
      RECT 0.7350 68.6400 100.2800 68.9800 ;
      RECT 0.0000 67.3600 100.2800 68.6400 ;
      RECT 0.7350 66.9400 100.2800 67.3600 ;
      RECT 0.0000 66.3400 100.2800 66.9400 ;
      RECT 0.0000 66.0000 99.5450 66.3400 ;
      RECT 0.7350 65.9200 99.5450 66.0000 ;
      RECT 0.7350 65.5800 100.2800 65.9200 ;
      RECT 0.0000 64.6400 100.2800 65.5800 ;
      RECT 0.7350 64.2200 100.2800 64.6400 ;
      RECT 0.0000 63.6200 100.2800 64.2200 ;
      RECT 0.0000 63.2000 99.5450 63.6200 ;
      RECT 0.0000 62.6000 100.2800 63.2000 ;
      RECT 0.7350 62.1800 100.2800 62.6000 ;
      RECT 0.0000 61.5800 100.2800 62.1800 ;
      RECT 0.7350 61.1600 100.2800 61.5800 ;
      RECT 0.0000 60.5600 100.2800 61.1600 ;
      RECT 0.0000 60.2200 99.5450 60.5600 ;
      RECT 0.7350 60.1400 99.5450 60.2200 ;
      RECT 0.7350 59.8000 100.2800 60.1400 ;
      RECT 0.0000 58.5200 100.2800 59.8000 ;
      RECT 0.7350 58.1000 100.2800 58.5200 ;
      RECT 0.0000 57.5000 100.2800 58.1000 ;
      RECT 0.0000 57.1600 99.5450 57.5000 ;
      RECT 0.7350 57.0800 99.5450 57.1600 ;
      RECT 0.7350 56.7400 100.2800 57.0800 ;
      RECT 0.0000 55.8000 100.2800 56.7400 ;
      RECT 0.7350 55.3800 100.2800 55.8000 ;
      RECT 0.0000 54.7800 100.2800 55.3800 ;
      RECT 0.0000 54.3600 99.5450 54.7800 ;
      RECT 0.0000 54.1000 100.2800 54.3600 ;
      RECT 0.7350 53.6800 100.2800 54.1000 ;
      RECT 0.0000 52.7400 100.2800 53.6800 ;
      RECT 0.7350 52.3200 100.2800 52.7400 ;
      RECT 0.0000 51.7200 100.2800 52.3200 ;
      RECT 0.0000 51.3800 99.5450 51.7200 ;
      RECT 0.7350 51.3000 99.5450 51.3800 ;
      RECT 0.7350 50.9600 100.2800 51.3000 ;
      RECT 0.0000 49.6800 100.2800 50.9600 ;
      RECT 0.7350 49.2600 100.2800 49.6800 ;
      RECT 0.0000 48.6600 100.2800 49.2600 ;
      RECT 0.0000 48.3200 99.5450 48.6600 ;
      RECT 0.7350 48.2400 99.5450 48.3200 ;
      RECT 0.7350 47.9000 100.2800 48.2400 ;
      RECT 0.0000 46.9600 100.2800 47.9000 ;
      RECT 0.7350 46.5400 100.2800 46.9600 ;
      RECT 0.0000 45.6000 100.2800 46.5400 ;
      RECT 0.0000 45.2600 99.5450 45.6000 ;
      RECT 0.7350 45.1800 99.5450 45.2600 ;
      RECT 0.7350 44.8400 100.2800 45.1800 ;
      RECT 0.0000 43.9000 100.2800 44.8400 ;
      RECT 0.7350 43.4800 100.2800 43.9000 ;
      RECT 0.0000 42.8800 100.2800 43.4800 ;
      RECT 0.0000 42.5400 99.5450 42.8800 ;
      RECT 0.7350 42.4600 99.5450 42.5400 ;
      RECT 0.7350 42.1200 100.2800 42.4600 ;
      RECT 0.0000 40.8400 100.2800 42.1200 ;
      RECT 0.7350 40.4200 100.2800 40.8400 ;
      RECT 0.0000 39.8200 100.2800 40.4200 ;
      RECT 0.0000 39.4800 99.5450 39.8200 ;
      RECT 0.7350 39.4000 99.5450 39.4800 ;
      RECT 0.7350 39.0600 100.2800 39.4000 ;
      RECT 0.0000 38.1200 100.2800 39.0600 ;
      RECT 0.7350 37.7000 100.2800 38.1200 ;
      RECT 0.0000 36.7600 100.2800 37.7000 ;
      RECT 0.0000 36.4200 99.5450 36.7600 ;
      RECT 0.7350 36.3400 99.5450 36.4200 ;
      RECT 0.7350 36.0000 100.2800 36.3400 ;
      RECT 0.0000 35.0600 100.2800 36.0000 ;
      RECT 0.7350 34.6400 100.2800 35.0600 ;
      RECT 0.0000 33.7000 100.2800 34.6400 ;
      RECT 0.7350 33.2800 99.5450 33.7000 ;
      RECT 0.0000 32.0000 100.2800 33.2800 ;
      RECT 0.7350 31.5800 100.2800 32.0000 ;
      RECT 0.0000 30.9800 100.2800 31.5800 ;
      RECT 0.0000 30.6400 99.5450 30.9800 ;
      RECT 0.7350 30.5600 99.5450 30.6400 ;
      RECT 0.7350 30.2200 100.2800 30.5600 ;
      RECT 0.0000 29.2800 100.2800 30.2200 ;
      RECT 0.7350 28.8600 100.2800 29.2800 ;
      RECT 0.0000 27.9200 100.2800 28.8600 ;
      RECT 0.0000 27.5800 99.5450 27.9200 ;
      RECT 0.7350 27.5000 99.5450 27.5800 ;
      RECT 0.7350 27.1600 100.2800 27.5000 ;
      RECT 0.0000 26.2200 100.2800 27.1600 ;
      RECT 0.7350 25.8000 100.2800 26.2200 ;
      RECT 0.0000 24.8600 100.2800 25.8000 ;
      RECT 0.7350 24.4400 99.5450 24.8600 ;
      RECT 0.0000 23.1600 100.2800 24.4400 ;
      RECT 0.7350 22.7400 100.2800 23.1600 ;
      RECT 0.0000 21.8000 100.2800 22.7400 ;
      RECT 0.7350 21.3800 99.5450 21.8000 ;
      RECT 0.0000 20.4400 100.2800 21.3800 ;
      RECT 0.7350 20.0200 100.2800 20.4400 ;
      RECT 0.0000 19.0800 100.2800 20.0200 ;
      RECT 0.0000 18.7400 99.5450 19.0800 ;
      RECT 0.7350 18.6600 99.5450 18.7400 ;
      RECT 0.7350 18.3200 100.2800 18.6600 ;
      RECT 0.0000 17.3800 100.2800 18.3200 ;
      RECT 0.7350 16.9600 100.2800 17.3800 ;
      RECT 0.0000 16.0200 100.2800 16.9600 ;
      RECT 0.7350 15.6000 99.5450 16.0200 ;
      RECT 0.0000 14.3200 100.2800 15.6000 ;
      RECT 0.7350 13.9000 100.2800 14.3200 ;
      RECT 0.0000 12.9600 100.2800 13.9000 ;
      RECT 0.7350 12.5400 99.5450 12.9600 ;
      RECT 0.0000 11.6000 100.2800 12.5400 ;
      RECT 0.7350 11.1800 100.2800 11.6000 ;
      RECT 0.0000 10.2400 100.2800 11.1800 ;
      RECT 0.7350 9.8200 99.5450 10.2400 ;
      RECT 0.0000 0.0000 100.2800 9.8200 ;
    LAYER met2 ;
      RECT 97.9600 219.0150 100.2800 219.6400 ;
      RECT 97.0400 219.0150 97.5400 219.6400 ;
      RECT 96.1200 219.0150 96.6200 219.6400 ;
      RECT 95.2000 219.0150 95.7000 219.6400 ;
      RECT 94.2800 219.0150 94.7800 219.6400 ;
      RECT 93.8200 219.0150 93.8600 219.6400 ;
      RECT 92.9000 219.0150 93.4000 219.6400 ;
      RECT 91.9800 219.0150 92.4800 219.6400 ;
      RECT 91.0600 219.0150 91.5600 219.6400 ;
      RECT 90.1400 219.0150 90.6400 219.6400 ;
      RECT 89.6800 219.0150 89.7200 219.6400 ;
      RECT 88.7600 219.0150 89.2600 219.6400 ;
      RECT 87.8400 219.0150 88.3400 219.6400 ;
      RECT 86.9200 219.0150 87.4200 219.6400 ;
      RECT 86.0000 219.0150 86.5000 219.6400 ;
      RECT 85.5400 219.0150 85.5800 219.6400 ;
      RECT 84.1600 219.0150 85.1200 219.6400 ;
      RECT 83.7000 219.0150 83.7400 219.6400 ;
      RECT 83.2400 219.0150 83.2800 219.6400 ;
      RECT 82.3200 219.0150 82.8200 219.6400 ;
      RECT 0.0000 219.0150 81.9000 219.6400 ;
      RECT 0.0000 0.6250 100.2800 219.0150 ;
      RECT 97.5000 0.0000 100.2800 0.6250 ;
      RECT 97.0400 0.0000 97.0800 0.6250 ;
      RECT 96.1200 0.0000 96.6200 0.6250 ;
      RECT 95.2000 0.0000 95.7000 0.6250 ;
      RECT 94.7400 0.0000 94.7800 0.6250 ;
      RECT 92.9000 0.0000 94.3200 0.6250 ;
      RECT 92.4400 0.0000 92.4800 0.6250 ;
      RECT 91.5200 0.0000 92.0200 0.6250 ;
      RECT 90.6000 0.0000 91.1000 0.6250 ;
      RECT 89.6800 0.0000 90.1800 0.6250 ;
      RECT 89.2200 0.0000 89.2600 0.6250 ;
      RECT 88.3000 0.0000 88.8000 0.6250 ;
      RECT 87.3800 0.0000 87.8800 0.6250 ;
      RECT 86.9200 0.0000 86.9600 0.6250 ;
      RECT 86.0000 0.0000 86.5000 0.6250 ;
      RECT 85.0800 0.0000 85.5800 0.6250 ;
      RECT 84.6200 0.0000 84.6600 0.6250 ;
      RECT 83.7000 0.0000 84.2000 0.6250 ;
      RECT 82.7800 0.0000 83.2800 0.6250 ;
      RECT 82.3200 0.0000 82.3600 0.6250 ;
      RECT 0.0000 0.0000 81.9000 0.6250 ;
    LAYER met3 ;
      RECT 0.0000 216.3300 100.2800 219.6400 ;
      RECT 97.5200 214.2300 100.2800 216.3300 ;
      RECT 0.0000 214.2300 2.7600 216.3300 ;
      RECT 0.0000 213.8300 100.2800 214.2300 ;
      RECT 95.0200 211.7300 100.2800 213.8300 ;
      RECT 0.0000 211.7300 5.2600 213.8300 ;
      RECT 0.0000 209.9500 100.2800 211.7300 ;
      RECT 1.1000 209.0500 99.1800 209.9500 ;
      RECT 0.0000 208.9600 100.2800 209.0500 ;
      RECT 95.0200 208.1200 100.2800 208.9600 ;
      RECT 0.0000 208.1200 5.2600 208.9600 ;
      RECT 95.0200 207.8800 99.1800 208.1200 ;
      RECT 7.3600 207.8800 92.9200 208.9600 ;
      RECT 1.1000 207.8800 5.2600 208.1200 ;
      RECT 1.1000 207.2200 99.1800 207.8800 ;
      RECT 0.0000 206.2900 100.2800 207.2200 ;
      RECT 1.1000 206.2400 99.1800 206.2900 ;
      RECT 97.5200 205.3900 99.1800 206.2400 ;
      RECT 1.1000 205.3900 2.7600 206.2400 ;
      RECT 97.5200 205.1600 100.2800 205.3900 ;
      RECT 4.8600 205.1600 95.4200 206.2400 ;
      RECT 0.0000 205.1600 2.7600 205.3900 ;
      RECT 0.0000 204.4600 100.2800 205.1600 ;
      RECT 1.1000 203.5600 99.1800 204.4600 ;
      RECT 0.0000 203.5200 100.2800 203.5600 ;
      RECT 95.0200 202.6300 100.2800 203.5200 ;
      RECT 0.0000 202.6300 5.2600 203.5200 ;
      RECT 95.0200 202.4400 99.1800 202.6300 ;
      RECT 7.3600 202.4400 92.9200 203.5200 ;
      RECT 1.1000 202.4400 5.2600 202.6300 ;
      RECT 1.1000 201.7300 99.1800 202.4400 ;
      RECT 0.0000 200.8000 100.2800 201.7300 ;
      RECT 97.5200 199.9000 99.1800 200.8000 ;
      RECT 1.1000 199.9000 2.7600 200.8000 ;
      RECT 97.5200 199.7200 100.2800 199.9000 ;
      RECT 4.8600 199.7200 95.4200 200.8000 ;
      RECT 0.0000 199.7200 2.7600 199.9000 ;
      RECT 0.0000 198.9700 100.2800 199.7200 ;
      RECT 1.1000 198.0800 99.1800 198.9700 ;
      RECT 95.0200 198.0700 99.1800 198.0800 ;
      RECT 1.1000 198.0700 5.2600 198.0800 ;
      RECT 95.0200 197.1400 100.2800 198.0700 ;
      RECT 0.0000 197.1400 5.2600 198.0700 ;
      RECT 95.0200 197.0000 99.1800 197.1400 ;
      RECT 7.3600 197.0000 92.9200 198.0800 ;
      RECT 1.1000 197.0000 5.2600 197.1400 ;
      RECT 1.1000 196.2400 99.1800 197.0000 ;
      RECT 0.0000 195.9200 100.2800 196.2400 ;
      RECT 1.1000 195.3600 99.1800 195.9200 ;
      RECT 97.5200 195.0200 99.1800 195.3600 ;
      RECT 1.1000 195.0200 2.7600 195.3600 ;
      RECT 97.5200 194.2800 100.2800 195.0200 ;
      RECT 4.8600 194.2800 95.4200 195.3600 ;
      RECT 0.0000 194.2800 2.7600 195.0200 ;
      RECT 0.0000 194.0900 100.2800 194.2800 ;
      RECT 1.1000 193.1900 99.1800 194.0900 ;
      RECT 0.0000 192.6400 100.2800 193.1900 ;
      RECT 95.0200 192.2600 100.2800 192.6400 ;
      RECT 0.0000 192.2600 5.2600 192.6400 ;
      RECT 95.0200 191.5600 99.1800 192.2600 ;
      RECT 7.3600 191.5600 92.9200 192.6400 ;
      RECT 1.1000 191.5600 5.2600 192.2600 ;
      RECT 1.1000 191.3600 99.1800 191.5600 ;
      RECT 0.0000 190.4300 100.2800 191.3600 ;
      RECT 1.1000 189.9200 99.1800 190.4300 ;
      RECT 97.5200 189.5300 99.1800 189.9200 ;
      RECT 1.1000 189.5300 2.7600 189.9200 ;
      RECT 97.5200 188.8400 100.2800 189.5300 ;
      RECT 4.8600 188.8400 95.4200 189.9200 ;
      RECT 0.0000 188.8400 2.7600 189.5300 ;
      RECT 0.0000 188.6000 100.2800 188.8400 ;
      RECT 1.1000 187.7000 99.1800 188.6000 ;
      RECT 0.0000 187.2000 100.2800 187.7000 ;
      RECT 95.0200 186.7700 100.2800 187.2000 ;
      RECT 0.0000 186.7700 5.2600 187.2000 ;
      RECT 95.0200 186.1200 99.1800 186.7700 ;
      RECT 7.3600 186.1200 92.9200 187.2000 ;
      RECT 1.1000 186.1200 5.2600 186.7700 ;
      RECT 1.1000 185.8700 99.1800 186.1200 ;
      RECT 0.0000 184.9400 100.2800 185.8700 ;
      RECT 1.1000 184.4800 99.1800 184.9400 ;
      RECT 97.5200 184.0400 99.1800 184.4800 ;
      RECT 1.1000 184.0400 2.7600 184.4800 ;
      RECT 97.5200 183.4000 100.2800 184.0400 ;
      RECT 4.8600 183.4000 95.4200 184.4800 ;
      RECT 0.0000 183.4000 2.7600 184.0400 ;
      RECT 0.0000 183.1100 100.2800 183.4000 ;
      RECT 1.1000 182.2100 99.1800 183.1100 ;
      RECT 0.0000 181.8900 100.2800 182.2100 ;
      RECT 1.1000 181.7600 99.1800 181.8900 ;
      RECT 95.0200 180.9900 99.1800 181.7600 ;
      RECT 1.1000 180.9900 5.2600 181.7600 ;
      RECT 95.0200 180.6800 100.2800 180.9900 ;
      RECT 7.3600 180.6800 92.9200 181.7600 ;
      RECT 0.0000 180.6800 5.2600 180.9900 ;
      RECT 0.0000 180.0600 100.2800 180.6800 ;
      RECT 1.1000 179.1600 99.1800 180.0600 ;
      RECT 0.0000 179.0400 100.2800 179.1600 ;
      RECT 97.5200 178.2300 100.2800 179.0400 ;
      RECT 0.0000 178.2300 2.7600 179.0400 ;
      RECT 97.5200 177.9600 99.1800 178.2300 ;
      RECT 4.8600 177.9600 95.4200 179.0400 ;
      RECT 1.1000 177.9600 2.7600 178.2300 ;
      RECT 1.1000 177.3300 99.1800 177.9600 ;
      RECT 0.0000 176.4000 100.2800 177.3300 ;
      RECT 1.1000 176.3200 99.1800 176.4000 ;
      RECT 95.0200 175.5000 99.1800 176.3200 ;
      RECT 1.1000 175.5000 5.2600 176.3200 ;
      RECT 95.0200 175.2400 100.2800 175.5000 ;
      RECT 7.3600 175.2400 92.9200 176.3200 ;
      RECT 0.0000 175.2400 5.2600 175.5000 ;
      RECT 0.0000 174.5700 100.2800 175.2400 ;
      RECT 1.1000 173.6700 99.1800 174.5700 ;
      RECT 0.0000 173.6000 100.2800 173.6700 ;
      RECT 97.5200 172.7400 100.2800 173.6000 ;
      RECT 0.0000 172.7400 2.7600 173.6000 ;
      RECT 97.5200 172.5200 99.1800 172.7400 ;
      RECT 4.8600 172.5200 95.4200 173.6000 ;
      RECT 1.1000 172.5200 2.7600 172.7400 ;
      RECT 1.1000 171.8400 99.1800 172.5200 ;
      RECT 0.0000 170.9100 100.2800 171.8400 ;
      RECT 1.1000 170.8800 99.1800 170.9100 ;
      RECT 95.0200 170.0100 99.1800 170.8800 ;
      RECT 1.1000 170.0100 5.2600 170.8800 ;
      RECT 95.0200 169.8000 100.2800 170.0100 ;
      RECT 7.3600 169.8000 92.9200 170.8800 ;
      RECT 0.0000 169.8000 5.2600 170.0100 ;
      RECT 0.0000 169.0800 100.2800 169.8000 ;
      RECT 1.1000 168.1800 99.1800 169.0800 ;
      RECT 0.0000 168.1600 100.2800 168.1800 ;
      RECT 97.5200 167.8600 100.2800 168.1600 ;
      RECT 0.0000 167.8600 2.7600 168.1600 ;
      RECT 97.5200 167.0800 99.1800 167.8600 ;
      RECT 4.8600 167.0800 95.4200 168.1600 ;
      RECT 1.1000 167.0800 2.7600 167.8600 ;
      RECT 1.1000 166.9600 99.1800 167.0800 ;
      RECT 0.0000 166.0300 100.2800 166.9600 ;
      RECT 1.1000 165.4400 99.1800 166.0300 ;
      RECT 95.0200 165.1300 99.1800 165.4400 ;
      RECT 1.1000 165.1300 5.2600 165.4400 ;
      RECT 95.0200 164.3600 100.2800 165.1300 ;
      RECT 7.3600 164.3600 92.9200 165.4400 ;
      RECT 0.0000 164.3600 5.2600 165.1300 ;
      RECT 0.0000 164.2000 100.2800 164.3600 ;
      RECT 1.1000 163.3000 99.1800 164.2000 ;
      RECT 0.0000 162.7200 100.2800 163.3000 ;
      RECT 97.5200 162.3700 100.2800 162.7200 ;
      RECT 0.0000 162.3700 2.7600 162.7200 ;
      RECT 97.5200 161.6400 99.1800 162.3700 ;
      RECT 4.8600 161.6400 95.4200 162.7200 ;
      RECT 1.1000 161.6400 2.7600 162.3700 ;
      RECT 1.1000 161.4700 99.1800 161.6400 ;
      RECT 0.0000 160.5400 100.2800 161.4700 ;
      RECT 1.1000 160.0000 99.1800 160.5400 ;
      RECT 95.0200 159.6400 99.1800 160.0000 ;
      RECT 1.1000 159.6400 5.2600 160.0000 ;
      RECT 95.0200 158.9200 100.2800 159.6400 ;
      RECT 7.3600 158.9200 92.9200 160.0000 ;
      RECT 0.0000 158.9200 5.2600 159.6400 ;
      RECT 0.0000 158.7100 100.2800 158.9200 ;
      RECT 1.1000 158.1000 100.2800 158.7100 ;
      RECT 1.1000 157.8100 99.1800 158.1000 ;
      RECT 0.0000 157.2800 99.1800 157.8100 ;
      RECT 97.5200 157.2000 99.1800 157.2800 ;
      RECT 97.5200 156.8800 100.2800 157.2000 ;
      RECT 0.0000 156.8800 2.7600 157.2800 ;
      RECT 97.5200 156.2000 99.1800 156.8800 ;
      RECT 4.8600 156.2000 95.4200 157.2800 ;
      RECT 1.1000 156.2000 2.7600 156.8800 ;
      RECT 1.1000 155.9800 99.1800 156.2000 ;
      RECT 0.0000 155.6600 100.2800 155.9800 ;
      RECT 1.1000 154.7600 99.1800 155.6600 ;
      RECT 0.0000 154.5600 100.2800 154.7600 ;
      RECT 95.0200 153.4800 100.2800 154.5600 ;
      RECT 7.3600 153.4800 92.9200 154.5600 ;
      RECT 0.0000 153.4800 5.2600 154.5600 ;
      RECT 0.0000 151.8400 100.2800 153.4800 ;
      RECT 97.5200 150.7600 100.2800 151.8400 ;
      RECT 4.8600 150.7600 95.4200 151.8400 ;
      RECT 0.0000 150.7600 2.7600 151.8400 ;
      RECT 0.0000 149.1200 100.2800 150.7600 ;
      RECT 95.0200 148.0400 100.2800 149.1200 ;
      RECT 7.3600 148.0400 92.9200 149.1200 ;
      RECT 0.0000 148.0400 5.2600 149.1200 ;
      RECT 0.0000 146.4000 100.2800 148.0400 ;
      RECT 97.5200 145.3200 100.2800 146.4000 ;
      RECT 4.8600 145.3200 95.4200 146.4000 ;
      RECT 0.0000 145.3200 2.7600 146.4000 ;
      RECT 0.0000 143.6800 100.2800 145.3200 ;
      RECT 95.0200 142.6000 100.2800 143.6800 ;
      RECT 7.3600 142.6000 92.9200 143.6800 ;
      RECT 0.0000 142.6000 5.2600 143.6800 ;
      RECT 0.0000 140.9600 100.2800 142.6000 ;
      RECT 97.5200 139.8800 100.2800 140.9600 ;
      RECT 4.8600 139.8800 95.4200 140.9600 ;
      RECT 0.0000 139.8800 2.7600 140.9600 ;
      RECT 0.0000 138.2400 100.2800 139.8800 ;
      RECT 95.0200 137.1600 100.2800 138.2400 ;
      RECT 7.3600 137.1600 92.9200 138.2400 ;
      RECT 0.0000 137.1600 5.2600 138.2400 ;
      RECT 0.0000 135.5200 100.2800 137.1600 ;
      RECT 97.5200 134.4400 100.2800 135.5200 ;
      RECT 4.8600 134.4400 95.4200 135.5200 ;
      RECT 0.0000 134.4400 2.7600 135.5200 ;
      RECT 0.0000 132.8000 100.2800 134.4400 ;
      RECT 95.0200 131.7200 100.2800 132.8000 ;
      RECT 7.3600 131.7200 92.9200 132.8000 ;
      RECT 0.0000 131.7200 5.2600 132.8000 ;
      RECT 0.0000 130.0800 100.2800 131.7200 ;
      RECT 97.5200 129.0000 100.2800 130.0800 ;
      RECT 4.8600 129.0000 95.4200 130.0800 ;
      RECT 0.0000 129.0000 2.7600 130.0800 ;
      RECT 0.0000 127.3600 100.2800 129.0000 ;
      RECT 95.0200 126.2800 100.2800 127.3600 ;
      RECT 7.3600 126.2800 92.9200 127.3600 ;
      RECT 0.0000 126.2800 5.2600 127.3600 ;
      RECT 0.0000 124.6400 100.2800 126.2800 ;
      RECT 97.5200 123.5600 100.2800 124.6400 ;
      RECT 4.8600 123.5600 95.4200 124.6400 ;
      RECT 0.0000 123.5600 2.7600 124.6400 ;
      RECT 0.0000 121.9200 100.2800 123.5600 ;
      RECT 95.0200 120.8400 100.2800 121.9200 ;
      RECT 7.3600 120.8400 92.9200 121.9200 ;
      RECT 0.0000 120.8400 5.2600 121.9200 ;
      RECT 0.0000 119.2000 100.2800 120.8400 ;
      RECT 97.5200 118.1200 100.2800 119.2000 ;
      RECT 4.8600 118.1200 95.4200 119.2000 ;
      RECT 0.0000 118.1200 2.7600 119.2000 ;
      RECT 0.0000 116.4800 100.2800 118.1200 ;
      RECT 95.0200 115.4000 100.2800 116.4800 ;
      RECT 7.3600 115.4000 92.9200 116.4800 ;
      RECT 0.0000 115.4000 5.2600 116.4800 ;
      RECT 0.0000 113.7600 100.2800 115.4000 ;
      RECT 97.5200 112.6800 100.2800 113.7600 ;
      RECT 4.8600 112.6800 95.4200 113.7600 ;
      RECT 0.0000 112.6800 2.7600 113.7600 ;
      RECT 0.0000 111.0400 100.2800 112.6800 ;
      RECT 95.0200 109.9600 100.2800 111.0400 ;
      RECT 7.3600 109.9600 92.9200 111.0400 ;
      RECT 0.0000 109.9600 5.2600 111.0400 ;
      RECT 0.0000 108.3200 100.2800 109.9600 ;
      RECT 97.5200 107.2400 100.2800 108.3200 ;
      RECT 4.8600 107.2400 95.4200 108.3200 ;
      RECT 0.0000 107.2400 2.7600 108.3200 ;
      RECT 0.0000 105.6000 100.2800 107.2400 ;
      RECT 95.0200 104.5200 100.2800 105.6000 ;
      RECT 7.3600 104.5200 92.9200 105.6000 ;
      RECT 0.0000 104.5200 5.2600 105.6000 ;
      RECT 0.0000 102.8800 100.2800 104.5200 ;
      RECT 97.5200 101.8000 100.2800 102.8800 ;
      RECT 4.8600 101.8000 95.4200 102.8800 ;
      RECT 0.0000 101.8000 2.7600 102.8800 ;
      RECT 0.0000 100.1600 100.2800 101.8000 ;
      RECT 95.0200 99.0800 100.2800 100.1600 ;
      RECT 7.3600 99.0800 92.9200 100.1600 ;
      RECT 0.0000 99.0800 5.2600 100.1600 ;
      RECT 0.0000 97.4400 100.2800 99.0800 ;
      RECT 97.5200 96.3600 100.2800 97.4400 ;
      RECT 4.8600 96.3600 95.4200 97.4400 ;
      RECT 0.0000 96.3600 2.7600 97.4400 ;
      RECT 0.0000 94.7200 100.2800 96.3600 ;
      RECT 95.0200 93.6400 100.2800 94.7200 ;
      RECT 7.3600 93.6400 92.9200 94.7200 ;
      RECT 0.0000 93.6400 5.2600 94.7200 ;
      RECT 0.0000 92.0000 100.2800 93.6400 ;
      RECT 97.5200 90.9200 100.2800 92.0000 ;
      RECT 4.8600 90.9200 95.4200 92.0000 ;
      RECT 0.0000 90.9200 2.7600 92.0000 ;
      RECT 0.0000 89.2800 100.2800 90.9200 ;
      RECT 95.0200 88.2000 100.2800 89.2800 ;
      RECT 7.3600 88.2000 92.9200 89.2800 ;
      RECT 0.0000 88.2000 5.2600 89.2800 ;
      RECT 0.0000 86.5600 100.2800 88.2000 ;
      RECT 97.5200 85.4800 100.2800 86.5600 ;
      RECT 4.8600 85.4800 95.4200 86.5600 ;
      RECT 0.0000 85.4800 2.7600 86.5600 ;
      RECT 0.0000 83.8400 100.2800 85.4800 ;
      RECT 95.0200 82.7600 100.2800 83.8400 ;
      RECT 7.3600 82.7600 92.9200 83.8400 ;
      RECT 0.0000 82.7600 5.2600 83.8400 ;
      RECT 0.0000 81.1200 100.2800 82.7600 ;
      RECT 97.5200 80.0400 100.2800 81.1200 ;
      RECT 4.8600 80.0400 95.4200 81.1200 ;
      RECT 0.0000 80.0400 2.7600 81.1200 ;
      RECT 0.0000 78.4000 100.2800 80.0400 ;
      RECT 95.0200 77.3200 100.2800 78.4000 ;
      RECT 7.3600 77.3200 92.9200 78.4000 ;
      RECT 0.0000 77.3200 5.2600 78.4000 ;
      RECT 0.0000 75.6800 100.2800 77.3200 ;
      RECT 97.5200 74.6000 100.2800 75.6800 ;
      RECT 4.8600 74.6000 95.4200 75.6800 ;
      RECT 0.0000 74.6000 2.7600 75.6800 ;
      RECT 0.0000 72.9600 100.2800 74.6000 ;
      RECT 95.0200 71.8800 100.2800 72.9600 ;
      RECT 7.3600 71.8800 92.9200 72.9600 ;
      RECT 0.0000 71.8800 5.2600 72.9600 ;
      RECT 0.0000 70.2400 100.2800 71.8800 ;
      RECT 97.5200 69.1600 100.2800 70.2400 ;
      RECT 4.8600 69.1600 95.4200 70.2400 ;
      RECT 0.0000 69.1600 2.7600 70.2400 ;
      RECT 0.0000 67.5200 100.2800 69.1600 ;
      RECT 95.0200 66.4400 100.2800 67.5200 ;
      RECT 7.3600 66.4400 92.9200 67.5200 ;
      RECT 0.0000 66.4400 5.2600 67.5200 ;
      RECT 0.0000 64.8000 100.2800 66.4400 ;
      RECT 97.5200 63.7200 100.2800 64.8000 ;
      RECT 4.8600 63.7200 95.4200 64.8000 ;
      RECT 0.0000 63.7200 2.7600 64.8000 ;
      RECT 0.0000 62.0800 100.2800 63.7200 ;
      RECT 95.0200 61.0000 100.2800 62.0800 ;
      RECT 7.3600 61.0000 92.9200 62.0800 ;
      RECT 0.0000 61.0000 5.2600 62.0800 ;
      RECT 0.0000 59.3600 100.2800 61.0000 ;
      RECT 97.5200 58.2800 100.2800 59.3600 ;
      RECT 4.8600 58.2800 95.4200 59.3600 ;
      RECT 0.0000 58.2800 2.7600 59.3600 ;
      RECT 0.0000 56.6400 100.2800 58.2800 ;
      RECT 95.0200 55.5600 100.2800 56.6400 ;
      RECT 7.3600 55.5600 92.9200 56.6400 ;
      RECT 0.0000 55.5600 5.2600 56.6400 ;
      RECT 0.0000 53.9200 100.2800 55.5600 ;
      RECT 97.5200 52.8400 100.2800 53.9200 ;
      RECT 4.8600 52.8400 95.4200 53.9200 ;
      RECT 0.0000 52.8400 2.7600 53.9200 ;
      RECT 0.0000 51.2000 100.2800 52.8400 ;
      RECT 95.0200 50.1200 100.2800 51.2000 ;
      RECT 7.3600 50.1200 92.9200 51.2000 ;
      RECT 0.0000 50.1200 5.2600 51.2000 ;
      RECT 0.0000 48.4800 100.2800 50.1200 ;
      RECT 97.5200 47.4000 100.2800 48.4800 ;
      RECT 4.8600 47.4000 95.4200 48.4800 ;
      RECT 0.0000 47.4000 2.7600 48.4800 ;
      RECT 0.0000 45.7600 100.2800 47.4000 ;
      RECT 95.0200 44.6800 100.2800 45.7600 ;
      RECT 7.3600 44.6800 92.9200 45.7600 ;
      RECT 0.0000 44.6800 5.2600 45.7600 ;
      RECT 0.0000 43.0400 100.2800 44.6800 ;
      RECT 97.5200 41.9600 100.2800 43.0400 ;
      RECT 4.8600 41.9600 95.4200 43.0400 ;
      RECT 0.0000 41.9600 2.7600 43.0400 ;
      RECT 0.0000 40.3200 100.2800 41.9600 ;
      RECT 95.0200 39.2400 100.2800 40.3200 ;
      RECT 7.3600 39.2400 92.9200 40.3200 ;
      RECT 0.0000 39.2400 5.2600 40.3200 ;
      RECT 0.0000 37.6000 100.2800 39.2400 ;
      RECT 97.5200 36.5200 100.2800 37.6000 ;
      RECT 4.8600 36.5200 95.4200 37.6000 ;
      RECT 0.0000 36.5200 2.7600 37.6000 ;
      RECT 0.0000 34.8800 100.2800 36.5200 ;
      RECT 95.0200 33.8000 100.2800 34.8800 ;
      RECT 7.3600 33.8000 92.9200 34.8800 ;
      RECT 0.0000 33.8000 5.2600 34.8800 ;
      RECT 0.0000 32.1600 100.2800 33.8000 ;
      RECT 97.5200 31.0800 100.2800 32.1600 ;
      RECT 4.8600 31.0800 95.4200 32.1600 ;
      RECT 0.0000 31.0800 2.7600 32.1600 ;
      RECT 0.0000 29.4400 100.2800 31.0800 ;
      RECT 95.0200 28.3600 100.2800 29.4400 ;
      RECT 7.3600 28.3600 92.9200 29.4400 ;
      RECT 0.0000 28.3600 5.2600 29.4400 ;
      RECT 0.0000 26.7200 100.2800 28.3600 ;
      RECT 97.5200 25.6400 100.2800 26.7200 ;
      RECT 4.8600 25.6400 95.4200 26.7200 ;
      RECT 0.0000 25.6400 2.7600 26.7200 ;
      RECT 0.0000 24.0000 100.2800 25.6400 ;
      RECT 95.0200 22.9200 100.2800 24.0000 ;
      RECT 7.3600 22.9200 92.9200 24.0000 ;
      RECT 0.0000 22.9200 5.2600 24.0000 ;
      RECT 0.0000 21.2800 100.2800 22.9200 ;
      RECT 97.5200 20.2000 100.2800 21.2800 ;
      RECT 4.8600 20.2000 95.4200 21.2800 ;
      RECT 0.0000 20.2000 2.7600 21.2800 ;
      RECT 0.0000 18.5600 100.2800 20.2000 ;
      RECT 95.0200 17.4800 100.2800 18.5600 ;
      RECT 7.3600 17.4800 92.9200 18.5600 ;
      RECT 0.0000 17.4800 5.2600 18.5600 ;
      RECT 0.0000 15.8400 100.2800 17.4800 ;
      RECT 97.5200 14.7600 100.2800 15.8400 ;
      RECT 4.8600 14.7600 95.4200 15.8400 ;
      RECT 0.0000 14.7600 2.7600 15.8400 ;
      RECT 0.0000 13.1200 100.2800 14.7600 ;
      RECT 95.0200 12.0400 100.2800 13.1200 ;
      RECT 7.3600 12.0400 92.9200 13.1200 ;
      RECT 0.0000 12.0400 5.2600 13.1200 ;
      RECT 0.0000 10.4000 100.2800 12.0400 ;
      RECT 97.5200 9.3200 100.2800 10.4000 ;
      RECT 4.8600 9.3200 95.4200 10.4000 ;
      RECT 0.0000 9.3200 2.7600 10.4000 ;
      RECT 0.0000 7.2300 100.2800 9.3200 ;
      RECT 95.0200 5.1300 100.2800 7.2300 ;
      RECT 0.0000 5.1300 5.2600 7.2300 ;
      RECT 0.0000 4.7300 100.2800 5.1300 ;
      RECT 97.5200 2.6300 100.2800 4.7300 ;
      RECT 0.0000 2.6300 2.7600 4.7300 ;
      RECT 0.0000 1.1000 100.2800 2.6300 ;
      RECT 81.1800 0.0000 100.2800 1.1000 ;
      RECT 0.0000 0.0000 80.2800 1.1000 ;
    LAYER met4 ;
      RECT 0.0000 216.3300 100.2800 219.6400 ;
      RECT 4.8600 213.8300 95.4200 216.3300 ;
      RECT 95.0200 5.1300 95.4200 213.8300 ;
      RECT 7.3600 5.1300 92.9200 213.8300 ;
      RECT 4.8600 5.1300 5.2600 213.8300 ;
      RECT 97.5200 2.6300 100.2800 216.3300 ;
      RECT 4.8600 2.6300 95.4200 5.1300 ;
      RECT 0.0000 2.6300 2.7600 216.3300 ;
      RECT 0.0000 0.0000 100.2800 2.6300 ;
  END
END RAM_IO

END LIBRARY
