magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< locali >>
rect 567 1431 601 1447
rect 567 1381 601 1397
rect 567 17 601 33
rect 567 -33 601 -17
<< viali >>
rect 567 1397 601 1431
rect 567 -17 601 17
<< metal1 >>
rect 552 1388 558 1440
rect 610 1388 616 1440
rect 552 -26 558 26
rect 610 -26 616 26
<< via1 >>
rect 558 1431 610 1440
rect 558 1397 567 1431
rect 567 1397 601 1431
rect 601 1397 610 1431
rect 558 1388 610 1397
rect 558 17 610 26
rect 558 -17 567 17
rect 567 -17 601 17
rect 601 -17 610 17
rect 558 -26 610 -17
<< metal2 >>
rect 556 1442 612 1451
rect 137 538 203 590
rect 369 345 397 1414
rect 556 1377 612 1386
rect 1082 609 1148 661
rect 368 336 424 345
rect 368 271 424 280
rect 369 0 397 271
rect 556 28 612 37
rect 556 -37 612 -28
<< via2 >>
rect 556 1440 612 1442
rect 556 1388 558 1440
rect 558 1388 610 1440
rect 610 1388 612 1440
rect 556 1386 612 1388
rect 368 280 424 336
rect 556 26 612 28
rect 556 -26 558 26
rect 558 -26 610 26
rect 610 -26 612 26
rect 556 -28 612 -26
<< metal3 >>
rect 535 1442 633 1463
rect 535 1386 556 1442
rect 612 1386 633 1442
rect 535 1365 633 1386
rect 363 338 429 341
rect 0 336 1168 338
rect 0 280 368 336
rect 424 280 1168 336
rect 0 278 1168 280
rect 363 275 429 278
rect 535 28 633 49
rect 535 -28 556 28
rect 612 -28 633 28
rect 535 -49 633 -28
use contact_7  contact_7_0
timestamp 1707688321
transform 1 0 555 0 1 -33
box 0 0 1 1
use contact_7  contact_7_1
timestamp 1707688321
transform 1 0 555 0 1 1381
box 0 0 1 1
use contact_8  contact_8_0
timestamp 1707688321
transform 1 0 552 0 1 -32
box 0 0 1 1
use contact_8  contact_8_1
timestamp 1707688321
transform 1 0 552 0 1 1382
box 0 0 1 1
use contact_9  contact_9_0
timestamp 1707688321
transform 1 0 363 0 1 271
box 0 0 1 1
use contact_9  contact_9_1
timestamp 1707688321
transform 1 0 551 0 1 -37
box 0 0 1 1
use contact_9  contact_9_2
timestamp 1707688321
transform 1 0 551 0 1 1377
box 0 0 1 1
use dff  dff_0
timestamp 1707688321
transform 1 0 0 0 1 0
box -8 -43 1176 1467
<< labels >>
rlabel metal2 s 170 564 170 564 4 din_0
port 1 nsew
rlabel metal2 s 1115 635 1115 635 4 dout_0
port 2 nsew
rlabel metal3 s 584 0 584 0 4 gnd
port 5 nsew
rlabel metal3 s 584 1414 584 1414 4 vdd
port 4 nsew
rlabel metal3 s 584 308 584 308 4 clk
port 3 nsew
<< properties >>
string FIXED_BBOX 551 -37 617 0
string GDS_END 5302684
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 5301352
<< end >>
