magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -54 139 204 164
rect -59 -29 209 139
rect -54 -54 204 -29
<< scpmos >>
rect 60 0 90 110
<< pdiff >>
rect 0 72 60 110
rect 0 38 8 72
rect 42 38 60 72
rect 0 0 60 38
rect 90 72 150 110
rect 90 38 108 72
rect 142 38 150 72
rect 90 0 150 38
<< pdiffc >>
rect 8 38 42 72
rect 108 38 142 72
<< poly >>
rect 60 110 90 136
rect 60 -26 90 0
<< locali >>
rect 8 72 42 88
rect 8 22 42 38
rect 108 72 142 88
rect 108 22 142 38
use contact_11  contact_11_0
timestamp 1707688321
transform 1 0 100 0 1 22
box 0 0 1 1
use contact_11  contact_11_1
timestamp 1707688321
transform 1 0 0 0 1 22
box 0 0 1 1
<< labels >>
rlabel locali s 125 55 125 55 4 D
port 1 nsew
rlabel locali s 25 55 25 55 4 S
port 2 nsew
rlabel poly s 75 55 75 55 4 G
port 3 nsew
<< properties >>
string FIXED_BBOX -54 -54 204 -29
string GDS_END 37124
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 36308
<< end >>
