magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -84 2850 139 3672
rect 8029 2850 8341 3672
rect 169 557 529 778
rect -53 -8 529 557
<< pwell >>
rect -43 2702 124 2790
rect 9427 2702 9507 2790
rect -43 1248 44 2702
rect -43 617 43 896
<< psubdiff >>
rect -17 820 17 870
rect -17 701 17 786
rect -17 643 17 667
<< nsubdiff >>
rect -17 497 17 521
rect -17 429 17 463
rect -17 361 17 395
rect -17 293 17 327
rect -17 224 17 259
rect -17 155 17 190
rect -17 86 17 121
rect 17 52 56 62
rect -17 28 56 52
rect 90 28 129 62
rect 163 28 201 62
rect 235 28 259 62
<< mvpsubdiff >>
rect -17 2728 98 2764
rect 9453 2728 9481 2764
rect -17 2720 18 2728
rect 17 2686 18 2720
rect -17 2650 18 2686
rect 17 2616 18 2650
rect -17 2582 18 2616
rect 17 2548 18 2582
rect -17 2514 18 2548
rect 17 2480 18 2514
rect -17 2378 18 2480
rect 17 2344 18 2378
rect -17 2309 18 2344
rect 17 2275 18 2309
rect -17 2240 18 2275
rect 17 2206 18 2240
rect -17 2171 18 2206
rect 17 2137 18 2171
rect -17 2102 18 2137
rect 17 2068 18 2102
rect -17 2032 18 2068
rect 17 1998 18 2032
rect -17 1962 18 1998
rect 17 1928 18 1962
rect -17 1892 18 1928
rect 17 1858 18 1892
rect -17 1822 18 1858
rect 17 1788 18 1822
rect -17 1752 18 1788
rect 17 1718 18 1752
rect -17 1682 18 1718
rect 17 1648 18 1682
rect -17 1612 18 1648
rect 17 1578 18 1612
rect -17 1542 18 1578
rect 17 1508 18 1542
rect -17 1472 18 1508
rect 17 1438 18 1472
rect -17 1402 18 1438
rect 17 1368 18 1402
rect -17 1332 18 1368
rect 17 1298 18 1332
rect -17 1274 18 1298
<< mvnsubdiff >>
rect -17 3522 18 3606
rect 17 3488 18 3522
rect -17 3454 18 3488
rect 17 3420 18 3454
rect -17 3386 18 3420
rect 17 3352 18 3386
rect -17 3318 18 3352
rect 17 3284 18 3318
rect -17 3248 18 3284
rect 17 3214 18 3248
rect -17 3180 18 3214
rect 17 3146 18 3180
rect -17 3112 18 3146
rect 17 3078 18 3112
rect -17 3044 18 3078
rect 17 3010 18 3044
rect -17 2974 18 3010
rect 17 2952 18 2974
rect 17 2940 113 2952
rect -17 2916 113 2940
rect 9453 2916 9481 2952
<< psubdiffcont >>
rect -17 786 17 820
rect -17 667 17 701
<< nsubdiffcont >>
rect -17 463 17 497
rect -17 395 17 429
rect -17 327 17 361
rect -17 259 17 293
rect -17 190 17 224
rect -17 121 17 155
rect -17 52 17 86
rect 56 28 90 62
rect 129 28 163 62
rect 201 28 235 62
<< mvpsubdiffcont >>
rect -17 2686 17 2720
rect -17 2616 17 2650
rect -17 2548 17 2582
rect -17 2480 17 2514
rect -17 2344 17 2378
rect -17 2275 17 2309
rect -17 2206 17 2240
rect -17 2137 17 2171
rect -17 2068 17 2102
rect -17 1998 17 2032
rect -17 1928 17 1962
rect -17 1858 17 1892
rect -17 1788 17 1822
rect -17 1718 17 1752
rect -17 1648 17 1682
rect -17 1578 17 1612
rect -17 1508 17 1542
rect -17 1438 17 1472
rect -17 1368 17 1402
rect -17 1298 17 1332
<< mvnsubdiffcont >>
rect -17 3488 17 3522
rect -17 3420 17 3454
rect -17 3352 17 3386
rect -17 3284 17 3318
rect -17 3214 17 3248
rect -17 3146 17 3180
rect -17 3078 17 3112
rect -17 3010 17 3044
rect -17 2940 17 2974
<< locali >>
rect 2666 3698 2704 3732
rect 2401 3624 2439 3658
rect -17 3522 17 3604
rect 1555 3544 1593 3578
rect -17 3454 17 3488
rect 223 3464 257 3502
rect 643 3430 677 3468
rect -17 3386 17 3420
rect 1947 3432 1981 3470
rect 2653 3430 2727 3698
rect 4577 3624 4615 3658
rect 5796 3639 5901 3704
rect 6201 3654 6235 3704
rect 6904 3639 6991 3704
rect 9604 3698 9642 3732
rect 9676 3698 9757 3704
rect 9668 3638 9757 3698
rect 10754 3638 10875 3704
rect 5019 3544 5057 3578
rect 5473 3555 5507 3604
rect 7277 3555 7311 3604
rect 6362 3504 6396 3542
rect 7631 3504 7665 3542
rect 8839 3556 8873 3605
rect 10061 3555 10095 3604
rect 10413 3555 10447 3604
rect 7739 3504 7773 3542
rect 10849 3470 10887 3504
rect 7847 3430 7881 3468
rect 2687 3396 2727 3430
rect -17 3318 17 3352
rect 2653 3358 2727 3396
rect -17 3248 17 3284
rect 563 3272 597 3310
rect 1003 3272 1037 3310
rect 1212 3278 1246 3316
rect 2687 3324 2727 3358
rect 2869 3358 2903 3396
rect 2231 3272 2265 3310
rect 8752 3278 8786 3316
rect 3147 3238 3185 3272
rect 4241 3238 4279 3272
rect 8932 3278 8966 3316
rect 9953 3278 9987 3316
rect 10521 3278 10555 3316
rect -17 3180 17 3214
rect -17 3112 17 3146
rect -17 3044 17 3078
rect -17 2974 17 3010
rect 17 2934 55 2968
rect -17 2902 17 2934
rect 10989 2902 11096 2968
rect 115 2820 149 2858
rect 745 2860 783 2894
rect 1841 2860 1879 2894
rect 5927 2860 5965 2894
rect 6707 2860 6745 2894
rect 6779 2860 6817 2894
rect 291 2820 325 2858
rect 2067 2812 2105 2846
rect 5107 2822 5141 2860
rect 6533 2812 6571 2846
rect 7153 2812 7191 2846
rect 8485 2820 8519 2858
rect -17 2746 17 2784
rect 10997 2712 11120 2778
rect -17 2650 17 2686
rect -17 2582 17 2616
rect -17 2514 17 2548
rect -17 2378 17 2480
rect 6001 2450 6077 2484
rect 361 2404 399 2438
rect 1374 2398 1412 2432
rect 3377 2378 3415 2412
rect 4010 2378 4048 2412
rect 5191 2378 5229 2412
rect 6043 2407 6077 2450
rect 5558 2373 5596 2407
rect 6049 2373 6087 2407
rect -17 2309 17 2344
rect -17 2240 17 2275
rect 233 2254 267 2288
rect 421 2264 459 2298
rect 735 2254 769 2288
rect -17 2171 17 2206
rect -17 2102 17 2137
rect -17 2032 17 2068
rect -17 1972 17 1998
rect -17 1900 17 1928
rect -17 1828 17 1858
rect -17 1756 17 1788
rect -17 1684 17 1718
rect -17 1612 17 1648
rect -17 1542 17 1578
rect -17 1472 17 1508
rect -17 1402 17 1438
rect -17 1332 17 1368
rect -17 1274 17 1291
rect -17 823 17 870
rect -17 751 17 786
rect -17 701 17 717
rect -17 643 17 645
rect -17 497 17 521
rect -17 429 17 463
rect -17 361 17 395
rect -17 293 17 327
rect -17 224 17 259
rect -17 155 17 190
rect -17 86 17 121
rect -17 28 17 52
rect 32 28 56 62
rect 90 28 129 62
rect 163 28 201 62
rect 235 28 259 62
<< viali >>
rect 2632 3698 2666 3732
rect 2704 3698 2738 3732
rect 2367 3624 2401 3658
rect 2439 3624 2473 3658
rect 1521 3544 1555 3578
rect 1593 3544 1627 3578
rect 223 3502 257 3536
rect 223 3430 257 3464
rect 643 3468 677 3502
rect 643 3396 677 3430
rect 1947 3470 1981 3504
rect 1947 3398 1981 3432
rect 4543 3624 4577 3658
rect 4615 3624 4649 3658
rect 9570 3698 9604 3732
rect 9642 3698 9676 3732
rect 9294 3622 9328 3656
rect 4985 3544 5019 3578
rect 5057 3544 5091 3578
rect 6362 3542 6396 3576
rect 6362 3470 6396 3504
rect 7631 3542 7665 3576
rect 7631 3470 7665 3504
rect 7739 3542 7773 3576
rect 7739 3470 7773 3504
rect 7847 3468 7881 3502
rect 10815 3470 10849 3504
rect 10887 3470 10921 3504
rect 2653 3396 2687 3430
rect 563 3310 597 3344
rect 563 3238 597 3272
rect 1003 3310 1037 3344
rect 1003 3238 1037 3272
rect 1212 3316 1246 3350
rect 1212 3244 1246 3278
rect 2231 3310 2265 3344
rect 2653 3324 2687 3358
rect 2869 3396 2903 3430
rect 7847 3396 7881 3430
rect 9107 3396 9141 3430
rect 2869 3324 2903 3358
rect 4015 3320 4049 3354
rect 8752 3316 8786 3350
rect 2231 3238 2265 3272
rect 3113 3238 3147 3272
rect 3185 3238 3219 3272
rect 4207 3238 4241 3272
rect 4279 3238 4313 3272
rect 8752 3244 8786 3278
rect 8932 3316 8966 3350
rect 8932 3244 8966 3278
rect 9953 3316 9987 3350
rect 9953 3244 9987 3278
rect 10521 3316 10555 3350
rect 10521 3244 10555 3278
rect -17 2940 17 2968
rect -17 2934 17 2940
rect 55 2934 89 2968
rect 115 2858 149 2892
rect -17 2784 17 2818
rect 115 2786 149 2820
rect 291 2858 325 2892
rect 711 2860 745 2894
rect 783 2860 817 2894
rect 1807 2860 1841 2894
rect 1879 2860 1913 2894
rect 5107 2860 5141 2894
rect 5893 2860 5927 2894
rect 5965 2860 5999 2894
rect 6673 2860 6707 2894
rect 6745 2860 6779 2894
rect 6817 2860 6851 2894
rect 291 2786 325 2820
rect 2033 2812 2067 2846
rect 2105 2812 2139 2846
rect 8485 2858 8519 2892
rect 5107 2788 5141 2822
rect 6499 2812 6533 2846
rect 6571 2812 6605 2846
rect 7119 2812 7153 2846
rect 7191 2812 7225 2846
rect 8485 2786 8519 2820
rect -17 2720 17 2746
rect -17 2712 17 2720
rect 327 2404 361 2438
rect 399 2404 433 2438
rect 1340 2398 1374 2432
rect 1412 2398 1446 2432
rect 3343 2378 3377 2412
rect 3415 2378 3449 2412
rect 3976 2378 4010 2412
rect 4048 2378 4082 2412
rect 5157 2378 5191 2412
rect 5229 2378 5263 2412
rect 5524 2373 5558 2407
rect 5596 2373 5630 2407
rect 6015 2373 6049 2407
rect 6087 2373 6121 2407
rect 387 2264 421 2298
rect 459 2264 493 2298
rect -17 1962 17 1972
rect -17 1938 17 1962
rect -17 1892 17 1900
rect -17 1866 17 1892
rect -17 1822 17 1828
rect -17 1794 17 1822
rect -17 1752 17 1756
rect -17 1722 17 1752
rect -17 1682 17 1684
rect -17 1650 17 1682
rect -17 1578 17 1612
rect -17 1298 17 1325
rect -17 1291 17 1298
rect -17 820 17 823
rect -17 789 17 820
rect -17 717 17 751
rect -17 667 17 679
rect -17 645 17 667
<< metal1 >>
rect 2620 3732 9688 3738
rect 2620 3698 2632 3732
rect 2666 3698 2704 3732
rect 2738 3698 9570 3732
rect 9604 3698 9642 3732
rect 9676 3698 9688 3732
rect 2620 3692 9688 3698
rect 2355 3662 6433 3664
tri 6433 3662 6435 3664 sw
rect 2355 3658 6435 3662
rect 2355 3624 2367 3658
rect 2401 3624 2439 3658
rect 2473 3624 4543 3658
rect 4577 3624 4615 3658
rect 4649 3656 6435 3658
tri 6435 3656 6441 3662 sw
tri 8344 3656 8350 3662 se
rect 8350 3656 9345 3662
rect 4649 3654 6441 3656
tri 6441 3654 6443 3656 sw
tri 8342 3654 8344 3656 se
rect 4649 3642 6443 3654
tri 6443 3642 6455 3654 sw
rect 4649 3624 6455 3642
rect 2355 3622 6455 3624
tri 6455 3622 6475 3642 sw
rect 2355 3618 6475 3622
tri 6475 3618 6479 3622 sw
tri 6413 3584 6447 3618 ne
rect 6447 3584 6479 3618
tri 6479 3584 6513 3618 sw
rect 7619 3610 8292 3654
rect 211 3578 5103 3584
tri 6447 3582 6449 3584 ne
rect 6449 3582 6513 3584
tri 6513 3582 6515 3584 sw
rect 211 3544 1521 3578
rect 1555 3544 1593 3578
rect 1627 3544 4985 3578
rect 5019 3544 5057 3578
rect 5091 3544 5103 3578
rect 211 3538 5103 3544
rect 6350 3576 6408 3582
tri 6449 3576 6455 3582 ne
rect 6455 3576 6515 3582
tri 6515 3576 6521 3582 sw
rect 7619 3576 7677 3610
tri 7677 3585 7702 3610 nw
tri 8261 3585 8286 3610 ne
rect 8286 3602 8292 3610
rect 8344 3622 9294 3656
rect 9328 3622 9345 3656
rect 8344 3616 9345 3622
rect 8344 3602 8350 3616
rect 8286 3590 8350 3602
rect 6350 3542 6362 3576
rect 6396 3542 6408 3576
tri 6455 3542 6489 3576 ne
rect 6489 3542 6521 3576
tri 6521 3542 6555 3576 sw
rect 7619 3542 7631 3576
rect 7665 3542 7677 3576
rect 211 3536 291 3538
rect 211 3502 223 3536
rect 257 3535 291 3536
tri 291 3535 294 3538 nw
rect 257 3502 269 3535
tri 269 3513 291 3535 nw
tri 6328 3513 6350 3535 se
rect 6350 3513 6408 3542
tri 6325 3510 6328 3513 se
rect 6328 3510 6408 3513
tri 6489 3510 6521 3542 ne
rect 6521 3510 6555 3542
tri 6555 3510 6587 3542 sw
tri 7594 3510 7619 3535 se
rect 7619 3510 7677 3542
rect 211 3464 269 3502
rect 211 3430 223 3464
rect 257 3430 269 3464
rect 211 3424 269 3430
rect 631 3502 689 3508
rect 631 3468 643 3502
rect 677 3470 689 3502
rect 1935 3504 6408 3510
tri 6521 3504 6527 3510 ne
rect 6527 3504 7677 3510
tri 689 3470 692 3473 sw
rect 1935 3470 1947 3504
rect 1981 3470 6362 3504
rect 6396 3470 6408 3504
tri 6527 3470 6561 3504 ne
rect 6561 3470 7631 3504
rect 7665 3470 7677 3504
rect 677 3468 692 3470
tri 692 3468 694 3470 sw
rect 631 3448 694 3468
tri 694 3448 714 3468 sw
rect 1935 3464 6408 3470
tri 6561 3468 6563 3470 ne
rect 6563 3468 7677 3470
tri 6563 3464 6567 3468 ne
rect 6567 3464 7677 3468
rect 7727 3576 7927 3582
tri 7927 3576 7933 3582 sw
rect 7727 3542 7739 3576
rect 7773 3542 7933 3576
rect 7727 3538 7933 3542
tri 7933 3538 7971 3576 sw
rect 8286 3538 8292 3590
rect 8344 3538 8350 3590
tri 8350 3582 8384 3616 nw
rect 7727 3536 7971 3538
tri 7971 3536 7973 3538 sw
rect 7727 3504 7785 3536
tri 7785 3511 7810 3536 nw
tri 7907 3511 7932 3536 ne
rect 7932 3511 7973 3536
tri 7973 3511 7998 3536 sw
tri 7932 3510 7933 3511 ne
rect 7933 3510 7998 3511
tri 7998 3510 7999 3511 sw
tri 7933 3508 7935 3510 ne
rect 7935 3508 10933 3510
rect 7727 3470 7739 3504
rect 7773 3470 7785 3504
rect 7727 3464 7785 3470
rect 7835 3502 7893 3508
tri 7935 3504 7939 3508 ne
rect 7939 3504 10933 3508
rect 7835 3468 7847 3502
rect 7881 3468 7893 3502
tri 7939 3470 7973 3504 ne
rect 7973 3470 10815 3504
rect 10849 3470 10887 3504
rect 10921 3470 10933 3504
rect 1935 3461 2015 3464
tri 2015 3461 2018 3464 nw
rect 631 3432 1822 3448
tri 1822 3432 1838 3448 sw
rect 1935 3432 1993 3461
tri 1993 3439 2015 3461 nw
tri 7813 3439 7835 3461 se
rect 7835 3439 7893 3468
tri 7973 3464 7979 3470 ne
rect 7979 3464 9325 3470
tri 9325 3464 9331 3470 nw
tri 10119 3464 10125 3470 ne
rect 10125 3464 10933 3470
tri 7810 3436 7813 3439 se
rect 7813 3436 7893 3439
tri 7893 3436 7918 3461 sw
rect 631 3430 1838 3432
rect 631 3396 643 3430
rect 677 3398 1838 3430
tri 1838 3398 1872 3432 sw
rect 1935 3398 1947 3432
rect 1981 3398 1993 3432
tri 2148 3430 2154 3436 se
rect 2154 3430 2699 3436
rect 677 3396 1872 3398
tri 1872 3396 1874 3398 sw
rect 631 3392 1874 3396
tri 1874 3392 1878 3396 sw
rect 1935 3392 1993 3398
tri 2114 3396 2148 3430 se
rect 2148 3396 2653 3430
rect 2687 3396 2699 3430
tri 2110 3392 2114 3396 se
rect 2114 3392 2699 3396
rect 631 3390 1878 3392
tri 1878 3390 1880 3392 sw
tri 2108 3390 2110 3392 se
rect 2110 3390 2699 3392
tri 1798 3362 1826 3390 ne
rect 1826 3378 1880 3390
tri 1880 3378 1892 3390 sw
tri 2096 3378 2108 3390 se
rect 2108 3378 2699 3390
rect 1826 3362 1892 3378
rect 1206 3350 1465 3362
tri 1826 3358 1830 3362 ne
rect 1830 3359 1892 3362
tri 1892 3359 1911 3378 sw
tri 2077 3359 2096 3378 se
rect 2096 3359 2159 3378
tri 2159 3359 2178 3378 nw
tri 2616 3359 2635 3378 ne
rect 2635 3359 2699 3378
rect 1830 3358 1911 3359
tri 1911 3358 1912 3359 sw
tri 2076 3358 2077 3359 se
rect 2077 3358 2158 3359
tri 2158 3358 2159 3359 nw
tri 2635 3358 2636 3359 ne
rect 2636 3358 2699 3359
tri 1830 3350 1838 3358 ne
rect 1838 3350 1912 3358
rect 551 3344 609 3350
rect 551 3310 563 3344
rect 597 3310 609 3344
rect 991 3344 1049 3350
tri 609 3310 614 3315 sw
tri 986 3310 991 3315 se
rect 991 3310 1003 3344
rect 1037 3310 1049 3344
rect 551 3290 614 3310
tri 614 3290 634 3310 sw
tri 966 3290 986 3310 se
rect 986 3290 1049 3310
rect 551 3272 1049 3290
rect 551 3238 563 3272
rect 597 3238 1003 3272
rect 1037 3238 1049 3272
rect 551 3232 1049 3238
rect 1206 3316 1212 3350
rect 1246 3316 1465 3350
tri 1838 3344 1844 3350 ne
rect 1844 3344 1912 3350
tri 1912 3344 1926 3358 sw
tri 2062 3344 2076 3358 se
rect 2076 3350 2150 3358
tri 2150 3350 2158 3358 nw
tri 2636 3353 2641 3358 ne
rect 2076 3344 2144 3350
tri 2144 3344 2150 3350 nw
rect 2219 3344 2277 3350
rect 1206 3278 1465 3316
tri 1844 3310 1878 3344 ne
rect 1878 3335 1926 3344
tri 1926 3335 1935 3344 sw
tri 2053 3335 2062 3344 se
rect 2062 3335 2110 3344
rect 1878 3310 2110 3335
tri 2110 3310 2144 3344 nw
rect 2219 3310 2231 3344
rect 2265 3310 2277 3344
rect 2641 3324 2653 3358
rect 2687 3324 2699 3358
rect 2641 3318 2699 3324
rect 2857 3430 9172 3436
rect 2857 3396 2869 3430
rect 2903 3396 7847 3430
rect 7881 3396 9107 3430
rect 9141 3396 9172 3430
rect 2857 3390 9172 3396
rect 2857 3358 2915 3390
tri 2915 3365 2940 3390 nw
rect 2857 3324 2869 3358
rect 2903 3324 2915 3358
rect 2857 3318 2915 3324
rect 4003 3354 5670 3360
rect 4003 3320 4015 3354
rect 4049 3352 5670 3354
tri 5670 3352 5678 3360 sw
rect 8746 3352 8792 3362
rect 4049 3350 8792 3352
rect 4049 3321 8752 3350
rect 4049 3320 4064 3321
rect 4003 3316 4064 3320
tri 4064 3316 4069 3321 nw
tri 5649 3316 5654 3321 ne
rect 5654 3316 8752 3321
rect 8786 3316 8792 3350
rect 4003 3314 4062 3316
tri 4062 3314 4064 3316 nw
tri 5654 3314 5656 3316 ne
rect 5656 3314 8792 3316
tri 1878 3308 1880 3310 ne
rect 1880 3308 2108 3310
tri 2108 3308 2110 3310 nw
tri 1880 3278 1910 3308 ne
rect 1910 3278 2078 3308
tri 2078 3278 2108 3308 nw
rect 2219 3284 2277 3310
tri 5656 3306 5664 3314 ne
rect 5664 3306 8792 3314
tri 2277 3284 2296 3303 sw
rect 2219 3278 2296 3284
tri 2296 3278 2302 3284 sw
rect 1206 3244 1212 3278
rect 1246 3244 1465 3278
tri 1910 3277 1911 3278 ne
rect 1911 3277 2077 3278
tri 2077 3277 2078 3278 nw
rect 1206 3232 1465 3244
rect 2219 3272 3231 3278
rect 2219 3238 2231 3272
rect 2265 3238 3113 3272
rect 3147 3238 3185 3272
rect 3219 3238 3231 3272
rect 2219 3232 3231 3238
rect 4195 3272 4761 3284
rect 4195 3238 4207 3272
rect 4241 3238 4279 3272
rect 4313 3238 4761 3272
rect 4195 3232 4761 3238
rect 4813 3232 4825 3284
rect 4877 3232 4883 3284
rect 8746 3278 8792 3306
rect 8746 3244 8752 3278
rect 8786 3244 8792 3278
rect 8746 3232 8792 3244
rect 8915 3350 9199 3362
rect 8915 3316 8932 3350
rect 8966 3316 9199 3350
rect 8915 3278 9199 3316
rect 8915 3244 8932 3278
rect 8966 3244 9199 3278
rect 8915 3232 9199 3244
rect 9735 3350 9993 3362
rect 9735 3316 9953 3350
rect 9987 3316 9993 3350
rect 9735 3278 9993 3316
rect 9735 3244 9953 3278
rect 9987 3244 9993 3278
rect 9735 3232 9993 3244
rect 10515 3350 10773 3362
rect 10515 3316 10521 3350
rect 10555 3316 10773 3350
rect 10515 3278 10773 3316
rect 10515 3244 10521 3278
rect 10555 3244 10773 3278
rect 10515 3232 10773 3244
rect -29 3002 154 3204
rect 836 3002 946 3204
rect 1678 3002 1788 3204
rect 2492 3002 2602 3204
rect 3658 3002 3768 3204
rect 4824 3002 4934 3204
rect 6018 3002 6128 3204
rect 6656 3002 6766 3204
rect 7499 3002 8386 3204
rect 8570 3002 8680 3204
rect 9412 3002 9522 3204
rect -29 2974 11132 3002
rect -29 2968 154 2974
rect -29 2934 -17 2968
rect 17 2934 55 2968
rect 89 2934 154 2968
rect -29 2928 154 2934
rect 836 2928 946 2974
rect 1678 2928 1788 2974
rect 2492 2928 2602 2974
rect 3658 2928 3768 2974
rect 4824 2928 4934 2974
rect 6018 2928 6128 2974
rect 6656 2928 6766 2974
rect 7499 2928 8383 2974
rect 8570 2928 8680 2974
rect 9412 2928 9522 2974
rect 103 2894 829 2900
tri 1194 2894 1200 2900 se
rect 1200 2894 1925 2900
rect 103 2892 711 2894
rect 103 2858 115 2892
rect 149 2858 291 2892
rect 325 2860 711 2892
rect 745 2860 783 2894
rect 817 2860 829 2894
tri 1160 2860 1194 2894 se
rect 1194 2860 1807 2894
rect 1841 2860 1879 2894
rect 1913 2860 1925 2894
rect 325 2858 829 2860
tri 1158 2858 1160 2860 se
rect 1160 2858 1925 2860
rect 103 2854 829 2858
tri 1154 2854 1158 2858 se
rect 1158 2854 1925 2858
rect 5095 2894 6011 2900
rect 5095 2860 5107 2894
rect 5141 2860 5893 2894
rect 5927 2860 5965 2894
rect 5999 2860 6011 2894
rect 5095 2854 6011 2860
rect 6661 2894 6863 2900
rect 6661 2860 6673 2894
rect 6707 2860 6745 2894
rect 6779 2860 6817 2894
rect 6851 2860 6863 2894
rect 6661 2854 6863 2860
rect 8473 2892 8531 2898
rect 8473 2858 8485 2892
rect 8519 2858 8531 2892
rect 103 2852 429 2854
tri 429 2852 431 2854 nw
tri 1152 2852 1154 2854 se
rect 1154 2852 1218 2854
tri 1218 2852 1220 2854 nw
rect 5095 2852 5176 2854
tri 5176 2852 5178 2854 nw
rect 103 2846 423 2852
tri 423 2846 429 2852 nw
tri 1151 2851 1152 2852 se
rect 1152 2851 1212 2852
tri 1146 2846 1151 2851 se
rect 1151 2846 1212 2851
tri 1212 2846 1218 2852 nw
rect 2021 2846 2287 2852
tri 2287 2846 2293 2852 sw
rect 5095 2846 5170 2852
tri 5170 2846 5176 2852 nw
tri 6327 2846 6333 2852 se
rect 6333 2846 6617 2852
tri 6965 2846 6971 2852 se
rect 6971 2846 7237 2852
rect 103 2826 403 2846
tri 403 2826 423 2846 nw
tri 1134 2834 1146 2846 se
rect 1146 2834 1200 2846
tri 1200 2834 1212 2846 nw
tri 1126 2826 1134 2834 se
rect 1134 2826 1192 2834
tri 1192 2826 1200 2834 nw
rect -29 2818 29 2824
rect -29 2784 -17 2818
rect 17 2784 29 2818
tri -54 2752 -29 2777 se
rect -29 2752 29 2784
rect 103 2822 399 2826
tri 399 2822 403 2826 nw
tri 1122 2822 1126 2826 se
rect 1126 2822 1188 2826
tri 1188 2822 1192 2826 nw
rect 103 2820 389 2822
rect 103 2786 115 2820
rect 149 2809 291 2820
rect 149 2786 161 2809
rect 103 2780 161 2786
rect 279 2786 291 2809
rect 325 2812 389 2820
tri 389 2812 399 2822 nw
tri 1113 2813 1122 2822 se
rect 1122 2813 1179 2822
tri 1179 2813 1188 2822 nw
rect 1113 2812 1178 2813
tri 1178 2812 1179 2813 nw
rect 325 2809 386 2812
tri 386 2809 389 2812 nw
tri 1113 2809 1116 2812 ne
rect 1116 2809 1154 2812
rect 325 2788 365 2809
tri 365 2788 386 2809 nw
tri 1116 2788 1137 2809 ne
rect 1137 2788 1154 2809
tri 1154 2788 1178 2812 nw
rect 325 2786 363 2788
tri 363 2786 365 2788 nw
tri 1137 2786 1139 2788 ne
rect 1139 2786 1152 2788
tri 1152 2786 1154 2788 nw
rect 279 2780 357 2786
tri 357 2780 363 2786 nw
tri 1139 2780 1145 2786 ne
rect 1145 2780 1146 2786
tri 1146 2780 1152 2786 nw
tri 29 2752 54 2777 sw
tri 1419 2752 1444 2777 se
rect -54 2746 154 2752
rect -54 2712 -17 2746
rect 17 2712 154 2746
rect -54 2706 154 2712
rect 836 2706 946 2752
rect 1444 2706 1450 2822
rect 1566 2706 1572 2822
rect 2021 2812 2033 2846
rect 2067 2812 2105 2846
rect 2139 2826 2293 2846
tri 2293 2826 2313 2846 sw
rect 2139 2812 2287 2826
rect 2021 2806 2287 2812
tri 2261 2788 2279 2806 ne
rect 2279 2788 2287 2806
tri 2279 2786 2281 2788 ne
rect 2281 2786 2287 2788
tri 2281 2782 2285 2786 ne
rect 2285 2782 2287 2786
rect 5095 2822 5153 2846
tri 5153 2829 5170 2846 nw
tri 6310 2829 6327 2846 se
rect 6327 2829 6499 2846
tri 6307 2826 6310 2829 se
rect 6310 2826 6499 2829
rect 5095 2788 5107 2822
rect 5141 2788 5153 2822
rect 5095 2782 5153 2788
rect 6333 2812 6499 2826
rect 6533 2812 6571 2846
rect 6605 2812 6617 2846
tri 6945 2826 6965 2846 se
rect 6965 2826 7119 2846
rect 6333 2806 6617 2812
rect 6971 2812 7119 2826
rect 7153 2812 7191 2846
rect 7225 2812 7237 2846
rect 6971 2806 7237 2812
rect 8473 2826 8531 2858
tri 8531 2826 8556 2851 sw
rect 8473 2820 8651 2826
rect 6333 2786 6339 2806
tri 6339 2786 6359 2806 nw
rect 6971 2786 6977 2806
tri 6977 2786 6997 2806 nw
rect 8473 2786 8485 2820
rect 8519 2786 8651 2820
rect 6333 2782 6335 2786
tri 6335 2782 6339 2786 nw
rect 6971 2782 6973 2786
tri 6973 2782 6977 2786 nw
tri 2285 2780 2287 2782 ne
tri 6333 2780 6335 2782 nw
tri 6971 2780 6973 2782 nw
rect 8473 2780 8651 2786
tri 1572 2752 1597 2777 sw
rect 1678 2706 1788 2752
rect 2492 2706 2602 2752
rect 3658 2706 3768 2752
rect 4824 2706 4934 2752
rect 6018 2706 6128 2752
rect 6656 2706 6766 2752
rect 7499 2706 8415 2752
rect 8570 2706 8680 2752
rect 9412 2706 9522 2752
rect -29 2476 154 2678
rect 530 2476 536 2656
rect 652 2476 658 2656
rect 836 2476 946 2678
rect 1678 2476 1788 2678
rect 2492 2476 2602 2678
rect 3658 2476 3768 2678
rect 4824 2476 4934 2678
rect 6018 2476 6128 2678
rect 6656 2476 6766 2678
rect 7499 2476 8383 2678
rect 8570 2476 8680 2678
rect 9412 2476 9522 2678
rect 315 2438 1288 2444
tri 1288 2438 1294 2444 sw
rect 315 2404 327 2438
rect 361 2404 399 2438
rect 433 2432 1458 2438
rect 433 2404 1340 2432
rect 315 2398 1340 2404
rect 1374 2398 1412 2432
rect 1446 2398 1458 2432
tri 1268 2392 1274 2398 ne
rect 1274 2392 1458 2398
rect 3331 2412 4094 2418
rect 3331 2378 3343 2412
rect 3377 2378 3415 2412
rect 3449 2378 3976 2412
rect 4010 2378 4048 2412
rect 4082 2378 4094 2412
rect 3331 2372 4094 2378
rect 4831 2366 4837 2418
rect 4889 2366 4901 2418
rect 4953 2412 5275 2418
rect 4953 2378 5157 2412
rect 5191 2378 5229 2412
rect 5263 2378 5275 2412
rect 4953 2366 5275 2378
rect 5512 2407 6133 2413
rect 5512 2373 5524 2407
rect 5558 2373 5596 2407
rect 5630 2373 6015 2407
rect 6049 2373 6087 2407
rect 6121 2373 6133 2407
rect 5512 2367 6133 2373
rect 375 2298 536 2304
rect 375 2264 387 2298
rect 421 2264 459 2298
rect 493 2264 536 2298
rect 375 2252 536 2264
rect 588 2252 600 2304
rect 652 2252 658 2304
rect 2085 2012 2125 2214
rect -51 1972 106 1984
rect -51 1938 -17 1972
rect 17 1938 106 1972
rect -51 1900 106 1938
rect -51 1866 -17 1900
rect 17 1866 106 1900
rect -51 1854 106 1866
rect 1444 1864 1450 1980
rect 1566 1864 1572 1980
rect 2102 1854 2125 1984
tri -51 1829 -26 1854 ne
rect -23 1828 23 1854
tri 26 1829 51 1854 nw
rect -23 1794 -17 1828
rect 17 1794 23 1828
rect -23 1756 23 1794
rect -23 1722 -17 1756
rect 17 1722 23 1756
rect -23 1684 23 1722
rect -23 1650 -17 1684
rect 17 1650 23 1684
rect -23 1612 23 1650
rect -23 1578 -17 1612
rect 17 1578 23 1612
tri -51 1415 -26 1440 se
rect -23 1415 23 1578
rect 542 1639 658 1645
rect 1747 1607 1781 1641
rect 542 1517 658 1523
tri 26 1415 51 1440 sw
rect -51 1363 53 1415
tri -51 1338 -26 1363 ne
rect -23 1325 23 1363
tri 26 1338 51 1363 nw
rect -23 1291 -17 1325
rect 17 1291 23 1325
rect -23 1201 23 1291
rect 99 1221 133 1255
tri -51 1145 -26 1170 se
tri 26 1145 51 1170 sw
rect -51 1093 51 1145
rect 542 1055 658 1061
rect 542 869 658 875
rect 2102 863 2125 1065
rect -26 824 26 835
rect 1873 795 1907 829
rect -26 760 26 772
rect -26 696 26 708
rect -26 633 26 644
rect 2074 218 2097 420
rect 2102 72 2125 190
<< via1 >>
rect 8292 3602 8344 3654
rect 8292 3538 8344 3590
rect 4761 3232 4813 3284
rect 4825 3232 4877 3284
rect 1450 2706 1566 2822
rect 536 2476 652 2656
rect 4837 2366 4889 2418
rect 4901 2366 4953 2418
rect 536 2252 588 2304
rect 600 2252 652 2304
rect 1450 1864 1566 1980
rect 542 1523 658 1639
rect 542 875 658 1055
rect -26 823 26 824
rect -26 789 -17 823
rect -17 789 17 823
rect 17 789 26 823
rect -26 772 26 789
rect -26 751 26 760
rect -26 717 -17 751
rect -17 717 17 751
rect 17 717 26 751
rect -26 708 26 717
rect -26 679 26 696
rect -26 645 -17 679
rect -17 645 17 679
rect 17 645 26 679
rect -26 644 26 645
<< metal2 >>
rect 8286 3602 8292 3654
rect 8344 3602 8350 3654
rect 8286 3590 8350 3602
rect 8286 3538 8292 3590
rect 8344 3538 8350 3590
rect 4755 3232 4761 3284
rect 4813 3232 4825 3284
rect 4877 3232 4883 3284
rect 1444 2706 1450 2822
rect 1566 2706 1572 2822
rect 530 2476 536 2656
rect 652 2476 658 2656
rect 530 2304 658 2476
rect 530 2252 536 2304
rect 588 2252 600 2304
rect 652 2252 658 2304
rect -26 824 26 1978
rect 530 1639 658 2252
rect 1444 1980 1572 2706
rect 1600 2214 1856 3010
rect 4755 2418 4883 3232
tri 4883 2418 4908 2443 sw
rect 4755 2366 4837 2418
rect 4889 2366 4901 2418
rect 4953 2366 4959 2418
rect 1444 1864 1450 1980
rect 1566 1864 1572 1980
rect 530 1523 542 1639
rect 530 1055 658 1523
rect 1461 1220 1491 1250
rect 530 875 542 1055
rect 530 869 658 875
rect -26 760 26 772
rect -26 696 26 708
rect -26 638 26 644
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1707688321
transform -1 0 7773 0 1 3470
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_1
timestamp 1707688321
transform -1 0 597 0 1 3238
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_2
timestamp 1707688321
transform -1 0 257 0 1 3430
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_3
timestamp 1707688321
transform -1 0 1981 0 1 3398
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_4
timestamp 1707688321
transform -1 0 1037 0 1 3238
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_5
timestamp 1707688321
transform -1 0 677 0 1 3396
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_6
timestamp 1707688321
transform -1 0 5141 0 -1 2894
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_7
timestamp 1707688321
transform 1 0 2869 0 -1 3430
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_8
timestamp 1707688321
transform 1 0 6362 0 -1 3576
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_9
timestamp 1707688321
transform 1 0 115 0 1 2786
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_10
timestamp 1707688321
transform 1 0 2231 0 1 3238
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_11
timestamp 1707688321
transform 1 0 7631 0 1 3470
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_12
timestamp 1707688321
transform 1 0 8485 0 1 2786
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_13
timestamp 1707688321
transform 1 0 7847 0 1 3396
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_14
timestamp 1707688321
transform 1 0 2653 0 1 3324
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_15
timestamp 1707688321
transform 1 0 -17 0 1 2712
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_16
timestamp 1707688321
transform 1 0 291 0 1 2786
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1707688321
transform 0 -1 9987 -1 0 3350
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1707688321
transform 0 -1 10555 -1 0 3350
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1707688321
transform -1 0 817 0 1 2860
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1707688321
transform -1 0 7225 0 1 2812
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1707688321
transform -1 0 6605 0 1 2812
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1707688321
transform -1 0 1446 0 1 2398
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1707688321
transform -1 0 1627 0 1 3544
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1707688321
transform -1 0 433 0 1 2404
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1707688321
transform -1 0 4649 0 1 3624
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_9
timestamp 1707688321
transform -1 0 3219 0 1 3238
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_10
timestamp 1707688321
transform -1 0 493 0 1 2264
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_11
timestamp 1707688321
transform -1 0 1913 0 -1 2894
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_12
timestamp 1707688321
transform -1 0 5091 0 -1 3578
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_13
timestamp 1707688321
transform 0 1 1212 1 0 3244
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_14
timestamp 1707688321
transform 0 -1 8786 1 0 3244
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_15
timestamp 1707688321
transform 0 -1 8966 1 0 3244
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_16
timestamp 1707688321
transform 1 0 3343 0 -1 2412
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_17
timestamp 1707688321
transform 1 0 3976 0 -1 2412
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_18
timestamp 1707688321
transform 1 0 -17 0 -1 2968
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_19
timestamp 1707688321
transform 1 0 5157 0 -1 2412
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_20
timestamp 1707688321
transform 1 0 2033 0 1 2812
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_21
timestamp 1707688321
transform 1 0 5524 0 1 2373
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_22
timestamp 1707688321
transform 1 0 10815 0 1 3470
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_23
timestamp 1707688321
transform 1 0 5893 0 1 2860
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_24
timestamp 1707688321
transform 1 0 6015 0 1 2373
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_25
timestamp 1707688321
transform 1 0 2367 0 1 3624
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_26
timestamp 1707688321
transform 1 0 2632 0 1 3698
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_27
timestamp 1707688321
transform 1 0 9570 0 1 3698
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_28
timestamp 1707688321
transform 1 0 4207 0 1 3238
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1707688321
transform 0 -1 17 1 0 645
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1707688321
transform 1 0 6673 0 -1 2894
box 0 0 1 1
use L1M1_CDNS_52468879185308  L1M1_CDNS_52468879185308_0
timestamp 1707688321
transform 0 -1 17 -1 0 1972
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_0
timestamp 1707688321
transform 0 -1 17 -1 0 1325
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_1
timestamp 1707688321
transform 1 0 4015 0 1 3320
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_2
timestamp 1707688321
transform 1 0 9107 0 1 3396
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_3
timestamp 1707688321
transform 1 0 9294 0 1 3622
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1707688321
transform -1 0 658 0 -1 2304
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1707688321
transform 1 0 4755 0 1 3232
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1707688321
transform 1 0 4831 0 1 2366
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_0
timestamp 1707688321
transform 0 -1 658 -1 0 1061
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_0
timestamp 1707688321
transform 0 -1 658 -1 0 1645
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_1
timestamp 1707688321
transform -1 0 1572 0 1 1864
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_2
timestamp 1707688321
transform -1 0 1572 0 1 2706
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_0
timestamp 1707688321
transform -1 0 658 0 1 2476
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_0
timestamp 1707688321
transform 0 -1 26 1 0 638
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_0
timestamp 1707688321
transform -1 0 8350 0 -1 3654
box 0 0 1 1
use M1M2_CDNS_524688791851023  M1M2_CDNS_524688791851023_0
timestamp 1707688321
transform 0 -1 26 -1 0 1978
box 0 0 832 52
use M1M2_CDNS_524688791851081  M1M2_CDNS_524688791851081_0
timestamp 1707688321
transform 1 0 1600 0 1 2034
box 0 0 256 180
use M1M2_CDNS_524688791851150  M1M2_CDNS_524688791851150_0
timestamp 1707688321
transform 1 0 1600 0 -1 3190
box 0 0 256 244
use sky130_fd_io__sio_com_ctl_ls  sky130_fd_io__sio_com_ctl_ls_0
timestamp 1707688321
transform -1 0 2102 0 -1 2304
box -91 0 2150 2319
use sky130_fd_io__sio_hvsbt_diff_space  sky130_fd_io__sio_hvsbt_diff_space_0
timestamp 1707688321
transform -1 0 9522 0 1 2335
box 0 0 1 1
use sky130_fd_io__sio_hvsbt_diff_space  sky130_fd_io__sio_hvsbt_diff_space_1
timestamp 1707688321
transform -1 0 8680 0 1 2335
box 0 0 1 1
use sky130_fd_io__sio_hvsbt_diff_space  sky130_fd_io__sio_hvsbt_diff_space_2
timestamp 1707688321
transform 1 0 1678 0 1 2335
box 0 0 1 1
use sky130_fd_io__sio_hvsbt_diff_space  sky130_fd_io__sio_hvsbt_diff_space_3
timestamp 1707688321
transform 1 0 2492 0 1 2335
box 0 0 1 1
use sky130_fd_io__sio_hvsbt_diff_space  sky130_fd_io__sio_hvsbt_diff_space_4
timestamp 1707688321
transform 1 0 4824 0 1 2335
box 0 0 1 1
use sky130_fd_io__sio_hvsbt_diff_space  sky130_fd_io__sio_hvsbt_diff_space_5
timestamp 1707688321
transform 1 0 6018 0 1 2335
box 0 0 1 1
use sky130_fd_io__sio_hvsbt_diff_space  sky130_fd_io__sio_hvsbt_diff_space_6
timestamp 1707688321
transform 1 0 6656 0 1 2335
box 0 0 1 1
use sky130_fd_io__sio_hvsbt_diff_space  sky130_fd_io__sio_hvsbt_diff_space_7
timestamp 1707688321
transform 1 0 836 0 1 2335
box 0 0 1 1
use sky130_fd_io__sio_hvsbt_diff_space  sky130_fd_io__sio_hvsbt_diff_space_8
timestamp 1707688321
transform 1 0 3658 0 1 2335
box 0 0 1 1
use sky130_fd_io__sio_hvsbt_endcap  sky130_fd_io__sio_hvsbt_endcap_0
timestamp 1707688321
transform -1 0 11103 0 1 2335
box -84 93 164 1337
use sky130_fd_io__sio_hvsbt_inv_x1  sky130_fd_io__sio_hvsbt_inv_x1_0
timestamp 1707688321
transform 1 0 8394 0 1 2335
box -107 21 267 1369
use sky130_fd_io__sio_hvsbt_inv_x1  sky130_fd_io__sio_hvsbt_inv_x1_1
timestamp 1707688321
transform 1 0 6480 0 1 2335
box -107 21 267 1369
use sky130_fd_io__sio_hvsbt_inv_x2  sky130_fd_io__sio_hvsbt_inv_x2_0
timestamp 1707688321
transform 1 0 5314 0 1 2335
box -107 21 459 1369
use sky130_fd_io__sio_hvsbt_inv_x2  sky130_fd_io__sio_hvsbt_inv_x2_1
timestamp 1707688321
transform 1 0 7118 0 1 2335
box -107 21 459 1369
use sky130_fd_io__sio_hvsbt_inv_x2  sky130_fd_io__sio_hvsbt_inv_x2_2
timestamp 1707688321
transform 1 0 10254 0 1 2335
box -107 21 459 1369
use sky130_fd_io__sio_hvsbt_inv_x2  sky130_fd_io__sio_hvsbt_inv_x2_3
timestamp 1707688321
transform 1 0 9902 0 1 2335
box -107 21 459 1369
use sky130_fd_io__sio_hvsbt_nand2  sky130_fd_io__sio_hvsbt_nand2_0
timestamp 1707688321
transform -1 0 9032 0 1 2335
box -107 21 459 1369
use sky130_fd_io__sio_hvsbt_nand2  sky130_fd_io__sio_hvsbt_nand2_1
timestamp 1707688321
transform -1 0 1298 0 1 2335
box -107 21 459 1369
use sky130_fd_io__sio_hvsbt_nand2  sky130_fd_io__sio_hvsbt_nand2_2
timestamp 1707688321
transform -1 0 6480 0 1 2335
box -107 21 459 1369
use sky130_fd_io__sio_hvsbt_nand2  sky130_fd_io__sio_hvsbt_nand2_3
timestamp 1707688321
transform -1 0 2140 0 1 2335
box -107 21 459 1369
use sky130_fd_io__sio_hvsbt_nand2  sky130_fd_io__sio_hvsbt_nand2_4
timestamp 1707688321
transform -1 0 7118 0 1 2335
box -107 21 459 1369
use sky130_fd_io__sio_hvsbt_nand2  sky130_fd_io__sio_hvsbt_nand2_5
timestamp 1707688321
transform -1 0 7932 0 1 2335
box -107 21 459 1369
use sky130_fd_io__sio_hvsbt_nand2  sky130_fd_io__sio_hvsbt_nand2_6
timestamp 1707688321
transform -1 0 484 0 1 2335
box -107 21 459 1369
use sky130_fd_io__sio_hvsbt_nand2  sky130_fd_io__sio_hvsbt_nand2_7
timestamp 1707688321
transform 1 0 5666 0 1 2335
box -107 21 459 1369
use sky130_fd_io__sio_hvsbt_nand2  sky130_fd_io__sio_hvsbt_nand2_8
timestamp 1707688321
transform 1 0 2140 0 1 2335
box -107 21 459 1369
use sky130_fd_io__sio_hvsbt_nand2  sky130_fd_io__sio_hvsbt_nand2_9
timestamp 1707688321
transform 1 0 484 0 1 2335
box -107 21 459 1369
use sky130_fd_io__sio_hvsbt_nor  sky130_fd_io__sio_hvsbt_nor_0
timestamp 1707688321
transform -1 0 9902 0 1 2335
box -107 21 487 1369
use sky130_fd_io__sio_hvsbt_nor  sky130_fd_io__sio_hvsbt_nor_1
timestamp 1707688321
transform 1 0 9032 0 1 2335
box -107 21 487 1369
use sky130_fd_io__sio_hvsbt_nor  sky130_fd_io__sio_hvsbt_nor_2
timestamp 1707688321
transform 1 0 1298 0 1 2335
box -107 21 487 1369
use sky130_fd_io__sio_hvsbt_nor  sky130_fd_io__sio_hvsbt_nor_3
timestamp 1707688321
transform 1 0 10606 0 1 2335
box -107 21 487 1369
use sky130_fd_io__sio_hvsbt_nor_a  sky130_fd_io__sio_hvsbt_nor_a_0
timestamp 1707688321
transform -1 0 5314 0 1 2335
box -107 21 487 1369
use sky130_fd_io__sio_hvsbt_xor  sky130_fd_io__sio_hvsbt_xor_0
timestamp 1707688321
transform -1 0 3658 0 1 2335
box -91 21 1147 1369
use sky130_fd_io__sio_hvsbt_xor  sky130_fd_io__sio_hvsbt_xor_1
timestamp 1707688321
transform 1 0 3768 0 1 2335
box -91 21 1147 1369
<< labels >>
flabel comment s 60 2942 60 2942 0 FreeSans 200 180 0 0 vpb
flabel comment s 60 3038 60 3038 0 FreeSans 200 180 0 0 vpwr
flabel comment s 60 2564 60 2564 0 FreeSans 200 180 0 0 vgnd
flabel comment s 60 2735 60 2735 0 FreeSans 200 180 0 0 vnb
flabel comment s 9700 3338 9700 3338 0 FreeSans 400 0 0 0 pden_h1
flabel comment s 6705 3642 6705 3642 0 FreeSans 200 180 0 0 dm_h<0>
flabel comment s 888 2407 888 2407 0 FreeSans 200 0 0 0 dm_h_n<2>
flabel comment s 6099 3491 6099 3491 0 FreeSans 200 180 0 0 puen_2or1_h
flabel comment s 864 3567 864 3567 0 FreeSans 200 0 0 0 dm_h_n<1>
flabel comment s 892 3268 892 3268 0 FreeSans 200 180 0 0 dm_h_n<0>
flabel comment s 449 2877 449 2877 0 FreeSans 200 180 0 0 n<4>
flabel comment s 5315 2878 5315 2878 0 FreeSans 200 180 0 0 puen_0_h
flabel comment s 5830 2387 5830 2387 0 FreeSans 200 0 0 0 puen_h0_n
flabel comment s 7085 2829 7085 2829 0 FreeSans 200 180 0 0 puen_h1_n
flabel comment s 6774 2890 6774 2890 0 FreeSans 200 180 0 0 n<2>
flabel comment s 6433 2826 6433 2826 0 FreeSans 200 0 0 0 n<5>
flabel comment s 1862 3726 1862 3726 0 FreeSans 200 180 0 0 n<0>
flabel comment s 2133 2847 2133 2847 0 FreeSans 200 180 0 0 n<1>
flabel comment s 1306 3323 1306 3323 0 FreeSans 200 180 0 0 n<9>
flabel comment s 10780 3602 10780 3602 0 FreeSans 200 270 0 0 pden_h0
flabel comment s 10436 3602 10436 3602 0 FreeSans 200 270 0 0 pden_h_n<0>
flabel comment s 10087 3602 10087 3602 0 FreeSans 200 270 0 0 pden_h_n<1>
flabel comment s 9691 3616 9691 3616 0 FreeSans 200 270 0 0 pden_h1
flabel comment s 299 3620 299 3620 0 FreeSans 200 270 0 0 n<4>
flabel comment s 5499 3551 5499 3551 0 FreeSans 200 270 0 0 puen_h<0>
flabel comment s 7238 3551 7238 3551 0 FreeSans 200 270 0 0 puen_h<1>
flabel comment s 6952 3551 6952 3551 0 FreeSans 200 270 0 0 puen_h1_n
flabel comment s 6287 3651 6287 3651 0 FreeSans 200 270 0 0 n<5>
flabel comment s 6640 3655 6640 3655 0 FreeSans 200 270 0 0 n<2>
flabel comment s 5844 3622 5844 3622 0 FreeSans 200 270 0 0 puen_h0_n
flabel comment s 5107 3622 5107 3622 0 FreeSans 200 270 0 0 puen_0_h
flabel comment s 4280 3676 4280 3676 0 FreeSans 200 270 0 0 n<8>
flabel comment s 3112 3653 3112 3653 0 FreeSans 200 270 0 0 n<10>
flabel comment s 2295 3648 2295 3648 0 FreeSans 200 270 0 0 n<1>
flabel comment s 1948 3648 1948 3648 0 FreeSans 200 270 0 0 puen_20r1_h
flabel comment s 1111 3648 1111 3648 0 FreeSans 200 270 0 0 n<0>
flabel comment s 1475 3531 1475 3531 0 FreeSans 200 270 0 0 n<9>
flabel comment s 7841 3731 7841 3731 0 FreeSans 200 180 0 0 dm_h<1>
flabel comment s 7630 3731 7630 3731 0 FreeSans 200 180 0 0 dm_h<0>
flabel comment s 10879 3732 10879 3732 0 FreeSans 200 180 0 0 n<3>
flabel comment s 10676 3732 10676 3732 0 FreeSans 200 180 0 0 pd_dis_h
flabel comment s 10386 3732 10386 3732 0 FreeSans 200 180 0 0 pden_h0
flabel comment s 10058 3732 10058 3732 0 FreeSans 200 180 0 0 pden_h1
flabel comment s 9783 3732 9783 3732 0 FreeSans 200 180 0 0 pd_dis_h
flabel comment s 738 3732 738 3732 0 FreeSans 200 180 0 0 n<4>
flabel comment s 594 3732 594 3732 0 FreeSans 200 180 0 0 dm_h_n<0>
flabel comment s 8500 3735 8500 3735 0 FreeSans 200 0 0 0 frc_lohi_comb
flabel comment s 8720 3735 8720 3735 0 FreeSans 200 0 0 0 force_lo_h_n
flabel comment s 161 3732 161 3732 0 FreeSans 200 0 0 0 dm_h_n<1>
flabel comment s 401 3732 401 3732 0 FreeSans 200 0 0 0 dm_h_n<2>
flabel comment s 5524 3732 5524 3732 0 FreeSans 200 180 0 0 puen_h0_n
flabel comment s 7261 3732 7261 3732 0 FreeSans 200 180 0 0 puen_h1_n
flabel comment s 6831 3732 6831 3732 0 FreeSans 200 180 0 0 n<2>
flabel comment s 6553 3732 6553 3732 0 FreeSans 200 180 0 0 n<5>
flabel comment s 6401 3732 6401 3732 0 FreeSans 200 180 0 0 puen_2or1_h
flabel comment s 6181 3732 6181 3732 0 FreeSans 200 180 0 0 vreg_en_h_n
flabel comment s 5921 3732 5921 3732 0 FreeSans 200 180 0 0 puen_0_h
flabel comment s 5736 3732 5736 3732 0 FreeSans 200 180 0 0 pu_dis_h_n
flabel comment s 5203 3732 5203 3732 0 FreeSans 200 180 0 0 n<8>
flabel comment s 5007 3732 5007 3732 0 FreeSans 200 180 0 0 dm_h_n<1>
flabel comment s 4550 3732 4550 3732 0 FreeSans 200 180 0 0 dm_h<0>
flabel comment s 3977 3732 3977 3732 0 FreeSans 200 180 0 0 dm_h<2>
flabel comment s 3384 3732 3384 3732 0 FreeSans 200 180 0 0 dm_h<2>
flabel comment s 2833 3717 2833 3717 0 FreeSans 200 180 0 0 dm_h<1>
flabel comment s 2374 3732 2374 3732 0 FreeSans 200 180 0 0 dm_h<0>
flabel comment s 2229 3732 2229 3732 0 FreeSans 200 180 0 0 n<10>
flabel comment s 2038 3732 2038 3732 0 FreeSans 200 180 0 0 n<1>
flabel comment s 944 2855 944 2855 0 FreeSans 200 0 0 0 n<0>
flabel comment s 1196 3732 1196 3732 0 FreeSans 200 0 0 0 n<9>
flabel comment s 1384 3732 1384 3732 0 FreeSans 200 0 0 0 dm_h_n<2>
flabel comment s 1581 3732 1581 3732 0 FreeSans 200 0 0 0 dm_h_n<1>
flabel comment s 1015 3732 1015 3732 0 FreeSans 200 0 0 0 dm_h_n<0>
flabel metal1 s 10635 3491 10635 3491 3 FreeSans 400 0 0 0 n<3>
flabel metal1 s 7154 2838 7154 2838 0 FreeSans 400 0 0 0 puen_h1_n
flabel metal1 s 5841 2803 5841 2803 0 FreeSans 400 0 0 0 puen_h0_n
flabel metal1 s 10793 3335 10793 3335 0 FreeSans 400 0 0 0 pden_h0
flabel metal1 s 2560 3259 2560 3259 3 FreeSans 400 0 0 0 n<10>
flabel metal1 s 1483 3334 1483 3334 0 FreeSans 400 0 0 0 n<9>
flabel metal1 s 4664 3262 4664 3262 0 FreeSans 400 0 0 0 n<8>
flabel metal1 s 6491 2834 6491 2834 0 FreeSans 400 0 0 0 n<5>
flabel metal1 s 731 2876 731 2876 0 FreeSans 400 0 0 0 n<4>
flabel metal1 s 6826 2876 6826 2876 0 FreeSans 400 0 0 0 n<2>
flabel metal1 s 2048 2830 2048 2830 0 FreeSans 400 0 0 0 n<1>
flabel metal1 s 1119 2803 1119 2803 0 FreeSans 400 0 0 0 n<0>
flabel metal1 s 132 2706 144 2752 3 FreeSans 400 0 0 0 vgnd
port 2 nsew
flabel metal1 s 3669 2378 3703 2412 3 FreeSans 400 0 0 0 dm_h<2>
port 3 nsew
flabel metal1 s 2074 218 2097 420 3 FreeSans 400 180 0 0 vpwr
port 4 nsew
flabel metal1 s 2102 72 2125 190 3 FreeSans 400 180 0 0 vpb
port 5 nsew
flabel metal1 s 2102 1854 2125 1984 3 FreeSans 400 180 0 0 vgnd
port 2 nsew
flabel metal1 s 132 2476 144 2678 3 FreeSans 400 0 0 0 vgnd
port 2 nsew
flabel metal1 s 132 3002 144 3204 3 FreeSans 400 0 0 0 vcc_io
port 6 nsew
flabel metal1 s 1747 1607 1781 1641 0 FreeSans 400 0 0 0 slow_h_n
port 7 nsew
flabel metal1 s 99 1221 133 1255 0 FreeSans 400 0 0 0 slow
port 8 nsew
flabel metal1 s 6362 3470 6395 3505 0 FreeSans 400 0 0 0 puen_2or1_h
port 9 nsew
flabel metal1 s 5893 2860 5927 2894 0 FreeSans 400 0 0 0 puen_0_h
port 10 nsew
flabel metal1 s 2102 863 2125 1065 3 FreeSans 400 180 0 0 vgnd
port 2 nsew
flabel metal1 s 2085 2012 2125 2214 3 FreeSans 400 180 0 0 vcc_io
port 6 nsew
flabel metal1 s 1873 795 1907 829 0 FreeSans 400 0 0 0 hld_i_vpwr
port 11 nsew
flabel metal1 s 363 2404 397 2438 0 FreeSans 400 0 0 0 dm_h_n<2>
port 12 nsew
flabel metal1 s 223 3501 257 3536 3 FreeSans 400 0 0 0 dm_h_n<1>
port 13 nsew
flabel metal1 s 563 3310 597 3344 0 FreeSans 400 0 0 0 dm_h_n<0>
port 14 nsew
flabel metal1 s 2869 3396 2903 3430 3 FreeSans 400 0 0 0 dm_h<1>
port 15 nsew
flabel metal1 s 2401 3618 2436 3652 0 FreeSans 400 0 0 0 dm_h<0>
port 16 nsew
flabel locali s 735 2254 769 2288 0 FreeSans 200 0 0 0 hld_i_h_n
port 17 nsew
flabel locali s 6201 3654 6235 3704 3 FreeSans 400 0 0 0 vreg_en_h_n
port 18 nsew
flabel locali s 7277 3555 7311 3604 0 FreeSans 400 0 0 0 puen_h<1>
port 19 nsew
flabel locali s 5473 3555 5507 3604 0 FreeSans 400 0 0 0 puen_h<0>
port 20 nsew
flabel locali s 10061 3555 10095 3604 0 FreeSans 400 0 0 0 pden_h_n<1>
port 21 nsew
flabel locali s 10413 3555 10447 3604 0 FreeSans 400 0 0 0 pden_h_n<0>
port 22 nsew
flabel locali s 233 2254 267 2288 3 FreeSans 400 0 0 0 od_h
port 23 nsew
flabel locali s 8839 3556 8873 3605 0 FreeSans 400 0 0 0 pden_h_n<2>
port 24 nsew
flabel metal2 s 1461 1220 1491 1250 0 FreeSans 400 0 0 0 slow_h
port 25 nsew
<< properties >>
string GDS_END 87702204
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87675040
string path 0.000 0.050 0.000 13.675 
<< end >>
