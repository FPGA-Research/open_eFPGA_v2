magic
tech sky130A
timestamp 1707688321
<< locali >>
rect 17 0 36 17
rect 53 0 72 17
rect 89 0 108 17
rect 125 0 144 17
rect 161 0 180 17
rect 197 0 216 17
rect 233 0 252 17
rect 269 0 288 17
rect 305 0 324 17
rect 341 0 360 17
rect 377 0 396 17
rect 413 0 432 17
rect 449 0 468 17
rect 485 0 504 17
rect 521 0 540 17
rect 557 0 576 17
rect 593 0 612 17
rect 629 0 648 17
rect 665 0 684 17
rect 701 0 720 17
rect 737 0 756 17
rect 773 0 792 17
rect 809 0 828 17
rect 845 0 864 17
rect 881 0 900 17
rect 917 0 936 17
rect 953 0 972 17
rect 989 0 1008 17
rect 1025 0 1044 17
rect 1061 0 1080 17
rect 1097 0 1116 17
rect 1133 0 1152 17
rect 1169 0 1188 17
rect 1205 0 1224 17
rect 1241 0 1260 17
rect 1277 0 1296 17
rect 1313 0 1332 17
rect 1349 0 1368 17
rect 1385 0 1404 17
rect 1421 0 1440 17
rect 1457 0 1476 17
rect 1493 0 1512 17
rect 1529 0 1548 17
rect 1565 0 1584 17
rect 1601 0 1620 17
rect 1637 0 1656 17
rect 1673 0 1692 17
rect 1709 0 1728 17
rect 1745 0 1764 17
rect 1781 0 1800 17
rect 1817 0 1836 17
rect 1853 0 1872 17
rect 1889 0 1908 17
rect 1925 0 1944 17
rect 1961 0 1980 17
rect 1997 0 2016 17
rect 2033 0 2052 17
rect 2069 0 2088 17
rect 2105 0 2124 17
rect 2141 0 2160 17
rect 2177 0 2196 17
rect 2213 0 2232 17
rect 2249 0 2268 17
rect 2285 0 2304 17
rect 2321 0 2340 17
rect 2357 0 2376 17
rect 2393 0 2412 17
rect 2429 0 2448 17
rect 2465 0 2484 17
rect 2501 0 2520 17
rect 2537 0 2556 17
rect 2573 0 2592 17
rect 2609 0 2628 17
rect 2645 0 2664 17
rect 2681 0 2700 17
rect 2717 0 2736 17
rect 2753 0 2772 17
rect 2789 0 2808 17
rect 2825 0 2844 17
rect 2861 0 2880 17
rect 2897 0 2916 17
rect 2933 0 2952 17
rect 2969 0 2988 17
rect 3005 0 3024 17
rect 3041 0 3060 17
rect 3077 0 3096 17
rect 3113 0 3132 17
rect 3149 0 3168 17
rect 3185 0 3204 17
rect 3221 0 3240 17
rect 3257 0 3276 17
rect 3293 0 3312 17
rect 3329 0 3348 17
rect 3365 0 3384 17
rect 3401 0 3420 17
rect 3437 0 3456 17
rect 3473 0 3492 17
rect 3509 0 3528 17
rect 3545 0 3564 17
rect 3581 0 3600 17
rect 3617 0 3636 17
rect 3653 0 3672 17
rect 3689 0 3708 17
rect 3725 0 3744 17
rect 3761 0 3780 17
rect 3797 0 3816 17
rect 3833 0 3852 17
rect 3869 0 3888 17
rect 3905 0 3924 17
rect 3941 0 3960 17
rect 3977 0 3996 17
rect 4013 0 4032 17
rect 4049 0 4068 17
rect 4085 0 4104 17
rect 4121 0 4140 17
rect 4157 0 4176 17
rect 4193 0 4212 17
rect 4229 0 4248 17
rect 4265 0 4284 17
rect 4301 0 4320 17
rect 4337 0 4356 17
rect 4373 0 4392 17
rect 4409 0 4428 17
rect 4445 0 4464 17
rect 4481 0 4500 17
rect 4517 0 4536 17
rect 4553 0 4572 17
rect 4589 0 4608 17
rect 4625 0 4644 17
rect 4661 0 4680 17
rect 4697 0 4716 17
rect 4733 0 4752 17
rect 4769 0 4788 17
rect 4805 0 4824 17
rect 4841 0 4860 17
rect 4877 0 4896 17
rect 4913 0 4932 17
rect 4949 0 4968 17
rect 4985 0 5004 17
rect 5021 0 5040 17
rect 5057 0 5076 17
rect 5093 0 5112 17
rect 5129 0 5148 17
rect 5165 0 5184 17
rect 5201 0 5220 17
rect 5237 0 5256 17
rect 5273 0 5292 17
rect 5309 0 5328 17
rect 5345 0 5364 17
rect 5381 0 5400 17
rect 5417 0 5436 17
rect 5453 0 5472 17
rect 5489 0 5508 17
rect 5525 0 5544 17
rect 5561 0 5580 17
rect 5597 0 5616 17
rect 5633 0 5652 17
rect 5669 0 5688 17
rect 5705 0 5724 17
rect 5741 0 5760 17
rect 5777 0 5796 17
rect 5813 0 5832 17
rect 5849 0 5868 17
rect 5885 0 5904 17
rect 5921 0 5940 17
rect 5957 0 5976 17
rect 5993 0 6012 17
rect 6029 0 6048 17
rect 6065 0 6084 17
rect 6101 0 6120 17
rect 6137 0 6156 17
rect 6173 0 6192 17
rect 6209 0 6228 17
rect 6245 0 6264 17
rect 6281 0 6300 17
rect 6317 0 6336 17
rect 6353 0 6372 17
rect 6389 0 6408 17
rect 6425 0 6444 17
rect 6461 0 6480 17
rect 6497 0 6516 17
rect 6533 0 6552 17
rect 6569 0 6588 17
rect 6605 0 6624 17
rect 6641 0 6660 17
rect 6677 0 6696 17
rect 6713 0 6732 17
rect 6749 0 6768 17
rect 6785 0 6804 17
rect 6821 0 6840 17
rect 6857 0 6876 17
rect 6893 0 6912 17
rect 6929 0 6948 17
rect 6965 0 6984 17
rect 7001 0 7020 17
rect 7037 0 7056 17
rect 7073 0 7092 17
rect 7109 0 7128 17
rect 7145 0 7164 17
rect 7181 0 7200 17
rect 7217 0 7236 17
rect 7253 0 7272 17
rect 7289 0 7308 17
rect 7325 0 7344 17
rect 7361 0 7380 17
rect 7397 0 7416 17
rect 7433 0 7452 17
rect 7469 0 7488 17
rect 7505 0 7524 17
rect 7541 0 7560 17
rect 7577 0 7596 17
rect 7613 0 7632 17
rect 7649 0 7668 17
rect 7685 0 7704 17
rect 7721 0 7740 17
rect 7757 0 7776 17
rect 7793 0 7812 17
rect 7829 0 7848 17
rect 7865 0 7884 17
rect 7901 0 7920 17
rect 7937 0 7956 17
rect 7973 0 7992 17
rect 8009 0 8028 17
rect 8045 0 8064 17
rect 8081 0 8100 17
rect 8117 0 8136 17
rect 8153 0 8172 17
rect 8189 0 8208 17
rect 8225 0 8244 17
rect 8261 0 8280 17
rect 8297 0 8316 17
rect 8333 0 8352 17
rect 8369 0 8388 17
rect 8405 0 8424 17
rect 8441 0 8460 17
rect 8477 0 8496 17
rect 8513 0 8532 17
rect 8549 0 8568 17
rect 8585 0 8604 17
rect 8621 0 8640 17
rect 8657 0 8676 17
rect 8693 0 8712 17
rect 8729 0 8748 17
rect 8765 0 8784 17
rect 8801 0 8820 17
rect 8837 0 8856 17
rect 8873 0 8892 17
rect 8909 0 8928 17
rect 8945 0 8964 17
rect 8981 0 9000 17
rect 9017 0 9036 17
rect 9053 0 9072 17
rect 9089 0 9108 17
rect 9125 0 9144 17
rect 9161 0 9180 17
rect 9197 0 9216 17
rect 9233 0 9252 17
rect 9269 0 9288 17
rect 9305 0 9324 17
rect 9341 0 9360 17
rect 9377 0 9396 17
rect 9413 0 9432 17
rect 9449 0 9468 17
rect 9485 0 9504 17
rect 9521 0 9540 17
rect 9557 0 9576 17
rect 9593 0 9612 17
rect 9629 0 9648 17
rect 9665 0 9684 17
rect 9701 0 9720 17
rect 9737 0 9756 17
rect 9773 0 9792 17
rect 9809 0 9828 17
rect 9845 0 9864 17
rect 9881 0 9900 17
rect 9917 0 9936 17
rect 9953 0 9972 17
rect 9989 0 10008 17
rect 10025 0 10044 17
rect 10061 0 10080 17
rect 10097 0 10116 17
rect 10133 0 10152 17
rect 10169 0 10188 17
rect 10205 0 10224 17
rect 10241 0 10260 17
rect 10277 0 10296 17
rect 10313 0 10332 17
<< viali >>
rect 0 0 17 17
rect 36 0 53 17
rect 72 0 89 17
rect 108 0 125 17
rect 144 0 161 17
rect 180 0 197 17
rect 216 0 233 17
rect 252 0 269 17
rect 288 0 305 17
rect 324 0 341 17
rect 360 0 377 17
rect 396 0 413 17
rect 432 0 449 17
rect 468 0 485 17
rect 504 0 521 17
rect 540 0 557 17
rect 576 0 593 17
rect 612 0 629 17
rect 648 0 665 17
rect 684 0 701 17
rect 720 0 737 17
rect 756 0 773 17
rect 792 0 809 17
rect 828 0 845 17
rect 864 0 881 17
rect 900 0 917 17
rect 936 0 953 17
rect 972 0 989 17
rect 1008 0 1025 17
rect 1044 0 1061 17
rect 1080 0 1097 17
rect 1116 0 1133 17
rect 1152 0 1169 17
rect 1188 0 1205 17
rect 1224 0 1241 17
rect 1260 0 1277 17
rect 1296 0 1313 17
rect 1332 0 1349 17
rect 1368 0 1385 17
rect 1404 0 1421 17
rect 1440 0 1457 17
rect 1476 0 1493 17
rect 1512 0 1529 17
rect 1548 0 1565 17
rect 1584 0 1601 17
rect 1620 0 1637 17
rect 1656 0 1673 17
rect 1692 0 1709 17
rect 1728 0 1745 17
rect 1764 0 1781 17
rect 1800 0 1817 17
rect 1836 0 1853 17
rect 1872 0 1889 17
rect 1908 0 1925 17
rect 1944 0 1961 17
rect 1980 0 1997 17
rect 2016 0 2033 17
rect 2052 0 2069 17
rect 2088 0 2105 17
rect 2124 0 2141 17
rect 2160 0 2177 17
rect 2196 0 2213 17
rect 2232 0 2249 17
rect 2268 0 2285 17
rect 2304 0 2321 17
rect 2340 0 2357 17
rect 2376 0 2393 17
rect 2412 0 2429 17
rect 2448 0 2465 17
rect 2484 0 2501 17
rect 2520 0 2537 17
rect 2556 0 2573 17
rect 2592 0 2609 17
rect 2628 0 2645 17
rect 2664 0 2681 17
rect 2700 0 2717 17
rect 2736 0 2753 17
rect 2772 0 2789 17
rect 2808 0 2825 17
rect 2844 0 2861 17
rect 2880 0 2897 17
rect 2916 0 2933 17
rect 2952 0 2969 17
rect 2988 0 3005 17
rect 3024 0 3041 17
rect 3060 0 3077 17
rect 3096 0 3113 17
rect 3132 0 3149 17
rect 3168 0 3185 17
rect 3204 0 3221 17
rect 3240 0 3257 17
rect 3276 0 3293 17
rect 3312 0 3329 17
rect 3348 0 3365 17
rect 3384 0 3401 17
rect 3420 0 3437 17
rect 3456 0 3473 17
rect 3492 0 3509 17
rect 3528 0 3545 17
rect 3564 0 3581 17
rect 3600 0 3617 17
rect 3636 0 3653 17
rect 3672 0 3689 17
rect 3708 0 3725 17
rect 3744 0 3761 17
rect 3780 0 3797 17
rect 3816 0 3833 17
rect 3852 0 3869 17
rect 3888 0 3905 17
rect 3924 0 3941 17
rect 3960 0 3977 17
rect 3996 0 4013 17
rect 4032 0 4049 17
rect 4068 0 4085 17
rect 4104 0 4121 17
rect 4140 0 4157 17
rect 4176 0 4193 17
rect 4212 0 4229 17
rect 4248 0 4265 17
rect 4284 0 4301 17
rect 4320 0 4337 17
rect 4356 0 4373 17
rect 4392 0 4409 17
rect 4428 0 4445 17
rect 4464 0 4481 17
rect 4500 0 4517 17
rect 4536 0 4553 17
rect 4572 0 4589 17
rect 4608 0 4625 17
rect 4644 0 4661 17
rect 4680 0 4697 17
rect 4716 0 4733 17
rect 4752 0 4769 17
rect 4788 0 4805 17
rect 4824 0 4841 17
rect 4860 0 4877 17
rect 4896 0 4913 17
rect 4932 0 4949 17
rect 4968 0 4985 17
rect 5004 0 5021 17
rect 5040 0 5057 17
rect 5076 0 5093 17
rect 5112 0 5129 17
rect 5148 0 5165 17
rect 5184 0 5201 17
rect 5220 0 5237 17
rect 5256 0 5273 17
rect 5292 0 5309 17
rect 5328 0 5345 17
rect 5364 0 5381 17
rect 5400 0 5417 17
rect 5436 0 5453 17
rect 5472 0 5489 17
rect 5508 0 5525 17
rect 5544 0 5561 17
rect 5580 0 5597 17
rect 5616 0 5633 17
rect 5652 0 5669 17
rect 5688 0 5705 17
rect 5724 0 5741 17
rect 5760 0 5777 17
rect 5796 0 5813 17
rect 5832 0 5849 17
rect 5868 0 5885 17
rect 5904 0 5921 17
rect 5940 0 5957 17
rect 5976 0 5993 17
rect 6012 0 6029 17
rect 6048 0 6065 17
rect 6084 0 6101 17
rect 6120 0 6137 17
rect 6156 0 6173 17
rect 6192 0 6209 17
rect 6228 0 6245 17
rect 6264 0 6281 17
rect 6300 0 6317 17
rect 6336 0 6353 17
rect 6372 0 6389 17
rect 6408 0 6425 17
rect 6444 0 6461 17
rect 6480 0 6497 17
rect 6516 0 6533 17
rect 6552 0 6569 17
rect 6588 0 6605 17
rect 6624 0 6641 17
rect 6660 0 6677 17
rect 6696 0 6713 17
rect 6732 0 6749 17
rect 6768 0 6785 17
rect 6804 0 6821 17
rect 6840 0 6857 17
rect 6876 0 6893 17
rect 6912 0 6929 17
rect 6948 0 6965 17
rect 6984 0 7001 17
rect 7020 0 7037 17
rect 7056 0 7073 17
rect 7092 0 7109 17
rect 7128 0 7145 17
rect 7164 0 7181 17
rect 7200 0 7217 17
rect 7236 0 7253 17
rect 7272 0 7289 17
rect 7308 0 7325 17
rect 7344 0 7361 17
rect 7380 0 7397 17
rect 7416 0 7433 17
rect 7452 0 7469 17
rect 7488 0 7505 17
rect 7524 0 7541 17
rect 7560 0 7577 17
rect 7596 0 7613 17
rect 7632 0 7649 17
rect 7668 0 7685 17
rect 7704 0 7721 17
rect 7740 0 7757 17
rect 7776 0 7793 17
rect 7812 0 7829 17
rect 7848 0 7865 17
rect 7884 0 7901 17
rect 7920 0 7937 17
rect 7956 0 7973 17
rect 7992 0 8009 17
rect 8028 0 8045 17
rect 8064 0 8081 17
rect 8100 0 8117 17
rect 8136 0 8153 17
rect 8172 0 8189 17
rect 8208 0 8225 17
rect 8244 0 8261 17
rect 8280 0 8297 17
rect 8316 0 8333 17
rect 8352 0 8369 17
rect 8388 0 8405 17
rect 8424 0 8441 17
rect 8460 0 8477 17
rect 8496 0 8513 17
rect 8532 0 8549 17
rect 8568 0 8585 17
rect 8604 0 8621 17
rect 8640 0 8657 17
rect 8676 0 8693 17
rect 8712 0 8729 17
rect 8748 0 8765 17
rect 8784 0 8801 17
rect 8820 0 8837 17
rect 8856 0 8873 17
rect 8892 0 8909 17
rect 8928 0 8945 17
rect 8964 0 8981 17
rect 9000 0 9017 17
rect 9036 0 9053 17
rect 9072 0 9089 17
rect 9108 0 9125 17
rect 9144 0 9161 17
rect 9180 0 9197 17
rect 9216 0 9233 17
rect 9252 0 9269 17
rect 9288 0 9305 17
rect 9324 0 9341 17
rect 9360 0 9377 17
rect 9396 0 9413 17
rect 9432 0 9449 17
rect 9468 0 9485 17
rect 9504 0 9521 17
rect 9540 0 9557 17
rect 9576 0 9593 17
rect 9612 0 9629 17
rect 9648 0 9665 17
rect 9684 0 9701 17
rect 9720 0 9737 17
rect 9756 0 9773 17
rect 9792 0 9809 17
rect 9828 0 9845 17
rect 9864 0 9881 17
rect 9900 0 9917 17
rect 9936 0 9953 17
rect 9972 0 9989 17
rect 10008 0 10025 17
rect 10044 0 10061 17
rect 10080 0 10097 17
rect 10116 0 10133 17
rect 10152 0 10169 17
rect 10188 0 10205 17
rect 10224 0 10241 17
rect 10260 0 10277 17
rect 10296 0 10313 17
rect 10332 0 10349 17
<< metal1 >>
rect -6 17 10355 20
rect -6 0 0 17
rect 17 0 36 17
rect 53 0 72 17
rect 89 0 108 17
rect 125 0 144 17
rect 161 0 180 17
rect 197 0 216 17
rect 233 0 252 17
rect 269 0 288 17
rect 305 0 324 17
rect 341 0 360 17
rect 377 0 396 17
rect 413 0 432 17
rect 449 0 468 17
rect 485 0 504 17
rect 521 0 540 17
rect 557 0 576 17
rect 593 0 612 17
rect 629 0 648 17
rect 665 0 684 17
rect 701 0 720 17
rect 737 0 756 17
rect 773 0 792 17
rect 809 0 828 17
rect 845 0 864 17
rect 881 0 900 17
rect 917 0 936 17
rect 953 0 972 17
rect 989 0 1008 17
rect 1025 0 1044 17
rect 1061 0 1080 17
rect 1097 0 1116 17
rect 1133 0 1152 17
rect 1169 0 1188 17
rect 1205 0 1224 17
rect 1241 0 1260 17
rect 1277 0 1296 17
rect 1313 0 1332 17
rect 1349 0 1368 17
rect 1385 0 1404 17
rect 1421 0 1440 17
rect 1457 0 1476 17
rect 1493 0 1512 17
rect 1529 0 1548 17
rect 1565 0 1584 17
rect 1601 0 1620 17
rect 1637 0 1656 17
rect 1673 0 1692 17
rect 1709 0 1728 17
rect 1745 0 1764 17
rect 1781 0 1800 17
rect 1817 0 1836 17
rect 1853 0 1872 17
rect 1889 0 1908 17
rect 1925 0 1944 17
rect 1961 0 1980 17
rect 1997 0 2016 17
rect 2033 0 2052 17
rect 2069 0 2088 17
rect 2105 0 2124 17
rect 2141 0 2160 17
rect 2177 0 2196 17
rect 2213 0 2232 17
rect 2249 0 2268 17
rect 2285 0 2304 17
rect 2321 0 2340 17
rect 2357 0 2376 17
rect 2393 0 2412 17
rect 2429 0 2448 17
rect 2465 0 2484 17
rect 2501 0 2520 17
rect 2537 0 2556 17
rect 2573 0 2592 17
rect 2609 0 2628 17
rect 2645 0 2664 17
rect 2681 0 2700 17
rect 2717 0 2736 17
rect 2753 0 2772 17
rect 2789 0 2808 17
rect 2825 0 2844 17
rect 2861 0 2880 17
rect 2897 0 2916 17
rect 2933 0 2952 17
rect 2969 0 2988 17
rect 3005 0 3024 17
rect 3041 0 3060 17
rect 3077 0 3096 17
rect 3113 0 3132 17
rect 3149 0 3168 17
rect 3185 0 3204 17
rect 3221 0 3240 17
rect 3257 0 3276 17
rect 3293 0 3312 17
rect 3329 0 3348 17
rect 3365 0 3384 17
rect 3401 0 3420 17
rect 3437 0 3456 17
rect 3473 0 3492 17
rect 3509 0 3528 17
rect 3545 0 3564 17
rect 3581 0 3600 17
rect 3617 0 3636 17
rect 3653 0 3672 17
rect 3689 0 3708 17
rect 3725 0 3744 17
rect 3761 0 3780 17
rect 3797 0 3816 17
rect 3833 0 3852 17
rect 3869 0 3888 17
rect 3905 0 3924 17
rect 3941 0 3960 17
rect 3977 0 3996 17
rect 4013 0 4032 17
rect 4049 0 4068 17
rect 4085 0 4104 17
rect 4121 0 4140 17
rect 4157 0 4176 17
rect 4193 0 4212 17
rect 4229 0 4248 17
rect 4265 0 4284 17
rect 4301 0 4320 17
rect 4337 0 4356 17
rect 4373 0 4392 17
rect 4409 0 4428 17
rect 4445 0 4464 17
rect 4481 0 4500 17
rect 4517 0 4536 17
rect 4553 0 4572 17
rect 4589 0 4608 17
rect 4625 0 4644 17
rect 4661 0 4680 17
rect 4697 0 4716 17
rect 4733 0 4752 17
rect 4769 0 4788 17
rect 4805 0 4824 17
rect 4841 0 4860 17
rect 4877 0 4896 17
rect 4913 0 4932 17
rect 4949 0 4968 17
rect 4985 0 5004 17
rect 5021 0 5040 17
rect 5057 0 5076 17
rect 5093 0 5112 17
rect 5129 0 5148 17
rect 5165 0 5184 17
rect 5201 0 5220 17
rect 5237 0 5256 17
rect 5273 0 5292 17
rect 5309 0 5328 17
rect 5345 0 5364 17
rect 5381 0 5400 17
rect 5417 0 5436 17
rect 5453 0 5472 17
rect 5489 0 5508 17
rect 5525 0 5544 17
rect 5561 0 5580 17
rect 5597 0 5616 17
rect 5633 0 5652 17
rect 5669 0 5688 17
rect 5705 0 5724 17
rect 5741 0 5760 17
rect 5777 0 5796 17
rect 5813 0 5832 17
rect 5849 0 5868 17
rect 5885 0 5904 17
rect 5921 0 5940 17
rect 5957 0 5976 17
rect 5993 0 6012 17
rect 6029 0 6048 17
rect 6065 0 6084 17
rect 6101 0 6120 17
rect 6137 0 6156 17
rect 6173 0 6192 17
rect 6209 0 6228 17
rect 6245 0 6264 17
rect 6281 0 6300 17
rect 6317 0 6336 17
rect 6353 0 6372 17
rect 6389 0 6408 17
rect 6425 0 6444 17
rect 6461 0 6480 17
rect 6497 0 6516 17
rect 6533 0 6552 17
rect 6569 0 6588 17
rect 6605 0 6624 17
rect 6641 0 6660 17
rect 6677 0 6696 17
rect 6713 0 6732 17
rect 6749 0 6768 17
rect 6785 0 6804 17
rect 6821 0 6840 17
rect 6857 0 6876 17
rect 6893 0 6912 17
rect 6929 0 6948 17
rect 6965 0 6984 17
rect 7001 0 7020 17
rect 7037 0 7056 17
rect 7073 0 7092 17
rect 7109 0 7128 17
rect 7145 0 7164 17
rect 7181 0 7200 17
rect 7217 0 7236 17
rect 7253 0 7272 17
rect 7289 0 7308 17
rect 7325 0 7344 17
rect 7361 0 7380 17
rect 7397 0 7416 17
rect 7433 0 7452 17
rect 7469 0 7488 17
rect 7505 0 7524 17
rect 7541 0 7560 17
rect 7577 0 7596 17
rect 7613 0 7632 17
rect 7649 0 7668 17
rect 7685 0 7704 17
rect 7721 0 7740 17
rect 7757 0 7776 17
rect 7793 0 7812 17
rect 7829 0 7848 17
rect 7865 0 7884 17
rect 7901 0 7920 17
rect 7937 0 7956 17
rect 7973 0 7992 17
rect 8009 0 8028 17
rect 8045 0 8064 17
rect 8081 0 8100 17
rect 8117 0 8136 17
rect 8153 0 8172 17
rect 8189 0 8208 17
rect 8225 0 8244 17
rect 8261 0 8280 17
rect 8297 0 8316 17
rect 8333 0 8352 17
rect 8369 0 8388 17
rect 8405 0 8424 17
rect 8441 0 8460 17
rect 8477 0 8496 17
rect 8513 0 8532 17
rect 8549 0 8568 17
rect 8585 0 8604 17
rect 8621 0 8640 17
rect 8657 0 8676 17
rect 8693 0 8712 17
rect 8729 0 8748 17
rect 8765 0 8784 17
rect 8801 0 8820 17
rect 8837 0 8856 17
rect 8873 0 8892 17
rect 8909 0 8928 17
rect 8945 0 8964 17
rect 8981 0 9000 17
rect 9017 0 9036 17
rect 9053 0 9072 17
rect 9089 0 9108 17
rect 9125 0 9144 17
rect 9161 0 9180 17
rect 9197 0 9216 17
rect 9233 0 9252 17
rect 9269 0 9288 17
rect 9305 0 9324 17
rect 9341 0 9360 17
rect 9377 0 9396 17
rect 9413 0 9432 17
rect 9449 0 9468 17
rect 9485 0 9504 17
rect 9521 0 9540 17
rect 9557 0 9576 17
rect 9593 0 9612 17
rect 9629 0 9648 17
rect 9665 0 9684 17
rect 9701 0 9720 17
rect 9737 0 9756 17
rect 9773 0 9792 17
rect 9809 0 9828 17
rect 9845 0 9864 17
rect 9881 0 9900 17
rect 9917 0 9936 17
rect 9953 0 9972 17
rect 9989 0 10008 17
rect 10025 0 10044 17
rect 10061 0 10080 17
rect 10097 0 10116 17
rect 10133 0 10152 17
rect 10169 0 10188 17
rect 10205 0 10224 17
rect 10241 0 10260 17
rect 10277 0 10296 17
rect 10313 0 10332 17
rect 10349 0 10355 17
rect -6 -3 10355 0
<< properties >>
string GDS_END 78601546
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 78582982
<< end >>
