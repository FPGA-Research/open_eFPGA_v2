magic
tech sky130B
timestamp 1707688321
<< locali >>
rect 0 3509 17 3528
rect 0 3473 17 3492
rect 0 3437 17 3456
rect 0 3401 17 3420
rect 0 3365 17 3384
rect 0 3329 17 3348
rect 0 3293 17 3312
rect 0 3257 17 3276
rect 0 3221 17 3240
rect 0 3185 17 3204
rect 0 3149 17 3168
rect 0 3113 17 3132
rect 0 3077 17 3096
rect 0 3041 17 3060
rect 0 3005 17 3024
rect 0 2969 17 2988
rect 0 2933 17 2952
rect 0 2897 17 2916
rect 0 2861 17 2880
rect 0 2825 17 2844
rect 0 2789 17 2808
rect 0 2753 17 2772
rect 0 2717 17 2736
rect 0 2681 17 2700
rect 0 2645 17 2664
rect 0 2609 17 2628
rect 0 2573 17 2592
rect 0 2537 17 2556
rect 0 2501 17 2520
rect 0 2465 17 2484
rect 0 2429 17 2448
rect 0 2393 17 2412
rect 0 2357 17 2376
rect 0 2321 17 2340
rect 0 2285 17 2304
rect 0 2249 17 2268
rect 0 2213 17 2232
rect 0 2177 17 2196
rect 0 2141 17 2160
rect 0 2105 17 2124
rect 0 2069 17 2088
rect 0 2033 17 2052
rect 0 1997 17 2016
rect 0 1961 17 1980
rect 0 1925 17 1944
rect 0 1889 17 1908
rect 0 1853 17 1872
rect 0 1817 17 1836
rect 0 1781 17 1800
rect 0 1745 17 1764
rect 0 1709 17 1728
rect 0 1673 17 1692
rect 0 1637 17 1656
rect 0 1601 17 1620
rect 0 1565 17 1584
rect 0 1529 17 1548
rect 0 1493 17 1512
rect 0 1457 17 1476
rect 0 1421 17 1440
rect 0 1385 17 1404
rect 0 1349 17 1368
rect 0 1313 17 1332
rect 0 1277 17 1296
rect 0 1241 17 1260
rect 0 1205 17 1224
rect 0 1169 17 1188
rect 0 1133 17 1152
rect 0 1097 17 1116
rect 0 1061 17 1080
rect 0 1025 17 1044
rect 0 989 17 1008
rect 0 953 17 972
rect 0 917 17 936
rect 0 881 17 900
rect 0 845 17 864
rect 0 809 17 828
rect 0 773 17 792
rect 0 737 17 756
rect 0 701 17 720
rect 0 665 17 684
rect 0 629 17 648
rect 0 593 17 612
rect 0 557 17 576
rect 0 521 17 540
rect 0 485 17 504
rect 0 449 17 468
rect 0 413 17 432
rect 0 377 17 396
rect 0 341 17 360
rect 0 305 17 324
rect 0 269 17 288
rect 0 233 17 252
rect 0 197 17 216
rect 0 161 17 180
rect 0 125 17 144
rect 0 89 17 108
rect 0 53 17 72
rect 0 17 17 36
<< viali >>
rect 0 3528 17 3545
rect 0 3492 17 3509
rect 0 3456 17 3473
rect 0 3420 17 3437
rect 0 3384 17 3401
rect 0 3348 17 3365
rect 0 3312 17 3329
rect 0 3276 17 3293
rect 0 3240 17 3257
rect 0 3204 17 3221
rect 0 3168 17 3185
rect 0 3132 17 3149
rect 0 3096 17 3113
rect 0 3060 17 3077
rect 0 3024 17 3041
rect 0 2988 17 3005
rect 0 2952 17 2969
rect 0 2916 17 2933
rect 0 2880 17 2897
rect 0 2844 17 2861
rect 0 2808 17 2825
rect 0 2772 17 2789
rect 0 2736 17 2753
rect 0 2700 17 2717
rect 0 2664 17 2681
rect 0 2628 17 2645
rect 0 2592 17 2609
rect 0 2556 17 2573
rect 0 2520 17 2537
rect 0 2484 17 2501
rect 0 2448 17 2465
rect 0 2412 17 2429
rect 0 2376 17 2393
rect 0 2340 17 2357
rect 0 2304 17 2321
rect 0 2268 17 2285
rect 0 2232 17 2249
rect 0 2196 17 2213
rect 0 2160 17 2177
rect 0 2124 17 2141
rect 0 2088 17 2105
rect 0 2052 17 2069
rect 0 2016 17 2033
rect 0 1980 17 1997
rect 0 1944 17 1961
rect 0 1908 17 1925
rect 0 1872 17 1889
rect 0 1836 17 1853
rect 0 1800 17 1817
rect 0 1764 17 1781
rect 0 1728 17 1745
rect 0 1692 17 1709
rect 0 1656 17 1673
rect 0 1620 17 1637
rect 0 1584 17 1601
rect 0 1548 17 1565
rect 0 1512 17 1529
rect 0 1476 17 1493
rect 0 1440 17 1457
rect 0 1404 17 1421
rect 0 1368 17 1385
rect 0 1332 17 1349
rect 0 1296 17 1313
rect 0 1260 17 1277
rect 0 1224 17 1241
rect 0 1188 17 1205
rect 0 1152 17 1169
rect 0 1116 17 1133
rect 0 1080 17 1097
rect 0 1044 17 1061
rect 0 1008 17 1025
rect 0 972 17 989
rect 0 936 17 953
rect 0 900 17 917
rect 0 864 17 881
rect 0 828 17 845
rect 0 792 17 809
rect 0 756 17 773
rect 0 720 17 737
rect 0 684 17 701
rect 0 648 17 665
rect 0 612 17 629
rect 0 576 17 593
rect 0 540 17 557
rect 0 504 17 521
rect 0 468 17 485
rect 0 432 17 449
rect 0 396 17 413
rect 0 360 17 377
rect 0 324 17 341
rect 0 288 17 305
rect 0 252 17 269
rect 0 216 17 233
rect 0 180 17 197
rect 0 144 17 161
rect 0 108 17 125
rect 0 72 17 89
rect 0 36 17 53
rect 0 0 17 17
<< metal1 >>
rect -6 3545 23 3548
rect -6 3528 0 3545
rect 17 3528 23 3545
rect -6 3509 23 3528
rect -6 3492 0 3509
rect 17 3492 23 3509
rect -6 3473 23 3492
rect -6 3456 0 3473
rect 17 3456 23 3473
rect -6 3437 23 3456
rect -6 3420 0 3437
rect 17 3420 23 3437
rect -6 3401 23 3420
rect -6 3384 0 3401
rect 17 3384 23 3401
rect -6 3365 23 3384
rect -6 3348 0 3365
rect 17 3348 23 3365
rect -6 3329 23 3348
rect -6 3312 0 3329
rect 17 3312 23 3329
rect -6 3293 23 3312
rect -6 3276 0 3293
rect 17 3276 23 3293
rect -6 3257 23 3276
rect -6 3240 0 3257
rect 17 3240 23 3257
rect -6 3221 23 3240
rect -6 3204 0 3221
rect 17 3204 23 3221
rect -6 3185 23 3204
rect -6 3168 0 3185
rect 17 3168 23 3185
rect -6 3149 23 3168
rect -6 3132 0 3149
rect 17 3132 23 3149
rect -6 3113 23 3132
rect -6 3096 0 3113
rect 17 3096 23 3113
rect -6 3077 23 3096
rect -6 3060 0 3077
rect 17 3060 23 3077
rect -6 3041 23 3060
rect -6 3024 0 3041
rect 17 3024 23 3041
rect -6 3005 23 3024
rect -6 2988 0 3005
rect 17 2988 23 3005
rect -6 2969 23 2988
rect -6 2952 0 2969
rect 17 2952 23 2969
rect -6 2933 23 2952
rect -6 2916 0 2933
rect 17 2916 23 2933
rect -6 2897 23 2916
rect -6 2880 0 2897
rect 17 2880 23 2897
rect -6 2861 23 2880
rect -6 2844 0 2861
rect 17 2844 23 2861
rect -6 2825 23 2844
rect -6 2808 0 2825
rect 17 2808 23 2825
rect -6 2789 23 2808
rect -6 2772 0 2789
rect 17 2772 23 2789
rect -6 2753 23 2772
rect -6 2736 0 2753
rect 17 2736 23 2753
rect -6 2717 23 2736
rect -6 2700 0 2717
rect 17 2700 23 2717
rect -6 2681 23 2700
rect -6 2664 0 2681
rect 17 2664 23 2681
rect -6 2645 23 2664
rect -6 2628 0 2645
rect 17 2628 23 2645
rect -6 2609 23 2628
rect -6 2592 0 2609
rect 17 2592 23 2609
rect -6 2573 23 2592
rect -6 2556 0 2573
rect 17 2556 23 2573
rect -6 2537 23 2556
rect -6 2520 0 2537
rect 17 2520 23 2537
rect -6 2501 23 2520
rect -6 2484 0 2501
rect 17 2484 23 2501
rect -6 2465 23 2484
rect -6 2448 0 2465
rect 17 2448 23 2465
rect -6 2429 23 2448
rect -6 2412 0 2429
rect 17 2412 23 2429
rect -6 2393 23 2412
rect -6 2376 0 2393
rect 17 2376 23 2393
rect -6 2357 23 2376
rect -6 2340 0 2357
rect 17 2340 23 2357
rect -6 2321 23 2340
rect -6 2304 0 2321
rect 17 2304 23 2321
rect -6 2285 23 2304
rect -6 2268 0 2285
rect 17 2268 23 2285
rect -6 2249 23 2268
rect -6 2232 0 2249
rect 17 2232 23 2249
rect -6 2213 23 2232
rect -6 2196 0 2213
rect 17 2196 23 2213
rect -6 2177 23 2196
rect -6 2160 0 2177
rect 17 2160 23 2177
rect -6 2141 23 2160
rect -6 2124 0 2141
rect 17 2124 23 2141
rect -6 2105 23 2124
rect -6 2088 0 2105
rect 17 2088 23 2105
rect -6 2069 23 2088
rect -6 2052 0 2069
rect 17 2052 23 2069
rect -6 2033 23 2052
rect -6 2016 0 2033
rect 17 2016 23 2033
rect -6 1997 23 2016
rect -6 1980 0 1997
rect 17 1980 23 1997
rect -6 1961 23 1980
rect -6 1944 0 1961
rect 17 1944 23 1961
rect -6 1925 23 1944
rect -6 1908 0 1925
rect 17 1908 23 1925
rect -6 1889 23 1908
rect -6 1872 0 1889
rect 17 1872 23 1889
rect -6 1853 23 1872
rect -6 1836 0 1853
rect 17 1836 23 1853
rect -6 1817 23 1836
rect -6 1800 0 1817
rect 17 1800 23 1817
rect -6 1781 23 1800
rect -6 1764 0 1781
rect 17 1764 23 1781
rect -6 1745 23 1764
rect -6 1728 0 1745
rect 17 1728 23 1745
rect -6 1709 23 1728
rect -6 1692 0 1709
rect 17 1692 23 1709
rect -6 1673 23 1692
rect -6 1656 0 1673
rect 17 1656 23 1673
rect -6 1637 23 1656
rect -6 1620 0 1637
rect 17 1620 23 1637
rect -6 1601 23 1620
rect -6 1584 0 1601
rect 17 1584 23 1601
rect -6 1565 23 1584
rect -6 1548 0 1565
rect 17 1548 23 1565
rect -6 1529 23 1548
rect -6 1512 0 1529
rect 17 1512 23 1529
rect -6 1493 23 1512
rect -6 1476 0 1493
rect 17 1476 23 1493
rect -6 1457 23 1476
rect -6 1440 0 1457
rect 17 1440 23 1457
rect -6 1421 23 1440
rect -6 1404 0 1421
rect 17 1404 23 1421
rect -6 1385 23 1404
rect -6 1368 0 1385
rect 17 1368 23 1385
rect -6 1349 23 1368
rect -6 1332 0 1349
rect 17 1332 23 1349
rect -6 1313 23 1332
rect -6 1296 0 1313
rect 17 1296 23 1313
rect -6 1277 23 1296
rect -6 1260 0 1277
rect 17 1260 23 1277
rect -6 1241 23 1260
rect -6 1224 0 1241
rect 17 1224 23 1241
rect -6 1205 23 1224
rect -6 1188 0 1205
rect 17 1188 23 1205
rect -6 1169 23 1188
rect -6 1152 0 1169
rect 17 1152 23 1169
rect -6 1133 23 1152
rect -6 1116 0 1133
rect 17 1116 23 1133
rect -6 1097 23 1116
rect -6 1080 0 1097
rect 17 1080 23 1097
rect -6 1061 23 1080
rect -6 1044 0 1061
rect 17 1044 23 1061
rect -6 1025 23 1044
rect -6 1008 0 1025
rect 17 1008 23 1025
rect -6 989 23 1008
rect -6 972 0 989
rect 17 972 23 989
rect -6 953 23 972
rect -6 936 0 953
rect 17 936 23 953
rect -6 917 23 936
rect -6 900 0 917
rect 17 900 23 917
rect -6 881 23 900
rect -6 864 0 881
rect 17 864 23 881
rect -6 845 23 864
rect -6 828 0 845
rect 17 828 23 845
rect -6 809 23 828
rect -6 792 0 809
rect 17 792 23 809
rect -6 773 23 792
rect -6 756 0 773
rect 17 756 23 773
rect -6 737 23 756
rect -6 720 0 737
rect 17 720 23 737
rect -6 701 23 720
rect -6 684 0 701
rect 17 684 23 701
rect -6 665 23 684
rect -6 648 0 665
rect 17 648 23 665
rect -6 629 23 648
rect -6 612 0 629
rect 17 612 23 629
rect -6 593 23 612
rect -6 576 0 593
rect 17 576 23 593
rect -6 557 23 576
rect -6 540 0 557
rect 17 540 23 557
rect -6 521 23 540
rect -6 504 0 521
rect 17 504 23 521
rect -6 485 23 504
rect -6 468 0 485
rect 17 468 23 485
rect -6 449 23 468
rect -6 432 0 449
rect 17 432 23 449
rect -6 413 23 432
rect -6 396 0 413
rect 17 396 23 413
rect -6 377 23 396
rect -6 360 0 377
rect 17 360 23 377
rect -6 341 23 360
rect -6 324 0 341
rect 17 324 23 341
rect -6 305 23 324
rect -6 288 0 305
rect 17 288 23 305
rect -6 269 23 288
rect -6 252 0 269
rect 17 252 23 269
rect -6 233 23 252
rect -6 216 0 233
rect 17 216 23 233
rect -6 197 23 216
rect -6 180 0 197
rect 17 180 23 197
rect -6 161 23 180
rect -6 144 0 161
rect 17 144 23 161
rect -6 125 23 144
rect -6 108 0 125
rect 17 108 23 125
rect -6 89 23 108
rect -6 72 0 89
rect 17 72 23 89
rect -6 53 23 72
rect -6 36 0 53
rect 17 36 23 53
rect -6 17 23 36
rect -6 0 0 17
rect 17 0 23 17
rect -6 -3 23 0
<< properties >>
string GDS_END 80287718
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 80281250
<< end >>
