magic
tech sky130B
timestamp 1707688321
<< metal1 >>
rect 0 0 3 122
rect 125 0 128 122
<< via1 >>
rect 3 0 125 122
<< metal2 >>
rect 0 0 3 122
rect 125 0 128 122
<< properties >>
string GDS_END 79747674
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 79746518
<< end >>
