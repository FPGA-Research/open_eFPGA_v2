magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< viali >>
rect -89 -17 17 4913
<< metal1 >>
rect -101 4913 29 4925
rect -101 -17 -89 4913
rect 17 -17 29 4913
rect -101 -29 29 -17
<< properties >>
string GDS_END 13753890
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 13744926
<< end >>
