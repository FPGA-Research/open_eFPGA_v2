magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect 832 1425 1387 1467
rect 802 1293 1387 1425
rect 832 1251 1387 1293
<< mvnsubdiff >>
rect 838 1376 1121 1389
rect 838 1342 862 1376
rect 896 1342 930 1376
rect 964 1342 998 1376
rect 1032 1342 1121 1376
rect 838 1329 1121 1342
<< mvnsubdiffcont >>
rect 862 1342 896 1376
rect 930 1342 964 1376
rect 998 1342 1032 1376
<< poly >>
rect 403 1483 537 1499
rect 403 1449 419 1483
rect 453 1449 487 1483
rect 521 1449 537 1483
rect 403 1433 537 1449
rect 593 1269 727 1285
rect 593 1235 609 1269
rect 643 1235 677 1269
rect 711 1235 727 1269
rect 593 1219 727 1235
rect 107 1118 403 1134
rect 107 1084 123 1118
rect 157 1084 200 1118
rect 234 1084 277 1118
rect 311 1084 353 1118
rect 387 1084 403 1118
rect 107 1068 403 1084
rect 459 1118 755 1134
rect 459 1084 475 1118
rect 509 1084 552 1118
rect 586 1084 629 1118
rect 663 1084 705 1118
rect 739 1084 755 1118
rect 459 1068 755 1084
rect 1942 814 2238 830
rect 1942 780 1958 814
rect 1992 780 2034 814
rect 2068 780 2111 814
rect 2145 780 2188 814
rect 2222 780 2238 814
rect 1942 764 2238 780
rect 1942 372 2062 764
<< polycont >>
rect 419 1449 453 1483
rect 487 1449 521 1483
rect 609 1235 643 1269
rect 677 1235 711 1269
rect 123 1084 157 1118
rect 200 1084 234 1118
rect 277 1084 311 1118
rect 353 1084 387 1118
rect 475 1084 509 1118
rect 552 1084 586 1118
rect 629 1084 663 1118
rect 705 1084 739 1118
rect 1958 780 1992 814
rect 2034 780 2068 814
rect 2111 780 2145 814
rect 2188 780 2222 814
<< locali >>
rect 403 1489 793 1519
rect 403 1455 404 1489
rect 438 1483 476 1489
rect 510 1483 793 1489
rect 453 1455 476 1483
rect 403 1449 419 1455
rect 453 1449 487 1455
rect 521 1449 793 1483
rect 341 1362 432 1379
rect 341 1328 357 1362
rect 391 1328 432 1362
rect 341 1290 432 1328
rect 548 1340 582 1378
rect 686 1313 793 1449
rect 1776 1432 1820 1466
rect 1854 1432 1898 1466
rect 1742 1394 1932 1432
rect 838 1376 1121 1389
rect 896 1342 921 1376
rect 964 1342 998 1376
rect 1038 1342 1087 1376
rect 838 1329 1121 1342
rect 1776 1360 1820 1394
rect 1854 1360 1898 1394
rect 1742 1322 1932 1360
rect 341 1256 357 1290
rect 391 1269 432 1290
rect 1776 1288 1820 1322
rect 1854 1288 1898 1322
rect 391 1256 609 1269
rect 341 1235 609 1256
rect 643 1235 677 1269
rect 711 1235 727 1269
rect 1742 1250 1932 1288
rect 1776 1216 1820 1250
rect 1854 1216 1898 1250
rect 2249 1394 2283 1432
rect 2249 1322 2283 1360
rect 2249 1250 2283 1288
rect 107 1164 741 1198
rect 775 1164 813 1198
rect 107 1118 403 1164
rect 107 1084 123 1118
rect 157 1084 200 1118
rect 234 1084 277 1118
rect 311 1084 353 1118
rect 387 1084 403 1118
rect 459 1084 475 1118
rect 509 1084 552 1118
rect 586 1084 629 1118
rect 673 1084 705 1118
rect 745 1084 755 1118
rect 2073 958 2107 996
rect 238 769 272 811
rect 238 693 272 735
rect 238 617 272 659
rect 238 541 272 583
rect 590 766 624 811
rect 1935 780 1958 814
rect 2007 780 2034 814
rect 2068 780 2111 814
rect 2145 780 2188 814
rect 2222 780 2238 814
rect 590 687 624 732
rect 590 607 624 653
rect 238 464 272 507
rect 62 210 96 248
rect 62 138 96 176
rect 62 66 96 104
rect 414 210 448 248
rect 414 138 448 176
rect 414 66 448 104
rect 766 210 800 248
rect 766 138 800 176
rect 766 66 800 104
rect 1821 248 1897 282
rect 1787 210 1931 248
rect 1821 176 1897 210
rect 1787 138 1931 176
rect 1821 104 1897 138
rect 2073 144 2107 182
rect 1787 66 1931 104
rect 1821 32 1897 66
<< viali >>
rect 404 1483 438 1489
rect 476 1483 510 1489
rect 404 1455 419 1483
rect 419 1455 438 1483
rect 476 1455 487 1483
rect 487 1455 510 1483
rect 357 1328 391 1362
rect 548 1378 582 1412
rect 548 1306 582 1340
rect 1742 1432 1776 1466
rect 1820 1432 1854 1466
rect 1898 1432 1932 1466
rect 838 1342 862 1376
rect 862 1342 872 1376
rect 921 1342 930 1376
rect 930 1342 955 1376
rect 1004 1342 1032 1376
rect 1032 1342 1038 1376
rect 1087 1342 1121 1376
rect 1742 1360 1776 1394
rect 1820 1360 1854 1394
rect 1898 1360 1932 1394
rect 357 1256 391 1290
rect 1742 1288 1776 1322
rect 1820 1288 1854 1322
rect 1898 1288 1932 1322
rect 1742 1216 1776 1250
rect 1820 1216 1854 1250
rect 1898 1216 1932 1250
rect 2249 1432 2283 1466
rect 2249 1360 2283 1394
rect 2249 1288 2283 1322
rect 2249 1216 2283 1250
rect 741 1164 775 1198
rect 813 1164 847 1198
rect 639 1084 663 1118
rect 663 1084 673 1118
rect 711 1084 739 1118
rect 739 1084 745 1118
rect 2073 996 2107 1030
rect 2073 924 2107 958
rect 238 811 272 845
rect 238 735 272 769
rect 238 659 272 693
rect 238 583 272 617
rect 590 811 624 845
rect 1901 780 1935 814
rect 1973 780 1992 814
rect 1992 780 2007 814
rect 590 732 624 766
rect 590 653 624 687
rect 590 573 624 607
rect 238 507 272 541
rect 238 430 272 464
rect 62 248 96 282
rect 62 176 96 210
rect 62 104 96 138
rect 62 32 96 66
rect 414 248 448 282
rect 414 176 448 210
rect 414 104 448 138
rect 414 32 448 66
rect 766 248 800 282
rect 766 176 800 210
rect 766 104 800 138
rect 766 32 800 66
rect 1787 248 1821 282
rect 1897 248 1931 282
rect 1787 176 1821 210
rect 1897 176 1931 210
rect 1787 104 1821 138
rect 1897 104 1931 138
rect 2073 182 2107 216
rect 2073 110 2107 144
rect 1787 32 1821 66
rect 1897 32 1931 66
<< metal1 >>
rect 392 1489 522 1495
rect 392 1455 404 1489
rect 438 1455 476 1489
rect 510 1455 522 1489
tri 1146 1466 1158 1478 se
rect 1158 1466 2289 1478
rect 392 1449 522 1455
tri 1129 1449 1146 1466 se
rect 1146 1449 1742 1466
rect 351 1362 397 1376
rect 351 1328 357 1362
rect 391 1328 397 1362
rect 351 1290 397 1328
rect 351 1256 357 1290
rect 391 1256 397 1290
tri 331 1044 351 1064 se
rect 351 1044 397 1256
tri 317 1030 331 1044 se
rect 331 1030 383 1044
tri 383 1030 397 1044 nw
rect 464 1053 510 1449
tri 1112 1432 1129 1449 se
rect 1129 1432 1742 1449
rect 1776 1432 1820 1466
rect 1854 1432 1898 1466
rect 1932 1432 2249 1466
rect 2283 1432 2289 1466
tri 1104 1424 1112 1432 se
rect 1112 1424 2289 1432
rect 542 1412 2289 1424
rect 542 1378 548 1412
rect 582 1394 2289 1412
rect 582 1378 1742 1394
rect 542 1376 1742 1378
rect 542 1342 838 1376
rect 872 1342 921 1376
rect 955 1342 1004 1376
rect 1038 1342 1087 1376
rect 1121 1360 1742 1376
rect 1776 1360 1820 1394
rect 1854 1360 1898 1394
rect 1932 1360 2249 1394
rect 2283 1360 2289 1394
rect 1121 1342 2289 1360
rect 542 1340 2289 1342
rect 542 1306 548 1340
rect 582 1322 2289 1340
rect 582 1306 1742 1322
rect 542 1294 1742 1306
tri 1068 1288 1074 1294 ne
rect 1074 1288 1742 1294
rect 1776 1288 1820 1322
rect 1854 1288 1898 1322
rect 1932 1288 2249 1322
rect 2283 1288 2289 1322
tri 1074 1250 1112 1288 ne
rect 1112 1250 2289 1288
tri 1112 1216 1146 1250 ne
rect 1146 1216 1742 1250
rect 1776 1216 1820 1250
rect 1854 1216 1898 1250
rect 1932 1216 2249 1250
rect 2283 1216 2289 1250
tri 1146 1204 1158 1216 ne
rect 1158 1204 2289 1216
rect 729 1198 859 1204
rect 729 1164 741 1198
rect 775 1164 813 1198
rect 847 1164 859 1198
rect 729 1158 859 1164
rect 627 1118 757 1124
rect 627 1084 639 1118
rect 673 1084 711 1118
rect 745 1084 757 1118
rect 627 1078 757 1084
tri 464 1030 487 1053 ne
rect 487 1030 510 1053
tri 510 1030 553 1073 sw
rect 2067 1030 2113 1042
tri 283 996 317 1030 se
rect 317 1019 372 1030
tri 372 1019 383 1030 nw
tri 487 1019 498 1030 ne
rect 498 1019 553 1030
tri 553 1019 564 1030 sw
rect 317 1007 360 1019
tri 360 1007 372 1019 nw
tri 498 1007 510 1019 ne
rect 510 1007 564 1019
rect 317 996 349 1007
tri 349 996 360 1007 nw
tri 510 996 521 1007 ne
rect 521 996 564 1007
tri 564 996 587 1019 sw
rect 2067 996 2073 1030
rect 2107 996 2113 1030
tri 278 991 283 996 se
rect 283 991 344 996
tri 344 991 349 996 nw
tri 521 991 526 996 ne
rect 526 991 587 996
tri 245 958 278 991 se
rect 278 958 311 991
tri 311 958 344 991 nw
tri 526 958 559 991 ne
rect 559 958 587 991
tri 587 958 625 996 sw
rect 2067 958 2113 996
tri 232 945 245 958 se
rect 245 953 306 958
tri 306 953 311 958 nw
tri 559 953 564 958 ne
rect 564 953 625 958
tri 625 953 630 958 sw
rect 245 945 286 953
rect 232 933 286 945
tri 286 933 306 953 nw
tri 564 933 584 953 ne
rect 232 845 278 933
tri 278 925 286 933 nw
rect 232 811 238 845
rect 272 811 278 845
rect 232 769 278 811
rect 232 735 238 769
rect 272 735 278 769
rect 232 693 278 735
rect 232 659 238 693
rect 272 659 278 693
rect 232 617 278 659
rect 232 583 238 617
rect 272 583 278 617
rect 232 541 278 583
rect 584 845 630 953
rect 584 811 590 845
rect 624 811 630 845
rect 2067 924 2073 958
rect 2107 924 2113 958
tri 1658 814 1664 820 se
rect 1664 814 2019 820
rect 584 766 630 811
tri 1624 780 1658 814 se
rect 1658 780 1901 814
rect 1935 780 1973 814
rect 2007 780 2019 814
rect 584 732 590 766
rect 624 732 630 766
tri 1598 754 1624 780 se
rect 1624 774 2019 780
rect 1624 754 1664 774
tri 1664 754 1684 774 nw
rect 584 687 630 732
rect 584 653 590 687
rect 624 653 630 687
rect 584 607 630 653
rect 584 573 590 607
rect 624 573 630 607
rect 584 561 630 573
tri 1580 736 1598 754 se
rect 1598 736 1646 754
tri 1646 736 1664 754 nw
rect 232 507 238 541
rect 272 507 278 541
rect 232 464 278 507
rect 232 430 238 464
rect 272 430 278 464
tri 1514 431 1580 497 se
rect 1580 477 1626 736
tri 1626 716 1646 736 nw
tri 1580 431 1626 477 nw
rect 232 419 278 430
tri 1502 419 1514 431 se
rect 1514 419 1568 431
tri 1568 419 1580 431 nw
rect 232 373 1522 419
tri 1522 373 1568 419 nw
rect 48 282 1937 294
rect 48 248 62 282
rect 96 248 414 282
rect 448 248 766 282
rect 800 248 1787 282
rect 1821 248 1897 282
rect 1931 248 1937 282
rect 48 210 1937 248
rect 48 176 62 210
rect 96 176 414 210
rect 448 176 766 210
rect 800 176 1787 210
rect 1821 176 1897 210
rect 1931 176 1937 210
rect 48 138 1937 176
rect 48 104 62 138
rect 96 104 414 138
rect 448 104 766 138
rect 800 104 1787 138
rect 1821 104 1897 138
rect 1931 104 1937 138
rect 48 66 1937 104
rect 2067 216 2113 924
rect 2067 182 2073 216
rect 2107 182 2113 216
rect 2067 144 2113 182
rect 2067 110 2073 144
rect 2107 110 2113 144
rect 2067 98 2113 110
rect 48 32 62 66
rect 96 32 414 66
rect 448 32 766 66
rect 800 32 1787 66
rect 1821 32 1897 66
rect 1931 32 1937 66
rect 48 20 1937 32
use nfet_CDNS_52468879185919  nfet_CDNS_52468879185919_0
timestamp 1707688321
transform 1 0 459 0 1 36
box -79 -32 522 1032
use nfet_CDNS_52468879185921  nfet_CDNS_52468879185921_0
timestamp 1707688321
transform 1 0 107 0 1 36
box -79 -32 375 1032
use nfet_CDNS_52468879185922  nfet_CDNS_52468879185922_0
timestamp 1707688321
transform -1 0 2062 0 1 -260
box -79 -32 346 632
use pfet_CDNS_52468879185918  pfet_CDNS_52468879185918_0
timestamp 1707688321
transform -1 0 537 0 1 1317
box -119 -66 239 150
use pfet_CDNS_52468879185918  pfet_CDNS_52468879185918_1
timestamp 1707688321
transform 1 0 593 0 1 1317
box -119 -66 239 150
use pfet_CDNS_52468879185925  pfet_CDNS_52468879185925_0
timestamp 1707688321
transform -1 0 2238 0 -1 1462
box -266 -66 562 666
<< labels >>
flabel metal1 s 1721 1309 1857 1430 0 FreeSans 200 0 0 0 vswitch
port 1 nsew
flabel metal1 s 695 123 766 209 0 FreeSans 200 0 0 0 vssa
port 2 nsew
flabel metal1 s 2072 638 2109 707 0 FreeSans 200 90 0 0 out_h
port 3 nsew
<< properties >>
string GDS_END 80531114
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 80520896
string path 20.300 33.975 28.675 33.975 
<< end >>
