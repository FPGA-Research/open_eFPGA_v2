magic
tech sky130A
timestamp 1707688321
<< properties >>
string GDS_END 17354026
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 17353638
<< end >>
