magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< pwell >>
rect 39 123 335 799
rect 1587 663 2190 799
rect 2700 663 2999 799
rect 1587 349 1883 663
rect 1587 123 2190 349
rect 2500 123 2799 349
rect 39 37 3376 123
<< mvndiff >>
rect 65 173 283 773
rect 1639 173 1857 773
rect 1917 735 2138 773
rect 1917 701 2104 735
rect 1917 689 2138 701
rect 2752 735 2973 773
rect 2786 701 2973 735
rect 2752 689 2973 701
rect 1917 173 2138 323
rect 2552 173 2773 323
<< mvndiffc >>
rect 2104 701 2138 735
rect 2752 701 2786 735
<< mvpsubdiff >>
rect 65 63 89 97
rect 123 63 158 97
rect 192 63 227 97
rect 261 63 296 97
rect 330 63 365 97
rect 399 63 434 97
rect 468 63 503 97
rect 537 63 572 97
rect 606 63 640 97
rect 674 63 708 97
rect 742 63 776 97
rect 810 63 844 97
rect 878 63 912 97
rect 946 63 980 97
rect 1014 63 1048 97
rect 1082 63 1116 97
rect 1150 63 1184 97
rect 1218 63 1252 97
rect 1286 63 1320 97
rect 1354 63 1388 97
rect 1422 63 1456 97
rect 1490 63 1524 97
rect 1558 63 1592 97
rect 1626 63 1660 97
rect 1694 63 1728 97
rect 1762 63 1796 97
rect 1830 63 1864 97
rect 1898 63 1932 97
rect 1966 63 2000 97
rect 2034 63 2068 97
rect 2102 63 2136 97
rect 2170 63 2204 97
rect 2238 63 2272 97
rect 2306 63 2340 97
rect 2374 63 2408 97
rect 2442 63 2476 97
rect 2510 63 2544 97
rect 2578 63 2612 97
rect 2646 63 2680 97
rect 2714 63 2748 97
rect 2782 63 2816 97
rect 2850 63 2884 97
rect 2918 63 2952 97
rect 2986 63 3020 97
rect 3054 63 3088 97
rect 3122 63 3156 97
rect 3190 63 3224 97
rect 3258 63 3292 97
rect 3326 63 3350 97
<< mvpsubdiffcont >>
rect 89 63 123 97
rect 158 63 192 97
rect 227 63 261 97
rect 296 63 330 97
rect 365 63 399 97
rect 434 63 468 97
rect 503 63 537 97
rect 572 63 606 97
rect 640 63 674 97
rect 708 63 742 97
rect 776 63 810 97
rect 844 63 878 97
rect 912 63 946 97
rect 980 63 1014 97
rect 1048 63 1082 97
rect 1116 63 1150 97
rect 1184 63 1218 97
rect 1252 63 1286 97
rect 1320 63 1354 97
rect 1388 63 1422 97
rect 1456 63 1490 97
rect 1524 63 1558 97
rect 1592 63 1626 97
rect 1660 63 1694 97
rect 1728 63 1762 97
rect 1796 63 1830 97
rect 1864 63 1898 97
rect 1932 63 1966 97
rect 2000 63 2034 97
rect 2068 63 2102 97
rect 2136 63 2170 97
rect 2204 63 2238 97
rect 2272 63 2306 97
rect 2340 63 2374 97
rect 2408 63 2442 97
rect 2476 63 2510 97
rect 2544 63 2578 97
rect 2612 63 2646 97
rect 2680 63 2714 97
rect 2748 63 2782 97
rect 2816 63 2850 97
rect 2884 63 2918 97
rect 2952 63 2986 97
rect 3020 63 3054 97
rect 3088 63 3122 97
rect 3156 63 3190 97
rect 3224 63 3258 97
rect 3292 63 3326 97
<< poly >>
rect 365 855 777 871
rect 365 821 381 855
rect 415 821 451 855
rect 485 821 520 855
rect 554 821 589 855
rect 623 821 658 855
rect 692 821 727 855
rect 761 821 777 855
rect 365 805 777 821
rect 833 855 1089 871
rect 833 821 849 855
rect 883 821 944 855
rect 978 821 1039 855
rect 1073 821 1089 855
rect 833 805 1089 821
rect 1145 855 1557 871
rect 1145 821 1161 855
rect 1195 821 1231 855
rect 1265 821 1300 855
rect 1334 821 1369 855
rect 1403 821 1438 855
rect 1472 821 1507 855
rect 1541 821 1557 855
rect 1145 805 1557 821
rect 3086 855 3246 871
rect 3086 821 3102 855
rect 3136 821 3196 855
rect 3230 821 3246 855
rect 3086 805 3246 821
rect 2217 641 2417 657
rect 2217 607 2233 641
rect 2267 607 2367 641
rect 2401 607 2417 641
rect 2217 591 2417 607
rect 2473 641 2673 657
rect 2473 607 2489 641
rect 2523 607 2623 641
rect 2657 607 2673 641
rect 2473 591 2673 607
rect 2183 405 2317 421
rect 2183 371 2199 405
rect 2233 371 2267 405
rect 2301 371 2317 405
rect 2183 355 2317 371
rect 2373 405 2507 421
rect 2373 371 2389 405
rect 2423 371 2457 405
rect 2491 371 2507 405
rect 2373 355 2507 371
rect 2997 405 3131 421
rect 2997 371 3013 405
rect 3047 371 3081 405
rect 3115 371 3131 405
rect 2997 355 3131 371
rect 3187 405 3321 421
rect 3187 371 3203 405
rect 3237 371 3271 405
rect 3305 371 3321 405
rect 3187 355 3321 371
<< polycont >>
rect 381 821 415 855
rect 451 821 485 855
rect 520 821 554 855
rect 589 821 623 855
rect 658 821 692 855
rect 727 821 761 855
rect 849 821 883 855
rect 944 821 978 855
rect 1039 821 1073 855
rect 1161 821 1195 855
rect 1231 821 1265 855
rect 1300 821 1334 855
rect 1369 821 1403 855
rect 1438 821 1472 855
rect 1507 821 1541 855
rect 3102 821 3136 855
rect 3196 821 3230 855
rect 2233 607 2267 641
rect 2367 607 2401 641
rect 2489 607 2523 641
rect 2623 607 2657 641
rect 2199 371 2233 405
rect 2267 371 2301 405
rect 2389 371 2423 405
rect 2457 371 2491 405
rect 3013 371 3047 405
rect 3081 371 3115 405
rect 3203 371 3237 405
rect 3271 371 3305 405
<< locali >>
rect 365 821 381 855
rect 436 821 451 855
rect 512 821 520 855
rect 588 821 589 855
rect 623 821 630 855
rect 692 821 707 855
rect 761 821 777 855
rect 833 821 849 855
rect 889 821 936 855
rect 978 821 1016 855
rect 1073 821 1089 855
rect 1145 821 1161 855
rect 1214 821 1231 855
rect 1290 821 1300 855
rect 1366 821 1369 855
rect 1403 821 1407 855
rect 1472 821 1482 855
rect 1541 821 1557 855
rect 3086 821 3102 855
rect 3140 821 3178 855
rect 3230 821 3246 855
rect 2128 767 2166 801
rect 2200 767 2206 801
rect 320 673 354 715
rect 320 597 354 639
rect 632 672 666 715
rect 320 521 354 563
rect 320 445 354 487
rect 320 369 354 411
rect 320 292 354 335
rect 320 215 354 258
rect 476 551 510 595
rect 476 472 510 517
rect 476 393 510 438
rect 476 314 510 359
rect 632 595 666 638
rect 632 518 666 561
rect 632 441 666 484
rect 632 363 666 407
rect 788 686 822 727
rect 788 611 822 652
rect 788 536 822 577
rect 788 461 822 502
rect 788 386 822 427
rect 476 235 510 280
rect 788 311 822 352
rect 788 235 822 277
rect 944 670 978 709
rect 944 597 978 636
rect 944 524 978 563
rect 944 451 978 490
rect 944 378 978 417
rect 944 305 978 344
rect 944 231 978 271
rect 1100 686 1134 727
rect 1100 611 1134 652
rect 1100 535 1134 577
rect 1100 459 1134 501
rect 1100 383 1134 425
rect 1256 670 1290 715
rect 1256 590 1290 636
rect 1568 673 1602 715
rect 2104 735 2206 767
rect 2138 701 2206 735
rect 2104 685 2206 701
rect 2428 723 2462 761
rect 2684 751 2718 761
rect 2684 735 2786 751
rect 2684 723 2752 735
rect 2718 701 2752 723
rect 2718 689 2786 701
rect 2706 685 2786 689
rect 1256 510 1290 556
rect 1256 430 1290 476
rect 1412 556 1446 595
rect 1412 483 1446 522
rect 1412 410 1446 449
rect 1100 307 1134 349
rect 1100 231 1134 273
rect 1412 337 1446 376
rect 1412 263 1446 303
rect 1412 189 1446 229
rect 1568 597 1602 639
rect 2217 607 2233 641
rect 2297 607 2335 641
rect 2401 607 2417 641
rect 2473 607 2489 641
rect 2523 607 2532 641
rect 2566 607 2604 641
rect 2657 607 2673 641
rect 3041 619 3075 727
rect 3257 619 3291 727
rect 1568 521 1602 563
rect 1568 445 1602 487
rect 1568 369 1602 411
rect 3043 405 3081 406
rect 2183 371 2193 405
rect 2233 371 2265 405
rect 2301 371 2317 405
rect 2373 371 2385 405
rect 2423 371 2457 405
rect 2491 371 2507 405
rect 2997 372 3009 405
rect 2997 371 3013 372
rect 3047 371 3081 405
rect 3115 371 3131 405
rect 3187 371 3199 405
rect 3237 371 3271 405
rect 3305 371 3321 405
rect 1568 292 1602 335
rect 1568 215 1602 258
rect 2172 207 2206 245
rect 2328 207 2362 245
rect 2484 207 2518 245
rect 2986 207 3020 245
rect 3142 207 3176 245
rect 3298 207 3332 245
rect 123 63 138 97
rect 192 63 211 97
rect 261 63 284 97
rect 330 63 357 97
rect 399 63 430 97
rect 468 63 503 97
rect 537 63 572 97
rect 610 63 640 97
rect 683 63 708 97
rect 756 63 776 97
rect 829 63 844 97
rect 902 63 912 97
rect 974 63 980 97
rect 1046 63 1048 97
rect 1082 63 1084 97
rect 1150 63 1156 97
rect 1218 63 1228 97
rect 1286 63 1300 97
rect 1354 63 1372 97
rect 1422 63 1444 97
rect 1490 63 1516 97
rect 1558 63 1588 97
rect 1626 63 1660 97
rect 1694 63 1728 97
rect 1766 63 1796 97
rect 1838 63 1864 97
rect 1910 63 1932 97
rect 1982 63 2000 97
rect 2054 63 2068 97
rect 2126 63 2136 97
rect 2198 63 2204 97
rect 2270 63 2272 97
rect 2306 63 2308 97
rect 2374 63 2380 97
rect 2442 63 2452 97
rect 2510 63 2524 97
rect 2578 63 2596 97
rect 2646 63 2668 97
rect 2714 63 2740 97
rect 2782 63 2812 97
rect 2850 63 2884 97
rect 2918 63 2952 97
rect 2990 63 3020 97
rect 3062 63 3088 97
rect 3134 63 3156 97
rect 3206 63 3224 97
rect 3278 63 3292 97
<< viali >>
rect 402 821 415 855
rect 415 821 436 855
rect 478 821 485 855
rect 485 821 512 855
rect 554 821 588 855
rect 630 821 658 855
rect 658 821 664 855
rect 707 821 727 855
rect 727 821 741 855
rect 855 821 883 855
rect 883 821 889 855
rect 936 821 944 855
rect 944 821 970 855
rect 1016 821 1039 855
rect 1039 821 1050 855
rect 1180 821 1195 855
rect 1195 821 1214 855
rect 1256 821 1265 855
rect 1265 821 1290 855
rect 1332 821 1334 855
rect 1334 821 1366 855
rect 1407 821 1438 855
rect 1438 821 1441 855
rect 1482 821 1507 855
rect 1507 821 1516 855
rect 3106 821 3136 855
rect 3136 821 3140 855
rect 3178 821 3196 855
rect 3196 821 3212 855
rect 2094 767 2128 801
rect 2166 767 2200 801
rect 320 715 354 749
rect 320 639 354 673
rect 632 715 666 749
rect 632 638 666 672
rect 320 563 354 597
rect 320 487 354 521
rect 320 411 354 445
rect 320 335 354 369
rect 320 258 354 292
rect 320 181 354 215
rect 476 595 510 629
rect 476 517 510 551
rect 476 438 510 472
rect 476 359 510 393
rect 632 561 666 595
rect 632 484 666 518
rect 632 407 666 441
rect 632 329 666 363
rect 788 727 822 761
rect 788 652 822 686
rect 788 577 822 611
rect 788 502 822 536
rect 788 427 822 461
rect 788 352 822 386
rect 476 280 510 314
rect 476 201 510 235
rect 788 277 822 311
rect 788 201 822 235
rect 944 709 978 743
rect 944 636 978 670
rect 944 563 978 597
rect 944 490 978 524
rect 944 417 978 451
rect 944 344 978 378
rect 944 271 978 305
rect 944 197 978 231
rect 1100 727 1134 761
rect 1100 652 1134 686
rect 1100 577 1134 611
rect 1100 501 1134 535
rect 1100 425 1134 459
rect 1256 715 1290 749
rect 1256 636 1290 670
rect 1568 715 1602 749
rect 2428 761 2462 795
rect 2428 689 2462 723
rect 2684 761 2718 795
rect 2684 689 2718 723
rect 3041 727 3075 761
rect 1568 639 1602 673
rect 1256 556 1290 590
rect 1256 476 1290 510
rect 1256 396 1290 430
rect 1412 595 1446 629
rect 1412 522 1446 556
rect 1412 449 1446 483
rect 1100 349 1134 383
rect 1100 273 1134 307
rect 1100 197 1134 231
rect 1412 376 1446 410
rect 1412 303 1446 337
rect 1412 229 1446 263
rect 1412 155 1446 189
rect 2263 607 2267 641
rect 2267 607 2297 641
rect 2335 607 2367 641
rect 2367 607 2369 641
rect 2532 607 2566 641
rect 2604 607 2623 641
rect 2623 607 2638 641
rect 1568 563 1602 597
rect 3041 585 3075 619
rect 3257 727 3291 761
rect 3257 585 3291 619
rect 1568 487 1602 521
rect 1568 411 1602 445
rect 3009 405 3043 406
rect 3081 405 3115 406
rect 2193 371 2199 405
rect 2199 371 2227 405
rect 2265 371 2267 405
rect 2267 371 2299 405
rect 2385 371 2389 405
rect 2389 371 2419 405
rect 2457 371 2491 405
rect 3009 372 3013 405
rect 3013 372 3043 405
rect 3081 372 3115 405
rect 3199 371 3203 405
rect 3203 371 3233 405
rect 3271 371 3305 405
rect 1568 335 1602 369
rect 1568 258 1602 292
rect 1568 181 1602 215
rect 2172 245 2206 279
rect 2172 173 2206 207
rect 2328 245 2362 279
rect 2328 173 2362 207
rect 2484 245 2518 279
rect 2484 173 2518 207
rect 2986 245 3020 279
rect 2986 173 3020 207
rect 3142 245 3176 279
rect 3142 173 3176 207
rect 3298 245 3332 279
rect 3298 173 3332 207
rect 65 63 89 97
rect 89 63 99 97
rect 138 63 158 97
rect 158 63 172 97
rect 211 63 227 97
rect 227 63 245 97
rect 284 63 296 97
rect 296 63 318 97
rect 357 63 365 97
rect 365 63 391 97
rect 430 63 434 97
rect 434 63 464 97
rect 503 63 537 97
rect 576 63 606 97
rect 606 63 610 97
rect 649 63 674 97
rect 674 63 683 97
rect 722 63 742 97
rect 742 63 756 97
rect 795 63 810 97
rect 810 63 829 97
rect 868 63 878 97
rect 878 63 902 97
rect 940 63 946 97
rect 946 63 974 97
rect 1012 63 1014 97
rect 1014 63 1046 97
rect 1084 63 1116 97
rect 1116 63 1118 97
rect 1156 63 1184 97
rect 1184 63 1190 97
rect 1228 63 1252 97
rect 1252 63 1262 97
rect 1300 63 1320 97
rect 1320 63 1334 97
rect 1372 63 1388 97
rect 1388 63 1406 97
rect 1444 63 1456 97
rect 1456 63 1478 97
rect 1516 63 1524 97
rect 1524 63 1550 97
rect 1588 63 1592 97
rect 1592 63 1622 97
rect 1660 63 1694 97
rect 1732 63 1762 97
rect 1762 63 1766 97
rect 1804 63 1830 97
rect 1830 63 1838 97
rect 1876 63 1898 97
rect 1898 63 1910 97
rect 1948 63 1966 97
rect 1966 63 1982 97
rect 2020 63 2034 97
rect 2034 63 2054 97
rect 2092 63 2102 97
rect 2102 63 2126 97
rect 2164 63 2170 97
rect 2170 63 2198 97
rect 2236 63 2238 97
rect 2238 63 2270 97
rect 2308 63 2340 97
rect 2340 63 2342 97
rect 2380 63 2408 97
rect 2408 63 2414 97
rect 2452 63 2476 97
rect 2476 63 2486 97
rect 2524 63 2544 97
rect 2544 63 2558 97
rect 2596 63 2612 97
rect 2612 63 2630 97
rect 2668 63 2680 97
rect 2680 63 2702 97
rect 2740 63 2748 97
rect 2748 63 2774 97
rect 2812 63 2816 97
rect 2816 63 2846 97
rect 2884 63 2918 97
rect 2956 63 2986 97
rect 2986 63 2990 97
rect 3028 63 3054 97
rect 3054 63 3062 97
rect 3100 63 3122 97
rect 3122 63 3134 97
rect 3172 63 3190 97
rect 3190 63 3206 97
rect 3244 63 3258 97
rect 3258 63 3278 97
rect 3316 63 3326 97
rect 3326 63 3350 97
<< metal1 >>
rect 390 855 753 861
rect 390 821 402 855
rect 436 821 478 855
rect 512 821 554 855
rect 588 821 630 855
rect 664 821 707 855
rect 741 821 753 855
rect 390 815 753 821
rect 843 855 1066 861
rect 843 821 855 855
rect 889 821 936 855
rect 970 821 1016 855
rect 1050 821 1066 855
rect 843 815 1066 821
tri 667 801 681 815 ne
rect 681 801 753 815
tri 980 801 994 815 ne
rect 994 801 1066 815
tri 681 781 701 801 ne
rect 314 749 672 761
rect 314 715 320 749
rect 354 725 632 749
rect 354 715 550 725
rect 314 673 550 715
rect 602 673 614 725
rect 666 673 672 749
rect 314 639 320 673
rect 354 672 393 673
tri 393 672 394 673 nw
tri 592 672 593 673 ne
rect 593 672 672 673
rect 354 639 360 672
tri 360 639 393 672 nw
tri 593 641 624 672 ne
rect 624 641 632 672
rect 314 597 360 639
rect 314 563 320 597
rect 354 563 360 597
rect 314 521 360 563
rect 314 487 320 521
rect 354 487 360 521
rect 314 445 360 487
rect 314 411 320 445
rect 354 411 360 445
rect 314 369 360 411
rect 314 335 320 369
rect 354 335 360 369
rect 314 292 360 335
rect 314 258 320 292
rect 354 258 360 292
rect 314 215 360 258
rect 314 181 320 215
rect 354 181 360 215
rect 470 629 516 641
tri 624 639 626 641 ne
rect 470 595 476 629
rect 510 595 516 629
rect 470 551 516 595
rect 470 517 476 551
rect 510 517 516 551
rect 470 472 516 517
rect 470 438 476 472
rect 510 438 516 472
rect 470 393 516 438
rect 470 359 476 393
rect 510 359 516 393
rect 470 314 516 359
rect 626 638 632 641
rect 666 638 672 672
rect 626 595 672 638
rect 626 561 632 595
rect 666 561 672 595
rect 626 518 672 561
rect 626 484 632 518
rect 666 484 672 518
rect 626 441 672 484
rect 626 407 632 441
rect 666 407 672 441
rect 626 363 672 407
rect 626 329 632 363
rect 666 329 672 363
rect 701 484 753 801
tri 994 781 1014 801 ne
rect 701 420 753 432
rect 701 362 753 368
rect 782 761 828 773
rect 782 727 788 761
rect 822 727 828 761
rect 782 686 828 727
rect 782 652 788 686
rect 822 652 828 686
rect 782 611 828 652
rect 782 577 788 611
rect 822 577 828 611
rect 782 536 828 577
rect 782 502 788 536
rect 822 502 828 536
rect 782 461 828 502
rect 782 427 788 461
rect 822 427 828 461
rect 782 386 828 427
rect 470 280 476 314
rect 510 311 516 314
tri 516 311 528 323 sw
rect 626 317 672 329
rect 782 352 788 386
rect 822 352 828 386
tri 776 317 782 323 se
rect 782 317 828 352
tri 770 311 776 317 se
rect 776 311 828 317
rect 510 289 528 311
tri 528 289 550 311 sw
tri 748 289 770 311 se
rect 770 289 788 311
rect 510 280 788 289
rect 470 277 788 280
rect 822 277 828 311
rect 470 235 828 277
rect 470 201 476 235
rect 510 201 788 235
rect 822 201 828 235
rect 470 189 828 201
rect 938 743 984 755
rect 938 709 944 743
rect 978 709 984 743
rect 938 670 984 709
rect 938 636 944 670
rect 978 636 984 670
rect 938 597 984 636
rect 938 563 944 597
rect 978 563 984 597
rect 938 524 984 563
rect 938 490 944 524
rect 978 490 984 524
rect 938 451 984 490
rect 938 417 944 451
rect 978 417 984 451
rect 1014 567 1066 801
rect 1168 855 1528 861
rect 1168 821 1180 855
rect 1214 821 1256 855
rect 1290 821 1332 855
rect 1366 821 1407 855
rect 1441 821 1482 855
rect 1516 821 1528 855
rect 1168 815 1528 821
rect 3094 855 3224 861
rect 3094 821 3106 855
rect 3140 821 3178 855
rect 3212 821 3224 855
rect 3094 815 3224 821
rect 1168 801 1240 815
tri 1240 801 1254 815 nw
tri 3109 807 3117 815 ne
rect 3117 807 3195 815
rect 1014 503 1066 515
rect 1014 445 1066 451
rect 1094 761 1140 773
rect 1094 727 1100 761
rect 1134 727 1140 761
rect 1094 686 1140 727
rect 1094 652 1100 686
rect 1134 652 1140 686
rect 1094 611 1140 652
rect 1094 577 1100 611
rect 1134 577 1140 611
rect 1094 535 1140 577
rect 1094 501 1100 535
rect 1134 501 1140 535
rect 1094 459 1140 501
rect 938 378 984 417
rect 938 344 944 378
rect 978 344 984 378
rect 938 305 984 344
rect 938 271 944 305
rect 978 271 984 305
rect 938 231 984 271
rect 938 197 944 231
rect 978 197 984 231
rect 314 169 360 181
tri 904 103 938 137 se
rect 938 103 984 197
rect 1094 425 1100 459
rect 1134 425 1140 459
rect 1094 383 1140 425
rect 1094 349 1100 383
rect 1134 349 1140 383
rect 1094 307 1140 349
rect 1094 273 1100 307
rect 1134 273 1140 307
rect 1094 231 1140 273
rect 1168 337 1220 801
tri 1220 781 1240 801 nw
rect 1250 749 1608 761
rect 2082 755 2090 807
rect 2142 755 2154 807
rect 2206 755 2212 807
rect 2422 795 2468 807
rect 2422 761 2428 795
rect 2462 761 2468 795
tri 2420 755 2422 757 se
rect 2422 755 2468 761
rect 1250 675 1256 749
rect 1290 727 1568 749
rect 1308 675 1353 727
rect 1405 675 1450 727
rect 1502 675 1546 727
rect 1602 715 1608 749
tri 2392 727 2420 755 se
rect 2420 727 2468 755
tri 2388 723 2392 727 se
rect 2392 723 2468 727
rect 1598 675 1608 715
tri 1745 689 1779 723 se
rect 1779 689 2428 723
rect 2462 689 2468 723
tri 1733 677 1745 689 se
rect 1745 677 2468 689
rect 2516 755 2522 807
rect 2574 755 2586 807
rect 2638 755 2650 807
rect 1250 673 1608 675
rect 1250 670 1296 673
rect 1250 636 1256 670
rect 1290 636 1296 670
tri 1296 639 1330 673 nw
tri 1528 641 1560 673 ne
rect 1560 641 1568 673
rect 1250 590 1296 636
rect 1250 556 1256 590
rect 1290 556 1296 590
rect 1250 510 1296 556
rect 1250 476 1256 510
rect 1290 476 1296 510
rect 1250 430 1296 476
rect 1250 396 1256 430
rect 1290 396 1296 430
rect 1250 384 1296 396
rect 1406 629 1452 641
tri 1560 639 1562 641 ne
rect 1562 639 1568 641
rect 1602 639 1608 673
rect 1406 595 1412 629
rect 1446 595 1452 629
rect 1406 556 1452 595
rect 1406 522 1412 556
rect 1446 522 1452 556
rect 1406 483 1452 522
rect 1406 449 1412 483
rect 1446 449 1452 483
rect 1406 410 1452 449
rect 1406 376 1412 410
rect 1446 376 1452 410
tri 1220 337 1240 357 sw
rect 1406 337 1452 376
rect 1168 323 1240 337
tri 1240 323 1254 337 sw
rect 1168 271 1174 323
rect 1226 271 1238 323
rect 1290 271 1296 323
rect 1406 303 1412 337
rect 1446 303 1452 337
rect 1406 263 1452 303
rect 1094 197 1100 231
rect 1134 229 1140 231
tri 1140 229 1169 258 sw
tri 1377 229 1406 258 se
rect 1406 229 1412 263
rect 1446 229 1452 263
rect 1134 224 1169 229
tri 1169 224 1174 229 sw
tri 1372 224 1377 229 se
rect 1377 224 1452 229
rect 1134 197 1452 224
rect 1094 189 1452 197
rect 1094 155 1412 189
rect 1446 155 1452 189
rect 1562 597 1608 639
rect 1562 563 1568 597
rect 1602 563 1608 597
rect 1562 521 1608 563
rect 1562 487 1568 521
rect 1602 487 1608 521
rect 1562 445 1608 487
rect 1562 411 1568 445
rect 1602 411 1608 445
rect 1562 369 1608 411
rect 1562 335 1568 369
rect 1602 335 1608 369
rect 1562 292 1608 335
rect 1562 258 1568 292
rect 1602 258 1608 292
rect 1562 215 1608 258
rect 1562 181 1568 215
rect 1602 181 1608 215
rect 1562 169 1608 181
tri 1724 668 1733 677 se
rect 1733 668 1770 677
rect 1094 143 1452 155
tri 984 103 1018 137 sw
tri 1690 103 1724 137 se
rect 1724 103 1770 668
tri 1770 648 1799 677 nw
rect 2251 597 2257 649
rect 2309 597 2321 649
rect 2373 597 2381 649
rect 2516 641 2650 755
rect 2678 795 2724 807
rect 2678 761 2684 795
rect 2718 761 2724 795
rect 2678 727 2724 761
tri 2724 727 2758 761 sw
rect 2850 755 2856 807
rect 2908 755 2920 807
rect 2972 755 2978 807
tri 3117 781 3143 807 ne
rect 3032 761 3084 773
tri 2850 727 2878 755 ne
rect 2878 727 2942 755
tri 2942 727 2970 755 nw
rect 3032 727 3041 761
rect 3075 727 3084 761
rect 2678 675 2684 727
rect 2736 675 2748 727
rect 2800 675 2806 727
tri 2878 721 2884 727 ne
rect 2516 607 2532 641
rect 2566 607 2604 641
rect 2638 607 2650 641
rect 2516 601 2650 607
rect 1908 362 1914 414
rect 1966 362 1978 414
rect 2030 362 2036 414
rect 2181 405 2311 411
rect 2181 371 2193 405
rect 2227 371 2265 405
rect 2299 371 2311 405
rect 2181 365 2311 371
rect 2373 362 2379 414
rect 2431 362 2443 414
rect 2495 362 2503 414
rect 2884 412 2936 727
tri 2936 721 2942 727 nw
rect 3032 721 3084 727
rect 3032 657 3084 669
rect 3032 585 3041 605
rect 3075 585 3084 605
rect 3032 573 3084 585
rect 3143 585 3195 807
tri 3195 786 3224 815 nw
rect 3251 761 3297 773
rect 3251 727 3257 761
rect 3291 727 3297 761
rect 3251 639 3297 727
tri 3297 639 3331 673 sw
rect 3251 619 3429 639
tri 3195 585 3198 588 sw
rect 3251 585 3257 619
rect 3291 585 3429 619
rect 3143 566 3198 585
tri 3143 544 3165 566 ne
rect 3165 544 3198 566
tri 3198 544 3239 585 sw
rect 3251 573 3429 585
tri 3165 522 3187 544 ne
tri 2936 412 2970 446 sw
rect 2884 406 3127 412
rect 2884 372 3009 406
rect 3043 372 3081 406
rect 3115 372 3127 406
rect 2884 366 3127 372
rect 3187 411 3239 544
tri 3335 539 3369 573 ne
tri 3239 411 3273 445 sw
rect 3187 405 3317 411
rect 3187 371 3199 405
rect 3233 371 3271 405
rect 3305 371 3317 405
rect 3187 365 3317 371
rect 1908 243 2036 362
rect 2084 271 2090 323
rect 2142 271 2154 323
tri 2132 245 2158 271 ne
rect 2158 245 2172 271
rect 2206 245 2212 323
rect 1908 191 1914 243
rect 1966 191 1978 243
rect 2030 191 2036 243
tri 2158 237 2166 245 ne
rect 2166 207 2212 245
rect 2166 173 2172 207
rect 2206 173 2212 207
rect 2166 161 2212 173
rect 2322 279 2368 291
rect 2322 245 2328 279
rect 2362 245 2368 279
rect 2322 207 2368 245
rect 2322 173 2328 207
rect 2362 173 2368 207
tri 1770 103 1804 137 sw
tri 2288 103 2322 137 se
rect 2322 103 2368 173
rect 2478 279 2524 291
rect 2478 245 2484 279
rect 2518 275 2524 279
rect 2980 279 3026 291
tri 2524 275 2526 277 sw
rect 2518 271 2526 275
tri 2526 271 2530 275 sw
rect 2518 245 2530 271
tri 2530 245 2556 271 sw
rect 2980 245 2986 279
rect 3020 245 3026 279
rect 2478 243 2556 245
tri 2556 243 2558 245 sw
rect 2478 173 2484 243
rect 2536 191 2548 243
rect 2600 191 2606 243
rect 2980 207 3026 245
rect 2518 173 2536 191
tri 2536 173 2554 191 nw
rect 2980 173 2986 207
rect 3020 173 3026 207
rect 2478 161 2524 173
tri 2524 161 2536 173 nw
rect 2980 161 3026 173
rect 3136 279 3182 291
rect 3136 245 3142 279
rect 3176 245 3182 279
rect 3210 275 3216 327
rect 3268 275 3280 327
tri 3258 271 3262 275 ne
rect 3262 271 3298 275
tri 3262 245 3288 271 ne
rect 3288 245 3298 271
rect 3332 245 3338 327
rect 3136 207 3182 245
tri 3288 241 3292 245 ne
rect 3136 173 3142 207
rect 3176 173 3182 207
tri 2368 103 2402 137 sw
tri 3102 103 3136 137 se
rect 3136 103 3182 173
rect 3292 207 3338 245
rect 3292 173 3298 207
rect 3332 173 3338 207
rect 3292 161 3338 173
tri 3182 103 3216 137 sw
tri 3335 103 3369 137 se
rect 3369 103 3429 573
rect 53 97 3429 103
rect 53 63 65 97
rect 99 63 138 97
rect 172 63 211 97
rect 245 63 284 97
rect 318 63 357 97
rect 391 63 430 97
rect 464 63 503 97
rect 537 63 576 97
rect 610 63 649 97
rect 683 63 722 97
rect 756 63 795 97
rect 829 63 868 97
rect 902 63 940 97
rect 974 63 1012 97
rect 1046 63 1084 97
rect 1118 63 1156 97
rect 1190 63 1228 97
rect 1262 63 1300 97
rect 1334 63 1372 97
rect 1406 63 1444 97
rect 1478 63 1516 97
rect 1550 63 1588 97
rect 1622 63 1660 97
rect 1694 63 1732 97
rect 1766 63 1804 97
rect 1838 63 1876 97
rect 1910 63 1948 97
rect 1982 63 2020 97
rect 2054 63 2092 97
rect 2126 63 2164 97
rect 2198 63 2236 97
rect 2270 63 2308 97
rect 2342 63 2380 97
rect 2414 63 2452 97
rect 2486 63 2524 97
rect 2558 63 2596 97
rect 2630 63 2668 97
rect 2702 63 2740 97
rect 2774 63 2812 97
rect 2846 63 2884 97
rect 2918 63 2956 97
rect 2990 63 3028 97
rect 3062 63 3100 97
rect 3134 63 3172 97
rect 3206 63 3244 97
rect 3278 63 3316 97
rect 3350 63 3429 97
rect 53 45 3429 63
tri 3338 29 3354 45 ne
rect 3354 29 3429 45
<< via1 >>
rect 550 673 602 725
rect 614 715 632 725
rect 632 715 666 725
rect 614 673 666 715
rect 701 432 753 484
rect 701 368 753 420
rect 1014 515 1066 567
rect 1014 451 1066 503
rect 2090 801 2142 807
rect 2090 767 2094 801
rect 2094 767 2128 801
rect 2128 767 2142 801
rect 2090 755 2142 767
rect 2154 801 2206 807
rect 2154 767 2166 801
rect 2166 767 2200 801
rect 2200 767 2206 801
rect 2154 755 2206 767
rect 1256 715 1290 727
rect 1290 715 1308 727
rect 1256 675 1308 715
rect 1353 675 1405 727
rect 1450 675 1502 727
rect 1546 715 1568 727
rect 1568 715 1598 727
rect 1546 675 1598 715
rect 2522 755 2574 807
rect 2586 755 2638 807
rect 1174 271 1226 323
rect 1238 271 1290 323
rect 2257 641 2309 649
rect 2257 607 2263 641
rect 2263 607 2297 641
rect 2297 607 2309 641
rect 2257 597 2309 607
rect 2321 641 2373 649
rect 2321 607 2335 641
rect 2335 607 2369 641
rect 2369 607 2373 641
rect 2321 597 2373 607
rect 2856 755 2908 807
rect 2920 755 2972 807
rect 2684 723 2736 727
rect 2684 689 2718 723
rect 2718 689 2736 723
rect 2684 675 2736 689
rect 2748 675 2800 727
rect 1914 362 1966 414
rect 1978 362 2030 414
rect 2379 405 2431 414
rect 2379 371 2385 405
rect 2385 371 2419 405
rect 2419 371 2431 405
rect 2379 362 2431 371
rect 2443 405 2495 414
rect 2443 371 2457 405
rect 2457 371 2491 405
rect 2491 371 2495 405
rect 2443 362 2495 371
rect 3032 669 3084 721
rect 3032 619 3084 657
rect 3032 605 3041 619
rect 3041 605 3075 619
rect 3075 605 3084 619
rect 2090 271 2142 323
rect 2154 279 2206 323
rect 2154 271 2172 279
rect 2172 271 2206 279
rect 1914 191 1966 243
rect 1978 191 2030 243
rect 2484 207 2536 243
rect 2484 191 2518 207
rect 2518 191 2536 207
rect 2548 191 2600 243
rect 3216 275 3268 327
rect 3280 279 3332 327
rect 3280 275 3298 279
rect 3298 275 3332 279
<< metal2 >>
rect 544 755 2090 807
rect 2142 755 2154 807
rect 2206 755 2522 807
rect 2574 755 2586 807
rect 2638 755 2856 807
rect 2908 755 2920 807
rect 2972 755 2978 807
rect 544 727 678 755
tri 678 727 706 755 nw
rect 544 725 672 727
rect 544 673 550 725
rect 602 673 614 725
rect 666 673 672 725
tri 672 721 678 727 nw
rect 1246 675 1256 727
rect 1308 675 1353 727
rect 1405 675 1450 727
rect 1502 675 1546 727
rect 1598 675 2684 727
rect 2736 675 2748 727
rect 2800 721 3084 727
rect 2800 675 3032 721
tri 2217 673 2219 675 ne
rect 2219 673 2407 675
tri 2219 669 2223 673 ne
rect 2223 669 2407 673
tri 2407 669 2413 675 nw
tri 2998 669 3004 675 ne
rect 3004 669 3032 675
tri 2223 657 2235 669 ne
rect 2235 657 2395 669
tri 2395 657 2407 669 nw
tri 3004 657 3016 669 ne
rect 3016 657 3084 669
tri 2235 649 2243 657 ne
rect 2243 649 2379 657
tri 2243 641 2251 649 ne
rect 2251 597 2257 649
rect 2309 597 2321 649
rect 2373 597 2379 649
tri 2379 641 2395 657 nw
tri 3016 641 3032 657 ne
rect 3032 599 3084 605
rect 1014 567 1066 573
tri 998 515 1014 531 se
tri 986 503 998 515 se
rect 998 503 1066 515
tri 980 497 986 503 se
rect 986 497 1014 503
rect 701 484 753 490
rect 839 451 1014 497
tri 1066 497 1100 531 sw
rect 1066 451 2668 497
rect 701 420 753 432
tri 753 414 787 448 sw
rect 839 445 2668 451
tri 2582 414 2613 445 ne
rect 2613 414 2668 445
rect 753 368 1914 414
rect 701 362 1914 368
rect 1966 362 1978 414
rect 2030 362 2036 414
rect 2373 362 2379 414
rect 2431 362 2443 414
rect 2495 362 2501 414
tri 2613 411 2616 414 ne
tri 2343 327 2373 357 se
rect 2373 327 2501 362
tri 2339 323 2343 327 se
rect 2343 323 2501 327
rect 1168 271 1174 323
rect 1226 271 1238 323
rect 1290 271 2090 323
rect 2142 271 2154 323
rect 2206 271 2501 323
rect 2616 327 2668 414
tri 2668 327 2702 361 sw
rect 2616 275 3216 327
rect 3268 275 3280 327
rect 3332 275 3341 327
rect 1908 191 1914 243
rect 1966 191 1978 243
rect 2030 191 2484 243
rect 2536 191 2548 243
rect 2600 191 2606 243
use DFL1_CDNS_52468879185881  DFL1_CDNS_52468879185881_0
timestamp 1707688321
transform 1 0 2744 0 1 689
box 0 0 1 1
use DFL1_CDNS_52468879185881  DFL1_CDNS_52468879185881_1
timestamp 1707688321
transform 1 0 2096 0 1 689
box 0 0 1 1
use nfet_CDNS_52468879185783  nfet_CDNS_52468879185783_0
timestamp 1707688321
transform 1 0 3086 0 1 573
box -79 -32 239 232
use nfet_CDNS_52468879185871  nfet_CDNS_52468879185871_0
timestamp 1707688321
transform 1 0 2217 0 1 173
box -79 -32 179 182
use nfet_CDNS_52468879185871  nfet_CDNS_52468879185871_1
timestamp 1707688321
transform 1 0 3187 0 1 173
box -79 -32 179 182
use nfet_CDNS_52468879185871  nfet_CDNS_52468879185871_2
timestamp 1707688321
transform 1 0 3031 0 1 173
box -79 -32 179 182
use nfet_CDNS_52468879185871  nfet_CDNS_52468879185871_3
timestamp 1707688321
transform 1 0 2373 0 1 173
box -79 -32 179 182
use nfet_CDNS_52468879185882  nfet_CDNS_52468879185882_0
timestamp 1707688321
transform 1 0 1145 0 1 173
box -82 -32 494 632
use nfet_CDNS_52468879185883  nfet_CDNS_52468879185883_0
timestamp 1707688321
transform -1 0 933 0 1 173
box -82 -32 182 632
use nfet_CDNS_52468879185883  nfet_CDNS_52468879185883_1
timestamp 1707688321
transform -1 0 1089 0 1 173
box -82 -32 182 632
use nfet_CDNS_52468879185884  nfet_CDNS_52468879185884_0
timestamp 1707688321
transform 1 0 365 0 1 173
box -82 -32 494 632
use nfet_CDNS_52468879185885  nfet_CDNS_52468879185885_0
timestamp 1707688321
transform 1 0 2217 0 1 689
box -79 -32 279 116
use nfet_CDNS_52468879185885  nfet_CDNS_52468879185885_1
timestamp 1707688321
transform 1 0 2473 0 1 689
box -79 -32 279 116
<< properties >>
string GDS_END 7597022
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7565376
string path 52.100 19.525 55.300 19.525 
<< end >>
