magic
tech sky130B
timestamp 1707688321
<< properties >>
string GDS_END 30560338
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 30555918
<< end >>
