magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< obsli1 >>
rect 214 200 14555 39939
<< metal1 >>
rect 621 7763 1123 8496
rect 621 7749 1109 7763
rect 621 7735 1095 7749
rect 621 7721 1081 7735
rect 621 7707 1067 7721
rect 621 7693 1053 7707
rect 621 7679 1039 7693
rect 621 7665 1025 7679
rect 621 7651 1011 7665
rect 621 7637 997 7651
rect 621 7623 983 7637
rect 621 7609 969 7623
rect 621 7595 955 7609
rect 621 5831 941 7595
rect 620 4781 2366 5518
rect 620 4767 2352 4781
rect 620 4753 2338 4767
rect 620 4739 2324 4753
rect 620 4725 2310 4739
rect 9537 4792 10263 8496
rect 620 4711 2296 4725
rect 620 4697 2282 4711
rect 620 4683 2268 4697
rect 620 4669 2254 4683
rect 620 4655 2240 4669
rect 620 4641 2226 4655
rect 620 4627 2212 4641
rect 620 4613 2198 4627
rect 620 4599 2184 4613
rect 620 4585 2170 4599
rect 620 4571 2156 4585
rect 620 4557 2142 4571
rect 620 4543 2128 4557
rect 620 4529 2114 4543
rect 620 4515 2100 4529
rect 620 4501 2086 4515
rect 620 4487 2072 4501
rect 620 4473 2058 4487
rect 620 4459 2044 4473
rect 620 4445 2030 4459
rect 620 4431 2016 4445
rect 620 4417 2002 4431
rect 620 4403 1988 4417
rect 620 4389 1974 4403
rect 620 4375 1960 4389
rect 620 4361 1946 4375
rect 620 4347 1932 4361
rect 620 4333 1918 4347
rect 620 4319 1904 4333
rect 620 4305 1890 4319
rect 620 4291 1876 4305
rect 620 4277 1862 4291
rect 620 4263 1848 4277
rect 620 4249 1834 4263
rect 620 4235 1820 4249
rect 620 4221 1806 4235
rect 620 4207 1792 4221
rect 620 4193 1778 4207
rect 620 4179 1764 4193
rect 620 4165 1750 4179
rect 620 4151 1736 4165
rect 620 4137 1722 4151
rect 620 4123 1708 4137
rect 620 4109 1694 4123
rect 620 4095 1680 4109
rect 620 2 1666 4095
<< obsm1 >>
rect 0 8524 15000 40000
rect 0 5803 593 8524
rect 1179 7707 9481 8524
rect 1165 7693 9481 7707
rect 1151 7679 9481 7693
rect 1137 7665 9481 7679
rect 1123 7651 9481 7665
rect 1109 7637 9481 7651
rect 1095 7623 9481 7637
rect 1081 7609 9481 7623
rect 1067 7595 9481 7609
rect 1053 7581 9481 7595
rect 1039 7567 9481 7581
rect 1025 7553 9481 7567
rect 1011 7539 9481 7553
rect 997 5803 9481 7539
rect 0 5546 9481 5803
rect 0 0 592 5546
rect 2422 4736 9481 5546
rect 10319 4736 15000 8524
rect 2422 4725 15000 4736
rect 2408 4711 15000 4725
rect 2394 4697 15000 4711
rect 2380 4683 15000 4697
rect 2366 4669 15000 4683
rect 2352 4655 15000 4669
rect 2338 4641 15000 4655
rect 2324 4627 15000 4641
rect 2310 4613 15000 4627
rect 2296 4599 15000 4613
rect 2282 4585 15000 4599
rect 2268 4571 15000 4585
rect 2254 4557 15000 4571
rect 2240 4543 15000 4557
rect 2226 4529 15000 4543
rect 2212 4515 15000 4529
rect 2198 4501 15000 4515
rect 2184 4487 15000 4501
rect 2170 4473 15000 4487
rect 2156 4459 15000 4473
rect 2142 4445 15000 4459
rect 2128 4431 15000 4445
rect 2114 4417 15000 4431
rect 2100 4403 15000 4417
rect 2086 4389 15000 4403
rect 2072 4375 15000 4389
rect 2058 4361 15000 4375
rect 2044 4347 15000 4361
rect 2030 4333 15000 4347
rect 2016 4319 15000 4333
rect 2002 4305 15000 4319
rect 1988 4291 15000 4305
rect 1974 4277 15000 4291
rect 1960 4263 15000 4277
rect 1946 4249 15000 4263
rect 1932 4235 15000 4249
rect 1918 4221 15000 4235
rect 1904 4207 15000 4221
rect 1890 4193 15000 4207
rect 1876 4179 15000 4193
rect 1862 4165 15000 4179
rect 1848 4151 15000 4165
rect 1834 4137 15000 4151
rect 1820 4123 15000 4137
rect 1806 4109 15000 4123
rect 1792 4095 15000 4109
rect 1778 4081 15000 4095
rect 1764 4067 15000 4081
rect 1750 4053 15000 4067
rect 1736 4039 15000 4053
rect 1722 0 15000 4039
<< metal2 >>
rect 187 8390 2824 39015
rect 187 3698 3041 8390
rect 10934 7223 11383 7933
rect 12222 6182 14858 38003
rect 12213 6168 14858 6182
rect 12199 6154 14858 6168
rect 12185 6140 14858 6154
rect 12171 6126 14858 6140
rect 12157 6112 14858 6126
rect 12143 6098 14858 6112
rect 12129 6084 14858 6098
rect 12115 6070 14858 6084
rect 12101 6056 14858 6070
rect 12087 6042 14858 6056
rect 12073 6028 14858 6042
rect 12059 6014 14858 6028
rect 12045 6000 14858 6014
rect 12031 5986 14858 6000
rect 12017 5972 14858 5986
rect 12003 5958 14858 5972
rect 11989 5944 14858 5958
rect 11975 5930 14858 5944
rect 11961 5916 14858 5930
rect 11947 5902 14858 5916
rect 11933 5888 14858 5902
rect 11919 5874 14858 5888
rect 11905 5860 14858 5874
rect 11891 5846 14858 5860
rect 11877 5832 14858 5846
rect 11863 5818 14858 5832
rect 11849 5804 14858 5818
rect 11835 5790 14858 5804
rect 11821 5776 14858 5790
rect 11807 5762 14858 5776
rect 11793 5748 14858 5762
rect 11779 5734 14858 5748
rect 11765 5720 14858 5734
rect 11751 5706 14858 5720
rect 11737 5692 14858 5706
rect 11723 5678 14858 5692
rect 11709 5664 14858 5678
rect 11695 5650 14858 5664
rect 11681 5636 14858 5650
rect 11667 5622 14858 5636
rect 11653 5608 14858 5622
rect 11639 5594 14858 5608
rect 11625 5580 14858 5594
rect 11611 5566 14858 5580
rect 11597 5552 14858 5566
rect 11583 5538 14858 5552
rect 11569 5524 14858 5538
rect 11555 5510 14858 5524
rect 11541 5496 14858 5510
rect 11527 5482 14858 5496
rect 11513 5468 14858 5482
rect 11499 5454 14858 5468
rect 11485 5440 14858 5454
rect 11471 5426 14858 5440
rect 11457 5412 14858 5426
rect 11443 5398 14858 5412
rect 11429 5384 14858 5398
rect 11415 5370 14858 5384
rect 11401 5356 14858 5370
rect 11387 5342 14858 5356
rect 11373 5328 14858 5342
rect 11359 5314 14858 5328
rect 11345 5300 14858 5314
rect 11331 5286 14858 5300
rect 11317 5272 14858 5286
rect 11303 5258 14858 5272
rect 11289 5244 14858 5258
rect 11275 5230 14858 5244
rect 11261 5216 14858 5230
rect 11247 5202 14858 5216
rect 11233 5188 14858 5202
rect 11219 5174 14858 5188
rect 11205 5160 14858 5174
rect 11191 5146 14858 5160
rect 11177 5132 14858 5146
rect 187 411 4879 3698
rect 99 0 4879 411
rect 5179 0 5579 384
rect 10078 0 14858 5132
<< obsm2 >>
rect 0 39071 15000 40000
rect 0 434 131 39071
rect 2880 38059 15000 39071
rect 2880 8446 12166 38059
rect 3097 7989 12166 8446
rect 3097 7167 10878 7989
rect 11439 7167 12166 7989
rect 3097 6238 12166 7167
rect 3097 6224 12157 6238
rect 3097 6210 12143 6224
rect 3097 6196 12129 6210
rect 3097 6182 12115 6196
rect 3097 6168 12101 6182
rect 3097 6154 12087 6168
rect 3097 6140 12073 6154
rect 3097 6126 12059 6140
rect 3097 6112 12045 6126
rect 3097 6098 12031 6112
rect 3097 6084 12017 6098
rect 3097 6070 12003 6084
rect 3097 6056 11989 6070
rect 3097 6042 11975 6056
rect 3097 6028 11961 6042
rect 3097 6014 11947 6028
rect 3097 6000 11933 6014
rect 3097 5986 11919 6000
rect 3097 5972 11905 5986
rect 3097 5958 11891 5972
rect 3097 5944 11877 5958
rect 3097 5930 11863 5944
rect 3097 5916 11849 5930
rect 3097 5902 11835 5916
rect 3097 5888 11821 5902
rect 3097 5874 11807 5888
rect 3097 5860 11793 5874
rect 3097 5846 11779 5860
rect 3097 5832 11765 5846
rect 3097 5818 11751 5832
rect 3097 5804 11737 5818
rect 3097 5790 11723 5804
rect 3097 5776 11709 5790
rect 3097 5762 11695 5776
rect 3097 5748 11681 5762
rect 3097 5734 11667 5748
rect 3097 5720 11653 5734
rect 3097 5706 11639 5720
rect 3097 5692 11625 5706
rect 3097 5678 11611 5692
rect 3097 5664 11597 5678
rect 3097 5650 11583 5664
rect 3097 5636 11569 5650
rect 3097 5622 11555 5636
rect 3097 5608 11541 5622
rect 3097 5594 11527 5608
rect 3097 5580 11513 5594
rect 3097 5566 11499 5580
rect 3097 5552 11485 5566
rect 3097 5538 11471 5552
rect 3097 5524 11457 5538
rect 3097 5510 11443 5524
rect 3097 5496 11429 5510
rect 3097 5482 11415 5496
rect 3097 5468 11401 5482
rect 3097 5454 11387 5468
rect 3097 5440 11373 5454
rect 3097 5426 11359 5440
rect 3097 5412 11345 5426
rect 3097 5398 11331 5412
rect 3097 5384 11317 5398
rect 3097 5370 11303 5384
rect 3097 5356 11289 5370
rect 3097 5342 11275 5356
rect 3097 5328 11261 5342
rect 3097 5314 11247 5328
rect 3097 5300 11233 5314
rect 3097 5286 11219 5300
rect 3097 5272 11205 5286
rect 3097 5258 11191 5272
rect 3097 5244 11177 5258
rect 3097 5230 11163 5244
rect 3097 5216 11149 5230
rect 3097 5202 11135 5216
rect 3097 5188 11121 5202
rect 3097 3754 10022 5188
rect 0 0 43 434
rect 4935 440 10022 3754
rect 4935 0 5123 440
rect 5635 0 10022 440
rect 14914 0 15000 38059
<< metal3 >>
rect 3100 34528 5002 39015
rect 3100 34516 4990 34528
rect 3100 34486 4960 34516
rect 3100 34456 4930 34486
rect 3100 34426 4900 34456
rect 3100 34396 4870 34426
rect 3100 34366 4840 34396
rect 3100 34336 4810 34366
rect 3100 34306 4780 34336
rect 3100 34276 4750 34306
rect 3100 34246 4720 34276
rect 3100 34216 4690 34246
rect 3100 34186 4660 34216
rect 3100 34156 4630 34186
rect 3100 34126 4600 34156
rect 3100 34096 4570 34126
rect 3100 34066 4540 34096
rect 3100 34036 4510 34066
rect 3100 34006 4480 34036
rect 3100 33976 4450 34006
rect 3100 33946 4420 33976
rect 3100 33916 4390 33946
rect 3100 33886 4360 33916
rect 3100 33856 4330 33886
rect 3100 20440 4300 33856
rect 5186 35070 7364 39015
rect 5186 35052 7346 35070
rect 5186 35022 7316 35052
rect 5186 34992 7286 35022
rect 5186 34962 7256 34992
rect 5186 34932 7226 34962
rect 5186 34902 7196 34932
rect 5186 34872 7166 34902
rect 5186 34842 7136 34872
rect 5186 34812 7106 34842
rect 5186 34782 7076 34812
rect 5186 34752 7046 34782
rect 5186 34722 7016 34752
rect 5186 34692 6986 34722
rect 5186 34662 6956 34692
rect 5186 34632 6926 34662
rect 5186 34602 6896 34632
rect 5186 34572 6866 34602
rect 5186 34542 6836 34572
rect 5186 34512 6806 34542
rect 5186 34482 6776 34512
rect 5186 34452 6746 34482
rect 5186 34422 6716 34452
rect 5186 34392 6686 34422
rect 5186 34362 6656 34392
rect 5186 34332 6626 34362
rect 5186 34302 6596 34332
rect 5186 34272 6566 34302
rect 5186 34242 6536 34272
rect 5186 34212 6506 34242
rect 5186 34182 6476 34212
rect 5186 34152 6446 34182
rect 5186 34122 6416 34152
rect 5186 20478 6386 34122
rect 8571 21630 9771 38004
rect 8077 21611 9752 21630
rect 8058 21581 9722 21611
rect 8028 21551 9692 21581
rect 10657 21592 11857 38008
rect 10161 21581 11846 21592
rect 7998 21521 9662 21551
rect 10150 21551 11816 21581
rect 7968 21491 9632 21521
rect 10120 21521 11786 21551
rect 7938 21461 9602 21491
rect 10090 21491 11756 21521
rect 7908 21431 9572 21461
rect 10060 21461 11726 21491
rect 7878 21401 9542 21431
rect 10030 21431 11696 21461
rect 7848 21371 9512 21401
rect 10000 21401 11666 21431
rect 7818 21341 9482 21371
rect 9970 21371 11636 21401
rect 7788 21311 9452 21341
rect 9940 21341 11606 21371
rect 7758 21281 9422 21311
rect 9910 21311 11576 21341
rect 7728 21251 9392 21281
rect 9880 21281 11546 21311
rect 7698 21221 9362 21251
rect 9850 21251 11516 21281
rect 7668 21191 9332 21221
rect 9820 21221 11486 21251
rect 7638 21161 9302 21191
rect 9790 21191 11456 21221
rect 7608 21131 9272 21161
rect 9760 21161 11426 21191
rect 3129 20411 4796 20440
rect 5205 20459 6880 20478
rect 3159 20381 4825 20411
rect 5235 20429 6899 20459
rect 5265 20399 6929 20429
rect 3189 20351 4855 20381
rect 3219 20321 4885 20351
rect 5295 20369 6959 20399
rect 3249 20291 4915 20321
rect 5325 20339 6989 20369
rect 3279 20261 4945 20291
rect 5355 20309 7019 20339
rect 3309 20231 4975 20261
rect 5385 20279 7049 20309
rect 3339 20201 5005 20231
rect 5415 20249 7079 20279
rect 3369 20171 5035 20201
rect 5445 20219 7109 20249
rect 3399 20141 5065 20171
rect 5475 20189 7139 20219
rect 3429 20111 5095 20141
rect 5505 20159 7169 20189
rect 3459 20081 5125 20111
rect 5535 20129 7199 20159
rect 3489 20051 5155 20081
rect 5565 20099 7229 20129
rect 3519 20021 5185 20051
rect 5595 20069 7259 20099
rect 3549 19991 5215 20021
rect 5625 20039 7289 20069
rect 3579 19961 5245 19991
rect 5655 20009 7319 20039
rect 3609 19931 5275 19961
rect 5685 19979 7349 20009
rect 5699 19965 7379 19979
rect 3639 19901 5305 19931
rect 5729 19935 7379 19965
rect 3669 19871 5335 19901
rect 5759 19905 7379 19935
rect 3699 19841 5365 19871
rect 5789 19875 7379 19905
rect 3729 19811 5395 19841
rect 5819 19845 7379 19875
rect 3759 19781 5425 19811
rect 5849 19815 7379 19845
rect 3789 19751 5455 19781
rect 5879 19785 7379 19815
rect 3819 19721 5485 19751
rect 5909 19755 7379 19785
rect 3849 19691 5515 19721
rect 5939 19725 7379 19755
rect 3879 19661 5545 19691
rect 5969 19695 7379 19725
rect 3909 19631 5575 19661
rect 5999 19665 7379 19695
rect 3939 19601 5605 19631
rect 6029 19635 7379 19665
rect 3969 19571 5635 19601
rect 6059 19605 7379 19635
rect 3999 19541 5665 19571
rect 6089 19575 7379 19605
rect 4029 19511 5695 19541
rect 6119 19545 7379 19575
rect 4059 19481 5725 19511
rect 6149 19515 7379 19545
rect 4089 19451 5755 19481
rect 6179 19485 7379 19515
rect 4119 19421 5785 19451
rect 6209 19455 7379 19485
rect 4149 19391 5815 19421
rect 6239 19425 7379 19455
rect 4179 19361 5845 19391
rect 6269 19395 7379 19425
rect 4209 19331 5875 19361
rect 6299 19365 7379 19395
rect 4239 19301 5905 19331
rect 4269 19271 5905 19301
rect 4299 19241 5905 19271
rect 4329 19211 5905 19241
rect 4359 19181 5905 19211
rect 4389 19151 5905 19181
rect 4419 19121 5905 19151
rect 4449 19091 5905 19121
rect 4479 19061 5905 19091
rect 4509 19031 5905 19061
rect 4539 19001 5905 19031
rect 4569 18971 5905 19001
rect 4599 18941 5905 18971
rect 4629 18911 5905 18941
rect 4659 18881 5905 18911
rect 4689 18851 5905 18881
rect 4719 18821 5905 18851
rect 4749 18508 5905 18821
rect 6329 19335 7379 19365
rect 6359 19305 7379 19335
rect 4764 18493 6017 18508
rect 4779 18478 6032 18493
rect 6389 0 7379 19305
rect 7578 21117 9258 21131
rect 9730 21131 11396 21161
rect 7578 21087 9228 21117
rect 9700 21101 11366 21131
rect 7578 21057 9198 21087
rect 9670 21071 11336 21101
rect 7578 21027 9168 21057
rect 9640 21041 11306 21071
rect 7578 20997 9138 21027
rect 9610 21011 11276 21041
rect 7578 20967 9108 20997
rect 9580 20981 11246 21011
rect 7578 20937 9078 20967
rect 9550 20951 11216 20981
rect 7578 20907 9048 20937
rect 9520 20921 11186 20951
rect 7578 20877 9018 20907
rect 9490 20891 11156 20921
rect 7578 20847 8988 20877
rect 9460 20861 11126 20891
rect 7578 20817 8958 20847
rect 9430 20831 11096 20861
rect 7578 20787 8928 20817
rect 9400 20801 11066 20831
rect 7578 20757 8898 20787
rect 9370 20771 11036 20801
rect 7578 20727 8868 20757
rect 9340 20741 11006 20771
rect 7578 20697 8838 20727
rect 9310 20711 10976 20741
rect 7578 20667 8808 20697
rect 9280 20681 10946 20711
rect 7578 20637 8778 20667
rect 9250 20651 10916 20681
rect 7578 20607 8748 20637
rect 9220 20621 10886 20651
rect 7578 20577 8718 20607
rect 9190 20591 10856 20621
rect 7578 20547 8688 20577
rect 9160 20561 10826 20591
rect 7578 20517 8658 20547
rect 9130 20531 10796 20561
rect 7578 20487 8628 20517
rect 9100 20501 10766 20531
rect 7578 20457 8598 20487
rect 7578 0 8568 20457
rect 9070 20033 10298 20501
rect 9057 20003 10268 20033
rect 9027 19973 10238 20003
rect 8997 19943 10208 19973
rect 8967 19660 10208 19943
<< obsm3 >>
rect 2525 20360 3020 39015
rect 5082 34448 5106 39015
rect 5070 34436 5106 34448
rect 5040 34406 5106 34436
rect 5010 34376 5106 34406
rect 4980 34346 5106 34376
rect 4950 34316 5106 34346
rect 4920 34286 5106 34316
rect 4890 34256 5106 34286
rect 4860 34226 5106 34256
rect 4830 34196 5106 34226
rect 4800 34166 5106 34196
rect 4770 34136 5106 34166
rect 4740 34106 5106 34136
rect 4710 34076 5106 34106
rect 4680 34046 5106 34076
rect 4650 34016 5106 34046
rect 4620 33986 5106 34016
rect 4590 33956 5106 33986
rect 4560 33926 5106 33956
rect 4530 33896 5106 33926
rect 4500 33866 5106 33896
rect 4470 33836 5106 33866
rect 4440 33806 5106 33836
rect 4410 33776 5106 33806
rect 4380 20520 5106 33776
rect 4876 20491 5106 20520
rect 4905 20461 5106 20491
rect 7444 38088 12298 39015
rect 7444 38084 10577 38088
rect 7444 34990 8491 38084
rect 7426 34972 8491 34990
rect 7396 34942 8491 34972
rect 7366 34912 8491 34942
rect 7336 34882 8491 34912
rect 7306 34852 8491 34882
rect 7276 34822 8491 34852
rect 7246 34792 8491 34822
rect 7216 34762 8491 34792
rect 7186 34732 8491 34762
rect 7156 34702 8491 34732
rect 7126 34672 8491 34702
rect 7096 34642 8491 34672
rect 7066 34612 8491 34642
rect 7036 34582 8491 34612
rect 7006 34552 8491 34582
rect 6976 34522 8491 34552
rect 6946 34492 8491 34522
rect 6916 34462 8491 34492
rect 6886 34432 8491 34462
rect 6856 34402 8491 34432
rect 6826 34372 8491 34402
rect 6796 34342 8491 34372
rect 6766 34312 8491 34342
rect 6736 34282 8491 34312
rect 6706 34252 8491 34282
rect 6676 34222 8491 34252
rect 6646 34192 8491 34222
rect 6616 34162 8491 34192
rect 6586 34132 8491 34162
rect 6556 34102 8491 34132
rect 6526 34072 8491 34102
rect 6496 34042 8491 34072
rect 6466 21710 8491 34042
rect 6466 21691 7997 21710
rect 6466 21661 7978 21691
rect 6466 21631 7948 21661
rect 6466 21601 7918 21631
rect 9851 21672 10577 38084
rect 9851 21661 10081 21672
rect 9851 21631 10070 21661
rect 6466 21571 7888 21601
rect 9851 21601 10040 21631
rect 6466 21541 7858 21571
rect 9851 21571 10010 21601
rect 6466 21511 7828 21541
rect 9851 21550 9980 21571
rect 9832 21541 9980 21550
rect 9832 21531 9950 21541
rect 6466 21481 7798 21511
rect 9802 21511 9950 21531
rect 9802 21501 9920 21511
rect 6466 21451 7768 21481
rect 9772 21481 9920 21501
rect 11937 21512 12298 38088
rect 11926 21501 12298 21512
rect 9772 21471 9890 21481
rect 6466 21421 7738 21451
rect 9742 21451 9890 21471
rect 11896 21471 12298 21501
rect 9742 21441 9860 21451
rect 6466 21391 7708 21421
rect 9712 21421 9860 21441
rect 11866 21441 12298 21471
rect 9712 21411 9830 21421
rect 6466 21361 7678 21391
rect 9682 21391 9830 21411
rect 11836 21411 12298 21441
rect 9682 21381 9800 21391
rect 6466 21331 7648 21361
rect 9652 21361 9800 21381
rect 11806 21381 12298 21411
rect 9652 21351 9770 21361
rect 6466 21301 7618 21331
rect 9622 21331 9770 21351
rect 11776 21351 12298 21381
rect 9622 21321 9740 21331
rect 6466 21271 7588 21301
rect 9592 21301 9740 21321
rect 11746 21321 12298 21351
rect 9592 21291 9710 21301
rect 6466 21241 7558 21271
rect 9562 21271 9710 21291
rect 11716 21291 12298 21321
rect 9562 21261 9680 21271
rect 6466 21211 7528 21241
rect 9532 21241 9680 21261
rect 11686 21261 12298 21291
rect 9532 21231 9650 21241
rect 6466 20558 7498 21211
rect 9502 21211 9650 21231
rect 11656 21231 12298 21261
rect 9502 21201 9620 21211
rect 9472 21181 9620 21201
rect 11626 21201 12298 21231
rect 9472 21171 9590 21181
rect 9442 21151 9590 21171
rect 11596 21171 12298 21201
rect 9442 21141 9560 21151
rect 6960 20539 7498 20558
rect 6979 20509 7498 20539
rect 7009 20479 7498 20509
rect 4935 20431 5106 20461
rect 4965 20401 5106 20431
rect 7039 20449 7498 20479
rect 4995 20398 5106 20401
rect 7069 20419 7498 20449
rect 2525 20331 3049 20360
rect 4995 20379 5125 20398
rect 4995 20371 5155 20379
rect 2525 20301 3079 20331
rect 5025 20349 5155 20371
rect 7099 20389 7498 20419
rect 5025 20341 5185 20349
rect 2525 20271 3109 20301
rect 5055 20319 5185 20341
rect 7129 20359 7498 20389
rect 5055 20311 5215 20319
rect 2525 20241 3139 20271
rect 5085 20289 5215 20311
rect 7159 20329 7498 20359
rect 5085 20281 5245 20289
rect 2525 20211 3169 20241
rect 5115 20259 5245 20281
rect 7189 20299 7498 20329
rect 5115 20251 5275 20259
rect 2525 20181 3199 20211
rect 5145 20229 5275 20251
rect 7219 20269 7498 20299
rect 5145 20221 5305 20229
rect 2525 20151 3229 20181
rect 5175 20199 5305 20221
rect 7249 20239 7498 20269
rect 5175 20191 5335 20199
rect 2525 20121 3259 20151
rect 5205 20169 5335 20191
rect 7279 20209 7498 20239
rect 5205 20161 5365 20169
rect 2525 20091 3289 20121
rect 5235 20139 5365 20161
rect 7309 20179 7498 20209
rect 5235 20131 5395 20139
rect 2525 20061 3319 20091
rect 5265 20109 5395 20131
rect 7339 20149 7498 20179
rect 5265 20101 5425 20109
rect 2525 20031 3349 20061
rect 5295 20079 5425 20101
rect 7369 20119 7498 20149
rect 5295 20071 5455 20079
rect 2525 20001 3379 20031
rect 5325 20049 5455 20071
rect 7399 20089 7498 20119
rect 5325 20041 5485 20049
rect 2525 19971 3409 20001
rect 5355 20019 5485 20041
rect 7429 20059 7498 20089
rect 5355 20011 5515 20019
rect 2525 19941 3439 19971
rect 5385 19989 5515 20011
rect 5385 19981 5545 19989
rect 2525 19911 3469 19941
rect 5415 19959 5545 19981
rect 5415 19951 5575 19959
rect 2525 19881 3499 19911
rect 5445 19929 5575 19951
rect 5445 19921 5605 19929
rect 2525 19851 3529 19881
rect 5475 19899 5605 19921
rect 5475 19891 5619 19899
rect 5505 19885 5619 19891
rect 2525 19821 3559 19851
rect 5505 19861 5649 19885
rect 5535 19855 5649 19861
rect 2525 19791 3589 19821
rect 5535 19831 5679 19855
rect 5565 19825 5679 19831
rect 2525 19761 3619 19791
rect 5565 19801 5709 19825
rect 5595 19795 5709 19801
rect 2525 19731 3649 19761
rect 5595 19771 5739 19795
rect 5625 19765 5739 19771
rect 2525 19701 3679 19731
rect 5625 19741 5769 19765
rect 5655 19735 5769 19741
rect 2525 19671 3709 19701
rect 5655 19711 5799 19735
rect 5685 19705 5799 19711
rect 2525 19641 3739 19671
rect 5685 19681 5829 19705
rect 5715 19675 5829 19681
rect 2525 19611 3769 19641
rect 5715 19651 5859 19675
rect 5745 19645 5859 19651
rect 2525 19581 3799 19611
rect 5745 19621 5889 19645
rect 5775 19615 5889 19621
rect 2525 19551 3829 19581
rect 5775 19591 5919 19615
rect 5805 19585 5919 19591
rect 2525 19521 3859 19551
rect 5805 19561 5949 19585
rect 5835 19555 5949 19561
rect 2525 19491 3889 19521
rect 5835 19531 5979 19555
rect 5865 19525 5979 19531
rect 2525 19461 3919 19491
rect 5865 19501 6009 19525
rect 5895 19495 6009 19501
rect 2525 19431 3949 19461
rect 5895 19471 6039 19495
rect 5925 19465 6039 19471
rect 2525 19401 3979 19431
rect 5925 19441 6069 19465
rect 5955 19435 6069 19441
rect 2525 19371 4009 19401
rect 5955 19411 6099 19435
rect 5985 19405 6099 19411
rect 2525 19341 4039 19371
rect 5985 19375 6129 19405
rect 2525 19311 4069 19341
rect 5985 19345 6159 19375
rect 2525 19281 4099 19311
rect 2525 19251 4129 19281
rect 2525 19221 4159 19251
rect 2525 19191 4189 19221
rect 2525 19161 4219 19191
rect 2525 19131 4249 19161
rect 2525 19101 4279 19131
rect 2525 19071 4309 19101
rect 2525 19041 4339 19071
rect 2525 19011 4369 19041
rect 2525 18981 4399 19011
rect 2525 18951 4429 18981
rect 2525 18921 4459 18951
rect 2525 18891 4489 18921
rect 2525 18861 4519 18891
rect 2525 18831 4549 18861
rect 2525 18801 4579 18831
rect 2525 18771 4609 18801
rect 2525 18741 4639 18771
rect 2525 18428 4669 18741
rect 5985 19315 6189 19345
rect 5985 19285 6219 19315
rect 5985 19255 6249 19285
rect 5985 19225 6279 19255
rect 5985 18588 6309 19225
rect 6097 18573 6309 18588
rect 2525 18413 4684 18428
rect 2525 18398 4699 18413
rect 6112 18398 6309 18573
rect 2525 0 6309 18398
rect 7459 0 7498 20059
rect 9412 21121 9560 21141
rect 11566 21141 12298 21171
rect 9412 21111 9530 21121
rect 9382 21091 9530 21111
rect 11536 21111 12298 21141
rect 9382 21081 9500 21091
rect 9352 21061 9500 21081
rect 11506 21081 12298 21111
rect 9352 21051 9470 21061
rect 9338 21037 9470 21051
rect 11476 21051 12298 21081
rect 9308 21031 9470 21037
rect 9308 21007 9440 21031
rect 11446 21021 12298 21051
rect 9278 21001 9440 21007
rect 9278 20977 9410 21001
rect 11416 20991 12298 21021
rect 9248 20971 9410 20977
rect 9248 20947 9380 20971
rect 11386 20961 12298 20991
rect 9218 20941 9380 20947
rect 9218 20917 9350 20941
rect 11356 20931 12298 20961
rect 9188 20911 9350 20917
rect 9188 20887 9320 20911
rect 11326 20901 12298 20931
rect 9158 20881 9320 20887
rect 9158 20857 9290 20881
rect 11296 20871 12298 20901
rect 9128 20851 9290 20857
rect 9128 20827 9260 20851
rect 11266 20841 12298 20871
rect 9098 20821 9260 20827
rect 9098 20797 9230 20821
rect 11236 20811 12298 20841
rect 9068 20791 9230 20797
rect 9068 20767 9200 20791
rect 11206 20781 12298 20811
rect 9038 20761 9200 20767
rect 9038 20737 9170 20761
rect 11176 20751 12298 20781
rect 9008 20731 9170 20737
rect 9008 20707 9140 20731
rect 11146 20721 12298 20751
rect 8978 20701 9140 20707
rect 8978 20677 9110 20701
rect 11116 20691 12298 20721
rect 8948 20671 9110 20677
rect 8948 20647 9080 20671
rect 11086 20661 12298 20691
rect 8918 20641 9080 20647
rect 8918 20617 9050 20641
rect 11056 20631 12298 20661
rect 8888 20611 9050 20617
rect 8888 20587 9020 20611
rect 11026 20601 12298 20631
rect 8858 20581 9020 20587
rect 8858 20557 8990 20581
rect 10996 20571 12298 20601
rect 8828 20527 8990 20557
rect 10966 20541 12298 20571
rect 8798 20497 8990 20527
rect 10936 20511 12298 20541
rect 8768 20467 8990 20497
rect 8738 20437 8990 20467
rect 8708 20407 8990 20437
rect 8678 20377 8990 20407
rect 8648 20113 8990 20377
rect 8648 20083 8977 20113
rect 8648 20053 8947 20083
rect 8648 20023 8917 20053
rect 10906 20481 12298 20511
rect 10876 20451 12298 20481
rect 10846 20421 12298 20451
rect 8648 19580 8887 20023
rect 10378 19953 12298 20421
rect 10348 19923 12298 19953
rect 10318 19893 12298 19923
rect 10288 19580 12298 19893
rect 8648 0 12298 19580
<< labels >>
rlabel metal1 s 9537 4792 10263 8496 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 621 7763 1123 8496 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 621 7749 1109 7763 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 621 7735 1095 7749 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 621 7721 1081 7735 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 621 7707 1067 7721 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 621 7693 1053 7707 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 621 7679 1039 7693 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 621 7665 1025 7679 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 621 7651 1011 7665 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 621 7637 997 7651 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 621 7623 983 7637 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 621 7609 969 7623 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 621 7595 955 7609 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 621 5831 941 7595 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4781 2366 5518 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4767 2352 4781 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4753 2338 4767 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4739 2324 4753 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4725 2310 4739 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4711 2296 4725 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4697 2282 4711 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4683 2268 4697 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4669 2254 4683 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4655 2240 4669 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4641 2226 4655 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4627 2212 4641 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4613 2198 4627 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4599 2184 4613 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4585 2170 4599 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4571 2156 4585 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4557 2142 4571 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4543 2128 4557 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4529 2114 4543 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4515 2100 4529 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4501 2086 4515 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4487 2072 4501 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4473 2058 4487 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4459 2044 4473 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4445 2030 4459 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4431 2016 4445 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4417 2002 4431 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4403 1988 4417 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4389 1974 4403 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4375 1960 4389 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4361 1946 4375 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4347 1932 4361 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4333 1918 4347 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4319 1904 4333 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4305 1890 4319 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4291 1876 4305 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4277 1862 4291 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4263 1848 4277 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4249 1834 4263 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4235 1820 4249 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4221 1806 4235 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4207 1792 4221 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4193 1778 4207 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4179 1764 4193 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4165 1750 4179 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4151 1736 4165 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4137 1722 4151 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4123 1708 4137 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4109 1694 4123 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 4095 1680 4109 6 vssd
port 1 nsew ground bidirectional
rlabel metal1 s 620 2 1666 4095 6 vssd
port 1 nsew ground bidirectional
rlabel metal2 s 5179 0 5579 384 6 ogc_hvc
port 2 nsew power bidirectional
rlabel metal3 s 3100 34528 5002 39015 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34516 4990 34528 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34486 4960 34516 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34456 4930 34486 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34426 4900 34456 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34396 4870 34426 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34366 4840 34396 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34336 4810 34366 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34306 4780 34336 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34276 4750 34306 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34246 4720 34276 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34216 4690 34246 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34186 4660 34216 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34156 4630 34186 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34126 4600 34156 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34096 4570 34126 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34066 4540 34096 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34036 4510 34066 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 34006 4480 34036 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 33976 4450 34006 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 33946 4420 33976 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 33916 4390 33946 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 33886 4360 33916 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 33856 4330 33886 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3100 20440 4300 33856 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 35070 7364 39015 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 35052 7346 35070 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 35022 7316 35052 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34992 7286 35022 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34962 7256 34992 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34932 7226 34962 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34902 7196 34932 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34872 7166 34902 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34842 7136 34872 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34812 7106 34842 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34782 7076 34812 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34752 7046 34782 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34722 7016 34752 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34692 6986 34722 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34662 6956 34692 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34632 6926 34662 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34602 6896 34632 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34572 6866 34602 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34542 6836 34572 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34512 6806 34542 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34482 6776 34512 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34452 6746 34482 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34422 6716 34452 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34392 6686 34422 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34362 6656 34392 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34332 6626 34362 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34302 6596 34332 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34272 6566 34302 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34242 6536 34272 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34212 6506 34242 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34182 6476 34212 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34152 6446 34182 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 34122 6416 34152 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5186 20478 6386 34122 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3129 20411 4796 20440 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3159 20381 4825 20411 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3189 20351 4855 20381 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3219 20321 4885 20351 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3249 20291 4915 20321 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3279 20261 4945 20291 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3309 20231 4975 20261 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3339 20201 5005 20231 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3369 20171 5035 20201 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3399 20141 5065 20171 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3429 20111 5095 20141 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3459 20081 5125 20111 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3489 20051 5155 20081 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3519 20021 5185 20051 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3549 19991 5215 20021 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3579 19961 5245 19991 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3609 19931 5275 19961 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3639 19901 5305 19931 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3669 19871 5335 19901 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3699 19841 5365 19871 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3729 19811 5395 19841 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3759 19781 5425 19811 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3789 19751 5455 19781 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3819 19721 5485 19751 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3849 19691 5515 19721 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3879 19661 5545 19691 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3909 19631 5575 19661 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3939 19601 5605 19631 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3969 19571 5635 19601 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 3999 19541 5665 19571 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4029 19511 5695 19541 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4059 19481 5725 19511 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4089 19451 5755 19481 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4119 19421 5785 19451 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4149 19391 5815 19421 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4179 19361 5845 19391 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4209 19331 5875 19361 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4239 19301 5905 19331 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4269 19271 5905 19301 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4299 19241 5905 19271 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4329 19211 5905 19241 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4359 19181 5905 19211 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4389 19151 5905 19181 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4419 19121 5905 19151 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4449 19091 5905 19121 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4479 19061 5905 19091 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4509 19031 5905 19061 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4539 19001 5905 19031 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4569 18971 5905 19001 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4599 18941 5905 18971 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4629 18911 5905 18941 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4659 18881 5905 18911 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4689 18851 5905 18881 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4719 18821 5905 18851 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4749 18508 5905 18821 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5205 20459 6880 20478 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5235 20429 6899 20459 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5265 20399 6929 20429 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5295 20369 6959 20399 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5325 20339 6989 20369 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5355 20309 7019 20339 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5385 20279 7049 20309 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5415 20249 7079 20279 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5445 20219 7109 20249 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5475 20189 7139 20219 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5505 20159 7169 20189 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5535 20129 7199 20159 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5565 20099 7229 20129 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5595 20069 7259 20099 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5625 20039 7289 20069 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5655 20009 7319 20039 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5685 19979 7349 20009 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5699 19965 7379 19979 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5729 19935 7379 19965 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5759 19905 7379 19935 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5789 19875 7379 19905 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5819 19845 7379 19875 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5849 19815 7379 19845 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5879 19785 7379 19815 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5909 19755 7379 19785 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5939 19725 7379 19755 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5969 19695 7379 19725 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 5999 19665 7379 19695 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 6029 19635 7379 19665 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 6059 19605 7379 19635 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 6089 19575 7379 19605 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 6119 19545 7379 19575 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 6149 19515 7379 19545 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 6179 19485 7379 19515 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 6209 19455 7379 19485 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 6239 19425 7379 19455 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 6269 19395 7379 19425 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 6299 19365 7379 19395 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 6329 19335 7379 19365 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 6359 19305 7379 19335 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 6389 0 7379 19305 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4764 18493 6017 18508 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 4779 18478 6032 18493 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 99 0 4879 411 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 411 4879 3698 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 3698 3041 8390 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 10934 7223 11383 7933 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal2 s 187 8390 2824 39015 6 src_bdy_hvc
port 3 nsew ground bidirectional
rlabel metal3 s 8571 21630 9771 38004 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10657 21592 11857 38008 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8077 21611 9752 21630 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8058 21581 9722 21611 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8028 21551 9692 21581 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7998 21521 9662 21551 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7968 21491 9632 21521 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7938 21461 9602 21491 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7908 21431 9572 21461 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7878 21401 9542 21431 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7848 21371 9512 21401 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7818 21341 9482 21371 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7788 21311 9452 21341 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7758 21281 9422 21311 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7728 21251 9392 21281 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7698 21221 9362 21251 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7668 21191 9332 21221 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7638 21161 9302 21191 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7608 21131 9272 21161 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10161 21581 11846 21592 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10150 21551 11816 21581 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10120 21521 11786 21551 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10090 21491 11756 21521 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10060 21461 11726 21491 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10030 21431 11696 21461 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 10000 21401 11666 21431 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9970 21371 11636 21401 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9940 21341 11606 21371 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9910 21311 11576 21341 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9880 21281 11546 21311 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9850 21251 11516 21281 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9820 21221 11486 21251 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9790 21191 11456 21221 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9760 21161 11426 21191 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9730 21131 11396 21161 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9700 21101 11366 21131 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9670 21071 11336 21101 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9640 21041 11306 21071 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9610 21011 11276 21041 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9580 20981 11246 21011 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9550 20951 11216 20981 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9520 20921 11186 20951 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9490 20891 11156 20921 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9460 20861 11126 20891 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9430 20831 11096 20861 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9400 20801 11066 20831 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9370 20771 11036 20801 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9340 20741 11006 20771 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9310 20711 10976 20741 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9280 20681 10946 20711 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9250 20651 10916 20681 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9220 20621 10886 20651 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9190 20591 10856 20621 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9160 20561 10826 20591 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9130 20531 10796 20561 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9100 20501 10766 20531 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 21117 9258 21131 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 21087 9228 21117 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 21057 9198 21087 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 21027 9168 21057 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20997 9138 21027 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20967 9108 20997 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20937 9078 20967 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20907 9048 20937 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20877 9018 20907 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20847 8988 20877 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20817 8958 20847 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20787 8928 20817 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20757 8898 20787 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20727 8868 20757 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20697 8838 20727 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20667 8808 20697 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20637 8778 20667 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20607 8748 20637 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20577 8718 20607 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20547 8688 20577 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20517 8658 20547 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20487 8628 20517 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 20457 8598 20487 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 7578 0 8568 20457 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8967 19660 10208 19943 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9070 20033 10298 20501 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9057 20003 10268 20033 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 9027 19973 10238 20003 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal3 s 8997 19943 10208 19973 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 10078 0 14858 5132 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11177 5132 14858 5146 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11191 5146 14858 5160 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11205 5160 14858 5174 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11219 5174 14858 5188 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11233 5188 14858 5202 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11247 5202 14858 5216 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11261 5216 14858 5230 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11275 5230 14858 5244 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11289 5244 14858 5258 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11303 5258 14858 5272 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11317 5272 14858 5286 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11331 5286 14858 5300 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11345 5300 14858 5314 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11359 5314 14858 5328 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11373 5328 14858 5342 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11387 5342 14858 5356 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11401 5356 14858 5370 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11415 5370 14858 5384 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11429 5384 14858 5398 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11443 5398 14858 5412 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11457 5412 14858 5426 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11471 5426 14858 5440 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11485 5440 14858 5454 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11499 5454 14858 5468 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11513 5468 14858 5482 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11527 5482 14858 5496 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11541 5496 14858 5510 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11555 5510 14858 5524 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11569 5524 14858 5538 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11583 5538 14858 5552 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11597 5552 14858 5566 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11611 5566 14858 5580 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11625 5580 14858 5594 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11639 5594 14858 5608 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11653 5608 14858 5622 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11667 5622 14858 5636 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11681 5636 14858 5650 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11695 5650 14858 5664 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11709 5664 14858 5678 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11723 5678 14858 5692 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11737 5692 14858 5706 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11751 5706 14858 5720 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11765 5720 14858 5734 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11779 5734 14858 5748 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11793 5748 14858 5762 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11807 5762 14858 5776 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11821 5776 14858 5790 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11835 5790 14858 5804 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11849 5804 14858 5818 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11863 5818 14858 5832 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11877 5832 14858 5846 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11891 5846 14858 5860 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11905 5860 14858 5874 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11919 5874 14858 5888 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11933 5888 14858 5902 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11947 5902 14858 5916 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11961 5916 14858 5930 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11975 5930 14858 5944 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 11989 5944 14858 5958 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12003 5958 14858 5972 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12017 5972 14858 5986 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12031 5986 14858 6000 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12045 6000 14858 6014 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12059 6014 14858 6028 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12073 6028 14858 6042 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12087 6042 14858 6056 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12101 6056 14858 6070 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12115 6070 14858 6084 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12129 6084 14858 6098 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12143 6098 14858 6112 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12157 6112 14858 6126 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12171 6126 14858 6140 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12185 6140 14858 6154 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12199 6154 14858 6168 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12213 6168 14858 6182 6 drn_hvc
port 4 nsew power bidirectional
rlabel metal2 s 12222 6182 14858 38003 6 drn_hvc
port 4 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 40000
string LEFclass BLOCK
string LEFsymmetry R90
string LEFview TRUE
<< end >>
