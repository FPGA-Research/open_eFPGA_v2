magic
tech sky130B
magscale 1 2
timestamp 1707688321
<< nwell >>
rect -36 679 404 1471
<< pwell >>
rect 232 25 334 159
<< psubdiff >>
rect 258 109 308 133
rect 258 75 266 109
rect 300 75 308 109
rect 258 51 308 75
<< nsubdiff >>
rect 258 1339 308 1363
rect 258 1305 266 1339
rect 300 1305 308 1339
rect 258 1281 308 1305
<< psubdiffcont >>
rect 266 75 300 109
<< nsubdiffcont >>
rect 266 1305 300 1339
<< poly >>
rect 114 742 144 1007
rect 48 726 144 742
rect 48 692 64 726
rect 98 692 144 726
rect 48 676 144 692
rect 114 413 144 676
<< polycont >>
rect 64 692 98 726
<< locali >>
rect 0 1397 368 1431
rect 62 1165 96 1397
rect 266 1339 300 1397
rect 266 1289 300 1305
rect 64 726 98 742
rect 64 676 98 692
rect 162 726 196 1231
rect 162 692 213 726
rect 162 186 196 692
rect 62 17 96 186
rect 266 109 300 125
rect 266 17 300 75
rect 0 -17 368 17
use contact_12  contact_12_0
timestamp 1707688321
transform 1 0 48 0 1 676
box 0 0 1 1
use contact_23  contact_23_0
timestamp 1707688321
transform 1 0 258 0 1 1281
box 0 0 1 1
use contact_24  contact_24_0
timestamp 1707688321
transform 1 0 258 0 1 51
box 0 0 1 1
use nmos_m3_w1_680_sli_dli_da_p  nmos_m3_w1_680_sli_dli_da_p_0
timestamp 1707688321
transform 1 0 54 0 1 51
box -26 -26 176 362
use pmos_m3_w1_650_sli_dli_da_p  pmos_m3_w1_650_sli_dli_da_p_0
timestamp 1707688321
transform 1 0 54 0 1 1033
box -59 -54 209 384
<< labels >>
rlabel locali s 196 709 196 709 4 Z
port 2 nsew
rlabel locali s 81 709 81 709 4 A
port 1 nsew
rlabel locali s 184 1414 184 1414 4 vdd
port 3 nsew
rlabel locali s 184 0 184 0 4 gnd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 368 1414
string GDS_END 55114
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 53396
<< end >>
