magic
tech sky130A
magscale 1 2
timestamp 1707688321
<< metal2 >>
rect 0 1185 536 1194
rect 0 0 536 9
<< via2 >>
rect 0 9 536 1185
<< metal3 >>
rect -5 1185 541 1190
rect -5 9 0 1185
rect 536 9 541 1185
rect -5 4 541 9
<< properties >>
string GDS_END 93494200
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 93487348
<< end >>
